magic
tech scmos
timestamp 1732943601
<< metal1 >>
rect 880 2103 882 2107
rect 886 2103 889 2107
rect 893 2103 896 2107
rect 1912 2103 1914 2107
rect 1918 2103 1921 2107
rect 1925 2103 1928 2107
rect 614 2068 625 2071
rect 1294 2068 1297 2078
rect 1726 2068 1734 2071
rect 2294 2068 2302 2071
rect 262 2058 281 2061
rect 614 2061 617 2068
rect 574 2058 593 2061
rect 598 2058 617 2061
rect 854 2058 873 2061
rect 886 2058 902 2061
rect 1134 2058 1153 2061
rect 1190 2058 1198 2061
rect 1358 2058 1378 2061
rect 1542 2058 1561 2061
rect 1726 2058 1745 2061
rect 1906 2058 1913 2061
rect 1986 2058 1993 2061
rect 2054 2058 2073 2061
rect 2154 2058 2169 2061
rect 278 2048 281 2058
rect 574 2048 577 2058
rect 870 2048 873 2058
rect 1134 2048 1137 2058
rect 1542 2048 1545 2058
rect 1726 2048 1729 2058
rect 1830 2052 1834 2057
rect 2054 2048 2057 2058
rect 1083 2038 1086 2042
rect 1218 2038 1219 2042
rect 1491 2038 1494 2042
rect 376 2003 378 2007
rect 382 2003 385 2007
rect 389 2003 392 2007
rect 1392 2003 1394 2007
rect 1398 2003 1401 2007
rect 1405 2003 1408 2007
rect 181 1988 182 1992
rect 754 1988 755 1992
rect 1770 1988 1771 1992
rect 149 1968 150 1972
rect 213 1968 214 1972
rect 475 1968 478 1972
rect 882 1968 883 1972
rect 1058 1968 1059 1972
rect 1282 1968 1283 1972
rect 1930 1968 1937 1971
rect 2082 1968 2089 1971
rect 106 1948 113 1951
rect 214 1948 230 1951
rect 262 1951 265 1961
rect 234 1948 241 1951
rect 246 1948 265 1951
rect 438 1948 454 1951
rect 766 1951 769 1961
rect 894 1958 910 1961
rect 766 1948 785 1951
rect 1206 1948 1214 1951
rect 1294 1951 1297 1961
rect 1294 1948 1313 1951
rect 1366 1951 1369 1961
rect 1378 1958 1382 1962
rect 1322 1948 1345 1951
rect 1350 1948 1369 1951
rect 1630 1951 1633 1961
rect 1630 1948 1649 1951
rect 1714 1948 1721 1951
rect 1782 1951 1785 1961
rect 1782 1948 1801 1951
rect 1886 1951 1889 1961
rect 1886 1948 1905 1951
rect 2054 1951 2057 1961
rect 2054 1948 2073 1951
rect 2258 1948 2273 1951
rect 222 1938 230 1941
rect 834 1938 841 1941
rect 1330 1938 1337 1941
rect 1654 1938 1666 1941
rect 1886 1938 1894 1941
rect 1910 1938 1926 1941
rect 1662 1936 1666 1938
rect 557 1918 558 1922
rect 1837 1918 1838 1922
rect 880 1903 882 1907
rect 886 1903 889 1907
rect 893 1903 896 1907
rect 1912 1903 1914 1907
rect 1918 1903 1921 1907
rect 1925 1903 1928 1907
rect 2050 1878 2051 1882
rect 1686 1872 1690 1877
rect 318 1868 326 1871
rect 710 1868 718 1871
rect 730 1868 737 1871
rect 894 1868 902 1871
rect 982 1868 990 1871
rect 1038 1868 1057 1871
rect 2194 1868 2201 1871
rect 38 1858 46 1861
rect 130 1858 145 1861
rect 286 1858 305 1861
rect 310 1858 334 1861
rect 454 1858 470 1861
rect 542 1858 561 1861
rect 690 1858 697 1861
rect 886 1858 894 1861
rect 1038 1861 1041 1868
rect 1030 1858 1041 1861
rect 1050 1858 1057 1861
rect 1122 1858 1129 1861
rect 1174 1858 1193 1861
rect 1274 1858 1281 1861
rect 1382 1858 1390 1861
rect 1454 1858 1470 1861
rect 1606 1858 1625 1861
rect 1702 1858 1710 1861
rect 1774 1858 1793 1861
rect 1854 1858 1862 1861
rect 2062 1858 2070 1861
rect 2182 1858 2201 1861
rect 2238 1858 2257 1861
rect 286 1848 289 1858
rect 542 1848 545 1858
rect 1190 1848 1193 1858
rect 1622 1848 1625 1858
rect 1790 1848 1793 1858
rect 2198 1848 2201 1858
rect 2254 1848 2257 1858
rect 885 1838 886 1842
rect 338 1818 339 1822
rect 397 1818 398 1822
rect 1418 1818 1419 1822
rect 1954 1818 1955 1822
rect 2002 1818 2003 1822
rect 376 1803 378 1807
rect 382 1803 385 1807
rect 389 1803 392 1807
rect 1392 1803 1394 1807
rect 1398 1803 1401 1807
rect 1405 1803 1408 1807
rect 1906 1788 1907 1792
rect 1707 1768 1710 1772
rect 278 1748 286 1751
rect 346 1748 353 1751
rect 470 1748 478 1751
rect 558 1751 561 1761
rect 558 1748 577 1751
rect 738 1748 745 1751
rect 806 1748 822 1751
rect 894 1751 897 1761
rect 894 1748 929 1751
rect 1070 1751 1073 1761
rect 1146 1758 1150 1762
rect 1406 1758 1414 1761
rect 1054 1748 1073 1751
rect 1254 1751 1258 1753
rect 982 1738 990 1741
rect 1006 1741 1009 1748
rect 1254 1748 1273 1751
rect 1338 1748 1345 1751
rect 1398 1748 1422 1751
rect 1482 1748 1489 1751
rect 1550 1751 1553 1761
rect 1550 1748 1569 1751
rect 1606 1751 1609 1761
rect 1958 1758 1977 1761
rect 1606 1748 1625 1751
rect 998 1738 1009 1741
rect 1382 1738 1385 1748
rect 1918 1748 1942 1751
rect 2050 1748 2065 1751
rect 2278 1751 2281 1761
rect 2262 1748 2281 1751
rect 1606 1738 1614 1741
rect 1810 1738 1817 1741
rect 2118 1738 2126 1741
rect 413 1718 414 1722
rect 1826 1718 1827 1722
rect 1850 1718 1851 1722
rect 2146 1718 2147 1722
rect 880 1703 882 1707
rect 886 1703 889 1707
rect 893 1703 896 1707
rect 1912 1703 1914 1707
rect 1918 1703 1921 1707
rect 1925 1703 1928 1707
rect 682 1678 683 1682
rect 2034 1678 2035 1682
rect 2078 1672 2082 1677
rect 190 1668 198 1671
rect 886 1668 910 1671
rect 1190 1668 1209 1671
rect 1466 1668 1467 1672
rect 1698 1668 1705 1671
rect 126 1658 145 1661
rect 258 1658 265 1661
rect 310 1658 329 1661
rect 342 1658 366 1661
rect 406 1658 422 1661
rect 462 1658 478 1661
rect 542 1658 561 1661
rect 578 1658 585 1661
rect 706 1658 721 1661
rect 726 1658 745 1661
rect 898 1658 929 1661
rect 1026 1658 1033 1661
rect 1206 1661 1209 1668
rect 1206 1658 1217 1661
rect 1306 1658 1313 1661
rect 1562 1658 1569 1661
rect 1686 1658 1705 1661
rect 1786 1658 1793 1661
rect 2046 1658 2066 1661
rect 2166 1658 2185 1661
rect 142 1648 145 1658
rect 326 1648 329 1658
rect 462 1657 466 1658
rect 542 1648 545 1658
rect 742 1648 745 1658
rect 1702 1648 1705 1658
rect 2062 1657 2066 1658
rect 2182 1648 2185 1658
rect 294 1638 302 1641
rect 1670 1638 1678 1641
rect 493 1618 494 1622
rect 1010 1618 1011 1622
rect 1229 1618 1230 1622
rect 1277 1618 1278 1622
rect 1373 1618 1374 1622
rect 376 1603 378 1607
rect 382 1603 385 1607
rect 389 1603 392 1607
rect 1392 1603 1394 1607
rect 1398 1603 1401 1607
rect 1405 1603 1408 1607
rect 21 1588 22 1592
rect 2018 1588 2019 1592
rect 442 1568 443 1572
rect 611 1568 614 1572
rect 955 1568 958 1572
rect 990 1568 998 1571
rect 1379 1568 1382 1572
rect 1586 1568 1593 1571
rect 1858 1568 1865 1571
rect 22 1548 38 1551
rect 350 1548 358 1551
rect 454 1551 457 1561
rect 650 1558 654 1562
rect 454 1548 473 1551
rect 498 1548 505 1551
rect 574 1548 582 1551
rect 662 1551 665 1561
rect 1454 1561 1457 1568
rect 1990 1566 1994 1568
rect 1446 1558 1457 1561
rect 1714 1558 1718 1562
rect 662 1548 681 1551
rect 774 1548 790 1551
rect 918 1548 926 1551
rect 1342 1548 1358 1551
rect 78 1538 86 1541
rect 710 1541 713 1548
rect 690 1538 697 1541
rect 710 1538 721 1541
rect 982 1541 985 1548
rect 1766 1548 1782 1551
rect 1830 1551 1833 1561
rect 1830 1548 1849 1551
rect 1906 1548 1921 1551
rect 2102 1551 2105 1561
rect 2102 1548 2121 1551
rect 2138 1548 2145 1551
rect 982 1538 993 1541
rect 1486 1538 1505 1541
rect 1578 1538 1585 1541
rect 1802 1538 1809 1541
rect 1854 1538 1866 1541
rect 2050 1538 2057 1541
rect 2290 1538 2302 1541
rect 42 1528 46 1532
rect 694 1528 697 1538
rect 1862 1536 1866 1538
rect 1410 1528 1425 1531
rect 1045 1518 1046 1522
rect 1754 1518 1755 1522
rect 1986 1518 1987 1522
rect 880 1503 882 1507
rect 886 1503 889 1507
rect 893 1503 896 1507
rect 1912 1503 1914 1507
rect 1918 1503 1921 1507
rect 1925 1503 1928 1507
rect 902 1488 910 1491
rect 1004 1488 1006 1492
rect 1060 1488 1062 1492
rect 1318 1472 1321 1481
rect 1366 1478 1374 1482
rect 2266 1478 2282 1481
rect 1366 1472 1369 1478
rect 2278 1474 2282 1478
rect 154 1468 161 1471
rect 262 1468 273 1471
rect 358 1468 366 1471
rect 126 1458 145 1461
rect 166 1458 174 1461
rect 246 1458 257 1461
rect 454 1461 457 1471
rect 706 1468 713 1471
rect 1074 1468 1081 1471
rect 1382 1468 1390 1471
rect 1685 1468 1686 1472
rect 1930 1468 1953 1471
rect 2074 1468 2082 1471
rect 450 1458 457 1461
rect 510 1458 518 1461
rect 582 1458 590 1461
rect 670 1458 689 1461
rect 698 1458 721 1461
rect 774 1458 782 1461
rect 798 1458 806 1461
rect 1118 1458 1126 1461
rect 1146 1458 1153 1461
rect 1206 1458 1225 1461
rect 1302 1458 1318 1461
rect 1350 1458 1358 1461
rect 1430 1458 1449 1461
rect 1458 1458 1465 1461
rect 1554 1458 1561 1461
rect 1766 1458 1785 1461
rect 1842 1458 1857 1461
rect 1910 1458 1934 1461
rect 2190 1458 2198 1461
rect 126 1448 129 1458
rect 254 1452 257 1458
rect 670 1448 673 1458
rect 918 1448 926 1451
rect 982 1448 990 1451
rect 1038 1448 1046 1451
rect 1206 1448 1209 1458
rect 1278 1451 1281 1458
rect 1270 1448 1281 1451
rect 1430 1448 1433 1458
rect 1766 1448 1769 1458
rect 1918 1448 1926 1451
rect 293 1438 294 1442
rect 902 1438 918 1441
rect 1534 1438 1542 1441
rect 1794 1438 1801 1441
rect 402 1418 403 1422
rect 722 1418 723 1422
rect 1621 1418 1622 1422
rect 376 1403 378 1407
rect 382 1403 385 1407
rect 389 1403 392 1407
rect 1392 1403 1394 1407
rect 1398 1403 1401 1407
rect 1405 1403 1408 1407
rect 1829 1388 1830 1392
rect 94 1368 102 1371
rect 1058 1368 1073 1371
rect 1846 1366 1850 1368
rect 126 1351 129 1361
rect 110 1348 129 1351
rect 190 1348 206 1351
rect 318 1348 326 1351
rect 402 1348 409 1351
rect 422 1351 425 1361
rect 618 1358 625 1361
rect 1142 1358 1150 1361
rect 1182 1358 1190 1361
rect 1426 1358 1430 1362
rect 1478 1358 1486 1361
rect 1714 1358 1718 1362
rect 422 1348 441 1351
rect 670 1348 678 1351
rect 738 1348 745 1351
rect 122 1338 129 1341
rect 214 1332 217 1342
rect 338 1338 339 1342
rect 486 1341 489 1348
rect 966 1348 977 1351
rect 1278 1348 1289 1351
rect 1574 1348 1582 1351
rect 1686 1348 1702 1351
rect 1758 1351 1761 1361
rect 1814 1351 1817 1361
rect 1758 1348 1777 1351
rect 1798 1348 1817 1351
rect 1930 1348 1945 1351
rect 2054 1351 2057 1361
rect 2066 1358 2070 1362
rect 2038 1348 2057 1351
rect 2270 1351 2274 1353
rect 2270 1348 2281 1351
rect 966 1342 969 1348
rect 1278 1342 1281 1348
rect 486 1338 497 1341
rect 798 1338 812 1341
rect 1090 1338 1097 1341
rect 1526 1338 1534 1341
rect 1630 1341 1633 1348
rect 1622 1338 1633 1341
rect 1660 1338 1662 1342
rect 2022 1338 2030 1341
rect 2174 1338 2186 1341
rect 2294 1338 2302 1341
rect 798 1332 801 1338
rect 1550 1328 1561 1331
rect 2022 1328 2025 1338
rect 1044 1318 1046 1322
rect 1076 1318 1078 1322
rect 1122 1318 1124 1322
rect 1162 1318 1169 1321
rect 1254 1318 1262 1321
rect 1853 1318 1854 1322
rect 880 1303 882 1307
rect 886 1303 889 1307
rect 893 1303 896 1307
rect 1912 1303 1914 1307
rect 1918 1303 1921 1307
rect 1925 1303 1928 1307
rect 414 1288 422 1291
rect 946 1288 953 1291
rect 1142 1288 1150 1291
rect 1418 1288 1425 1291
rect 1698 1288 1699 1292
rect 566 1271 569 1278
rect 742 1277 746 1278
rect 1166 1272 1169 1281
rect 1518 1272 1521 1281
rect 2046 1278 2057 1281
rect 2106 1278 2107 1282
rect 558 1268 569 1271
rect 574 1268 585 1271
rect 1174 1268 1182 1271
rect 1470 1268 1481 1271
rect 1502 1268 1513 1271
rect 1918 1268 1934 1271
rect 1958 1268 1969 1271
rect 2126 1268 2134 1271
rect 182 1258 190 1261
rect 286 1258 305 1261
rect 458 1258 465 1261
rect 534 1258 553 1261
rect 606 1258 625 1261
rect 686 1258 694 1261
rect 706 1258 713 1261
rect 806 1258 825 1261
rect 1470 1262 1473 1268
rect 1286 1258 1294 1261
rect 1390 1258 1422 1261
rect 1734 1258 1742 1261
rect 1766 1258 1785 1261
rect 1842 1258 1857 1261
rect 1966 1261 1969 1268
rect 1966 1258 1977 1261
rect 2126 1261 2129 1268
rect 2118 1258 2129 1261
rect 2142 1258 2161 1261
rect 2174 1258 2182 1261
rect 18 1248 22 1252
rect 286 1248 289 1258
rect 534 1248 537 1258
rect 606 1248 609 1258
rect 806 1248 809 1258
rect 1142 1248 1153 1251
rect 1418 1248 1425 1251
rect 1766 1248 1769 1258
rect 2158 1248 2161 1258
rect 1142 1246 1146 1248
rect 614 1242 618 1244
rect 1150 1242 1153 1248
rect 754 1238 761 1241
rect 2210 1238 2213 1242
rect 594 1218 595 1222
rect 376 1203 378 1207
rect 382 1203 385 1207
rect 389 1203 392 1207
rect 1392 1203 1394 1207
rect 1398 1203 1401 1207
rect 1405 1203 1408 1207
rect 698 1188 699 1192
rect 410 1168 411 1172
rect 1030 1168 1041 1171
rect 1022 1166 1026 1168
rect 1038 1162 1041 1168
rect 166 1151 169 1161
rect 166 1148 185 1151
rect 342 1148 350 1151
rect 494 1151 497 1161
rect 478 1148 497 1151
rect 578 1148 585 1151
rect 710 1151 713 1161
rect 710 1148 729 1151
rect 862 1148 870 1151
rect 966 1151 969 1161
rect 950 1148 969 1151
rect 1042 1148 1049 1151
rect 1070 1151 1073 1161
rect 1222 1158 1230 1161
rect 1070 1148 1089 1151
rect 1446 1151 1449 1161
rect 1746 1158 1750 1162
rect 1810 1158 1814 1162
rect 294 1138 305 1141
rect 930 1138 945 1141
rect 1046 1138 1049 1148
rect 1430 1148 1449 1151
rect 1486 1148 1505 1151
rect 1726 1148 1734 1151
rect 1750 1148 1769 1151
rect 1790 1148 1798 1151
rect 1878 1148 1886 1151
rect 1902 1148 1926 1151
rect 1206 1138 1217 1141
rect 1526 1138 1534 1141
rect 1910 1138 1918 1141
rect 2034 1138 2041 1141
rect 1198 1128 1201 1138
rect 1214 1132 1217 1138
rect 1878 1128 1889 1131
rect 1174 1118 1182 1121
rect 1261 1118 1262 1122
rect 1541 1118 1542 1122
rect 2090 1118 2091 1122
rect 880 1103 882 1107
rect 886 1103 889 1107
rect 893 1103 896 1107
rect 1912 1103 1914 1107
rect 1918 1103 1921 1107
rect 1925 1103 1928 1107
rect 13 1088 14 1092
rect 1850 1088 1851 1092
rect 422 1074 426 1078
rect 22 1068 33 1071
rect 758 1068 769 1071
rect 882 1068 890 1071
rect 942 1068 945 1078
rect 1230 1068 1238 1071
rect 1446 1071 1449 1081
rect 1538 1078 1550 1081
rect 1442 1068 1449 1071
rect 1518 1068 1529 1071
rect 1610 1068 1617 1071
rect 30 1062 33 1068
rect 38 1058 49 1061
rect 54 1058 73 1061
rect 86 1058 94 1061
rect 134 1058 150 1061
rect 222 1058 241 1061
rect 318 1061 321 1068
rect 310 1058 321 1061
rect 510 1058 526 1061
rect 598 1058 617 1061
rect 766 1061 769 1068
rect 1782 1062 1785 1071
rect 1934 1071 1938 1074
rect 1910 1068 1938 1071
rect 2190 1068 2202 1071
rect 766 1058 782 1061
rect 822 1058 841 1061
rect 1006 1058 1025 1061
rect 1378 1058 1385 1061
rect 1406 1058 1433 1061
rect 1454 1058 1462 1061
rect 1490 1058 1505 1061
rect 1558 1058 1566 1061
rect 1602 1058 1609 1061
rect 1630 1058 1638 1061
rect 1790 1058 1809 1061
rect 1886 1058 1905 1061
rect 1978 1058 1993 1061
rect 2086 1058 2094 1061
rect 2154 1058 2161 1061
rect 46 1052 49 1058
rect 70 1048 73 1058
rect 82 1048 86 1052
rect 222 1048 225 1058
rect 614 1048 617 1058
rect 838 1048 841 1058
rect 994 1048 998 1052
rect 1006 1048 1009 1058
rect 1258 1048 1262 1052
rect 1406 1051 1409 1058
rect 1398 1048 1409 1051
rect 1474 1048 1478 1052
rect 1586 1048 1590 1052
rect 1806 1048 1809 1058
rect 1886 1048 1889 1058
rect 582 1038 590 1041
rect 1682 1038 1689 1041
rect 266 1018 267 1022
rect 326 1018 334 1021
rect 1653 1018 1654 1022
rect 1922 1018 1937 1021
rect 376 1003 378 1007
rect 382 1003 385 1007
rect 389 1003 392 1007
rect 1392 1003 1394 1007
rect 1398 1003 1401 1007
rect 1405 1003 1408 1007
rect 1525 988 1526 992
rect 330 968 337 971
rect 494 968 502 971
rect 534 968 545 971
rect 651 968 654 972
rect 670 968 678 971
rect 1810 968 1811 972
rect 1902 968 1918 971
rect 2219 968 2222 972
rect 2286 968 2294 971
rect 526 966 530 968
rect 542 962 545 968
rect 1902 966 1906 968
rect 126 951 129 961
rect 110 948 129 951
rect 182 951 185 961
rect 449 958 454 962
rect 182 948 201 951
rect 702 951 705 961
rect 1318 958 1337 961
rect 686 948 705 951
rect 782 948 790 951
rect 1098 948 1105 951
rect 1190 948 1198 951
rect 1250 948 1257 951
rect 1330 948 1345 951
rect 1350 948 1358 951
rect 1414 948 1422 951
rect 1482 948 1489 951
rect 1570 948 1577 951
rect 45 938 46 942
rect 182 938 190 941
rect 414 941 417 948
rect 1734 948 1742 951
rect 1822 951 1825 961
rect 1802 948 1809 951
rect 1822 948 1841 951
rect 1922 948 1929 951
rect 1950 948 1958 951
rect 1974 948 1982 951
rect 2014 948 2022 951
rect 358 938 385 941
rect 406 938 417 941
rect 422 938 433 941
rect 494 938 505 941
rect 698 938 705 941
rect 898 938 913 941
rect 1062 938 1070 941
rect 1246 938 1254 941
rect 1534 938 1542 941
rect 1990 941 1993 948
rect 2238 951 2242 953
rect 2238 948 2249 951
rect 1922 938 1937 941
rect 1982 938 1993 941
rect 654 932 658 936
rect 1950 928 1961 931
rect 2014 928 2025 931
rect 1149 918 1150 922
rect 1237 918 1238 922
rect 1898 918 1899 922
rect 880 903 882 907
rect 886 903 889 907
rect 893 903 896 907
rect 1912 903 1914 907
rect 1918 903 1921 907
rect 1925 903 1928 907
rect 1485 888 1486 892
rect 2290 888 2291 892
rect 418 878 425 882
rect 422 872 425 878
rect 158 868 166 871
rect 226 868 233 871
rect 582 871 585 881
rect 1550 872 1553 881
rect 1838 878 1846 882
rect 1838 872 1841 878
rect 578 868 585 871
rect 38 858 46 861
rect 106 858 113 861
rect 118 858 126 861
rect 150 858 174 861
rect 182 858 201 861
rect 246 858 254 861
rect 678 862 681 871
rect 550 858 569 861
rect 638 858 646 861
rect 982 862 985 871
rect 1146 868 1153 871
rect 1410 868 1425 871
rect 1442 868 1449 871
rect 1950 868 1958 871
rect 1982 871 1986 874
rect 2142 872 2146 877
rect 1978 868 1986 871
rect 1102 858 1121 861
rect 1142 858 1161 861
rect 1266 858 1273 861
rect 1430 858 1449 861
rect 1582 858 1593 861
rect 1758 858 1766 861
rect 1906 858 1926 861
rect 1950 858 1969 861
rect 2110 858 2130 861
rect 2230 858 2249 861
rect 198 848 201 858
rect 274 848 278 852
rect 550 848 553 858
rect 914 848 918 852
rect 1446 848 1449 858
rect 1498 848 1505 851
rect 1686 848 1689 858
rect 1754 848 1758 852
rect 1950 848 1953 858
rect 2126 857 2130 858
rect 2246 848 2249 858
rect 938 838 945 841
rect 2146 838 2149 842
rect 213 818 214 822
rect 621 818 622 822
rect 1885 818 1886 822
rect 2098 818 2099 822
rect 376 803 378 807
rect 382 803 385 807
rect 389 803 392 807
rect 1392 803 1394 807
rect 1398 803 1401 807
rect 1405 803 1408 807
rect 450 788 451 792
rect 1114 788 1115 792
rect 1874 788 1875 792
rect 1933 788 1934 792
rect 114 768 115 772
rect 38 748 46 751
rect 126 751 129 761
rect 126 748 145 751
rect 182 751 185 761
rect 182 748 201 751
rect 550 748 558 751
rect 566 751 569 761
rect 574 758 582 761
rect 562 748 569 751
rect 678 751 681 761
rect 678 748 697 751
rect 754 748 769 751
rect 810 748 817 751
rect 822 748 830 751
rect 854 751 857 761
rect 854 748 873 751
rect 1198 751 1201 758
rect 1190 748 1201 751
rect 1286 748 1302 751
rect 1354 748 1361 751
rect 1374 751 1377 761
rect 1374 748 1393 751
rect 1446 751 1449 761
rect 1830 758 1841 761
rect 1446 748 1465 751
rect 58 738 59 742
rect 342 738 353 741
rect 394 738 401 741
rect 518 738 526 741
rect 614 738 617 748
rect 1702 751 1706 753
rect 1830 752 1833 758
rect 1702 748 1713 751
rect 1970 748 1977 751
rect 2182 751 2185 761
rect 2166 748 2185 751
rect 702 738 714 741
rect 854 738 862 741
rect 878 738 894 741
rect 1030 738 1038 741
rect 1082 738 1089 741
rect 1226 738 1233 741
rect 1942 738 1953 741
rect 2018 738 2025 741
rect 2178 738 2185 741
rect 710 736 714 738
rect 918 732 922 736
rect 374 718 382 721
rect 898 718 905 721
rect 880 703 882 707
rect 886 703 889 707
rect 893 703 896 707
rect 1912 703 1914 707
rect 1918 703 1921 707
rect 1925 703 1928 707
rect 870 688 878 691
rect 949 688 950 692
rect 1130 688 1131 692
rect 1874 688 1875 692
rect 174 672 177 681
rect 1702 678 1713 681
rect 2274 678 2290 681
rect 2286 674 2290 678
rect 182 668 193 671
rect 214 662 217 671
rect 342 668 353 671
rect 638 668 649 671
rect 1026 668 1033 671
rect 350 662 353 668
rect 78 658 86 661
rect 146 658 153 661
rect 274 658 281 661
rect 646 662 649 668
rect 750 658 769 661
rect 1286 662 1289 671
rect 1394 668 1417 671
rect 2206 668 2218 671
rect 882 658 905 661
rect 994 658 1001 661
rect 1022 658 1030 661
rect 1150 658 1169 661
rect 1214 658 1233 661
rect 1254 658 1273 661
rect 1346 658 1353 661
rect 1574 658 1585 661
rect 2090 658 2097 661
rect 478 648 486 651
rect 750 648 753 658
rect 962 648 969 651
rect 978 648 982 652
rect 1134 648 1142 651
rect 1166 648 1169 658
rect 2054 648 2073 651
rect 502 642 506 644
rect 670 642 674 644
rect 1314 638 1317 642
rect 1430 638 1457 641
rect 2138 638 2141 642
rect 917 618 918 622
rect 1522 618 1523 622
rect 376 603 378 607
rect 382 603 385 607
rect 389 603 392 607
rect 1392 603 1394 607
rect 1398 603 1401 607
rect 1405 603 1408 607
rect 322 588 323 592
rect 538 588 539 592
rect 845 588 846 592
rect 1109 588 1110 592
rect 1477 588 1478 592
rect 1866 588 1867 592
rect 170 568 171 572
rect 570 568 571 572
rect 1062 568 1070 571
rect 1326 568 1337 571
rect 1653 568 1654 572
rect 1326 562 1329 568
rect 182 551 185 561
rect 334 558 342 561
rect 182 548 201 551
rect 390 548 398 551
rect 458 548 465 551
rect 478 551 481 561
rect 1050 558 1057 561
rect 1246 558 1254 561
rect 478 548 497 551
rect 518 548 526 551
rect 30 541 33 548
rect 22 538 33 541
rect 206 538 209 548
rect 862 548 886 551
rect 1150 548 1158 551
rect 1190 548 1198 551
rect 1638 551 1641 561
rect 1622 548 1641 551
rect 814 541 817 548
rect 746 538 753 541
rect 806 538 817 541
rect 1150 541 1153 548
rect 1878 548 1894 551
rect 1934 551 1937 561
rect 1902 548 1937 551
rect 2094 548 2110 551
rect 2158 548 2166 551
rect 2226 548 2233 551
rect 1142 538 1153 541
rect 1574 532 1577 542
rect 2286 538 2294 541
rect 1370 528 1371 532
rect 2034 528 2035 532
rect 762 518 763 522
rect 1501 518 1502 522
rect 1690 518 1691 522
rect 880 503 882 507
rect 886 503 889 507
rect 893 503 896 507
rect 1912 503 1914 507
rect 1918 503 1921 507
rect 1925 503 1928 507
rect 346 488 347 492
rect 1221 488 1222 492
rect 1461 488 1462 492
rect 1834 488 1835 492
rect 1702 474 1706 478
rect 94 471 98 474
rect 94 468 105 471
rect 270 471 274 474
rect 270 468 278 471
rect 778 468 785 471
rect 838 471 842 474
rect 830 468 842 471
rect 926 468 942 471
rect 974 468 982 471
rect 1654 468 1662 471
rect 1686 471 1690 474
rect 2206 472 2210 474
rect 1678 468 1690 471
rect 102 462 105 468
rect 110 458 129 461
rect 214 458 222 461
rect 286 458 305 461
rect 318 458 326 461
rect 494 458 513 461
rect 686 458 694 461
rect 754 458 761 461
rect 806 458 825 461
rect 882 458 897 461
rect 974 458 993 461
rect 1198 458 1206 461
rect 1366 458 1385 461
rect 1654 458 1673 461
rect 1718 458 1726 461
rect 1970 458 1977 461
rect 2094 458 2113 461
rect 2182 458 2190 461
rect 2250 458 2257 461
rect 126 448 129 458
rect 302 448 305 458
rect 494 448 497 458
rect 806 448 809 458
rect 974 448 977 458
rect 1234 448 1241 451
rect 1382 448 1385 458
rect 1654 448 1657 458
rect 2110 448 2113 458
rect 443 438 446 442
rect 1141 428 1142 432
rect 376 403 378 407
rect 382 403 385 407
rect 389 403 392 407
rect 1392 403 1394 407
rect 1398 403 1401 407
rect 1405 403 1408 407
rect 141 388 142 392
rect 293 388 294 392
rect 434 388 441 391
rect 565 388 566 392
rect 693 388 694 392
rect 730 388 731 392
rect 853 388 854 392
rect 1186 388 1187 392
rect 1229 388 1230 392
rect 395 368 398 372
rect 1029 368 1030 372
rect 1634 368 1641 371
rect 2202 368 2209 371
rect 766 366 770 368
rect 70 351 73 361
rect 70 348 89 351
rect 294 348 313 351
rect 358 348 374 351
rect 478 351 481 361
rect 462 348 481 351
rect 546 348 553 351
rect 638 351 641 361
rect 742 358 761 361
rect 638 348 657 351
rect 670 348 678 351
rect 798 351 801 361
rect 798 348 817 351
rect 834 348 841 351
rect 1014 351 1017 361
rect 22 338 33 341
rect 94 338 105 341
rect 110 338 121 341
rect 450 338 457 341
rect 670 341 673 348
rect 998 348 1017 351
rect 1030 348 1038 351
rect 1142 351 1145 361
rect 1126 348 1145 351
rect 1202 348 1217 351
rect 1286 348 1294 351
rect 1374 351 1377 361
rect 1386 358 1390 362
rect 1358 348 1377 351
rect 1562 348 1569 351
rect 1598 348 1606 351
rect 1646 351 1649 358
rect 1646 348 1665 351
rect 1726 348 1734 351
rect 1758 351 1761 361
rect 1742 348 1761 351
rect 1822 348 1830 351
rect 2022 351 2025 361
rect 2022 348 2041 351
rect 2174 351 2177 361
rect 2174 348 2193 351
rect 2238 348 2246 351
rect 662 338 673 341
rect 1114 338 1121 341
rect 2174 338 2182 341
rect 30 332 33 338
rect 102 332 105 338
rect 246 331 250 333
rect 246 328 257 331
rect 446 328 449 338
rect 1053 318 1054 322
rect 1618 318 1619 322
rect 880 303 882 307
rect 886 303 889 307
rect 893 303 896 307
rect 1912 303 1914 307
rect 1918 303 1921 307
rect 1925 303 1928 307
rect 1989 288 1990 292
rect 810 268 817 271
rect 978 268 985 271
rect 1862 268 1890 271
rect 2062 268 2070 271
rect 2094 271 2098 274
rect 2086 268 2098 271
rect 2133 268 2134 272
rect 178 258 193 261
rect 254 258 273 261
rect 550 258 569 261
rect 630 258 638 261
rect 798 258 817 261
rect 830 258 846 261
rect 914 258 921 261
rect 1446 258 1465 261
rect 1526 258 1534 261
rect 1646 258 1665 261
rect 1730 258 1737 261
rect 1818 258 1833 261
rect 2062 258 2081 261
rect 18 248 22 252
rect 270 248 273 258
rect 510 248 529 251
rect 566 248 569 258
rect 814 248 817 258
rect 1002 248 1009 251
rect 1462 248 1465 258
rect 1474 248 1478 252
rect 1646 248 1649 258
rect 2062 248 2065 258
rect 58 238 61 242
rect 376 203 378 207
rect 382 203 385 207
rect 389 203 392 207
rect 1392 203 1394 207
rect 1398 203 1401 207
rect 1405 203 1408 207
rect 1341 188 1342 192
rect 1461 188 1462 192
rect 2285 188 2286 192
rect 1670 168 1678 171
rect 1803 168 1806 172
rect 1938 168 1941 172
rect 58 148 65 151
rect 278 148 286 151
rect 346 148 353 151
rect 358 148 374 151
rect 394 148 401 151
rect 502 148 518 151
rect 590 151 593 161
rect 590 148 609 151
rect 662 151 665 161
rect 662 148 681 151
rect 462 141 465 148
rect 846 151 849 161
rect 1114 158 1118 162
rect 846 148 865 151
rect 1126 151 1129 161
rect 1106 148 1113 151
rect 1126 148 1145 151
rect 1230 151 1233 161
rect 1230 148 1249 151
rect 1406 151 1409 161
rect 1374 148 1409 151
rect 1442 148 1449 151
rect 1518 148 1526 151
rect 1702 151 1705 161
rect 1686 148 1705 151
rect 1718 148 1726 151
rect 1962 148 1977 151
rect 2086 151 2089 161
rect 2046 148 2065 151
rect 2070 148 2089 151
rect 2142 151 2145 161
rect 2270 151 2273 161
rect 2142 148 2161 151
rect 2254 148 2273 151
rect 454 138 465 141
rect 618 138 625 141
rect 662 138 670 141
rect 846 138 854 141
rect 870 138 886 141
rect 1366 138 1369 148
rect 2062 142 2065 148
rect 1698 138 1705 141
rect 1846 138 1857 141
rect 1898 138 1922 141
rect 2114 138 2121 141
rect 78 131 82 136
rect 66 128 82 131
rect 206 131 210 136
rect 194 128 210 131
rect 222 131 226 133
rect 222 128 233 131
rect 622 128 625 138
rect 766 133 770 138
rect 1854 132 1857 138
rect 1918 136 1922 138
rect 1306 118 1307 122
rect 880 103 882 107
rect 886 103 889 107
rect 893 103 896 107
rect 1912 103 1914 107
rect 1918 103 1921 107
rect 1925 103 1928 107
rect 141 88 142 92
rect 402 88 417 91
rect 2197 88 2198 92
rect 838 78 857 81
rect 862 78 873 81
rect 1754 78 1769 81
rect 30 68 38 71
rect 62 68 73 71
rect 226 68 233 71
rect 582 68 594 71
rect 646 68 649 78
rect 862 72 865 78
rect 870 68 881 71
rect 906 68 913 71
rect 1582 68 1590 71
rect 1646 71 1650 74
rect 1846 72 1849 81
rect 1638 68 1650 71
rect 1806 68 1814 71
rect 1894 71 1897 81
rect 1894 68 1913 71
rect 1966 71 1969 81
rect 1938 68 1953 71
rect 1966 68 1985 71
rect 62 62 65 68
rect 22 58 41 61
rect 46 58 54 61
rect 86 58 106 61
rect 194 58 201 61
rect 334 58 350 61
rect 446 58 465 61
rect 870 62 873 68
rect 718 58 726 61
rect 806 58 814 61
rect 886 58 902 61
rect 934 58 953 61
rect 1134 58 1142 61
rect 1542 58 1561 61
rect 1586 58 1601 61
rect 1614 58 1633 61
rect 1782 58 1801 61
rect 1814 58 1817 68
rect 1918 58 1926 61
rect 2138 58 2153 61
rect 38 52 41 58
rect 462 48 465 58
rect 934 48 937 58
rect 1558 48 1561 58
rect 1614 48 1617 58
rect 1758 42 1762 44
rect 376 3 378 7
rect 382 3 385 7
rect 389 3 392 7
rect 1392 3 1394 7
rect 1398 3 1401 7
rect 1405 3 1408 7
<< m2contact >>
rect 882 2103 886 2107
rect 889 2103 893 2107
rect 1914 2103 1918 2107
rect 1921 2103 1925 2107
rect 1510 2088 1514 2092
rect 1846 2088 1850 2092
rect 2110 2088 2114 2092
rect 1294 2078 1298 2082
rect 6 2068 10 2072
rect 78 2068 82 2072
rect 142 2068 146 2072
rect 158 2068 162 2072
rect 246 2068 250 2072
rect 302 2068 306 2072
rect 318 2068 322 2072
rect 350 2068 354 2072
rect 462 2068 466 2072
rect 550 2068 554 2072
rect 566 2068 570 2072
rect 606 2068 610 2072
rect 670 2068 674 2072
rect 822 2068 826 2072
rect 838 2068 842 2072
rect 894 2068 898 2072
rect 926 2068 930 2072
rect 1022 2068 1026 2072
rect 1110 2068 1114 2072
rect 1166 2068 1170 2072
rect 1174 2068 1178 2072
rect 1206 2068 1210 2072
rect 1246 2068 1250 2072
rect 1366 2068 1370 2072
rect 1430 2068 1434 2072
rect 1518 2068 1522 2072
rect 1566 2068 1570 2072
rect 1686 2068 1690 2072
rect 1702 2068 1706 2072
rect 1734 2068 1738 2072
rect 1750 2068 1754 2072
rect 1886 2068 1890 2072
rect 1974 2068 1978 2072
rect 2030 2068 2034 2072
rect 2054 2068 2058 2072
rect 2078 2068 2082 2072
rect 2086 2068 2090 2072
rect 2166 2068 2170 2072
rect 2222 2068 2226 2072
rect 2230 2068 2234 2072
rect 2302 2068 2306 2072
rect 182 2058 186 2062
rect 254 2058 258 2062
rect 286 2058 290 2062
rect 294 2058 298 2062
rect 334 2059 338 2063
rect 446 2058 450 2062
rect 486 2058 490 2062
rect 558 2058 562 2062
rect 638 2058 642 2062
rect 678 2058 682 2062
rect 774 2058 778 2062
rect 806 2059 810 2063
rect 846 2058 850 2062
rect 878 2058 882 2062
rect 902 2058 906 2062
rect 942 2059 946 2063
rect 974 2058 978 2062
rect 1046 2058 1050 2062
rect 1118 2058 1122 2062
rect 1126 2058 1130 2062
rect 1158 2058 1162 2062
rect 1182 2058 1186 2062
rect 1198 2058 1202 2062
rect 1214 2058 1218 2062
rect 1262 2059 1266 2063
rect 1454 2058 1458 2062
rect 1526 2058 1530 2062
rect 1534 2058 1538 2062
rect 1574 2058 1578 2062
rect 1670 2059 1674 2063
rect 1710 2058 1714 2062
rect 1782 2059 1786 2063
rect 1814 2058 1818 2062
rect 1902 2058 1906 2062
rect 1982 2058 1986 2062
rect 2014 2058 2018 2062
rect 2022 2058 2026 2062
rect 2038 2058 2042 2062
rect 2150 2058 2154 2062
rect 2238 2058 2242 2062
rect 2246 2058 2250 2062
rect 1142 2048 1146 2052
rect 1198 2048 1202 2052
rect 1550 2048 1554 2052
rect 1734 2048 1738 2052
rect 1830 2048 1834 2052
rect 2062 2048 2066 2052
rect 2102 2048 2106 2052
rect 2206 2048 2210 2052
rect 2254 2048 2258 2052
rect 270 2038 274 2042
rect 430 2038 434 2042
rect 542 2038 546 2042
rect 582 2038 586 2042
rect 862 2038 866 2042
rect 1086 2038 1090 2042
rect 1102 2038 1106 2042
rect 1214 2038 1218 2042
rect 1230 2038 1234 2042
rect 1326 2038 1330 2042
rect 1494 2038 1498 2042
rect 398 2028 402 2032
rect 1006 2028 1010 2032
rect 62 2018 66 2022
rect 238 2018 242 2022
rect 622 2018 626 2022
rect 734 2018 738 2022
rect 742 2018 746 2022
rect 1342 2018 1346 2022
rect 1390 2018 1394 2022
rect 1590 2018 1594 2022
rect 1606 2018 1610 2022
rect 1862 2018 1866 2022
rect 1998 2018 2002 2022
rect 2094 2018 2098 2022
rect 2214 2018 2218 2022
rect 2270 2018 2274 2022
rect 378 2003 382 2007
rect 385 2003 389 2007
rect 1394 2003 1398 2007
rect 1401 2003 1405 2007
rect 182 1988 186 1992
rect 750 1988 754 1992
rect 1766 1988 1770 1992
rect 6 1978 10 1982
rect 134 1968 138 1972
rect 150 1968 154 1972
rect 198 1968 202 1972
rect 214 1968 218 1972
rect 254 1968 258 1972
rect 382 1968 386 1972
rect 478 1968 482 1972
rect 774 1968 778 1972
rect 878 1968 882 1972
rect 1054 1968 1058 1972
rect 1262 1968 1266 1972
rect 1278 1968 1282 1972
rect 1358 1968 1362 1972
rect 1414 1968 1418 1972
rect 1926 1968 1930 1972
rect 2078 1968 2082 1972
rect 102 1958 106 1962
rect 166 1958 170 1962
rect 70 1947 74 1951
rect 102 1948 106 1952
rect 118 1948 122 1952
rect 150 1948 154 1952
rect 182 1948 186 1952
rect 230 1948 234 1952
rect 502 1958 506 1962
rect 606 1958 610 1962
rect 734 1958 738 1962
rect 278 1948 282 1952
rect 318 1947 322 1951
rect 350 1948 354 1952
rect 454 1948 458 1952
rect 518 1948 522 1952
rect 542 1948 546 1952
rect 566 1948 570 1952
rect 574 1948 578 1952
rect 590 1948 594 1952
rect 638 1947 642 1951
rect 718 1948 722 1952
rect 750 1948 754 1952
rect 806 1958 810 1962
rect 862 1958 866 1962
rect 910 1958 914 1962
rect 1038 1958 1042 1962
rect 1070 1958 1074 1962
rect 790 1948 794 1952
rect 814 1948 818 1952
rect 822 1948 826 1952
rect 846 1948 850 1952
rect 878 1948 882 1952
rect 942 1947 946 1951
rect 974 1948 978 1952
rect 1022 1948 1026 1952
rect 1054 1948 1058 1952
rect 1102 1947 1106 1951
rect 1214 1948 1218 1952
rect 1278 1948 1282 1952
rect 1302 1958 1306 1962
rect 1318 1948 1322 1952
rect 1382 1958 1386 1962
rect 1382 1948 1386 1952
rect 1470 1948 1474 1952
rect 1574 1947 1578 1951
rect 1614 1948 1618 1952
rect 1638 1958 1642 1962
rect 1710 1948 1714 1952
rect 1766 1948 1770 1952
rect 1790 1958 1794 1962
rect 1822 1948 1826 1952
rect 1846 1948 1850 1952
rect 1854 1948 1858 1952
rect 1870 1948 1874 1952
rect 1894 1958 1898 1962
rect 1966 1948 1970 1952
rect 1990 1948 1994 1952
rect 2038 1948 2042 1952
rect 2062 1958 2066 1962
rect 2206 1958 2210 1962
rect 2118 1948 2122 1952
rect 2142 1948 2146 1952
rect 2190 1948 2194 1952
rect 2246 1948 2250 1952
rect 2254 1948 2258 1952
rect 62 1938 66 1942
rect 126 1938 130 1942
rect 158 1938 162 1942
rect 190 1938 194 1942
rect 230 1938 234 1942
rect 270 1938 274 1942
rect 286 1938 290 1942
rect 414 1938 418 1942
rect 502 1938 506 1942
rect 526 1938 530 1942
rect 582 1938 586 1942
rect 606 1938 610 1942
rect 622 1938 626 1942
rect 710 1938 714 1942
rect 726 1938 730 1942
rect 742 1938 746 1942
rect 798 1938 802 1942
rect 830 1938 834 1942
rect 862 1938 866 1942
rect 870 1938 874 1942
rect 1014 1938 1018 1942
rect 1038 1938 1042 1942
rect 1046 1938 1050 1942
rect 1086 1938 1090 1942
rect 1270 1938 1274 1942
rect 1326 1938 1330 1942
rect 1390 1938 1394 1942
rect 1494 1938 1498 1942
rect 1590 1938 1594 1942
rect 1606 1938 1610 1942
rect 1630 1938 1634 1942
rect 1710 1938 1714 1942
rect 1758 1938 1762 1942
rect 1806 1938 1810 1942
rect 1862 1938 1866 1942
rect 1894 1938 1898 1942
rect 1926 1938 1930 1942
rect 2030 1938 2034 1942
rect 2054 1938 2058 1942
rect 2078 1938 2082 1942
rect 2166 1938 2170 1942
rect 2182 1938 2186 1942
rect 1198 1928 1202 1932
rect 494 1918 498 1922
rect 558 1918 562 1922
rect 702 1918 706 1922
rect 1006 1918 1010 1922
rect 1166 1918 1170 1922
rect 1510 1918 1514 1922
rect 1662 1918 1666 1922
rect 1838 1918 1842 1922
rect 2206 1918 2210 1922
rect 2214 1918 2218 1922
rect 882 1903 886 1907
rect 889 1903 893 1907
rect 1914 1903 1918 1907
rect 1921 1903 1925 1907
rect 582 1888 586 1892
rect 662 1888 666 1892
rect 1142 1888 1146 1892
rect 1326 1888 1330 1892
rect 1622 1888 1626 1892
rect 2078 1888 2082 1892
rect 2254 1888 2258 1892
rect 838 1878 842 1882
rect 1102 1878 1106 1882
rect 1286 1878 1290 1882
rect 1526 1878 1530 1882
rect 1662 1878 1666 1882
rect 1790 1878 1794 1882
rect 2046 1878 2050 1882
rect 102 1868 106 1872
rect 126 1868 130 1872
rect 158 1868 162 1872
rect 262 1868 266 1872
rect 278 1868 282 1872
rect 326 1868 330 1872
rect 462 1868 466 1872
rect 518 1868 522 1872
rect 574 1868 578 1872
rect 606 1868 610 1872
rect 686 1868 690 1872
rect 718 1868 722 1872
rect 726 1868 730 1872
rect 902 1868 906 1872
rect 918 1868 922 1872
rect 942 1868 946 1872
rect 990 1868 994 1872
rect 1158 1868 1162 1872
rect 1190 1868 1194 1872
rect 1214 1868 1218 1872
rect 1318 1868 1322 1872
rect 1406 1868 1410 1872
rect 1438 1868 1442 1872
rect 1470 1868 1474 1872
rect 1494 1868 1498 1872
rect 1598 1868 1602 1872
rect 1646 1868 1650 1872
rect 1686 1868 1690 1872
rect 1766 1868 1770 1872
rect 1814 1868 1818 1872
rect 1854 1868 1858 1872
rect 2174 1868 2178 1872
rect 2190 1868 2194 1872
rect 2222 1868 2226 1872
rect 2230 1868 2234 1872
rect 2278 1868 2282 1872
rect 46 1858 50 1862
rect 62 1858 66 1862
rect 118 1858 122 1862
rect 126 1858 130 1862
rect 150 1858 154 1862
rect 198 1858 202 1862
rect 222 1858 226 1862
rect 270 1858 274 1862
rect 334 1858 338 1862
rect 382 1858 386 1862
rect 406 1858 410 1862
rect 414 1858 418 1862
rect 470 1858 474 1862
rect 526 1858 530 1862
rect 534 1858 538 1862
rect 566 1858 570 1862
rect 598 1858 602 1862
rect 614 1858 618 1862
rect 622 1858 626 1862
rect 646 1858 650 1862
rect 678 1858 682 1862
rect 686 1858 690 1862
rect 734 1858 738 1862
rect 758 1858 762 1862
rect 766 1858 770 1862
rect 838 1859 842 1863
rect 894 1858 898 1862
rect 934 1858 938 1862
rect 950 1858 954 1862
rect 958 1858 962 1862
rect 982 1858 986 1862
rect 998 1858 1002 1862
rect 1006 1858 1010 1862
rect 1046 1858 1050 1862
rect 1078 1858 1082 1862
rect 1086 1858 1090 1862
rect 1118 1858 1122 1862
rect 1166 1858 1170 1862
rect 1206 1858 1210 1862
rect 1270 1858 1274 1862
rect 1350 1858 1354 1862
rect 1374 1858 1378 1862
rect 1390 1858 1394 1862
rect 1414 1858 1418 1862
rect 1446 1858 1450 1862
rect 1470 1858 1474 1862
rect 1478 1858 1482 1862
rect 1526 1859 1530 1863
rect 1638 1858 1642 1862
rect 1710 1858 1714 1862
rect 1734 1859 1738 1863
rect 1806 1858 1810 1862
rect 1822 1858 1826 1862
rect 1830 1858 1834 1862
rect 1862 1858 1866 1862
rect 1870 1858 1874 1862
rect 1878 1858 1882 1862
rect 1902 1858 1906 1862
rect 1934 1858 1938 1862
rect 1942 1858 1946 1862
rect 1966 1858 1970 1862
rect 1982 1858 1986 1862
rect 1990 1858 1994 1862
rect 2014 1858 2018 1862
rect 2030 1858 2034 1862
rect 2038 1858 2042 1862
rect 2070 1858 2074 1862
rect 2110 1858 2114 1862
rect 2142 1859 2146 1863
rect 2214 1858 2218 1862
rect 2270 1858 2274 1862
rect 102 1848 106 1852
rect 550 1848 554 1852
rect 582 1848 586 1852
rect 662 1848 666 1852
rect 870 1848 874 1852
rect 918 1848 922 1852
rect 1182 1848 1186 1852
rect 1462 1848 1466 1852
rect 1494 1848 1498 1852
rect 1614 1848 1618 1852
rect 1782 1848 1786 1852
rect 2190 1848 2194 1852
rect 2246 1848 2250 1852
rect 94 1838 98 1842
rect 134 1838 138 1842
rect 254 1838 258 1842
rect 294 1838 298 1842
rect 350 1838 354 1842
rect 774 1838 778 1842
rect 886 1838 890 1842
rect 1222 1838 1226 1842
rect 1430 1838 1434 1842
rect 1590 1838 1594 1842
rect 1022 1828 1026 1832
rect 334 1818 338 1822
rect 398 1818 402 1822
rect 510 1818 514 1822
rect 638 1818 642 1822
rect 710 1818 714 1822
rect 1358 1818 1362 1822
rect 1414 1818 1418 1822
rect 1654 1818 1658 1822
rect 1670 1818 1674 1822
rect 1894 1818 1898 1822
rect 1950 1818 1954 1822
rect 1998 1818 2002 1822
rect 378 1803 382 1807
rect 385 1803 389 1807
rect 1394 1803 1398 1807
rect 1401 1803 1405 1807
rect 62 1788 66 1792
rect 334 1788 338 1792
rect 622 1788 626 1792
rect 758 1788 762 1792
rect 974 1788 978 1792
rect 1430 1788 1434 1792
rect 1758 1788 1762 1792
rect 1902 1788 1906 1792
rect 2158 1778 2162 1782
rect 526 1768 530 1772
rect 862 1768 866 1772
rect 1158 1768 1162 1772
rect 1254 1768 1258 1772
rect 1710 1768 1714 1772
rect 1726 1768 1730 1772
rect 342 1758 346 1762
rect 110 1748 114 1752
rect 142 1747 146 1751
rect 286 1748 290 1752
rect 342 1748 346 1752
rect 358 1748 362 1752
rect 398 1748 402 1752
rect 422 1748 426 1752
rect 430 1748 434 1752
rect 478 1748 482 1752
rect 542 1748 546 1752
rect 550 1748 554 1752
rect 566 1758 570 1762
rect 582 1748 586 1752
rect 598 1748 602 1752
rect 606 1748 610 1752
rect 630 1748 634 1752
rect 654 1748 658 1752
rect 662 1748 666 1752
rect 678 1748 682 1752
rect 686 1748 690 1752
rect 694 1748 698 1752
rect 702 1748 706 1752
rect 726 1748 730 1752
rect 734 1748 738 1752
rect 822 1748 826 1752
rect 878 1748 882 1752
rect 886 1748 890 1752
rect 918 1758 922 1762
rect 1006 1758 1010 1762
rect 1062 1758 1066 1762
rect 934 1748 938 1752
rect 1006 1748 1010 1752
rect 1046 1748 1050 1752
rect 1126 1758 1130 1762
rect 1142 1758 1146 1762
rect 1310 1758 1314 1762
rect 1414 1758 1418 1762
rect 1086 1748 1090 1752
rect 1110 1748 1114 1752
rect 1142 1748 1146 1752
rect 6 1738 10 1742
rect 174 1738 178 1742
rect 254 1738 258 1742
rect 366 1738 370 1742
rect 462 1738 466 1742
rect 534 1738 538 1742
rect 590 1738 594 1742
rect 782 1738 786 1742
rect 870 1738 874 1742
rect 942 1738 946 1742
rect 990 1738 994 1742
rect 1190 1747 1194 1751
rect 1294 1748 1298 1752
rect 1302 1748 1306 1752
rect 1334 1748 1338 1752
rect 1366 1748 1370 1752
rect 1374 1748 1378 1752
rect 1382 1748 1386 1752
rect 1390 1748 1394 1752
rect 1422 1748 1426 1752
rect 1462 1748 1466 1752
rect 1478 1748 1482 1752
rect 1534 1748 1538 1752
rect 1558 1758 1562 1762
rect 1590 1748 1594 1752
rect 1614 1758 1618 1762
rect 1830 1758 1834 1762
rect 1854 1758 1858 1762
rect 1862 1758 1866 1762
rect 1950 1758 1954 1762
rect 2150 1758 2154 1762
rect 2270 1758 2274 1762
rect 1014 1738 1018 1742
rect 1038 1738 1042 1742
rect 1078 1738 1082 1742
rect 1094 1738 1098 1742
rect 1102 1738 1106 1742
rect 1126 1738 1130 1742
rect 1134 1738 1138 1742
rect 1198 1738 1202 1742
rect 1318 1738 1322 1742
rect 1326 1738 1330 1742
rect 1662 1747 1666 1751
rect 1734 1748 1738 1752
rect 1742 1748 1746 1752
rect 1766 1748 1770 1752
rect 1782 1748 1786 1752
rect 1886 1748 1890 1752
rect 1894 1748 1898 1752
rect 1942 1748 1946 1752
rect 1982 1748 1986 1752
rect 1990 1748 1994 1752
rect 2046 1748 2050 1752
rect 2102 1748 2106 1752
rect 2190 1748 2194 1752
rect 2222 1747 2226 1751
rect 2294 1748 2298 1752
rect 1526 1738 1530 1742
rect 1542 1738 1546 1742
rect 1574 1738 1578 1742
rect 1582 1738 1586 1742
rect 1614 1738 1618 1742
rect 1630 1738 1634 1742
rect 1806 1738 1810 1742
rect 1838 1738 1842 1742
rect 1878 1738 1882 1742
rect 1966 1738 1970 1742
rect 1998 1738 2002 1742
rect 2086 1738 2090 1742
rect 2126 1738 2130 1742
rect 2134 1738 2138 1742
rect 2254 1738 2258 1742
rect 2278 1738 2282 1742
rect 2302 1738 2306 1742
rect 1662 1728 1666 1732
rect 62 1718 66 1722
rect 78 1718 82 1722
rect 230 1718 234 1722
rect 414 1718 418 1722
rect 718 1718 722 1722
rect 1022 1718 1026 1722
rect 1278 1718 1282 1722
rect 1350 1718 1354 1722
rect 1798 1718 1802 1722
rect 1822 1718 1826 1722
rect 1846 1718 1850 1722
rect 1862 1718 1866 1722
rect 2006 1718 2010 1722
rect 2142 1718 2146 1722
rect 882 1703 886 1707
rect 889 1703 893 1707
rect 1914 1703 1918 1707
rect 1921 1703 1925 1707
rect 142 1688 146 1692
rect 862 1688 866 1692
rect 1150 1688 1154 1692
rect 1502 1688 1506 1692
rect 1942 1688 1946 1692
rect 102 1678 106 1682
rect 326 1678 330 1682
rect 542 1678 546 1682
rect 678 1678 682 1682
rect 1518 1678 1522 1682
rect 2030 1678 2034 1682
rect 118 1668 122 1672
rect 166 1668 170 1672
rect 198 1668 202 1672
rect 302 1668 306 1672
rect 350 1668 354 1672
rect 518 1668 522 1672
rect 574 1668 578 1672
rect 710 1668 714 1672
rect 766 1668 770 1672
rect 782 1668 786 1672
rect 910 1668 914 1672
rect 942 1668 946 1672
rect 998 1668 1002 1672
rect 1046 1668 1050 1672
rect 1422 1668 1426 1672
rect 1462 1668 1466 1672
rect 1550 1668 1554 1672
rect 1558 1668 1562 1672
rect 1590 1668 1594 1672
rect 1678 1668 1682 1672
rect 1694 1668 1698 1672
rect 1726 1668 1730 1672
rect 1766 1668 1770 1672
rect 1822 1668 1826 1672
rect 1846 1668 1850 1672
rect 1894 1668 1898 1672
rect 2078 1668 2082 1672
rect 2110 1668 2114 1672
rect 2158 1668 2162 1672
rect 2182 1668 2186 1672
rect 2206 1668 2210 1672
rect 2214 1668 2218 1672
rect 2238 1668 2242 1672
rect 30 1659 34 1663
rect 62 1658 66 1662
rect 158 1658 162 1662
rect 174 1658 178 1662
rect 238 1658 242 1662
rect 254 1658 258 1662
rect 366 1658 370 1662
rect 422 1658 426 1662
rect 430 1658 434 1662
rect 478 1658 482 1662
rect 502 1658 506 1662
rect 510 1658 514 1662
rect 526 1658 530 1662
rect 566 1658 570 1662
rect 574 1658 578 1662
rect 614 1658 618 1662
rect 622 1658 626 1662
rect 646 1658 650 1662
rect 662 1658 666 1662
rect 670 1658 674 1662
rect 694 1658 698 1662
rect 702 1658 706 1662
rect 750 1658 754 1662
rect 758 1658 762 1662
rect 798 1659 802 1663
rect 870 1658 874 1662
rect 894 1658 898 1662
rect 934 1658 938 1662
rect 950 1658 954 1662
rect 958 1658 962 1662
rect 982 1658 986 1662
rect 1006 1658 1010 1662
rect 1022 1658 1026 1662
rect 1086 1659 1090 1663
rect 1118 1658 1122 1662
rect 1158 1658 1162 1662
rect 1166 1658 1170 1662
rect 1190 1658 1194 1662
rect 1238 1658 1242 1662
rect 1246 1658 1250 1662
rect 1262 1658 1266 1662
rect 1286 1658 1290 1662
rect 1294 1658 1298 1662
rect 1302 1658 1306 1662
rect 1334 1658 1338 1662
rect 1342 1658 1346 1662
rect 1358 1658 1362 1662
rect 1382 1658 1386 1662
rect 1390 1658 1394 1662
rect 1446 1658 1450 1662
rect 1534 1658 1538 1662
rect 1542 1658 1546 1662
rect 1558 1658 1562 1662
rect 1614 1658 1618 1662
rect 1718 1658 1722 1662
rect 1750 1658 1754 1662
rect 1774 1658 1778 1662
rect 1782 1658 1786 1662
rect 1830 1658 1834 1662
rect 1878 1659 1882 1663
rect 1966 1658 1970 1662
rect 1974 1658 1978 1662
rect 1998 1658 2002 1662
rect 2014 1658 2018 1662
rect 2022 1658 2026 1662
rect 2126 1659 2130 1663
rect 2198 1658 2202 1662
rect 134 1648 138 1652
rect 318 1648 322 1652
rect 550 1648 554 1652
rect 598 1648 602 1652
rect 734 1648 738 1652
rect 918 1648 922 1652
rect 974 1648 978 1652
rect 1022 1648 1026 1652
rect 1318 1648 1322 1652
rect 1526 1648 1530 1652
rect 1574 1648 1578 1652
rect 1694 1648 1698 1652
rect 1758 1648 1762 1652
rect 1782 1648 1786 1652
rect 1846 1648 1850 1652
rect 1990 1648 1994 1652
rect 2174 1648 2178 1652
rect 2230 1648 2234 1652
rect 302 1638 306 1642
rect 1678 1638 1682 1642
rect 1742 1638 1746 1642
rect 94 1618 98 1622
rect 110 1618 114 1622
rect 494 1618 498 1622
rect 638 1618 642 1622
rect 1006 1618 1010 1622
rect 1230 1618 1234 1622
rect 1278 1618 1282 1622
rect 1374 1618 1378 1622
rect 1510 1618 1514 1622
rect 1750 1618 1754 1622
rect 1806 1618 1810 1622
rect 2222 1618 2226 1622
rect 2294 1618 2298 1622
rect 378 1603 382 1607
rect 385 1603 389 1607
rect 1394 1603 1398 1607
rect 1401 1603 1405 1607
rect 22 1588 26 1592
rect 830 1588 834 1592
rect 974 1588 978 1592
rect 1294 1588 1298 1592
rect 2014 1588 2018 1592
rect 2166 1588 2170 1592
rect 438 1568 442 1572
rect 614 1568 618 1572
rect 630 1568 634 1572
rect 958 1568 962 1572
rect 998 1568 1002 1572
rect 1382 1568 1386 1572
rect 1454 1568 1458 1572
rect 1582 1568 1586 1572
rect 1606 1568 1610 1572
rect 1854 1568 1858 1572
rect 1990 1568 1994 1572
rect 6 1558 10 1562
rect 38 1558 42 1562
rect 118 1558 122 1562
rect 38 1548 42 1552
rect 62 1548 66 1552
rect 102 1548 106 1552
rect 150 1547 154 1551
rect 182 1548 186 1552
rect 254 1548 258 1552
rect 278 1548 282 1552
rect 358 1548 362 1552
rect 438 1548 442 1552
rect 462 1558 466 1562
rect 646 1558 650 1562
rect 478 1548 482 1552
rect 494 1548 498 1552
rect 526 1548 530 1552
rect 534 1548 538 1552
rect 582 1548 586 1552
rect 646 1548 650 1552
rect 670 1558 674 1562
rect 862 1558 866 1562
rect 982 1558 986 1562
rect 1006 1558 1010 1562
rect 1038 1558 1042 1562
rect 1286 1558 1290 1562
rect 1438 1558 1442 1562
rect 1486 1558 1490 1562
rect 1574 1558 1578 1562
rect 1598 1558 1602 1562
rect 1702 1558 1706 1562
rect 1718 1558 1722 1562
rect 1798 1558 1802 1562
rect 710 1548 714 1552
rect 734 1548 738 1552
rect 790 1548 794 1552
rect 846 1548 850 1552
rect 854 1548 858 1552
rect 926 1548 930 1552
rect 982 1548 986 1552
rect 1014 1548 1018 1552
rect 1022 1548 1026 1552
rect 1094 1548 1098 1552
rect 1118 1548 1122 1552
rect 1190 1548 1194 1552
rect 1214 1548 1218 1552
rect 1278 1548 1282 1552
rect 1358 1548 1362 1552
rect 1470 1548 1474 1552
rect 1494 1548 1498 1552
rect 1550 1548 1554 1552
rect 1566 1548 1570 1552
rect 30 1538 34 1542
rect 54 1538 58 1542
rect 86 1538 90 1542
rect 94 1538 98 1542
rect 118 1538 122 1542
rect 166 1538 170 1542
rect 326 1538 330 1542
rect 430 1538 434 1542
rect 486 1538 490 1542
rect 550 1538 554 1542
rect 582 1538 586 1542
rect 638 1538 642 1542
rect 686 1538 690 1542
rect 750 1538 754 1542
rect 798 1538 802 1542
rect 838 1538 842 1542
rect 894 1538 898 1542
rect 1670 1547 1674 1551
rect 1718 1548 1722 1552
rect 1734 1548 1738 1552
rect 1742 1548 1746 1552
rect 1782 1548 1786 1552
rect 1814 1548 1818 1552
rect 1838 1558 1842 1562
rect 1902 1548 1906 1552
rect 1998 1548 2002 1552
rect 2006 1548 2010 1552
rect 2030 1548 2034 1552
rect 2070 1548 2074 1552
rect 2086 1548 2090 1552
rect 2110 1558 2114 1562
rect 2134 1558 2138 1562
rect 2262 1558 2266 1562
rect 2134 1548 2138 1552
rect 2150 1548 2154 1552
rect 2222 1548 2226 1552
rect 2278 1548 2282 1552
rect 998 1538 1002 1542
rect 1030 1538 1034 1542
rect 1054 1538 1058 1542
rect 1086 1538 1090 1542
rect 1166 1538 1170 1542
rect 1198 1538 1202 1542
rect 1302 1538 1306 1542
rect 1318 1538 1322 1542
rect 1454 1538 1458 1542
rect 1462 1538 1466 1542
rect 1558 1538 1562 1542
rect 1574 1538 1578 1542
rect 1686 1538 1690 1542
rect 1726 1538 1730 1542
rect 1782 1538 1786 1542
rect 1798 1538 1802 1542
rect 1830 1538 1834 1542
rect 1942 1538 1946 1542
rect 1974 1538 1978 1542
rect 2046 1538 2050 1542
rect 2078 1538 2082 1542
rect 2126 1538 2130 1542
rect 2158 1538 2162 1542
rect 2246 1538 2250 1542
rect 2270 1538 2274 1542
rect 2286 1538 2290 1542
rect 2302 1538 2306 1542
rect 38 1528 42 1532
rect 1406 1528 1410 1532
rect 1430 1528 1434 1532
rect 1518 1528 1522 1532
rect 214 1518 218 1522
rect 310 1518 314 1522
rect 406 1518 410 1522
rect 510 1518 514 1522
rect 702 1518 706 1522
rect 1046 1518 1050 1522
rect 1150 1518 1154 1522
rect 1246 1518 1250 1522
rect 1262 1518 1266 1522
rect 1398 1518 1402 1522
rect 1510 1518 1514 1522
rect 1534 1518 1538 1522
rect 1750 1518 1754 1522
rect 1798 1518 1802 1522
rect 1982 1518 1986 1522
rect 2102 1518 2106 1522
rect 882 1503 886 1507
rect 889 1503 893 1507
rect 1914 1503 1918 1507
rect 1921 1503 1925 1507
rect 94 1488 98 1492
rect 182 1488 186 1492
rect 230 1488 234 1492
rect 422 1488 426 1492
rect 846 1488 850 1492
rect 910 1488 914 1492
rect 966 1488 970 1492
rect 1006 1488 1010 1492
rect 1062 1488 1066 1492
rect 1134 1488 1138 1492
rect 1206 1488 1210 1492
rect 1238 1488 1242 1492
rect 1334 1488 1338 1492
rect 1646 1488 1650 1492
rect 2054 1488 2058 1492
rect 2166 1488 2170 1492
rect 238 1478 242 1482
rect 254 1478 258 1482
rect 814 1478 818 1482
rect 1030 1478 1034 1482
rect 1102 1478 1106 1482
rect 1142 1478 1146 1482
rect 1174 1478 1178 1482
rect 1542 1478 1546 1482
rect 1990 1478 1994 1482
rect 2070 1478 2074 1482
rect 2262 1478 2266 1482
rect 46 1468 50 1472
rect 102 1468 106 1472
rect 150 1468 154 1472
rect 198 1468 202 1472
rect 206 1468 210 1472
rect 302 1468 306 1472
rect 334 1468 338 1472
rect 366 1468 370 1472
rect 390 1468 394 1472
rect 446 1468 450 1472
rect 38 1458 42 1462
rect 110 1458 114 1462
rect 118 1458 122 1462
rect 174 1458 178 1462
rect 214 1458 218 1462
rect 278 1458 282 1462
rect 294 1458 298 1462
rect 318 1458 322 1462
rect 326 1458 330 1462
rect 342 1458 346 1462
rect 398 1458 402 1462
rect 438 1458 442 1462
rect 446 1458 450 1462
rect 478 1468 482 1472
rect 534 1468 538 1472
rect 574 1468 578 1472
rect 582 1468 586 1472
rect 646 1468 650 1472
rect 702 1468 706 1472
rect 774 1468 778 1472
rect 790 1468 794 1472
rect 822 1468 826 1472
rect 870 1468 874 1472
rect 958 1468 962 1472
rect 1070 1468 1074 1472
rect 1166 1468 1170 1472
rect 1182 1468 1186 1472
rect 1230 1468 1234 1472
rect 1254 1468 1258 1472
rect 1278 1468 1282 1472
rect 1286 1468 1290 1472
rect 1318 1468 1322 1472
rect 1358 1468 1362 1472
rect 1366 1468 1370 1472
rect 1390 1468 1394 1472
rect 1406 1468 1410 1472
rect 1422 1468 1426 1472
rect 1454 1468 1458 1472
rect 1470 1468 1474 1472
rect 1478 1468 1482 1472
rect 1486 1468 1490 1472
rect 1686 1468 1690 1472
rect 1726 1468 1730 1472
rect 1742 1468 1746 1472
rect 1790 1468 1794 1472
rect 1878 1468 1882 1472
rect 1894 1468 1898 1472
rect 1926 1468 1930 1472
rect 1958 1468 1962 1472
rect 2070 1468 2074 1472
rect 2174 1468 2178 1472
rect 2238 1468 2242 1472
rect 2246 1468 2250 1472
rect 470 1458 474 1462
rect 518 1458 522 1462
rect 590 1458 594 1462
rect 654 1458 658 1462
rect 662 1458 666 1462
rect 694 1458 698 1462
rect 742 1458 746 1462
rect 750 1458 754 1462
rect 782 1458 786 1462
rect 806 1458 810 1462
rect 862 1458 866 1462
rect 910 1458 914 1462
rect 934 1458 938 1462
rect 990 1458 994 1462
rect 1014 1458 1018 1462
rect 1046 1458 1050 1462
rect 1094 1458 1098 1462
rect 1126 1458 1130 1462
rect 1142 1458 1146 1462
rect 1190 1458 1194 1462
rect 1278 1458 1282 1462
rect 1294 1458 1298 1462
rect 1318 1458 1322 1462
rect 1358 1458 1362 1462
rect 1414 1458 1418 1462
rect 1454 1458 1458 1462
rect 1494 1458 1498 1462
rect 1510 1458 1514 1462
rect 1550 1458 1554 1462
rect 1566 1458 1570 1462
rect 1582 1458 1586 1462
rect 1590 1458 1594 1462
rect 1606 1458 1610 1462
rect 1630 1458 1634 1462
rect 1638 1458 1642 1462
rect 1710 1459 1714 1463
rect 1750 1458 1754 1462
rect 1758 1458 1762 1462
rect 1838 1458 1842 1462
rect 1902 1458 1906 1462
rect 1934 1458 1938 1462
rect 1990 1459 1994 1463
rect 2022 1458 2026 1462
rect 2102 1459 2106 1463
rect 2134 1458 2138 1462
rect 2182 1458 2186 1462
rect 2198 1458 2202 1462
rect 2230 1459 2234 1463
rect 134 1448 138 1452
rect 174 1448 178 1452
rect 182 1448 186 1452
rect 230 1448 234 1452
rect 254 1448 258 1452
rect 310 1448 314 1452
rect 414 1448 418 1452
rect 422 1448 426 1452
rect 454 1448 458 1452
rect 678 1448 682 1452
rect 734 1448 738 1452
rect 846 1448 850 1452
rect 926 1448 930 1452
rect 990 1448 994 1452
rect 1022 1448 1026 1452
rect 1046 1448 1050 1452
rect 1134 1448 1138 1452
rect 1214 1448 1218 1452
rect 1238 1448 1242 1452
rect 1262 1448 1266 1452
rect 1310 1448 1314 1452
rect 1334 1448 1338 1452
rect 1366 1448 1370 1452
rect 1438 1448 1442 1452
rect 1502 1448 1506 1452
rect 1774 1448 1778 1452
rect 1926 1448 1930 1452
rect 1942 1448 1946 1452
rect 2198 1448 2202 1452
rect 294 1438 298 1442
rect 638 1438 642 1442
rect 838 1438 842 1442
rect 918 1438 922 1442
rect 942 1438 946 1442
rect 998 1438 1002 1442
rect 1054 1438 1058 1442
rect 1518 1438 1522 1442
rect 1542 1438 1546 1442
rect 1790 1438 1794 1442
rect 1118 1428 1122 1432
rect 398 1418 402 1422
rect 494 1418 498 1422
rect 718 1418 722 1422
rect 910 1418 914 1422
rect 934 1418 938 1422
rect 1006 1418 1010 1422
rect 1326 1418 1330 1422
rect 1526 1418 1530 1422
rect 1622 1418 1626 1422
rect 2062 1418 2066 1422
rect 2294 1418 2298 1422
rect 378 1403 382 1407
rect 385 1403 389 1407
rect 1394 1403 1398 1407
rect 1401 1403 1405 1407
rect 246 1388 250 1392
rect 726 1388 730 1392
rect 998 1388 1002 1392
rect 1174 1388 1178 1392
rect 1206 1388 1210 1392
rect 1230 1388 1234 1392
rect 1534 1388 1538 1392
rect 1830 1388 1834 1392
rect 374 1378 378 1382
rect 102 1368 106 1372
rect 806 1368 810 1372
rect 1038 1368 1042 1372
rect 1054 1368 1058 1372
rect 1126 1368 1130 1372
rect 1166 1368 1170 1372
rect 1198 1368 1202 1372
rect 1222 1368 1226 1372
rect 1254 1368 1258 1372
rect 1654 1368 1658 1372
rect 1846 1368 1850 1372
rect 1886 1368 1890 1372
rect 2086 1368 2090 1372
rect 118 1358 122 1362
rect 38 1348 42 1352
rect 278 1358 282 1362
rect 142 1348 146 1352
rect 206 1348 210 1352
rect 262 1348 266 1352
rect 270 1348 274 1352
rect 326 1348 330 1352
rect 398 1348 402 1352
rect 414 1348 418 1352
rect 430 1358 434 1362
rect 462 1358 466 1362
rect 614 1358 618 1362
rect 630 1358 634 1362
rect 734 1358 738 1362
rect 766 1358 770 1362
rect 790 1358 794 1362
rect 846 1358 850 1362
rect 1022 1358 1026 1362
rect 1054 1358 1058 1362
rect 1150 1358 1154 1362
rect 1190 1358 1194 1362
rect 1238 1358 1242 1362
rect 1270 1358 1274 1362
rect 1310 1358 1314 1362
rect 1350 1358 1354 1362
rect 1414 1358 1418 1362
rect 1430 1358 1434 1362
rect 1470 1358 1474 1362
rect 1486 1358 1490 1362
rect 1558 1358 1562 1362
rect 1606 1358 1610 1362
rect 1630 1358 1634 1362
rect 1638 1358 1642 1362
rect 1670 1358 1674 1362
rect 1710 1358 1714 1362
rect 1726 1358 1730 1362
rect 446 1348 450 1352
rect 486 1348 490 1352
rect 510 1348 514 1352
rect 550 1348 554 1352
rect 574 1348 578 1352
rect 678 1348 682 1352
rect 734 1348 738 1352
rect 750 1348 754 1352
rect 798 1348 802 1352
rect 830 1348 834 1352
rect 838 1348 842 1352
rect 46 1338 50 1342
rect 102 1338 106 1342
rect 118 1338 122 1342
rect 150 1338 154 1342
rect 166 1338 170 1342
rect 254 1338 258 1342
rect 294 1338 298 1342
rect 334 1338 338 1342
rect 398 1338 402 1342
rect 454 1338 458 1342
rect 478 1338 482 1342
rect 894 1347 898 1351
rect 982 1348 986 1352
rect 1014 1348 1018 1352
rect 1030 1348 1034 1352
rect 1062 1348 1066 1352
rect 1110 1348 1114 1352
rect 1134 1348 1138 1352
rect 1158 1348 1162 1352
rect 1190 1348 1194 1352
rect 1230 1348 1234 1352
rect 1262 1348 1266 1352
rect 1294 1348 1298 1352
rect 1326 1348 1330 1352
rect 1366 1348 1370 1352
rect 1382 1348 1386 1352
rect 1430 1348 1434 1352
rect 1454 1348 1458 1352
rect 1534 1348 1538 1352
rect 1582 1348 1586 1352
rect 1630 1348 1634 1352
rect 1646 1348 1650 1352
rect 1702 1348 1706 1352
rect 1710 1348 1714 1352
rect 1742 1348 1746 1352
rect 1766 1358 1770 1362
rect 1806 1358 1810 1362
rect 1982 1358 1986 1362
rect 2046 1358 2050 1362
rect 1830 1348 1834 1352
rect 1926 1348 1930 1352
rect 1998 1348 2002 1352
rect 2070 1358 2074 1362
rect 2070 1348 2074 1352
rect 2142 1348 2146 1352
rect 2214 1348 2218 1352
rect 2238 1348 2242 1352
rect 614 1338 618 1342
rect 646 1338 650 1342
rect 758 1338 762 1342
rect 782 1338 786 1342
rect 822 1338 826 1342
rect 878 1338 882 1342
rect 966 1338 970 1342
rect 1086 1338 1090 1342
rect 1278 1338 1282 1342
rect 1334 1338 1338 1342
rect 1358 1338 1362 1342
rect 1390 1338 1394 1342
rect 1438 1338 1442 1342
rect 1446 1338 1450 1342
rect 1462 1338 1466 1342
rect 1534 1338 1538 1342
rect 1582 1338 1586 1342
rect 1590 1338 1594 1342
rect 1614 1338 1618 1342
rect 1662 1338 1666 1342
rect 1694 1338 1698 1342
rect 1702 1338 1706 1342
rect 1734 1338 1738 1342
rect 1758 1338 1762 1342
rect 1782 1338 1786 1342
rect 1790 1338 1794 1342
rect 1838 1338 1842 1342
rect 1862 1338 1866 1342
rect 1950 1338 1954 1342
rect 1966 1338 1970 1342
rect 2006 1338 2010 1342
rect 2030 1338 2034 1342
rect 2078 1338 2082 1342
rect 2134 1338 2138 1342
rect 2302 1338 2306 1342
rect 182 1328 186 1332
rect 214 1328 218 1332
rect 798 1328 802 1332
rect 966 1328 970 1332
rect 1278 1328 1282 1332
rect 1486 1328 1490 1332
rect 462 1318 466 1322
rect 606 1318 610 1322
rect 726 1318 730 1322
rect 766 1318 770 1322
rect 958 1318 962 1322
rect 1046 1318 1050 1322
rect 1078 1318 1082 1322
rect 1118 1318 1122 1322
rect 1158 1318 1162 1322
rect 1262 1318 1266 1322
rect 1350 1318 1354 1322
rect 1382 1318 1386 1322
rect 1502 1318 1506 1322
rect 1606 1318 1610 1322
rect 1670 1318 1674 1322
rect 1854 1318 1858 1322
rect 1982 1318 1986 1322
rect 2014 1318 2018 1322
rect 2270 1318 2274 1322
rect 882 1303 886 1307
rect 889 1303 893 1307
rect 1914 1303 1918 1307
rect 1921 1303 1925 1307
rect 422 1288 426 1292
rect 534 1288 538 1292
rect 942 1288 946 1292
rect 1150 1288 1154 1292
rect 1342 1288 1346 1292
rect 1414 1288 1418 1292
rect 1526 1288 1530 1292
rect 1694 1288 1698 1292
rect 1718 1288 1722 1292
rect 1798 1288 1802 1292
rect 1894 1288 1898 1292
rect 1958 1288 1962 1292
rect 2038 1288 2042 1292
rect 2190 1288 2194 1292
rect 134 1278 138 1282
rect 246 1278 250 1282
rect 446 1278 450 1282
rect 566 1278 570 1282
rect 638 1278 642 1282
rect 742 1278 746 1282
rect 750 1278 754 1282
rect 766 1278 770 1282
rect 774 1278 778 1282
rect 990 1278 994 1282
rect 1086 1278 1090 1282
rect 30 1268 34 1272
rect 118 1268 122 1272
rect 182 1268 186 1272
rect 262 1268 266 1272
rect 318 1268 322 1272
rect 334 1268 338 1272
rect 478 1268 482 1272
rect 502 1268 506 1272
rect 510 1268 514 1272
rect 2102 1278 2106 1282
rect 630 1268 634 1272
rect 782 1268 786 1272
rect 806 1268 810 1272
rect 830 1268 834 1272
rect 870 1268 874 1272
rect 966 1268 970 1272
rect 982 1268 986 1272
rect 1062 1268 1066 1272
rect 1094 1268 1098 1272
rect 1166 1268 1170 1272
rect 1182 1268 1186 1272
rect 1286 1268 1290 1272
rect 1374 1268 1378 1272
rect 1382 1268 1386 1272
rect 1446 1268 1450 1272
rect 1454 1268 1458 1272
rect 1518 1268 1522 1272
rect 1622 1268 1626 1272
rect 1646 1268 1650 1272
rect 1686 1268 1690 1272
rect 1742 1268 1746 1272
rect 1766 1268 1770 1272
rect 1790 1268 1794 1272
rect 1878 1268 1882 1272
rect 1934 1268 1938 1272
rect 2030 1268 2034 1272
rect 2078 1268 2082 1272
rect 2134 1268 2138 1272
rect 2182 1268 2186 1272
rect 2238 1268 2242 1272
rect 22 1258 26 1262
rect 94 1258 98 1262
rect 190 1258 194 1262
rect 270 1258 274 1262
rect 278 1258 282 1262
rect 310 1258 314 1262
rect 358 1258 362 1262
rect 454 1258 458 1262
rect 470 1258 474 1262
rect 518 1258 522 1262
rect 590 1258 594 1262
rect 694 1258 698 1262
rect 702 1258 706 1262
rect 790 1258 794 1262
rect 862 1259 866 1263
rect 974 1258 978 1262
rect 1014 1258 1018 1262
rect 1038 1258 1042 1262
rect 1070 1258 1074 1262
rect 1086 1258 1090 1262
rect 1118 1258 1122 1262
rect 1150 1258 1154 1262
rect 1182 1258 1186 1262
rect 1198 1258 1202 1262
rect 1246 1258 1250 1262
rect 1294 1258 1298 1262
rect 1358 1258 1362 1262
rect 1366 1258 1370 1262
rect 1422 1258 1426 1262
rect 1438 1258 1442 1262
rect 1470 1258 1474 1262
rect 1494 1258 1498 1262
rect 1558 1258 1562 1262
rect 1590 1259 1594 1263
rect 1638 1258 1642 1262
rect 1670 1258 1674 1262
rect 1742 1258 1746 1262
rect 1750 1258 1754 1262
rect 1838 1258 1842 1262
rect 1910 1258 1914 1262
rect 1942 1258 1946 1262
rect 1982 1258 1986 1262
rect 1998 1258 2002 1262
rect 2006 1258 2010 1262
rect 2022 1258 2026 1262
rect 2070 1258 2074 1262
rect 2086 1258 2090 1262
rect 2094 1258 2098 1262
rect 2166 1258 2170 1262
rect 2182 1258 2186 1262
rect 2246 1258 2250 1262
rect 2286 1258 2290 1262
rect 6 1248 10 1252
rect 22 1248 26 1252
rect 294 1248 298 1252
rect 454 1248 458 1252
rect 542 1248 546 1252
rect 814 1248 818 1252
rect 950 1248 954 1252
rect 1022 1248 1026 1252
rect 1054 1248 1058 1252
rect 1126 1248 1130 1252
rect 1158 1248 1162 1252
rect 1190 1248 1194 1252
rect 1350 1248 1354 1252
rect 1398 1248 1402 1252
rect 1414 1248 1418 1252
rect 1470 1248 1474 1252
rect 1478 1248 1482 1252
rect 1622 1248 1626 1252
rect 1678 1248 1682 1252
rect 1702 1248 1706 1252
rect 1774 1248 1778 1252
rect 1894 1248 1898 1252
rect 2054 1248 2058 1252
rect 2150 1248 2154 1252
rect 614 1238 618 1242
rect 750 1238 754 1242
rect 1006 1238 1010 1242
rect 1038 1238 1042 1242
rect 1110 1238 1114 1242
rect 1150 1238 1154 1242
rect 1206 1238 1210 1242
rect 1662 1238 1666 1242
rect 2206 1238 2210 1242
rect 2302 1238 2306 1242
rect 38 1218 42 1222
rect 142 1218 146 1222
rect 238 1218 242 1222
rect 254 1218 258 1222
rect 438 1218 442 1222
rect 494 1218 498 1222
rect 590 1218 594 1222
rect 646 1218 650 1222
rect 742 1218 746 1222
rect 926 1218 930 1222
rect 1014 1218 1018 1222
rect 1046 1218 1050 1222
rect 1118 1218 1122 1222
rect 1134 1218 1138 1222
rect 1198 1218 1202 1222
rect 1230 1218 1234 1222
rect 1462 1218 1466 1222
rect 1654 1218 1658 1222
rect 378 1203 382 1207
rect 385 1203 389 1207
rect 1394 1203 1398 1207
rect 1401 1203 1405 1207
rect 14 1188 18 1192
rect 446 1188 450 1192
rect 694 1188 698 1192
rect 814 1188 818 1192
rect 1102 1188 1106 1192
rect 1142 1188 1146 1192
rect 1246 1188 1250 1192
rect 1622 1188 1626 1192
rect 2102 1188 2106 1192
rect 134 1168 138 1172
rect 174 1168 178 1172
rect 406 1168 410 1172
rect 718 1168 722 1172
rect 830 1168 834 1172
rect 1022 1168 1026 1172
rect 1174 1168 1178 1172
rect 1238 1168 1242 1172
rect 1310 1168 1314 1172
rect 2022 1168 2026 1172
rect 78 1148 82 1152
rect 102 1148 106 1152
rect 150 1148 154 1152
rect 158 1148 162 1152
rect 374 1158 378 1162
rect 422 1158 426 1162
rect 486 1158 490 1162
rect 190 1148 194 1152
rect 230 1148 234 1152
rect 246 1148 250 1152
rect 270 1148 274 1152
rect 286 1148 290 1152
rect 350 1148 354 1152
rect 358 1148 362 1152
rect 406 1148 410 1152
rect 430 1148 434 1152
rect 470 1148 474 1152
rect 502 1148 506 1152
rect 510 1148 514 1152
rect 574 1148 578 1152
rect 654 1148 658 1152
rect 694 1148 698 1152
rect 958 1158 962 1162
rect 734 1148 738 1152
rect 758 1148 762 1152
rect 774 1148 778 1152
rect 790 1148 794 1152
rect 870 1148 874 1152
rect 1014 1158 1018 1162
rect 1038 1158 1042 1162
rect 894 1147 898 1151
rect 982 1148 986 1152
rect 1038 1148 1042 1152
rect 1054 1148 1058 1152
rect 1078 1158 1082 1162
rect 1118 1158 1122 1162
rect 1190 1158 1194 1162
rect 1230 1158 1234 1162
rect 1254 1158 1258 1162
rect 1438 1158 1442 1162
rect 1142 1148 1146 1152
rect 1182 1148 1186 1152
rect 1214 1148 1218 1152
rect 1230 1148 1234 1152
rect 1278 1148 1282 1152
rect 1534 1158 1538 1162
rect 1558 1158 1562 1162
rect 1606 1158 1610 1162
rect 1630 1158 1634 1162
rect 1662 1158 1666 1162
rect 1734 1158 1738 1162
rect 1750 1158 1754 1162
rect 1806 1158 1810 1162
rect 1822 1158 1826 1162
rect 1830 1158 1834 1162
rect 1886 1158 1890 1162
rect 2094 1158 2098 1162
rect 6 1138 10 1142
rect 142 1138 146 1142
rect 198 1138 202 1142
rect 222 1138 226 1142
rect 254 1138 258 1142
rect 262 1138 266 1142
rect 350 1138 354 1142
rect 398 1138 402 1142
rect 462 1138 466 1142
rect 518 1138 522 1142
rect 606 1138 610 1142
rect 622 1138 626 1142
rect 638 1138 642 1142
rect 686 1138 690 1142
rect 742 1138 746 1142
rect 750 1138 754 1142
rect 782 1138 786 1142
rect 806 1138 810 1142
rect 926 1138 930 1142
rect 966 1138 970 1142
rect 990 1138 994 1142
rect 998 1138 1002 1142
rect 1038 1138 1042 1142
rect 1374 1147 1378 1151
rect 1462 1148 1466 1152
rect 1518 1148 1522 1152
rect 1574 1148 1578 1152
rect 1638 1148 1642 1152
rect 1670 1148 1674 1152
rect 1734 1148 1738 1152
rect 1798 1148 1802 1152
rect 1806 1148 1810 1152
rect 1854 1148 1858 1152
rect 1886 1148 1890 1152
rect 1926 1148 1930 1152
rect 1958 1147 1962 1151
rect 2038 1148 2042 1152
rect 2062 1148 2066 1152
rect 2070 1148 2074 1152
rect 2166 1147 2170 1151
rect 2230 1148 2234 1152
rect 1094 1138 1098 1142
rect 1134 1138 1138 1142
rect 1198 1138 1202 1142
rect 1270 1138 1274 1142
rect 1390 1138 1394 1142
rect 1422 1138 1426 1142
rect 1446 1138 1450 1142
rect 1470 1138 1474 1142
rect 1494 1138 1498 1142
rect 1534 1138 1538 1142
rect 1550 1138 1554 1142
rect 1566 1138 1570 1142
rect 1582 1138 1586 1142
rect 1590 1138 1594 1142
rect 1614 1138 1618 1142
rect 1646 1138 1650 1142
rect 1678 1138 1682 1142
rect 1758 1138 1762 1142
rect 1782 1138 1786 1142
rect 1798 1138 1802 1142
rect 1846 1138 1850 1142
rect 1862 1138 1866 1142
rect 1918 1138 1922 1142
rect 1966 1138 1970 1142
rect 2030 1138 2034 1142
rect 2078 1138 2082 1142
rect 206 1128 210 1132
rect 310 1128 314 1132
rect 326 1128 330 1132
rect 646 1128 650 1132
rect 774 1128 778 1132
rect 798 1128 802 1132
rect 1110 1128 1114 1132
rect 1158 1128 1162 1132
rect 1214 1128 1218 1132
rect 1478 1128 1482 1132
rect 1662 1128 1666 1132
rect 1694 1128 1698 1132
rect 1766 1128 1770 1132
rect 2166 1128 2170 1132
rect 2222 1128 2226 1132
rect 214 1118 218 1122
rect 230 1118 234 1122
rect 270 1118 274 1122
rect 374 1118 378 1122
rect 526 1118 530 1122
rect 670 1118 674 1122
rect 1014 1118 1018 1122
rect 1070 1118 1074 1122
rect 1118 1118 1122 1122
rect 1182 1118 1186 1122
rect 1262 1118 1266 1122
rect 1294 1118 1298 1122
rect 1518 1118 1522 1122
rect 1542 1118 1546 1122
rect 1606 1118 1610 1122
rect 1686 1118 1690 1122
rect 1710 1118 1714 1122
rect 1830 1118 1834 1122
rect 2086 1118 2090 1122
rect 2286 1118 2290 1122
rect 882 1103 886 1107
rect 889 1103 893 1107
rect 1914 1103 1918 1107
rect 1921 1103 1925 1107
rect 14 1088 18 1092
rect 190 1088 194 1092
rect 294 1088 298 1092
rect 566 1088 570 1092
rect 974 1088 978 1092
rect 1126 1088 1130 1092
rect 1142 1088 1146 1092
rect 1190 1088 1194 1092
rect 1670 1088 1674 1092
rect 1846 1088 1850 1092
rect 2102 1088 2106 1092
rect 2286 1088 2290 1092
rect 30 1078 34 1082
rect 318 1078 322 1082
rect 422 1078 426 1082
rect 574 1078 578 1082
rect 942 1078 946 1082
rect 1174 1078 1178 1082
rect 46 1068 50 1072
rect 94 1068 98 1072
rect 110 1068 114 1072
rect 198 1068 202 1072
rect 246 1068 250 1072
rect 254 1068 258 1072
rect 318 1068 322 1072
rect 486 1068 490 1072
rect 590 1068 594 1072
rect 614 1068 618 1072
rect 638 1068 642 1072
rect 654 1068 658 1072
rect 702 1068 706 1072
rect 774 1068 778 1072
rect 806 1068 810 1072
rect 838 1068 842 1072
rect 862 1068 866 1072
rect 878 1068 882 1072
rect 982 1068 986 1072
rect 1030 1068 1034 1072
rect 1062 1068 1066 1072
rect 1134 1068 1138 1072
rect 1238 1068 1242 1072
rect 1270 1068 1274 1072
rect 1286 1068 1290 1072
rect 1374 1068 1378 1072
rect 1390 1068 1394 1072
rect 1438 1068 1442 1072
rect 1550 1078 1554 1082
rect 1566 1078 1570 1082
rect 1630 1078 1634 1082
rect 1678 1078 1682 1082
rect 2166 1078 2170 1082
rect 1486 1068 1490 1072
rect 1494 1068 1498 1072
rect 1598 1068 1602 1072
rect 1606 1068 1610 1072
rect 1662 1068 1666 1072
rect 1750 1068 1754 1072
rect 30 1058 34 1062
rect 94 1058 98 1062
rect 150 1058 154 1062
rect 206 1058 210 1062
rect 214 1058 218 1062
rect 262 1058 266 1062
rect 374 1059 378 1063
rect 406 1058 410 1062
rect 446 1058 450 1062
rect 526 1058 530 1062
rect 630 1058 634 1062
rect 678 1058 682 1062
rect 742 1058 746 1062
rect 1806 1068 1810 1072
rect 1830 1068 1834 1072
rect 1838 1068 1842 1072
rect 1862 1068 1866 1072
rect 1886 1068 1890 1072
rect 2014 1068 2018 1072
rect 2030 1068 2034 1072
rect 2070 1068 2074 1072
rect 2206 1068 2210 1072
rect 782 1058 786 1062
rect 790 1058 794 1062
rect 814 1058 818 1062
rect 854 1058 858 1062
rect 918 1058 922 1062
rect 990 1058 994 1062
rect 1070 1058 1074 1062
rect 1158 1058 1162 1062
rect 1206 1058 1210 1062
rect 1214 1058 1218 1062
rect 1262 1058 1266 1062
rect 1310 1058 1314 1062
rect 1374 1058 1378 1062
rect 1462 1058 1466 1062
rect 1478 1058 1482 1062
rect 1486 1058 1490 1062
rect 1550 1058 1554 1062
rect 1566 1058 1570 1062
rect 1590 1058 1594 1062
rect 1598 1058 1602 1062
rect 1638 1058 1642 1062
rect 1654 1058 1658 1062
rect 1742 1058 1746 1062
rect 1782 1058 1786 1062
rect 1822 1058 1826 1062
rect 1870 1058 1874 1062
rect 1974 1058 1978 1062
rect 2046 1058 2050 1062
rect 2078 1058 2082 1062
rect 2094 1058 2098 1062
rect 2150 1058 2154 1062
rect 2230 1058 2234 1062
rect 6 1048 10 1052
rect 46 1048 50 1052
rect 62 1048 66 1052
rect 86 1048 90 1052
rect 230 1048 234 1052
rect 278 1048 282 1052
rect 606 1048 610 1052
rect 830 1048 834 1052
rect 990 1048 994 1052
rect 1014 1048 1018 1052
rect 1246 1048 1250 1052
rect 1262 1048 1266 1052
rect 1422 1048 1426 1052
rect 1462 1048 1466 1052
rect 1478 1048 1482 1052
rect 1518 1048 1522 1052
rect 1542 1048 1546 1052
rect 1574 1048 1578 1052
rect 1590 1048 1594 1052
rect 1638 1048 1642 1052
rect 1798 1048 1802 1052
rect 1854 1048 1858 1052
rect 1894 1048 1898 1052
rect 2094 1048 2098 1052
rect 590 1038 594 1042
rect 734 1038 738 1042
rect 798 1038 802 1042
rect 1366 1038 1370 1042
rect 1678 1038 1682 1042
rect 262 1018 266 1022
rect 334 1018 338 1022
rect 438 1018 442 1022
rect 462 1018 466 1022
rect 1142 1018 1146 1022
rect 1158 1018 1162 1022
rect 1654 1018 1658 1022
rect 1918 1018 1922 1022
rect 378 1003 382 1007
rect 385 1003 389 1007
rect 1394 1003 1398 1007
rect 1401 1003 1405 1007
rect 6 988 10 992
rect 742 988 746 992
rect 798 988 802 992
rect 950 988 954 992
rect 974 988 978 992
rect 1206 988 1210 992
rect 1294 988 1298 992
rect 1526 988 1530 992
rect 1590 988 1594 992
rect 302 968 306 972
rect 326 968 330 972
rect 502 968 506 972
rect 526 968 530 972
rect 654 968 658 972
rect 678 968 682 972
rect 942 968 946 972
rect 1806 968 1810 972
rect 1918 968 1922 972
rect 2142 968 2146 972
rect 2222 968 2226 972
rect 2238 968 2242 972
rect 2294 968 2298 972
rect 118 958 122 962
rect 70 947 74 951
rect 134 948 138 952
rect 142 948 146 952
rect 166 948 170 952
rect 190 958 194 962
rect 342 958 346 962
rect 406 958 410 962
rect 454 958 458 962
rect 494 958 498 962
rect 518 958 522 962
rect 542 958 546 962
rect 574 958 578 962
rect 694 958 698 962
rect 238 947 242 951
rect 390 948 394 952
rect 414 948 418 952
rect 438 948 442 952
rect 454 948 458 952
rect 478 948 482 952
rect 558 948 562 952
rect 614 948 618 952
rect 638 948 642 952
rect 790 958 794 962
rect 926 958 930 962
rect 958 958 962 962
rect 966 958 970 962
rect 1006 958 1010 962
rect 1014 958 1018 962
rect 1046 958 1050 962
rect 1070 958 1074 962
rect 1142 958 1146 962
rect 1230 958 1234 962
rect 1310 958 1314 962
rect 1478 958 1482 962
rect 1510 958 1514 962
rect 718 948 722 952
rect 758 948 762 952
rect 774 948 778 952
rect 790 948 794 952
rect 854 948 858 952
rect 950 948 954 952
rect 1022 948 1026 952
rect 1030 948 1034 952
rect 1094 948 1098 952
rect 1126 948 1130 952
rect 1134 948 1138 952
rect 1198 948 1202 952
rect 1222 948 1226 952
rect 1246 948 1250 952
rect 1286 948 1290 952
rect 1326 948 1330 952
rect 1358 948 1362 952
rect 1422 948 1426 952
rect 1438 948 1442 952
rect 1478 948 1482 952
rect 1494 948 1498 952
rect 1526 948 1530 952
rect 1566 948 1570 952
rect 46 938 50 942
rect 86 938 90 942
rect 102 938 106 942
rect 150 938 154 942
rect 158 938 162 942
rect 190 938 194 942
rect 206 938 210 942
rect 246 938 250 942
rect 326 938 330 942
rect 1630 947 1634 951
rect 1662 948 1666 952
rect 1742 948 1746 952
rect 1758 948 1762 952
rect 1798 948 1802 952
rect 1830 958 1834 962
rect 1958 958 1962 962
rect 2022 958 2026 962
rect 1878 948 1882 952
rect 1918 948 1922 952
rect 1958 948 1962 952
rect 1982 948 1986 952
rect 1990 948 1994 952
rect 2022 948 2026 952
rect 2038 948 2042 952
rect 462 938 466 942
rect 470 938 474 942
rect 542 938 546 942
rect 550 938 554 942
rect 678 938 682 942
rect 694 938 698 942
rect 726 938 730 942
rect 766 938 770 942
rect 854 938 858 942
rect 878 938 882 942
rect 894 938 898 942
rect 982 938 986 942
rect 990 938 994 942
rect 1038 938 1042 942
rect 1070 938 1074 942
rect 1086 938 1090 942
rect 1102 938 1106 942
rect 1158 938 1162 942
rect 1254 938 1258 942
rect 1262 938 1266 942
rect 1278 938 1282 942
rect 1326 938 1330 942
rect 1358 938 1362 942
rect 1502 938 1506 942
rect 1542 938 1546 942
rect 1798 938 1802 942
rect 1846 938 1850 942
rect 1886 938 1890 942
rect 1918 938 1922 942
rect 2078 947 2082 951
rect 2110 948 2114 952
rect 2174 947 2178 951
rect 2206 948 2210 952
rect 2270 948 2274 952
rect 1998 938 2002 942
rect 2046 938 2050 942
rect 2062 938 2066 942
rect 2158 938 2162 942
rect 2262 938 2266 942
rect 310 928 314 932
rect 318 928 322 932
rect 350 928 354 932
rect 414 928 418 932
rect 574 928 578 932
rect 654 928 658 932
rect 1302 928 1306 932
rect 518 918 522 922
rect 798 918 802 922
rect 926 918 930 922
rect 1006 918 1010 922
rect 1046 918 1050 922
rect 1070 918 1074 922
rect 1150 918 1154 922
rect 1174 918 1178 922
rect 1206 918 1210 922
rect 1238 918 1242 922
rect 1270 918 1274 922
rect 1470 918 1474 922
rect 1550 918 1554 922
rect 1694 918 1698 922
rect 1790 918 1794 922
rect 1862 918 1866 922
rect 1894 918 1898 922
rect 882 903 886 907
rect 889 903 893 907
rect 1914 903 1918 907
rect 1921 903 1925 907
rect 94 888 98 892
rect 382 888 386 892
rect 518 888 522 892
rect 694 888 698 892
rect 790 888 794 892
rect 1078 888 1082 892
rect 1206 888 1210 892
rect 1302 888 1306 892
rect 1310 888 1314 892
rect 1486 888 1490 892
rect 1606 888 1610 892
rect 1654 888 1658 892
rect 1830 888 1834 892
rect 2246 888 2250 892
rect 2286 888 2290 892
rect 46 868 50 872
rect 126 868 130 872
rect 166 868 170 872
rect 222 868 226 872
rect 262 868 266 872
rect 302 868 306 872
rect 406 868 410 872
rect 422 868 426 872
rect 438 868 442 872
rect 486 868 490 872
rect 526 868 530 872
rect 574 868 578 872
rect 646 878 650 882
rect 854 878 858 882
rect 1142 878 1146 882
rect 1582 878 1586 882
rect 1614 878 1618 882
rect 1646 878 1650 882
rect 1686 878 1690 882
rect 1774 878 1778 882
rect 598 868 602 872
rect 630 868 634 872
rect 654 868 658 872
rect 46 858 50 862
rect 62 858 66 862
rect 102 858 106 862
rect 126 858 130 862
rect 142 858 146 862
rect 174 858 178 862
rect 214 858 218 862
rect 238 858 242 862
rect 254 858 258 862
rect 270 858 274 862
rect 318 859 322 863
rect 750 868 754 872
rect 902 868 906 872
rect 934 868 938 872
rect 958 868 962 872
rect 462 858 466 862
rect 534 858 538 862
rect 542 858 546 862
rect 606 858 610 862
rect 622 858 626 862
rect 646 858 650 862
rect 662 858 666 862
rect 678 858 682 862
rect 766 858 770 862
rect 822 858 826 862
rect 854 859 858 863
rect 1086 868 1090 872
rect 1126 868 1130 872
rect 1142 868 1146 872
rect 1182 868 1186 872
rect 1406 868 1410 872
rect 1438 868 1442 872
rect 1470 868 1474 872
rect 1494 868 1498 872
rect 1518 868 1522 872
rect 1534 868 1538 872
rect 1550 868 1554 872
rect 1566 868 1570 872
rect 1598 868 1602 872
rect 1630 868 1634 872
rect 1678 868 1682 872
rect 1710 868 1714 872
rect 1766 868 1770 872
rect 1790 868 1794 872
rect 1806 868 1810 872
rect 1838 868 1842 872
rect 1854 868 1858 872
rect 1926 868 1930 872
rect 1958 868 1962 872
rect 1974 868 1978 872
rect 2014 868 2018 872
rect 2062 868 2066 872
rect 2142 868 2146 872
rect 2206 868 2210 872
rect 2222 868 2226 872
rect 2270 868 2274 872
rect 2278 868 2282 872
rect 910 858 914 862
rect 966 858 970 862
rect 982 858 986 862
rect 1014 859 1018 863
rect 1046 858 1050 862
rect 1094 858 1098 862
rect 1166 858 1170 862
rect 1190 858 1194 862
rect 1246 858 1250 862
rect 1262 858 1266 862
rect 1342 858 1346 862
rect 1374 859 1378 863
rect 1462 858 1466 862
rect 1526 858 1530 862
rect 1558 858 1562 862
rect 1622 858 1626 862
rect 1670 858 1674 862
rect 1686 858 1690 862
rect 1702 858 1706 862
rect 1718 858 1722 862
rect 1766 858 1770 862
rect 1782 858 1786 862
rect 1798 858 1802 862
rect 1814 858 1818 862
rect 1870 858 1874 862
rect 1894 858 1898 862
rect 1902 858 1906 862
rect 1926 858 1930 862
rect 1934 858 1938 862
rect 2038 858 2042 862
rect 2078 858 2082 862
rect 2086 858 2090 862
rect 2190 859 2194 863
rect 2262 858 2266 862
rect 102 848 106 852
rect 134 848 138 852
rect 254 848 258 852
rect 270 848 274 852
rect 286 848 290 852
rect 422 848 426 852
rect 558 848 562 852
rect 678 848 682 852
rect 758 848 762 852
rect 910 848 914 852
rect 926 848 930 852
rect 950 848 954 852
rect 982 848 986 852
rect 1110 848 1114 852
rect 1174 848 1178 852
rect 1206 848 1210 852
rect 1438 848 1442 852
rect 1478 848 1482 852
rect 1494 848 1498 852
rect 1550 848 1554 852
rect 1654 848 1658 852
rect 1742 848 1746 852
rect 1758 848 1762 852
rect 1830 848 1834 852
rect 1838 848 1842 852
rect 1958 848 1962 852
rect 2238 848 2242 852
rect 2294 848 2298 852
rect 190 838 194 842
rect 774 838 778 842
rect 934 838 938 842
rect 1734 838 1738 842
rect 2142 838 2146 842
rect 214 818 218 822
rect 590 818 594 822
rect 622 818 626 822
rect 694 818 698 822
rect 766 818 770 822
rect 790 818 794 822
rect 1510 818 1514 822
rect 1646 818 1650 822
rect 1886 818 1890 822
rect 2094 818 2098 822
rect 378 803 382 807
rect 385 803 389 807
rect 1394 803 1398 807
rect 1401 803 1405 807
rect 302 788 306 792
rect 446 788 450 792
rect 1110 788 1114 792
rect 1142 788 1146 792
rect 1174 788 1178 792
rect 1598 788 1602 792
rect 1702 788 1706 792
rect 1782 788 1786 792
rect 1814 788 1818 792
rect 1870 788 1874 792
rect 1934 788 1938 792
rect 2270 788 2274 792
rect 94 768 98 772
rect 110 768 114 772
rect 1062 768 1066 772
rect 1150 768 1154 772
rect 1726 768 1730 772
rect 1806 768 1810 772
rect 2062 768 2066 772
rect 46 748 50 752
rect 62 748 66 752
rect 110 748 114 752
rect 134 758 138 762
rect 166 748 170 752
rect 190 758 194 762
rect 462 758 466 762
rect 494 758 498 762
rect 534 758 538 762
rect 238 747 242 751
rect 270 748 274 752
rect 318 748 322 752
rect 334 748 338 752
rect 406 748 410 752
rect 422 748 426 752
rect 446 748 450 752
rect 478 748 482 752
rect 502 748 506 752
rect 558 748 562 752
rect 582 758 586 762
rect 614 758 618 762
rect 622 758 626 762
rect 598 748 602 752
rect 614 748 618 752
rect 638 748 642 752
rect 662 748 666 752
rect 686 758 690 762
rect 742 748 746 752
rect 750 748 754 752
rect 806 748 810 752
rect 830 748 834 752
rect 838 748 842 752
rect 862 758 866 762
rect 1046 758 1050 762
rect 1078 758 1082 762
rect 1126 758 1130 762
rect 1134 758 1138 762
rect 1198 758 1202 762
rect 1214 758 1218 762
rect 934 748 938 752
rect 958 748 962 752
rect 998 748 1002 752
rect 1006 748 1010 752
rect 1030 748 1034 752
rect 1054 748 1058 752
rect 1110 748 1114 752
rect 1142 748 1146 752
rect 1246 748 1250 752
rect 1302 748 1306 752
rect 1310 748 1314 752
rect 1350 748 1354 752
rect 1366 748 1370 752
rect 1382 758 1386 762
rect 1430 748 1434 752
rect 1438 748 1442 752
rect 1454 758 1458 762
rect 1734 758 1738 762
rect 1822 758 1826 762
rect 1846 758 1850 762
rect 1918 758 1922 762
rect 2174 758 2178 762
rect 54 738 58 742
rect 102 738 106 742
rect 150 738 154 742
rect 158 738 162 742
rect 182 738 186 742
rect 206 738 210 742
rect 310 738 314 742
rect 326 738 330 742
rect 390 738 394 742
rect 414 738 418 742
rect 430 738 434 742
rect 438 738 442 742
rect 470 738 474 742
rect 526 738 530 742
rect 558 738 562 742
rect 582 738 586 742
rect 590 738 594 742
rect 1502 747 1506 751
rect 1646 748 1650 752
rect 1742 748 1746 752
rect 1750 748 1754 752
rect 1766 748 1770 752
rect 1814 748 1818 752
rect 1830 748 1834 752
rect 1854 748 1858 752
rect 1862 748 1866 752
rect 1886 748 1890 752
rect 1934 748 1938 752
rect 1966 748 1970 752
rect 1998 748 2002 752
rect 2006 748 2010 752
rect 2022 748 2026 752
rect 2046 748 2050 752
rect 2054 748 2058 752
rect 2126 747 2130 751
rect 2198 748 2202 752
rect 2286 748 2290 752
rect 646 738 650 742
rect 654 738 658 742
rect 678 738 682 742
rect 830 738 834 742
rect 862 738 866 742
rect 894 738 898 742
rect 1038 738 1042 742
rect 1078 738 1082 742
rect 1094 738 1098 742
rect 1102 738 1106 742
rect 1198 738 1202 742
rect 1222 738 1226 742
rect 1262 738 1266 742
rect 1350 738 1354 742
rect 1398 738 1402 742
rect 1422 738 1426 742
rect 1470 738 1474 742
rect 1486 738 1490 742
rect 1606 738 1610 742
rect 1654 738 1658 742
rect 1758 738 1762 742
rect 1830 738 1834 742
rect 1974 738 1978 742
rect 2014 738 2018 742
rect 2142 738 2146 742
rect 2158 738 2162 742
rect 2174 738 2178 742
rect 2206 738 2210 742
rect 2214 738 2218 742
rect 2302 738 2306 742
rect 358 728 362 732
rect 366 728 370 732
rect 806 728 810 732
rect 918 728 922 732
rect 1958 728 1962 732
rect 382 718 386 722
rect 494 718 498 722
rect 534 718 538 722
rect 622 718 626 722
rect 710 718 714 722
rect 894 718 898 722
rect 1062 718 1066 722
rect 1174 718 1178 722
rect 1214 718 1218 722
rect 1342 718 1346 722
rect 1566 718 1570 722
rect 1582 718 1586 722
rect 882 703 886 707
rect 889 703 893 707
rect 1914 703 1918 707
rect 1921 703 1925 707
rect 134 688 138 692
rect 310 688 314 692
rect 398 688 402 692
rect 502 688 506 692
rect 598 688 602 692
rect 670 688 674 692
rect 878 688 882 692
rect 950 688 954 692
rect 1086 688 1090 692
rect 1094 688 1098 692
rect 1126 688 1130 692
rect 1294 688 1298 692
rect 1494 688 1498 692
rect 1646 688 1650 692
rect 1694 688 1698 692
rect 1830 688 1834 692
rect 1838 688 1842 692
rect 1870 688 1874 692
rect 2118 688 2122 692
rect 358 678 362 682
rect 1022 678 1026 682
rect 1254 678 1258 682
rect 1430 678 1434 682
rect 1574 678 1578 682
rect 1606 678 1610 682
rect 1638 678 1642 682
rect 2270 678 2274 682
rect 6 668 10 672
rect 54 668 58 672
rect 78 668 82 672
rect 166 668 170 672
rect 174 668 178 672
rect 318 668 322 672
rect 422 668 426 672
rect 462 668 466 672
rect 486 668 490 672
rect 622 668 626 672
rect 630 668 634 672
rect 654 668 658 672
rect 726 668 730 672
rect 750 668 754 672
rect 774 668 778 672
rect 822 668 826 672
rect 958 668 962 672
rect 990 668 994 672
rect 1006 668 1010 672
rect 1022 668 1026 672
rect 1054 668 1058 672
rect 1062 668 1066 672
rect 1110 668 1114 672
rect 1118 668 1122 672
rect 1142 668 1146 672
rect 1174 668 1178 672
rect 1190 668 1194 672
rect 1198 668 1202 672
rect 1238 668 1242 672
rect 1262 668 1266 672
rect 86 658 90 662
rect 142 658 146 662
rect 158 658 162 662
rect 198 658 202 662
rect 214 658 218 662
rect 254 658 258 662
rect 270 658 274 662
rect 326 658 330 662
rect 350 658 354 662
rect 374 658 378 662
rect 414 658 418 662
rect 430 658 434 662
rect 534 659 538 663
rect 566 658 570 662
rect 646 658 650 662
rect 678 658 682 662
rect 686 658 690 662
rect 710 658 714 662
rect 734 658 738 662
rect 806 659 810 663
rect 1390 668 1394 672
rect 1470 668 1474 672
rect 1558 668 1562 672
rect 1590 668 1594 672
rect 1622 668 1626 672
rect 1670 668 1674 672
rect 1686 668 1690 672
rect 1734 668 1738 672
rect 1774 668 1778 672
rect 1854 668 1858 672
rect 1862 668 1866 672
rect 2014 668 2018 672
rect 2030 668 2034 672
rect 2062 668 2066 672
rect 2110 668 2114 672
rect 2254 668 2258 672
rect 878 658 882 662
rect 926 658 930 662
rect 934 658 938 662
rect 982 658 986 662
rect 990 658 994 662
rect 1030 658 1034 662
rect 1046 658 1050 662
rect 1070 658 1074 662
rect 1182 658 1186 662
rect 1206 658 1210 662
rect 1286 658 1290 662
rect 1326 658 1330 662
rect 1342 658 1346 662
rect 1406 658 1410 662
rect 1446 658 1450 662
rect 1478 658 1482 662
rect 1502 658 1506 662
rect 1510 658 1514 662
rect 1534 658 1538 662
rect 1550 658 1554 662
rect 1614 658 1618 662
rect 1662 658 1666 662
rect 1678 658 1682 662
rect 1726 658 1730 662
rect 1766 659 1770 663
rect 1886 658 1890 662
rect 1998 659 2002 663
rect 2038 658 2042 662
rect 2046 658 2050 662
rect 2086 658 2090 662
rect 2102 658 2106 662
rect 2174 658 2178 662
rect 2246 658 2250 662
rect 142 648 146 652
rect 214 648 218 652
rect 342 648 346 652
rect 398 648 402 652
rect 486 648 490 652
rect 606 648 610 652
rect 646 648 650 652
rect 758 648 762 652
rect 942 648 946 652
rect 958 648 962 652
rect 982 648 986 652
rect 1030 648 1034 652
rect 1086 648 1090 652
rect 1094 648 1098 652
rect 1142 648 1146 652
rect 1158 648 1162 652
rect 1222 648 1226 652
rect 1286 648 1290 652
rect 1438 648 1442 652
rect 1462 648 1466 652
rect 1494 648 1498 652
rect 1646 648 1650 652
rect 1710 648 1714 652
rect 1838 648 1842 652
rect 1878 648 1882 652
rect 2078 648 2082 652
rect 2086 648 2090 652
rect 30 638 34 642
rect 502 638 506 642
rect 670 638 674 642
rect 1310 638 1314 642
rect 1638 638 1642 642
rect 2134 638 2138 642
rect 134 618 138 622
rect 446 618 450 622
rect 470 618 474 622
rect 614 618 618 622
rect 702 618 706 622
rect 918 618 922 622
rect 1518 618 1522 622
rect 1606 618 1610 622
rect 1902 618 1906 622
rect 1934 618 1938 622
rect 2302 618 2306 622
rect 378 603 382 607
rect 385 603 389 607
rect 1394 603 1398 607
rect 1401 603 1405 607
rect 142 588 146 592
rect 270 588 274 592
rect 294 588 298 592
rect 318 588 322 592
rect 534 588 538 592
rect 710 588 714 592
rect 846 588 850 592
rect 910 588 914 592
rect 1038 588 1042 592
rect 1086 588 1090 592
rect 1110 588 1114 592
rect 1222 588 1226 592
rect 1318 588 1322 592
rect 1414 588 1418 592
rect 1430 588 1434 592
rect 1478 588 1482 592
rect 1606 588 1610 592
rect 1862 588 1866 592
rect 1982 588 1986 592
rect 1998 588 2002 592
rect 1806 578 1810 582
rect 126 568 130 572
rect 166 568 170 572
rect 446 568 450 572
rect 566 568 570 572
rect 1022 568 1026 572
rect 1070 568 1074 572
rect 1182 568 1186 572
rect 1214 568 1218 572
rect 1310 568 1314 572
rect 1654 568 1658 572
rect 150 558 154 562
rect 6 548 10 552
rect 30 548 34 552
rect 70 548 74 552
rect 166 548 170 552
rect 190 558 194 562
rect 302 558 306 562
rect 342 558 346 562
rect 206 548 210 552
rect 278 548 282 552
rect 318 548 322 552
rect 398 548 402 552
rect 454 548 458 552
rect 470 548 474 552
rect 486 558 490 562
rect 550 558 554 562
rect 582 558 586 562
rect 614 558 618 562
rect 766 558 770 562
rect 1030 558 1034 562
rect 1046 558 1050 562
rect 1094 558 1098 562
rect 1230 558 1234 562
rect 1238 558 1242 562
rect 1254 558 1258 562
rect 1294 558 1298 562
rect 1326 558 1330 562
rect 1342 558 1346 562
rect 1462 558 1466 562
rect 1494 558 1498 562
rect 1630 558 1634 562
rect 526 548 530 552
rect 534 548 538 552
rect 566 548 570 552
rect 598 548 602 552
rect 78 538 82 542
rect 134 538 138 542
rect 158 538 162 542
rect 646 547 650 551
rect 718 548 722 552
rect 774 548 778 552
rect 782 548 786 552
rect 806 548 810 552
rect 814 548 818 552
rect 830 548 834 552
rect 854 548 858 552
rect 886 548 890 552
rect 894 548 898 552
rect 918 548 922 552
rect 966 548 970 552
rect 1110 548 1114 552
rect 1126 548 1130 552
rect 1158 548 1162 552
rect 1166 548 1170 552
rect 1198 548 1202 552
rect 1222 548 1226 552
rect 1262 548 1266 552
rect 1302 548 1306 552
rect 1350 548 1354 552
rect 1358 548 1362 552
rect 1382 548 1386 552
rect 1478 548 1482 552
rect 1550 548 1554 552
rect 1910 558 1914 562
rect 1654 548 1658 552
rect 1670 548 1674 552
rect 1678 548 1682 552
rect 1702 548 1706 552
rect 214 538 218 542
rect 286 538 290 542
rect 310 538 314 542
rect 366 538 370 542
rect 454 538 458 542
rect 502 538 506 542
rect 526 538 530 542
rect 558 538 562 542
rect 590 538 594 542
rect 614 538 618 542
rect 662 538 666 542
rect 742 538 746 542
rect 942 538 946 542
rect 1046 538 1050 542
rect 1070 538 1074 542
rect 1118 538 1122 542
rect 1742 547 1746 551
rect 1774 548 1778 552
rect 1838 548 1842 552
rect 1846 548 1850 552
rect 1854 548 1858 552
rect 1894 548 1898 552
rect 2166 558 2170 562
rect 1950 548 1954 552
rect 1966 548 1970 552
rect 2014 548 2018 552
rect 2022 548 2026 552
rect 2046 548 2050 552
rect 2062 548 2066 552
rect 2070 548 2074 552
rect 2086 548 2090 552
rect 2110 548 2114 552
rect 2134 548 2138 552
rect 2150 548 2154 552
rect 2166 548 2170 552
rect 2222 548 2226 552
rect 2270 548 2274 552
rect 1254 538 1258 542
rect 1326 538 1330 542
rect 1446 538 1450 542
rect 1486 538 1490 542
rect 1510 538 1514 542
rect 1614 538 1618 542
rect 1662 538 1666 542
rect 1726 538 1730 542
rect 1822 538 1826 542
rect 1894 538 1898 542
rect 1942 538 1946 542
rect 1958 538 1962 542
rect 2142 538 2146 542
rect 2254 538 2258 542
rect 2294 538 2298 542
rect 510 528 514 532
rect 1078 528 1082 532
rect 1366 528 1370 532
rect 1422 528 1426 532
rect 1454 528 1458 532
rect 1542 528 1546 532
rect 1574 528 1578 532
rect 2006 528 2010 532
rect 2030 528 2034 532
rect 734 518 738 522
rect 758 518 762 522
rect 1278 518 1282 522
rect 1502 518 1506 522
rect 1606 518 1610 522
rect 1686 518 1690 522
rect 2118 518 2122 522
rect 2174 518 2178 522
rect 882 503 886 507
rect 889 503 893 507
rect 1914 503 1918 507
rect 1921 503 1925 507
rect 174 488 178 492
rect 342 488 346 492
rect 462 488 466 492
rect 742 488 746 492
rect 1094 488 1098 492
rect 1110 488 1114 492
rect 1222 488 1226 492
rect 1238 488 1242 492
rect 1382 488 1386 492
rect 1438 488 1442 492
rect 1462 488 1466 492
rect 1598 488 1602 492
rect 1790 488 1794 492
rect 1830 488 1834 492
rect 1862 488 1866 492
rect 2014 488 2018 492
rect 2158 488 2162 492
rect 2198 488 2202 492
rect 126 478 130 482
rect 302 478 306 482
rect 1102 478 1106 482
rect 1702 478 1706 482
rect 150 468 154 472
rect 158 468 162 472
rect 214 468 218 472
rect 278 468 282 472
rect 326 468 330 472
rect 334 468 338 472
rect 398 468 402 472
rect 470 468 474 472
rect 518 468 522 472
rect 646 468 650 472
rect 662 468 666 472
rect 774 468 778 472
rect 806 468 810 472
rect 902 468 906 472
rect 942 468 946 472
rect 950 468 954 472
rect 982 468 986 472
rect 998 468 1002 472
rect 1014 468 1018 472
rect 1198 468 1202 472
rect 1230 468 1234 472
rect 1254 468 1258 472
rect 1342 468 1346 472
rect 1358 468 1362 472
rect 1406 468 1410 472
rect 1430 468 1434 472
rect 1470 468 1474 472
rect 1478 468 1482 472
rect 1518 468 1522 472
rect 1542 468 1546 472
rect 1630 468 1634 472
rect 1662 468 1666 472
rect 1918 468 1922 472
rect 2046 468 2050 472
rect 2086 468 2090 472
rect 2134 468 2138 472
rect 2142 468 2146 472
rect 2166 468 2170 472
rect 2206 468 2210 472
rect 2254 468 2258 472
rect 38 458 42 462
rect 62 458 66 462
rect 102 458 106 462
rect 142 458 146 462
rect 222 458 226 462
rect 326 458 330 462
rect 406 458 410 462
rect 478 458 482 462
rect 486 458 490 462
rect 558 458 562 462
rect 590 459 594 463
rect 630 458 634 462
rect 638 458 642 462
rect 694 458 698 462
rect 710 458 714 462
rect 750 458 754 462
rect 766 458 770 462
rect 790 458 794 462
rect 878 458 882 462
rect 958 458 962 462
rect 1030 459 1034 463
rect 1126 458 1130 462
rect 1150 458 1154 462
rect 1158 458 1162 462
rect 1166 458 1170 462
rect 1174 458 1178 462
rect 1206 458 1210 462
rect 1318 458 1322 462
rect 1398 458 1402 462
rect 1486 458 1490 462
rect 1494 458 1498 462
rect 1534 459 1538 463
rect 1606 458 1610 462
rect 1638 458 1642 462
rect 1726 458 1730 462
rect 1742 458 1746 462
rect 1806 458 1810 462
rect 1814 458 1818 462
rect 1822 458 1826 462
rect 1846 458 1850 462
rect 1926 459 1930 463
rect 1966 458 1970 462
rect 2030 458 2034 462
rect 2046 458 2050 462
rect 2070 458 2074 462
rect 2078 458 2082 462
rect 2118 458 2122 462
rect 2126 458 2130 462
rect 2174 458 2178 462
rect 2190 458 2194 462
rect 2246 458 2250 462
rect 118 448 122 452
rect 174 448 178 452
rect 294 448 298 452
rect 350 448 354 452
rect 502 448 506 452
rect 622 448 626 452
rect 750 448 754 452
rect 814 448 818 452
rect 982 448 986 452
rect 1214 448 1218 452
rect 1230 448 1234 452
rect 1374 448 1378 452
rect 1454 448 1458 452
rect 1502 448 1506 452
rect 1662 448 1666 452
rect 2102 448 2106 452
rect 2158 448 2162 452
rect 2190 448 2194 452
rect 446 438 450 442
rect 1262 438 1266 442
rect 1142 428 1146 432
rect 526 418 530 422
rect 838 418 842 422
rect 1622 418 1626 422
rect 1990 418 1994 422
rect 378 403 382 407
rect 385 403 389 407
rect 1394 403 1398 407
rect 1401 403 1405 407
rect 142 388 146 392
rect 262 388 266 392
rect 294 388 298 392
rect 430 388 434 392
rect 566 388 570 392
rect 598 388 602 392
rect 694 388 698 392
rect 726 388 730 392
rect 854 388 858 392
rect 1094 388 1098 392
rect 1182 388 1186 392
rect 1230 388 1234 392
rect 1326 388 1330 392
rect 1534 388 1538 392
rect 1574 388 1578 392
rect 1686 388 1690 392
rect 1838 388 1842 392
rect 2054 388 2058 392
rect 398 368 402 372
rect 414 368 418 372
rect 766 368 770 372
rect 894 368 898 372
rect 1030 368 1034 372
rect 1422 368 1426 372
rect 1630 368 1634 372
rect 2198 368 2202 372
rect 6 358 10 362
rect 54 348 58 352
rect 78 358 82 362
rect 470 358 474 362
rect 126 348 130 352
rect 142 348 146 352
rect 190 348 194 352
rect 214 348 218 352
rect 278 348 282 352
rect 374 348 378 352
rect 606 358 610 362
rect 494 348 498 352
rect 510 348 514 352
rect 542 348 546 352
rect 574 348 578 352
rect 582 348 586 352
rect 622 348 626 352
rect 646 358 650 362
rect 678 348 682 352
rect 702 348 706 352
rect 710 348 714 352
rect 726 348 730 352
rect 782 348 786 352
rect 806 358 810 362
rect 1006 358 1010 362
rect 830 348 834 352
rect 862 348 866 352
rect 870 348 874 352
rect 1046 358 1050 362
rect 1134 358 1138 362
rect 38 338 42 342
rect 46 338 50 342
rect 150 338 154 342
rect 270 338 274 342
rect 302 338 306 342
rect 334 338 338 342
rect 446 338 450 342
rect 478 338 482 342
rect 502 338 506 342
rect 526 338 530 342
rect 590 338 594 342
rect 614 338 618 342
rect 958 347 962 351
rect 1038 348 1042 352
rect 1070 348 1074 352
rect 1078 348 1082 352
rect 1102 348 1106 352
rect 1198 358 1202 362
rect 1366 358 1370 362
rect 1158 348 1162 352
rect 1182 348 1186 352
rect 1198 348 1202 352
rect 1238 348 1242 352
rect 1246 348 1250 352
rect 1254 348 1258 352
rect 1262 348 1266 352
rect 1294 348 1298 352
rect 1302 348 1306 352
rect 1310 348 1314 352
rect 1334 348 1338 352
rect 1390 358 1394 362
rect 1622 358 1626 362
rect 1646 358 1650 362
rect 1678 358 1682 362
rect 1750 358 1754 362
rect 1390 348 1394 352
rect 1454 348 1458 352
rect 1478 348 1482 352
rect 1526 348 1530 352
rect 1542 348 1546 352
rect 1558 348 1562 352
rect 1590 348 1594 352
rect 1606 348 1610 352
rect 1734 348 1738 352
rect 1990 358 1994 362
rect 1774 348 1778 352
rect 1790 348 1794 352
rect 1798 348 1802 352
rect 1830 348 1834 352
rect 1910 348 1914 352
rect 1974 348 1978 352
rect 1982 348 1986 352
rect 2006 348 2010 352
rect 2030 358 2034 362
rect 2118 347 2122 351
rect 2158 348 2162 352
rect 2182 358 2186 362
rect 2246 348 2250 352
rect 2262 348 2266 352
rect 718 338 722 342
rect 750 338 754 342
rect 774 338 778 342
rect 822 338 826 342
rect 974 338 978 342
rect 990 338 994 342
rect 1038 338 1042 342
rect 1062 338 1066 342
rect 1110 338 1114 342
rect 1166 338 1170 342
rect 1174 338 1178 342
rect 1286 338 1290 342
rect 1350 338 1354 342
rect 1398 338 1402 342
rect 1502 338 1506 342
rect 1518 338 1522 342
rect 1550 338 1554 342
rect 1606 338 1610 342
rect 1630 338 1634 342
rect 1654 338 1658 342
rect 1710 338 1714 342
rect 1734 338 1738 342
rect 1782 338 1786 342
rect 1822 338 1826 342
rect 1918 338 1922 342
rect 1934 338 1938 342
rect 1966 338 1970 342
rect 1998 338 2002 342
rect 2046 338 2050 342
rect 2134 338 2138 342
rect 2150 338 2154 342
rect 2182 338 2186 342
rect 2198 338 2202 342
rect 30 328 34 332
rect 102 328 106 332
rect 318 328 322 332
rect 1678 328 1682 332
rect 1694 328 1698 332
rect 1846 328 1850 332
rect 6 318 10 322
rect 70 318 74 322
rect 246 318 250 322
rect 638 318 642 322
rect 798 318 802 322
rect 1054 318 1058 322
rect 1142 318 1146 322
rect 1614 318 1618 322
rect 1758 318 1762 322
rect 1854 318 1858 322
rect 2022 318 2026 322
rect 882 303 886 307
rect 889 303 893 307
rect 1914 303 1918 307
rect 1921 303 1925 307
rect 38 288 42 292
rect 134 288 138 292
rect 238 288 242 292
rect 270 288 274 292
rect 390 288 394 292
rect 686 288 690 292
rect 694 288 698 292
rect 862 288 866 292
rect 974 288 978 292
rect 998 288 1002 292
rect 1006 288 1010 292
rect 1150 288 1154 292
rect 1158 288 1162 292
rect 1254 288 1258 292
rect 1494 288 1498 292
rect 1678 288 1682 292
rect 1774 288 1778 292
rect 1990 288 1994 292
rect 2022 288 2026 292
rect 2094 288 2098 292
rect 2190 288 2194 292
rect 2214 288 2218 292
rect 230 278 234 282
rect 30 268 34 272
rect 118 268 122 272
rect 190 268 194 272
rect 214 268 218 272
rect 246 268 250 272
rect 294 268 298 272
rect 366 268 370 272
rect 470 268 474 272
rect 486 268 490 272
rect 502 268 506 272
rect 518 268 522 272
rect 542 268 546 272
rect 590 268 594 272
rect 606 268 610 272
rect 790 268 794 272
rect 806 268 810 272
rect 838 268 842 272
rect 918 268 922 272
rect 958 268 962 272
rect 974 268 978 272
rect 1022 268 1026 272
rect 1030 268 1034 272
rect 1070 268 1074 272
rect 1222 268 1226 272
rect 1270 268 1274 272
rect 1278 268 1282 272
rect 1342 268 1346 272
rect 1350 268 1354 272
rect 1438 268 1442 272
rect 1486 268 1490 272
rect 1590 268 1594 272
rect 1606 268 1610 272
rect 1622 268 1626 272
rect 1646 268 1650 272
rect 1670 268 1674 272
rect 1998 268 2002 272
rect 2038 268 2042 272
rect 2070 268 2074 272
rect 2134 268 2138 272
rect 2158 268 2162 272
rect 2206 268 2210 272
rect 22 258 26 262
rect 94 258 98 262
rect 174 258 178 262
rect 286 258 290 262
rect 302 258 306 262
rect 422 258 426 262
rect 454 259 458 263
rect 494 258 498 262
rect 574 258 578 262
rect 582 258 586 262
rect 638 258 642 262
rect 726 258 730 262
rect 758 259 762 263
rect 846 258 850 262
rect 894 258 898 262
rect 910 258 914 262
rect 1038 258 1042 262
rect 1046 258 1050 262
rect 1086 259 1090 263
rect 1118 258 1122 262
rect 1214 258 1218 262
rect 1478 258 1482 262
rect 1534 258 1538 262
rect 1550 258 1554 262
rect 1598 258 1602 262
rect 1630 258 1634 262
rect 1710 258 1714 262
rect 1726 258 1730 262
rect 1806 258 1810 262
rect 1814 258 1818 262
rect 1910 259 1914 263
rect 2006 258 2010 262
rect 2046 258 2050 262
rect 2150 258 2154 262
rect 2246 258 2250 262
rect 2270 258 2274 262
rect 6 248 10 252
rect 22 248 26 252
rect 262 248 266 252
rect 534 248 538 252
rect 558 248 562 252
rect 806 248 810 252
rect 974 248 978 252
rect 998 248 1002 252
rect 1054 248 1058 252
rect 1254 248 1258 252
rect 1454 248 1458 252
rect 1478 248 1482 252
rect 1614 248 1618 252
rect 1654 248 1658 252
rect 1982 248 1986 252
rect 2070 248 2074 252
rect 2190 248 2194 252
rect 54 238 58 242
rect 1974 238 1978 242
rect 1406 218 1410 222
rect 378 203 382 207
rect 385 203 389 207
rect 1394 203 1398 207
rect 1401 203 1405 207
rect 94 188 98 192
rect 238 188 242 192
rect 406 188 410 192
rect 558 188 562 192
rect 630 188 634 192
rect 782 188 786 192
rect 798 188 802 192
rect 814 188 818 192
rect 998 188 1002 192
rect 1094 188 1098 192
rect 1182 188 1186 192
rect 1278 188 1282 192
rect 1342 188 1346 192
rect 1462 188 1466 192
rect 1574 188 1578 192
rect 1870 188 1874 192
rect 2038 188 2042 192
rect 2286 188 2290 192
rect 982 168 986 172
rect 1678 168 1682 172
rect 1806 168 1810 172
rect 1934 168 1938 172
rect 126 158 130 162
rect 342 158 346 162
rect 30 147 34 151
rect 54 148 58 152
rect 110 148 114 152
rect 158 147 162 151
rect 190 148 194 152
rect 286 148 290 152
rect 302 148 306 152
rect 342 148 346 152
rect 374 148 378 152
rect 390 148 394 152
rect 422 148 426 152
rect 430 148 434 152
rect 438 148 442 152
rect 462 148 466 152
rect 518 148 522 152
rect 574 148 578 152
rect 598 158 602 162
rect 646 148 650 152
rect 670 158 674 162
rect 102 138 106 142
rect 126 138 130 142
rect 366 138 370 142
rect 718 147 722 151
rect 830 148 834 152
rect 854 158 858 162
rect 1110 158 1114 162
rect 926 148 930 152
rect 1038 148 1042 152
rect 1062 148 1066 152
rect 1102 148 1106 152
rect 1134 158 1138 162
rect 1158 148 1162 152
rect 1166 148 1170 152
rect 1190 148 1194 152
rect 1214 148 1218 152
rect 1238 158 1242 162
rect 1310 158 1314 162
rect 1382 158 1386 162
rect 1262 148 1266 152
rect 1326 148 1330 152
rect 1350 148 1354 152
rect 1358 148 1362 152
rect 1366 148 1370 152
rect 1694 158 1698 162
rect 1422 148 1426 152
rect 1438 148 1442 152
rect 1470 148 1474 152
rect 1478 148 1482 152
rect 1526 148 1530 152
rect 1614 148 1618 152
rect 2078 158 2082 162
rect 1726 148 1730 152
rect 1766 148 1770 152
rect 1870 148 1874 152
rect 1958 148 1962 152
rect 2014 148 2018 152
rect 2022 148 2026 152
rect 2102 148 2106 152
rect 2126 148 2130 152
rect 2150 158 2154 162
rect 2262 158 2266 162
rect 2286 148 2290 152
rect 478 138 482 142
rect 566 138 570 142
rect 614 138 618 142
rect 638 138 642 142
rect 670 138 674 142
rect 686 138 690 142
rect 726 138 730 142
rect 766 138 770 142
rect 790 138 794 142
rect 806 138 810 142
rect 822 138 826 142
rect 854 138 858 142
rect 886 138 890 142
rect 918 138 922 142
rect 1102 138 1106 142
rect 1150 138 1154 142
rect 1206 138 1210 142
rect 1254 138 1258 142
rect 1294 138 1298 142
rect 1430 138 1434 142
rect 1494 138 1498 142
rect 1606 138 1610 142
rect 1678 138 1682 142
rect 1694 138 1698 142
rect 1726 138 1730 142
rect 1742 138 1746 142
rect 1894 138 1898 142
rect 2062 138 2066 142
rect 2110 138 2114 142
rect 2166 138 2170 142
rect 2174 138 2178 142
rect 2246 138 2250 142
rect 2294 138 2298 142
rect 62 128 66 132
rect 190 128 194 132
rect 718 128 722 132
rect 990 128 994 132
rect 1854 128 1858 132
rect 1982 128 1986 132
rect 334 118 338 122
rect 590 118 594 122
rect 798 118 802 122
rect 814 118 818 122
rect 1230 118 1234 122
rect 1278 118 1282 122
rect 1302 118 1306 122
rect 1406 118 1410 122
rect 1822 118 1826 122
rect 1838 118 1842 122
rect 1886 118 1890 122
rect 2086 118 2090 122
rect 2142 118 2146 122
rect 2230 118 2234 122
rect 882 103 886 107
rect 889 103 893 107
rect 1914 103 1918 107
rect 1921 103 1925 107
rect 6 88 10 92
rect 118 88 122 92
rect 142 88 146 92
rect 182 88 186 92
rect 214 88 218 92
rect 390 88 394 92
rect 398 88 402 92
rect 494 88 498 92
rect 678 88 682 92
rect 774 88 778 92
rect 1054 88 1058 92
rect 1086 88 1090 92
rect 1190 88 1194 92
rect 1286 88 1290 92
rect 1326 88 1330 92
rect 1438 88 1442 92
rect 1646 88 1650 92
rect 1774 88 1778 92
rect 1830 88 1834 92
rect 1854 88 1858 92
rect 1958 88 1962 92
rect 2086 88 2090 92
rect 2094 88 2098 92
rect 2198 88 2202 92
rect 2214 88 2218 92
rect 646 78 650 82
rect 782 78 786 82
rect 1222 78 1226 82
rect 1710 78 1714 82
rect 1838 78 1842 82
rect 38 68 42 72
rect 54 68 58 72
rect 94 68 98 72
rect 150 68 154 72
rect 158 68 162 72
rect 222 68 226 72
rect 294 68 298 72
rect 310 68 314 72
rect 358 68 362 72
rect 430 68 434 72
rect 438 68 442 72
rect 462 68 466 72
rect 486 68 490 72
rect 694 68 698 72
rect 718 68 722 72
rect 798 68 802 72
rect 822 68 826 72
rect 862 68 866 72
rect 902 68 906 72
rect 934 68 938 72
rect 958 68 962 72
rect 1006 68 1010 72
rect 1094 68 1098 72
rect 1142 68 1146 72
rect 1238 68 1242 72
rect 1294 68 1298 72
rect 1318 68 1322 72
rect 1374 68 1378 72
rect 1494 68 1498 72
rect 1534 68 1538 72
rect 1558 68 1562 72
rect 1590 68 1594 72
rect 1614 68 1618 72
rect 1742 68 1746 72
rect 1814 68 1818 72
rect 1822 68 1826 72
rect 1846 68 1850 72
rect 1878 68 1882 72
rect 1902 78 1906 82
rect 1934 68 1938 72
rect 1974 78 1978 82
rect 2158 78 2162 82
rect 2174 68 2178 72
rect 2206 68 2210 72
rect 54 58 58 62
rect 62 58 66 62
rect 190 58 194 62
rect 350 58 354 62
rect 478 58 482 62
rect 526 58 530 62
rect 558 59 562 63
rect 622 58 626 62
rect 726 58 730 62
rect 814 58 818 62
rect 830 58 834 62
rect 846 58 850 62
rect 870 58 874 62
rect 902 58 906 62
rect 918 58 922 62
rect 990 59 994 63
rect 1142 58 1146 62
rect 1230 58 1234 62
rect 1310 58 1314 62
rect 1390 59 1394 63
rect 1502 59 1506 63
rect 1574 58 1578 62
rect 1582 58 1586 62
rect 1702 58 1706 62
rect 1862 58 1866 62
rect 1870 58 1874 62
rect 1926 58 1930 62
rect 1942 58 1946 62
rect 1990 58 1994 62
rect 2022 59 2026 63
rect 2054 58 2058 62
rect 2134 58 2138 62
rect 2246 58 2250 62
rect 2270 58 2274 62
rect 6 48 10 52
rect 38 48 42 52
rect 134 48 138 52
rect 414 48 418 52
rect 454 48 458 52
rect 782 48 786 52
rect 942 48 946 52
rect 1294 48 1298 52
rect 1550 48 1554 52
rect 1622 48 1626 52
rect 1790 48 1794 52
rect 1894 48 1898 52
rect 2190 48 2194 52
rect 1758 38 1762 42
rect 378 3 382 7
rect 385 3 389 7
rect 1394 3 1398 7
rect 1401 3 1405 7
<< metal2 >>
rect 1382 2128 1386 2132
rect 1870 2128 1874 2132
rect 880 2103 882 2107
rect 886 2103 889 2107
rect 893 2103 896 2107
rect 246 2072 249 2088
rect 318 2072 321 2078
rect 462 2072 465 2078
rect 606 2072 609 2088
rect 822 2072 825 2078
rect 838 2072 841 2088
rect 1382 2082 1385 2128
rect 1514 2088 1518 2091
rect 926 2072 929 2078
rect 1166 2072 1169 2078
rect 1206 2072 1209 2078
rect 1294 2072 1297 2078
rect 1366 2072 1369 2078
rect 1566 2072 1569 2088
rect 1846 2082 1849 2088
rect 1870 2082 1873 2128
rect 1912 2103 1914 2107
rect 1918 2103 1921 2107
rect 1925 2103 1928 2107
rect 1750 2072 1753 2078
rect 1886 2072 1889 2078
rect 570 2068 574 2071
rect 2058 2068 2062 2071
rect 6 2052 9 2068
rect 78 2052 81 2068
rect 142 2062 145 2068
rect 158 2062 161 2068
rect 10 1978 14 1981
rect 62 1942 65 2018
rect 182 1992 185 2058
rect 134 1972 137 1978
rect 198 1972 201 2018
rect 154 1968 158 1971
rect 218 1968 222 1971
rect 102 1962 105 1968
rect 70 1951 73 1958
rect 106 1948 110 1951
rect 62 1932 65 1938
rect 118 1922 121 1948
rect 126 1942 129 1958
rect 126 1872 129 1938
rect 134 1872 137 1968
rect 166 1962 169 1968
rect 230 1952 233 2038
rect 238 2012 241 2018
rect 154 1948 158 1951
rect 102 1862 105 1868
rect 150 1862 153 1948
rect 162 1938 166 1941
rect 158 1872 161 1938
rect 182 1922 185 1948
rect 190 1912 193 1938
rect 230 1902 233 1938
rect 198 1862 201 1878
rect 238 1862 241 2008
rect 246 1942 249 2068
rect 302 2062 305 2068
rect 282 2058 286 2061
rect 254 2042 257 2058
rect 294 2052 297 2058
rect 334 2052 337 2059
rect 270 2032 273 2038
rect 258 1968 262 1971
rect 282 1948 286 1951
rect 318 1942 321 1947
rect 266 1938 270 1941
rect 262 1872 265 1908
rect 270 1862 273 1918
rect 286 1912 289 1938
rect 278 1872 281 1878
rect 326 1872 329 1898
rect 334 1862 337 2038
rect 350 1952 353 2068
rect 446 2052 449 2058
rect 430 2042 433 2048
rect 394 2028 398 2031
rect 376 2003 378 2007
rect 382 2003 385 2007
rect 389 2003 392 2007
rect 378 1968 382 1971
rect 454 1942 457 1948
rect 414 1932 417 1938
rect 462 1922 465 2068
rect 486 2062 489 2068
rect 550 2052 553 2068
rect 546 2038 550 2041
rect 478 1972 481 2018
rect 498 1958 502 1961
rect 542 1952 545 2038
rect 558 1952 561 2058
rect 582 2042 585 2048
rect 566 1952 569 1968
rect 602 1958 606 1961
rect 622 1952 625 2018
rect 638 1972 641 2058
rect 514 1948 518 1951
rect 578 1948 582 1951
rect 590 1942 593 1948
rect 638 1942 641 1947
rect 506 1938 510 1941
rect 518 1938 526 1941
rect 578 1938 582 1941
rect 602 1938 606 1941
rect 50 1858 54 1861
rect 114 1858 118 1861
rect 62 1792 65 1858
rect 126 1852 129 1858
rect 106 1848 110 1851
rect 134 1842 137 1848
rect 98 1838 102 1841
rect 134 1782 137 1838
rect 6 1712 9 1738
rect 62 1722 65 1748
rect 110 1742 113 1748
rect 62 1662 65 1718
rect 78 1672 81 1718
rect 142 1692 145 1747
rect 222 1742 225 1858
rect 258 1838 262 1841
rect 254 1742 257 1748
rect 174 1712 177 1738
rect 102 1672 105 1678
rect 198 1672 201 1728
rect 114 1668 118 1671
rect 170 1668 174 1671
rect 194 1668 198 1671
rect 30 1621 33 1659
rect 178 1658 182 1661
rect 158 1652 161 1658
rect 130 1648 134 1651
rect 22 1618 33 1621
rect 90 1618 94 1621
rect 22 1592 25 1618
rect 6 1532 9 1558
rect 6 1181 9 1248
rect 14 1192 17 1568
rect 38 1552 41 1558
rect 54 1542 57 1618
rect 62 1552 65 1568
rect 102 1542 105 1548
rect 34 1538 38 1541
rect 82 1538 86 1541
rect 42 1528 46 1531
rect 54 1502 57 1538
rect 86 1482 89 1538
rect 94 1522 97 1538
rect 98 1488 102 1491
rect 38 1462 41 1468
rect 38 1342 41 1348
rect 46 1342 49 1468
rect 30 1272 33 1298
rect 46 1282 49 1338
rect 26 1258 30 1261
rect 22 1242 25 1248
rect 6 1178 17 1181
rect 6 1142 9 1148
rect 14 1092 17 1178
rect 30 1092 33 1258
rect 6 1052 9 1088
rect 26 1078 30 1081
rect 6 1042 9 1048
rect 14 991 17 1078
rect 38 1072 41 1218
rect 78 1152 81 1158
rect 86 1082 89 1478
rect 102 1472 105 1478
rect 110 1472 113 1618
rect 174 1572 177 1658
rect 230 1622 233 1718
rect 238 1662 241 1678
rect 254 1662 257 1738
rect 270 1732 273 1858
rect 294 1842 297 1848
rect 334 1802 337 1818
rect 350 1792 353 1838
rect 338 1788 342 1791
rect 358 1772 361 1828
rect 338 1758 342 1761
rect 358 1752 361 1768
rect 290 1748 294 1751
rect 346 1748 350 1751
rect 366 1742 369 1908
rect 462 1872 465 1918
rect 382 1862 385 1868
rect 402 1858 406 1861
rect 414 1822 417 1858
rect 376 1803 378 1807
rect 382 1803 385 1807
rect 389 1803 392 1807
rect 398 1791 401 1818
rect 398 1788 409 1791
rect 398 1752 401 1778
rect 406 1692 409 1788
rect 422 1752 425 1788
rect 430 1752 433 1818
rect 462 1742 465 1868
rect 474 1858 478 1861
rect 494 1852 497 1918
rect 518 1872 521 1938
rect 510 1802 513 1818
rect 518 1812 521 1868
rect 558 1862 561 1918
rect 582 1892 585 1928
rect 622 1922 625 1938
rect 578 1868 582 1871
rect 610 1868 614 1871
rect 538 1858 542 1861
rect 526 1832 529 1858
rect 550 1802 553 1848
rect 566 1832 569 1858
rect 482 1748 486 1751
rect 326 1682 329 1688
rect 254 1582 257 1658
rect 118 1552 121 1558
rect 150 1542 153 1547
rect 174 1541 177 1558
rect 182 1552 185 1578
rect 254 1552 257 1568
rect 278 1552 281 1668
rect 302 1642 305 1668
rect 350 1662 353 1668
rect 366 1652 369 1658
rect 322 1648 326 1651
rect 302 1562 305 1638
rect 326 1542 329 1578
rect 174 1538 185 1541
rect 118 1532 121 1538
rect 150 1472 153 1488
rect 122 1458 126 1461
rect 110 1442 113 1458
rect 134 1442 137 1448
rect 102 1342 105 1368
rect 118 1352 121 1358
rect 122 1338 126 1341
rect 102 1292 105 1338
rect 134 1322 137 1438
rect 146 1348 150 1351
rect 166 1342 169 1538
rect 182 1492 185 1538
rect 358 1532 361 1548
rect 210 1518 214 1521
rect 314 1518 318 1521
rect 198 1472 201 1518
rect 366 1502 369 1648
rect 376 1603 378 1607
rect 382 1603 385 1607
rect 389 1603 392 1607
rect 414 1552 417 1718
rect 422 1662 425 1678
rect 430 1662 433 1668
rect 462 1662 465 1738
rect 510 1711 513 1798
rect 574 1772 577 1868
rect 626 1858 630 1861
rect 586 1848 590 1851
rect 598 1832 601 1858
rect 526 1762 529 1768
rect 570 1758 574 1761
rect 554 1748 558 1751
rect 542 1742 545 1748
rect 534 1722 537 1738
rect 502 1708 513 1711
rect 502 1662 505 1708
rect 518 1672 521 1718
rect 582 1712 585 1748
rect 590 1742 593 1768
rect 606 1752 609 1848
rect 614 1802 617 1858
rect 646 1852 649 1858
rect 598 1742 601 1748
rect 538 1678 542 1681
rect 526 1662 529 1668
rect 566 1662 569 1708
rect 590 1672 593 1738
rect 578 1668 582 1671
rect 614 1662 617 1798
rect 622 1792 625 1848
rect 630 1752 633 1758
rect 622 1662 625 1688
rect 514 1658 518 1661
rect 422 1541 425 1608
rect 462 1572 465 1658
rect 478 1652 481 1658
rect 566 1652 569 1658
rect 546 1648 550 1651
rect 442 1568 446 1571
rect 442 1548 449 1551
rect 414 1538 425 1541
rect 434 1538 438 1541
rect 406 1512 409 1518
rect 230 1482 233 1488
rect 238 1482 241 1498
rect 206 1472 209 1478
rect 254 1471 257 1478
rect 366 1472 369 1478
rect 390 1472 393 1488
rect 254 1468 265 1471
rect 306 1468 310 1471
rect 338 1468 342 1471
rect 362 1468 366 1471
rect 178 1458 182 1461
rect 174 1442 177 1448
rect 182 1442 185 1448
rect 150 1312 153 1338
rect 134 1282 137 1288
rect 118 1272 121 1278
rect 182 1272 185 1328
rect 198 1282 201 1468
rect 210 1458 214 1461
rect 254 1452 257 1458
rect 262 1452 265 1468
rect 290 1458 294 1461
rect 226 1448 230 1451
rect 246 1392 249 1448
rect 278 1442 281 1458
rect 306 1448 310 1451
rect 290 1438 294 1441
rect 206 1352 209 1358
rect 262 1352 265 1388
rect 278 1362 281 1368
rect 270 1352 273 1358
rect 254 1342 257 1348
rect 214 1332 217 1338
rect 254 1332 257 1338
rect 242 1278 246 1281
rect 262 1281 265 1348
rect 294 1342 297 1348
rect 262 1278 273 1281
rect 194 1258 198 1261
rect 94 1252 97 1258
rect 262 1252 265 1268
rect 270 1262 273 1278
rect 310 1262 313 1378
rect 318 1362 321 1458
rect 326 1382 329 1458
rect 342 1372 345 1458
rect 398 1442 401 1458
rect 414 1452 417 1538
rect 422 1492 425 1528
rect 446 1492 449 1548
rect 462 1532 465 1558
rect 494 1552 497 1618
rect 534 1552 537 1588
rect 522 1548 526 1551
rect 478 1542 481 1548
rect 550 1542 553 1568
rect 462 1522 465 1528
rect 486 1481 489 1538
rect 574 1522 577 1658
rect 602 1648 606 1651
rect 614 1592 617 1658
rect 638 1632 641 1818
rect 654 1752 657 2028
rect 670 2022 673 2068
rect 682 2058 686 2061
rect 734 2012 737 2018
rect 742 2001 745 2018
rect 734 1998 745 2001
rect 734 1962 737 1998
rect 750 1992 753 2058
rect 774 2022 777 2058
rect 774 1972 777 2008
rect 806 1971 809 2059
rect 882 2058 886 2061
rect 806 1968 817 1971
rect 662 1892 665 1958
rect 710 1942 713 1948
rect 718 1942 721 1948
rect 726 1942 729 1948
rect 702 1882 705 1918
rect 662 1852 665 1878
rect 690 1868 694 1871
rect 714 1868 718 1871
rect 662 1782 665 1848
rect 662 1752 665 1758
rect 670 1751 673 1838
rect 678 1832 681 1858
rect 686 1792 689 1858
rect 694 1782 697 1798
rect 694 1752 697 1778
rect 702 1752 705 1758
rect 670 1748 678 1751
rect 686 1742 689 1748
rect 646 1662 649 1678
rect 662 1662 665 1668
rect 670 1662 673 1738
rect 682 1678 686 1681
rect 710 1672 713 1818
rect 726 1752 729 1868
rect 734 1862 737 1958
rect 790 1952 793 1958
rect 754 1948 758 1951
rect 806 1942 809 1958
rect 814 1952 817 1968
rect 822 1952 825 1988
rect 742 1912 745 1938
rect 798 1931 801 1938
rect 798 1928 809 1931
rect 742 1872 745 1908
rect 806 1902 809 1928
rect 806 1892 809 1898
rect 754 1858 758 1861
rect 766 1852 769 1858
rect 774 1842 777 1858
rect 822 1842 825 1948
rect 758 1792 761 1838
rect 822 1802 825 1838
rect 822 1752 825 1768
rect 734 1732 737 1748
rect 690 1658 694 1661
rect 702 1652 705 1658
rect 638 1592 641 1618
rect 614 1572 617 1578
rect 718 1572 721 1718
rect 766 1702 769 1718
rect 734 1662 737 1688
rect 766 1672 769 1698
rect 782 1672 785 1738
rect 830 1702 833 1938
rect 838 1882 841 2018
rect 846 1962 849 2058
rect 894 2042 897 2068
rect 946 2059 950 2062
rect 974 2062 977 2068
rect 1022 2062 1025 2068
rect 1050 2058 1054 2061
rect 902 2052 905 2058
rect 862 2032 865 2038
rect 878 1972 881 1978
rect 862 1962 865 1968
rect 850 1948 854 1951
rect 870 1942 873 1958
rect 858 1938 862 1941
rect 878 1922 881 1948
rect 880 1903 882 1907
rect 886 1903 889 1907
rect 893 1903 896 1907
rect 902 1872 905 1958
rect 910 1902 913 1958
rect 942 1942 945 1947
rect 918 1862 921 1868
rect 942 1862 945 1868
rect 958 1862 961 2008
rect 974 1952 977 2058
rect 1102 2042 1105 2048
rect 1110 2042 1113 2068
rect 1130 2058 1134 2061
rect 1002 2028 1006 2031
rect 998 1912 1001 2028
rect 1086 2012 1089 2038
rect 1058 1968 1062 1971
rect 1038 1962 1041 1968
rect 1022 1952 1025 1958
rect 1018 1938 1022 1941
rect 1038 1932 1041 1938
rect 1046 1932 1049 1938
rect 1054 1922 1057 1948
rect 1070 1922 1073 1958
rect 1086 1942 1089 2008
rect 1102 1942 1105 1947
rect 982 1862 985 1908
rect 1006 1902 1009 1918
rect 990 1862 993 1868
rect 838 1842 841 1859
rect 1010 1858 1014 1861
rect 870 1852 873 1858
rect 886 1832 889 1838
rect 862 1762 865 1768
rect 870 1742 873 1808
rect 886 1752 889 1768
rect 878 1742 881 1748
rect 894 1742 897 1858
rect 918 1842 921 1848
rect 934 1802 937 1858
rect 950 1842 953 1858
rect 978 1788 982 1791
rect 998 1782 1001 1858
rect 1018 1828 1022 1831
rect 922 1758 926 1761
rect 1010 1758 1017 1761
rect 934 1742 937 1748
rect 870 1722 873 1738
rect 880 1703 882 1707
rect 886 1703 889 1707
rect 893 1703 896 1707
rect 858 1688 862 1691
rect 750 1662 753 1668
rect 734 1652 737 1658
rect 758 1642 761 1658
rect 634 1568 638 1571
rect 650 1558 654 1561
rect 674 1558 678 1561
rect 582 1552 585 1558
rect 650 1548 654 1551
rect 686 1542 689 1568
rect 734 1552 737 1598
rect 710 1542 713 1548
rect 482 1478 489 1481
rect 478 1472 481 1478
rect 450 1468 454 1471
rect 474 1458 478 1461
rect 426 1448 430 1451
rect 438 1432 441 1458
rect 446 1452 449 1458
rect 458 1448 462 1451
rect 376 1403 378 1407
rect 382 1403 385 1407
rect 389 1403 392 1407
rect 398 1402 401 1418
rect 378 1378 382 1381
rect 330 1348 334 1351
rect 334 1272 337 1338
rect 342 1301 345 1368
rect 398 1362 401 1388
rect 430 1362 433 1378
rect 438 1362 441 1428
rect 466 1358 473 1361
rect 398 1352 401 1358
rect 410 1348 414 1351
rect 430 1342 433 1358
rect 450 1348 454 1351
rect 394 1338 398 1341
rect 458 1338 462 1341
rect 342 1298 353 1301
rect 318 1262 321 1268
rect 282 1258 286 1261
rect 242 1218 246 1221
rect 142 1182 145 1218
rect 138 1168 142 1171
rect 174 1162 177 1168
rect 162 1148 166 1151
rect 102 1111 105 1148
rect 150 1142 153 1148
rect 190 1142 193 1148
rect 102 1108 113 1111
rect 110 1072 113 1108
rect 42 1068 46 1071
rect 90 1068 94 1071
rect 30 1062 33 1068
rect 46 1052 49 1058
rect 82 1048 86 1051
rect 62 1012 65 1048
rect 94 1022 97 1058
rect 10 988 17 991
rect 14 962 17 988
rect 66 948 70 951
rect 102 942 105 958
rect 110 942 113 1068
rect 142 1032 145 1138
rect 150 1062 153 1068
rect 122 958 126 961
rect 130 948 134 951
rect 146 948 150 951
rect 158 942 161 1078
rect 166 952 169 958
rect 46 872 49 938
rect 86 932 89 938
rect 150 931 153 938
rect 146 928 153 931
rect 94 882 97 888
rect 50 858 54 861
rect 106 858 110 861
rect 46 752 49 768
rect 62 752 65 858
rect 106 848 110 851
rect 94 762 97 768
rect 102 742 105 838
rect 110 772 113 778
rect 54 672 57 738
rect 6 652 9 668
rect 34 638 38 641
rect 6 552 9 638
rect 70 552 73 568
rect 30 542 33 548
rect 78 542 81 668
rect 90 658 94 661
rect 102 651 105 738
rect 110 722 113 748
rect 94 648 105 651
rect 38 462 41 478
rect 62 422 65 458
rect 10 358 14 361
rect 86 361 89 548
rect 94 542 97 648
rect 102 462 105 468
rect 118 462 121 888
rect 126 872 129 908
rect 134 882 137 898
rect 126 712 129 858
rect 134 852 137 878
rect 142 852 145 858
rect 150 842 153 928
rect 158 852 161 938
rect 166 892 169 948
rect 174 892 177 1138
rect 198 1132 201 1138
rect 206 1132 209 1158
rect 230 1152 233 1178
rect 254 1161 257 1218
rect 270 1162 273 1258
rect 294 1222 297 1248
rect 310 1232 313 1258
rect 294 1172 297 1218
rect 254 1158 265 1161
rect 250 1148 254 1151
rect 262 1151 265 1158
rect 262 1148 270 1151
rect 226 1138 230 1141
rect 266 1138 270 1141
rect 254 1122 257 1138
rect 218 1118 222 1121
rect 230 1092 233 1118
rect 190 1072 193 1088
rect 198 1072 201 1078
rect 242 1068 246 1071
rect 254 1062 257 1068
rect 262 1062 265 1088
rect 218 1058 222 1061
rect 206 1052 209 1058
rect 230 1042 233 1048
rect 190 962 193 1038
rect 190 942 193 948
rect 166 872 169 878
rect 174 862 177 888
rect 134 722 137 758
rect 150 742 153 758
rect 158 742 161 848
rect 190 782 193 838
rect 166 752 169 768
rect 190 762 193 768
rect 134 682 137 688
rect 166 681 169 748
rect 182 742 185 748
rect 158 678 169 681
rect 158 662 161 678
rect 174 672 177 678
rect 138 658 142 661
rect 126 562 129 568
rect 134 542 137 618
rect 142 592 145 648
rect 158 561 161 658
rect 166 602 169 668
rect 198 662 201 1018
rect 206 942 209 968
rect 242 947 246 950
rect 218 868 222 871
rect 210 858 214 861
rect 238 852 241 858
rect 246 832 249 938
rect 262 922 265 1018
rect 270 901 273 1118
rect 278 1042 281 1048
rect 286 992 289 1148
rect 310 1132 313 1168
rect 350 1152 353 1298
rect 426 1288 430 1291
rect 446 1282 449 1338
rect 470 1322 473 1358
rect 494 1352 497 1418
rect 510 1382 513 1518
rect 518 1462 521 1518
rect 534 1462 537 1468
rect 542 1412 545 1498
rect 582 1472 585 1538
rect 638 1491 641 1538
rect 702 1502 705 1518
rect 734 1512 737 1548
rect 750 1542 753 1618
rect 766 1542 769 1668
rect 782 1582 785 1668
rect 910 1662 913 1668
rect 934 1662 937 1698
rect 942 1672 945 1738
rect 946 1668 950 1671
rect 958 1662 961 1758
rect 1006 1742 1009 1748
rect 1014 1742 1017 1758
rect 1038 1742 1041 1878
rect 1046 1862 1049 1898
rect 1054 1851 1057 1918
rect 1098 1878 1102 1881
rect 1110 1871 1113 2038
rect 1118 1982 1121 2058
rect 1158 2052 1161 2058
rect 1142 2042 1145 2048
rect 1142 2002 1145 2038
rect 1158 1932 1161 2048
rect 1166 1942 1169 2068
rect 1174 2062 1177 2068
rect 1202 2058 1206 2061
rect 1182 1942 1185 2058
rect 1214 2052 1217 2058
rect 1198 2042 1201 2048
rect 1230 2042 1233 2048
rect 1214 2032 1217 2038
rect 1246 2012 1249 2068
rect 1262 2063 1265 2068
rect 1430 2062 1433 2068
rect 1458 2058 1462 2061
rect 1322 2038 1326 2041
rect 1274 1968 1278 1971
rect 1214 1952 1217 1968
rect 1262 1962 1265 1968
rect 1274 1948 1278 1951
rect 1158 1912 1161 1928
rect 1170 1918 1177 1921
rect 1142 1892 1145 1908
rect 1102 1868 1113 1871
rect 1158 1872 1161 1878
rect 1046 1848 1057 1851
rect 1078 1852 1081 1858
rect 1046 1752 1049 1848
rect 1086 1822 1089 1858
rect 802 1659 806 1661
rect 798 1658 806 1659
rect 930 1658 934 1661
rect 830 1592 833 1638
rect 790 1552 793 1558
rect 854 1552 857 1558
rect 862 1552 865 1558
rect 842 1548 846 1551
rect 842 1538 846 1541
rect 798 1532 801 1538
rect 638 1488 646 1491
rect 646 1472 649 1488
rect 702 1472 705 1478
rect 510 1352 513 1368
rect 486 1342 489 1348
rect 362 1258 366 1261
rect 450 1258 454 1261
rect 462 1251 465 1318
rect 470 1262 473 1318
rect 478 1312 481 1338
rect 478 1292 481 1308
rect 478 1272 481 1278
rect 486 1272 489 1338
rect 474 1258 481 1261
rect 458 1248 465 1251
rect 376 1203 378 1207
rect 382 1203 385 1207
rect 389 1203 392 1207
rect 406 1172 409 1178
rect 374 1162 377 1168
rect 358 1152 361 1158
rect 410 1148 414 1151
rect 402 1138 406 1141
rect 326 1132 329 1138
rect 350 1132 353 1138
rect 294 1092 297 1098
rect 314 1078 318 1081
rect 318 1062 321 1068
rect 374 1063 377 1118
rect 422 1082 425 1158
rect 430 1122 433 1148
rect 438 1071 441 1218
rect 446 1192 449 1248
rect 462 1142 465 1178
rect 470 1152 473 1228
rect 478 1112 481 1258
rect 486 1182 489 1268
rect 494 1232 497 1348
rect 510 1302 513 1348
rect 534 1282 537 1288
rect 486 1122 489 1158
rect 494 1131 497 1218
rect 502 1182 505 1268
rect 510 1251 513 1268
rect 542 1262 545 1408
rect 574 1352 577 1468
rect 694 1462 697 1468
rect 750 1462 753 1528
rect 870 1522 873 1658
rect 894 1562 897 1658
rect 918 1642 921 1648
rect 950 1612 953 1658
rect 974 1652 977 1658
rect 982 1642 985 1658
rect 974 1592 977 1618
rect 990 1582 993 1738
rect 1014 1732 1017 1738
rect 1038 1732 1041 1738
rect 1022 1712 1025 1718
rect 1002 1668 1006 1671
rect 1002 1658 1006 1661
rect 1014 1658 1022 1661
rect 958 1562 961 1568
rect 982 1562 985 1578
rect 998 1572 1001 1618
rect 1006 1562 1009 1618
rect 1014 1602 1017 1658
rect 1022 1642 1025 1648
rect 1030 1602 1033 1718
rect 1038 1672 1041 1728
rect 1046 1702 1049 1748
rect 1062 1692 1065 1758
rect 1046 1662 1049 1668
rect 930 1548 934 1551
rect 1010 1548 1014 1551
rect 982 1542 985 1548
rect 1022 1542 1025 1548
rect 1030 1542 1033 1598
rect 1038 1562 1041 1568
rect 894 1532 897 1538
rect 998 1532 1001 1538
rect 1054 1532 1057 1538
rect 846 1492 849 1518
rect 880 1503 882 1507
rect 886 1503 889 1507
rect 893 1503 896 1507
rect 910 1492 913 1518
rect 810 1478 814 1481
rect 774 1472 777 1478
rect 782 1462 785 1468
rect 790 1462 793 1468
rect 594 1458 598 1461
rect 666 1458 670 1461
rect 642 1438 646 1441
rect 654 1432 657 1458
rect 726 1448 734 1451
rect 678 1442 681 1448
rect 718 1362 721 1418
rect 726 1392 729 1448
rect 742 1442 745 1458
rect 618 1358 622 1361
rect 730 1358 734 1361
rect 630 1352 633 1358
rect 750 1352 753 1428
rect 682 1348 686 1351
rect 730 1348 734 1351
rect 550 1292 553 1348
rect 574 1342 577 1348
rect 646 1342 649 1348
rect 750 1342 753 1348
rect 758 1342 761 1418
rect 766 1362 769 1398
rect 790 1362 793 1398
rect 806 1372 809 1458
rect 822 1422 825 1468
rect 870 1462 873 1468
rect 858 1458 862 1461
rect 910 1452 913 1458
rect 934 1452 937 1458
rect 842 1448 846 1451
rect 838 1432 841 1438
rect 810 1368 814 1371
rect 850 1358 854 1361
rect 802 1348 806 1351
rect 842 1348 846 1351
rect 782 1342 785 1348
rect 830 1342 833 1348
rect 898 1348 902 1351
rect 602 1318 606 1321
rect 566 1282 569 1318
rect 614 1312 617 1338
rect 798 1332 801 1338
rect 822 1332 825 1338
rect 730 1318 734 1321
rect 634 1278 638 1281
rect 634 1268 638 1271
rect 522 1258 526 1261
rect 594 1258 598 1261
rect 542 1252 545 1258
rect 510 1248 521 1251
rect 510 1152 513 1158
rect 502 1142 505 1148
rect 518 1142 521 1248
rect 494 1128 505 1131
rect 430 1068 441 1071
rect 406 1062 409 1068
rect 374 1058 377 1059
rect 334 982 337 1018
rect 298 968 302 971
rect 330 968 334 971
rect 302 942 305 968
rect 342 962 345 1008
rect 376 1003 378 1007
rect 382 1003 385 1007
rect 389 1003 392 1007
rect 346 958 350 961
rect 322 938 326 941
rect 322 928 326 931
rect 310 902 313 928
rect 270 898 281 901
rect 262 872 265 878
rect 270 862 273 878
rect 258 858 262 861
rect 258 848 262 851
rect 270 842 273 848
rect 278 842 281 898
rect 286 852 289 888
rect 302 832 305 868
rect 322 859 326 862
rect 206 742 209 788
rect 214 772 217 818
rect 242 748 246 751
rect 214 662 217 668
rect 254 662 257 768
rect 270 752 273 828
rect 350 792 353 928
rect 378 888 382 891
rect 390 852 393 948
rect 398 882 401 1008
rect 406 962 409 968
rect 414 942 417 948
rect 406 872 409 918
rect 414 892 417 928
rect 430 892 433 1068
rect 442 1058 446 1061
rect 466 1018 470 1021
rect 438 1002 441 1018
rect 438 952 441 988
rect 446 951 449 978
rect 458 958 481 961
rect 478 952 481 958
rect 446 948 454 951
rect 438 902 441 948
rect 470 942 473 948
rect 462 912 465 938
rect 422 872 425 878
rect 486 872 489 1068
rect 502 1042 505 1128
rect 518 1102 521 1138
rect 530 1118 534 1121
rect 542 1101 545 1248
rect 534 1098 545 1101
rect 526 1062 529 1068
rect 502 972 505 1038
rect 526 972 529 998
rect 518 962 521 968
rect 494 922 497 958
rect 518 912 521 918
rect 522 888 526 891
rect 534 882 537 1098
rect 542 962 545 968
rect 558 952 561 1258
rect 590 1182 593 1218
rect 614 1172 617 1238
rect 570 1148 574 1151
rect 566 1092 569 1098
rect 574 1082 577 1118
rect 590 1092 593 1168
rect 606 1102 609 1138
rect 622 1132 625 1138
rect 590 1072 593 1088
rect 610 1068 614 1071
rect 630 1062 633 1248
rect 646 1152 649 1218
rect 662 1151 665 1298
rect 742 1282 745 1288
rect 750 1282 753 1318
rect 766 1302 769 1318
rect 762 1278 766 1281
rect 774 1272 777 1278
rect 782 1272 785 1328
rect 878 1321 881 1338
rect 870 1318 881 1321
rect 790 1262 793 1318
rect 870 1272 873 1318
rect 880 1303 882 1307
rect 886 1303 889 1307
rect 893 1303 896 1307
rect 810 1268 814 1271
rect 694 1192 697 1258
rect 658 1148 665 1151
rect 690 1148 694 1151
rect 638 1132 641 1138
rect 686 1132 689 1138
rect 646 1122 649 1128
rect 670 1122 673 1128
rect 654 1072 657 1098
rect 630 1052 633 1058
rect 610 1048 614 1051
rect 574 962 577 968
rect 542 942 545 948
rect 550 932 553 938
rect 422 822 425 848
rect 438 832 441 868
rect 466 858 470 861
rect 376 803 378 807
rect 382 803 385 807
rect 389 803 392 807
rect 446 792 449 818
rect 306 788 310 791
rect 314 748 318 751
rect 338 748 342 751
rect 166 572 169 578
rect 154 558 161 561
rect 150 552 153 558
rect 162 548 166 551
rect 154 538 158 541
rect 126 482 129 488
rect 150 472 153 508
rect 174 492 177 648
rect 190 562 193 568
rect 190 552 193 558
rect 198 532 201 658
rect 210 648 214 651
rect 206 552 209 558
rect 206 542 209 548
rect 214 502 217 538
rect 158 472 161 478
rect 142 462 145 468
rect 138 458 142 461
rect 118 452 121 458
rect 170 448 174 451
rect 142 392 145 438
rect 214 422 217 468
rect 222 462 225 478
rect 82 358 89 361
rect 6 252 9 318
rect 22 262 25 358
rect 78 352 81 358
rect 58 348 62 351
rect 130 348 134 351
rect 38 342 41 348
rect 142 342 145 348
rect 30 291 33 328
rect 30 288 38 291
rect 46 272 49 338
rect 70 312 73 318
rect 102 292 105 328
rect 150 322 153 338
rect 130 288 134 291
rect 118 272 121 278
rect 34 268 38 271
rect 26 258 30 261
rect 22 242 25 248
rect 30 92 33 147
rect 46 112 49 268
rect 174 262 177 308
rect 94 252 97 258
rect 54 152 57 238
rect 98 188 102 191
rect 110 152 113 168
rect 122 158 126 161
rect 102 132 105 138
rect 10 88 14 91
rect 46 72 49 108
rect 62 81 65 128
rect 54 78 65 81
rect 54 72 57 78
rect 42 68 46 71
rect 62 62 65 68
rect 50 58 54 61
rect 6 52 9 58
rect 42 48 46 51
rect 94 -19 97 68
rect 110 52 113 148
rect 126 142 129 148
rect 142 92 145 158
rect 158 142 161 147
rect 182 92 185 358
rect 214 352 217 418
rect 262 392 265 748
rect 270 662 273 748
rect 306 738 310 741
rect 314 688 318 691
rect 314 668 318 671
rect 326 662 329 738
rect 358 732 361 778
rect 462 762 465 788
rect 366 732 369 758
rect 422 752 425 758
rect 478 752 481 838
rect 494 762 497 778
rect 502 752 505 758
rect 386 738 390 741
rect 358 692 361 728
rect 386 718 390 721
rect 398 692 401 728
rect 406 722 409 748
rect 430 742 433 748
rect 446 742 449 748
rect 418 738 422 741
rect 510 741 513 768
rect 502 738 513 741
rect 526 742 529 868
rect 534 862 537 878
rect 542 852 545 858
rect 538 758 542 761
rect 438 732 441 738
rect 414 718 422 721
rect 362 678 366 681
rect 350 662 353 668
rect 414 662 417 718
rect 458 668 462 671
rect 270 592 273 658
rect 294 592 297 628
rect 318 592 321 658
rect 342 582 345 648
rect 374 642 377 658
rect 398 632 401 648
rect 376 603 378 607
rect 382 603 385 607
rect 389 603 392 607
rect 274 548 278 551
rect 282 538 286 541
rect 278 461 281 468
rect 274 458 281 461
rect 286 352 289 528
rect 294 462 297 568
rect 302 562 305 568
rect 302 482 305 488
rect 294 452 297 458
rect 294 392 297 418
rect 282 348 286 351
rect 190 332 193 348
rect 214 282 217 348
rect 266 338 270 341
rect 298 338 302 341
rect 238 292 241 338
rect 214 272 217 278
rect 190 152 193 268
rect 214 132 217 158
rect 122 88 126 91
rect 150 72 153 78
rect 138 48 142 51
rect 110 -19 114 -18
rect 94 -22 114 -19
rect 158 -19 161 68
rect 182 61 185 88
rect 190 72 193 128
rect 214 92 217 128
rect 222 72 225 198
rect 230 192 233 278
rect 238 192 241 278
rect 246 272 249 318
rect 270 292 273 328
rect 294 322 297 338
rect 286 262 289 308
rect 310 282 313 538
rect 318 532 321 548
rect 326 512 329 538
rect 326 472 329 508
rect 342 492 345 558
rect 334 462 337 468
rect 322 458 326 461
rect 350 452 353 568
rect 402 548 406 551
rect 366 542 369 548
rect 414 532 417 658
rect 422 652 425 668
rect 470 662 473 738
rect 486 672 489 738
rect 430 642 433 658
rect 494 651 497 718
rect 502 692 505 738
rect 526 702 529 738
rect 534 663 537 718
rect 490 648 497 651
rect 430 592 433 638
rect 470 622 473 628
rect 446 602 449 618
rect 502 572 505 638
rect 534 592 537 648
rect 550 582 553 918
rect 558 891 561 948
rect 574 932 577 938
rect 558 888 569 891
rect 558 852 561 878
rect 558 752 561 848
rect 566 842 569 888
rect 574 872 577 888
rect 590 871 593 1038
rect 606 902 609 1038
rect 618 948 622 951
rect 590 868 598 871
rect 606 862 609 898
rect 630 892 633 1048
rect 638 1022 641 1068
rect 638 972 641 1018
rect 654 972 657 1068
rect 674 1058 678 1061
rect 686 1032 689 1128
rect 686 1022 689 1028
rect 694 982 697 1108
rect 702 1072 705 1258
rect 790 1252 793 1258
rect 818 1248 822 1251
rect 742 1172 745 1218
rect 718 1162 721 1168
rect 734 1072 737 1148
rect 750 1142 753 1238
rect 814 1192 817 1238
rect 830 1202 833 1268
rect 862 1263 865 1268
rect 862 1258 865 1259
rect 830 1162 833 1168
rect 790 1152 793 1158
rect 778 1148 782 1151
rect 742 1122 745 1138
rect 742 1062 745 1108
rect 746 1058 753 1061
rect 734 1042 737 1048
rect 750 1012 753 1058
rect 758 1042 761 1148
rect 782 1132 785 1138
rect 798 1132 801 1158
rect 870 1152 873 1268
rect 810 1138 817 1141
rect 770 1128 774 1131
rect 774 1072 777 1118
rect 806 1072 809 1118
rect 814 1072 817 1138
rect 782 1062 785 1068
rect 814 1062 817 1068
rect 838 1062 841 1068
rect 854 1062 857 1078
rect 870 1071 873 1148
rect 890 1147 894 1150
rect 880 1103 882 1107
rect 886 1103 889 1107
rect 893 1103 896 1107
rect 870 1068 878 1071
rect 742 992 745 1008
rect 750 991 753 1008
rect 758 1002 761 1038
rect 750 988 761 991
rect 638 932 641 948
rect 678 942 681 968
rect 694 962 697 978
rect 718 952 721 978
rect 694 942 697 948
rect 726 942 729 968
rect 758 952 761 988
rect 766 942 769 1018
rect 774 972 777 988
rect 774 952 777 968
rect 790 962 793 1058
rect 830 1042 833 1048
rect 798 992 801 1038
rect 862 1022 865 1068
rect 786 948 790 951
rect 806 942 809 958
rect 654 881 657 928
rect 694 892 697 928
rect 650 878 657 881
rect 630 872 633 878
rect 650 868 654 871
rect 678 862 681 868
rect 626 858 630 861
rect 642 858 646 861
rect 666 858 670 861
rect 578 758 582 761
rect 590 742 593 818
rect 598 782 601 838
rect 618 818 622 821
rect 598 752 601 778
rect 614 762 617 768
rect 558 732 561 738
rect 558 712 561 728
rect 582 692 585 738
rect 594 688 598 691
rect 562 658 566 661
rect 606 652 609 758
rect 622 752 625 758
rect 638 752 641 818
rect 662 792 665 858
rect 670 848 678 851
rect 662 752 665 758
rect 614 742 617 748
rect 658 738 662 741
rect 622 702 625 718
rect 450 568 454 571
rect 318 292 321 328
rect 334 272 337 338
rect 366 272 369 498
rect 376 403 378 407
rect 382 403 385 407
rect 389 403 392 407
rect 398 372 401 468
rect 410 458 414 461
rect 430 392 433 568
rect 490 558 494 561
rect 454 552 457 558
rect 466 548 470 551
rect 502 542 505 568
rect 534 552 537 568
rect 550 562 553 578
rect 566 572 569 578
rect 582 562 585 628
rect 522 548 526 551
rect 562 548 566 551
rect 590 542 593 598
rect 598 552 601 558
rect 606 551 609 648
rect 622 642 625 668
rect 630 652 633 668
rect 638 651 641 698
rect 646 682 649 738
rect 670 692 673 848
rect 686 762 689 888
rect 750 832 753 868
rect 758 852 761 928
rect 798 912 801 918
rect 766 852 769 858
rect 686 752 689 758
rect 694 752 697 818
rect 742 752 745 758
rect 750 742 753 748
rect 758 742 761 848
rect 774 842 777 908
rect 794 888 798 891
rect 682 738 686 741
rect 646 662 649 668
rect 638 648 646 651
rect 614 562 617 618
rect 654 572 657 668
rect 678 662 681 718
rect 686 662 689 688
rect 710 662 713 718
rect 726 672 729 728
rect 602 548 609 551
rect 614 542 617 548
rect 646 542 649 547
rect 662 542 665 658
rect 670 642 673 648
rect 702 612 705 618
rect 710 592 713 638
rect 726 602 729 668
rect 750 662 753 668
rect 734 652 737 658
rect 754 648 758 651
rect 766 632 769 818
rect 774 672 777 678
rect 790 602 793 818
rect 806 752 809 938
rect 830 862 833 878
rect 822 772 825 858
rect 822 762 825 768
rect 830 752 833 858
rect 838 762 841 968
rect 854 952 857 958
rect 878 942 881 1068
rect 894 942 897 948
rect 854 882 857 938
rect 880 903 882 907
rect 886 903 889 907
rect 893 903 896 907
rect 902 872 905 988
rect 910 972 913 1418
rect 918 1242 921 1438
rect 926 1432 929 1448
rect 942 1442 945 1528
rect 966 1492 969 1498
rect 1006 1492 1009 1528
rect 1046 1492 1049 1518
rect 1062 1492 1065 1508
rect 1030 1472 1033 1478
rect 1070 1472 1073 1778
rect 1086 1752 1089 1778
rect 1102 1752 1105 1868
rect 1118 1792 1121 1858
rect 1166 1802 1169 1858
rect 1158 1762 1161 1768
rect 1130 1758 1134 1761
rect 1146 1758 1150 1761
rect 1102 1742 1105 1748
rect 1082 1738 1089 1741
rect 1086 1663 1089 1738
rect 1086 1658 1089 1659
rect 1094 1622 1097 1738
rect 1110 1702 1113 1748
rect 1126 1742 1129 1748
rect 1134 1712 1137 1738
rect 1142 1732 1145 1748
rect 1174 1732 1177 1918
rect 1182 1902 1185 1938
rect 1190 1862 1193 1868
rect 1182 1852 1185 1858
rect 1190 1742 1193 1747
rect 1198 1742 1201 1928
rect 1206 1862 1209 1948
rect 1270 1932 1273 1938
rect 1214 1872 1217 1898
rect 1270 1872 1273 1928
rect 1286 1882 1289 2008
rect 1302 1962 1305 1968
rect 1086 1542 1089 1558
rect 1094 1552 1097 1558
rect 1110 1542 1113 1698
rect 1154 1688 1158 1691
rect 1118 1552 1121 1658
rect 1118 1542 1121 1548
rect 1134 1492 1137 1678
rect 1190 1662 1193 1728
rect 1154 1658 1158 1661
rect 1142 1492 1145 1658
rect 1166 1652 1169 1658
rect 1166 1542 1169 1548
rect 1190 1542 1193 1548
rect 1198 1542 1201 1738
rect 1206 1712 1209 1858
rect 1214 1652 1217 1868
rect 1266 1858 1270 1861
rect 1222 1842 1225 1848
rect 1250 1768 1254 1771
rect 1302 1761 1305 1958
rect 1318 1912 1321 1948
rect 1326 1892 1329 1938
rect 1318 1841 1321 1868
rect 1294 1758 1305 1761
rect 1310 1838 1321 1841
rect 1310 1762 1313 1838
rect 1294 1752 1297 1758
rect 1302 1742 1305 1748
rect 1278 1672 1281 1718
rect 1238 1662 1241 1668
rect 1286 1662 1289 1698
rect 1294 1662 1297 1668
rect 1302 1662 1305 1688
rect 1310 1682 1313 1758
rect 1334 1752 1337 2038
rect 1390 2022 1393 2028
rect 1394 2018 1398 2021
rect 1342 1982 1345 2018
rect 1392 2003 1394 2007
rect 1398 2003 1401 2007
rect 1405 2003 1408 2007
rect 1342 1952 1345 1978
rect 1350 1862 1353 1998
rect 1410 1968 1414 1971
rect 1358 1962 1361 1968
rect 1374 1862 1377 1968
rect 1386 1958 1390 1961
rect 1470 1952 1473 1958
rect 1386 1948 1390 1951
rect 1390 1932 1393 1938
rect 1390 1891 1393 1928
rect 1382 1888 1393 1891
rect 1342 1741 1345 1848
rect 1334 1738 1345 1741
rect 1318 1732 1321 1738
rect 1246 1652 1249 1658
rect 1262 1652 1265 1658
rect 1154 1518 1158 1521
rect 1206 1492 1209 1558
rect 1214 1552 1217 1558
rect 1230 1552 1233 1618
rect 1238 1602 1241 1648
rect 1318 1642 1321 1648
rect 1142 1482 1145 1488
rect 962 1468 966 1471
rect 994 1458 1001 1461
rect 998 1452 1001 1458
rect 926 1402 929 1428
rect 934 1392 937 1418
rect 942 1392 945 1438
rect 990 1432 993 1448
rect 998 1432 1001 1438
rect 990 1421 993 1428
rect 990 1418 1001 1421
rect 942 1372 945 1388
rect 942 1292 945 1358
rect 966 1342 969 1348
rect 950 1312 953 1338
rect 974 1332 977 1418
rect 998 1392 1001 1418
rect 986 1348 990 1351
rect 970 1328 974 1331
rect 950 1252 953 1308
rect 958 1251 961 1318
rect 990 1282 993 1288
rect 986 1268 990 1271
rect 966 1252 969 1268
rect 1006 1262 1009 1418
rect 1014 1372 1017 1458
rect 1022 1452 1025 1458
rect 1030 1442 1033 1468
rect 1042 1458 1046 1461
rect 1094 1452 1097 1458
rect 1038 1372 1041 1428
rect 1022 1352 1025 1358
rect 1030 1352 1033 1358
rect 1046 1352 1049 1448
rect 1054 1422 1057 1438
rect 1054 1372 1057 1418
rect 1054 1352 1057 1358
rect 1062 1352 1065 1358
rect 1014 1342 1017 1348
rect 1014 1262 1017 1268
rect 958 1248 966 1251
rect 926 1202 929 1218
rect 974 1212 977 1258
rect 1022 1252 1025 1348
rect 1030 1272 1033 1348
rect 1038 1262 1041 1268
rect 926 1142 929 1158
rect 958 1132 961 1158
rect 966 1142 969 1148
rect 982 1132 985 1148
rect 998 1142 1001 1248
rect 1006 1242 1009 1248
rect 1038 1242 1041 1248
rect 1046 1242 1049 1318
rect 1054 1252 1057 1348
rect 1086 1342 1089 1348
rect 1062 1272 1065 1278
rect 1070 1262 1073 1328
rect 1034 1238 1038 1241
rect 1014 1182 1017 1218
rect 1022 1172 1025 1198
rect 1038 1162 1041 1168
rect 1046 1162 1049 1218
rect 1018 1158 1022 1161
rect 1054 1152 1057 1158
rect 1034 1148 1038 1151
rect 1042 1138 1049 1141
rect 942 1072 945 1078
rect 918 1052 921 1058
rect 942 972 945 1028
rect 950 992 953 1018
rect 958 982 961 1128
rect 990 1112 993 1138
rect 1010 1118 1014 1121
rect 978 1088 982 1091
rect 990 1082 993 1108
rect 1030 1072 1033 1088
rect 982 1062 985 1068
rect 994 1058 998 1061
rect 994 1048 998 1051
rect 1018 1048 1022 1051
rect 974 992 977 998
rect 1006 972 1009 1018
rect 1046 992 1049 1138
rect 1054 1102 1057 1148
rect 1070 1131 1073 1258
rect 1078 1212 1081 1318
rect 1094 1282 1097 1438
rect 1086 1272 1089 1278
rect 1094 1272 1097 1278
rect 1086 1222 1089 1258
rect 1102 1242 1105 1478
rect 1174 1472 1177 1478
rect 1182 1472 1185 1478
rect 1230 1472 1233 1518
rect 1238 1492 1241 1598
rect 1250 1518 1254 1521
rect 1262 1472 1265 1518
rect 1186 1468 1190 1471
rect 1270 1471 1273 1608
rect 1278 1561 1281 1618
rect 1294 1592 1297 1628
rect 1326 1622 1329 1738
rect 1334 1662 1337 1738
rect 1350 1702 1353 1718
rect 1358 1672 1361 1818
rect 1366 1752 1369 1778
rect 1382 1752 1385 1888
rect 1406 1872 1409 1878
rect 1414 1862 1417 1908
rect 1438 1872 1441 1908
rect 1470 1872 1473 1898
rect 1478 1862 1481 1948
rect 1494 1942 1497 2038
rect 1518 1962 1521 2068
rect 1534 2062 1537 2068
rect 1526 2052 1529 2058
rect 1518 1952 1521 1958
rect 1494 1882 1497 1938
rect 1494 1862 1497 1868
rect 1510 1862 1513 1918
rect 1526 1882 1529 1888
rect 1526 1863 1529 1868
rect 1394 1858 1398 1861
rect 1526 1858 1529 1859
rect 1392 1803 1394 1807
rect 1398 1803 1401 1807
rect 1405 1803 1408 1807
rect 1414 1762 1417 1818
rect 1430 1792 1433 1838
rect 1446 1792 1449 1858
rect 1470 1852 1473 1858
rect 1458 1848 1462 1851
rect 1490 1848 1494 1851
rect 1462 1842 1465 1848
rect 1430 1782 1433 1788
rect 1422 1752 1425 1758
rect 1478 1752 1481 1758
rect 1278 1558 1286 1561
rect 1282 1548 1286 1551
rect 1302 1542 1305 1548
rect 1318 1542 1321 1558
rect 1342 1542 1345 1658
rect 1358 1652 1361 1658
rect 1374 1652 1377 1748
rect 1382 1742 1385 1748
rect 1390 1742 1393 1748
rect 1462 1682 1465 1748
rect 1510 1721 1513 1858
rect 1550 1812 1553 2048
rect 1566 2012 1569 2068
rect 1686 2062 1689 2068
rect 1574 2002 1577 2058
rect 1670 2042 1673 2059
rect 1590 1972 1593 2018
rect 1606 1982 1609 2018
rect 1702 1992 1705 2068
rect 1734 2062 1737 2068
rect 1814 2062 1817 2068
rect 1710 2052 1713 2058
rect 1782 2052 1785 2059
rect 1906 2058 1910 2061
rect 1730 2048 1734 2051
rect 1766 1992 1769 2038
rect 1642 1958 1646 1961
rect 1538 1748 1542 1751
rect 1530 1738 1534 1741
rect 1510 1718 1521 1721
rect 1502 1692 1505 1698
rect 1518 1682 1521 1718
rect 1462 1672 1465 1678
rect 1542 1672 1545 1738
rect 1550 1672 1553 1798
rect 1558 1762 1561 1928
rect 1574 1892 1577 1947
rect 1590 1942 1593 1948
rect 1606 1942 1609 1958
rect 1614 1952 1617 1958
rect 1706 1948 1710 1951
rect 1630 1942 1633 1948
rect 1758 1942 1761 1988
rect 1618 1888 1622 1891
rect 1662 1882 1665 1918
rect 1642 1868 1646 1871
rect 1682 1868 1686 1871
rect 1598 1862 1601 1868
rect 1710 1862 1713 1938
rect 1766 1932 1769 1948
rect 1734 1863 1737 1878
rect 1766 1872 1769 1878
rect 1634 1858 1638 1861
rect 1734 1858 1737 1859
rect 1614 1852 1617 1858
rect 1586 1838 1590 1841
rect 1558 1752 1561 1758
rect 1590 1752 1593 1808
rect 1614 1792 1617 1848
rect 1654 1802 1657 1818
rect 1614 1752 1617 1758
rect 1582 1742 1585 1748
rect 1574 1702 1577 1738
rect 1590 1722 1593 1748
rect 1630 1742 1633 1768
rect 1662 1742 1665 1747
rect 1610 1738 1614 1741
rect 1662 1682 1665 1728
rect 1590 1672 1593 1678
rect 1562 1668 1566 1671
rect 1382 1662 1385 1668
rect 1394 1658 1398 1661
rect 1370 1618 1374 1621
rect 1392 1603 1394 1607
rect 1398 1603 1401 1607
rect 1405 1603 1408 1607
rect 1422 1582 1425 1668
rect 1446 1662 1449 1668
rect 1614 1662 1617 1668
rect 1670 1662 1673 1818
rect 1710 1772 1713 1858
rect 1758 1792 1761 1808
rect 1722 1768 1726 1771
rect 1766 1752 1769 1768
rect 1774 1751 1777 2018
rect 1790 1952 1793 1958
rect 1790 1932 1793 1948
rect 1806 1942 1809 1978
rect 1822 1952 1825 2008
rect 1786 1878 1790 1881
rect 1806 1872 1809 1938
rect 1814 1872 1817 1918
rect 1830 1902 1833 2048
rect 1862 2002 1865 2018
rect 1926 1962 1929 1968
rect 1966 1962 1969 2058
rect 1846 1952 1849 1958
rect 1894 1952 1897 1958
rect 1866 1948 1870 1951
rect 1854 1942 1857 1948
rect 1926 1942 1929 1958
rect 1966 1952 1969 1958
rect 1890 1938 1894 1941
rect 1862 1922 1865 1938
rect 1838 1882 1841 1918
rect 1912 1903 1914 1907
rect 1918 1903 1921 1907
rect 1925 1903 1928 1907
rect 1850 1868 1854 1871
rect 1802 1858 1806 1861
rect 1782 1852 1785 1858
rect 1774 1748 1782 1751
rect 1726 1672 1729 1678
rect 1698 1668 1702 1671
rect 1554 1658 1558 1661
rect 1526 1652 1529 1658
rect 1382 1572 1385 1578
rect 1438 1562 1441 1618
rect 1510 1572 1513 1618
rect 1454 1562 1457 1568
rect 1358 1552 1361 1558
rect 1302 1532 1305 1538
rect 1334 1492 1337 1538
rect 1402 1528 1406 1531
rect 1390 1522 1393 1528
rect 1286 1472 1289 1478
rect 1318 1472 1321 1478
rect 1270 1468 1278 1471
rect 1130 1458 1142 1461
rect 1114 1428 1118 1431
rect 1126 1372 1129 1428
rect 1134 1422 1137 1448
rect 1166 1442 1169 1468
rect 1190 1452 1193 1458
rect 1214 1452 1217 1458
rect 1230 1452 1233 1468
rect 1238 1452 1241 1458
rect 1134 1382 1137 1418
rect 1174 1392 1177 1418
rect 1206 1412 1209 1428
rect 1206 1392 1209 1408
rect 1230 1382 1233 1388
rect 1198 1372 1201 1378
rect 1254 1372 1257 1468
rect 1262 1452 1265 1458
rect 1270 1382 1273 1468
rect 1298 1458 1302 1461
rect 1278 1452 1281 1458
rect 1318 1452 1321 1458
rect 1334 1452 1337 1478
rect 1366 1472 1369 1478
rect 1390 1472 1393 1518
rect 1398 1512 1401 1518
rect 1422 1472 1425 1558
rect 1486 1552 1489 1558
rect 1474 1548 1478 1551
rect 1454 1542 1457 1548
rect 1462 1532 1465 1538
rect 1430 1522 1433 1528
rect 1354 1468 1358 1471
rect 1402 1468 1406 1471
rect 1358 1452 1361 1458
rect 1306 1448 1310 1451
rect 1362 1448 1366 1451
rect 1218 1368 1222 1371
rect 1166 1362 1169 1368
rect 1194 1358 1198 1361
rect 1242 1358 1246 1361
rect 1150 1352 1153 1358
rect 1234 1348 1238 1351
rect 1110 1342 1113 1348
rect 1134 1342 1137 1348
rect 1158 1342 1161 1348
rect 1190 1342 1193 1348
rect 1254 1342 1257 1368
rect 1274 1358 1278 1361
rect 1294 1352 1297 1378
rect 1326 1372 1329 1418
rect 1310 1362 1313 1368
rect 1350 1352 1353 1358
rect 1266 1348 1270 1351
rect 1278 1342 1281 1348
rect 1122 1318 1126 1321
rect 1134 1302 1137 1338
rect 1158 1312 1161 1318
rect 1118 1262 1121 1298
rect 1150 1292 1153 1298
rect 1166 1282 1169 1308
rect 1166 1272 1169 1278
rect 1178 1268 1182 1271
rect 1150 1262 1153 1268
rect 1198 1262 1201 1268
rect 1118 1252 1121 1258
rect 1182 1252 1185 1258
rect 1110 1242 1113 1248
rect 1126 1222 1129 1248
rect 1102 1192 1105 1218
rect 1118 1182 1121 1218
rect 1134 1202 1137 1218
rect 1142 1192 1145 1248
rect 1150 1242 1153 1248
rect 1158 1222 1161 1248
rect 1118 1162 1121 1168
rect 1082 1158 1086 1161
rect 1134 1142 1137 1178
rect 1158 1172 1161 1218
rect 1174 1172 1177 1248
rect 1190 1172 1193 1248
rect 1206 1242 1209 1258
rect 1214 1252 1217 1278
rect 1238 1262 1241 1338
rect 1282 1328 1286 1331
rect 1246 1322 1249 1328
rect 1246 1262 1249 1318
rect 1190 1162 1193 1168
rect 1198 1162 1201 1218
rect 1214 1152 1217 1248
rect 1230 1172 1233 1218
rect 1238 1172 1241 1258
rect 1246 1232 1249 1248
rect 1262 1232 1265 1318
rect 1278 1292 1281 1328
rect 1294 1282 1297 1348
rect 1326 1322 1329 1348
rect 1358 1342 1361 1368
rect 1366 1342 1369 1348
rect 1334 1291 1337 1338
rect 1334 1288 1342 1291
rect 1342 1282 1345 1288
rect 1246 1192 1249 1228
rect 1262 1192 1265 1228
rect 1230 1162 1233 1168
rect 1254 1162 1257 1168
rect 1146 1148 1153 1151
rect 1138 1138 1145 1141
rect 1094 1132 1097 1138
rect 1070 1128 1081 1131
rect 1106 1128 1110 1131
rect 1062 1102 1065 1128
rect 1062 1072 1065 1078
rect 1070 1062 1073 1118
rect 926 962 929 968
rect 1006 962 1009 968
rect 1014 962 1017 978
rect 926 952 929 958
rect 950 952 953 958
rect 910 862 913 948
rect 854 852 857 859
rect 926 852 929 918
rect 934 872 937 888
rect 950 882 953 948
rect 958 932 961 958
rect 966 952 969 958
rect 990 942 993 948
rect 982 932 985 938
rect 1014 922 1017 958
rect 1022 952 1025 988
rect 1046 962 1049 968
rect 1070 962 1073 1008
rect 1078 1002 1081 1128
rect 1030 942 1033 948
rect 1086 942 1089 978
rect 1094 952 1097 1088
rect 1118 1012 1121 1118
rect 1126 1092 1129 1128
rect 1142 1092 1145 1138
rect 1150 1122 1153 1148
rect 1182 1142 1185 1148
rect 1230 1142 1233 1148
rect 1270 1142 1273 1178
rect 1278 1152 1281 1158
rect 1198 1132 1201 1138
rect 1214 1132 1217 1138
rect 1162 1128 1166 1131
rect 1182 1102 1185 1118
rect 1174 1072 1177 1078
rect 1134 1002 1137 1068
rect 1158 1042 1161 1058
rect 1162 1018 1166 1021
rect 1038 922 1041 938
rect 1070 931 1073 938
rect 1070 928 1078 931
rect 1006 911 1009 918
rect 1002 908 1009 911
rect 1046 882 1049 918
rect 954 868 958 871
rect 982 862 985 868
rect 1014 863 1017 868
rect 970 858 974 861
rect 1046 862 1049 868
rect 914 848 918 851
rect 954 848 958 851
rect 978 848 982 851
rect 938 838 942 841
rect 858 758 862 761
rect 838 752 841 758
rect 934 752 937 768
rect 954 748 958 751
rect 862 742 865 748
rect 806 732 809 738
rect 830 732 833 738
rect 894 722 897 738
rect 810 659 814 661
rect 806 658 814 659
rect 718 552 721 588
rect 458 538 462 541
rect 562 538 566 541
rect 514 528 521 531
rect 518 492 521 528
rect 466 488 470 491
rect 518 472 521 488
rect 446 442 449 448
rect 374 342 377 348
rect 394 288 398 291
rect 262 252 265 258
rect 286 252 289 258
rect 266 248 270 251
rect 294 182 297 268
rect 302 262 305 268
rect 294 162 297 178
rect 302 152 305 258
rect 366 202 369 268
rect 376 203 378 207
rect 382 203 385 207
rect 389 203 392 207
rect 406 192 409 388
rect 470 382 473 468
rect 478 462 481 468
rect 490 458 494 461
rect 502 452 505 468
rect 526 442 529 538
rect 558 452 561 458
rect 418 368 422 371
rect 446 342 449 368
rect 470 352 473 358
rect 510 352 513 358
rect 526 352 529 418
rect 498 348 502 351
rect 474 338 478 341
rect 522 338 526 341
rect 502 332 505 338
rect 518 272 521 288
rect 506 268 510 271
rect 422 262 425 268
rect 454 263 457 268
rect 470 222 473 268
rect 486 262 489 268
rect 534 262 537 428
rect 566 392 569 518
rect 662 472 665 538
rect 586 459 590 461
rect 586 458 593 459
rect 626 458 630 461
rect 622 422 625 448
rect 598 392 601 418
rect 570 348 574 351
rect 542 272 545 348
rect 582 342 585 348
rect 590 342 593 348
rect 598 331 601 378
rect 606 352 609 358
rect 590 328 601 331
rect 614 342 617 358
rect 622 352 625 358
rect 638 352 641 458
rect 646 452 649 468
rect 698 458 702 461
rect 646 382 649 448
rect 710 442 713 458
rect 694 392 697 408
rect 726 392 729 578
rect 734 482 737 518
rect 742 492 745 538
rect 766 532 769 558
rect 774 552 777 558
rect 782 542 785 548
rect 750 462 753 468
rect 758 451 761 518
rect 766 462 769 528
rect 754 448 761 451
rect 774 452 777 468
rect 790 462 793 588
rect 806 552 809 598
rect 814 542 817 548
rect 810 468 814 471
rect 790 452 793 458
rect 810 448 814 451
rect 822 442 825 668
rect 846 592 849 598
rect 766 372 769 398
rect 650 358 654 361
rect 726 352 729 368
rect 806 362 809 418
rect 830 392 833 548
rect 854 542 857 548
rect 838 402 841 418
rect 806 352 809 358
rect 786 348 790 351
rect 614 332 617 338
rect 590 272 593 328
rect 614 302 617 328
rect 498 258 502 261
rect 534 252 537 258
rect 346 158 350 161
rect 290 148 294 151
rect 346 148 350 151
rect 338 118 342 121
rect 366 112 369 138
rect 358 72 361 88
rect 294 62 297 68
rect 310 62 313 68
rect 350 62 353 68
rect 374 62 377 148
rect 390 92 393 148
rect 398 92 401 158
rect 430 152 433 158
rect 438 152 441 188
rect 470 171 473 218
rect 470 168 481 171
rect 422 141 425 148
rect 462 142 465 148
rect 478 142 481 168
rect 518 152 521 248
rect 542 192 545 268
rect 574 252 577 258
rect 558 242 561 248
rect 582 242 585 258
rect 554 188 558 191
rect 578 148 582 151
rect 590 142 593 268
rect 606 222 609 268
rect 630 192 633 328
rect 638 262 641 318
rect 678 291 681 348
rect 702 292 705 348
rect 710 342 713 348
rect 822 342 825 348
rect 718 332 721 338
rect 750 332 753 338
rect 678 288 686 291
rect 698 288 702 291
rect 758 263 761 268
rect 598 152 601 158
rect 638 142 641 178
rect 670 162 673 238
rect 646 152 649 158
rect 422 138 433 141
rect 562 138 566 141
rect 678 141 681 158
rect 718 151 721 158
rect 726 142 729 258
rect 774 182 777 338
rect 802 318 806 321
rect 790 272 793 288
rect 810 268 814 271
rect 810 248 814 251
rect 830 242 833 348
rect 838 272 841 298
rect 846 262 849 528
rect 854 392 857 398
rect 870 352 873 718
rect 880 703 882 707
rect 886 703 889 707
rect 893 703 896 707
rect 878 672 881 688
rect 878 662 881 668
rect 918 661 921 728
rect 950 692 953 728
rect 958 672 961 678
rect 982 662 985 788
rect 998 752 1001 788
rect 1070 771 1073 918
rect 1078 892 1081 928
rect 1086 872 1089 918
rect 1094 902 1097 938
rect 1094 862 1097 898
rect 1094 792 1097 858
rect 1066 768 1073 771
rect 1102 762 1105 938
rect 1110 792 1113 848
rect 1030 752 1033 758
rect 1006 742 1009 748
rect 1038 742 1041 748
rect 1046 732 1049 758
rect 1078 752 1081 758
rect 1118 752 1121 988
rect 1134 952 1137 988
rect 1142 982 1145 1018
rect 1182 982 1185 1098
rect 1190 1092 1193 1118
rect 1262 1092 1265 1118
rect 1234 1068 1238 1071
rect 1206 1052 1209 1058
rect 1206 992 1209 1038
rect 1142 962 1145 968
rect 1158 962 1161 978
rect 1126 932 1129 948
rect 1126 842 1129 868
rect 1134 812 1137 948
rect 1158 942 1161 958
rect 1142 882 1145 888
rect 1142 792 1145 868
rect 1150 772 1153 918
rect 1114 748 1118 751
rect 1054 742 1057 748
rect 1082 738 1086 741
rect 1094 732 1097 738
rect 1026 678 1030 681
rect 994 668 998 671
rect 1010 668 1014 671
rect 918 658 926 661
rect 886 552 889 658
rect 934 652 937 658
rect 990 651 993 658
rect 986 648 993 651
rect 910 592 913 628
rect 918 552 921 618
rect 942 602 945 648
rect 958 582 961 648
rect 1022 582 1025 668
rect 1046 662 1049 688
rect 1054 672 1057 708
rect 1062 672 1065 718
rect 1094 692 1097 718
rect 1086 682 1089 688
rect 1034 658 1038 661
rect 1050 658 1057 661
rect 1066 658 1070 661
rect 1034 648 1041 651
rect 1038 592 1041 648
rect 966 552 969 578
rect 1026 568 1030 571
rect 1046 562 1049 568
rect 1054 562 1057 658
rect 1082 648 1086 651
rect 1086 592 1089 638
rect 1094 632 1097 648
rect 1102 642 1105 738
rect 1110 672 1113 698
rect 1126 692 1129 758
rect 1134 722 1137 758
rect 1146 748 1150 751
rect 1122 668 1126 671
rect 1110 592 1113 608
rect 1074 568 1078 571
rect 1094 562 1097 568
rect 1118 562 1121 668
rect 1034 558 1038 561
rect 894 542 897 548
rect 880 503 882 507
rect 886 503 889 507
rect 893 503 896 507
rect 942 502 945 538
rect 942 472 945 498
rect 950 482 953 508
rect 950 472 953 478
rect 998 472 1001 488
rect 1014 472 1017 498
rect 978 468 982 471
rect 878 462 881 468
rect 902 442 905 468
rect 1030 463 1033 468
rect 962 458 966 461
rect 982 452 985 458
rect 894 352 897 368
rect 862 292 865 348
rect 870 342 873 348
rect 880 303 882 307
rect 886 303 889 307
rect 893 303 896 307
rect 902 262 905 438
rect 982 392 985 448
rect 958 351 961 368
rect 990 352 993 438
rect 1038 432 1041 558
rect 1046 542 1049 558
rect 1070 542 1073 558
rect 1126 552 1129 658
rect 1114 548 1118 551
rect 1110 538 1118 541
rect 1078 492 1081 528
rect 1110 492 1113 538
rect 1090 488 1094 491
rect 1134 482 1137 698
rect 1142 672 1145 698
rect 1158 682 1161 918
rect 1174 902 1177 918
rect 1166 852 1169 858
rect 1174 852 1177 888
rect 1182 841 1185 868
rect 1190 862 1193 978
rect 1198 942 1201 948
rect 1214 942 1217 1058
rect 1222 972 1225 1058
rect 1246 1052 1249 1088
rect 1286 1082 1289 1268
rect 1298 1258 1302 1261
rect 1350 1252 1353 1318
rect 1374 1272 1377 1438
rect 1414 1422 1417 1458
rect 1438 1422 1441 1448
rect 1392 1403 1394 1407
rect 1398 1403 1401 1407
rect 1405 1403 1408 1407
rect 1430 1362 1433 1368
rect 1410 1358 1414 1361
rect 1438 1352 1441 1418
rect 1446 1382 1449 1518
rect 1454 1472 1457 1508
rect 1478 1472 1481 1478
rect 1486 1472 1489 1528
rect 1494 1502 1497 1548
rect 1534 1532 1537 1658
rect 1542 1622 1545 1658
rect 1574 1652 1577 1658
rect 1550 1552 1553 1648
rect 1678 1642 1681 1668
rect 1718 1652 1721 1658
rect 1690 1648 1694 1651
rect 1558 1542 1561 1638
rect 1678 1602 1681 1638
rect 1586 1568 1590 1571
rect 1606 1562 1609 1568
rect 1702 1562 1705 1568
rect 1718 1562 1721 1568
rect 1566 1552 1569 1558
rect 1574 1542 1577 1558
rect 1598 1552 1601 1558
rect 1670 1551 1673 1558
rect 1554 1538 1558 1541
rect 1518 1522 1521 1528
rect 1494 1482 1497 1498
rect 1466 1468 1470 1471
rect 1510 1471 1513 1518
rect 1534 1492 1537 1518
rect 1542 1482 1545 1488
rect 1510 1468 1521 1471
rect 1490 1458 1494 1461
rect 1506 1458 1510 1461
rect 1454 1452 1457 1458
rect 1498 1448 1502 1451
rect 1518 1442 1521 1468
rect 1550 1462 1553 1508
rect 1566 1452 1569 1458
rect 1530 1418 1534 1421
rect 1470 1362 1473 1408
rect 1534 1392 1537 1398
rect 1482 1358 1486 1361
rect 1386 1348 1390 1351
rect 1386 1338 1390 1341
rect 1430 1332 1433 1348
rect 1446 1342 1449 1358
rect 1438 1332 1441 1338
rect 1382 1312 1385 1318
rect 1418 1288 1422 1291
rect 1382 1272 1385 1278
rect 1358 1262 1361 1268
rect 1366 1252 1369 1258
rect 1310 1152 1313 1168
rect 1294 1102 1297 1118
rect 1286 1072 1289 1078
rect 1262 1062 1265 1068
rect 1262 1042 1265 1048
rect 1270 1012 1273 1068
rect 1310 1062 1313 1078
rect 1294 992 1297 1008
rect 1222 952 1225 968
rect 1230 962 1233 978
rect 1246 952 1249 958
rect 1286 952 1289 958
rect 1278 942 1281 948
rect 1206 922 1209 928
rect 1210 888 1214 891
rect 1238 882 1241 918
rect 1254 892 1257 938
rect 1262 932 1265 938
rect 1302 922 1305 928
rect 1206 852 1209 878
rect 1246 862 1249 888
rect 1262 862 1265 868
rect 1174 838 1185 841
rect 1174 792 1177 838
rect 1174 722 1177 728
rect 1170 668 1174 671
rect 1142 652 1145 668
rect 1182 662 1185 768
rect 1210 758 1214 761
rect 1198 752 1201 758
rect 1242 748 1246 751
rect 1262 742 1265 858
rect 1270 792 1273 918
rect 1310 911 1313 958
rect 1326 952 1329 958
rect 1326 932 1329 938
rect 1302 908 1313 911
rect 1302 892 1305 908
rect 1318 892 1321 918
rect 1298 888 1302 891
rect 1314 888 1318 891
rect 1342 862 1345 868
rect 1302 752 1305 758
rect 1350 752 1353 1198
rect 1358 1032 1361 1068
rect 1366 1061 1369 1248
rect 1374 1212 1377 1268
rect 1430 1262 1433 1328
rect 1454 1312 1457 1348
rect 1446 1272 1449 1278
rect 1454 1272 1457 1288
rect 1438 1262 1441 1268
rect 1394 1248 1398 1251
rect 1414 1242 1417 1248
rect 1422 1242 1425 1258
rect 1462 1251 1465 1338
rect 1470 1332 1473 1358
rect 1534 1342 1537 1348
rect 1486 1302 1489 1328
rect 1498 1318 1502 1321
rect 1526 1292 1529 1298
rect 1518 1272 1521 1278
rect 1470 1262 1473 1268
rect 1462 1248 1470 1251
rect 1478 1242 1481 1248
rect 1392 1203 1394 1207
rect 1398 1203 1401 1207
rect 1405 1203 1408 1207
rect 1374 1151 1377 1168
rect 1390 1132 1393 1138
rect 1374 1072 1377 1098
rect 1414 1092 1417 1238
rect 1438 1162 1441 1218
rect 1462 1192 1465 1218
rect 1422 1142 1425 1148
rect 1446 1142 1449 1168
rect 1462 1152 1465 1158
rect 1494 1152 1497 1258
rect 1534 1202 1537 1338
rect 1530 1158 1534 1161
rect 1514 1148 1518 1151
rect 1470 1102 1473 1138
rect 1478 1132 1481 1148
rect 1490 1138 1494 1141
rect 1542 1141 1545 1438
rect 1558 1362 1561 1368
rect 1558 1212 1561 1258
rect 1538 1138 1545 1141
rect 1550 1142 1553 1178
rect 1558 1162 1561 1168
rect 1574 1152 1577 1508
rect 1590 1462 1593 1468
rect 1582 1442 1585 1458
rect 1598 1361 1601 1548
rect 1714 1548 1718 1551
rect 1726 1542 1729 1668
rect 1734 1642 1737 1748
rect 1742 1702 1745 1748
rect 1750 1652 1753 1658
rect 1758 1652 1761 1678
rect 1742 1632 1745 1638
rect 1742 1552 1745 1598
rect 1638 1501 1641 1518
rect 1630 1498 1641 1501
rect 1630 1462 1633 1498
rect 1646 1492 1649 1498
rect 1642 1488 1646 1491
rect 1686 1472 1689 1538
rect 1734 1512 1737 1548
rect 1750 1532 1753 1618
rect 1766 1532 1769 1668
rect 1782 1662 1785 1748
rect 1798 1672 1801 1718
rect 1774 1652 1777 1658
rect 1786 1648 1790 1651
rect 1806 1642 1809 1738
rect 1814 1672 1817 1868
rect 1830 1862 1833 1868
rect 1862 1862 1865 1898
rect 1878 1862 1881 1878
rect 1942 1862 1945 1868
rect 1966 1862 1969 1868
rect 1822 1822 1825 1858
rect 1870 1852 1873 1858
rect 1830 1762 1833 1788
rect 1854 1762 1857 1768
rect 1862 1762 1865 1838
rect 1862 1752 1865 1758
rect 1886 1752 1889 1818
rect 1894 1762 1897 1818
rect 1902 1792 1905 1858
rect 1934 1852 1937 1858
rect 1822 1682 1825 1718
rect 1818 1668 1822 1671
rect 1830 1662 1833 1748
rect 1878 1742 1881 1748
rect 1838 1732 1841 1738
rect 1846 1712 1849 1718
rect 1846 1662 1849 1668
rect 1774 1541 1777 1638
rect 1806 1582 1809 1618
rect 1830 1592 1833 1658
rect 1862 1652 1865 1718
rect 1886 1702 1889 1748
rect 1894 1742 1897 1748
rect 1894 1672 1897 1728
rect 1934 1722 1937 1848
rect 1974 1832 1977 2068
rect 1986 2058 1990 2061
rect 1990 1942 1993 1948
rect 1998 1872 2001 2018
rect 2014 1982 2017 2058
rect 2022 2052 2025 2058
rect 2030 1992 2033 2068
rect 2078 2062 2081 2068
rect 2038 2052 2041 2058
rect 2066 2048 2070 2051
rect 2030 1942 2033 1988
rect 2078 1972 2081 1978
rect 2062 1952 2065 1958
rect 2042 1948 2046 1951
rect 2050 1938 2054 1941
rect 2014 1862 2017 1868
rect 2038 1862 2041 1878
rect 2046 1872 2049 1878
rect 2026 1858 2030 1861
rect 1982 1852 1985 1858
rect 1942 1752 1945 1778
rect 1950 1772 1953 1818
rect 1990 1812 1993 1858
rect 2062 1842 2065 1948
rect 2078 1942 2081 1968
rect 2070 1862 2073 1898
rect 2078 1882 2081 1888
rect 1998 1792 2001 1818
rect 1950 1752 1953 1758
rect 1982 1752 1985 1768
rect 1990 1752 1993 1758
rect 2046 1752 2049 1768
rect 2086 1762 2089 2068
rect 2110 2062 2113 2088
rect 2218 2068 2222 2071
rect 2234 2068 2238 2071
rect 2150 2062 2153 2068
rect 2102 2022 2105 2048
rect 2094 1771 2097 2018
rect 2118 1952 2121 1958
rect 2166 1952 2169 2068
rect 2238 2052 2241 2058
rect 2246 2052 2249 2058
rect 2302 2052 2305 2068
rect 2258 2048 2262 2051
rect 2206 2041 2209 2048
rect 2198 2038 2209 2041
rect 2198 1951 2201 2038
rect 2266 2018 2270 2021
rect 2214 1961 2217 2018
rect 2210 1958 2217 1961
rect 2194 1948 2201 1951
rect 2246 1952 2249 1958
rect 2118 1861 2121 1948
rect 2142 1942 2145 1948
rect 2166 1942 2169 1948
rect 2174 1872 2177 1888
rect 2114 1858 2121 1861
rect 2142 1863 2145 1868
rect 2094 1768 2102 1771
rect 2102 1752 2105 1758
rect 1912 1703 1914 1707
rect 1918 1703 1921 1707
rect 1925 1703 1928 1707
rect 1942 1692 1945 1738
rect 1878 1663 1881 1668
rect 1842 1648 1846 1651
rect 1782 1552 1785 1568
rect 1838 1562 1841 1638
rect 1850 1568 1854 1571
rect 1802 1558 1806 1561
rect 1838 1552 1841 1558
rect 1814 1542 1817 1548
rect 1774 1538 1782 1541
rect 1794 1538 1798 1541
rect 1834 1538 1838 1541
rect 1754 1518 1758 1521
rect 1726 1472 1729 1488
rect 1782 1482 1785 1538
rect 1790 1472 1793 1498
rect 1638 1462 1641 1468
rect 1706 1459 1710 1461
rect 1706 1458 1713 1459
rect 1606 1452 1609 1458
rect 1742 1422 1745 1468
rect 1762 1458 1766 1461
rect 1750 1452 1753 1458
rect 1770 1448 1774 1451
rect 1598 1358 1606 1361
rect 1622 1361 1625 1418
rect 1638 1362 1641 1378
rect 1622 1358 1630 1361
rect 1582 1352 1585 1358
rect 1582 1332 1585 1338
rect 1590 1302 1593 1338
rect 1598 1312 1601 1358
rect 1630 1342 1633 1348
rect 1646 1342 1649 1348
rect 1610 1338 1614 1341
rect 1590 1263 1593 1268
rect 1606 1252 1609 1318
rect 1626 1268 1630 1271
rect 1638 1262 1641 1308
rect 1654 1302 1657 1368
rect 1670 1362 1673 1418
rect 1702 1358 1710 1361
rect 1702 1352 1705 1358
rect 1666 1338 1670 1341
rect 1690 1338 1694 1341
rect 1702 1332 1705 1338
rect 1710 1322 1713 1348
rect 1670 1312 1673 1318
rect 1694 1292 1697 1298
rect 1718 1292 1721 1418
rect 1726 1362 1729 1368
rect 1738 1348 1742 1351
rect 1734 1332 1737 1338
rect 1742 1272 1745 1328
rect 1650 1268 1654 1271
rect 1686 1262 1689 1268
rect 1750 1262 1753 1448
rect 1766 1352 1769 1358
rect 1782 1342 1785 1358
rect 1790 1342 1793 1438
rect 1798 1372 1801 1518
rect 1806 1352 1809 1358
rect 1762 1338 1766 1341
rect 1798 1281 1801 1288
rect 1794 1278 1801 1281
rect 1790 1272 1793 1278
rect 1770 1268 1774 1271
rect 1622 1252 1625 1258
rect 1670 1242 1673 1258
rect 1682 1248 1686 1251
rect 1706 1248 1710 1251
rect 1658 1238 1662 1241
rect 1622 1192 1625 1198
rect 1602 1158 1606 1161
rect 1634 1158 1638 1161
rect 1562 1138 1566 1141
rect 1574 1132 1577 1148
rect 1590 1142 1593 1148
rect 1638 1142 1641 1148
rect 1646 1142 1649 1188
rect 1654 1152 1657 1218
rect 1666 1158 1670 1161
rect 1726 1158 1734 1161
rect 1670 1142 1673 1148
rect 1486 1082 1489 1118
rect 1518 1112 1521 1118
rect 1542 1112 1545 1118
rect 1390 1072 1393 1078
rect 1486 1072 1489 1078
rect 1494 1072 1497 1108
rect 1366 1058 1374 1061
rect 1374 1052 1377 1058
rect 1418 1048 1422 1051
rect 1370 1038 1374 1041
rect 1358 952 1361 1028
rect 1392 1003 1394 1007
rect 1398 1003 1401 1007
rect 1405 1003 1408 1007
rect 1422 962 1425 1048
rect 1438 1042 1441 1068
rect 1458 1058 1462 1061
rect 1474 1058 1478 1061
rect 1458 1048 1462 1051
rect 1486 1051 1489 1058
rect 1482 1048 1489 1051
rect 1438 952 1441 978
rect 1482 958 1489 961
rect 1426 948 1430 951
rect 1474 948 1478 951
rect 1358 922 1361 938
rect 1470 892 1473 918
rect 1406 872 1409 888
rect 1470 872 1473 878
rect 1442 868 1446 871
rect 1374 863 1377 868
rect 1458 858 1462 861
rect 1438 852 1441 858
rect 1478 852 1481 898
rect 1486 892 1489 958
rect 1494 952 1497 1008
rect 1494 902 1497 948
rect 1502 942 1505 1098
rect 1518 1052 1521 1088
rect 1550 1082 1553 1118
rect 1582 1092 1585 1138
rect 1614 1132 1617 1138
rect 1566 1072 1569 1078
rect 1606 1072 1609 1118
rect 1594 1068 1598 1071
rect 1586 1058 1590 1061
rect 1538 1048 1542 1051
rect 1518 1032 1521 1048
rect 1526 992 1529 1048
rect 1510 962 1513 988
rect 1550 972 1553 1058
rect 1566 962 1569 1058
rect 1598 1051 1601 1058
rect 1594 1048 1601 1051
rect 1574 1042 1577 1048
rect 1566 952 1569 958
rect 1522 948 1526 951
rect 1494 872 1497 888
rect 1518 872 1521 908
rect 1534 872 1537 888
rect 1494 852 1497 868
rect 1392 803 1394 807
rect 1398 803 1401 807
rect 1405 803 1408 807
rect 1366 752 1369 758
rect 1382 752 1385 758
rect 1430 752 1433 778
rect 1438 752 1441 758
rect 1194 738 1198 741
rect 1226 738 1230 741
rect 1198 672 1201 678
rect 1214 672 1217 718
rect 1254 682 1257 708
rect 1294 692 1297 698
rect 1234 668 1238 671
rect 1158 652 1161 658
rect 1158 592 1161 648
rect 1158 552 1161 578
rect 1166 552 1169 598
rect 1178 568 1182 571
rect 1030 372 1033 378
rect 1046 362 1049 388
rect 1010 358 1014 361
rect 990 342 993 348
rect 974 322 977 338
rect 1006 332 1009 358
rect 1038 352 1041 358
rect 1034 338 1038 341
rect 910 262 913 318
rect 974 292 977 308
rect 998 292 1001 298
rect 1010 288 1014 291
rect 1046 281 1049 358
rect 1062 342 1065 458
rect 1094 392 1097 448
rect 1102 442 1105 478
rect 1158 462 1161 548
rect 1126 452 1129 458
rect 1138 428 1142 431
rect 1150 402 1153 458
rect 1166 392 1169 458
rect 1174 452 1177 458
rect 1182 392 1185 538
rect 1190 512 1193 668
rect 1206 582 1209 658
rect 1222 642 1225 648
rect 1262 632 1265 668
rect 1278 652 1281 678
rect 1286 662 1289 668
rect 1282 648 1286 651
rect 1310 642 1313 748
rect 1346 738 1350 741
rect 1418 738 1422 741
rect 1398 722 1401 738
rect 1346 718 1350 721
rect 1430 682 1433 708
rect 1426 678 1430 681
rect 1338 658 1342 661
rect 1326 631 1329 658
rect 1390 641 1393 668
rect 1446 662 1449 788
rect 1454 762 1457 778
rect 1478 772 1481 848
rect 1510 762 1513 818
rect 1486 742 1489 758
rect 1518 752 1521 868
rect 1526 862 1529 868
rect 1542 861 1545 938
rect 1550 891 1553 918
rect 1550 888 1561 891
rect 1550 872 1553 878
rect 1558 872 1561 888
rect 1582 882 1585 1008
rect 1590 992 1593 1038
rect 1614 1012 1617 1128
rect 1626 1078 1630 1081
rect 1638 1072 1641 1138
rect 1658 1128 1662 1131
rect 1678 1122 1681 1138
rect 1690 1128 1694 1131
rect 1674 1088 1678 1091
rect 1678 1072 1681 1078
rect 1666 1068 1670 1071
rect 1634 1058 1638 1061
rect 1650 1058 1654 1061
rect 1630 922 1633 947
rect 1606 892 1609 918
rect 1614 882 1617 888
rect 1578 878 1582 881
rect 1570 868 1574 871
rect 1534 858 1545 861
rect 1558 862 1561 868
rect 1534 852 1537 858
rect 1546 848 1550 851
rect 1506 748 1510 751
rect 1470 732 1473 738
rect 1498 688 1502 691
rect 1410 658 1414 661
rect 1462 652 1465 658
rect 1382 638 1393 641
rect 1430 648 1438 651
rect 1326 628 1337 631
rect 1222 592 1225 628
rect 1322 588 1326 591
rect 1206 562 1209 578
rect 1214 572 1217 578
rect 1314 568 1318 571
rect 1238 562 1241 568
rect 1294 562 1297 568
rect 1326 562 1329 568
rect 1258 558 1273 561
rect 1230 551 1233 558
rect 1230 548 1241 551
rect 1198 472 1201 548
rect 1222 492 1225 548
rect 1230 472 1233 518
rect 1238 492 1241 548
rect 1206 442 1209 458
rect 1214 432 1217 448
rect 1230 392 1233 448
rect 1070 352 1073 358
rect 1102 352 1105 378
rect 1134 362 1137 368
rect 1166 362 1169 388
rect 1246 372 1249 558
rect 1262 542 1265 548
rect 1270 542 1273 558
rect 1302 542 1305 548
rect 1254 532 1257 538
rect 1326 522 1329 538
rect 1278 502 1281 518
rect 1334 511 1337 628
rect 1382 612 1385 638
rect 1392 603 1394 607
rect 1398 603 1401 607
rect 1405 603 1408 607
rect 1414 592 1417 648
rect 1430 592 1433 648
rect 1342 542 1345 558
rect 1350 552 1353 558
rect 1358 552 1361 568
rect 1382 542 1385 548
rect 1366 532 1369 538
rect 1422 532 1425 578
rect 1334 508 1345 511
rect 1254 472 1257 478
rect 1318 462 1321 488
rect 1342 472 1345 508
rect 1378 488 1382 491
rect 1406 472 1409 498
rect 1430 472 1433 528
rect 1438 522 1441 558
rect 1446 542 1449 638
rect 1470 592 1473 668
rect 1510 662 1513 718
rect 1518 702 1521 748
rect 1558 742 1561 858
rect 1550 738 1558 741
rect 1534 722 1537 738
rect 1534 662 1537 718
rect 1550 662 1553 738
rect 1582 731 1585 878
rect 1630 872 1633 908
rect 1594 868 1598 871
rect 1622 852 1625 858
rect 1638 842 1641 1048
rect 1678 1042 1681 1068
rect 1654 912 1657 1018
rect 1662 952 1665 978
rect 1686 962 1689 1118
rect 1694 1092 1697 1128
rect 1710 1102 1713 1118
rect 1726 1052 1729 1158
rect 1742 1151 1745 1258
rect 1750 1232 1753 1258
rect 1774 1232 1777 1248
rect 1738 1148 1745 1151
rect 1798 1158 1806 1161
rect 1734 1012 1737 1148
rect 1750 1142 1753 1158
rect 1798 1152 1801 1158
rect 1758 1142 1761 1148
rect 1766 1082 1769 1128
rect 1782 1122 1785 1138
rect 1798 1132 1801 1138
rect 1806 1082 1809 1148
rect 1742 1052 1745 1058
rect 1750 981 1753 1068
rect 1766 991 1769 1078
rect 1814 1072 1817 1538
rect 1830 1458 1838 1461
rect 1830 1392 1833 1458
rect 1846 1362 1849 1368
rect 1826 1348 1830 1351
rect 1862 1342 1865 1618
rect 1894 1492 1897 1668
rect 1950 1642 1953 1748
rect 1970 1738 1977 1741
rect 2002 1738 2006 1741
rect 1974 1722 1977 1738
rect 1966 1662 1969 1718
rect 1974 1662 1977 1668
rect 1966 1562 1969 1658
rect 1990 1652 1993 1658
rect 1998 1652 2001 1658
rect 2006 1642 2009 1718
rect 2014 1662 2017 1688
rect 2030 1672 2033 1678
rect 1990 1572 1993 1638
rect 2014 1592 2017 1648
rect 2022 1572 2025 1658
rect 2070 1552 2073 1748
rect 2086 1732 2089 1738
rect 2110 1732 2113 1858
rect 2182 1822 2185 1938
rect 2190 1862 2193 1868
rect 2190 1842 2193 1848
rect 2154 1778 2158 1781
rect 2150 1752 2153 1758
rect 2122 1738 2126 1741
rect 2078 1672 2081 1678
rect 2110 1672 2113 1728
rect 2134 1702 2137 1738
rect 2190 1732 2193 1748
rect 2126 1652 2129 1659
rect 2110 1552 2113 1558
rect 1994 1548 1998 1551
rect 2090 1548 2094 1551
rect 1902 1542 1905 1548
rect 1912 1503 1914 1507
rect 1918 1503 1921 1507
rect 1925 1503 1928 1507
rect 1942 1492 1945 1538
rect 1878 1472 1881 1488
rect 1894 1472 1897 1478
rect 1882 1368 1886 1371
rect 1834 1338 1838 1341
rect 1830 1171 1833 1288
rect 1838 1262 1841 1268
rect 1854 1252 1857 1318
rect 1822 1168 1833 1171
rect 1822 1162 1825 1168
rect 1830 1152 1833 1158
rect 1838 1131 1841 1238
rect 1862 1202 1865 1338
rect 1894 1332 1897 1468
rect 1902 1452 1905 1458
rect 1926 1452 1929 1468
rect 1938 1458 1942 1461
rect 1926 1352 1929 1358
rect 1942 1332 1945 1448
rect 1950 1342 1953 1488
rect 1958 1472 1961 1528
rect 1974 1372 1977 1538
rect 2006 1532 2009 1548
rect 2030 1532 2033 1548
rect 2050 1538 2054 1541
rect 2074 1538 2078 1541
rect 1982 1512 1985 1518
rect 2006 1492 2009 1528
rect 1990 1482 1993 1488
rect 2046 1482 2049 1538
rect 2054 1492 2057 1498
rect 2070 1482 2073 1488
rect 1990 1463 1993 1468
rect 2022 1462 2025 1468
rect 2070 1462 2073 1468
rect 2102 1463 2105 1518
rect 2102 1458 2105 1459
rect 1982 1362 1985 1368
rect 1998 1352 2001 1408
rect 1912 1303 1914 1307
rect 1918 1303 1921 1307
rect 1925 1303 1928 1307
rect 1894 1282 1897 1288
rect 1878 1272 1881 1278
rect 1934 1272 1937 1318
rect 1958 1292 1961 1308
rect 1966 1272 1969 1338
rect 1982 1271 1985 1318
rect 1998 1302 2001 1348
rect 2006 1342 2009 1358
rect 2030 1342 2033 1368
rect 2062 1362 2065 1418
rect 2110 1392 2113 1548
rect 2126 1542 2129 1568
rect 2142 1561 2145 1718
rect 2158 1672 2161 1678
rect 2166 1592 2169 1698
rect 2174 1652 2177 1658
rect 2182 1652 2185 1668
rect 2198 1662 2201 1948
rect 2206 1912 2209 1918
rect 2214 1902 2217 1918
rect 2230 1872 2233 1898
rect 2254 1892 2257 1948
rect 2274 1868 2278 1871
rect 2214 1842 2217 1858
rect 2222 1812 2225 1868
rect 2270 1852 2273 1858
rect 2250 1848 2254 1851
rect 2206 1742 2209 1808
rect 2218 1748 2222 1751
rect 2254 1742 2257 1778
rect 2270 1762 2273 1848
rect 2266 1758 2270 1761
rect 2294 1752 2297 1758
rect 2278 1742 2281 1748
rect 2302 1742 2305 1818
rect 2206 1672 2209 1738
rect 2234 1668 2238 1671
rect 2166 1582 2169 1588
rect 2138 1558 2145 1561
rect 2138 1548 2142 1551
rect 2150 1522 2153 1548
rect 2158 1542 2161 1548
rect 2166 1492 2169 1568
rect 2174 1472 2177 1538
rect 2198 1522 2201 1658
rect 2206 1542 2209 1668
rect 2214 1562 2217 1668
rect 2234 1648 2238 1651
rect 2222 1562 2225 1618
rect 2262 1562 2265 1568
rect 2278 1552 2281 1648
rect 2218 1548 2222 1551
rect 2246 1542 2249 1548
rect 2246 1472 2249 1538
rect 2230 1463 2233 1468
rect 2178 1458 2182 1461
rect 2194 1458 2198 1461
rect 2082 1368 2086 1371
rect 2074 1358 2078 1361
rect 2046 1352 2049 1358
rect 2066 1348 2070 1351
rect 2078 1342 2081 1348
rect 2134 1342 2137 1458
rect 2142 1352 2145 1358
rect 2014 1322 2017 1328
rect 2038 1292 2041 1328
rect 1974 1268 1985 1271
rect 1906 1258 1910 1261
rect 1894 1242 1897 1248
rect 1846 1142 1849 1178
rect 1886 1172 1889 1218
rect 1886 1162 1889 1168
rect 1926 1152 1929 1168
rect 1858 1148 1862 1151
rect 1882 1148 1886 1151
rect 1858 1138 1862 1141
rect 1838 1128 1849 1131
rect 1834 1118 1838 1121
rect 1838 1072 1841 1108
rect 1846 1092 1849 1128
rect 1918 1122 1921 1138
rect 1912 1103 1914 1107
rect 1918 1103 1921 1107
rect 1925 1103 1928 1107
rect 1862 1072 1865 1098
rect 1890 1068 1894 1071
rect 1782 1062 1785 1068
rect 1798 1052 1801 1058
rect 1806 1052 1809 1068
rect 1830 1062 1833 1068
rect 1818 1058 1822 1061
rect 1766 988 1777 991
rect 1750 978 1758 981
rect 1742 952 1745 968
rect 1758 952 1761 978
rect 1694 912 1697 918
rect 1658 888 1662 891
rect 1650 878 1654 881
rect 1670 862 1673 908
rect 1774 882 1777 988
rect 1810 968 1814 971
rect 1830 952 1833 958
rect 1802 948 1806 951
rect 1790 922 1793 938
rect 1798 902 1801 938
rect 1830 892 1833 918
rect 1838 902 1841 1068
rect 1870 1062 1873 1068
rect 1886 1058 1894 1061
rect 1870 1052 1873 1058
rect 1858 1048 1862 1051
rect 1874 948 1878 951
rect 1886 942 1889 1058
rect 1898 1048 1902 1051
rect 1850 938 1854 941
rect 1878 938 1886 941
rect 1690 878 1694 881
rect 1766 872 1769 878
rect 1790 872 1793 878
rect 1838 872 1841 878
rect 1682 868 1686 871
rect 1714 868 1718 871
rect 1810 868 1825 871
rect 1786 858 1790 861
rect 1810 858 1814 861
rect 1658 848 1662 851
rect 1670 842 1673 858
rect 1686 852 1689 858
rect 1598 792 1601 838
rect 1638 812 1641 838
rect 1646 752 1649 818
rect 1602 738 1606 741
rect 1574 728 1585 731
rect 1562 718 1566 721
rect 1574 682 1577 728
rect 1582 712 1585 718
rect 1606 701 1609 738
rect 1654 722 1657 738
rect 1686 702 1689 848
rect 1702 792 1705 858
rect 1718 842 1721 858
rect 1754 848 1758 851
rect 1730 838 1734 841
rect 1730 768 1734 771
rect 1730 758 1734 761
rect 1742 752 1745 848
rect 1766 842 1769 858
rect 1798 852 1801 858
rect 1822 851 1825 868
rect 1838 852 1841 858
rect 1814 848 1825 851
rect 1782 792 1785 818
rect 1814 792 1817 848
rect 1830 812 1833 848
rect 1854 832 1857 868
rect 1862 842 1865 918
rect 1870 862 1873 938
rect 1802 768 1806 771
rect 1846 762 1849 768
rect 1862 762 1865 838
rect 1870 792 1873 848
rect 1878 822 1881 938
rect 1894 902 1897 918
rect 1894 862 1897 878
rect 1902 862 1905 988
rect 1918 972 1921 1018
rect 1918 952 1921 958
rect 1942 952 1945 1258
rect 1958 1151 1961 1158
rect 1966 1142 1969 1268
rect 1974 1182 1977 1268
rect 2006 1262 2009 1278
rect 2030 1272 2033 1288
rect 2070 1262 2073 1318
rect 2078 1262 2081 1268
rect 2086 1262 2089 1308
rect 2106 1278 2110 1281
rect 2134 1272 2137 1288
rect 1994 1258 1998 1261
rect 2026 1258 2030 1261
rect 2098 1258 2102 1261
rect 1982 1252 1985 1258
rect 2018 1168 2022 1171
rect 2030 1142 2033 1248
rect 2038 1102 2041 1148
rect 2046 1122 2049 1258
rect 2054 1222 2057 1248
rect 2058 1148 2062 1151
rect 2030 1082 2033 1088
rect 2030 1072 2033 1078
rect 1974 1062 1977 1068
rect 2014 982 2017 1068
rect 2046 1062 2049 1118
rect 2070 1092 2073 1148
rect 2078 1142 2081 1148
rect 2086 1142 2089 1258
rect 2102 1192 2105 1258
rect 2150 1252 2153 1458
rect 2198 1442 2201 1448
rect 2214 1332 2217 1348
rect 2186 1288 2190 1291
rect 2178 1268 2182 1271
rect 2170 1258 2174 1261
rect 2182 1252 2185 1258
rect 2154 1248 2158 1251
rect 2098 1158 2102 1161
rect 2166 1151 2169 1158
rect 2074 1068 2078 1071
rect 1962 958 1966 961
rect 1982 952 1985 968
rect 1954 948 1958 951
rect 1994 948 1998 951
rect 1918 922 1921 938
rect 1912 903 1914 907
rect 1918 903 1921 907
rect 1925 903 1928 907
rect 1926 872 1929 888
rect 1974 872 1977 878
rect 1990 872 1993 948
rect 2002 938 2006 941
rect 2014 872 2017 978
rect 2026 958 2030 961
rect 2038 952 2041 958
rect 2046 952 2049 1058
rect 2078 1052 2081 1058
rect 2086 1051 2089 1118
rect 2102 1092 2105 1148
rect 2166 1082 2169 1128
rect 2098 1058 2102 1061
rect 2146 1058 2150 1061
rect 2086 1048 2094 1051
rect 2138 968 2142 971
rect 2022 942 2025 948
rect 2046 942 2049 948
rect 2082 947 2086 950
rect 2110 942 2113 948
rect 2174 942 2177 947
rect 1958 862 1961 868
rect 1854 758 1862 761
rect 1814 752 1817 758
rect 1822 752 1825 758
rect 1830 752 1833 758
rect 1854 752 1857 758
rect 1886 752 1889 818
rect 1926 781 1929 858
rect 1934 852 1937 858
rect 1958 842 1961 848
rect 1934 792 1937 828
rect 1926 778 1937 781
rect 1918 762 1921 768
rect 1934 752 1937 778
rect 1866 748 1870 751
rect 1750 742 1753 748
rect 1758 732 1761 738
rect 1766 712 1769 748
rect 1830 732 1833 738
rect 1606 698 1617 701
rect 1574 672 1577 678
rect 1590 672 1593 688
rect 1606 682 1609 688
rect 1562 668 1566 671
rect 1614 662 1617 698
rect 1650 688 1654 691
rect 1698 688 1702 691
rect 1638 672 1641 678
rect 1686 672 1689 688
rect 1674 668 1678 671
rect 1498 658 1502 661
rect 1478 592 1481 658
rect 1490 648 1494 651
rect 1622 622 1625 668
rect 1650 648 1654 651
rect 1638 642 1641 648
rect 1518 572 1521 618
rect 1606 602 1609 618
rect 1446 532 1449 538
rect 1454 522 1457 528
rect 1438 492 1441 518
rect 1462 492 1465 558
rect 1478 542 1481 548
rect 1486 542 1489 548
rect 1494 531 1497 558
rect 1550 552 1553 598
rect 1610 588 1614 591
rect 1614 542 1617 578
rect 1630 562 1633 628
rect 1662 592 1665 658
rect 1678 642 1681 658
rect 1710 652 1713 698
rect 1718 661 1721 698
rect 1774 672 1777 718
rect 1830 692 1833 698
rect 1838 692 1841 748
rect 1874 688 1878 691
rect 1854 672 1857 678
rect 1862 672 1865 678
rect 1730 668 1734 671
rect 1766 663 1769 668
rect 1718 658 1726 661
rect 1658 568 1662 571
rect 1630 552 1633 558
rect 1650 548 1654 551
rect 1742 551 1745 568
rect 1774 552 1777 668
rect 1886 662 1889 708
rect 1912 703 1914 707
rect 1918 703 1921 707
rect 1925 703 1928 707
rect 1830 648 1838 651
rect 1802 578 1806 581
rect 1486 528 1497 531
rect 1470 472 1473 478
rect 1478 472 1481 498
rect 1258 438 1262 441
rect 1326 392 1329 448
rect 1202 358 1209 361
rect 1134 352 1137 358
rect 1182 352 1185 358
rect 1082 348 1086 351
rect 1154 348 1158 351
rect 1110 342 1113 348
rect 1162 338 1166 341
rect 1038 278 1049 281
rect 958 272 961 278
rect 898 258 902 261
rect 846 252 849 258
rect 782 192 785 238
rect 798 192 801 208
rect 814 192 817 218
rect 822 142 825 178
rect 830 152 833 168
rect 854 162 857 168
rect 854 142 857 148
rect 674 138 681 141
rect 770 138 774 141
rect 794 138 798 141
rect 810 138 814 141
rect 430 122 433 138
rect 390 72 393 88
rect 430 72 433 118
rect 438 72 441 78
rect 458 68 462 71
rect 478 62 481 108
rect 486 72 489 98
rect 494 92 497 98
rect 590 92 593 118
rect 614 102 617 138
rect 686 132 689 138
rect 682 88 686 91
rect 526 62 529 88
rect 558 63 561 88
rect 646 72 649 78
rect 694 72 697 78
rect 718 72 721 128
rect 774 92 777 98
rect 790 92 793 138
rect 182 58 190 61
rect 726 62 729 78
rect 782 72 785 78
rect 798 72 801 118
rect 806 102 809 138
rect 886 132 889 138
rect 818 118 825 121
rect 814 62 817 78
rect 822 72 825 118
rect 880 103 882 107
rect 886 103 889 107
rect 893 103 896 107
rect 862 72 865 78
rect 902 72 905 178
rect 918 142 921 268
rect 974 252 977 268
rect 974 212 977 248
rect 998 222 1001 248
rect 998 192 1001 208
rect 1022 192 1025 268
rect 926 152 929 158
rect 982 132 985 168
rect 986 128 990 131
rect 942 92 945 118
rect 1030 102 1033 268
rect 1038 262 1041 278
rect 1046 262 1049 268
rect 1038 172 1041 258
rect 1054 252 1057 318
rect 1062 292 1065 338
rect 1110 322 1113 338
rect 1070 272 1073 318
rect 1142 302 1145 318
rect 1158 292 1161 318
rect 1146 288 1150 291
rect 1086 263 1089 268
rect 1118 252 1121 258
rect 1094 192 1097 198
rect 1038 152 1041 158
rect 1054 92 1057 138
rect 1050 88 1054 91
rect 870 62 873 68
rect 918 62 921 88
rect 934 62 937 68
rect 414 52 417 58
rect 478 52 481 58
rect 622 52 625 58
rect 458 48 462 51
rect 782 42 785 48
rect 376 3 378 7
rect 382 3 385 7
rect 389 3 392 7
rect 814 -18 817 58
rect 830 52 833 58
rect 174 -19 178 -18
rect 158 -22 178 -19
rect 814 -22 818 -18
rect 846 -19 849 58
rect 902 -18 905 58
rect 942 52 945 88
rect 958 72 961 88
rect 1062 82 1065 148
rect 1086 92 1089 178
rect 1102 152 1105 248
rect 1110 162 1113 168
rect 1134 152 1137 158
rect 1150 142 1153 188
rect 1166 162 1169 338
rect 1174 212 1177 338
rect 1198 222 1201 348
rect 1206 342 1209 358
rect 1246 352 1249 368
rect 1254 352 1257 358
rect 1302 352 1305 368
rect 1214 262 1217 288
rect 1182 192 1185 218
rect 1214 162 1217 238
rect 1158 152 1161 158
rect 1166 142 1169 148
rect 1190 142 1193 148
rect 1206 142 1209 158
rect 1214 152 1217 158
rect 1102 102 1105 138
rect 1190 92 1193 138
rect 1206 92 1209 138
rect 1222 82 1225 268
rect 1238 222 1241 348
rect 1254 292 1257 338
rect 1254 252 1257 268
rect 1262 192 1265 348
rect 1286 342 1289 348
rect 1270 272 1273 298
rect 1294 292 1297 348
rect 1310 342 1313 348
rect 1334 332 1337 348
rect 1342 342 1345 468
rect 1358 442 1361 468
rect 1394 458 1398 461
rect 1374 452 1377 458
rect 1392 403 1394 407
rect 1398 403 1401 407
rect 1405 403 1408 407
rect 1430 372 1433 468
rect 1486 462 1489 528
rect 1494 462 1497 468
rect 1450 448 1454 451
rect 1486 422 1489 458
rect 1502 452 1505 518
rect 1510 492 1513 538
rect 1574 532 1577 538
rect 1542 472 1545 528
rect 1594 488 1598 491
rect 1518 432 1521 468
rect 1606 462 1609 518
rect 1662 502 1665 538
rect 1670 532 1673 548
rect 1630 472 1633 498
rect 1534 452 1537 459
rect 1638 452 1641 458
rect 1418 368 1422 371
rect 1350 342 1353 368
rect 1394 358 1398 361
rect 1366 352 1369 358
rect 1394 348 1398 351
rect 1278 272 1281 278
rect 1342 272 1345 338
rect 1398 282 1401 338
rect 1430 312 1433 368
rect 1478 352 1481 358
rect 1454 342 1457 348
rect 1502 342 1505 428
rect 1534 392 1537 428
rect 1526 352 1529 388
rect 1542 352 1545 368
rect 1550 342 1553 398
rect 1574 392 1577 418
rect 1622 382 1625 418
rect 1522 338 1526 341
rect 1350 272 1353 278
rect 1342 252 1345 268
rect 1278 182 1281 188
rect 1310 162 1313 228
rect 1342 192 1345 218
rect 1350 182 1353 268
rect 1406 222 1409 228
rect 1234 158 1238 161
rect 1262 152 1265 158
rect 1290 138 1294 141
rect 1006 72 1009 78
rect 1142 72 1145 78
rect 990 52 993 59
rect 1094 12 1097 68
rect 1230 62 1233 118
rect 1254 112 1257 138
rect 1278 102 1281 118
rect 1286 92 1289 108
rect 1238 72 1241 78
rect 1294 62 1297 68
rect 1146 58 1150 61
rect 1302 51 1305 118
rect 1310 62 1313 158
rect 1358 152 1361 158
rect 1326 112 1329 148
rect 1350 142 1353 148
rect 1366 142 1369 148
rect 1350 102 1353 138
rect 1326 92 1329 98
rect 1318 72 1321 88
rect 1374 82 1377 218
rect 1392 203 1394 207
rect 1398 203 1401 207
rect 1405 203 1408 207
rect 1382 152 1385 158
rect 1422 152 1425 158
rect 1418 148 1422 151
rect 1430 142 1433 278
rect 1438 272 1441 288
rect 1454 252 1457 258
rect 1454 242 1457 248
rect 1462 192 1465 328
rect 1558 302 1561 348
rect 1590 332 1593 348
rect 1490 288 1494 291
rect 1474 258 1478 261
rect 1478 242 1481 248
rect 1486 242 1489 268
rect 1478 152 1481 228
rect 1486 192 1489 238
rect 1374 72 1377 78
rect 1298 48 1305 51
rect 1390 52 1393 59
rect 1406 52 1409 118
rect 1430 92 1433 138
rect 1438 92 1441 148
rect 1470 102 1473 148
rect 1494 142 1497 218
rect 1526 152 1529 268
rect 1534 222 1537 258
rect 1550 252 1553 258
rect 1574 192 1577 298
rect 1590 242 1593 268
rect 1598 262 1601 358
rect 1606 352 1609 378
rect 1634 368 1638 371
rect 1646 362 1649 368
rect 1618 358 1622 361
rect 1610 348 1617 351
rect 1614 342 1617 348
rect 1654 342 1657 498
rect 1678 492 1681 548
rect 1690 518 1694 521
rect 1702 482 1705 548
rect 1726 542 1729 548
rect 1822 542 1825 548
rect 1662 462 1665 468
rect 1726 462 1729 538
rect 1790 492 1793 528
rect 1830 492 1833 648
rect 1862 592 1865 638
rect 1838 552 1841 578
rect 1846 552 1849 558
rect 1790 462 1793 488
rect 1806 462 1809 468
rect 1814 462 1817 478
rect 1838 472 1841 548
rect 1854 542 1857 548
rect 1854 491 1857 538
rect 1878 532 1881 648
rect 1886 582 1889 658
rect 1902 622 1905 658
rect 1934 642 1937 748
rect 1958 732 1961 768
rect 1998 752 2001 788
rect 2022 771 2025 888
rect 2062 872 2065 938
rect 2158 932 2161 938
rect 2086 862 2089 898
rect 2138 868 2142 871
rect 2034 858 2038 861
rect 2078 852 2081 858
rect 2094 792 2097 818
rect 2022 768 2033 771
rect 2006 752 2009 758
rect 2022 752 2025 758
rect 1966 732 1969 748
rect 1974 742 1977 748
rect 1894 552 1897 598
rect 1902 562 1905 618
rect 1910 562 1913 608
rect 1934 602 1937 618
rect 1982 592 1985 738
rect 2014 732 2017 738
rect 2030 672 2033 768
rect 1998 652 2001 659
rect 2014 642 2017 668
rect 1998 592 2001 628
rect 2030 572 2033 668
rect 2038 662 2041 778
rect 2066 768 2070 771
rect 2046 702 2049 748
rect 1910 552 1913 558
rect 1946 548 1950 551
rect 1890 538 1894 541
rect 1912 503 1914 507
rect 1918 503 1921 507
rect 1925 503 1928 507
rect 1942 492 1945 538
rect 1950 502 1953 548
rect 1958 542 1961 568
rect 2010 548 2014 551
rect 2026 548 2030 551
rect 1854 488 1862 491
rect 1738 458 1742 461
rect 1666 448 1670 451
rect 1662 352 1665 448
rect 1686 392 1689 398
rect 1806 372 1809 458
rect 1678 362 1681 368
rect 1734 352 1737 368
rect 1746 358 1750 361
rect 1774 352 1777 358
rect 1786 348 1790 351
rect 1710 342 1713 348
rect 1798 341 1801 348
rect 1790 338 1801 341
rect 1822 342 1825 458
rect 1846 442 1849 458
rect 1838 382 1841 388
rect 1910 352 1913 358
rect 1606 302 1609 338
rect 1630 332 1633 338
rect 1682 328 1689 331
rect 1614 302 1617 318
rect 1622 272 1625 278
rect 1610 268 1614 271
rect 1630 262 1633 308
rect 1646 252 1649 268
rect 1654 252 1657 308
rect 1678 292 1681 318
rect 1686 312 1689 328
rect 1694 322 1697 328
rect 1666 268 1670 271
rect 1610 248 1614 251
rect 1438 82 1441 88
rect 1494 72 1497 138
rect 1534 72 1537 78
rect 1502 52 1505 59
rect 1550 52 1553 58
rect 1558 52 1561 68
rect 1574 62 1577 138
rect 1582 62 1585 118
rect 1590 72 1593 238
rect 1606 142 1609 218
rect 1678 172 1681 238
rect 1710 222 1713 258
rect 1614 152 1617 168
rect 1614 62 1617 68
rect 1570 58 1574 61
rect 1582 52 1585 58
rect 1622 52 1625 148
rect 1678 142 1681 168
rect 1686 151 1689 168
rect 1698 158 1702 161
rect 1686 148 1697 151
rect 1694 142 1697 148
rect 1710 122 1713 218
rect 1718 141 1721 328
rect 1734 322 1737 338
rect 1782 332 1785 338
rect 1758 312 1761 318
rect 1726 262 1729 308
rect 1774 292 1777 318
rect 1790 242 1793 338
rect 1830 322 1833 348
rect 1918 342 1921 468
rect 1926 463 1929 488
rect 1966 472 1969 548
rect 2026 528 2030 531
rect 2006 522 2009 528
rect 2014 492 2017 508
rect 2038 492 2041 658
rect 2046 652 2049 658
rect 2046 472 2049 548
rect 2054 512 2057 748
rect 2062 602 2065 668
rect 2102 662 2105 718
rect 2110 672 2113 728
rect 2118 692 2121 758
rect 2126 751 2129 758
rect 2142 742 2145 838
rect 2158 742 2161 768
rect 2174 762 2177 798
rect 2174 742 2177 748
rect 2182 722 2185 1248
rect 2206 1072 2209 1238
rect 2230 1152 2233 1438
rect 2238 1352 2241 1468
rect 2238 1272 2241 1348
rect 2242 1258 2246 1261
rect 2222 972 2225 1128
rect 2230 1062 2233 1138
rect 2238 962 2241 968
rect 2190 863 2193 888
rect 2206 872 2209 948
rect 2242 888 2246 891
rect 2222 872 2225 878
rect 2190 858 2193 859
rect 2206 842 2209 868
rect 2254 862 2257 1518
rect 2262 1482 2265 1528
rect 2270 1502 2273 1538
rect 2278 1452 2281 1548
rect 2294 1542 2297 1618
rect 2302 1542 2305 1738
rect 2286 1342 2289 1538
rect 2266 1318 2270 1321
rect 2286 1172 2289 1258
rect 2294 1242 2297 1418
rect 2302 1342 2305 1348
rect 2302 1242 2305 1248
rect 2282 1118 2286 1121
rect 2286 1092 2289 1098
rect 2286 1078 2294 1081
rect 2270 952 2273 968
rect 2262 942 2265 948
rect 2278 872 2281 898
rect 2286 892 2289 1078
rect 2298 968 2302 971
rect 2258 858 2262 861
rect 2238 852 2241 858
rect 2270 852 2273 868
rect 2198 752 2201 798
rect 2238 782 2241 848
rect 2270 792 2273 838
rect 2206 732 2209 738
rect 2214 732 2217 738
rect 2270 682 2273 698
rect 2286 692 2289 748
rect 2090 658 2094 661
rect 2078 652 2081 658
rect 2090 648 2094 651
rect 2062 552 2065 558
rect 2090 548 2094 551
rect 2070 482 2073 548
rect 2102 502 2105 628
rect 2110 622 2113 668
rect 2170 658 2174 661
rect 2246 652 2249 658
rect 2130 638 2134 641
rect 2134 552 2137 558
rect 2110 502 2113 548
rect 2142 542 2145 618
rect 2150 552 2153 588
rect 2158 558 2166 561
rect 2142 532 2145 538
rect 1966 462 1969 468
rect 2030 462 2033 468
rect 1926 458 1929 459
rect 1990 372 1993 418
rect 1982 352 1985 358
rect 1846 311 1849 328
rect 1858 318 1862 321
rect 1846 308 1857 311
rect 1814 262 1817 308
rect 1854 292 1857 308
rect 1912 303 1914 307
rect 1918 303 1921 307
rect 1925 303 1928 307
rect 1806 172 1809 258
rect 1866 188 1870 191
rect 1726 152 1729 158
rect 1718 138 1726 141
rect 1742 122 1745 138
rect 1646 92 1649 98
rect 1710 82 1713 118
rect 1766 102 1769 148
rect 1774 92 1777 168
rect 1870 152 1873 158
rect 1854 122 1857 128
rect 1826 118 1830 121
rect 1838 112 1841 118
rect 1814 72 1817 78
rect 1822 72 1825 108
rect 1830 92 1833 98
rect 1838 82 1841 88
rect 1854 82 1857 88
rect 1846 72 1849 78
rect 1878 72 1881 278
rect 1910 252 1913 259
rect 1934 172 1937 338
rect 1966 332 1969 338
rect 1966 302 1969 328
rect 1966 241 1969 268
rect 1974 262 1977 348
rect 1990 292 1993 358
rect 2006 352 2009 358
rect 1998 342 2001 348
rect 1998 272 2001 318
rect 2006 262 2009 268
rect 1982 252 1985 258
rect 1966 238 1974 241
rect 2014 202 2017 368
rect 2030 362 2033 368
rect 2022 322 2025 328
rect 2022 292 2025 308
rect 1894 142 1897 158
rect 2014 152 2017 198
rect 1886 122 1889 128
rect 1890 118 1894 121
rect 1912 103 1914 107
rect 1918 103 1921 107
rect 1925 103 1928 107
rect 1742 62 1745 68
rect 1698 58 1702 61
rect 1790 52 1793 58
rect 1618 48 1622 51
rect 1078 -18 1081 8
rect 1392 3 1394 7
rect 1398 3 1401 7
rect 1405 3 1408 7
rect 1614 -18 1617 8
rect 854 -19 858 -18
rect 846 -22 858 -19
rect 902 -22 906 -18
rect 1078 -22 1082 -18
rect 1614 -22 1618 -18
rect 1750 -19 1754 -18
rect 1758 -19 1761 38
rect 1750 -22 1761 -19
rect 1798 -18 1801 58
rect 1814 -18 1817 68
rect 1902 62 1905 78
rect 1934 72 1937 118
rect 1958 92 1961 148
rect 1974 62 1977 78
rect 1982 62 1985 128
rect 2022 102 2025 148
rect 1874 58 1878 61
rect 1938 58 1942 61
rect 1798 -22 1802 -18
rect 1814 -22 1818 -18
rect 1854 -19 1858 -18
rect 1862 -19 1865 58
rect 1894 42 1897 48
rect 1854 -22 1865 -19
rect 1926 -19 1929 58
rect 1934 -19 1938 -18
rect 1926 -22 1938 -19
rect 1982 -19 1986 -18
rect 1990 -19 1993 58
rect 2022 52 2025 59
rect 2030 52 2033 358
rect 2038 302 2041 468
rect 2046 342 2049 458
rect 2054 392 2057 478
rect 2086 472 2089 478
rect 2102 462 2105 498
rect 2118 472 2121 518
rect 2142 472 2145 518
rect 2134 462 2137 468
rect 2082 458 2086 461
rect 2070 442 2073 458
rect 2102 452 2105 458
rect 2118 351 2121 458
rect 2126 452 2129 458
rect 2150 451 2153 548
rect 2158 492 2161 558
rect 2170 548 2174 551
rect 2218 548 2222 551
rect 2254 542 2257 668
rect 2294 632 2297 848
rect 2302 742 2305 748
rect 2270 552 2273 558
rect 2290 538 2294 541
rect 2170 518 2174 521
rect 2198 492 2201 498
rect 2150 448 2158 451
rect 2158 362 2161 408
rect 2158 352 2161 358
rect 2166 352 2169 468
rect 2174 462 2177 488
rect 2254 472 2257 538
rect 2194 458 2198 461
rect 2178 358 2182 361
rect 2150 342 2153 348
rect 2182 342 2185 348
rect 2046 312 2049 338
rect 2038 272 2041 298
rect 2094 282 2097 288
rect 2066 268 2070 271
rect 2042 258 2046 261
rect 2070 252 2073 258
rect 2038 192 2041 238
rect 2078 142 2081 158
rect 2102 142 2105 148
rect 2110 142 2113 298
rect 2134 272 2137 338
rect 2190 292 2193 448
rect 2198 372 2201 438
rect 2198 342 2201 368
rect 2150 262 2153 268
rect 2150 152 2153 158
rect 2122 148 2126 151
rect 2062 112 2065 138
rect 2090 118 2094 121
rect 2094 92 2097 108
rect 2082 88 2086 91
rect 2134 62 2137 118
rect 2142 72 2145 118
rect 2158 82 2161 268
rect 2190 252 2193 258
rect 2174 142 2177 178
rect 2166 102 2169 138
rect 2198 92 2201 328
rect 2206 272 2209 468
rect 2242 458 2246 461
rect 2254 351 2257 468
rect 2250 348 2257 351
rect 2214 292 2217 308
rect 2246 272 2249 348
rect 2262 342 2265 348
rect 2302 332 2305 618
rect 2246 262 2249 268
rect 2206 72 2209 258
rect 2254 251 2257 328
rect 2270 262 2273 318
rect 2246 248 2257 251
rect 2246 142 2249 248
rect 2286 192 2289 218
rect 2258 158 2262 161
rect 2286 152 2289 158
rect 2294 142 2297 268
rect 2214 92 2217 98
rect 2174 62 2177 68
rect 2230 62 2233 118
rect 2270 62 2273 68
rect 2050 58 2054 61
rect 2250 58 2254 61
rect 2190 42 2193 48
rect 1982 -22 1993 -19
<< m3contact >>
rect 882 2103 886 2107
rect 889 2103 893 2107
rect 246 2088 250 2092
rect 606 2088 610 2092
rect 838 2088 842 2092
rect 318 2078 322 2082
rect 462 2078 466 2082
rect 822 2078 826 2082
rect 1518 2088 1522 2092
rect 1566 2088 1570 2092
rect 926 2078 930 2082
rect 1166 2078 1170 2082
rect 1206 2078 1210 2082
rect 1366 2078 1370 2082
rect 1382 2078 1386 2082
rect 1914 2103 1918 2107
rect 1921 2103 1925 2107
rect 1750 2078 1754 2082
rect 1846 2078 1850 2082
rect 1870 2078 1874 2082
rect 1886 2078 1890 2082
rect 486 2068 490 2072
rect 574 2068 578 2072
rect 974 2068 978 2072
rect 1110 2068 1114 2072
rect 1262 2068 1266 2072
rect 1294 2068 1298 2072
rect 1534 2068 1538 2072
rect 1814 2068 1818 2072
rect 2062 2068 2066 2072
rect 142 2058 146 2062
rect 158 2058 162 2062
rect 6 2048 10 2052
rect 78 2048 82 2052
rect 14 1978 18 1982
rect 230 2038 234 2042
rect 198 2018 202 2022
rect 134 1978 138 1982
rect 102 1968 106 1972
rect 158 1968 162 1972
rect 166 1968 170 1972
rect 222 1968 226 1972
rect 70 1958 74 1962
rect 126 1958 130 1962
rect 110 1948 114 1952
rect 62 1928 66 1932
rect 118 1918 122 1922
rect 238 2008 242 2012
rect 158 1948 162 1952
rect 230 1948 234 1952
rect 134 1868 138 1872
rect 166 1938 170 1942
rect 182 1918 186 1922
rect 190 1908 194 1912
rect 230 1898 234 1902
rect 198 1878 202 1882
rect 278 2058 282 2062
rect 302 2058 306 2062
rect 294 2048 298 2052
rect 334 2048 338 2052
rect 254 2038 258 2042
rect 334 2038 338 2042
rect 270 2028 274 2032
rect 262 1968 266 1972
rect 286 1948 290 1952
rect 246 1938 250 1942
rect 262 1938 266 1942
rect 318 1938 322 1942
rect 270 1918 274 1922
rect 262 1908 266 1912
rect 286 1908 290 1912
rect 326 1898 330 1902
rect 278 1878 282 1882
rect 430 2048 434 2052
rect 446 2048 450 2052
rect 390 2028 394 2032
rect 378 2003 382 2007
rect 385 2003 389 2007
rect 374 1968 378 1972
rect 454 1938 458 1942
rect 414 1928 418 1932
rect 638 2058 642 2062
rect 550 2048 554 2052
rect 550 2038 554 2042
rect 478 2018 482 2022
rect 494 1958 498 1962
rect 582 2048 586 2052
rect 566 1968 570 1972
rect 598 1958 602 1962
rect 654 2028 658 2032
rect 638 1968 642 1972
rect 510 1948 514 1952
rect 558 1948 562 1952
rect 582 1948 586 1952
rect 622 1948 626 1952
rect 510 1938 514 1942
rect 526 1938 530 1942
rect 574 1938 578 1942
rect 590 1938 594 1942
rect 598 1938 602 1942
rect 638 1938 642 1942
rect 462 1918 466 1922
rect 366 1908 370 1912
rect 54 1858 58 1862
rect 102 1858 106 1862
rect 110 1858 114 1862
rect 238 1858 242 1862
rect 110 1848 114 1852
rect 126 1848 130 1852
rect 134 1848 138 1852
rect 102 1838 106 1842
rect 134 1778 138 1782
rect 62 1748 66 1752
rect 110 1738 114 1742
rect 6 1708 10 1712
rect 262 1838 266 1842
rect 254 1748 258 1752
rect 222 1738 226 1742
rect 198 1728 202 1732
rect 174 1708 178 1712
rect 78 1668 82 1672
rect 102 1668 106 1672
rect 110 1668 114 1672
rect 174 1668 178 1672
rect 190 1668 194 1672
rect 182 1658 186 1662
rect 126 1648 130 1652
rect 158 1648 162 1652
rect 54 1618 58 1622
rect 86 1618 90 1622
rect 14 1568 18 1572
rect 6 1528 10 1532
rect 38 1548 42 1552
rect 62 1568 66 1572
rect 38 1538 42 1542
rect 78 1538 82 1542
rect 102 1538 106 1542
rect 46 1528 50 1532
rect 54 1498 58 1502
rect 94 1518 98 1522
rect 102 1488 106 1492
rect 86 1478 90 1482
rect 102 1478 106 1482
rect 38 1468 42 1472
rect 38 1338 42 1342
rect 30 1298 34 1302
rect 46 1278 50 1282
rect 30 1258 34 1262
rect 22 1238 26 1242
rect 6 1148 10 1152
rect 6 1088 10 1092
rect 30 1088 34 1092
rect 14 1078 18 1082
rect 22 1078 26 1082
rect 6 1038 10 1042
rect 78 1158 82 1162
rect 238 1678 242 1682
rect 294 1848 298 1852
rect 334 1798 338 1802
rect 358 1828 362 1832
rect 342 1788 346 1792
rect 350 1788 354 1792
rect 358 1768 362 1772
rect 334 1758 338 1762
rect 294 1748 298 1752
rect 350 1748 354 1752
rect 382 1868 386 1872
rect 398 1858 402 1862
rect 414 1818 418 1822
rect 430 1818 434 1822
rect 378 1803 382 1807
rect 385 1803 389 1807
rect 398 1778 402 1782
rect 270 1728 274 1732
rect 422 1788 426 1792
rect 478 1858 482 1862
rect 582 1928 586 1932
rect 494 1848 498 1852
rect 622 1918 626 1922
rect 582 1868 586 1872
rect 614 1868 618 1872
rect 542 1858 546 1862
rect 558 1858 562 1862
rect 526 1828 530 1832
rect 518 1808 522 1812
rect 566 1828 570 1832
rect 510 1798 514 1802
rect 550 1798 554 1802
rect 486 1748 490 1752
rect 326 1688 330 1692
rect 406 1688 410 1692
rect 278 1668 282 1672
rect 230 1618 234 1622
rect 182 1578 186 1582
rect 254 1578 258 1582
rect 174 1568 178 1572
rect 174 1558 178 1562
rect 118 1548 122 1552
rect 150 1538 154 1542
rect 254 1568 258 1572
rect 350 1658 354 1662
rect 326 1648 330 1652
rect 366 1648 370 1652
rect 326 1578 330 1582
rect 302 1558 306 1562
rect 118 1528 122 1532
rect 150 1488 154 1492
rect 110 1468 114 1472
rect 126 1458 130 1462
rect 110 1438 114 1442
rect 134 1438 138 1442
rect 118 1348 122 1352
rect 126 1338 130 1342
rect 150 1348 154 1352
rect 358 1528 362 1532
rect 198 1518 202 1522
rect 206 1518 210 1522
rect 318 1518 322 1522
rect 378 1603 382 1607
rect 385 1603 389 1607
rect 422 1678 426 1682
rect 430 1668 434 1672
rect 630 1858 634 1862
rect 590 1848 594 1852
rect 606 1848 610 1852
rect 598 1828 602 1832
rect 574 1768 578 1772
rect 590 1768 594 1772
rect 526 1758 530 1762
rect 574 1758 578 1762
rect 558 1748 562 1752
rect 542 1738 546 1742
rect 518 1718 522 1722
rect 534 1718 538 1722
rect 622 1848 626 1852
rect 646 1848 650 1852
rect 614 1798 618 1802
rect 598 1738 602 1742
rect 566 1708 570 1712
rect 582 1708 586 1712
rect 534 1678 538 1682
rect 526 1668 530 1672
rect 582 1668 586 1672
rect 590 1668 594 1672
rect 630 1758 634 1762
rect 622 1688 626 1692
rect 462 1658 466 1662
rect 518 1658 522 1662
rect 422 1608 426 1612
rect 414 1548 418 1552
rect 478 1648 482 1652
rect 542 1648 546 1652
rect 566 1648 570 1652
rect 446 1568 450 1572
rect 462 1568 466 1572
rect 438 1538 442 1542
rect 406 1508 410 1512
rect 238 1498 242 1502
rect 366 1498 370 1502
rect 390 1488 394 1492
rect 206 1478 210 1482
rect 230 1478 234 1482
rect 366 1478 370 1482
rect 310 1468 314 1472
rect 342 1468 346 1472
rect 358 1468 362 1472
rect 182 1458 186 1462
rect 174 1438 178 1442
rect 182 1438 186 1442
rect 134 1318 138 1322
rect 150 1308 154 1312
rect 102 1288 106 1292
rect 134 1288 138 1292
rect 118 1278 122 1282
rect 206 1458 210 1462
rect 254 1458 258 1462
rect 286 1458 290 1462
rect 222 1448 226 1452
rect 246 1448 250 1452
rect 262 1448 266 1452
rect 302 1448 306 1452
rect 278 1438 282 1442
rect 286 1438 290 1442
rect 262 1388 266 1392
rect 206 1358 210 1362
rect 310 1378 314 1382
rect 278 1368 282 1372
rect 270 1358 274 1362
rect 254 1348 258 1352
rect 294 1348 298 1352
rect 214 1338 218 1342
rect 254 1328 258 1332
rect 198 1278 202 1282
rect 238 1278 242 1282
rect 182 1268 186 1272
rect 198 1258 202 1262
rect 326 1378 330 1382
rect 422 1528 426 1532
rect 534 1588 538 1592
rect 550 1568 554 1572
rect 518 1548 522 1552
rect 478 1538 482 1542
rect 462 1528 466 1532
rect 462 1518 466 1522
rect 446 1488 450 1492
rect 478 1478 482 1482
rect 606 1648 610 1652
rect 686 2058 690 2062
rect 750 2058 754 2062
rect 670 2018 674 2022
rect 734 2008 738 2012
rect 774 2018 778 2022
rect 774 2008 778 2012
rect 886 2058 890 2062
rect 838 2018 842 2022
rect 822 1988 826 1992
rect 662 1958 666 1962
rect 790 1958 794 1962
rect 710 1948 714 1952
rect 726 1948 730 1952
rect 718 1938 722 1942
rect 662 1878 666 1882
rect 702 1878 706 1882
rect 694 1868 698 1872
rect 710 1868 714 1872
rect 686 1858 690 1862
rect 670 1838 674 1842
rect 662 1778 666 1782
rect 662 1758 666 1762
rect 678 1828 682 1832
rect 694 1798 698 1802
rect 686 1788 690 1792
rect 694 1778 698 1782
rect 702 1758 706 1762
rect 670 1738 674 1742
rect 686 1738 690 1742
rect 646 1678 650 1682
rect 662 1668 666 1672
rect 686 1678 690 1682
rect 758 1948 762 1952
rect 806 1938 810 1942
rect 742 1908 746 1912
rect 806 1898 810 1902
rect 806 1888 810 1892
rect 742 1868 746 1872
rect 750 1858 754 1862
rect 774 1858 778 1862
rect 766 1848 770 1852
rect 758 1838 762 1842
rect 822 1838 826 1842
rect 822 1798 826 1802
rect 822 1768 826 1772
rect 734 1728 738 1732
rect 766 1718 770 1722
rect 686 1658 690 1662
rect 702 1648 706 1652
rect 638 1628 642 1632
rect 614 1588 618 1592
rect 638 1588 642 1592
rect 614 1578 618 1582
rect 766 1698 770 1702
rect 734 1688 738 1692
rect 950 2059 954 2063
rect 1022 2058 1026 2062
rect 1054 2058 1058 2062
rect 902 2048 906 2052
rect 894 2038 898 2042
rect 862 2028 866 2032
rect 958 2008 962 2012
rect 878 1978 882 1982
rect 862 1968 866 1972
rect 846 1958 850 1962
rect 870 1958 874 1962
rect 902 1958 906 1962
rect 854 1948 858 1952
rect 854 1938 858 1942
rect 878 1918 882 1922
rect 882 1903 886 1907
rect 889 1903 893 1907
rect 942 1938 946 1942
rect 910 1898 914 1902
rect 1102 2048 1106 2052
rect 1134 2058 1138 2062
rect 1110 2038 1114 2042
rect 998 2028 1002 2032
rect 1086 2008 1090 2012
rect 1038 1968 1042 1972
rect 1062 1968 1066 1972
rect 1022 1958 1026 1962
rect 1022 1938 1026 1942
rect 1038 1928 1042 1932
rect 1046 1928 1050 1932
rect 1102 1938 1106 1942
rect 1054 1918 1058 1922
rect 1070 1918 1074 1922
rect 982 1908 986 1912
rect 998 1908 1002 1912
rect 1006 1898 1010 1902
rect 1046 1898 1050 1902
rect 1038 1878 1042 1882
rect 870 1858 874 1862
rect 918 1858 922 1862
rect 942 1858 946 1862
rect 990 1858 994 1862
rect 1014 1858 1018 1862
rect 838 1838 842 1842
rect 886 1828 890 1832
rect 870 1808 874 1812
rect 862 1758 866 1762
rect 886 1768 890 1772
rect 918 1838 922 1842
rect 950 1838 954 1842
rect 934 1798 938 1802
rect 982 1788 986 1792
rect 1014 1828 1018 1832
rect 998 1778 1002 1782
rect 926 1758 930 1762
rect 958 1758 962 1762
rect 878 1738 882 1742
rect 894 1738 898 1742
rect 934 1738 938 1742
rect 870 1718 874 1722
rect 882 1703 886 1707
rect 889 1703 893 1707
rect 830 1698 834 1702
rect 934 1698 938 1702
rect 854 1688 858 1692
rect 750 1668 754 1672
rect 734 1658 738 1662
rect 758 1638 762 1642
rect 750 1618 754 1622
rect 734 1598 738 1602
rect 638 1568 642 1572
rect 686 1568 690 1572
rect 718 1568 722 1572
rect 582 1558 586 1562
rect 654 1558 658 1562
rect 678 1558 682 1562
rect 654 1548 658 1552
rect 710 1538 714 1542
rect 518 1518 522 1522
rect 574 1518 578 1522
rect 454 1468 458 1472
rect 478 1458 482 1462
rect 430 1448 434 1452
rect 398 1438 402 1442
rect 446 1448 450 1452
rect 462 1448 466 1452
rect 438 1428 442 1432
rect 378 1403 382 1407
rect 385 1403 389 1407
rect 398 1398 402 1402
rect 398 1388 402 1392
rect 382 1378 386 1382
rect 342 1368 346 1372
rect 318 1358 322 1362
rect 334 1348 338 1352
rect 430 1378 434 1382
rect 398 1358 402 1362
rect 438 1358 442 1362
rect 406 1348 410 1352
rect 454 1348 458 1352
rect 390 1338 394 1342
rect 430 1338 434 1342
rect 446 1338 450 1342
rect 462 1338 466 1342
rect 286 1258 290 1262
rect 318 1258 322 1262
rect 94 1248 98 1252
rect 262 1248 266 1252
rect 246 1218 250 1222
rect 142 1178 146 1182
rect 230 1178 234 1182
rect 142 1168 146 1172
rect 174 1158 178 1162
rect 206 1158 210 1162
rect 166 1148 170 1152
rect 150 1138 154 1142
rect 174 1138 178 1142
rect 190 1138 194 1142
rect 86 1078 90 1082
rect 30 1068 34 1072
rect 38 1068 42 1072
rect 86 1068 90 1072
rect 46 1058 50 1062
rect 78 1048 82 1052
rect 94 1018 98 1022
rect 62 1008 66 1012
rect 14 958 18 962
rect 102 958 106 962
rect 62 948 66 952
rect 158 1078 162 1082
rect 150 1068 154 1072
rect 142 1028 146 1032
rect 126 958 130 962
rect 126 948 130 952
rect 150 948 154 952
rect 166 958 170 962
rect 110 938 114 942
rect 86 928 90 932
rect 142 928 146 932
rect 126 908 130 912
rect 118 888 122 892
rect 94 878 98 882
rect 54 858 58 862
rect 110 858 114 862
rect 46 768 50 772
rect 110 848 114 852
rect 102 838 106 842
rect 94 758 98 762
rect 110 778 114 782
rect 6 648 10 652
rect 6 638 10 642
rect 38 638 42 642
rect 70 568 74 572
rect 94 658 98 662
rect 110 718 114 722
rect 86 548 90 552
rect 30 538 34 542
rect 38 478 42 482
rect 62 418 66 422
rect 14 358 18 362
rect 22 358 26 362
rect 94 538 98 542
rect 102 468 106 472
rect 134 898 138 902
rect 134 878 138 882
rect 126 868 130 872
rect 142 848 146 852
rect 310 1228 314 1232
rect 294 1218 298 1222
rect 294 1168 298 1172
rect 310 1168 314 1172
rect 270 1158 274 1162
rect 254 1148 258 1152
rect 286 1148 290 1152
rect 230 1138 234 1142
rect 270 1138 274 1142
rect 198 1128 202 1132
rect 222 1118 226 1122
rect 254 1118 258 1122
rect 230 1088 234 1092
rect 262 1088 266 1092
rect 198 1078 202 1082
rect 190 1068 194 1072
rect 238 1068 242 1072
rect 222 1058 226 1062
rect 254 1058 258 1062
rect 206 1048 210 1052
rect 190 1038 194 1042
rect 230 1038 234 1042
rect 198 1018 202 1022
rect 190 958 194 962
rect 190 948 194 952
rect 166 888 170 892
rect 174 888 178 892
rect 166 878 170 882
rect 158 848 162 852
rect 150 838 154 842
rect 150 758 154 762
rect 190 778 194 782
rect 166 768 170 772
rect 190 768 194 772
rect 182 748 186 752
rect 134 718 138 722
rect 126 708 130 712
rect 134 678 138 682
rect 174 678 178 682
rect 134 658 138 662
rect 126 558 130 562
rect 206 968 210 972
rect 246 947 250 951
rect 246 938 250 942
rect 214 868 218 872
rect 206 858 210 862
rect 238 848 242 852
rect 262 918 266 922
rect 278 1038 282 1042
rect 430 1288 434 1292
rect 542 1498 546 1502
rect 534 1468 538 1472
rect 534 1458 538 1462
rect 950 1668 954 1672
rect 1094 1878 1098 1882
rect 1158 2048 1162 2052
rect 1142 2038 1146 2042
rect 1142 1998 1146 2002
rect 1118 1978 1122 1982
rect 1174 2058 1178 2062
rect 1206 2058 1210 2062
rect 1214 2048 1218 2052
rect 1230 2048 1234 2052
rect 1198 2038 1202 2042
rect 1214 2028 1218 2032
rect 1430 2058 1434 2062
rect 1462 2058 1466 2062
rect 1318 2038 1322 2042
rect 1334 2038 1338 2042
rect 1246 2008 1250 2012
rect 1286 2008 1290 2012
rect 1214 1968 1218 1972
rect 1270 1968 1274 1972
rect 1262 1958 1266 1962
rect 1206 1948 1210 1952
rect 1270 1948 1274 1952
rect 1166 1938 1170 1942
rect 1182 1938 1186 1942
rect 1158 1928 1162 1932
rect 1166 1918 1170 1922
rect 1142 1908 1146 1912
rect 1158 1908 1162 1912
rect 1158 1878 1162 1882
rect 1078 1848 1082 1852
rect 1086 1818 1090 1822
rect 1070 1778 1074 1782
rect 1086 1778 1090 1782
rect 1006 1738 1010 1742
rect 806 1658 810 1662
rect 910 1658 914 1662
rect 926 1658 930 1662
rect 974 1658 978 1662
rect 830 1638 834 1642
rect 782 1578 786 1582
rect 790 1558 794 1562
rect 854 1558 858 1562
rect 838 1548 842 1552
rect 862 1548 866 1552
rect 766 1538 770 1542
rect 846 1538 850 1542
rect 750 1528 754 1532
rect 798 1528 802 1532
rect 734 1508 738 1512
rect 702 1498 706 1502
rect 646 1488 650 1492
rect 702 1478 706 1482
rect 694 1468 698 1472
rect 542 1408 546 1412
rect 510 1378 514 1382
rect 510 1368 514 1372
rect 494 1348 498 1352
rect 486 1338 490 1342
rect 470 1318 474 1322
rect 366 1258 370 1262
rect 446 1258 450 1262
rect 446 1248 450 1252
rect 478 1308 482 1312
rect 478 1288 482 1292
rect 478 1278 482 1282
rect 486 1268 490 1272
rect 378 1203 382 1207
rect 385 1203 389 1207
rect 406 1178 410 1182
rect 374 1168 378 1172
rect 358 1158 362 1162
rect 414 1148 418 1152
rect 326 1138 330 1142
rect 406 1138 410 1142
rect 350 1128 354 1132
rect 294 1098 298 1102
rect 310 1078 314 1082
rect 430 1118 434 1122
rect 406 1068 410 1072
rect 470 1228 474 1232
rect 462 1178 466 1182
rect 470 1148 474 1152
rect 462 1138 466 1142
rect 510 1298 514 1302
rect 534 1278 538 1282
rect 510 1268 514 1272
rect 494 1228 498 1232
rect 486 1178 490 1182
rect 918 1638 922 1642
rect 982 1638 986 1642
rect 974 1618 978 1622
rect 950 1608 954 1612
rect 1014 1728 1018 1732
rect 1038 1728 1042 1732
rect 1030 1718 1034 1722
rect 1022 1708 1026 1712
rect 1006 1668 1010 1672
rect 998 1658 1002 1662
rect 998 1618 1002 1622
rect 982 1578 986 1582
rect 990 1578 994 1582
rect 1022 1638 1026 1642
rect 1046 1698 1050 1702
rect 1062 1688 1066 1692
rect 1038 1668 1042 1672
rect 1046 1658 1050 1662
rect 1014 1598 1018 1602
rect 1030 1598 1034 1602
rect 894 1558 898 1562
rect 958 1558 962 1562
rect 934 1548 938 1552
rect 1006 1548 1010 1552
rect 1038 1568 1042 1572
rect 982 1538 986 1542
rect 1022 1538 1026 1542
rect 894 1528 898 1532
rect 942 1528 946 1532
rect 998 1528 1002 1532
rect 1006 1528 1010 1532
rect 1054 1528 1058 1532
rect 846 1518 850 1522
rect 870 1518 874 1522
rect 910 1518 914 1522
rect 882 1503 886 1507
rect 889 1503 893 1507
rect 774 1478 778 1482
rect 806 1478 810 1482
rect 782 1468 786 1472
rect 598 1458 602 1462
rect 670 1458 674 1462
rect 694 1458 698 1462
rect 790 1458 794 1462
rect 646 1438 650 1442
rect 678 1438 682 1442
rect 654 1428 658 1432
rect 742 1438 746 1442
rect 750 1428 754 1432
rect 622 1358 626 1362
rect 718 1358 722 1362
rect 726 1358 730 1362
rect 758 1418 762 1422
rect 630 1348 634 1352
rect 646 1348 650 1352
rect 686 1348 690 1352
rect 726 1348 730 1352
rect 766 1398 770 1402
rect 790 1398 794 1402
rect 854 1458 858 1462
rect 870 1458 874 1462
rect 838 1448 842 1452
rect 910 1448 914 1452
rect 934 1448 938 1452
rect 838 1428 842 1432
rect 822 1418 826 1422
rect 814 1368 818 1372
rect 854 1358 858 1362
rect 782 1348 786 1352
rect 806 1348 810 1352
rect 846 1348 850 1352
rect 902 1348 906 1352
rect 574 1338 578 1342
rect 750 1338 754 1342
rect 798 1338 802 1342
rect 830 1338 834 1342
rect 566 1318 570 1322
rect 598 1318 602 1322
rect 550 1288 554 1292
rect 782 1328 786 1332
rect 822 1328 826 1332
rect 734 1318 738 1322
rect 750 1318 754 1322
rect 614 1308 618 1312
rect 662 1298 666 1302
rect 630 1278 634 1282
rect 638 1268 642 1272
rect 526 1258 530 1262
rect 542 1258 546 1262
rect 558 1258 562 1262
rect 598 1258 602 1262
rect 502 1178 506 1182
rect 510 1158 514 1162
rect 502 1138 506 1142
rect 486 1118 490 1122
rect 478 1108 482 1112
rect 486 1068 490 1072
rect 318 1058 322 1062
rect 286 988 290 992
rect 342 1008 346 1012
rect 398 1008 402 1012
rect 334 978 338 982
rect 294 968 298 972
rect 334 968 338 972
rect 378 1003 382 1007
rect 385 1003 389 1007
rect 350 958 354 962
rect 302 938 306 942
rect 318 938 322 942
rect 326 928 330 932
rect 310 898 314 902
rect 262 878 266 882
rect 270 878 274 882
rect 262 858 266 862
rect 262 848 266 852
rect 286 888 290 892
rect 270 838 274 842
rect 278 838 282 842
rect 326 859 330 863
rect 246 828 250 832
rect 270 828 274 832
rect 302 828 306 832
rect 206 788 210 792
rect 214 768 218 772
rect 254 768 258 772
rect 246 748 250 752
rect 214 668 218 672
rect 374 888 378 892
rect 406 968 410 972
rect 414 938 418 942
rect 406 918 410 922
rect 398 878 402 882
rect 438 1058 442 1062
rect 470 1018 474 1022
rect 438 998 442 1002
rect 438 988 442 992
rect 446 978 450 982
rect 470 948 474 952
rect 462 908 466 912
rect 438 898 442 902
rect 414 888 418 892
rect 430 888 434 892
rect 422 878 426 882
rect 534 1118 538 1122
rect 518 1098 522 1102
rect 526 1068 530 1072
rect 502 1038 506 1042
rect 526 998 530 1002
rect 518 968 522 972
rect 494 918 498 922
rect 518 908 522 912
rect 526 888 530 892
rect 542 968 546 972
rect 630 1248 634 1252
rect 590 1178 594 1182
rect 590 1168 594 1172
rect 614 1168 618 1172
rect 566 1148 570 1152
rect 574 1118 578 1122
rect 566 1098 570 1102
rect 622 1128 626 1132
rect 606 1098 610 1102
rect 590 1088 594 1092
rect 606 1068 610 1072
rect 646 1148 650 1152
rect 742 1288 746 1292
rect 766 1298 770 1302
rect 758 1278 762 1282
rect 790 1318 794 1322
rect 774 1268 778 1272
rect 882 1303 886 1307
rect 889 1303 893 1307
rect 814 1268 818 1272
rect 862 1268 866 1272
rect 686 1148 690 1152
rect 638 1128 642 1132
rect 670 1128 674 1132
rect 686 1128 690 1132
rect 646 1118 650 1122
rect 654 1098 658 1102
rect 614 1048 618 1052
rect 630 1048 634 1052
rect 606 1038 610 1042
rect 574 968 578 972
rect 542 948 546 952
rect 550 928 554 932
rect 550 918 554 922
rect 534 878 538 882
rect 390 848 394 852
rect 470 858 474 862
rect 478 838 482 842
rect 438 828 442 832
rect 422 818 426 822
rect 446 818 450 822
rect 378 803 382 807
rect 385 803 389 807
rect 310 788 314 792
rect 350 788 354 792
rect 462 788 466 792
rect 358 778 362 782
rect 262 748 266 752
rect 310 748 314 752
rect 342 748 346 752
rect 174 648 178 652
rect 166 598 170 602
rect 166 578 170 582
rect 150 548 154 552
rect 158 548 162 552
rect 150 538 154 542
rect 150 508 154 512
rect 126 488 130 492
rect 190 568 194 572
rect 190 548 194 552
rect 206 648 210 652
rect 206 558 210 562
rect 206 538 210 542
rect 198 528 202 532
rect 214 498 218 502
rect 158 478 162 482
rect 222 478 226 482
rect 142 468 146 472
rect 118 458 122 462
rect 134 458 138 462
rect 166 448 170 452
rect 142 438 146 442
rect 214 418 218 422
rect 182 358 186 362
rect 38 348 42 352
rect 62 348 66 352
rect 78 348 82 352
rect 134 348 138 352
rect 142 338 146 342
rect 70 308 74 312
rect 150 318 154 322
rect 174 308 178 312
rect 102 288 106 292
rect 126 288 130 292
rect 118 278 122 282
rect 38 268 42 272
rect 46 268 50 272
rect 30 258 34 262
rect 22 238 26 242
rect 94 248 98 252
rect 102 188 106 192
rect 110 168 114 172
rect 118 158 122 162
rect 142 158 146 162
rect 126 148 130 152
rect 102 128 106 132
rect 46 108 50 112
rect 14 88 18 92
rect 30 88 34 92
rect 46 68 50 72
rect 62 68 66 72
rect 6 58 10 62
rect 46 58 50 62
rect 46 48 50 52
rect 158 138 162 142
rect 302 738 306 742
rect 318 688 322 692
rect 310 668 314 672
rect 366 758 370 762
rect 422 758 426 762
rect 494 778 498 782
rect 510 768 514 772
rect 502 758 506 762
rect 430 748 434 752
rect 382 738 386 742
rect 398 728 402 732
rect 390 718 394 722
rect 422 738 426 742
rect 446 738 450 742
rect 486 738 490 742
rect 542 848 546 852
rect 542 758 546 762
rect 438 728 442 732
rect 406 718 410 722
rect 422 718 426 722
rect 358 688 362 692
rect 366 678 370 682
rect 350 668 354 672
rect 454 668 458 672
rect 318 658 322 662
rect 294 628 298 632
rect 374 638 378 642
rect 398 628 402 632
rect 378 603 382 607
rect 385 603 389 607
rect 342 578 346 582
rect 294 568 298 572
rect 302 568 306 572
rect 350 568 354 572
rect 270 548 274 552
rect 278 538 282 542
rect 286 528 290 532
rect 270 458 274 462
rect 302 488 306 492
rect 294 458 298 462
rect 294 418 298 422
rect 286 348 290 352
rect 190 328 194 332
rect 238 338 242 342
rect 262 338 266 342
rect 294 338 298 342
rect 270 328 274 332
rect 214 278 218 282
rect 238 278 242 282
rect 222 198 226 202
rect 214 158 218 162
rect 214 128 218 132
rect 126 88 130 92
rect 150 78 154 82
rect 110 48 114 52
rect 142 48 146 52
rect 294 318 298 322
rect 286 308 290 312
rect 326 538 330 542
rect 318 528 322 532
rect 326 508 330 512
rect 318 458 322 462
rect 334 458 338 462
rect 366 548 370 552
rect 406 548 410 552
rect 470 658 474 662
rect 422 648 426 652
rect 526 698 530 702
rect 534 648 538 652
rect 430 638 434 642
rect 470 628 474 632
rect 446 598 450 602
rect 430 588 434 592
rect 574 938 578 942
rect 558 878 562 882
rect 574 888 578 892
rect 622 948 626 952
rect 606 898 610 902
rect 638 1018 642 1022
rect 670 1058 674 1062
rect 694 1108 698 1112
rect 686 1028 690 1032
rect 686 1018 690 1022
rect 790 1248 794 1252
rect 822 1248 826 1252
rect 814 1238 818 1242
rect 742 1168 746 1172
rect 718 1158 722 1162
rect 830 1198 834 1202
rect 790 1158 794 1162
rect 798 1158 802 1162
rect 830 1158 834 1162
rect 782 1148 786 1152
rect 742 1118 746 1122
rect 742 1108 746 1112
rect 734 1068 738 1072
rect 734 1048 738 1052
rect 766 1128 770 1132
rect 782 1128 786 1132
rect 774 1118 778 1122
rect 806 1118 810 1122
rect 854 1078 858 1082
rect 782 1068 786 1072
rect 814 1068 818 1072
rect 886 1147 890 1151
rect 882 1103 886 1107
rect 889 1103 893 1107
rect 838 1058 842 1062
rect 758 1038 762 1042
rect 742 1008 746 1012
rect 750 1008 754 1012
rect 766 1018 770 1022
rect 758 998 762 1002
rect 694 978 698 982
rect 718 978 722 982
rect 638 968 642 972
rect 726 968 730 972
rect 694 948 698 952
rect 774 988 778 992
rect 774 968 778 972
rect 830 1038 834 1042
rect 862 1018 866 1022
rect 838 968 842 972
rect 806 958 810 962
rect 782 948 786 952
rect 806 938 810 942
rect 638 928 642 932
rect 694 928 698 932
rect 758 928 762 932
rect 630 888 634 892
rect 630 878 634 882
rect 686 888 690 892
rect 646 868 650 872
rect 678 868 682 872
rect 630 858 634 862
rect 638 858 642 862
rect 670 858 674 862
rect 566 838 570 842
rect 598 838 602 842
rect 574 758 578 762
rect 614 818 618 822
rect 638 818 642 822
rect 598 778 602 782
rect 614 768 618 772
rect 606 758 610 762
rect 598 748 602 752
rect 558 728 562 732
rect 558 708 562 712
rect 582 688 586 692
rect 590 688 594 692
rect 558 658 562 662
rect 662 788 666 792
rect 662 758 666 762
rect 622 748 626 752
rect 614 738 618 742
rect 662 738 666 742
rect 622 698 626 702
rect 638 698 642 702
rect 582 628 586 632
rect 550 578 554 582
rect 566 578 570 582
rect 430 568 434 572
rect 454 568 458 572
rect 502 568 506 572
rect 534 568 538 572
rect 414 528 418 532
rect 366 498 370 502
rect 350 448 354 452
rect 318 288 322 292
rect 310 278 314 282
rect 378 403 382 407
rect 385 403 389 407
rect 414 458 418 462
rect 454 558 458 562
rect 494 558 498 562
rect 462 548 466 552
rect 590 598 594 602
rect 518 548 522 552
rect 558 548 562 552
rect 598 558 602 562
rect 630 648 634 652
rect 774 908 778 912
rect 798 908 802 912
rect 766 848 770 852
rect 750 828 754 832
rect 742 758 746 762
rect 686 748 690 752
rect 694 748 698 752
rect 798 888 802 892
rect 686 738 690 742
rect 750 738 754 742
rect 758 738 762 742
rect 726 728 730 732
rect 678 718 682 722
rect 646 678 650 682
rect 646 668 650 672
rect 622 638 626 642
rect 686 688 690 692
rect 662 658 666 662
rect 654 568 658 572
rect 614 548 618 552
rect 670 648 674 652
rect 710 638 714 642
rect 702 608 706 612
rect 750 658 754 662
rect 734 648 738 652
rect 750 648 754 652
rect 774 678 778 682
rect 766 628 770 632
rect 830 878 834 882
rect 830 858 834 862
rect 822 768 826 772
rect 822 758 826 762
rect 854 958 858 962
rect 902 988 906 992
rect 894 948 898 952
rect 882 903 886 907
rect 889 903 893 907
rect 966 1498 970 1502
rect 1062 1508 1066 1512
rect 1046 1488 1050 1492
rect 1166 1798 1170 1802
rect 1118 1788 1122 1792
rect 1134 1758 1138 1762
rect 1150 1758 1154 1762
rect 1158 1758 1162 1762
rect 1102 1748 1106 1752
rect 1126 1748 1130 1752
rect 1182 1898 1186 1902
rect 1182 1858 1186 1862
rect 1190 1858 1194 1862
rect 1270 1928 1274 1932
rect 1214 1898 1218 1902
rect 1302 1968 1306 1972
rect 1270 1868 1274 1872
rect 1190 1738 1194 1742
rect 1142 1728 1146 1732
rect 1174 1728 1178 1732
rect 1190 1728 1194 1732
rect 1134 1708 1138 1712
rect 1110 1698 1114 1702
rect 1094 1618 1098 1622
rect 1086 1558 1090 1562
rect 1094 1558 1098 1562
rect 1158 1688 1162 1692
rect 1134 1678 1138 1682
rect 1110 1538 1114 1542
rect 1118 1538 1122 1542
rect 1142 1658 1146 1662
rect 1150 1658 1154 1662
rect 1166 1648 1170 1652
rect 1166 1548 1170 1552
rect 1206 1708 1210 1712
rect 1262 1858 1266 1862
rect 1222 1848 1226 1852
rect 1246 1768 1250 1772
rect 1318 1908 1322 1912
rect 1326 1888 1330 1892
rect 1302 1738 1306 1742
rect 1286 1698 1290 1702
rect 1238 1668 1242 1672
rect 1278 1668 1282 1672
rect 1302 1688 1306 1692
rect 1294 1668 1298 1672
rect 1390 2028 1394 2032
rect 1398 2018 1402 2022
rect 1394 2003 1398 2007
rect 1401 2003 1405 2007
rect 1350 1998 1354 2002
rect 1342 1978 1346 1982
rect 1342 1948 1346 1952
rect 1374 1968 1378 1972
rect 1406 1968 1410 1972
rect 1358 1958 1362 1962
rect 1390 1958 1394 1962
rect 1470 1958 1474 1962
rect 1390 1948 1394 1952
rect 1478 1948 1482 1952
rect 1390 1928 1394 1932
rect 1414 1908 1418 1912
rect 1438 1908 1442 1912
rect 1342 1848 1346 1852
rect 1318 1728 1322 1732
rect 1310 1678 1314 1682
rect 1214 1648 1218 1652
rect 1238 1648 1242 1652
rect 1246 1648 1250 1652
rect 1262 1648 1266 1652
rect 1206 1558 1210 1562
rect 1214 1558 1218 1562
rect 1190 1538 1194 1542
rect 1158 1518 1162 1522
rect 1318 1638 1322 1642
rect 1294 1628 1298 1632
rect 1270 1608 1274 1612
rect 1238 1598 1242 1602
rect 1230 1548 1234 1552
rect 1230 1518 1234 1522
rect 1142 1488 1146 1492
rect 1182 1478 1186 1482
rect 966 1468 970 1472
rect 1030 1468 1034 1472
rect 1014 1458 1018 1462
rect 1022 1458 1026 1462
rect 998 1448 1002 1452
rect 926 1428 930 1432
rect 926 1398 930 1402
rect 990 1428 994 1432
rect 998 1428 1002 1432
rect 974 1418 978 1422
rect 934 1388 938 1392
rect 942 1388 946 1392
rect 942 1368 946 1372
rect 942 1358 946 1362
rect 966 1348 970 1352
rect 950 1338 954 1342
rect 990 1348 994 1352
rect 974 1328 978 1332
rect 950 1308 954 1312
rect 990 1288 994 1292
rect 990 1268 994 1272
rect 1038 1458 1042 1462
rect 1094 1448 1098 1452
rect 1030 1438 1034 1442
rect 1038 1428 1042 1432
rect 1014 1368 1018 1372
rect 1030 1358 1034 1362
rect 1094 1438 1098 1442
rect 1054 1418 1058 1422
rect 1062 1358 1066 1362
rect 1022 1348 1026 1352
rect 1046 1348 1050 1352
rect 1054 1348 1058 1352
rect 1086 1348 1090 1352
rect 1014 1338 1018 1342
rect 1014 1268 1018 1272
rect 1006 1258 1010 1262
rect 966 1248 970 1252
rect 918 1238 922 1242
rect 1030 1268 1034 1272
rect 1038 1268 1042 1272
rect 998 1248 1002 1252
rect 1006 1248 1010 1252
rect 1038 1248 1042 1252
rect 974 1208 978 1212
rect 926 1198 930 1202
rect 926 1158 930 1162
rect 966 1148 970 1152
rect 1070 1328 1074 1332
rect 1062 1278 1066 1282
rect 1030 1238 1034 1242
rect 1046 1238 1050 1242
rect 1022 1198 1026 1202
rect 1014 1178 1018 1182
rect 1038 1168 1042 1172
rect 1022 1158 1026 1162
rect 1046 1158 1050 1162
rect 1054 1158 1058 1162
rect 1030 1148 1034 1152
rect 1038 1138 1042 1142
rect 958 1128 962 1132
rect 982 1128 986 1132
rect 942 1068 946 1072
rect 918 1048 922 1052
rect 942 1028 946 1032
rect 950 1018 954 1022
rect 1006 1118 1010 1122
rect 990 1108 994 1112
rect 982 1088 986 1092
rect 1030 1088 1034 1092
rect 990 1078 994 1082
rect 982 1058 986 1062
rect 998 1058 1002 1062
rect 998 1048 1002 1052
rect 1022 1048 1026 1052
rect 1006 1018 1010 1022
rect 974 998 978 1002
rect 958 978 962 982
rect 1062 1128 1066 1132
rect 1094 1278 1098 1282
rect 1086 1268 1090 1272
rect 1254 1518 1258 1522
rect 1174 1468 1178 1472
rect 1190 1468 1194 1472
rect 1262 1468 1266 1472
rect 1350 1698 1354 1702
rect 1366 1778 1370 1782
rect 1406 1878 1410 1882
rect 1470 1898 1474 1902
rect 1526 2048 1530 2052
rect 1550 2048 1554 2052
rect 1518 1958 1522 1962
rect 1518 1948 1522 1952
rect 1494 1878 1498 1882
rect 1526 1888 1530 1892
rect 1526 1868 1530 1872
rect 1398 1858 1402 1862
rect 1494 1858 1498 1862
rect 1510 1858 1514 1862
rect 1394 1803 1398 1807
rect 1401 1803 1405 1807
rect 1454 1848 1458 1852
rect 1470 1848 1474 1852
rect 1486 1848 1490 1852
rect 1462 1838 1466 1842
rect 1446 1788 1450 1792
rect 1430 1778 1434 1782
rect 1422 1758 1426 1762
rect 1478 1758 1482 1762
rect 1358 1668 1362 1672
rect 1326 1618 1330 1622
rect 1318 1558 1322 1562
rect 1286 1548 1290 1552
rect 1302 1548 1306 1552
rect 1382 1738 1386 1742
rect 1390 1738 1394 1742
rect 1566 2008 1570 2012
rect 1686 2058 1690 2062
rect 1670 2038 1674 2042
rect 1574 1998 1578 2002
rect 1734 2058 1738 2062
rect 1910 2058 1914 2062
rect 1966 2058 1970 2062
rect 1710 2048 1714 2052
rect 1726 2048 1730 2052
rect 1782 2048 1786 2052
rect 1766 2038 1770 2042
rect 1774 2018 1778 2022
rect 1702 1988 1706 1992
rect 1758 1988 1762 1992
rect 1606 1978 1610 1982
rect 1590 1968 1594 1972
rect 1606 1958 1610 1962
rect 1614 1958 1618 1962
rect 1646 1958 1650 1962
rect 1590 1948 1594 1952
rect 1558 1928 1562 1932
rect 1550 1808 1554 1812
rect 1550 1798 1554 1802
rect 1542 1748 1546 1752
rect 1534 1738 1538 1742
rect 1502 1698 1506 1702
rect 1462 1678 1466 1682
rect 1630 1948 1634 1952
rect 1702 1948 1706 1952
rect 1710 1938 1714 1942
rect 1574 1888 1578 1892
rect 1614 1888 1618 1892
rect 1638 1868 1642 1872
rect 1678 1868 1682 1872
rect 1766 1928 1770 1932
rect 1734 1878 1738 1882
rect 1766 1878 1770 1882
rect 1598 1858 1602 1862
rect 1614 1858 1618 1862
rect 1630 1858 1634 1862
rect 1582 1838 1586 1842
rect 1590 1808 1594 1812
rect 1654 1798 1658 1802
rect 1614 1788 1618 1792
rect 1630 1768 1634 1772
rect 1558 1748 1562 1752
rect 1582 1748 1586 1752
rect 1590 1748 1594 1752
rect 1614 1748 1618 1752
rect 1606 1738 1610 1742
rect 1662 1738 1666 1742
rect 1590 1718 1594 1722
rect 1574 1698 1578 1702
rect 1590 1678 1594 1682
rect 1662 1678 1666 1682
rect 1382 1668 1386 1672
rect 1446 1668 1450 1672
rect 1542 1668 1546 1672
rect 1566 1668 1570 1672
rect 1614 1668 1618 1672
rect 1398 1658 1402 1662
rect 1358 1648 1362 1652
rect 1374 1648 1378 1652
rect 1366 1618 1370 1622
rect 1394 1603 1398 1607
rect 1401 1603 1405 1607
rect 1758 1808 1762 1812
rect 1718 1768 1722 1772
rect 1766 1768 1770 1772
rect 1822 2008 1826 2012
rect 1806 1978 1810 1982
rect 1790 1948 1794 1952
rect 1790 1928 1794 1932
rect 1782 1878 1786 1882
rect 1814 1918 1818 1922
rect 1862 1998 1866 2002
rect 1846 1958 1850 1962
rect 1926 1958 1930 1962
rect 1966 1958 1970 1962
rect 1862 1948 1866 1952
rect 1894 1948 1898 1952
rect 1854 1938 1858 1942
rect 1886 1938 1890 1942
rect 1862 1918 1866 1922
rect 1830 1898 1834 1902
rect 1914 1903 1918 1907
rect 1921 1903 1925 1907
rect 1862 1898 1866 1902
rect 1838 1878 1842 1882
rect 1806 1868 1810 1872
rect 1830 1868 1834 1872
rect 1846 1868 1850 1872
rect 1782 1858 1786 1862
rect 1798 1858 1802 1862
rect 1726 1678 1730 1682
rect 1702 1668 1706 1672
rect 1526 1658 1530 1662
rect 1550 1658 1554 1662
rect 1574 1658 1578 1662
rect 1670 1658 1674 1662
rect 1438 1618 1442 1622
rect 1382 1578 1386 1582
rect 1422 1578 1426 1582
rect 1510 1568 1514 1572
rect 1358 1558 1362 1562
rect 1422 1558 1426 1562
rect 1454 1558 1458 1562
rect 1334 1538 1338 1542
rect 1342 1538 1346 1542
rect 1302 1528 1306 1532
rect 1390 1528 1394 1532
rect 1398 1528 1402 1532
rect 1390 1518 1394 1522
rect 1286 1478 1290 1482
rect 1318 1478 1322 1482
rect 1334 1478 1338 1482
rect 1366 1478 1370 1482
rect 1110 1428 1114 1432
rect 1126 1428 1130 1432
rect 1214 1458 1218 1462
rect 1238 1458 1242 1462
rect 1190 1448 1194 1452
rect 1230 1448 1234 1452
rect 1166 1438 1170 1442
rect 1206 1428 1210 1432
rect 1134 1418 1138 1422
rect 1174 1418 1178 1422
rect 1206 1408 1210 1412
rect 1134 1378 1138 1382
rect 1198 1378 1202 1382
rect 1230 1378 1234 1382
rect 1262 1458 1266 1462
rect 1302 1458 1306 1462
rect 1398 1508 1402 1512
rect 1454 1548 1458 1552
rect 1478 1548 1482 1552
rect 1486 1548 1490 1552
rect 1462 1528 1466 1532
rect 1486 1528 1490 1532
rect 1430 1518 1434 1522
rect 1446 1518 1450 1522
rect 1350 1468 1354 1472
rect 1398 1468 1402 1472
rect 1278 1448 1282 1452
rect 1302 1448 1306 1452
rect 1318 1448 1322 1452
rect 1358 1448 1362 1452
rect 1374 1438 1378 1442
rect 1270 1378 1274 1382
rect 1294 1378 1298 1382
rect 1214 1368 1218 1372
rect 1166 1358 1170 1362
rect 1198 1358 1202 1362
rect 1246 1358 1250 1362
rect 1150 1348 1154 1352
rect 1238 1348 1242 1352
rect 1278 1358 1282 1362
rect 1310 1368 1314 1372
rect 1326 1368 1330 1372
rect 1358 1368 1362 1372
rect 1270 1348 1274 1352
rect 1278 1348 1282 1352
rect 1350 1348 1354 1352
rect 1110 1338 1114 1342
rect 1134 1338 1138 1342
rect 1158 1338 1162 1342
rect 1190 1338 1194 1342
rect 1238 1338 1242 1342
rect 1254 1338 1258 1342
rect 1126 1318 1130 1322
rect 1158 1308 1162 1312
rect 1166 1308 1170 1312
rect 1118 1298 1122 1302
rect 1134 1298 1138 1302
rect 1150 1298 1154 1302
rect 1166 1278 1170 1282
rect 1214 1278 1218 1282
rect 1150 1268 1154 1272
rect 1174 1268 1178 1272
rect 1198 1268 1202 1272
rect 1182 1258 1186 1262
rect 1206 1258 1210 1262
rect 1110 1248 1114 1252
rect 1118 1248 1122 1252
rect 1142 1248 1146 1252
rect 1150 1248 1154 1252
rect 1174 1248 1178 1252
rect 1182 1248 1186 1252
rect 1102 1238 1106 1242
rect 1086 1218 1090 1222
rect 1102 1218 1106 1222
rect 1126 1218 1130 1222
rect 1078 1208 1082 1212
rect 1134 1198 1138 1202
rect 1158 1218 1162 1222
rect 1118 1178 1122 1182
rect 1134 1178 1138 1182
rect 1118 1168 1122 1172
rect 1086 1158 1090 1162
rect 1246 1328 1250 1332
rect 1286 1328 1290 1332
rect 1246 1318 1250 1322
rect 1238 1258 1242 1262
rect 1214 1248 1218 1252
rect 1198 1218 1202 1222
rect 1158 1168 1162 1172
rect 1190 1168 1194 1172
rect 1198 1158 1202 1162
rect 1246 1248 1250 1252
rect 1278 1288 1282 1292
rect 1366 1338 1370 1342
rect 1326 1318 1330 1322
rect 1294 1278 1298 1282
rect 1342 1278 1346 1282
rect 1246 1228 1250 1232
rect 1262 1228 1266 1232
rect 1262 1188 1266 1192
rect 1270 1178 1274 1182
rect 1230 1168 1234 1172
rect 1254 1168 1258 1172
rect 1142 1148 1146 1152
rect 1094 1128 1098 1132
rect 1102 1128 1106 1132
rect 1126 1128 1130 1132
rect 1054 1098 1058 1102
rect 1062 1098 1066 1102
rect 1062 1078 1066 1082
rect 1070 1008 1074 1012
rect 1022 988 1026 992
rect 1046 988 1050 992
rect 1014 978 1018 982
rect 910 968 914 972
rect 926 968 930 972
rect 1006 968 1010 972
rect 950 958 954 962
rect 910 948 914 952
rect 926 948 930 952
rect 902 868 906 872
rect 910 858 914 862
rect 934 888 938 892
rect 966 948 970 952
rect 990 948 994 952
rect 958 928 962 932
rect 982 928 986 932
rect 1046 968 1050 972
rect 1094 1088 1098 1092
rect 1078 998 1082 1002
rect 1086 978 1090 982
rect 1214 1148 1218 1152
rect 1278 1158 1282 1162
rect 1182 1138 1186 1142
rect 1214 1138 1218 1142
rect 1230 1138 1234 1142
rect 1166 1128 1170 1132
rect 1198 1128 1202 1132
rect 1150 1118 1154 1122
rect 1190 1118 1194 1122
rect 1182 1098 1186 1102
rect 1174 1068 1178 1072
rect 1118 1008 1122 1012
rect 1158 1038 1162 1042
rect 1166 1018 1170 1022
rect 1134 998 1138 1002
rect 1118 988 1122 992
rect 1134 988 1138 992
rect 1030 938 1034 942
rect 1094 938 1098 942
rect 1078 928 1082 932
rect 1014 918 1018 922
rect 1038 918 1042 922
rect 998 908 1002 912
rect 950 878 954 882
rect 1046 878 1050 882
rect 950 868 954 872
rect 982 868 986 872
rect 1014 868 1018 872
rect 1046 868 1050 872
rect 974 858 978 862
rect 854 848 858 852
rect 918 848 922 852
rect 958 848 962 852
rect 974 848 978 852
rect 942 838 946 842
rect 982 788 986 792
rect 998 788 1002 792
rect 934 768 938 772
rect 838 758 842 762
rect 854 758 858 762
rect 862 748 866 752
rect 950 748 954 752
rect 806 738 810 742
rect 830 728 834 732
rect 950 728 954 732
rect 870 718 874 722
rect 814 658 818 662
rect 726 598 730 602
rect 790 598 794 602
rect 806 598 810 602
rect 718 588 722 592
rect 790 588 794 592
rect 726 578 730 582
rect 462 538 466 542
rect 566 538 570 542
rect 646 538 650 542
rect 470 488 474 492
rect 518 488 522 492
rect 478 468 482 472
rect 502 468 506 472
rect 446 448 450 452
rect 406 388 410 392
rect 374 338 378 342
rect 398 288 402 292
rect 302 268 306 272
rect 334 268 338 272
rect 262 258 266 262
rect 270 248 274 252
rect 286 248 290 252
rect 230 188 234 192
rect 294 178 298 182
rect 294 158 298 162
rect 378 203 382 207
rect 385 203 389 207
rect 366 198 370 202
rect 494 458 498 462
rect 566 518 570 522
rect 558 448 562 452
rect 526 438 530 442
rect 534 428 538 432
rect 470 378 474 382
rect 422 368 426 372
rect 446 368 450 372
rect 510 358 514 362
rect 470 348 474 352
rect 502 348 506 352
rect 526 348 530 352
rect 470 338 474 342
rect 518 338 522 342
rect 502 328 506 332
rect 518 288 522 292
rect 422 268 426 272
rect 454 268 458 272
rect 510 268 514 272
rect 582 458 586 462
rect 622 458 626 462
rect 598 418 602 422
rect 622 418 626 422
rect 598 378 602 382
rect 566 348 570 352
rect 590 348 594 352
rect 582 338 586 342
rect 614 358 618 362
rect 622 358 626 362
rect 606 348 610 352
rect 702 458 706 462
rect 646 448 650 452
rect 710 438 714 442
rect 694 408 698 412
rect 774 558 778 562
rect 742 538 746 542
rect 782 538 786 542
rect 766 528 770 532
rect 734 478 738 482
rect 750 468 754 472
rect 814 538 818 542
rect 814 468 818 472
rect 774 448 778 452
rect 790 448 794 452
rect 806 448 810 452
rect 846 598 850 602
rect 822 438 826 442
rect 806 418 810 422
rect 766 398 770 402
rect 646 378 650 382
rect 726 368 730 372
rect 654 358 658 362
rect 854 538 858 542
rect 846 528 850 532
rect 838 398 842 402
rect 830 388 834 392
rect 638 348 642 352
rect 790 348 794 352
rect 806 348 810 352
rect 822 348 826 352
rect 614 328 618 332
rect 630 328 634 332
rect 614 298 618 302
rect 486 258 490 262
rect 502 258 506 262
rect 534 258 538 262
rect 518 248 522 252
rect 470 218 474 222
rect 438 188 442 192
rect 350 158 354 162
rect 398 158 402 162
rect 430 158 434 162
rect 294 148 298 152
rect 350 148 354 152
rect 342 118 346 122
rect 366 108 370 112
rect 358 88 362 92
rect 190 68 194 72
rect 350 68 354 72
rect 574 248 578 252
rect 558 238 562 242
rect 582 238 586 242
rect 542 188 546 192
rect 550 188 554 192
rect 582 148 586 152
rect 606 218 610 222
rect 710 338 714 342
rect 718 328 722 332
rect 750 328 754 332
rect 702 288 706 292
rect 758 268 762 272
rect 726 258 730 262
rect 670 238 674 242
rect 638 178 642 182
rect 598 148 602 152
rect 646 158 650 162
rect 670 158 674 162
rect 678 158 682 162
rect 718 158 722 162
rect 462 138 466 142
rect 558 138 562 142
rect 590 138 594 142
rect 806 318 810 322
rect 790 288 794 292
rect 814 268 818 272
rect 814 248 818 252
rect 838 298 842 302
rect 854 398 858 402
rect 882 703 886 707
rect 889 703 893 707
rect 878 668 882 672
rect 886 658 890 662
rect 958 678 962 682
rect 1086 918 1090 922
rect 1094 898 1098 902
rect 1094 788 1098 792
rect 1030 758 1034 762
rect 1102 758 1106 762
rect 1038 748 1042 752
rect 1006 738 1010 742
rect 1246 1088 1250 1092
rect 1262 1088 1266 1092
rect 1230 1068 1234 1072
rect 1222 1058 1226 1062
rect 1206 1048 1210 1052
rect 1206 1038 1210 1042
rect 1142 978 1146 982
rect 1158 978 1162 982
rect 1182 978 1186 982
rect 1190 978 1194 982
rect 1142 968 1146 972
rect 1158 958 1162 962
rect 1126 928 1130 932
rect 1126 838 1130 842
rect 1158 918 1162 922
rect 1142 888 1146 892
rect 1134 808 1138 812
rect 1078 748 1082 752
rect 1118 748 1122 752
rect 1054 738 1058 742
rect 1086 738 1090 742
rect 1046 728 1050 732
rect 1094 728 1098 732
rect 1094 718 1098 722
rect 1054 708 1058 712
rect 1046 688 1050 692
rect 1030 678 1034 682
rect 998 668 1002 672
rect 1014 668 1018 672
rect 982 658 986 662
rect 934 648 938 652
rect 910 628 914 632
rect 942 598 946 602
rect 1086 678 1090 682
rect 1038 658 1042 662
rect 1062 658 1066 662
rect 958 578 962 582
rect 966 578 970 582
rect 1022 578 1026 582
rect 1030 568 1034 572
rect 1046 568 1050 572
rect 1078 648 1082 652
rect 1086 638 1090 642
rect 1110 698 1114 702
rect 1150 748 1154 752
rect 1134 718 1138 722
rect 1134 698 1138 702
rect 1142 698 1146 702
rect 1126 668 1130 672
rect 1102 638 1106 642
rect 1094 628 1098 632
rect 1110 608 1114 612
rect 1078 568 1082 572
rect 1094 568 1098 572
rect 1126 658 1130 662
rect 1038 558 1042 562
rect 1054 558 1058 562
rect 1070 558 1074 562
rect 1118 558 1122 562
rect 894 538 898 542
rect 882 503 886 507
rect 889 503 893 507
rect 950 508 954 512
rect 942 498 946 502
rect 1014 498 1018 502
rect 998 488 1002 492
rect 950 478 954 482
rect 878 468 882 472
rect 974 468 978 472
rect 1030 468 1034 472
rect 966 458 970 462
rect 982 458 986 462
rect 902 438 906 442
rect 862 348 866 352
rect 894 348 898 352
rect 870 338 874 342
rect 882 303 886 307
rect 889 303 893 307
rect 990 438 994 442
rect 982 388 986 392
rect 958 368 962 372
rect 1118 548 1122 552
rect 1078 488 1082 492
rect 1086 488 1090 492
rect 1174 898 1178 902
rect 1174 888 1178 892
rect 1166 848 1170 852
rect 1302 1258 1306 1262
rect 1414 1418 1418 1422
rect 1438 1418 1442 1422
rect 1394 1403 1398 1407
rect 1401 1403 1405 1407
rect 1430 1368 1434 1372
rect 1406 1358 1410 1362
rect 1454 1508 1458 1512
rect 1478 1478 1482 1482
rect 1550 1648 1554 1652
rect 1542 1618 1546 1622
rect 1686 1648 1690 1652
rect 1718 1648 1722 1652
rect 1558 1638 1562 1642
rect 1678 1598 1682 1602
rect 1590 1568 1594 1572
rect 1702 1568 1706 1572
rect 1718 1568 1722 1572
rect 1566 1558 1570 1562
rect 1574 1558 1578 1562
rect 1606 1558 1610 1562
rect 1670 1558 1674 1562
rect 1598 1548 1602 1552
rect 1550 1538 1554 1542
rect 1534 1528 1538 1532
rect 1518 1518 1522 1522
rect 1494 1498 1498 1502
rect 1494 1478 1498 1482
rect 1462 1468 1466 1472
rect 1550 1508 1554 1512
rect 1574 1508 1578 1512
rect 1534 1488 1538 1492
rect 1542 1488 1546 1492
rect 1486 1458 1490 1462
rect 1502 1458 1506 1462
rect 1454 1448 1458 1452
rect 1494 1448 1498 1452
rect 1566 1448 1570 1452
rect 1534 1418 1538 1422
rect 1470 1408 1474 1412
rect 1446 1378 1450 1382
rect 1534 1398 1538 1402
rect 1446 1358 1450 1362
rect 1478 1358 1482 1362
rect 1390 1348 1394 1352
rect 1438 1348 1442 1352
rect 1382 1338 1386 1342
rect 1430 1328 1434 1332
rect 1438 1328 1442 1332
rect 1382 1308 1386 1312
rect 1422 1288 1426 1292
rect 1382 1278 1386 1282
rect 1358 1268 1362 1272
rect 1366 1248 1370 1252
rect 1350 1198 1354 1202
rect 1310 1148 1314 1152
rect 1294 1098 1298 1102
rect 1286 1078 1290 1082
rect 1310 1078 1314 1082
rect 1262 1068 1266 1072
rect 1262 1038 1266 1042
rect 1270 1008 1274 1012
rect 1294 1008 1298 1012
rect 1230 978 1234 982
rect 1222 968 1226 972
rect 1246 958 1250 962
rect 1286 958 1290 962
rect 1326 958 1330 962
rect 1278 948 1282 952
rect 1198 938 1202 942
rect 1214 938 1218 942
rect 1206 928 1210 932
rect 1214 888 1218 892
rect 1262 928 1266 932
rect 1302 918 1306 922
rect 1246 888 1250 892
rect 1254 888 1258 892
rect 1206 878 1210 882
rect 1238 878 1242 882
rect 1262 868 1266 872
rect 1182 768 1186 772
rect 1174 728 1178 732
rect 1158 678 1162 682
rect 1166 668 1170 672
rect 1206 758 1210 762
rect 1198 748 1202 752
rect 1238 748 1242 752
rect 1326 928 1330 932
rect 1318 918 1322 922
rect 1294 888 1298 892
rect 1318 888 1322 892
rect 1342 868 1346 872
rect 1270 788 1274 792
rect 1302 758 1306 762
rect 1358 1068 1362 1072
rect 1454 1308 1458 1312
rect 1454 1288 1458 1292
rect 1446 1278 1450 1282
rect 1438 1268 1442 1272
rect 1430 1258 1434 1262
rect 1390 1248 1394 1252
rect 1470 1328 1474 1332
rect 1494 1318 1498 1322
rect 1486 1298 1490 1302
rect 1526 1298 1530 1302
rect 1518 1278 1522 1282
rect 1470 1268 1474 1272
rect 1494 1258 1498 1262
rect 1414 1238 1418 1242
rect 1422 1238 1426 1242
rect 1478 1238 1482 1242
rect 1374 1208 1378 1212
rect 1394 1203 1398 1207
rect 1401 1203 1405 1207
rect 1374 1168 1378 1172
rect 1390 1128 1394 1132
rect 1374 1098 1378 1102
rect 1438 1218 1442 1222
rect 1462 1188 1466 1192
rect 1446 1168 1450 1172
rect 1438 1158 1442 1162
rect 1422 1148 1426 1152
rect 1462 1158 1466 1162
rect 1534 1198 1538 1202
rect 1526 1158 1530 1162
rect 1478 1148 1482 1152
rect 1494 1148 1498 1152
rect 1510 1148 1514 1152
rect 1486 1138 1490 1142
rect 1558 1368 1562 1372
rect 1558 1208 1562 1212
rect 1550 1178 1554 1182
rect 1558 1168 1562 1172
rect 1590 1468 1594 1472
rect 1582 1438 1586 1442
rect 1582 1358 1586 1362
rect 1710 1548 1714 1552
rect 1742 1698 1746 1702
rect 1758 1678 1762 1682
rect 1750 1648 1754 1652
rect 1734 1638 1738 1642
rect 1742 1628 1746 1632
rect 1742 1598 1746 1602
rect 1726 1538 1730 1542
rect 1638 1518 1642 1522
rect 1646 1498 1650 1502
rect 1638 1488 1642 1492
rect 1806 1738 1810 1742
rect 1798 1668 1802 1672
rect 1774 1648 1778 1652
rect 1790 1648 1794 1652
rect 1878 1878 1882 1882
rect 1942 1868 1946 1872
rect 1966 1868 1970 1872
rect 1870 1848 1874 1852
rect 1862 1838 1866 1842
rect 1822 1818 1826 1822
rect 1830 1788 1834 1792
rect 1854 1768 1858 1772
rect 1886 1818 1890 1822
rect 1934 1848 1938 1852
rect 1894 1758 1898 1762
rect 1830 1748 1834 1752
rect 1862 1748 1866 1752
rect 1878 1748 1882 1752
rect 1822 1678 1826 1682
rect 1814 1668 1818 1672
rect 1838 1728 1842 1732
rect 1846 1708 1850 1712
rect 1846 1658 1850 1662
rect 1774 1638 1778 1642
rect 1806 1638 1810 1642
rect 1894 1738 1898 1742
rect 1894 1728 1898 1732
rect 1886 1698 1890 1702
rect 1990 2058 1994 2062
rect 1990 1938 1994 1942
rect 2022 2048 2026 2052
rect 2078 2058 2082 2062
rect 2038 2048 2042 2052
rect 2070 2048 2074 2052
rect 2030 1988 2034 1992
rect 2014 1978 2018 1982
rect 2078 1978 2082 1982
rect 2046 1948 2050 1952
rect 2062 1948 2066 1952
rect 2046 1938 2050 1942
rect 2038 1878 2042 1882
rect 1998 1868 2002 1872
rect 2014 1868 2018 1872
rect 2046 1868 2050 1872
rect 2022 1858 2026 1862
rect 1982 1848 1986 1852
rect 1974 1828 1978 1832
rect 1942 1778 1946 1782
rect 2070 1898 2074 1902
rect 2078 1878 2082 1882
rect 2062 1838 2066 1842
rect 1990 1808 1994 1812
rect 1998 1788 2002 1792
rect 1950 1768 1954 1772
rect 1982 1768 1986 1772
rect 2046 1768 2050 1772
rect 1990 1758 1994 1762
rect 2150 2068 2154 2072
rect 2214 2068 2218 2072
rect 2238 2068 2242 2072
rect 2110 2058 2114 2062
rect 2102 2018 2106 2022
rect 2118 1958 2122 1962
rect 2238 2048 2242 2052
rect 2246 2048 2250 2052
rect 2262 2048 2266 2052
rect 2302 2048 2306 2052
rect 2166 1948 2170 1952
rect 2262 2018 2266 2022
rect 2246 1958 2250 1962
rect 2142 1938 2146 1942
rect 2174 1888 2178 1892
rect 2142 1868 2146 1872
rect 2102 1768 2106 1772
rect 2086 1758 2090 1762
rect 2102 1758 2106 1762
rect 1950 1748 1954 1752
rect 2070 1748 2074 1752
rect 1942 1738 1946 1742
rect 1934 1718 1938 1722
rect 1914 1703 1918 1707
rect 1921 1703 1925 1707
rect 1878 1668 1882 1672
rect 1838 1648 1842 1652
rect 1862 1648 1866 1652
rect 1838 1638 1842 1642
rect 1830 1588 1834 1592
rect 1806 1578 1810 1582
rect 1782 1568 1786 1572
rect 1862 1618 1866 1622
rect 1846 1568 1850 1572
rect 1806 1558 1810 1562
rect 1814 1548 1818 1552
rect 1838 1548 1842 1552
rect 1790 1538 1794 1542
rect 1814 1538 1818 1542
rect 1838 1538 1842 1542
rect 1750 1528 1754 1532
rect 1766 1528 1770 1532
rect 1758 1518 1762 1522
rect 1734 1508 1738 1512
rect 1726 1488 1730 1492
rect 1790 1498 1794 1502
rect 1782 1478 1786 1482
rect 1638 1468 1642 1472
rect 1702 1458 1706 1462
rect 1606 1448 1610 1452
rect 1766 1458 1770 1462
rect 1750 1448 1754 1452
rect 1766 1448 1770 1452
rect 1670 1418 1674 1422
rect 1718 1418 1722 1422
rect 1742 1418 1746 1422
rect 1638 1378 1642 1382
rect 1582 1328 1586 1332
rect 1606 1338 1610 1342
rect 1630 1338 1634 1342
rect 1646 1338 1650 1342
rect 1598 1308 1602 1312
rect 1590 1298 1594 1302
rect 1590 1268 1594 1272
rect 1638 1308 1642 1312
rect 1630 1268 1634 1272
rect 1670 1338 1674 1342
rect 1686 1338 1690 1342
rect 1702 1328 1706 1332
rect 1710 1318 1714 1322
rect 1670 1308 1674 1312
rect 1654 1298 1658 1302
rect 1694 1298 1698 1302
rect 1726 1368 1730 1372
rect 1734 1348 1738 1352
rect 1734 1328 1738 1332
rect 1742 1328 1746 1332
rect 1654 1268 1658 1272
rect 1742 1268 1746 1272
rect 1790 1438 1794 1442
rect 1782 1358 1786 1362
rect 1766 1348 1770 1352
rect 1798 1368 1802 1372
rect 1806 1348 1810 1352
rect 1766 1338 1770 1342
rect 1790 1278 1794 1282
rect 1774 1268 1778 1272
rect 1622 1258 1626 1262
rect 1686 1258 1690 1262
rect 1606 1248 1610 1252
rect 1686 1248 1690 1252
rect 1710 1248 1714 1252
rect 1654 1238 1658 1242
rect 1670 1238 1674 1242
rect 1622 1198 1626 1202
rect 1646 1188 1650 1192
rect 1598 1158 1602 1162
rect 1638 1158 1642 1162
rect 1590 1148 1594 1152
rect 1558 1138 1562 1142
rect 1670 1158 1674 1162
rect 1654 1148 1658 1152
rect 1638 1138 1642 1142
rect 1670 1138 1674 1142
rect 1574 1128 1578 1132
rect 1486 1118 1490 1122
rect 1550 1118 1554 1122
rect 1470 1098 1474 1102
rect 1414 1088 1418 1092
rect 1494 1108 1498 1112
rect 1518 1108 1522 1112
rect 1542 1108 1546 1112
rect 1390 1078 1394 1082
rect 1486 1078 1490 1082
rect 1502 1098 1506 1102
rect 1374 1048 1378 1052
rect 1414 1048 1418 1052
rect 1374 1038 1378 1042
rect 1358 1028 1362 1032
rect 1394 1003 1398 1007
rect 1401 1003 1405 1007
rect 1454 1058 1458 1062
rect 1470 1058 1474 1062
rect 1454 1048 1458 1052
rect 1438 1038 1442 1042
rect 1494 1008 1498 1012
rect 1438 978 1442 982
rect 1422 958 1426 962
rect 1430 948 1434 952
rect 1470 948 1474 952
rect 1358 918 1362 922
rect 1478 898 1482 902
rect 1406 888 1410 892
rect 1470 888 1474 892
rect 1470 878 1474 882
rect 1374 868 1378 872
rect 1446 868 1450 872
rect 1438 858 1442 862
rect 1454 858 1458 862
rect 1518 1088 1522 1092
rect 1614 1128 1618 1132
rect 1582 1088 1586 1092
rect 1566 1068 1570 1072
rect 1590 1068 1594 1072
rect 1550 1058 1554 1062
rect 1582 1058 1586 1062
rect 1526 1048 1530 1052
rect 1534 1048 1538 1052
rect 1518 1028 1522 1032
rect 1510 988 1514 992
rect 1550 968 1554 972
rect 1574 1038 1578 1042
rect 1590 1038 1594 1042
rect 1582 1008 1586 1012
rect 1566 958 1570 962
rect 1518 948 1522 952
rect 1518 908 1522 912
rect 1494 898 1498 902
rect 1494 888 1498 892
rect 1534 888 1538 892
rect 1526 868 1530 872
rect 1394 803 1398 807
rect 1401 803 1405 807
rect 1446 788 1450 792
rect 1430 778 1434 782
rect 1366 758 1370 762
rect 1438 758 1442 762
rect 1350 748 1354 752
rect 1382 748 1386 752
rect 1190 738 1194 742
rect 1230 738 1234 742
rect 1198 678 1202 682
rect 1254 708 1258 712
rect 1294 698 1298 702
rect 1278 678 1282 682
rect 1214 668 1218 672
rect 1230 668 1234 672
rect 1158 658 1162 662
rect 1182 658 1186 662
rect 1166 598 1170 602
rect 1158 588 1162 592
rect 1158 578 1162 582
rect 1174 568 1178 572
rect 1134 478 1138 482
rect 1062 458 1066 462
rect 1038 428 1042 432
rect 1046 388 1050 392
rect 1030 378 1034 382
rect 1014 358 1018 362
rect 1038 358 1042 362
rect 990 348 994 352
rect 1030 338 1034 342
rect 1006 328 1010 332
rect 910 318 914 322
rect 974 318 978 322
rect 974 308 978 312
rect 998 298 1002 302
rect 1014 288 1018 292
rect 958 278 962 282
rect 1094 448 1098 452
rect 1182 538 1186 542
rect 1126 448 1130 452
rect 1102 438 1106 442
rect 1134 428 1138 432
rect 1150 398 1154 402
rect 1174 448 1178 452
rect 1222 638 1226 642
rect 1286 668 1290 672
rect 1278 648 1282 652
rect 1342 738 1346 742
rect 1414 738 1418 742
rect 1350 718 1354 722
rect 1398 718 1402 722
rect 1430 708 1434 712
rect 1422 678 1426 682
rect 1334 658 1338 662
rect 1222 628 1226 632
rect 1262 628 1266 632
rect 1454 778 1458 782
rect 1478 768 1482 772
rect 1486 758 1490 762
rect 1510 758 1514 762
rect 1550 878 1554 882
rect 1622 1078 1626 1082
rect 1654 1128 1658 1132
rect 1686 1128 1690 1132
rect 1678 1118 1682 1122
rect 1678 1088 1682 1092
rect 1638 1068 1642 1072
rect 1670 1068 1674 1072
rect 1678 1068 1682 1072
rect 1630 1058 1634 1062
rect 1646 1058 1650 1062
rect 1638 1048 1642 1052
rect 1614 1008 1618 1012
rect 1606 918 1610 922
rect 1630 918 1634 922
rect 1630 908 1634 912
rect 1614 888 1618 892
rect 1574 878 1578 882
rect 1558 868 1562 872
rect 1574 868 1578 872
rect 1534 848 1538 852
rect 1542 848 1546 852
rect 1510 748 1514 752
rect 1518 748 1522 752
rect 1470 728 1474 732
rect 1510 718 1514 722
rect 1502 688 1506 692
rect 1414 658 1418 662
rect 1462 658 1466 662
rect 1414 648 1418 652
rect 1326 588 1330 592
rect 1206 578 1210 582
rect 1214 578 1218 582
rect 1238 568 1242 572
rect 1294 568 1298 572
rect 1318 568 1322 572
rect 1326 568 1330 572
rect 1206 558 1210 562
rect 1246 558 1250 562
rect 1190 508 1194 512
rect 1230 518 1234 522
rect 1206 438 1210 442
rect 1214 428 1218 432
rect 1166 388 1170 392
rect 1102 378 1106 382
rect 1070 358 1074 362
rect 1134 368 1138 372
rect 1262 538 1266 542
rect 1270 538 1274 542
rect 1302 538 1306 542
rect 1254 528 1258 532
rect 1326 518 1330 522
rect 1382 608 1386 612
rect 1394 603 1398 607
rect 1401 603 1405 607
rect 1446 638 1450 642
rect 1422 578 1426 582
rect 1358 568 1362 572
rect 1350 558 1354 562
rect 1342 538 1346 542
rect 1366 538 1370 542
rect 1382 538 1386 542
rect 1438 558 1442 562
rect 1430 528 1434 532
rect 1278 498 1282 502
rect 1318 488 1322 492
rect 1254 478 1258 482
rect 1406 498 1410 502
rect 1374 488 1378 492
rect 1534 738 1538 742
rect 1558 738 1562 742
rect 1534 718 1538 722
rect 1518 698 1522 702
rect 1590 868 1594 872
rect 1622 848 1626 852
rect 1662 978 1666 982
rect 1710 1098 1714 1102
rect 1694 1088 1698 1092
rect 1750 1228 1754 1232
rect 1774 1228 1778 1232
rect 1726 1048 1730 1052
rect 1758 1148 1762 1152
rect 1750 1138 1754 1142
rect 1798 1128 1802 1132
rect 1782 1118 1786 1122
rect 1766 1078 1770 1082
rect 1806 1078 1810 1082
rect 1742 1048 1746 1052
rect 1734 1008 1738 1012
rect 1846 1358 1850 1362
rect 1822 1348 1826 1352
rect 2006 1738 2010 1742
rect 1966 1718 1970 1722
rect 1974 1718 1978 1722
rect 2006 1718 2010 1722
rect 1974 1668 1978 1672
rect 1990 1658 1994 1662
rect 1950 1638 1954 1642
rect 1998 1648 2002 1652
rect 2014 1688 2018 1692
rect 2030 1668 2034 1672
rect 2014 1648 2018 1652
rect 1990 1638 1994 1642
rect 2006 1638 2010 1642
rect 2022 1568 2026 1572
rect 1966 1558 1970 1562
rect 2190 1858 2194 1862
rect 2190 1838 2194 1842
rect 2182 1818 2186 1822
rect 2150 1778 2154 1782
rect 2150 1748 2154 1752
rect 2118 1738 2122 1742
rect 2086 1728 2090 1732
rect 2110 1728 2114 1732
rect 2078 1678 2082 1682
rect 2190 1728 2194 1732
rect 2134 1698 2138 1702
rect 2126 1648 2130 1652
rect 2126 1568 2130 1572
rect 1990 1548 1994 1552
rect 2094 1548 2098 1552
rect 2110 1548 2114 1552
rect 1902 1538 1906 1542
rect 1914 1503 1918 1507
rect 1921 1503 1925 1507
rect 1958 1528 1962 1532
rect 1878 1488 1882 1492
rect 1894 1488 1898 1492
rect 1942 1488 1946 1492
rect 1950 1488 1954 1492
rect 1894 1478 1898 1482
rect 1878 1368 1882 1372
rect 1830 1338 1834 1342
rect 1830 1288 1834 1292
rect 1838 1268 1842 1272
rect 1854 1248 1858 1252
rect 1838 1238 1842 1242
rect 1830 1148 1834 1152
rect 1942 1458 1946 1462
rect 1902 1448 1906 1452
rect 1942 1448 1946 1452
rect 1926 1358 1930 1362
rect 2054 1538 2058 1542
rect 2070 1538 2074 1542
rect 2006 1528 2010 1532
rect 2030 1528 2034 1532
rect 1982 1508 1986 1512
rect 1990 1488 1994 1492
rect 2006 1488 2010 1492
rect 2054 1498 2058 1502
rect 2070 1488 2074 1492
rect 2046 1478 2050 1482
rect 1990 1468 1994 1472
rect 2022 1468 2026 1472
rect 2070 1458 2074 1462
rect 1998 1408 2002 1412
rect 1974 1368 1978 1372
rect 1982 1368 1986 1372
rect 2030 1368 2034 1372
rect 2006 1358 2010 1362
rect 1894 1328 1898 1332
rect 1942 1328 1946 1332
rect 1934 1318 1938 1322
rect 1914 1303 1918 1307
rect 1921 1303 1925 1307
rect 1878 1278 1882 1282
rect 1894 1278 1898 1282
rect 1958 1308 1962 1312
rect 1966 1268 1970 1272
rect 2166 1698 2170 1702
rect 2158 1678 2162 1682
rect 2174 1658 2178 1662
rect 2206 1908 2210 1912
rect 2214 1898 2218 1902
rect 2230 1898 2234 1902
rect 2222 1868 2226 1872
rect 2270 1868 2274 1872
rect 2214 1838 2218 1842
rect 2254 1848 2258 1852
rect 2270 1848 2274 1852
rect 2206 1808 2210 1812
rect 2222 1808 2226 1812
rect 2254 1778 2258 1782
rect 2214 1748 2218 1752
rect 2302 1818 2306 1822
rect 2262 1758 2266 1762
rect 2294 1758 2298 1762
rect 2278 1748 2282 1752
rect 2206 1738 2210 1742
rect 2230 1668 2234 1672
rect 2198 1658 2202 1662
rect 2182 1648 2186 1652
rect 2166 1578 2170 1582
rect 2166 1568 2170 1572
rect 2142 1548 2146 1552
rect 2158 1548 2162 1552
rect 2150 1518 2154 1522
rect 2174 1538 2178 1542
rect 2238 1648 2242 1652
rect 2278 1648 2282 1652
rect 2262 1568 2266 1572
rect 2214 1558 2218 1562
rect 2222 1558 2226 1562
rect 2214 1548 2218 1552
rect 2246 1548 2250 1552
rect 2206 1538 2210 1542
rect 2198 1518 2202 1522
rect 2262 1528 2266 1532
rect 2254 1518 2258 1522
rect 2230 1468 2234 1472
rect 2150 1458 2154 1462
rect 2174 1458 2178 1462
rect 2190 1458 2194 1462
rect 2110 1388 2114 1392
rect 2078 1368 2082 1372
rect 2062 1358 2066 1362
rect 2078 1358 2082 1362
rect 2046 1348 2050 1352
rect 2062 1348 2066 1352
rect 2078 1348 2082 1352
rect 2142 1358 2146 1362
rect 2014 1328 2018 1332
rect 2038 1328 2042 1332
rect 1998 1298 2002 1302
rect 2070 1318 2074 1322
rect 2030 1288 2034 1292
rect 2006 1278 2010 1282
rect 1902 1258 1906 1262
rect 1894 1238 1898 1242
rect 1886 1218 1890 1222
rect 1862 1198 1866 1202
rect 1846 1178 1850 1182
rect 1886 1168 1890 1172
rect 1926 1168 1930 1172
rect 1862 1148 1866 1152
rect 1878 1148 1882 1152
rect 1854 1138 1858 1142
rect 1838 1118 1842 1122
rect 1838 1108 1842 1112
rect 1918 1118 1922 1122
rect 1914 1103 1918 1107
rect 1921 1103 1925 1107
rect 1862 1098 1866 1102
rect 1782 1068 1786 1072
rect 1814 1068 1818 1072
rect 1870 1068 1874 1072
rect 1894 1068 1898 1072
rect 1798 1058 1802 1062
rect 1814 1058 1818 1062
rect 1830 1058 1834 1062
rect 1806 1048 1810 1052
rect 1758 978 1762 982
rect 1742 968 1746 972
rect 1686 958 1690 962
rect 1654 908 1658 912
rect 1670 908 1674 912
rect 1694 908 1698 912
rect 1662 888 1666 892
rect 1654 878 1658 882
rect 1814 968 1818 972
rect 1806 948 1810 952
rect 1830 948 1834 952
rect 1790 938 1794 942
rect 1830 918 1834 922
rect 1798 898 1802 902
rect 1894 1058 1898 1062
rect 1862 1048 1866 1052
rect 1870 1048 1874 1052
rect 1870 948 1874 952
rect 1902 1048 1906 1052
rect 1902 988 1906 992
rect 1854 938 1858 942
rect 1870 938 1874 942
rect 1838 898 1842 902
rect 1694 878 1698 882
rect 1766 878 1770 882
rect 1790 878 1794 882
rect 1838 878 1842 882
rect 1686 868 1690 872
rect 1718 868 1722 872
rect 1790 858 1794 862
rect 1806 858 1810 862
rect 1662 848 1666 852
rect 1686 848 1690 852
rect 1598 838 1602 842
rect 1638 838 1642 842
rect 1670 838 1674 842
rect 1638 808 1642 812
rect 1598 738 1602 742
rect 1558 718 1562 722
rect 1582 708 1586 712
rect 1654 718 1658 722
rect 1750 848 1754 852
rect 1718 838 1722 842
rect 1726 838 1730 842
rect 1734 768 1738 772
rect 1726 758 1730 762
rect 1798 848 1802 852
rect 1838 858 1842 862
rect 1766 838 1770 842
rect 1782 818 1786 822
rect 1870 848 1874 852
rect 1862 838 1866 842
rect 1854 828 1858 832
rect 1830 808 1834 812
rect 1798 768 1802 772
rect 1846 768 1850 772
rect 1894 898 1898 902
rect 1894 878 1898 882
rect 1918 958 1922 962
rect 1958 1158 1962 1162
rect 2086 1308 2090 1312
rect 2134 1288 2138 1292
rect 2110 1278 2114 1282
rect 1990 1258 1994 1262
rect 2030 1258 2034 1262
rect 2046 1258 2050 1262
rect 2078 1258 2082 1262
rect 2102 1258 2106 1262
rect 1982 1248 1986 1252
rect 2030 1248 2034 1252
rect 1974 1178 1978 1182
rect 2014 1168 2018 1172
rect 2054 1218 2058 1222
rect 2054 1148 2058 1152
rect 2078 1148 2082 1152
rect 2046 1118 2050 1122
rect 2038 1098 2042 1102
rect 2030 1088 2034 1092
rect 2030 1078 2034 1082
rect 1974 1068 1978 1072
rect 2198 1438 2202 1442
rect 2230 1438 2234 1442
rect 2214 1328 2218 1332
rect 2182 1288 2186 1292
rect 2174 1268 2178 1272
rect 2174 1258 2178 1262
rect 2158 1248 2162 1252
rect 2182 1248 2186 1252
rect 2102 1158 2106 1162
rect 2166 1158 2170 1162
rect 2102 1148 2106 1152
rect 2086 1138 2090 1142
rect 2070 1088 2074 1092
rect 2078 1068 2082 1072
rect 2014 978 2018 982
rect 1982 968 1986 972
rect 1966 958 1970 962
rect 1942 948 1946 952
rect 1950 948 1954 952
rect 1998 948 2002 952
rect 1918 918 1922 922
rect 1914 903 1918 907
rect 1921 903 1925 907
rect 1926 888 1930 892
rect 1974 878 1978 882
rect 2006 938 2010 942
rect 2030 958 2034 962
rect 2038 958 2042 962
rect 2078 1048 2082 1052
rect 2102 1058 2106 1062
rect 2142 1058 2146 1062
rect 2134 968 2138 972
rect 2046 948 2050 952
rect 2086 947 2090 951
rect 2022 938 2026 942
rect 2110 938 2114 942
rect 2174 938 2178 942
rect 2022 888 2026 892
rect 1990 868 1994 872
rect 1958 858 1962 862
rect 1878 818 1882 822
rect 1814 758 1818 762
rect 1830 758 1834 762
rect 1862 758 1866 762
rect 1934 848 1938 852
rect 1958 838 1962 842
rect 1934 828 1938 832
rect 1998 788 2002 792
rect 1918 768 1922 772
rect 1958 768 1962 772
rect 1822 748 1826 752
rect 1838 748 1842 752
rect 1870 748 1874 752
rect 1750 738 1754 742
rect 1758 728 1762 732
rect 1830 728 1834 732
rect 1774 718 1778 722
rect 1766 708 1770 712
rect 1686 698 1690 702
rect 1710 698 1714 702
rect 1718 698 1722 702
rect 1590 688 1594 692
rect 1606 688 1610 692
rect 1566 668 1570 672
rect 1574 668 1578 672
rect 1654 688 1658 692
rect 1686 688 1690 692
rect 1702 688 1706 692
rect 1638 668 1642 672
rect 1678 668 1682 672
rect 1494 658 1498 662
rect 1486 648 1490 652
rect 1638 648 1642 652
rect 1654 648 1658 652
rect 1630 628 1634 632
rect 1622 618 1626 622
rect 1470 588 1474 592
rect 1550 598 1554 602
rect 1606 598 1610 602
rect 1518 568 1522 572
rect 1446 528 1450 532
rect 1438 518 1442 522
rect 1454 518 1458 522
rect 1486 548 1490 552
rect 1478 538 1482 542
rect 1614 588 1618 592
rect 1614 578 1618 582
rect 1830 698 1834 702
rect 1886 708 1890 712
rect 1878 688 1882 692
rect 1854 678 1858 682
rect 1862 678 1866 682
rect 1726 668 1730 672
rect 1766 668 1770 672
rect 1710 648 1714 652
rect 1678 638 1682 642
rect 1662 588 1666 592
rect 1662 568 1666 572
rect 1742 568 1746 572
rect 1630 548 1634 552
rect 1646 548 1650 552
rect 1726 548 1730 552
rect 1914 703 1918 707
rect 1921 703 1925 707
rect 1902 658 1906 662
rect 1798 578 1802 582
rect 1574 538 1578 542
rect 1478 498 1482 502
rect 1470 478 1474 482
rect 1326 448 1330 452
rect 1254 438 1258 442
rect 1246 368 1250 372
rect 1302 368 1306 372
rect 1166 358 1170 362
rect 1182 358 1186 362
rect 1086 348 1090 352
rect 1110 348 1114 352
rect 1134 348 1138 352
rect 1150 348 1154 352
rect 1158 338 1162 342
rect 902 258 906 262
rect 846 248 850 252
rect 782 238 786 242
rect 830 238 834 242
rect 814 218 818 222
rect 798 208 802 212
rect 774 178 778 182
rect 822 178 826 182
rect 902 178 906 182
rect 830 168 834 172
rect 854 168 858 172
rect 830 148 834 152
rect 854 148 858 152
rect 774 138 778 142
rect 798 138 802 142
rect 814 138 818 142
rect 430 118 434 122
rect 478 108 482 112
rect 438 78 442 82
rect 390 68 394 72
rect 454 68 458 72
rect 486 98 490 102
rect 494 98 498 102
rect 686 128 690 132
rect 614 98 618 102
rect 526 88 530 92
rect 558 88 562 92
rect 590 88 594 92
rect 686 88 690 92
rect 694 78 698 82
rect 774 98 778 102
rect 790 88 794 92
rect 726 78 730 82
rect 646 68 650 72
rect 294 58 298 62
rect 310 58 314 62
rect 374 58 378 62
rect 414 58 418 62
rect 886 128 890 132
rect 806 98 810 102
rect 814 78 818 82
rect 782 68 786 72
rect 882 103 886 107
rect 889 103 893 107
rect 862 78 866 82
rect 998 218 1002 222
rect 974 208 978 212
rect 998 208 1002 212
rect 1022 188 1026 192
rect 926 158 930 162
rect 982 128 986 132
rect 942 118 946 122
rect 1046 268 1050 272
rect 1070 318 1074 322
rect 1110 318 1114 322
rect 1158 318 1162 322
rect 1062 288 1066 292
rect 1142 298 1146 302
rect 1142 288 1146 292
rect 1086 268 1090 272
rect 1102 248 1106 252
rect 1118 248 1122 252
rect 1094 198 1098 202
rect 1086 178 1090 182
rect 1038 168 1042 172
rect 1038 158 1042 162
rect 1054 138 1058 142
rect 1030 98 1034 102
rect 918 88 922 92
rect 942 88 946 92
rect 958 88 962 92
rect 1046 88 1050 92
rect 870 68 874 72
rect 934 58 938 62
rect 462 48 466 52
rect 478 48 482 52
rect 622 48 626 52
rect 782 38 786 42
rect 378 3 382 7
rect 385 3 389 7
rect 830 48 834 52
rect 1150 188 1154 192
rect 1110 168 1114 172
rect 1102 148 1106 152
rect 1134 148 1138 152
rect 1254 358 1258 362
rect 1286 348 1290 352
rect 1206 338 1210 342
rect 1214 288 1218 292
rect 1214 238 1218 242
rect 1182 218 1186 222
rect 1198 218 1202 222
rect 1174 208 1178 212
rect 1158 158 1162 162
rect 1166 158 1170 162
rect 1206 158 1210 162
rect 1214 158 1218 162
rect 1166 138 1170 142
rect 1190 138 1194 142
rect 1102 98 1106 102
rect 1206 88 1210 92
rect 1254 338 1258 342
rect 1254 268 1258 272
rect 1238 218 1242 222
rect 1270 298 1274 302
rect 1310 338 1314 342
rect 1374 458 1378 462
rect 1390 458 1394 462
rect 1358 438 1362 442
rect 1394 403 1398 407
rect 1401 403 1405 407
rect 1494 468 1498 472
rect 1446 448 1450 452
rect 1510 488 1514 492
rect 1590 488 1594 492
rect 1670 528 1674 532
rect 1630 498 1634 502
rect 1654 498 1658 502
rect 1662 498 1666 502
rect 1534 448 1538 452
rect 1638 448 1642 452
rect 1502 428 1506 432
rect 1518 428 1522 432
rect 1534 428 1538 432
rect 1486 418 1490 422
rect 1350 368 1354 372
rect 1414 368 1418 372
rect 1430 368 1434 372
rect 1398 358 1402 362
rect 1366 348 1370 352
rect 1398 348 1402 352
rect 1342 338 1346 342
rect 1334 328 1338 332
rect 1294 288 1298 292
rect 1278 278 1282 282
rect 1478 358 1482 362
rect 1574 418 1578 422
rect 1550 398 1554 402
rect 1526 388 1530 392
rect 1542 368 1546 372
rect 1606 378 1610 382
rect 1622 378 1626 382
rect 1598 358 1602 362
rect 1454 338 1458 342
rect 1526 338 1530 342
rect 1462 328 1466 332
rect 1430 308 1434 312
rect 1438 288 1442 292
rect 1350 278 1354 282
rect 1398 278 1402 282
rect 1430 278 1434 282
rect 1342 248 1346 252
rect 1310 228 1314 232
rect 1262 188 1266 192
rect 1278 178 1282 182
rect 1342 218 1346 222
rect 1406 228 1410 232
rect 1374 218 1378 222
rect 1350 178 1354 182
rect 1230 158 1234 162
rect 1262 158 1266 162
rect 1358 158 1362 162
rect 1286 138 1290 142
rect 1006 78 1010 82
rect 1062 78 1066 82
rect 1142 78 1146 82
rect 990 48 994 52
rect 1254 108 1258 112
rect 1286 108 1290 112
rect 1278 98 1282 102
rect 1238 78 1242 82
rect 1150 58 1154 62
rect 1294 58 1298 62
rect 1350 138 1354 142
rect 1366 138 1370 142
rect 1326 108 1330 112
rect 1326 98 1330 102
rect 1350 98 1354 102
rect 1318 88 1322 92
rect 1394 203 1398 207
rect 1401 203 1405 207
rect 1422 158 1426 162
rect 1382 148 1386 152
rect 1414 148 1418 152
rect 1454 258 1458 262
rect 1454 238 1458 242
rect 1590 328 1594 332
rect 1558 298 1562 302
rect 1574 298 1578 302
rect 1486 288 1490 292
rect 1526 268 1530 272
rect 1470 258 1474 262
rect 1478 238 1482 242
rect 1486 238 1490 242
rect 1478 228 1482 232
rect 1494 218 1498 222
rect 1486 188 1490 192
rect 1374 78 1378 82
rect 1310 58 1314 62
rect 1550 248 1554 252
rect 1534 218 1538 222
rect 1638 368 1642 372
rect 1646 368 1650 372
rect 1614 358 1618 362
rect 1694 518 1698 522
rect 1678 488 1682 492
rect 1822 548 1826 552
rect 1790 528 1794 532
rect 1862 638 1866 642
rect 1838 578 1842 582
rect 1846 558 1850 562
rect 1814 478 1818 482
rect 1806 468 1810 472
rect 1854 538 1858 542
rect 2158 928 2162 932
rect 2086 898 2090 902
rect 2134 868 2138 872
rect 2030 858 2034 862
rect 2078 848 2082 852
rect 2094 788 2098 792
rect 2038 778 2042 782
rect 2006 758 2010 762
rect 2022 758 2026 762
rect 1974 748 1978 752
rect 1982 738 1986 742
rect 1966 728 1970 732
rect 1934 638 1938 642
rect 1894 598 1898 602
rect 1886 578 1890 582
rect 1910 608 1914 612
rect 1934 598 1938 602
rect 2014 728 2018 732
rect 1998 648 2002 652
rect 2014 638 2018 642
rect 1998 628 2002 632
rect 2070 768 2074 772
rect 2118 758 2122 762
rect 2126 758 2130 762
rect 2054 748 2058 752
rect 2046 698 2050 702
rect 2038 658 2042 662
rect 1958 568 1962 572
rect 2030 568 2034 572
rect 1902 558 1906 562
rect 1910 548 1914 552
rect 1942 548 1946 552
rect 1886 538 1890 542
rect 1878 528 1882 532
rect 1914 503 1918 507
rect 1921 503 1925 507
rect 2006 548 2010 552
rect 2030 548 2034 552
rect 1950 498 1954 502
rect 1926 488 1930 492
rect 1942 488 1946 492
rect 1838 468 1842 472
rect 1662 458 1666 462
rect 1734 458 1738 462
rect 1790 458 1794 462
rect 1670 448 1674 452
rect 1686 398 1690 402
rect 1678 368 1682 372
rect 1734 368 1738 372
rect 1806 368 1810 372
rect 1742 358 1746 362
rect 1774 358 1778 362
rect 1662 348 1666 352
rect 1710 348 1714 352
rect 1782 348 1786 352
rect 1614 338 1618 342
rect 1710 338 1714 342
rect 1846 438 1850 442
rect 1838 378 1842 382
rect 1910 358 1914 362
rect 1630 328 1634 332
rect 1678 318 1682 322
rect 1630 308 1634 312
rect 1654 308 1658 312
rect 1606 298 1610 302
rect 1614 298 1618 302
rect 1622 278 1626 282
rect 1614 268 1618 272
rect 1718 328 1722 332
rect 1694 318 1698 322
rect 1686 308 1690 312
rect 1662 268 1666 272
rect 1606 248 1610 252
rect 1646 248 1650 252
rect 1590 238 1594 242
rect 1678 238 1682 242
rect 1574 138 1578 142
rect 1470 98 1474 102
rect 1430 88 1434 92
rect 1438 78 1442 82
rect 1534 78 1538 82
rect 1550 58 1554 62
rect 1582 118 1586 122
rect 1606 218 1610 222
rect 1710 218 1714 222
rect 1614 168 1618 172
rect 1686 168 1690 172
rect 1622 148 1626 152
rect 1566 58 1570 62
rect 1614 58 1618 62
rect 1702 158 1706 162
rect 1782 328 1786 332
rect 1734 318 1738 322
rect 1774 318 1778 322
rect 1726 308 1730 312
rect 1758 308 1762 312
rect 2022 528 2026 532
rect 2006 518 2010 522
rect 2014 508 2018 512
rect 2046 648 2050 652
rect 2038 488 2042 492
rect 2110 728 2114 732
rect 2102 718 2106 722
rect 2174 798 2178 802
rect 2158 768 2162 772
rect 2174 748 2178 752
rect 2238 1258 2242 1262
rect 2230 1138 2234 1142
rect 2238 958 2242 962
rect 2190 888 2194 892
rect 2238 888 2242 892
rect 2222 878 2226 882
rect 2270 1498 2274 1502
rect 2294 1538 2298 1542
rect 2278 1448 2282 1452
rect 2286 1338 2290 1342
rect 2262 1318 2266 1322
rect 2302 1348 2306 1352
rect 2302 1248 2306 1252
rect 2294 1238 2298 1242
rect 2286 1168 2290 1172
rect 2278 1118 2282 1122
rect 2286 1098 2290 1102
rect 2294 1078 2298 1082
rect 2270 968 2274 972
rect 2262 948 2266 952
rect 2278 898 2282 902
rect 2302 968 2306 972
rect 2238 858 2242 862
rect 2254 858 2258 862
rect 2270 848 2274 852
rect 2206 838 2210 842
rect 2198 798 2202 802
rect 2270 838 2274 842
rect 2238 778 2242 782
rect 2206 728 2210 732
rect 2214 728 2218 732
rect 2182 718 2186 722
rect 2270 698 2274 702
rect 2286 688 2290 692
rect 2078 658 2082 662
rect 2094 658 2098 662
rect 2094 648 2098 652
rect 2102 628 2106 632
rect 2062 598 2066 602
rect 2062 558 2066 562
rect 2094 548 2098 552
rect 2054 508 2058 512
rect 2166 658 2170 662
rect 2246 648 2250 652
rect 2126 638 2130 642
rect 2110 618 2114 622
rect 2142 618 2146 622
rect 2134 558 2138 562
rect 2150 588 2154 592
rect 2142 528 2146 532
rect 2142 518 2146 522
rect 2102 498 2106 502
rect 2110 498 2114 502
rect 2054 478 2058 482
rect 2070 478 2074 482
rect 2086 478 2090 482
rect 1966 468 1970 472
rect 2030 468 2034 472
rect 2038 468 2042 472
rect 1990 368 1994 372
rect 2014 368 2018 372
rect 2030 368 2034 372
rect 1982 358 1986 362
rect 2006 358 2010 362
rect 1830 318 1834 322
rect 1814 308 1818 312
rect 1862 318 1866 322
rect 1914 303 1918 307
rect 1921 303 1925 307
rect 1854 288 1858 292
rect 1878 278 1882 282
rect 1790 238 1794 242
rect 1862 188 1866 192
rect 1774 168 1778 172
rect 1726 158 1730 162
rect 1710 118 1714 122
rect 1742 118 1746 122
rect 1646 98 1650 102
rect 1766 98 1770 102
rect 1870 158 1874 162
rect 1830 118 1834 122
rect 1854 118 1858 122
rect 1822 108 1826 112
rect 1838 108 1842 112
rect 1814 78 1818 82
rect 1830 98 1834 102
rect 1838 88 1842 92
rect 1846 78 1850 82
rect 1854 78 1858 82
rect 1910 248 1914 252
rect 1966 328 1970 332
rect 1966 298 1970 302
rect 1966 268 1970 272
rect 1998 348 2002 352
rect 1998 318 2002 322
rect 2006 268 2010 272
rect 1974 258 1978 262
rect 1982 258 1986 262
rect 2022 328 2026 332
rect 2022 308 2026 312
rect 2014 198 2018 202
rect 1894 158 1898 162
rect 1886 128 1890 132
rect 1894 118 1898 122
rect 1934 118 1938 122
rect 1914 103 1918 107
rect 1921 103 1925 107
rect 1694 58 1698 62
rect 1742 58 1746 62
rect 1790 58 1794 62
rect 1798 58 1802 62
rect 1390 48 1394 52
rect 1406 48 1410 52
rect 1502 48 1506 52
rect 1558 48 1562 52
rect 1582 48 1586 52
rect 1614 48 1618 52
rect 1078 8 1082 12
rect 1094 8 1098 12
rect 1614 8 1618 12
rect 1394 3 1398 7
rect 1401 3 1405 7
rect 2022 98 2026 102
rect 1878 58 1882 62
rect 1902 58 1906 62
rect 1934 58 1938 62
rect 1974 58 1978 62
rect 1982 58 1986 62
rect 1894 38 1898 42
rect 2118 468 2122 472
rect 2086 458 2090 462
rect 2102 458 2106 462
rect 2134 458 2138 462
rect 2070 438 2074 442
rect 2126 448 2130 452
rect 2174 548 2178 552
rect 2214 548 2218 552
rect 2302 748 2306 752
rect 2294 628 2298 632
rect 2270 558 2274 562
rect 2286 538 2290 542
rect 2166 518 2170 522
rect 2198 498 2202 502
rect 2174 488 2178 492
rect 2166 468 2170 472
rect 2158 408 2162 412
rect 2158 358 2162 362
rect 2198 458 2202 462
rect 2174 358 2178 362
rect 2150 348 2154 352
rect 2166 348 2170 352
rect 2182 348 2186 352
rect 2046 308 2050 312
rect 2038 298 2042 302
rect 2110 298 2114 302
rect 2094 278 2098 282
rect 2062 268 2066 272
rect 2038 258 2042 262
rect 2070 258 2074 262
rect 2038 238 2042 242
rect 2198 438 2202 442
rect 2198 328 2202 332
rect 2150 268 2154 272
rect 2158 268 2162 272
rect 2118 148 2122 152
rect 2150 148 2154 152
rect 2078 138 2082 142
rect 2102 138 2106 142
rect 2094 118 2098 122
rect 2134 118 2138 122
rect 2062 108 2066 112
rect 2094 108 2098 112
rect 2078 88 2082 92
rect 2190 258 2194 262
rect 2174 178 2178 182
rect 2166 98 2170 102
rect 2238 458 2242 462
rect 2214 308 2218 312
rect 2262 338 2266 342
rect 2254 328 2258 332
rect 2302 328 2306 332
rect 2246 268 2250 272
rect 2206 258 2210 262
rect 2270 318 2274 322
rect 2294 268 2298 272
rect 2286 218 2290 222
rect 2254 158 2258 162
rect 2286 158 2290 162
rect 2214 98 2218 102
rect 2142 68 2146 72
rect 2270 68 2274 72
rect 2046 58 2050 62
rect 2174 58 2178 62
rect 2230 58 2234 62
rect 2254 58 2258 62
rect 2022 48 2026 52
rect 2030 48 2034 52
rect 2190 38 2194 42
<< metal3 >>
rect 880 2103 882 2107
rect 886 2103 889 2107
rect 894 2103 896 2107
rect 1912 2103 1914 2107
rect 1918 2103 1921 2107
rect 1926 2103 1928 2107
rect 250 2088 606 2091
rect 610 2088 838 2091
rect 842 2088 1169 2091
rect 1522 2088 1566 2091
rect 1166 2082 1169 2088
rect 826 2078 926 2081
rect 1170 2078 1206 2081
rect 1370 2078 1382 2081
rect 1754 2078 1846 2081
rect 1874 2078 1886 2081
rect 318 2071 321 2078
rect 462 2071 465 2078
rect 142 2068 465 2071
rect 490 2068 574 2071
rect 978 2068 1025 2071
rect 1114 2068 1177 2071
rect 142 2062 145 2068
rect 158 2062 161 2068
rect 282 2058 289 2061
rect 306 2058 310 2061
rect 446 2058 638 2061
rect 690 2058 750 2061
rect 878 2058 886 2061
rect 890 2059 950 2061
rect 1022 2062 1025 2068
rect 1174 2062 1177 2068
rect 1298 2068 1433 2071
rect 890 2058 953 2059
rect 1058 2058 1134 2061
rect 1262 2061 1265 2068
rect 1210 2058 1265 2061
rect 1430 2062 1433 2068
rect 1686 2068 1814 2071
rect 2066 2068 2150 2071
rect 2218 2068 2222 2071
rect 2234 2068 2238 2071
rect 1534 2061 1537 2068
rect 1466 2058 1537 2061
rect 1686 2062 1689 2068
rect 1814 2061 1817 2068
rect 1738 2058 1785 2061
rect 1814 2058 1910 2061
rect 1914 2058 1966 2061
rect 1994 2058 2078 2061
rect 2082 2058 2110 2061
rect 2138 2058 2241 2061
rect 294 2052 297 2058
rect 334 2052 337 2058
rect 446 2052 449 2058
rect 1782 2052 1785 2058
rect 2238 2052 2241 2058
rect 2246 2052 2249 2058
rect -26 2051 -22 2052
rect -26 2048 6 2051
rect 10 2048 78 2051
rect 554 2048 574 2051
rect 906 2048 910 2051
rect 1106 2048 1145 2051
rect 1162 2048 1214 2051
rect 1530 2048 1550 2051
rect 1554 2048 1710 2051
rect 1714 2048 1726 2051
rect 2018 2048 2022 2051
rect 2042 2048 2070 2051
rect 2074 2048 2174 2051
rect 2266 2048 2286 2051
rect 2334 2051 2338 2052
rect 2306 2048 2338 2051
rect 234 2038 254 2041
rect 258 2038 334 2041
rect 430 2041 433 2048
rect 338 2038 433 2041
rect 582 2041 585 2048
rect 1142 2042 1145 2048
rect 554 2038 585 2041
rect 762 2038 894 2041
rect 898 2038 1110 2041
rect 1230 2041 1233 2048
rect 1202 2038 1217 2041
rect 1230 2038 1318 2041
rect 1322 2038 1334 2041
rect 1674 2038 1766 2041
rect 1214 2032 1217 2038
rect 274 2028 390 2031
rect 394 2028 654 2031
rect 866 2028 998 2031
rect 1282 2028 1390 2031
rect 202 2018 241 2021
rect 482 2018 670 2021
rect 674 2018 774 2021
rect 778 2018 838 2021
rect 1402 2018 1774 2021
rect 2106 2018 2110 2021
rect 2258 2018 2262 2021
rect 238 2012 241 2018
rect 738 2008 774 2011
rect 778 2008 958 2011
rect 1090 2008 1246 2011
rect 1250 2008 1286 2011
rect 1570 2008 1822 2011
rect 376 2003 378 2007
rect 382 2003 385 2007
rect 390 2003 392 2007
rect 1392 2003 1394 2007
rect 1398 2003 1401 2007
rect 1406 2003 1408 2007
rect 1146 1998 1350 2001
rect 1570 1998 1574 2001
rect 1578 1998 1862 2001
rect 1866 1998 2014 2001
rect 826 1988 1702 1991
rect 1706 1988 1758 1991
rect 1762 1988 2030 1991
rect 18 1978 134 1981
rect 1114 1978 1118 1981
rect 1122 1978 1342 1981
rect 1610 1978 1806 1981
rect 2018 1978 2078 1981
rect 106 1968 158 1971
rect 170 1968 222 1971
rect 254 1968 262 1971
rect 266 1968 374 1971
rect 378 1968 566 1971
rect 642 1968 646 1971
rect 878 1971 881 1978
rect 866 1968 881 1971
rect 1042 1968 1062 1971
rect 1218 1968 1270 1971
rect 1274 1968 1281 1971
rect 1358 1968 1374 1971
rect 1378 1968 1406 1971
rect 1594 1968 1606 1971
rect 130 1958 302 1961
rect 498 1958 502 1961
rect 602 1958 662 1961
rect 710 1958 790 1961
rect 794 1958 846 1961
rect 850 1958 870 1961
rect 874 1958 902 1961
rect 1026 1958 1225 1961
rect 1302 1961 1305 1968
rect 1266 1958 1305 1961
rect 1358 1962 1361 1968
rect 1382 1958 1390 1961
rect 1394 1958 1470 1961
rect 1522 1958 1606 1961
rect 1618 1958 1638 1961
rect 1642 1958 1646 1961
rect 1850 1958 1926 1961
rect 1970 1958 2118 1961
rect 70 1951 73 1958
rect 710 1952 713 1958
rect 1222 1952 1225 1958
rect 70 1948 110 1951
rect 162 1948 230 1951
rect 290 1948 510 1951
rect 514 1948 518 1951
rect 522 1948 558 1951
rect 578 1948 582 1951
rect 626 1948 710 1951
rect 762 1948 766 1951
rect 770 1948 854 1951
rect 858 1948 902 1951
rect 906 1948 1206 1951
rect 1226 1948 1270 1951
rect 1346 1948 1390 1951
rect 1394 1948 1478 1951
rect 1482 1948 1518 1951
rect 1634 1948 1702 1951
rect 1794 1948 1862 1951
rect 1866 1948 1894 1951
rect 2050 1948 2062 1951
rect 2246 1951 2249 1958
rect 2170 1948 2249 1951
rect 590 1942 593 1948
rect 170 1938 246 1941
rect 266 1938 318 1941
rect 458 1938 510 1941
rect 530 1938 574 1941
rect 602 1938 638 1941
rect 714 1938 718 1941
rect 726 1941 729 1948
rect 726 1938 806 1941
rect 858 1938 942 1941
rect 1038 1938 1102 1941
rect 1162 1938 1166 1941
rect 1186 1938 1414 1941
rect 1590 1941 1593 1948
rect 1590 1938 1710 1941
rect 1890 1938 1990 1941
rect 2050 1938 2142 1941
rect 1022 1932 1025 1938
rect 1038 1932 1041 1938
rect 1854 1932 1857 1938
rect 66 1928 414 1931
rect 506 1928 582 1931
rect 1050 1928 1158 1931
rect 1274 1928 1390 1931
rect 1562 1928 1766 1931
rect 1770 1928 1790 1931
rect 122 1918 182 1921
rect 186 1918 190 1921
rect 274 1918 294 1921
rect 466 1918 622 1921
rect 882 1918 1054 1921
rect 1074 1918 1166 1921
rect 1818 1918 1862 1921
rect 2194 1918 2209 1921
rect 2206 1912 2209 1918
rect 194 1908 262 1911
rect 266 1908 286 1911
rect 290 1908 366 1911
rect 370 1908 742 1911
rect 986 1908 998 1911
rect 1146 1908 1158 1911
rect 1162 1908 1318 1911
rect 1322 1908 1414 1911
rect 1418 1908 1438 1911
rect 880 1903 882 1907
rect 886 1903 889 1907
rect 894 1903 896 1907
rect 1912 1903 1914 1907
rect 1918 1903 1921 1907
rect 1926 1903 1928 1907
rect 234 1898 326 1901
rect 330 1898 806 1901
rect 914 1898 1006 1901
rect 1010 1898 1046 1901
rect 1066 1898 1182 1901
rect 1218 1898 1470 1901
rect 1834 1898 1862 1901
rect 2074 1898 2214 1901
rect 2218 1898 2230 1901
rect 810 1888 1326 1891
rect 1578 1888 1614 1891
rect 2078 1888 2174 1891
rect 202 1878 278 1881
rect 666 1878 702 1881
rect 1042 1878 1094 1881
rect 1098 1878 1158 1881
rect 1326 1881 1329 1888
rect 1326 1878 1406 1881
rect 1526 1881 1529 1888
rect 2078 1882 2081 1888
rect 1498 1878 1529 1881
rect 1738 1878 1750 1881
rect 1786 1878 1790 1881
rect 1842 1878 1878 1881
rect 2042 1878 2078 1881
rect 138 1868 382 1871
rect 586 1868 614 1871
rect 618 1868 694 1871
rect 698 1868 710 1871
rect 746 1868 1270 1871
rect 1494 1868 1526 1871
rect 1594 1868 1606 1871
rect 1610 1868 1638 1871
rect 1766 1871 1769 1878
rect 1682 1868 1769 1871
rect 1810 1868 1830 1871
rect 1850 1868 1942 1871
rect 1970 1868 1998 1871
rect 2018 1868 2046 1871
rect 2226 1868 2270 1871
rect 1494 1862 1497 1868
rect 58 1858 102 1861
rect 114 1858 118 1861
rect 242 1858 398 1861
rect 470 1858 478 1861
rect 482 1858 542 1861
rect 562 1858 630 1861
rect 642 1858 686 1861
rect 754 1858 774 1861
rect 778 1858 870 1861
rect 882 1858 918 1861
rect 946 1858 950 1861
rect 994 1858 1014 1861
rect 1194 1858 1262 1861
rect 1402 1858 1470 1861
rect 1514 1858 1598 1861
rect 1618 1858 1630 1861
rect 1634 1858 1782 1861
rect 1786 1858 1798 1861
rect 1858 1858 2022 1861
rect 2142 1861 2145 1868
rect 2142 1858 2190 1861
rect 114 1848 126 1851
rect 498 1848 590 1851
rect 594 1848 606 1851
rect 626 1848 646 1851
rect 770 1848 1054 1851
rect 1182 1851 1185 1858
rect 1082 1848 1222 1851
rect 1346 1848 1454 1851
rect 1474 1848 1486 1851
rect 1874 1848 1934 1851
rect 1938 1848 1982 1851
rect 2258 1848 2270 1851
rect 134 1841 137 1848
rect 106 1838 137 1841
rect 294 1841 297 1848
rect 266 1838 670 1841
rect 762 1838 822 1841
rect 842 1838 878 1841
rect 886 1838 918 1841
rect 954 1838 958 1841
rect 1466 1838 1582 1841
rect 1866 1838 2062 1841
rect 2066 1838 2190 1841
rect 2194 1838 2214 1841
rect 886 1832 889 1838
rect 362 1828 526 1831
rect 562 1828 566 1831
rect 570 1828 598 1831
rect 602 1828 678 1831
rect 1018 1828 1518 1831
rect 1978 1828 2198 1831
rect 418 1818 430 1821
rect 434 1818 638 1821
rect 642 1818 1086 1821
rect 1090 1818 1534 1821
rect 1554 1818 1822 1821
rect 1826 1818 1886 1821
rect 2186 1818 2302 1821
rect 522 1808 870 1811
rect 1554 1808 1590 1811
rect 1762 1808 1990 1811
rect 2210 1808 2222 1811
rect 376 1803 378 1807
rect 382 1803 385 1807
rect 390 1803 392 1807
rect 1392 1803 1394 1807
rect 1398 1803 1401 1807
rect 1406 1803 1408 1807
rect 338 1798 342 1801
rect 514 1798 550 1801
rect 618 1798 694 1801
rect 826 1798 934 1801
rect 986 1798 1166 1801
rect 1554 1798 1654 1801
rect 346 1788 350 1791
rect 354 1788 422 1791
rect 690 1788 982 1791
rect 986 1788 1118 1791
rect 1166 1791 1169 1798
rect 1166 1788 1446 1791
rect 1610 1788 1614 1791
rect 1834 1788 1998 1791
rect 138 1778 398 1781
rect 666 1778 670 1781
rect 698 1778 854 1781
rect 858 1778 998 1781
rect 1002 1778 1070 1781
rect 1090 1778 1110 1781
rect 1370 1778 1430 1781
rect 1946 1778 2150 1781
rect 2154 1778 2254 1781
rect 122 1768 358 1771
rect 578 1768 590 1771
rect 826 1768 886 1771
rect 1158 1768 1246 1771
rect 1634 1768 1718 1771
rect 1722 1768 1766 1771
rect 1858 1768 1950 1771
rect 1986 1768 2046 1771
rect 2098 1768 2102 1771
rect 1158 1762 1161 1768
rect 338 1758 342 1761
rect 530 1758 574 1761
rect 578 1758 630 1761
rect 866 1758 926 1761
rect 930 1758 958 1761
rect 1138 1758 1150 1761
rect 1426 1758 1478 1761
rect 1802 1758 1894 1761
rect 2034 1758 2086 1761
rect 2178 1758 2262 1761
rect 2266 1758 2294 1761
rect 66 1748 113 1751
rect 110 1742 113 1748
rect 298 1748 350 1751
rect 490 1748 558 1751
rect 662 1751 665 1758
rect 702 1751 705 1758
rect 662 1748 705 1751
rect 878 1748 1062 1751
rect 1130 1748 1193 1751
rect 1234 1748 1542 1751
rect 1546 1748 1558 1751
rect 1594 1748 1614 1751
rect 1834 1748 1862 1751
rect 1882 1748 1897 1751
rect 1990 1751 1993 1758
rect 1954 1748 1993 1751
rect 2018 1748 2070 1751
rect 2102 1751 2105 1758
rect 2074 1748 2105 1751
rect 2150 1752 2153 1758
rect 2218 1748 2278 1751
rect 114 1738 222 1741
rect 254 1741 257 1748
rect 598 1742 601 1748
rect 878 1742 881 1748
rect 226 1738 257 1741
rect 362 1738 518 1741
rect 522 1738 542 1741
rect 666 1738 670 1741
rect 690 1738 710 1741
rect 898 1738 934 1741
rect 938 1738 982 1741
rect 1102 1741 1105 1748
rect 1010 1738 1105 1741
rect 1190 1742 1193 1748
rect 1298 1738 1302 1741
rect 1318 1738 1382 1741
rect 1394 1738 1414 1741
rect 1418 1738 1534 1741
rect 1582 1741 1585 1748
rect 1894 1742 1897 1748
rect 1538 1738 1590 1741
rect 1610 1738 1662 1741
rect 1810 1738 1841 1741
rect 1898 1738 1942 1741
rect 2010 1738 2118 1741
rect 2122 1738 2206 1741
rect 1318 1732 1321 1738
rect 1838 1732 1841 1738
rect 202 1728 246 1731
rect 250 1728 270 1731
rect 282 1728 734 1731
rect 738 1728 862 1731
rect 1018 1728 1030 1731
rect 1042 1728 1142 1731
rect 1178 1728 1190 1731
rect 1898 1728 2086 1731
rect 2090 1728 2110 1731
rect 2114 1728 2190 1731
rect 522 1718 534 1721
rect 538 1718 766 1721
rect 874 1718 942 1721
rect 946 1718 1030 1721
rect 1050 1718 1590 1721
rect 1938 1718 1966 1721
rect 1978 1718 2006 1721
rect 10 1708 174 1711
rect 178 1708 462 1711
rect 570 1708 582 1711
rect 1026 1708 1134 1711
rect 1138 1708 1158 1711
rect 1210 1708 1678 1711
rect 1690 1708 1846 1711
rect 880 1703 882 1707
rect 886 1703 889 1707
rect 894 1703 896 1707
rect 1912 1703 1914 1707
rect 1918 1703 1921 1707
rect 1926 1703 1928 1707
rect 770 1698 830 1701
rect 938 1698 1046 1701
rect 1114 1698 1222 1701
rect 1290 1698 1350 1701
rect 1506 1698 1574 1701
rect 1578 1698 1742 1701
rect 1882 1698 1886 1701
rect 2138 1698 2166 1701
rect 410 1688 622 1691
rect 738 1688 854 1691
rect 1066 1688 1158 1691
rect 1162 1688 1302 1691
rect 1530 1688 2014 1691
rect 326 1681 329 1688
rect 242 1678 329 1681
rect 426 1678 534 1681
rect 650 1678 686 1681
rect 1138 1678 1310 1681
rect 1466 1678 1590 1681
rect 1594 1678 1662 1681
rect 1762 1678 1822 1681
rect 82 1668 102 1671
rect 106 1668 110 1671
rect 178 1668 190 1671
rect 282 1668 430 1671
rect 522 1668 526 1671
rect 586 1668 590 1671
rect 954 1668 1006 1671
rect 1010 1668 1038 1671
rect 1242 1668 1278 1671
rect 1362 1668 1382 1671
rect 1450 1668 1542 1671
rect 1562 1668 1566 1671
rect 1618 1668 1702 1671
rect 1726 1671 1729 1678
rect 1726 1668 1798 1671
rect 1802 1668 1814 1671
rect 1978 1668 2030 1671
rect 2078 1671 2081 1678
rect 2158 1671 2161 1678
rect 2078 1668 2161 1671
rect 2202 1668 2230 1671
rect 186 1658 278 1661
rect 354 1658 358 1661
rect 430 1661 433 1668
rect 430 1658 462 1661
rect 662 1661 665 1668
rect 522 1658 670 1661
rect 690 1658 734 1661
rect 750 1661 753 1668
rect 750 1658 806 1661
rect 914 1658 926 1661
rect 986 1658 998 1661
rect 1002 1658 1046 1661
rect 1058 1658 1142 1661
rect 1146 1658 1150 1661
rect 1294 1661 1297 1668
rect 1218 1658 1398 1661
rect 1530 1658 1550 1661
rect 1578 1658 1670 1661
rect 1750 1658 1777 1661
rect 1878 1661 1881 1668
rect 1850 1658 1881 1661
rect 2178 1658 2198 1661
rect 114 1648 126 1651
rect 130 1648 158 1651
rect 330 1648 366 1651
rect 482 1648 542 1651
rect 570 1648 606 1651
rect 610 1648 702 1651
rect 706 1648 718 1651
rect 974 1651 977 1658
rect 1246 1652 1249 1658
rect 1750 1652 1753 1658
rect 1774 1652 1777 1658
rect 974 1648 1006 1651
rect 1022 1648 1166 1651
rect 1218 1648 1238 1651
rect 1258 1648 1262 1651
rect 1318 1648 1358 1651
rect 1370 1648 1374 1651
rect 1554 1648 1574 1651
rect 1690 1648 1694 1651
rect 1698 1648 1718 1651
rect 1786 1648 1790 1651
rect 1842 1648 1862 1651
rect 1990 1651 1993 1658
rect 1874 1648 1993 1651
rect 2002 1648 2014 1651
rect 2130 1648 2182 1651
rect 2242 1648 2278 1651
rect 1022 1642 1025 1648
rect 1318 1642 1321 1648
rect 538 1638 590 1641
rect 594 1638 758 1641
rect 834 1638 918 1641
rect 922 1638 982 1641
rect 994 1638 1022 1641
rect 1562 1638 1734 1641
rect 1778 1638 1806 1641
rect 1842 1638 1950 1641
rect 1994 1638 2006 1641
rect 642 1628 1062 1631
rect 1298 1628 1742 1631
rect 58 1618 86 1621
rect 234 1618 750 1621
rect 978 1618 990 1621
rect 1002 1618 1022 1621
rect 1026 1618 1094 1621
rect 1242 1618 1326 1621
rect 1370 1618 1438 1621
rect 1538 1618 1542 1621
rect 1546 1618 1862 1621
rect 1866 1618 2022 1621
rect 426 1608 950 1611
rect 954 1608 1270 1611
rect 376 1603 378 1607
rect 382 1603 385 1607
rect 390 1603 392 1607
rect 1392 1603 1394 1607
rect 1398 1603 1401 1607
rect 1406 1603 1408 1607
rect 738 1598 1014 1601
rect 1034 1598 1238 1601
rect 1682 1598 1742 1601
rect 538 1588 614 1591
rect 642 1588 1006 1591
rect 1146 1588 1830 1591
rect 186 1578 254 1581
rect 258 1578 326 1581
rect 618 1578 782 1581
rect 986 1578 990 1581
rect 994 1578 1238 1581
rect 1386 1578 1422 1581
rect 1810 1578 1838 1581
rect 2074 1578 2166 1581
rect 18 1568 62 1571
rect 66 1568 174 1571
rect 258 1568 446 1571
rect 466 1568 550 1571
rect 642 1568 686 1571
rect 722 1568 1038 1571
rect 1442 1568 1510 1571
rect 1594 1568 1702 1571
rect 1786 1568 1846 1571
rect 2026 1568 2126 1571
rect 2130 1568 2166 1571
rect 118 1558 174 1561
rect 306 1558 558 1561
rect 586 1558 654 1561
rect 674 1558 678 1561
rect 794 1558 854 1561
rect 862 1558 894 1561
rect 962 1558 1086 1561
rect 1098 1558 1206 1561
rect 1218 1558 1318 1561
rect 1362 1558 1422 1561
rect 1458 1558 1542 1561
rect 1578 1558 1606 1561
rect 1718 1561 1721 1568
rect 1674 1558 1721 1561
rect 1802 1558 1806 1561
rect 2106 1558 2214 1561
rect 2262 1561 2265 1568
rect 2226 1558 2265 1561
rect 118 1552 121 1558
rect 862 1552 865 1558
rect 42 1548 102 1551
rect 418 1548 518 1551
rect 658 1548 670 1551
rect 842 1548 846 1551
rect 938 1548 1006 1551
rect 1234 1548 1254 1551
rect 1282 1548 1286 1551
rect 1306 1548 1454 1551
rect 1474 1548 1478 1551
rect 1566 1551 1569 1558
rect 1966 1552 1969 1558
rect 1490 1548 1569 1551
rect 1602 1548 1710 1551
rect 1818 1548 1838 1551
rect 2098 1548 2110 1551
rect 2114 1548 2134 1551
rect 2210 1548 2214 1551
rect 102 1542 105 1548
rect 42 1538 78 1541
rect 118 1538 150 1541
rect 482 1538 566 1541
rect 570 1538 710 1541
rect 770 1538 846 1541
rect 850 1538 982 1541
rect 1026 1538 1110 1541
rect 1166 1541 1169 1548
rect 1990 1542 1993 1548
rect 2142 1542 2145 1548
rect 1122 1538 1169 1541
rect 1194 1538 1334 1541
rect 1346 1538 1550 1541
rect 1730 1538 1790 1541
rect 1810 1538 1814 1541
rect 1842 1538 1902 1541
rect 2058 1538 2070 1541
rect 2074 1538 2078 1541
rect 2158 1541 2161 1548
rect 2158 1538 2174 1541
rect 2178 1538 2206 1541
rect 2246 1541 2249 1548
rect 2246 1538 2294 1541
rect 118 1532 121 1538
rect 438 1532 441 1538
rect 1550 1532 1553 1538
rect 10 1528 46 1531
rect 362 1528 422 1531
rect 466 1528 750 1531
rect 802 1528 894 1531
rect 946 1528 998 1531
rect 1010 1528 1046 1531
rect 1058 1528 1302 1531
rect 1394 1528 1398 1531
rect 1430 1528 1462 1531
rect 1490 1528 1534 1531
rect 1754 1528 1758 1531
rect 1770 1528 1806 1531
rect 1962 1528 2006 1531
rect 2034 1528 2262 1531
rect 1430 1522 1433 1528
rect 98 1518 118 1521
rect 202 1518 206 1521
rect 322 1518 462 1521
rect 522 1518 574 1521
rect 578 1518 846 1521
rect 850 1518 870 1521
rect 914 1518 1142 1521
rect 1162 1518 1230 1521
rect 1258 1518 1390 1521
rect 1450 1518 1518 1521
rect 1642 1518 1758 1521
rect 1802 1518 2150 1521
rect 2202 1518 2254 1521
rect 410 1508 454 1511
rect 738 1508 742 1511
rect 914 1508 1062 1511
rect 1066 1508 1230 1511
rect 1402 1508 1454 1511
rect 1458 1508 1550 1511
rect 1578 1508 1734 1511
rect 880 1503 882 1507
rect 886 1503 889 1507
rect 894 1503 896 1507
rect 1912 1503 1914 1507
rect 1918 1503 1921 1507
rect 1926 1503 1928 1507
rect 1982 1502 1985 1508
rect 58 1498 238 1501
rect 370 1498 542 1501
rect 706 1498 870 1501
rect 962 1498 966 1501
rect 970 1498 1494 1501
rect 1650 1498 1790 1501
rect 2170 1498 2270 1501
rect 106 1488 150 1491
rect 230 1488 390 1491
rect 450 1488 646 1491
rect 650 1488 817 1491
rect 1050 1488 1134 1491
rect 1146 1488 1158 1491
rect 1162 1488 1470 1491
rect 1482 1488 1534 1491
rect 1546 1488 1638 1491
rect 1730 1488 1878 1491
rect 1882 1488 1894 1491
rect 1946 1488 1950 1491
rect 1954 1488 1990 1491
rect 2054 1491 2057 1498
rect 2010 1488 2057 1491
rect 230 1482 233 1488
rect 90 1478 102 1481
rect 370 1478 478 1481
rect 482 1478 702 1481
rect 778 1478 806 1481
rect 814 1481 817 1488
rect 2070 1482 2073 1488
rect 814 1478 1182 1481
rect 1282 1478 1286 1481
rect 1306 1478 1318 1481
rect 1338 1478 1366 1481
rect 1498 1478 1782 1481
rect 1898 1478 2046 1481
rect 206 1471 209 1478
rect 114 1468 209 1471
rect 306 1468 310 1471
rect 346 1468 358 1471
rect 458 1468 478 1471
rect 538 1468 694 1471
rect 706 1468 782 1471
rect 802 1468 966 1471
rect 970 1468 1030 1471
rect 1058 1468 1174 1471
rect 1194 1468 1262 1471
rect 1266 1468 1350 1471
rect 1354 1468 1398 1471
rect 1478 1471 1481 1478
rect 1478 1468 1513 1471
rect 1530 1468 1590 1471
rect 1642 1468 1966 1471
rect 38 1461 41 1468
rect 1462 1462 1465 1468
rect 38 1458 126 1461
rect 186 1458 201 1461
rect 210 1458 214 1461
rect 258 1458 286 1461
rect 482 1458 534 1461
rect 602 1458 670 1461
rect 698 1458 790 1461
rect 874 1458 1014 1461
rect 1026 1458 1038 1461
rect 1094 1458 1126 1461
rect 1194 1458 1214 1461
rect 1242 1458 1246 1461
rect 1298 1458 1302 1461
rect 1306 1458 1374 1461
rect 1434 1458 1457 1461
rect 1490 1458 1494 1461
rect 1510 1461 1513 1468
rect 1506 1458 1513 1461
rect 1566 1458 1609 1461
rect 1706 1458 1766 1461
rect 1990 1461 1993 1468
rect 1946 1458 1993 1461
rect 2022 1461 2025 1468
rect 2022 1458 2070 1461
rect 2114 1458 2150 1461
rect 2154 1458 2174 1461
rect 2230 1461 2233 1468
rect 2194 1458 2233 1461
rect 198 1451 201 1458
rect 854 1452 857 1458
rect 106 1448 185 1451
rect 198 1448 222 1451
rect 250 1448 262 1451
rect 266 1448 302 1451
rect 434 1448 446 1451
rect 458 1448 462 1451
rect 578 1448 750 1451
rect 754 1448 838 1451
rect 914 1448 934 1451
rect 938 1448 998 1451
rect 1022 1451 1025 1458
rect 1002 1448 1025 1451
rect 1094 1452 1097 1458
rect 1190 1452 1193 1458
rect 1262 1451 1265 1458
rect 1454 1452 1457 1458
rect 1566 1452 1569 1458
rect 1606 1452 1609 1458
rect 1234 1448 1265 1451
rect 1282 1448 1302 1451
rect 1322 1448 1350 1451
rect 1498 1448 1502 1451
rect 1642 1448 1750 1451
rect 1754 1448 1766 1451
rect 1906 1448 1942 1451
rect 1946 1448 2278 1451
rect 182 1442 185 1448
rect 1358 1442 1361 1448
rect 114 1438 134 1441
rect 290 1438 398 1441
rect 650 1438 678 1441
rect 682 1438 702 1441
rect 714 1438 742 1441
rect 746 1438 790 1441
rect 838 1438 1022 1441
rect 1034 1438 1094 1441
rect 1170 1438 1214 1441
rect 1378 1438 1478 1441
rect 1586 1438 1790 1441
rect 2202 1438 2206 1441
rect 2234 1438 2246 1441
rect 174 1432 177 1438
rect 278 1432 281 1438
rect 838 1432 841 1438
rect 442 1428 654 1431
rect 658 1428 750 1431
rect 930 1428 990 1431
rect 1002 1428 1030 1431
rect 1034 1428 1038 1431
rect 1042 1428 1110 1431
rect 1114 1428 1126 1431
rect 1210 1428 1694 1431
rect 1698 1428 1798 1431
rect 762 1418 766 1421
rect 826 1418 974 1421
rect 1058 1418 1134 1421
rect 1178 1418 1414 1421
rect 1418 1418 1438 1421
rect 1526 1418 1534 1421
rect 1538 1418 1670 1421
rect 1682 1418 1718 1421
rect 1722 1418 1742 1421
rect 546 1408 1206 1411
rect 1474 1408 1558 1411
rect 1562 1408 1998 1411
rect 376 1403 378 1407
rect 382 1403 385 1407
rect 390 1403 392 1407
rect 1392 1403 1394 1407
rect 1398 1403 1401 1407
rect 1406 1403 1408 1407
rect 402 1398 518 1401
rect 770 1398 790 1401
rect 794 1398 926 1401
rect 1530 1398 1534 1401
rect 266 1388 398 1391
rect 770 1388 934 1391
rect 946 1388 1030 1391
rect 1230 1388 1614 1391
rect 1230 1382 1233 1388
rect 2110 1382 2113 1388
rect 314 1378 326 1381
rect 386 1378 430 1381
rect 514 1378 1118 1381
rect 1138 1378 1198 1381
rect 1298 1378 1446 1381
rect 1546 1378 1638 1381
rect 1270 1372 1273 1378
rect 346 1368 510 1371
rect 818 1368 942 1371
rect 1018 1368 1054 1371
rect 1174 1368 1214 1371
rect 1330 1368 1358 1371
rect 1458 1368 1542 1371
rect 1546 1368 1558 1371
rect 1730 1368 1798 1371
rect 1846 1368 1878 1371
rect 2034 1368 2078 1371
rect 210 1358 270 1361
rect 278 1361 281 1368
rect 622 1362 625 1368
rect 1174 1362 1177 1368
rect 278 1358 318 1361
rect 402 1358 438 1361
rect 722 1358 726 1361
rect 858 1358 942 1361
rect 1034 1358 1062 1361
rect 1170 1358 1174 1361
rect 1202 1358 1246 1361
rect 1250 1358 1278 1361
rect 1310 1361 1313 1368
rect 1282 1358 1313 1361
rect 1410 1358 1414 1361
rect 1430 1361 1433 1368
rect 1846 1362 1849 1368
rect 1974 1362 1977 1368
rect 1982 1362 1985 1368
rect 1430 1358 1446 1361
rect 1458 1358 1478 1361
rect 1570 1358 1582 1361
rect 1786 1358 1846 1361
rect 1866 1358 1926 1361
rect 2010 1358 2062 1361
rect 2070 1358 2078 1361
rect 2082 1358 2142 1361
rect 630 1352 633 1358
rect 122 1348 150 1351
rect 154 1348 230 1351
rect 250 1348 254 1351
rect 338 1348 406 1351
rect 458 1348 494 1351
rect 690 1348 726 1351
rect 786 1348 798 1351
rect 802 1348 806 1351
rect 850 1348 902 1351
rect 930 1348 966 1351
rect 994 1348 1014 1351
rect 1026 1348 1046 1351
rect 1050 1348 1054 1351
rect 1058 1348 1086 1351
rect 1198 1351 1201 1358
rect 1350 1352 1353 1358
rect 1154 1348 1201 1351
rect 1242 1348 1270 1351
rect 1274 1348 1278 1351
rect 1386 1348 1390 1351
rect 1442 1348 1510 1351
rect 1514 1348 1734 1351
rect 1738 1348 1766 1351
rect 1786 1348 1806 1351
rect 1810 1348 1822 1351
rect 1826 1348 2046 1351
rect 2050 1348 2062 1351
rect 2074 1348 2078 1351
rect 2334 1351 2338 1352
rect 2306 1348 2338 1351
rect 42 1338 126 1341
rect 294 1341 297 1348
rect 218 1338 297 1341
rect 362 1338 390 1341
rect 434 1338 446 1341
rect 466 1338 486 1341
rect 646 1341 649 1348
rect 1366 1342 1369 1348
rect 578 1338 649 1341
rect 754 1338 798 1341
rect 834 1338 950 1341
rect 1018 1338 1110 1341
rect 1138 1338 1158 1341
rect 1162 1338 1190 1341
rect 1242 1338 1254 1341
rect 1378 1338 1382 1341
rect 1386 1338 1414 1341
rect 1466 1338 1606 1341
rect 1634 1338 1646 1341
rect 1662 1338 1670 1341
rect 1674 1338 1686 1341
rect 1770 1338 1774 1341
rect 1834 1338 1838 1341
rect 1842 1338 2070 1341
rect 2074 1338 2182 1341
rect 2186 1338 2286 1341
rect 258 1328 782 1331
rect 786 1328 822 1331
rect 978 1328 1070 1331
rect 1074 1328 1102 1331
rect 1110 1331 1113 1338
rect 1438 1332 1441 1338
rect 1110 1328 1246 1331
rect 1290 1328 1430 1331
rect 1450 1328 1470 1331
rect 1578 1328 1582 1331
rect 1586 1328 1702 1331
rect 1738 1328 1742 1331
rect 1746 1328 1894 1331
rect 1946 1328 1958 1331
rect 2042 1328 2214 1331
rect 138 1318 190 1321
rect 194 1318 470 1321
rect 570 1318 598 1321
rect 738 1318 750 1321
rect 794 1318 1126 1321
rect 1130 1318 1182 1321
rect 1250 1318 1326 1321
rect 1330 1318 1494 1321
rect 1570 1318 1710 1321
rect 2014 1321 2017 1328
rect 1938 1318 2017 1321
rect 2074 1318 2262 1321
rect 482 1308 614 1311
rect 954 1308 1158 1311
rect 1170 1308 1374 1311
rect 1386 1308 1454 1311
rect 1478 1308 1598 1311
rect 1602 1308 1638 1311
rect 1674 1308 1902 1311
rect 1962 1308 1966 1311
rect 1978 1308 2086 1311
rect 150 1302 153 1308
rect 880 1303 882 1307
rect 886 1303 889 1307
rect 894 1303 896 1307
rect 34 1298 150 1301
rect 514 1298 662 1301
rect 666 1298 766 1301
rect 1122 1298 1134 1301
rect 1478 1301 1481 1308
rect 1912 1303 1914 1307
rect 1918 1303 1921 1307
rect 1926 1303 1928 1307
rect 1154 1298 1481 1301
rect 1490 1298 1526 1301
rect 1530 1298 1590 1301
rect 1658 1298 1694 1301
rect 2002 1298 2078 1301
rect 106 1288 134 1291
rect 434 1288 478 1291
rect 534 1288 550 1291
rect 994 1288 1278 1291
rect 1426 1288 1454 1291
rect 1834 1288 1897 1291
rect 1906 1288 2030 1291
rect 2138 1288 2182 1291
rect 534 1282 537 1288
rect 50 1278 118 1281
rect 202 1278 238 1281
rect 482 1278 486 1281
rect 562 1278 630 1281
rect 742 1281 745 1288
rect 1894 1282 1897 1288
rect 742 1278 758 1281
rect 774 1278 1062 1281
rect 1098 1278 1166 1281
rect 1218 1278 1294 1281
rect 1346 1278 1382 1281
rect 1522 1278 1790 1281
rect 2010 1278 2110 1281
rect 118 1271 121 1278
rect 774 1272 777 1278
rect 118 1268 182 1271
rect 318 1268 486 1271
rect 514 1268 534 1271
rect 546 1268 638 1271
rect 642 1268 646 1271
rect 818 1268 862 1271
rect 994 1268 1014 1271
rect 1018 1268 1030 1271
rect 1034 1268 1038 1271
rect 1090 1268 1142 1271
rect 1154 1268 1174 1271
rect 1178 1268 1198 1271
rect 1434 1268 1438 1271
rect 1446 1271 1449 1278
rect 1446 1268 1470 1271
rect 1594 1268 1630 1271
rect 1658 1268 1742 1271
rect 1778 1268 1838 1271
rect 1878 1271 1881 1278
rect 1878 1268 1966 1271
rect 2178 1268 2182 1271
rect 318 1262 321 1268
rect 34 1258 134 1261
rect 202 1258 286 1261
rect 370 1258 446 1261
rect 530 1258 542 1261
rect 562 1258 598 1261
rect 602 1258 606 1261
rect 930 1258 1006 1261
rect 1018 1258 1182 1261
rect 1202 1258 1206 1261
rect 1210 1258 1238 1261
rect 1358 1261 1361 1268
rect 2102 1262 2105 1268
rect 1306 1258 1361 1261
rect 1434 1258 1494 1261
rect 1690 1258 1806 1261
rect 1890 1258 1902 1261
rect 1914 1258 1990 1261
rect 1994 1258 2001 1261
rect 2034 1258 2046 1261
rect 2050 1258 2078 1261
rect 2166 1258 2174 1261
rect 2178 1258 2238 1261
rect 22 1248 94 1251
rect 122 1248 262 1251
rect 266 1248 446 1251
rect 634 1248 790 1251
rect 794 1248 822 1251
rect 970 1248 998 1251
rect 1010 1248 1030 1251
rect 1042 1248 1110 1251
rect 1122 1248 1142 1251
rect 1154 1248 1166 1251
rect 1170 1248 1174 1251
rect 1186 1248 1214 1251
rect 1250 1248 1350 1251
rect 1354 1248 1366 1251
rect 1386 1248 1390 1251
rect 1394 1248 1462 1251
rect 1622 1251 1625 1258
rect 1610 1248 1625 1251
rect 1690 1248 1694 1251
rect 1706 1248 1710 1251
rect 1858 1248 1897 1251
rect 1986 1248 2030 1251
rect 2162 1248 2182 1251
rect 2334 1251 2338 1252
rect 2306 1248 2338 1251
rect 22 1242 25 1248
rect 1894 1242 1897 1248
rect 818 1238 918 1241
rect 922 1238 1030 1241
rect 1050 1238 1070 1241
rect 1082 1238 1102 1241
rect 1106 1238 1414 1241
rect 1426 1238 1478 1241
rect 1658 1238 1662 1241
rect 1674 1238 1838 1241
rect 2258 1238 2294 1241
rect 314 1228 470 1231
rect 474 1228 494 1231
rect 674 1228 1246 1231
rect 1266 1228 1646 1231
rect 1650 1228 1750 1231
rect 1754 1228 1774 1231
rect 250 1218 294 1221
rect 1090 1218 1102 1221
rect 1130 1218 1158 1221
rect 1202 1218 1358 1221
rect 1362 1218 1438 1221
rect 1890 1218 2022 1221
rect 2026 1218 2054 1221
rect 978 1208 1054 1211
rect 1082 1208 1193 1211
rect 1202 1208 1374 1211
rect 1426 1208 1558 1211
rect 376 1203 378 1207
rect 382 1203 385 1207
rect 390 1203 392 1207
rect 834 1198 926 1201
rect 930 1198 1022 1201
rect 1090 1198 1134 1201
rect 1190 1201 1193 1208
rect 1392 1203 1394 1207
rect 1398 1203 1401 1207
rect 1406 1203 1408 1207
rect 1190 1198 1350 1201
rect 1538 1198 1622 1201
rect 1866 1198 1894 1201
rect 146 1188 1262 1191
rect 1466 1188 1646 1191
rect 146 1178 230 1181
rect 466 1178 486 1181
rect 594 1178 990 1181
rect 1114 1178 1118 1181
rect 1138 1178 1270 1181
rect 1274 1178 1542 1181
rect 1546 1178 1550 1181
rect 1850 1178 1974 1181
rect 146 1168 177 1171
rect 298 1168 310 1171
rect 406 1171 409 1178
rect 378 1168 409 1171
rect 502 1172 505 1178
rect 1014 1172 1017 1178
rect 594 1168 614 1171
rect 718 1168 742 1171
rect 1042 1168 1094 1171
rect 1122 1168 1126 1171
rect 1162 1168 1190 1171
rect 1194 1168 1230 1171
rect 1378 1168 1446 1171
rect 1638 1168 1886 1171
rect 1930 1168 2014 1171
rect 2018 1168 2286 1171
rect 174 1162 177 1168
rect 718 1162 721 1168
rect 1254 1162 1257 1168
rect 1558 1162 1561 1168
rect 1638 1162 1641 1168
rect 178 1158 206 1161
rect 274 1158 358 1161
rect 362 1158 510 1161
rect 802 1158 830 1161
rect 834 1158 926 1161
rect 1058 1158 1086 1161
rect 1090 1158 1198 1161
rect 1442 1158 1462 1161
rect 1522 1158 1526 1161
rect 1602 1158 1606 1161
rect 1662 1158 1670 1161
rect 1674 1158 1750 1161
rect 2106 1158 2110 1161
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 78 1151 81 1158
rect 78 1148 166 1151
rect 258 1148 278 1151
rect 282 1148 286 1151
rect 418 1148 470 1151
rect 502 1148 566 1151
rect 650 1148 654 1151
rect 690 1148 694 1151
rect 790 1151 793 1158
rect 1022 1152 1025 1158
rect 1046 1152 1049 1158
rect 1278 1152 1281 1158
rect 1638 1152 1641 1158
rect 1758 1152 1761 1158
rect 1830 1152 1833 1158
rect 786 1148 793 1151
rect 502 1142 505 1148
rect 890 1148 966 1151
rect 1034 1148 1038 1151
rect 1058 1148 1142 1151
rect 1178 1148 1214 1151
rect 1314 1148 1422 1151
rect 1426 1148 1478 1151
rect 1498 1148 1510 1151
rect 1514 1148 1518 1151
rect 1658 1148 1662 1151
rect 1850 1148 1862 1151
rect 1958 1151 1961 1158
rect 2166 1152 2169 1158
rect 1882 1148 1961 1151
rect 2058 1148 2078 1151
rect 2082 1148 2102 1151
rect 178 1138 190 1141
rect 234 1138 270 1141
rect 274 1138 302 1141
rect 410 1138 462 1141
rect 622 1138 689 1141
rect 150 1132 153 1138
rect 202 1128 262 1131
rect 326 1131 329 1138
rect 266 1128 329 1131
rect 350 1132 353 1138
rect 622 1132 625 1138
rect 686 1132 689 1138
rect 794 1138 1038 1141
rect 1186 1138 1214 1141
rect 1218 1138 1230 1141
rect 1418 1138 1486 1141
rect 1490 1138 1502 1141
rect 1590 1141 1593 1148
rect 1562 1138 1593 1141
rect 1642 1138 1670 1141
rect 1674 1138 1745 1141
rect 1754 1138 1854 1141
rect 2050 1138 2086 1141
rect 2194 1138 2230 1141
rect 782 1132 785 1138
rect 642 1128 646 1131
rect 770 1128 774 1131
rect 962 1128 982 1131
rect 986 1128 1062 1131
rect 1098 1128 1102 1131
rect 1106 1128 1126 1131
rect 1170 1128 1198 1131
rect 1394 1128 1422 1131
rect 1490 1128 1574 1131
rect 1618 1128 1654 1131
rect 1658 1128 1686 1131
rect 1742 1131 1745 1138
rect 1742 1128 1766 1131
rect 1770 1128 1798 1131
rect 214 1118 222 1121
rect 226 1118 254 1121
rect 490 1118 534 1121
rect 538 1118 574 1121
rect 670 1121 673 1128
rect 650 1118 742 1121
rect 746 1118 774 1121
rect 778 1118 806 1121
rect 1010 1118 1142 1121
rect 1154 1118 1190 1121
rect 1198 1121 1201 1128
rect 1198 1118 1486 1121
rect 1554 1118 1678 1121
rect 1786 1118 1838 1121
rect 1922 1118 2046 1121
rect 430 1112 433 1118
rect 2278 1112 2281 1118
rect 482 1108 694 1111
rect 738 1108 742 1111
rect 994 1108 1377 1111
rect 1498 1108 1518 1111
rect 1546 1108 1790 1111
rect 1810 1108 1838 1111
rect 880 1103 882 1107
rect 886 1103 889 1107
rect 894 1103 896 1107
rect 1374 1102 1377 1108
rect 1912 1103 1914 1107
rect 1918 1103 1921 1107
rect 1926 1103 1928 1107
rect 298 1098 518 1101
rect 610 1098 654 1101
rect 1042 1098 1054 1101
rect 1066 1098 1182 1101
rect 1186 1098 1190 1101
rect 1298 1098 1350 1101
rect 1378 1098 1470 1101
rect 1474 1098 1502 1101
rect 1506 1098 1710 1101
rect 1714 1098 1862 1101
rect 2042 1098 2222 1101
rect 2226 1098 2286 1101
rect 10 1088 30 1091
rect 234 1088 262 1091
rect 566 1091 569 1098
rect 566 1088 590 1091
rect 986 1088 1030 1091
rect 1034 1088 1094 1091
rect 1146 1088 1246 1091
rect 1266 1088 1286 1091
rect 1418 1088 1518 1091
rect 1586 1088 1678 1091
rect 1698 1088 2030 1091
rect 2074 1088 2078 1091
rect 18 1078 22 1081
rect 26 1078 33 1081
rect 90 1078 158 1081
rect 162 1078 198 1081
rect 246 1078 310 1081
rect 858 1078 990 1081
rect 1066 1078 1286 1081
rect 1314 1078 1390 1081
rect 1490 1078 1622 1081
rect 1626 1078 1766 1081
rect 2034 1078 2241 1081
rect 2290 1078 2294 1081
rect 34 1068 38 1071
rect 78 1068 86 1071
rect 194 1068 238 1071
rect 246 1071 249 1078
rect 242 1068 249 1071
rect 410 1068 486 1071
rect 530 1068 606 1071
rect 738 1068 782 1071
rect 786 1068 814 1071
rect 1062 1071 1065 1078
rect 1806 1072 1809 1078
rect 946 1068 1065 1071
rect 1178 1068 1214 1071
rect 1218 1068 1230 1071
rect 1266 1068 1358 1071
rect 1498 1068 1566 1071
rect 1570 1068 1582 1071
rect 1594 1068 1598 1071
rect 1602 1068 1638 1071
rect 1666 1068 1670 1071
rect 1682 1068 1782 1071
rect 1818 1068 1870 1071
rect 1898 1068 1974 1071
rect 2074 1068 2078 1071
rect 2238 1071 2241 1078
rect 2334 1071 2338 1072
rect 2238 1068 2338 1071
rect 78 1061 81 1068
rect 50 1058 81 1061
rect 150 1061 153 1068
rect 254 1062 257 1068
rect 1798 1062 1801 1068
rect 150 1058 222 1061
rect 322 1058 366 1061
rect 370 1058 438 1061
rect 674 1058 838 1061
rect 946 1058 982 1061
rect 1002 1058 1017 1061
rect 1014 1052 1017 1058
rect 1206 1058 1222 1061
rect 1458 1058 1470 1061
rect 1554 1058 1566 1061
rect 1578 1058 1582 1061
rect 1634 1058 1646 1061
rect 1802 1058 1814 1061
rect 1890 1058 1894 1061
rect 2106 1058 2142 1061
rect 1206 1052 1209 1058
rect 1830 1052 1833 1058
rect 82 1048 198 1051
rect 210 1048 230 1051
rect 618 1048 630 1051
rect 738 1048 833 1051
rect 922 1048 998 1051
rect 1018 1048 1022 1051
rect 1262 1048 1358 1051
rect 1378 1048 1414 1051
rect 1458 1048 1462 1051
rect 1530 1048 1534 1051
rect 1642 1048 1726 1051
rect 1746 1048 1806 1051
rect 1874 1048 1902 1051
rect 2082 1048 2110 1051
rect 230 1042 233 1048
rect 830 1042 833 1048
rect 1262 1042 1265 1048
rect 1574 1042 1577 1048
rect 1862 1042 1865 1048
rect 10 1038 190 1041
rect 282 1038 502 1041
rect 610 1038 758 1041
rect 1162 1038 1206 1041
rect 1378 1038 1438 1041
rect 1594 1038 1598 1041
rect 122 1028 142 1031
rect 146 1028 438 1031
rect 442 1028 686 1031
rect 830 1031 833 1038
rect 830 1028 942 1031
rect 1362 1028 1446 1031
rect 1522 1028 1630 1031
rect 98 1018 198 1021
rect 202 1018 214 1021
rect 462 1018 470 1021
rect 474 1018 638 1021
rect 690 1018 766 1021
rect 770 1018 862 1021
rect 954 1018 998 1021
rect 1010 1018 1166 1021
rect 1170 1018 1214 1021
rect 1218 1018 1606 1021
rect 66 1008 174 1011
rect 178 1008 342 1011
rect 402 1008 638 1011
rect 642 1008 742 1011
rect 754 1008 950 1011
rect 1010 1008 1070 1011
rect 1122 1008 1206 1011
rect 1274 1008 1294 1011
rect 1498 1008 1510 1011
rect 1586 1008 1614 1011
rect 1738 1008 2070 1011
rect 2074 1008 2262 1011
rect 376 1003 378 1007
rect 382 1003 385 1007
rect 390 1003 392 1007
rect 1392 1003 1394 1007
rect 1398 1003 1401 1007
rect 1406 1003 1408 1007
rect 442 998 526 1001
rect 762 998 974 1001
rect 978 998 1078 1001
rect 1082 998 1134 1001
rect 290 988 438 991
rect 778 988 902 991
rect 906 988 942 991
rect 954 988 1022 991
rect 1050 988 1118 991
rect 1138 988 1270 991
rect 1274 988 1486 991
rect 1514 988 1854 991
rect 1858 988 1902 991
rect 338 978 446 981
rect 698 978 718 981
rect 722 978 958 981
rect 1018 978 1078 981
rect 1090 978 1142 981
rect 1146 978 1158 981
rect 1186 978 1190 981
rect 1194 978 1230 981
rect 1426 978 1438 981
rect 1442 978 1486 981
rect 1490 978 1662 981
rect 1666 978 1758 981
rect 1762 978 2014 981
rect 210 968 294 971
rect 338 968 406 971
rect 514 968 518 971
rect 546 968 574 971
rect 642 968 726 971
rect 730 968 774 971
rect 842 968 910 971
rect 930 968 934 971
rect 954 968 1006 971
rect 1226 968 1457 971
rect 1482 968 1550 971
rect 1746 968 1814 971
rect 1986 968 2134 971
rect 2138 968 2270 971
rect 2334 971 2338 972
rect 2306 968 2338 971
rect 1046 962 1049 968
rect 18 958 102 961
rect 130 958 142 961
rect 170 958 190 961
rect 314 958 350 961
rect 354 958 630 961
rect 634 958 806 961
rect 822 958 854 961
rect 954 958 969 961
rect 1142 961 1145 968
rect 1066 958 1145 961
rect 1162 958 1246 961
rect 1290 958 1326 961
rect 1426 958 1446 961
rect 1454 961 1457 968
rect 1454 958 1566 961
rect 1690 958 1918 961
rect 1970 958 2022 961
rect 2026 958 2030 961
rect 2042 958 2238 961
rect 66 948 126 951
rect 146 948 150 951
rect 194 948 246 951
rect 626 948 694 951
rect 822 951 825 958
rect 966 952 969 958
rect 786 948 825 951
rect 834 948 894 951
rect 914 948 926 951
rect 986 948 990 951
rect 1022 948 1246 951
rect 1250 948 1278 951
rect 1282 948 1382 951
rect 1434 948 1470 951
rect 1522 948 1526 951
rect 1722 948 1806 951
rect 1810 948 1830 951
rect 1834 948 1854 951
rect 1874 948 1878 951
rect 1882 948 1942 951
rect 1954 948 1974 951
rect 2002 948 2046 951
rect 2066 948 2086 951
rect 86 938 110 941
rect 114 938 246 941
rect 306 938 318 941
rect 470 941 473 948
rect 542 942 545 948
rect 418 938 473 941
rect 490 938 542 941
rect 1022 941 1025 948
rect 2102 948 2177 951
rect 2334 951 2338 952
rect 2266 948 2338 951
rect 810 938 1025 941
rect 1034 938 1094 941
rect 1138 938 1198 941
rect 1202 938 1214 941
rect 1218 938 1542 941
rect 1794 938 1854 941
rect 1858 938 1870 941
rect 2002 938 2006 941
rect 2102 941 2105 948
rect 2174 942 2177 948
rect 2026 938 2105 941
rect 2114 938 2161 941
rect 86 932 89 938
rect 146 928 150 931
rect 318 928 326 931
rect 330 928 550 931
rect 574 931 577 938
rect 2158 932 2161 938
rect 574 928 622 931
rect 642 928 694 931
rect 762 928 958 931
rect 962 928 982 931
rect 1082 928 1126 931
rect 1258 928 1262 931
rect 1298 928 1326 931
rect 1330 928 2046 931
rect 266 918 406 921
rect 498 918 550 921
rect 554 918 1014 921
rect 1042 918 1086 921
rect 1090 918 1158 921
rect 1206 921 1209 928
rect 1162 918 1209 921
rect 1306 918 1318 921
rect 1362 918 1366 921
rect 1610 918 1630 921
rect 1834 918 1918 921
rect 122 908 126 911
rect 306 908 462 911
rect 522 908 758 911
rect 778 908 798 911
rect 1002 908 1006 911
rect 1522 908 1550 911
rect 1634 908 1654 911
rect 1674 908 1694 911
rect 880 903 882 907
rect 886 903 889 907
rect 894 903 896 907
rect 1912 903 1914 907
rect 1918 903 1921 907
rect 1926 903 1928 907
rect 138 898 310 901
rect 426 898 438 901
rect 442 898 606 901
rect 1098 898 1174 901
rect 1482 898 1494 901
rect 1546 898 1798 901
rect 1842 898 1846 901
rect 1898 898 1902 901
rect 2090 898 2278 901
rect 122 888 166 891
rect 178 888 273 891
rect 290 888 374 891
rect 378 888 414 891
rect 434 888 438 891
rect 530 888 574 891
rect 634 888 686 891
rect 802 888 830 891
rect 898 888 934 891
rect 1178 888 1182 891
rect 1206 888 1214 891
rect 1218 888 1246 891
rect 1258 888 1294 891
rect 1322 888 1406 891
rect 1474 888 1494 891
rect 1530 888 1534 891
rect 1618 888 1662 891
rect 1798 891 1801 898
rect 1798 888 1830 891
rect 1834 888 1926 891
rect 1930 888 2022 891
rect 2194 888 2238 891
rect 270 882 273 888
rect 98 878 134 881
rect 170 878 262 881
rect 274 878 398 881
rect 426 878 518 881
rect 538 878 558 881
rect 570 878 630 881
rect 634 878 782 881
rect 834 878 942 881
rect 946 878 950 881
rect 986 878 1046 881
rect 1142 881 1145 888
rect 1766 882 1769 888
rect 1142 878 1166 881
rect 1210 878 1238 881
rect 1354 878 1470 881
rect 1474 878 1542 881
rect 1554 878 1574 881
rect 1658 878 1694 881
rect 1794 878 1838 881
rect 1898 878 1974 881
rect 262 872 265 878
rect 130 868 214 871
rect 650 868 654 871
rect 682 868 894 871
rect 906 868 950 871
rect 986 868 1014 871
rect 1050 868 1262 871
rect 1266 868 1342 871
rect 1378 868 1446 871
rect 1530 868 1558 871
rect 1570 868 1574 871
rect 1594 868 1598 871
rect 1690 868 1718 871
rect 1722 868 1742 871
rect 1746 868 1990 871
rect 2222 871 2225 878
rect 2138 868 2225 871
rect 58 858 110 861
rect 178 858 206 861
rect 266 859 326 861
rect 266 858 329 859
rect 474 858 545 861
rect 634 858 638 861
rect 674 858 734 861
rect 766 858 830 861
rect 906 858 910 861
rect 978 858 1046 861
rect 1050 858 1102 861
rect 1114 858 1438 861
rect 1442 858 1454 861
rect 1458 858 1782 861
rect 1794 858 1806 861
rect 1962 858 2030 861
rect 2242 858 2254 861
rect 542 852 545 858
rect 766 852 769 858
rect 114 848 142 851
rect 162 848 238 851
rect 266 848 273 851
rect 394 848 414 851
rect 858 848 918 851
rect 954 848 958 851
rect 978 848 982 851
rect 1170 848 1526 851
rect 1546 848 1622 851
rect 1642 848 1662 851
rect 1666 848 1686 851
rect 1754 848 1798 851
rect 1838 851 1841 858
rect 2078 852 2081 858
rect 1826 848 1841 851
rect 1866 848 1870 851
rect 1938 848 1958 851
rect 2194 848 2230 851
rect 2234 848 2270 851
rect 2334 851 2338 852
rect 2306 848 2338 851
rect 270 842 273 848
rect 1534 842 1537 848
rect 1958 842 1961 848
rect 106 838 150 841
rect 282 838 478 841
rect 570 838 598 841
rect 946 838 1126 841
rect 1602 838 1638 841
rect 1674 838 1718 841
rect 1730 838 1758 841
rect 1770 838 1806 841
rect 1810 838 1862 841
rect 2210 838 2270 841
rect 250 828 270 831
rect 274 828 302 831
rect 306 828 438 831
rect 450 828 462 831
rect 466 828 750 831
rect 754 828 1078 831
rect 1858 828 1934 831
rect 426 818 446 821
rect 618 818 638 821
rect 1786 818 1878 821
rect 1034 808 1134 811
rect 1642 808 1830 811
rect 376 803 378 807
rect 382 803 385 807
rect 390 803 392 807
rect 1392 803 1394 807
rect 1398 803 1401 807
rect 1406 803 1408 807
rect 1802 798 2174 801
rect 2178 798 2198 801
rect 210 788 310 791
rect 314 788 350 791
rect 466 788 502 791
rect 506 788 662 791
rect 986 788 998 791
rect 1002 788 1094 791
rect 1274 788 1446 791
rect 2002 788 2094 791
rect 194 778 358 781
rect 498 778 598 781
rect 730 778 1070 781
rect 1074 778 1430 781
rect 1434 778 1454 781
rect 1458 778 2038 781
rect 2042 778 2238 781
rect 110 771 113 778
rect 50 768 113 771
rect 146 768 166 771
rect 170 768 190 771
rect 218 768 254 771
rect 514 768 614 771
rect 826 768 934 771
rect 1186 768 1374 771
rect 1378 768 1478 771
rect 1726 768 1734 771
rect 1738 768 1766 771
rect 1794 768 1798 771
rect 1850 768 1878 771
rect 1906 768 1918 771
rect 1962 768 2070 771
rect 2074 768 2158 771
rect 2334 771 2338 772
rect 2306 768 2338 771
rect 1486 762 1489 768
rect 98 758 150 761
rect 154 758 366 761
rect 434 758 502 761
rect 506 758 510 761
rect 546 758 574 761
rect 610 758 662 761
rect 746 758 822 761
rect 842 758 854 761
rect 1034 758 1102 761
rect 1210 758 1214 761
rect 1306 758 1366 761
rect 1514 758 1726 761
rect 1818 758 1830 761
rect 1866 758 2006 761
rect 2010 758 2014 761
rect 2026 758 2118 761
rect 422 752 425 758
rect 186 748 246 751
rect 266 748 310 751
rect 346 748 422 751
rect 434 748 438 751
rect 602 748 622 751
rect 662 751 665 758
rect 662 748 686 751
rect 742 751 745 758
rect 698 748 745 751
rect 866 748 950 751
rect 994 748 1009 751
rect 1042 748 1078 751
rect 1146 748 1150 751
rect 1202 748 1238 751
rect 1242 748 1262 751
rect 1354 748 1382 751
rect 1386 748 1430 751
rect 1438 751 1441 758
rect 1438 748 1510 751
rect 1522 748 1734 751
rect 1826 748 1838 751
rect 1866 748 1870 751
rect 1882 748 1974 751
rect 2022 751 2025 758
rect 2022 748 2030 751
rect 2050 748 2054 751
rect 2126 751 2129 758
rect 2126 748 2174 751
rect 2334 751 2338 752
rect 2306 748 2338 751
rect 1006 742 1009 748
rect 1118 742 1121 748
rect 298 738 302 741
rect 306 738 382 741
rect 414 738 422 741
rect 426 738 446 741
rect 490 738 494 741
rect 618 738 638 741
rect 658 738 662 741
rect 690 738 750 741
rect 762 738 790 741
rect 794 738 806 741
rect 1058 738 1086 741
rect 1194 738 1198 741
rect 1226 738 1230 741
rect 1234 738 1342 741
rect 1346 738 1414 741
rect 1470 738 1534 741
rect 1562 738 1598 741
rect 1754 738 1982 741
rect 1986 738 1990 741
rect 2202 738 2217 741
rect 1094 732 1097 738
rect 1470 732 1473 738
rect 2214 732 2217 738
rect 402 728 438 731
rect 562 728 654 731
rect 730 728 830 731
rect 954 728 1046 731
rect 1762 728 1774 731
rect 1834 728 1838 731
rect 1970 728 2014 731
rect 2114 728 2190 731
rect 2194 728 2206 731
rect 106 718 110 721
rect 114 718 134 721
rect 138 718 166 721
rect 394 718 406 721
rect 418 718 422 721
rect 682 718 870 721
rect 874 718 1022 721
rect 1098 718 1134 721
rect 1174 721 1177 728
rect 1142 718 1177 721
rect 1354 718 1398 721
rect 1402 718 1510 721
rect 1538 718 1558 721
rect 1658 718 1774 721
rect 1858 718 2030 721
rect 2034 718 2102 721
rect 2106 718 2182 721
rect 130 708 350 711
rect 354 708 558 711
rect 1058 708 1062 711
rect 1142 711 1145 718
rect 1066 708 1145 711
rect 1170 708 1254 711
rect 1434 708 1582 711
rect 1770 708 1886 711
rect 880 703 882 707
rect 886 703 889 707
rect 894 703 896 707
rect 1912 703 1914 707
rect 1918 703 1921 707
rect 1926 703 1928 707
rect 458 698 526 701
rect 626 698 638 701
rect 962 698 1110 701
rect 1114 698 1134 701
rect 1146 698 1294 701
rect 1306 698 1518 701
rect 1690 698 1710 701
rect 1722 698 1830 701
rect 1834 698 1905 701
rect 2050 698 2270 701
rect 322 688 358 691
rect 586 688 590 691
rect 594 688 686 691
rect 1050 688 1054 691
rect 1086 688 1486 691
rect 1494 688 1502 691
rect 1506 688 1574 691
rect 1586 688 1590 691
rect 1610 688 1654 691
rect 1682 688 1686 691
rect 1694 688 1702 691
rect 1706 688 1710 691
rect 1722 688 1878 691
rect 1902 691 1905 698
rect 1902 688 2286 691
rect 1086 682 1089 688
rect 138 678 174 681
rect 362 678 366 681
rect 594 678 646 681
rect 1026 678 1030 681
rect 1130 678 1158 681
rect 1162 678 1198 681
rect 1282 678 1422 681
rect 1458 678 1854 681
rect 218 668 310 671
rect 354 668 454 671
rect 758 671 761 678
rect 650 668 761 671
rect 774 671 777 678
rect 958 672 961 678
rect 998 672 1001 678
rect 774 668 878 671
rect 1010 668 1014 671
rect 1130 668 1158 671
rect 1170 668 1193 671
rect 1218 668 1230 671
rect 1290 668 1542 671
rect 1562 668 1566 671
rect 1578 668 1638 671
rect 1682 668 1726 671
rect 1730 668 1742 671
rect 1762 668 1766 671
rect 1862 671 1865 678
rect 1842 668 1865 671
rect 98 658 134 661
rect 322 658 470 661
rect 562 658 662 661
rect 754 658 814 661
rect 890 658 982 661
rect 1030 658 1038 661
rect 1042 658 1062 661
rect 1130 658 1134 661
rect 1162 658 1182 661
rect 1190 661 1193 668
rect 1190 658 1334 661
rect 1418 658 1422 661
rect 1426 658 1454 661
rect 1498 658 1894 661
rect 1898 658 1902 661
rect 2042 658 2078 661
rect 2098 658 2166 661
rect -26 651 -22 652
rect -26 648 6 651
rect 178 648 206 651
rect 426 648 430 651
rect 538 648 630 651
rect 690 648 734 651
rect 738 648 750 651
rect 754 648 766 651
rect 938 648 1030 651
rect 1034 648 1046 651
rect 1082 648 1174 651
rect 1178 648 1278 651
rect 1362 648 1414 651
rect 1462 651 1465 658
rect 2246 652 2249 658
rect 1462 648 1486 651
rect 1658 648 1710 651
rect 1714 648 1726 651
rect 2002 648 2046 651
rect 2098 648 2102 651
rect 10 638 38 641
rect 42 638 374 641
rect 378 638 430 641
rect 670 641 673 648
rect 626 638 710 641
rect 1090 638 1102 641
rect 1218 638 1222 641
rect 1450 638 1518 641
rect 1638 641 1641 648
rect 1862 642 1865 648
rect 1638 638 1678 641
rect 1938 638 1942 641
rect 2018 638 2126 641
rect 2130 638 2137 641
rect 298 628 398 631
rect 586 628 766 631
rect 914 628 1094 631
rect 1226 628 1262 631
rect 1450 628 1630 631
rect 1778 628 1998 631
rect 2106 628 2110 631
rect 2114 628 2294 631
rect 470 621 473 628
rect 470 618 1622 621
rect 2114 618 2142 621
rect 706 608 1105 611
rect 1114 608 1382 611
rect 1434 608 1910 611
rect 376 603 378 607
rect 382 603 385 607
rect 390 603 392 607
rect 170 598 174 601
rect 450 598 590 601
rect 594 598 614 601
rect 618 598 726 601
rect 794 598 806 601
rect 850 598 942 601
rect 1102 601 1105 608
rect 1392 603 1394 607
rect 1398 603 1401 607
rect 1406 603 1408 607
rect 1102 598 1166 601
rect 1554 598 1606 601
rect 1898 598 1934 601
rect 1938 598 2062 601
rect 434 588 718 591
rect 794 588 1158 591
rect 1318 588 1326 591
rect 1330 588 1470 591
rect 1618 588 1662 591
rect 1786 588 2150 591
rect 346 578 550 581
rect 730 578 958 581
rect 970 578 1022 581
rect 1162 578 1206 581
rect 1426 578 1614 581
rect 1618 578 1798 581
rect 1842 578 1886 581
rect 166 571 169 578
rect 74 568 169 571
rect 190 572 193 578
rect 194 568 294 571
rect 306 568 310 571
rect 314 568 350 571
rect 426 568 430 571
rect 458 568 502 571
rect 566 571 569 578
rect 538 568 569 571
rect 658 568 750 571
rect 1034 568 1046 571
rect 1082 568 1094 571
rect 1178 568 1190 571
rect 1214 571 1217 578
rect 1210 568 1217 571
rect 1234 568 1238 571
rect 1290 568 1294 571
rect 1322 568 1326 571
rect 1362 568 1518 571
rect 1654 568 1662 571
rect 1666 568 1742 571
rect 1962 568 2030 571
rect 130 558 206 561
rect 458 558 494 561
rect 498 558 598 561
rect 1042 558 1054 561
rect 1074 558 1118 561
rect 1122 558 1158 561
rect 1210 558 1246 561
rect 1250 558 1350 561
rect 1442 558 1838 561
rect 1906 558 2062 561
rect 2074 558 2134 561
rect 2138 558 2270 561
rect 90 548 150 551
rect 162 548 190 551
rect 274 548 366 551
rect 410 548 462 551
rect 522 548 558 551
rect 774 551 777 558
rect 774 548 1118 551
rect 1122 548 1414 551
rect 1634 548 1646 551
rect 1738 548 1822 551
rect 1846 551 1849 558
rect 1826 548 1849 551
rect 1914 548 1942 551
rect 2010 548 2014 551
rect 2034 548 2094 551
rect 2166 548 2174 551
rect 2178 548 2214 551
rect 34 538 94 541
rect 98 538 150 541
rect 210 538 278 541
rect 330 538 454 541
rect 458 538 462 541
rect 570 538 574 541
rect 614 541 617 548
rect 1478 542 1481 548
rect 614 538 646 541
rect 746 538 782 541
rect 818 538 854 541
rect 874 538 894 541
rect 1186 538 1222 541
rect 1258 538 1262 541
rect 1274 538 1302 541
rect 1346 538 1366 541
rect 1386 538 1462 541
rect 1486 541 1489 548
rect 1486 538 1494 541
rect 1726 541 1729 548
rect 1578 538 1729 541
rect 1858 538 1886 541
rect 2142 538 2286 541
rect 2142 532 2145 538
rect 202 528 286 531
rect 290 528 318 531
rect 322 528 414 531
rect 770 528 846 531
rect 850 528 910 531
rect 1250 528 1254 531
rect 1434 528 1446 531
rect 1454 528 1502 531
rect 1674 528 1790 531
rect 1882 528 2022 531
rect 2026 528 2033 531
rect 1454 522 1457 528
rect 570 518 990 521
rect 1098 518 1230 521
rect 1234 518 1326 521
rect 1330 518 1438 521
rect 1466 518 1694 521
rect 2010 518 2142 521
rect 2146 518 2166 521
rect 154 508 174 511
rect 178 508 326 511
rect 954 508 1190 511
rect 1194 508 1902 511
rect 2018 508 2054 511
rect 880 503 882 507
rect 886 503 889 507
rect 894 503 896 507
rect 1912 503 1914 507
rect 1918 503 1921 507
rect 1926 503 1928 507
rect 218 498 366 501
rect 370 498 446 501
rect 946 498 1014 501
rect 1034 498 1278 501
rect 1282 498 1406 501
rect 1410 498 1478 501
rect 1482 498 1630 501
rect 1634 498 1654 501
rect 1658 498 1662 501
rect 1954 498 2102 501
rect 2114 498 2198 501
rect 474 488 518 491
rect 1002 488 1078 491
rect 1082 488 1086 491
rect 1322 488 1374 491
rect 1514 488 1590 491
rect 1594 488 1678 491
rect 1930 488 1942 491
rect 2042 488 2174 491
rect 2178 488 2190 491
rect 126 481 129 488
rect 42 478 129 481
rect 134 478 158 481
rect 302 481 305 488
rect 226 478 305 481
rect 738 478 950 481
rect 1138 478 1254 481
rect 1258 478 1422 481
rect 1426 478 1470 481
rect 1818 478 2014 481
rect 2058 478 2070 481
rect 2074 478 2086 481
rect 134 471 137 478
rect 106 468 137 471
rect 146 468 478 471
rect 482 468 502 471
rect 818 468 878 471
rect 978 468 1030 471
rect 1810 468 1838 471
rect 1842 468 1966 471
rect 1970 468 2006 471
rect 2010 468 2030 471
rect 2042 468 2118 471
rect 2134 468 2166 471
rect 122 458 134 461
rect 274 458 278 461
rect 298 458 318 461
rect 330 458 334 461
rect 418 458 494 461
rect 586 458 622 461
rect 750 461 753 468
rect 1374 462 1377 468
rect 706 458 753 461
rect 970 458 982 461
rect 1066 458 1177 461
rect 1378 458 1390 461
rect 1394 458 1486 461
rect 1494 461 1497 468
rect 2134 462 2137 468
rect 1494 458 1537 461
rect 1666 458 1734 461
rect 1794 458 2078 461
rect 2082 458 2086 461
rect 2106 458 2129 461
rect 2202 458 2238 461
rect 1174 452 1177 458
rect 1534 452 1537 458
rect 2126 452 2129 458
rect 170 448 350 451
rect 450 448 558 451
rect 650 448 774 451
rect 794 448 806 451
rect 1098 448 1126 451
rect 1330 448 1446 451
rect 1642 448 1670 451
rect 1674 448 2030 451
rect 146 438 526 441
rect 714 438 822 441
rect 826 438 902 441
rect 994 438 1102 441
rect 1210 438 1254 441
rect 1258 438 1358 441
rect 1850 438 1854 441
rect 2074 438 2198 441
rect 1534 432 1537 438
rect 170 428 534 431
rect 538 428 1038 431
rect 1042 428 1126 431
rect 1138 428 1214 431
rect 1506 428 1518 431
rect 66 418 214 421
rect 298 418 590 421
rect 602 418 622 421
rect 810 418 982 421
rect 1106 418 1486 421
rect 1506 418 1574 421
rect 698 408 870 411
rect 1486 411 1489 418
rect 1486 408 1958 411
rect 1962 408 2158 411
rect 376 403 378 407
rect 382 403 385 407
rect 390 403 392 407
rect 1392 403 1394 407
rect 1398 403 1401 407
rect 1406 403 1408 407
rect 770 398 838 401
rect 858 398 1150 401
rect 1554 398 1686 401
rect 410 388 830 391
rect 986 388 1046 391
rect 1050 388 1110 391
rect 1170 388 1369 391
rect 1530 388 1841 391
rect 474 378 598 381
rect 602 378 646 381
rect 1366 381 1369 388
rect 1838 382 1841 388
rect 1106 378 1353 381
rect 1366 378 1606 381
rect 426 368 446 371
rect 730 368 734 371
rect 1030 371 1033 378
rect 1350 372 1353 378
rect 1622 372 1625 378
rect 1638 372 1641 378
rect 1646 372 1649 378
rect 962 368 1033 371
rect 1106 368 1134 371
rect 1250 368 1302 371
rect 1354 368 1414 371
rect 1434 368 1542 371
rect 1674 368 1678 371
rect 1738 368 1806 371
rect 1994 368 2014 371
rect 614 362 617 368
rect 1038 362 1041 368
rect 1614 362 1617 368
rect 2030 362 2033 368
rect 18 358 22 361
rect 186 358 510 361
rect 626 358 654 361
rect 658 358 902 361
rect 1018 358 1038 361
rect 1050 358 1070 361
rect 1074 358 1166 361
rect 1178 358 1182 361
rect 1186 358 1254 361
rect 1258 358 1302 361
rect 1390 358 1398 361
rect 1402 358 1478 361
rect 1602 358 1614 361
rect 1618 358 1742 361
rect 1746 358 1774 361
rect 2010 358 2030 361
rect 2162 358 2174 361
rect 2178 358 2262 361
rect 510 352 513 358
rect 66 348 78 351
rect 138 348 286 351
rect 290 348 326 351
rect 474 348 494 351
rect 498 348 502 351
rect 530 348 566 351
rect 570 348 590 351
rect 610 348 638 351
rect 642 348 790 351
rect 794 348 806 351
rect 826 348 862 351
rect 898 348 990 351
rect 1090 348 1110 351
rect 1138 348 1150 351
rect 1290 348 1313 351
rect 1370 348 1398 351
rect 1402 348 1662 351
rect 1714 348 1782 351
rect 1910 351 1913 358
rect 1982 351 1985 358
rect 1910 348 1985 351
rect 2154 348 2166 351
rect 2186 348 2265 351
rect 38 341 41 348
rect 1030 342 1033 348
rect 1310 342 1313 348
rect 38 338 142 341
rect 242 338 262 341
rect 298 338 302 341
rect 378 338 470 341
rect 522 338 566 341
rect 586 338 710 341
rect 714 338 870 341
rect 1050 338 1158 341
rect 1210 338 1254 341
rect 1346 338 1454 341
rect 1514 338 1526 341
rect 1618 338 1710 341
rect 1998 341 2001 348
rect 2150 341 2153 348
rect 1906 338 2153 341
rect 2262 342 2265 348
rect 194 328 270 331
rect 506 328 614 331
rect 634 328 718 331
rect 754 328 758 331
rect 770 328 1006 331
rect 1338 328 1462 331
rect 1594 328 1630 331
rect 1722 328 1782 331
rect 1786 328 1966 331
rect 2202 328 2206 331
rect 2258 328 2302 331
rect 154 318 294 321
rect 810 318 910 321
rect 978 318 1070 321
rect 1114 318 1158 321
rect 1630 321 1633 328
rect 1630 318 1678 321
rect 1698 318 1734 321
rect 1738 318 1774 321
rect 1834 318 1862 321
rect 1866 318 1998 321
rect 2022 321 2025 328
rect 2022 318 2270 321
rect 74 308 174 311
rect 290 308 766 311
rect 914 308 974 311
rect 978 308 1430 311
rect 1490 308 1630 311
rect 1634 308 1654 311
rect 1690 308 1726 311
rect 1762 308 1814 311
rect 1938 308 2022 311
rect 2050 308 2214 311
rect 880 303 882 307
rect 886 303 889 307
rect 894 303 896 307
rect 1912 303 1914 307
rect 1918 303 1921 307
rect 1926 303 1928 307
rect 618 298 838 301
rect 1002 298 1022 301
rect 1146 298 1169 301
rect 1178 298 1270 301
rect 1274 298 1422 301
rect 1562 298 1574 301
rect 1578 298 1606 301
rect 1970 298 2038 301
rect 2042 298 2110 301
rect 106 288 126 291
rect 322 288 398 291
rect 402 288 518 291
rect 706 288 790 291
rect 1018 288 1022 291
rect 1066 288 1142 291
rect 1166 291 1169 298
rect 1614 292 1617 298
rect 1166 288 1214 291
rect 1298 288 1438 291
rect 1442 288 1486 291
rect 1858 288 2097 291
rect 2094 282 2097 288
rect 242 278 310 281
rect 1082 278 1278 281
rect 1282 278 1350 281
rect 1402 278 1430 281
rect 1434 278 1622 281
rect 1634 278 1878 281
rect 42 268 46 271
rect 118 271 121 278
rect 214 271 217 278
rect 118 268 302 271
rect 306 268 334 271
rect 338 268 422 271
rect 458 268 510 271
rect 762 268 814 271
rect 958 271 961 278
rect 946 268 961 271
rect 1258 268 1510 271
rect 1530 268 1614 271
rect 1666 268 1670 271
rect 1674 268 1966 271
rect 2066 268 2150 271
rect 2162 268 2246 271
rect 2290 268 2294 271
rect 34 258 230 261
rect 234 258 262 261
rect 506 258 534 261
rect 730 258 902 261
rect 1046 261 1049 268
rect 1086 261 1089 268
rect 2006 262 2009 268
rect 1046 258 1089 261
rect 1458 258 1470 261
rect 1474 258 1974 261
rect 1978 258 1982 261
rect 2042 258 2046 261
rect 2050 258 2070 261
rect 2210 258 2254 261
rect 486 252 489 258
rect 2190 252 2193 258
rect 22 248 94 251
rect 274 248 286 251
rect 522 248 574 251
rect 818 248 846 251
rect 850 248 1102 251
rect 1122 248 1342 251
rect 1478 248 1550 251
rect 1610 248 1614 251
rect 1650 248 1910 251
rect 22 242 25 248
rect 1478 242 1481 248
rect 562 238 582 241
rect 586 238 670 241
rect 674 238 726 241
rect 786 238 830 241
rect 906 238 1214 241
rect 1218 238 1454 241
rect 1490 238 1590 241
rect 1682 238 1790 241
rect 1850 238 2038 241
rect 690 228 1310 231
rect 1426 228 1478 231
rect 1482 228 1934 231
rect 474 218 606 221
rect 818 218 998 221
rect 1186 218 1198 221
rect 1242 218 1342 221
rect 1406 221 1409 228
rect 1378 218 1494 221
rect 1498 218 1534 221
rect 1538 218 1606 221
rect 1610 218 1710 221
rect 2250 218 2286 221
rect 802 208 974 211
rect 1002 208 1174 211
rect 376 203 378 207
rect 382 203 385 207
rect 390 203 392 207
rect 1392 203 1394 207
rect 1398 203 1401 207
rect 1406 203 1408 207
rect 226 198 366 201
rect 1418 198 2014 201
rect 106 188 230 191
rect 242 188 366 191
rect 370 188 438 191
rect 546 188 550 191
rect 794 188 1022 191
rect 1094 191 1097 198
rect 1094 188 1150 191
rect 1154 188 1262 191
rect 1278 188 1486 191
rect 1866 188 1870 191
rect 1278 182 1281 188
rect 298 178 638 181
rect 642 178 774 181
rect 778 178 822 181
rect 826 178 902 181
rect 1090 178 1262 181
rect 1354 178 2174 181
rect 2178 178 2198 181
rect 114 168 494 171
rect 834 168 854 171
rect 858 168 1038 171
rect 1618 168 1686 171
rect 1730 168 1774 171
rect 122 158 142 161
rect 218 158 294 161
rect 354 158 398 161
rect 650 158 670 161
rect 682 158 718 161
rect 1110 161 1113 168
rect 1262 162 1265 168
rect 1042 158 1113 161
rect 1154 158 1158 161
rect 1170 158 1206 161
rect 1218 158 1230 161
rect 1362 158 1414 161
rect 1426 158 1702 161
rect 1706 158 1726 161
rect 1874 158 1894 161
rect 2258 158 2262 161
rect 2266 158 2286 161
rect 430 152 433 158
rect 298 148 350 151
rect 586 148 598 151
rect 602 148 830 151
rect 926 151 929 158
rect 858 148 929 151
rect 1106 148 1134 151
rect 1138 148 1382 151
rect 1386 148 1414 151
rect 1626 148 2118 151
rect 2122 148 2150 151
rect 126 141 129 148
rect 126 138 158 141
rect 466 138 558 141
rect 562 138 590 141
rect 686 138 774 141
rect 794 138 798 141
rect 818 138 942 141
rect 1058 138 1166 141
rect 1194 138 1286 141
rect 1354 138 1366 141
rect 1578 138 2078 141
rect 2082 138 2102 141
rect 2106 138 2174 141
rect 686 132 689 138
rect 106 128 214 131
rect 890 128 982 131
rect 1482 128 1886 131
rect 346 118 430 121
rect 946 118 1582 121
rect 1714 118 1742 121
rect 1822 118 1830 121
rect 1834 118 1854 121
rect 1898 118 1934 121
rect 2098 118 2134 121
rect 50 108 366 111
rect 482 108 686 111
rect 1258 108 1286 111
rect 1290 108 1326 111
rect 1498 108 1822 111
rect 1826 108 1838 111
rect 2066 108 2094 111
rect 366 101 369 108
rect 880 103 882 107
rect 886 103 889 107
rect 894 103 896 107
rect 1912 103 1914 107
rect 1918 103 1921 107
rect 1926 103 1928 107
rect 366 98 486 101
rect 498 98 614 101
rect 778 98 806 101
rect 1034 98 1102 101
rect 1106 98 1278 101
rect 1330 98 1350 101
rect 1474 98 1646 101
rect 1770 98 1830 101
rect 2026 98 2166 101
rect 2170 98 2214 101
rect 18 88 30 91
rect 130 88 238 91
rect 362 88 526 91
rect 562 88 590 91
rect 690 88 790 91
rect 858 88 918 91
rect 922 88 942 91
rect 962 88 1046 91
rect 1210 88 1318 91
rect 1322 88 1430 91
rect 1842 88 1857 91
rect 2010 88 2078 91
rect 1854 82 1857 88
rect 730 78 790 81
rect 818 78 862 81
rect 866 78 993 81
rect 1010 78 1062 81
rect 1066 78 1142 81
rect 1146 78 1238 81
rect 1242 78 1374 81
rect 1442 78 1534 81
rect 1818 78 1846 81
rect 50 68 62 71
rect 150 71 153 78
rect 150 68 190 71
rect 294 68 313 71
rect 354 68 374 71
rect 438 71 441 78
rect 394 68 441 71
rect 458 68 462 71
rect 694 71 697 78
rect 650 68 697 71
rect 786 68 870 71
rect 990 71 993 78
rect 990 68 1745 71
rect 2146 68 2270 71
rect 294 62 297 68
rect 310 62 313 68
rect 1742 62 1745 68
rect 10 58 46 61
rect 378 58 414 61
rect 418 58 854 61
rect 938 58 993 61
rect 1154 58 1294 61
rect 1314 58 1550 61
rect 1554 58 1566 61
rect 1618 58 1694 61
rect 1794 58 1798 61
rect 1802 58 1878 61
rect 1882 58 1902 61
rect 1906 58 1934 61
rect 1938 58 1974 61
rect 1986 58 2046 61
rect 2050 58 2174 61
rect 2178 58 2230 61
rect 2234 58 2254 61
rect 990 52 993 58
rect 50 48 110 51
rect 114 48 142 51
rect 466 48 478 51
rect 626 48 785 51
rect 794 48 830 51
rect 1394 48 1406 51
rect 1506 48 1558 51
rect 1586 48 1614 51
rect 1894 48 2022 51
rect 2034 48 2193 51
rect 782 42 785 48
rect 1894 42 1897 48
rect 2190 42 2193 48
rect 1082 8 1094 11
rect 1618 8 1622 11
rect 376 3 378 7
rect 382 3 385 7
rect 390 3 392 7
rect 1392 3 1394 7
rect 1398 3 1401 7
rect 1406 3 1408 7
<< m4contact >>
rect 882 2103 886 2107
rect 890 2103 893 2107
rect 893 2103 894 2107
rect 1914 2103 1918 2107
rect 1922 2103 1925 2107
rect 1925 2103 1926 2107
rect 278 2058 282 2062
rect 294 2058 298 2062
rect 310 2058 314 2062
rect 334 2058 338 2062
rect 2222 2068 2226 2072
rect 2230 2068 2234 2072
rect 2134 2058 2138 2062
rect 2246 2058 2250 2062
rect 6 2048 10 2052
rect 574 2048 578 2052
rect 910 2048 914 2052
rect 2014 2048 2018 2052
rect 2174 2048 2178 2052
rect 2286 2048 2290 2052
rect 758 2038 762 2042
rect 1278 2028 1282 2032
rect 2110 2018 2114 2022
rect 2254 2018 2258 2022
rect 378 2003 382 2007
rect 386 2003 389 2007
rect 389 2003 390 2007
rect 1394 2003 1398 2007
rect 1402 2003 1405 2007
rect 1405 2003 1406 2007
rect 1566 1998 1570 2002
rect 2014 1998 2018 2002
rect 1110 1978 1114 1982
rect 646 1968 650 1972
rect 1606 1968 1610 1972
rect 302 1958 306 1962
rect 502 1958 506 1962
rect 1638 1958 1642 1962
rect 518 1948 522 1952
rect 574 1948 578 1952
rect 590 1948 594 1952
rect 766 1948 770 1952
rect 902 1948 906 1952
rect 1222 1948 1226 1952
rect 710 1938 714 1942
rect 1158 1938 1162 1942
rect 1414 1938 1418 1942
rect 502 1928 506 1932
rect 1022 1928 1026 1932
rect 1854 1928 1858 1932
rect 190 1918 194 1922
rect 294 1918 298 1922
rect 2190 1918 2194 1922
rect 882 1903 886 1907
rect 890 1903 893 1907
rect 893 1903 894 1907
rect 1914 1903 1918 1907
rect 1922 1903 1925 1907
rect 1925 1903 1926 1907
rect 1062 1898 1066 1902
rect 1750 1878 1754 1882
rect 1790 1878 1794 1882
rect 1590 1868 1594 1872
rect 1606 1868 1610 1872
rect 118 1858 122 1862
rect 638 1858 642 1862
rect 878 1858 882 1862
rect 950 1858 954 1862
rect 1470 1858 1474 1862
rect 1854 1858 1858 1862
rect 1054 1848 1058 1852
rect 878 1838 882 1842
rect 958 1838 962 1842
rect 526 1828 530 1832
rect 558 1828 562 1832
rect 1518 1828 1522 1832
rect 2198 1828 2202 1832
rect 638 1818 642 1822
rect 1534 1818 1538 1822
rect 1550 1818 1554 1822
rect 378 1803 382 1807
rect 386 1803 389 1807
rect 389 1803 390 1807
rect 1394 1803 1398 1807
rect 1402 1803 1405 1807
rect 1405 1803 1406 1807
rect 342 1798 346 1802
rect 982 1798 986 1802
rect 1606 1788 1610 1792
rect 670 1778 674 1782
rect 854 1778 858 1782
rect 1110 1778 1114 1782
rect 118 1768 122 1772
rect 2094 1768 2098 1772
rect 342 1758 346 1762
rect 1798 1758 1802 1762
rect 2030 1758 2034 1762
rect 2150 1758 2154 1762
rect 2174 1758 2178 1762
rect 598 1748 602 1752
rect 1062 1748 1066 1752
rect 1230 1748 1234 1752
rect 2014 1748 2018 1752
rect 358 1738 362 1742
rect 518 1738 522 1742
rect 662 1738 666 1742
rect 710 1738 714 1742
rect 982 1738 986 1742
rect 1294 1738 1298 1742
rect 1414 1738 1418 1742
rect 1590 1738 1594 1742
rect 246 1728 250 1732
rect 278 1728 282 1732
rect 862 1728 866 1732
rect 1030 1728 1034 1732
rect 942 1718 946 1722
rect 1046 1718 1050 1722
rect 6 1708 10 1712
rect 462 1708 466 1712
rect 1158 1708 1162 1712
rect 1678 1708 1682 1712
rect 1686 1708 1690 1712
rect 882 1703 886 1707
rect 890 1703 893 1707
rect 893 1703 894 1707
rect 1914 1703 1918 1707
rect 1922 1703 1925 1707
rect 1925 1703 1926 1707
rect 1222 1698 1226 1702
rect 1878 1698 1882 1702
rect 1526 1688 1530 1692
rect 518 1668 522 1672
rect 1558 1668 1562 1672
rect 2198 1668 2202 1672
rect 278 1658 282 1662
rect 358 1658 362 1662
rect 670 1658 674 1662
rect 982 1658 986 1662
rect 1054 1658 1058 1662
rect 1214 1658 1218 1662
rect 110 1648 114 1652
rect 718 1648 722 1652
rect 1006 1648 1010 1652
rect 1254 1648 1258 1652
rect 1366 1648 1370 1652
rect 1574 1648 1578 1652
rect 1694 1648 1698 1652
rect 1782 1648 1786 1652
rect 1870 1648 1874 1652
rect 534 1638 538 1642
rect 590 1638 594 1642
rect 990 1638 994 1642
rect 1062 1628 1066 1632
rect 990 1618 994 1622
rect 1022 1618 1026 1622
rect 1238 1618 1242 1622
rect 1534 1618 1538 1622
rect 2022 1618 2026 1622
rect 378 1603 382 1607
rect 386 1603 389 1607
rect 389 1603 390 1607
rect 1394 1603 1398 1607
rect 1402 1603 1405 1607
rect 1405 1603 1406 1607
rect 1006 1588 1010 1592
rect 1142 1588 1146 1592
rect 1238 1578 1242 1582
rect 1838 1578 1842 1582
rect 2070 1578 2074 1582
rect 1438 1568 1442 1572
rect 558 1558 562 1562
rect 670 1558 674 1562
rect 1542 1558 1546 1562
rect 1798 1558 1802 1562
rect 2102 1558 2106 1562
rect 102 1548 106 1552
rect 670 1548 674 1552
rect 846 1548 850 1552
rect 1254 1548 1258 1552
rect 1278 1548 1282 1552
rect 1454 1548 1458 1552
rect 1470 1548 1474 1552
rect 1966 1548 1970 1552
rect 2134 1548 2138 1552
rect 2206 1548 2210 1552
rect 566 1538 570 1542
rect 1806 1538 1810 1542
rect 1990 1538 1994 1542
rect 2078 1538 2082 1542
rect 2142 1538 2146 1542
rect 438 1528 442 1532
rect 1046 1528 1050 1532
rect 1550 1528 1554 1532
rect 1758 1528 1762 1532
rect 1806 1528 1810 1532
rect 118 1518 122 1522
rect 1142 1518 1146 1522
rect 1798 1518 1802 1522
rect 2150 1518 2154 1522
rect 454 1508 458 1512
rect 742 1508 746 1512
rect 910 1508 914 1512
rect 1230 1508 1234 1512
rect 882 1503 886 1507
rect 890 1503 893 1507
rect 893 1503 894 1507
rect 1914 1503 1918 1507
rect 1922 1503 1925 1507
rect 1925 1503 1926 1507
rect 870 1498 874 1502
rect 958 1498 962 1502
rect 1982 1498 1986 1502
rect 2166 1498 2170 1502
rect 1134 1488 1138 1492
rect 1158 1488 1162 1492
rect 1470 1488 1474 1492
rect 1478 1488 1482 1492
rect 1278 1478 1282 1482
rect 1302 1478 1306 1482
rect 2070 1478 2074 1482
rect 302 1468 306 1472
rect 478 1468 482 1472
rect 702 1468 706 1472
rect 798 1468 802 1472
rect 1054 1468 1058 1472
rect 1526 1468 1530 1472
rect 1966 1468 1970 1472
rect 214 1458 218 1462
rect 1126 1458 1130 1462
rect 1190 1458 1194 1462
rect 1246 1458 1250 1462
rect 1294 1458 1298 1462
rect 1374 1458 1378 1462
rect 1430 1458 1434 1462
rect 1462 1458 1466 1462
rect 1494 1458 1498 1462
rect 2110 1458 2114 1462
rect 102 1448 106 1452
rect 454 1448 458 1452
rect 574 1448 578 1452
rect 750 1448 754 1452
rect 854 1448 858 1452
rect 1350 1448 1354 1452
rect 1502 1448 1506 1452
rect 1638 1448 1642 1452
rect 702 1438 706 1442
rect 710 1438 714 1442
rect 790 1438 794 1442
rect 1022 1438 1026 1442
rect 1214 1438 1218 1442
rect 1358 1438 1362 1442
rect 1478 1438 1482 1442
rect 2206 1438 2210 1442
rect 2246 1438 2250 1442
rect 174 1428 178 1432
rect 278 1428 282 1432
rect 1030 1428 1034 1432
rect 1694 1428 1698 1432
rect 1798 1428 1802 1432
rect 766 1418 770 1422
rect 1678 1418 1682 1422
rect 1558 1408 1562 1412
rect 378 1403 382 1407
rect 386 1403 389 1407
rect 389 1403 390 1407
rect 1394 1403 1398 1407
rect 1402 1403 1405 1407
rect 1405 1403 1406 1407
rect 518 1398 522 1402
rect 1526 1398 1530 1402
rect 766 1388 770 1392
rect 1030 1388 1034 1392
rect 1614 1388 1618 1392
rect 1118 1378 1122 1382
rect 1542 1378 1546 1382
rect 2110 1378 2114 1382
rect 622 1368 626 1372
rect 1054 1368 1058 1372
rect 1270 1368 1274 1372
rect 1454 1368 1458 1372
rect 1542 1368 1546 1372
rect 630 1358 634 1362
rect 1174 1358 1178 1362
rect 1350 1358 1354 1362
rect 1414 1358 1418 1362
rect 1454 1358 1458 1362
rect 1566 1358 1570 1362
rect 1862 1358 1866 1362
rect 1974 1358 1978 1362
rect 1982 1358 1986 1362
rect 230 1348 234 1352
rect 246 1348 250 1352
rect 798 1348 802 1352
rect 926 1348 930 1352
rect 1014 1348 1018 1352
rect 1366 1348 1370 1352
rect 1382 1348 1386 1352
rect 1510 1348 1514 1352
rect 1782 1348 1786 1352
rect 2070 1348 2074 1352
rect 358 1338 362 1342
rect 1374 1338 1378 1342
rect 1414 1338 1418 1342
rect 1438 1338 1442 1342
rect 1462 1338 1466 1342
rect 1774 1338 1778 1342
rect 1838 1338 1842 1342
rect 2070 1338 2074 1342
rect 2182 1338 2186 1342
rect 1102 1328 1106 1332
rect 1446 1328 1450 1332
rect 1574 1328 1578 1332
rect 1958 1328 1962 1332
rect 190 1318 194 1322
rect 1182 1318 1186 1322
rect 1566 1318 1570 1322
rect 1374 1308 1378 1312
rect 1902 1308 1906 1312
rect 1966 1308 1970 1312
rect 1974 1308 1978 1312
rect 882 1303 886 1307
rect 890 1303 893 1307
rect 893 1303 894 1307
rect 150 1298 154 1302
rect 1914 1303 1918 1307
rect 1922 1303 1925 1307
rect 1925 1303 1926 1307
rect 2078 1298 2082 1302
rect 1902 1288 1906 1292
rect 486 1278 490 1282
rect 558 1278 562 1282
rect 534 1268 538 1272
rect 542 1268 546 1272
rect 646 1268 650 1272
rect 1142 1268 1146 1272
rect 1430 1268 1434 1272
rect 2102 1268 2106 1272
rect 2182 1268 2186 1272
rect 134 1258 138 1262
rect 606 1258 610 1262
rect 926 1258 930 1262
rect 1014 1258 1018 1262
rect 1198 1258 1202 1262
rect 1806 1258 1810 1262
rect 1886 1258 1890 1262
rect 1910 1258 1914 1262
rect 118 1248 122 1252
rect 1030 1248 1034 1252
rect 1110 1248 1114 1252
rect 1166 1248 1170 1252
rect 1350 1248 1354 1252
rect 1382 1248 1386 1252
rect 1462 1248 1466 1252
rect 1694 1248 1698 1252
rect 1702 1248 1706 1252
rect 1070 1238 1074 1242
rect 1078 1238 1082 1242
rect 1662 1238 1666 1242
rect 2254 1238 2258 1242
rect 670 1228 674 1232
rect 1646 1228 1650 1232
rect 1358 1218 1362 1222
rect 2022 1218 2026 1222
rect 1054 1208 1058 1212
rect 1198 1208 1202 1212
rect 1422 1208 1426 1212
rect 378 1203 382 1207
rect 386 1203 389 1207
rect 389 1203 390 1207
rect 1086 1198 1090 1202
rect 1394 1203 1398 1207
rect 1402 1203 1405 1207
rect 1405 1203 1406 1207
rect 1894 1198 1898 1202
rect 142 1188 146 1192
rect 990 1178 994 1182
rect 1110 1178 1114 1182
rect 1542 1178 1546 1182
rect 502 1168 506 1172
rect 1014 1168 1018 1172
rect 1094 1168 1098 1172
rect 1126 1168 1130 1172
rect 1254 1158 1258 1162
rect 1518 1158 1522 1162
rect 1558 1158 1562 1162
rect 1606 1158 1610 1162
rect 1750 1158 1754 1162
rect 1758 1158 1762 1162
rect 1830 1158 1834 1162
rect 2110 1158 2114 1162
rect 278 1148 282 1152
rect 654 1148 658 1152
rect 694 1148 698 1152
rect 1022 1148 1026 1152
rect 1038 1148 1042 1152
rect 1046 1148 1050 1152
rect 1054 1148 1058 1152
rect 1174 1148 1178 1152
rect 1278 1148 1282 1152
rect 1518 1148 1522 1152
rect 1638 1148 1642 1152
rect 1662 1148 1666 1152
rect 1846 1148 1850 1152
rect 2166 1148 2170 1152
rect 302 1138 306 1142
rect 350 1138 354 1142
rect 150 1128 154 1132
rect 262 1128 266 1132
rect 782 1138 786 1142
rect 790 1138 794 1142
rect 1414 1138 1418 1142
rect 1502 1138 1506 1142
rect 2046 1138 2050 1142
rect 2190 1138 2194 1142
rect 646 1128 650 1132
rect 774 1128 778 1132
rect 1166 1128 1170 1132
rect 1422 1128 1426 1132
rect 1486 1128 1490 1132
rect 1766 1128 1770 1132
rect 1142 1118 1146 1122
rect 430 1108 434 1112
rect 734 1108 738 1112
rect 1790 1108 1794 1112
rect 1806 1108 1810 1112
rect 2278 1108 2282 1112
rect 882 1103 886 1107
rect 890 1103 893 1107
rect 893 1103 894 1107
rect 1914 1103 1918 1107
rect 1922 1103 1925 1107
rect 1925 1103 1926 1107
rect 1038 1098 1042 1102
rect 1190 1098 1194 1102
rect 1350 1098 1354 1102
rect 2222 1098 2226 1102
rect 1142 1088 1146 1092
rect 1286 1088 1290 1092
rect 2078 1088 2082 1092
rect 2286 1078 2290 1082
rect 254 1068 258 1072
rect 1214 1068 1218 1072
rect 1494 1068 1498 1072
rect 1582 1068 1586 1072
rect 1598 1068 1602 1072
rect 1662 1068 1666 1072
rect 1798 1068 1802 1072
rect 1806 1068 1810 1072
rect 2070 1068 2074 1072
rect 366 1058 370 1062
rect 942 1058 946 1062
rect 1566 1058 1570 1062
rect 1574 1058 1578 1062
rect 1886 1058 1890 1062
rect 198 1048 202 1052
rect 230 1048 234 1052
rect 1014 1048 1018 1052
rect 1358 1048 1362 1052
rect 1462 1048 1466 1052
rect 1574 1048 1578 1052
rect 1830 1048 1834 1052
rect 2110 1048 2114 1052
rect 1598 1038 1602 1042
rect 1862 1038 1866 1042
rect 118 1028 122 1032
rect 438 1028 442 1032
rect 1446 1028 1450 1032
rect 1630 1028 1634 1032
rect 214 1018 218 1022
rect 998 1018 1002 1022
rect 1214 1018 1218 1022
rect 1606 1018 1610 1022
rect 174 1008 178 1012
rect 638 1008 642 1012
rect 950 1008 954 1012
rect 1006 1008 1010 1012
rect 1206 1008 1210 1012
rect 1510 1008 1514 1012
rect 2070 1008 2074 1012
rect 2262 1008 2266 1012
rect 378 1003 382 1007
rect 386 1003 389 1007
rect 389 1003 390 1007
rect 1394 1003 1398 1007
rect 1402 1003 1405 1007
rect 1405 1003 1406 1007
rect 942 988 946 992
rect 950 988 954 992
rect 1270 988 1274 992
rect 1486 988 1490 992
rect 1854 988 1858 992
rect 1078 978 1082 982
rect 1422 978 1426 982
rect 1486 978 1490 982
rect 510 968 514 972
rect 934 968 938 972
rect 950 968 954 972
rect 1478 968 1482 972
rect 142 958 146 962
rect 310 958 314 962
rect 630 958 634 962
rect 1046 958 1050 962
rect 1062 958 1066 962
rect 1446 958 1450 962
rect 2022 958 2026 962
rect 142 948 146 952
rect 830 948 834 952
rect 982 948 986 952
rect 1246 948 1250 952
rect 1382 948 1386 952
rect 1526 948 1530 952
rect 1718 948 1722 952
rect 1854 948 1858 952
rect 1878 948 1882 952
rect 1974 948 1978 952
rect 2062 948 2066 952
rect 486 938 490 942
rect 542 938 546 942
rect 1134 938 1138 942
rect 1542 938 1546 942
rect 1998 938 2002 942
rect 150 928 154 932
rect 622 928 626 932
rect 1254 928 1258 932
rect 1294 928 1298 932
rect 2046 928 2050 932
rect 1366 918 1370 922
rect 118 908 122 912
rect 302 908 306 912
rect 758 908 762 912
rect 1006 908 1010 912
rect 1550 908 1554 912
rect 882 903 886 907
rect 890 903 893 907
rect 893 903 894 907
rect 1914 903 1918 907
rect 1922 903 1925 907
rect 1925 903 1926 907
rect 422 898 426 902
rect 1542 898 1546 902
rect 1846 898 1850 902
rect 1902 898 1906 902
rect 2278 898 2282 902
rect 438 888 442 892
rect 830 888 834 892
rect 894 888 898 892
rect 1182 888 1186 892
rect 1526 888 1530 892
rect 1766 888 1770 892
rect 1830 888 1834 892
rect 518 878 522 882
rect 566 878 570 882
rect 782 878 786 882
rect 942 878 946 882
rect 982 878 986 882
rect 1166 878 1170 882
rect 1350 878 1354 882
rect 1542 878 1546 882
rect 262 868 266 872
rect 654 868 658 872
rect 894 868 898 872
rect 1566 868 1570 872
rect 1598 868 1602 872
rect 1742 868 1746 872
rect 174 858 178 862
rect 734 858 738 862
rect 902 858 906 862
rect 1046 858 1050 862
rect 1102 858 1106 862
rect 1110 858 1114 862
rect 1782 858 1786 862
rect 2078 858 2082 862
rect 414 848 418 852
rect 950 848 954 852
rect 982 848 986 852
rect 1526 848 1530 852
rect 1638 848 1642 852
rect 1822 848 1826 852
rect 1862 848 1866 852
rect 1958 848 1962 852
rect 2190 848 2194 852
rect 2230 848 2234 852
rect 2302 848 2306 852
rect 1534 838 1538 842
rect 1758 838 1762 842
rect 1806 838 1810 842
rect 446 828 450 832
rect 462 828 466 832
rect 1078 828 1082 832
rect 1030 808 1034 812
rect 378 803 382 807
rect 386 803 389 807
rect 389 803 390 807
rect 1394 803 1398 807
rect 1402 803 1405 807
rect 1405 803 1406 807
rect 1798 798 1802 802
rect 502 788 506 792
rect 726 778 730 782
rect 1070 778 1074 782
rect 142 768 146 772
rect 1374 768 1378 772
rect 1486 768 1490 772
rect 1766 768 1770 772
rect 1790 768 1794 772
rect 1878 768 1882 772
rect 1902 768 1906 772
rect 2302 768 2306 772
rect 430 758 434 762
rect 510 758 514 762
rect 854 758 858 762
rect 1214 758 1218 762
rect 2014 758 2018 762
rect 422 748 426 752
rect 438 748 442 752
rect 990 748 994 752
rect 1142 748 1146 752
rect 1262 748 1266 752
rect 1430 748 1434 752
rect 1734 748 1738 752
rect 1862 748 1866 752
rect 1878 748 1882 752
rect 2030 748 2034 752
rect 2046 748 2050 752
rect 294 738 298 742
rect 494 738 498 742
rect 638 738 642 742
rect 654 738 658 742
rect 790 738 794 742
rect 1094 738 1098 742
rect 1118 738 1122 742
rect 1198 738 1202 742
rect 1222 738 1226 742
rect 1990 738 1994 742
rect 2198 738 2202 742
rect 654 728 658 732
rect 1774 728 1778 732
rect 1838 728 1842 732
rect 2190 728 2194 732
rect 102 718 106 722
rect 166 718 170 722
rect 414 718 418 722
rect 1022 718 1026 722
rect 1854 718 1858 722
rect 2030 718 2034 722
rect 350 708 354 712
rect 1062 708 1066 712
rect 1166 708 1170 712
rect 882 703 886 707
rect 890 703 893 707
rect 893 703 894 707
rect 1914 703 1918 707
rect 1922 703 1925 707
rect 1925 703 1926 707
rect 454 698 458 702
rect 958 698 962 702
rect 1302 698 1306 702
rect 1054 688 1058 692
rect 1486 688 1490 692
rect 1574 688 1578 692
rect 1582 688 1586 692
rect 1678 688 1682 692
rect 1710 688 1714 692
rect 1718 688 1722 692
rect 358 678 362 682
rect 590 678 594 682
rect 758 678 762 682
rect 998 678 1002 682
rect 1022 678 1026 682
rect 1126 678 1130 682
rect 1454 678 1458 682
rect 958 668 962 672
rect 1006 668 1010 672
rect 1158 668 1162 672
rect 1542 668 1546 672
rect 1558 668 1562 672
rect 1742 668 1746 672
rect 1758 668 1762 672
rect 1838 668 1842 672
rect 1134 658 1138 662
rect 1422 658 1426 662
rect 1454 658 1458 662
rect 1894 658 1898 662
rect 2246 658 2250 662
rect 430 648 434 652
rect 686 648 690 652
rect 766 648 770 652
rect 1030 648 1034 652
rect 1046 648 1050 652
rect 1174 648 1178 652
rect 1358 648 1362 652
rect 1726 648 1730 652
rect 1862 648 1866 652
rect 2102 648 2106 652
rect 1214 638 1218 642
rect 1518 638 1522 642
rect 1942 638 1946 642
rect 1446 628 1450 632
rect 1774 628 1778 632
rect 2110 628 2114 632
rect 1430 608 1434 612
rect 378 603 382 607
rect 386 603 389 607
rect 389 603 390 607
rect 174 598 178 602
rect 614 598 618 602
rect 1394 603 1398 607
rect 1402 603 1405 607
rect 1405 603 1406 607
rect 1782 588 1786 592
rect 190 578 194 582
rect 310 568 314 572
rect 422 568 426 572
rect 750 568 754 572
rect 1190 568 1194 572
rect 1206 568 1210 572
rect 1230 568 1234 572
rect 1286 568 1290 572
rect 1158 558 1162 562
rect 1838 558 1842 562
rect 2070 558 2074 562
rect 1118 548 1122 552
rect 1414 548 1418 552
rect 1478 548 1482 552
rect 1734 548 1738 552
rect 2014 548 2018 552
rect 454 538 458 542
rect 574 538 578 542
rect 870 538 874 542
rect 1222 538 1226 542
rect 1254 538 1258 542
rect 1462 538 1466 542
rect 1494 538 1498 542
rect 2286 538 2290 542
rect 910 528 914 532
rect 1246 528 1250 532
rect 1502 528 1506 532
rect 990 518 994 522
rect 1094 518 1098 522
rect 1462 518 1466 522
rect 174 508 178 512
rect 1902 508 1906 512
rect 882 503 886 507
rect 890 503 893 507
rect 893 503 894 507
rect 1914 503 1918 507
rect 1922 503 1925 507
rect 1925 503 1926 507
rect 446 498 450 502
rect 1030 498 1034 502
rect 2190 488 2194 492
rect 1422 478 1426 482
rect 2014 478 2018 482
rect 1374 468 1378 472
rect 2006 468 2010 472
rect 278 458 282 462
rect 326 458 330 462
rect 1486 458 1490 462
rect 2078 458 2082 462
rect 2030 448 2034 452
rect 1534 438 1538 442
rect 1854 438 1858 442
rect 166 428 170 432
rect 1126 428 1130 432
rect 590 418 594 422
rect 982 418 986 422
rect 1102 418 1106 422
rect 1502 418 1506 422
rect 870 408 874 412
rect 1958 408 1962 412
rect 378 403 382 407
rect 386 403 389 407
rect 389 403 390 407
rect 1394 403 1398 407
rect 1402 403 1405 407
rect 1405 403 1406 407
rect 1110 388 1114 392
rect 1638 378 1642 382
rect 1646 378 1650 382
rect 614 368 618 372
rect 734 368 738 372
rect 1038 368 1042 372
rect 1102 368 1106 372
rect 1614 368 1618 372
rect 1622 368 1626 372
rect 1670 368 1674 372
rect 902 358 906 362
rect 1046 358 1050 362
rect 1174 358 1178 362
rect 1302 358 1306 362
rect 2030 358 2034 362
rect 2262 358 2266 362
rect 326 348 330 352
rect 494 348 498 352
rect 510 348 514 352
rect 1030 348 1034 352
rect 302 338 306 342
rect 566 338 570 342
rect 1046 338 1050 342
rect 1510 338 1514 342
rect 1902 338 1906 342
rect 758 328 762 332
rect 766 328 770 332
rect 2206 328 2210 332
rect 766 308 770 312
rect 910 308 914 312
rect 1486 308 1490 312
rect 1934 308 1938 312
rect 882 303 886 307
rect 890 303 893 307
rect 893 303 894 307
rect 1914 303 1918 307
rect 1922 303 1925 307
rect 1925 303 1926 307
rect 1022 298 1026 302
rect 1174 298 1178 302
rect 1422 298 1426 302
rect 1022 288 1026 292
rect 1614 288 1618 292
rect 1078 278 1082 282
rect 1630 278 1634 282
rect 942 268 946 272
rect 1510 268 1514 272
rect 1670 268 1674 272
rect 2286 268 2290 272
rect 230 258 234 262
rect 2006 258 2010 262
rect 2046 258 2050 262
rect 2254 258 2258 262
rect 486 248 490 252
rect 1614 248 1618 252
rect 2190 248 2194 252
rect 726 238 730 242
rect 902 238 906 242
rect 1846 238 1850 242
rect 686 228 690 232
rect 1422 228 1426 232
rect 1934 228 1938 232
rect 2246 218 2250 222
rect 378 203 382 207
rect 386 203 389 207
rect 389 203 390 207
rect 1394 203 1398 207
rect 1402 203 1405 207
rect 1405 203 1406 207
rect 1414 198 1418 202
rect 238 188 242 192
rect 366 188 370 192
rect 790 188 794 192
rect 1870 188 1874 192
rect 1262 178 1266 182
rect 2198 178 2202 182
rect 110 168 114 172
rect 494 168 498 172
rect 1262 168 1266 172
rect 1726 168 1730 172
rect 1150 158 1154 162
rect 1414 158 1418 162
rect 2262 158 2266 162
rect 430 148 434 152
rect 790 138 794 142
rect 942 138 946 142
rect 2174 138 2178 142
rect 1478 128 1482 132
rect 686 108 690 112
rect 1494 108 1498 112
rect 882 103 886 107
rect 890 103 893 107
rect 893 103 894 107
rect 1914 103 1918 107
rect 1922 103 1925 107
rect 1925 103 1926 107
rect 486 98 490 102
rect 238 88 242 92
rect 854 88 858 92
rect 2006 88 2010 92
rect 790 78 794 82
rect 374 68 378 72
rect 462 68 466 72
rect 854 58 858 62
rect 790 48 794 52
rect 1622 8 1626 12
rect 378 3 382 7
rect 386 3 389 7
rect 389 3 390 7
rect 1394 3 1398 7
rect 1402 3 1405 7
rect 1405 3 1406 7
<< metal4 >>
rect 880 2103 882 2107
rect 886 2103 889 2107
rect 894 2103 896 2107
rect 1912 2103 1914 2107
rect 1918 2103 1921 2107
rect 1926 2103 1928 2107
rect 282 2058 286 2061
rect 302 2058 310 2061
rect 330 2058 334 2061
rect 6 1712 9 2048
rect 294 1922 297 2058
rect 302 2052 305 2058
rect 578 2048 582 2051
rect 902 2048 910 2051
rect 2018 2048 2025 2051
rect 302 1962 305 2048
rect 758 2042 761 2048
rect 376 2003 378 2007
rect 382 2003 385 2007
rect 390 2003 392 2007
rect 638 1968 646 1971
rect 502 1932 505 1958
rect 186 1918 190 1921
rect 118 1772 121 1858
rect 376 1803 378 1807
rect 382 1803 385 1807
rect 390 1803 392 1807
rect 102 1452 105 1548
rect 102 722 105 1448
rect 110 172 113 1648
rect 118 1522 121 1768
rect 342 1762 345 1798
rect 518 1742 521 1948
rect 562 1828 569 1831
rect 118 1252 121 1518
rect 138 1258 142 1261
rect 118 912 121 1028
rect 142 962 145 1188
rect 150 1132 153 1298
rect 142 952 145 958
rect 142 772 145 948
rect 150 932 153 1128
rect 174 1012 177 1428
rect 166 432 169 718
rect 174 602 177 858
rect 174 512 177 598
rect 190 582 193 1318
rect 198 1052 201 1068
rect 214 1022 217 1458
rect 246 1352 249 1728
rect 278 1662 281 1728
rect 358 1662 361 1738
rect 306 1468 310 1471
rect 230 1052 233 1348
rect 278 1152 281 1428
rect 302 1142 305 1468
rect 358 1342 361 1658
rect 376 1603 378 1607
rect 382 1603 385 1607
rect 390 1603 392 1607
rect 376 1403 378 1407
rect 382 1403 385 1407
rect 390 1403 392 1407
rect 250 1068 254 1071
rect 230 262 233 1048
rect 262 872 265 1128
rect 302 912 305 1138
rect 302 741 305 908
rect 298 738 305 741
rect 282 458 286 461
rect 302 342 305 738
rect 310 572 313 958
rect 350 712 353 1138
rect 358 682 361 1338
rect 376 1203 378 1207
rect 382 1203 385 1207
rect 390 1203 392 1207
rect 330 458 334 461
rect 330 348 334 351
rect 366 192 369 1058
rect 376 1003 378 1007
rect 382 1003 385 1007
rect 390 1003 392 1007
rect 376 803 378 807
rect 382 803 385 807
rect 390 803 392 807
rect 414 722 417 848
rect 422 752 425 898
rect 430 762 433 1108
rect 438 1032 441 1528
rect 454 1462 457 1508
rect 454 1452 457 1458
rect 438 752 441 888
rect 462 832 465 1708
rect 526 1671 529 1828
rect 522 1668 529 1671
rect 478 1281 481 1468
rect 478 1278 486 1281
rect 478 1152 481 1278
rect 422 648 430 651
rect 376 603 378 607
rect 382 603 385 607
rect 390 603 392 607
rect 422 572 425 648
rect 446 502 449 828
rect 486 741 489 938
rect 502 792 505 1168
rect 518 971 521 1398
rect 534 1272 537 1638
rect 558 1282 561 1558
rect 566 1542 569 1828
rect 574 1452 577 1948
rect 590 1922 593 1948
rect 590 1642 593 1918
rect 638 1862 641 1968
rect 902 1952 905 2048
rect 714 1938 721 1941
rect 598 1752 601 1838
rect 514 968 521 971
rect 542 942 545 1268
rect 598 1261 601 1748
rect 622 1362 625 1368
rect 598 1258 606 1261
rect 630 962 633 1358
rect 638 1271 641 1818
rect 662 1778 670 1781
rect 662 1742 665 1778
rect 674 1658 678 1661
rect 670 1552 673 1558
rect 638 1268 646 1271
rect 670 1262 673 1548
rect 702 1442 705 1468
rect 710 1442 713 1738
rect 718 1652 721 1938
rect 734 1508 742 1511
rect 670 1232 673 1258
rect 698 1148 702 1151
rect 638 1128 646 1131
rect 638 1012 641 1128
rect 626 928 630 931
rect 522 878 526 881
rect 486 738 494 741
rect 454 542 457 698
rect 376 403 378 407
rect 382 403 385 407
rect 390 403 392 407
rect 494 352 497 358
rect 510 352 513 758
rect 566 541 569 878
rect 654 872 657 1148
rect 734 1112 737 1508
rect 642 738 646 741
rect 654 732 657 738
rect 566 538 574 541
rect 590 422 593 678
rect 614 372 617 598
rect 376 203 378 207
rect 382 203 385 207
rect 390 203 392 207
rect 238 92 241 188
rect 434 148 438 151
rect 486 102 489 248
rect 494 172 497 348
rect 570 338 574 341
rect 686 232 689 648
rect 726 242 729 778
rect 734 372 737 858
rect 750 572 753 1448
rect 766 1422 769 1948
rect 880 1903 882 1907
rect 886 1903 889 1907
rect 894 1903 896 1907
rect 942 1858 950 1861
rect 878 1842 881 1858
rect 794 1468 798 1471
rect 758 892 761 908
rect 758 672 761 678
rect 766 652 769 1388
rect 790 1142 793 1438
rect 802 1348 806 1351
rect 846 1152 849 1548
rect 854 1452 857 1778
rect 862 1162 865 1728
rect 942 1722 945 1858
rect 954 1838 958 1841
rect 982 1742 985 1798
rect 880 1703 882 1707
rect 886 1703 889 1707
rect 894 1703 896 1707
rect 982 1662 985 1738
rect 1010 1648 1014 1651
rect 990 1622 993 1638
rect 1022 1622 1025 1928
rect 880 1503 882 1507
rect 886 1503 889 1507
rect 894 1503 896 1507
rect 870 1482 873 1498
rect 880 1303 882 1307
rect 886 1303 889 1307
rect 894 1303 896 1307
rect 782 1132 785 1138
rect 774 952 777 1128
rect 782 882 785 1128
rect 880 1103 882 1107
rect 886 1103 889 1107
rect 894 1103 896 1107
rect 830 892 833 948
rect 880 903 882 907
rect 886 903 889 907
rect 894 903 896 907
rect 894 872 897 888
rect 738 368 742 371
rect 750 332 753 568
rect 754 328 758 331
rect 766 312 769 328
rect 686 112 689 228
rect 790 192 793 738
rect 790 142 793 188
rect 854 92 857 758
rect 880 703 882 707
rect 886 703 889 707
rect 894 703 896 707
rect 870 412 873 538
rect 880 503 882 507
rect 886 503 889 507
rect 894 503 896 507
rect 902 362 905 858
rect 910 532 913 1508
rect 922 1348 926 1351
rect 926 971 929 1258
rect 942 992 945 1058
rect 950 992 953 1008
rect 926 968 934 971
rect 880 303 882 307
rect 886 303 889 307
rect 894 303 896 307
rect 902 242 905 358
rect 910 312 913 348
rect 942 272 945 878
rect 950 852 953 968
rect 958 702 961 1498
rect 990 951 993 1178
rect 998 1022 1001 1038
rect 1006 1012 1009 1588
rect 1022 1442 1025 1448
rect 1030 1432 1033 1728
rect 1046 1532 1049 1718
rect 1054 1662 1057 1848
rect 1062 1752 1065 1898
rect 1110 1782 1113 1978
rect 1158 1712 1161 1938
rect 1222 1702 1225 1948
rect 1014 1262 1017 1348
rect 1030 1252 1033 1388
rect 1054 1372 1057 1468
rect 1034 1248 1038 1251
rect 1054 1212 1057 1368
rect 1014 1052 1017 1168
rect 1054 1152 1057 1208
rect 1034 1148 1038 1151
rect 1022 1132 1025 1148
rect 1014 1032 1017 1048
rect 986 948 993 951
rect 982 852 985 878
rect 958 672 961 698
rect 990 522 993 748
rect 998 682 1001 688
rect 1006 672 1009 908
rect 1022 722 1025 1128
rect 1022 682 1025 708
rect 986 418 990 421
rect 1022 302 1025 678
rect 1030 652 1033 808
rect 1030 352 1033 498
rect 1038 372 1041 1098
rect 1046 962 1049 1148
rect 1046 862 1049 958
rect 1054 692 1057 978
rect 1062 962 1065 1628
rect 1142 1522 1145 1588
rect 1102 1332 1105 1348
rect 1110 1252 1113 1258
rect 1070 782 1073 1238
rect 1078 982 1081 1238
rect 1086 982 1089 1198
rect 1098 1168 1102 1171
rect 1110 862 1113 1178
rect 1118 1171 1121 1378
rect 1126 1231 1129 1458
rect 1134 1242 1137 1488
rect 1142 1272 1145 1278
rect 1126 1228 1137 1231
rect 1118 1168 1126 1171
rect 1134 942 1137 1228
rect 1142 1092 1145 1118
rect 1062 712 1065 728
rect 1046 362 1049 648
rect 1042 338 1046 341
rect 1018 288 1022 291
rect 1078 282 1081 828
rect 1094 522 1097 738
rect 1102 422 1105 858
rect 1102 372 1105 418
rect 1110 392 1113 858
rect 1118 552 1121 738
rect 1126 682 1129 688
rect 1134 662 1137 938
rect 1146 748 1150 751
rect 1158 672 1161 1488
rect 1166 1358 1174 1361
rect 1166 1252 1169 1358
rect 1182 1322 1185 1538
rect 1166 1132 1169 1138
rect 1166 882 1169 1128
rect 1174 891 1177 1148
rect 1190 1102 1193 1458
rect 1214 1442 1217 1658
rect 1202 1258 1206 1261
rect 1198 1152 1201 1208
rect 1214 1072 1217 1438
rect 1214 1062 1217 1068
rect 1174 888 1182 891
rect 1166 712 1169 878
rect 1174 652 1177 888
rect 1194 738 1198 741
rect 1206 572 1209 1008
rect 1214 762 1217 1018
rect 1222 742 1225 1698
rect 1230 1512 1233 1748
rect 1258 1648 1262 1651
rect 1238 1582 1241 1618
rect 1238 1461 1241 1578
rect 1278 1552 1281 2028
rect 1392 2003 1394 2007
rect 1398 2003 1401 2007
rect 1406 2003 1408 2007
rect 1570 1998 1577 2001
rect 1392 1803 1394 1807
rect 1398 1803 1401 1807
rect 1406 1803 1408 1807
rect 1414 1742 1417 1938
rect 1298 1738 1302 1741
rect 1370 1648 1377 1651
rect 1238 1458 1246 1461
rect 1246 1422 1249 1458
rect 1254 1162 1257 1548
rect 1282 1478 1286 1481
rect 1302 1462 1305 1478
rect 1374 1462 1377 1648
rect 1392 1603 1394 1607
rect 1398 1603 1401 1607
rect 1406 1603 1408 1607
rect 1426 1458 1430 1461
rect 1270 992 1273 1368
rect 1278 1152 1281 1158
rect 1294 1132 1297 1458
rect 1350 1452 1353 1458
rect 1350 1252 1353 1358
rect 1358 1222 1361 1438
rect 1392 1403 1394 1407
rect 1398 1403 1401 1407
rect 1406 1403 1408 1407
rect 1410 1358 1414 1361
rect 1386 1348 1390 1351
rect 1366 1342 1369 1348
rect 1438 1342 1441 1568
rect 1470 1552 1473 1858
rect 1474 1548 1478 1551
rect 1454 1372 1457 1548
rect 1470 1492 1473 1548
rect 1454 1352 1457 1358
rect 1462 1342 1465 1458
rect 1478 1442 1481 1488
rect 1498 1458 1502 1461
rect 1498 1448 1502 1451
rect 1374 1312 1377 1338
rect 1218 638 1225 641
rect 1194 568 1198 571
rect 1126 282 1129 428
rect 942 142 945 268
rect 1158 161 1161 558
rect 1222 542 1225 638
rect 1234 568 1238 571
rect 1246 532 1249 948
rect 1258 928 1262 931
rect 1262 541 1265 748
rect 1286 572 1289 1088
rect 1294 932 1297 1128
rect 1350 882 1353 1098
rect 1362 1048 1366 1051
rect 1382 952 1385 1248
rect 1392 1203 1394 1207
rect 1398 1203 1401 1207
rect 1406 1203 1408 1207
rect 1414 1142 1417 1338
rect 1434 1268 1438 1271
rect 1422 1132 1425 1208
rect 1392 1003 1394 1007
rect 1398 1003 1401 1007
rect 1406 1003 1408 1007
rect 1422 982 1425 1128
rect 1446 1032 1449 1328
rect 1462 1252 1465 1338
rect 1462 1042 1465 1048
rect 1486 992 1489 1128
rect 1358 918 1366 921
rect 1258 538 1265 541
rect 1174 362 1177 368
rect 1174 302 1177 328
rect 1262 182 1265 538
rect 1302 362 1305 698
rect 1358 652 1361 918
rect 1392 803 1394 807
rect 1398 803 1401 807
rect 1406 803 1408 807
rect 1374 472 1377 768
rect 1392 603 1394 607
rect 1398 603 1401 607
rect 1406 603 1408 607
rect 1392 403 1394 407
rect 1398 403 1401 407
rect 1406 403 1408 407
rect 1392 203 1394 207
rect 1398 203 1401 207
rect 1406 203 1408 207
rect 1414 202 1417 548
rect 1422 482 1425 658
rect 1430 612 1433 748
rect 1446 632 1449 958
rect 1454 662 1457 678
rect 1430 422 1433 608
rect 1478 552 1481 968
rect 1486 772 1489 978
rect 1486 692 1489 698
rect 1462 522 1465 538
rect 1422 232 1425 298
rect 1262 172 1265 178
rect 1154 158 1161 161
rect 1414 162 1417 198
rect 1150 152 1153 158
rect 1478 132 1481 548
rect 1494 542 1497 1068
rect 1502 561 1505 1138
rect 1510 1012 1513 1348
rect 1518 1162 1521 1828
rect 1550 1822 1553 1838
rect 1526 1692 1529 1738
rect 1526 1472 1529 1688
rect 1534 1622 1537 1818
rect 1558 1662 1561 1668
rect 1534 1401 1537 1418
rect 1530 1398 1537 1401
rect 1542 1382 1545 1558
rect 1542 1182 1545 1368
rect 1518 642 1521 1148
rect 1526 952 1529 958
rect 1542 942 1545 948
rect 1550 912 1553 1528
rect 1558 1412 1561 1658
rect 1574 1652 1577 1998
rect 1606 1872 1609 1968
rect 1590 1742 1593 1868
rect 1610 1788 1617 1791
rect 1614 1392 1617 1788
rect 1638 1452 1641 1958
rect 1754 1878 1758 1881
rect 1786 1878 1790 1881
rect 1854 1862 1857 1928
rect 1912 1903 1914 1907
rect 1918 1903 1921 1907
rect 1926 1903 1928 1907
rect 1678 1422 1681 1708
rect 1566 1322 1569 1358
rect 1578 1328 1585 1331
rect 1558 1162 1561 1168
rect 1566 1062 1569 1318
rect 1582 1072 1585 1328
rect 1578 1058 1582 1061
rect 1570 1048 1574 1051
rect 1598 1042 1601 1068
rect 1606 1022 1609 1158
rect 1530 888 1534 891
rect 1542 882 1545 898
rect 1566 872 1569 878
rect 1526 852 1529 868
rect 1502 558 1513 561
rect 1486 312 1489 458
rect 1494 112 1497 538
rect 1502 422 1505 528
rect 1510 342 1513 558
rect 1534 442 1537 838
rect 1574 692 1577 938
rect 1594 868 1598 871
rect 1586 688 1590 691
rect 1542 672 1545 678
rect 1554 668 1558 671
rect 1614 372 1617 1388
rect 1686 1251 1689 1708
rect 1786 1648 1790 1651
rect 1694 1432 1697 1648
rect 1798 1562 1801 1758
rect 1810 1538 1814 1541
rect 1686 1248 1694 1251
rect 1706 1248 1710 1251
rect 1658 1238 1662 1241
rect 1614 362 1617 368
rect 1510 292 1513 338
rect 1514 268 1518 271
rect 1614 252 1617 288
rect 880 103 882 107
rect 886 103 889 107
rect 894 103 896 107
rect 378 68 382 71
rect 458 68 462 71
rect 790 52 793 78
rect 854 62 857 88
rect 1622 12 1625 368
rect 1630 282 1633 1028
rect 1638 852 1641 1148
rect 1646 382 1649 1228
rect 1758 1162 1761 1528
rect 1798 1432 1801 1518
rect 1806 1462 1809 1528
rect 1770 1338 1774 1341
rect 1750 1152 1753 1158
rect 1662 1072 1665 1148
rect 1718 952 1721 1028
rect 1766 892 1769 1128
rect 1718 692 1721 748
rect 1682 688 1689 691
rect 1686 682 1689 688
rect 1710 672 1713 688
rect 1638 372 1641 378
rect 1674 368 1678 371
rect 1666 268 1670 271
rect 1726 172 1729 648
rect 1734 552 1737 748
rect 1742 672 1745 868
rect 1782 862 1785 1348
rect 1758 842 1761 848
rect 1770 768 1774 771
rect 1762 668 1766 671
rect 1774 632 1777 728
rect 1782 592 1785 858
rect 1790 772 1793 1108
rect 1798 1072 1801 1428
rect 1806 1262 1809 1458
rect 1838 1342 1841 1578
rect 1806 1112 1809 1258
rect 1826 1158 1830 1161
rect 1798 802 1801 1068
rect 1806 842 1809 1068
rect 1822 852 1825 1158
rect 1842 1148 1846 1151
rect 1830 892 1833 1048
rect 1854 992 1857 1858
rect 2014 1752 2017 1998
rect 1912 1703 1914 1707
rect 1918 1703 1921 1707
rect 1926 1703 1928 1707
rect 1870 1652 1873 1658
rect 1862 1342 1865 1358
rect 1878 1261 1881 1698
rect 2022 1622 2025 2048
rect 1912 1503 1914 1507
rect 1918 1503 1921 1507
rect 1926 1503 1928 1507
rect 1966 1472 1969 1548
rect 1990 1542 1993 1548
rect 1902 1292 1905 1308
rect 1912 1303 1914 1307
rect 1918 1303 1921 1307
rect 1926 1303 1928 1307
rect 1878 1258 1886 1261
rect 1886 1062 1889 1258
rect 1910 1252 1913 1258
rect 1838 898 1846 901
rect 1838 732 1841 898
rect 1838 672 1841 728
rect 1854 722 1857 948
rect 1862 852 1865 1038
rect 1874 948 1878 951
rect 1838 562 1841 668
rect 1862 652 1865 748
rect 1846 438 1854 441
rect 1846 242 1849 438
rect 1870 192 1873 948
rect 1878 752 1881 768
rect 1894 662 1897 1198
rect 1912 1103 1914 1107
rect 1918 1103 1921 1107
rect 1926 1103 1928 1107
rect 1912 903 1914 907
rect 1918 903 1921 907
rect 1926 903 1928 907
rect 1902 772 1905 898
rect 1958 852 1961 1328
rect 1966 1312 1969 1468
rect 1982 1362 1985 1498
rect 1974 1312 1977 1358
rect 1978 948 1982 951
rect 1912 703 1914 707
rect 1918 703 1921 707
rect 1926 703 1928 707
rect 1934 638 1942 641
rect 1902 342 1905 508
rect 1912 503 1914 507
rect 1918 503 1921 507
rect 1926 503 1928 507
rect 1934 312 1937 638
rect 1958 412 1961 848
rect 1990 742 1993 1538
rect 2022 962 2025 1218
rect 1998 932 2001 938
rect 2014 552 2017 758
rect 2030 752 2033 1758
rect 2070 1482 2073 1578
rect 2078 1351 2081 1538
rect 2074 1348 2081 1351
rect 2046 932 2049 1138
rect 2070 1072 2073 1338
rect 2078 1092 2081 1298
rect 2058 948 2062 951
rect 2046 752 2049 928
rect 2014 482 2017 548
rect 1912 303 1914 307
rect 1918 303 1921 307
rect 1926 303 1928 307
rect 1934 232 1937 308
rect 2006 262 2009 468
rect 2030 452 2033 718
rect 2070 562 2073 1008
rect 2078 862 2081 1088
rect 2078 462 2081 858
rect 2094 651 2097 1768
rect 2102 1272 2105 1558
rect 2110 1462 2113 2018
rect 2134 1552 2137 2058
rect 2174 1762 2177 2048
rect 2142 1542 2145 1548
rect 2150 1522 2153 1758
rect 2110 1162 2113 1378
rect 2110 1052 2113 1158
rect 2166 1152 2169 1498
rect 2094 648 2102 651
rect 2110 632 2113 1048
rect 2030 362 2033 448
rect 2046 262 2049 278
rect 1912 103 1914 107
rect 1918 103 1921 107
rect 1926 103 1928 107
rect 2006 92 2009 258
rect 2174 142 2177 1758
rect 2182 1272 2185 1338
rect 2190 1142 2193 1918
rect 2198 1672 2201 1828
rect 2190 732 2193 848
rect 2198 742 2201 1668
rect 2210 1548 2214 1551
rect 2190 252 2193 488
rect 2198 182 2201 738
rect 2206 332 2209 1438
rect 2222 1102 2225 2068
rect 2230 852 2233 2068
rect 2246 1442 2249 2058
rect 2258 2018 2265 2021
rect 2246 222 2249 658
rect 2254 262 2257 1238
rect 2262 1012 2265 2018
rect 2278 902 2281 1108
rect 2286 1082 2289 2048
rect 2298 848 2302 851
rect 2298 768 2302 771
rect 2262 162 2265 358
rect 2286 272 2289 538
rect 376 3 378 7
rect 382 3 385 7
rect 390 3 392 7
rect 1392 3 1394 7
rect 1398 3 1401 7
rect 1406 3 1408 7
<< m5contact >>
rect 882 2103 886 2107
rect 889 2103 890 2107
rect 890 2103 893 2107
rect 1914 2103 1918 2107
rect 1921 2103 1922 2107
rect 1922 2103 1925 2107
rect 286 2058 290 2062
rect 326 2058 330 2062
rect 302 2048 306 2052
rect 582 2048 586 2052
rect 758 2048 762 2052
rect 378 2003 382 2007
rect 385 2003 386 2007
rect 386 2003 389 2007
rect 182 1918 186 1922
rect 378 1803 382 1807
rect 385 1803 386 1807
rect 386 1803 389 1807
rect 142 1258 146 1262
rect 198 1068 202 1072
rect 310 1468 314 1472
rect 378 1603 382 1607
rect 385 1603 386 1607
rect 386 1603 389 1607
rect 378 1403 382 1407
rect 385 1403 386 1407
rect 386 1403 389 1407
rect 246 1068 250 1072
rect 286 458 290 462
rect 378 1203 382 1207
rect 385 1203 386 1207
rect 386 1203 389 1207
rect 334 458 338 462
rect 334 348 338 352
rect 378 1003 382 1007
rect 385 1003 386 1007
rect 386 1003 389 1007
rect 378 803 382 807
rect 385 803 386 807
rect 386 803 389 807
rect 454 1458 458 1462
rect 478 1148 482 1152
rect 378 603 382 607
rect 385 603 386 607
rect 386 603 389 607
rect 590 1918 594 1922
rect 598 1838 602 1842
rect 622 1358 626 1362
rect 710 1738 714 1742
rect 678 1658 682 1662
rect 670 1258 674 1262
rect 702 1148 706 1152
rect 630 928 634 932
rect 526 878 530 882
rect 378 403 382 407
rect 385 403 386 407
rect 386 403 389 407
rect 494 358 498 362
rect 646 738 650 742
rect 654 728 658 732
rect 378 203 382 207
rect 385 203 386 207
rect 386 203 389 207
rect 438 148 442 152
rect 574 338 578 342
rect 882 1903 886 1907
rect 889 1903 890 1907
rect 890 1903 893 1907
rect 790 1468 794 1472
rect 758 888 762 892
rect 758 668 762 672
rect 806 1348 810 1352
rect 950 1838 954 1842
rect 882 1703 886 1707
rect 889 1703 890 1707
rect 890 1703 893 1707
rect 1014 1648 1018 1652
rect 882 1503 886 1507
rect 889 1503 890 1507
rect 890 1503 893 1507
rect 870 1478 874 1482
rect 882 1303 886 1307
rect 889 1303 890 1307
rect 890 1303 893 1307
rect 862 1158 866 1162
rect 846 1148 850 1152
rect 782 1128 786 1132
rect 774 948 778 952
rect 882 1103 886 1107
rect 889 1103 890 1107
rect 890 1103 893 1107
rect 882 903 886 907
rect 889 903 890 907
rect 890 903 893 907
rect 742 368 746 372
rect 750 328 754 332
rect 882 703 886 707
rect 889 703 890 707
rect 890 703 893 707
rect 882 503 886 507
rect 889 503 890 507
rect 890 503 893 507
rect 918 1348 922 1352
rect 882 303 886 307
rect 889 303 890 307
rect 890 303 893 307
rect 910 348 914 352
rect 998 1038 1002 1042
rect 1022 1448 1026 1452
rect 1038 1248 1042 1252
rect 1030 1148 1034 1152
rect 1022 1128 1026 1132
rect 1014 1028 1018 1032
rect 998 688 1002 692
rect 1022 708 1026 712
rect 990 418 994 422
rect 1054 978 1058 982
rect 1182 1538 1186 1542
rect 1102 1348 1106 1352
rect 1110 1258 1114 1262
rect 1102 1168 1106 1172
rect 1086 978 1090 982
rect 1142 1278 1146 1282
rect 1134 1238 1138 1242
rect 1062 728 1066 732
rect 1038 338 1042 342
rect 1014 288 1018 292
rect 1126 688 1130 692
rect 1150 748 1154 752
rect 1166 1248 1170 1252
rect 1166 1138 1170 1142
rect 1206 1258 1210 1262
rect 1198 1148 1202 1152
rect 1214 1058 1218 1062
rect 1166 708 1170 712
rect 1190 738 1194 742
rect 1262 1648 1266 1652
rect 1394 2003 1398 2007
rect 1401 2003 1402 2007
rect 1402 2003 1405 2007
rect 1394 1803 1398 1807
rect 1401 1803 1402 1807
rect 1402 1803 1405 1807
rect 1302 1738 1306 1742
rect 1246 1418 1250 1422
rect 1286 1478 1290 1482
rect 1394 1603 1398 1607
rect 1401 1603 1402 1607
rect 1402 1603 1405 1607
rect 1302 1458 1306 1462
rect 1350 1458 1354 1462
rect 1422 1458 1426 1462
rect 1278 1158 1282 1162
rect 1394 1403 1398 1407
rect 1401 1403 1402 1407
rect 1402 1403 1405 1407
rect 1406 1358 1410 1362
rect 1390 1348 1394 1352
rect 1550 1838 1554 1842
rect 1478 1548 1482 1552
rect 1454 1348 1458 1352
rect 1502 1458 1506 1462
rect 1494 1448 1498 1452
rect 1366 1338 1370 1342
rect 1294 1128 1298 1132
rect 1198 568 1202 572
rect 1126 278 1130 282
rect 1238 568 1242 572
rect 1262 928 1266 932
rect 1366 1048 1370 1052
rect 1394 1203 1398 1207
rect 1401 1203 1402 1207
rect 1402 1203 1405 1207
rect 1438 1268 1442 1272
rect 1394 1003 1398 1007
rect 1401 1003 1402 1007
rect 1402 1003 1405 1007
rect 1462 1038 1466 1042
rect 1174 368 1178 372
rect 1174 328 1178 332
rect 1394 803 1398 807
rect 1401 803 1402 807
rect 1402 803 1405 807
rect 1394 603 1398 607
rect 1401 603 1402 607
rect 1402 603 1405 607
rect 1394 403 1398 407
rect 1401 403 1402 407
rect 1402 403 1405 407
rect 1394 203 1398 207
rect 1401 203 1402 207
rect 1402 203 1405 207
rect 1486 698 1490 702
rect 1430 418 1434 422
rect 1150 148 1154 152
rect 1526 1738 1530 1742
rect 1558 1658 1562 1662
rect 1534 1418 1538 1422
rect 1526 958 1530 962
rect 1542 948 1546 952
rect 1758 1878 1762 1882
rect 1782 1878 1786 1882
rect 1914 1903 1918 1907
rect 1921 1903 1922 1907
rect 1922 1903 1925 1907
rect 1558 1168 1562 1172
rect 1606 1158 1610 1162
rect 1582 1058 1586 1062
rect 1566 1048 1570 1052
rect 1574 938 1578 942
rect 1534 888 1538 892
rect 1566 878 1570 882
rect 1526 868 1530 872
rect 1590 868 1594 872
rect 1590 688 1594 692
rect 1542 678 1546 682
rect 1550 668 1554 672
rect 1790 1648 1794 1652
rect 1814 1538 1818 1542
rect 1710 1248 1714 1252
rect 1654 1238 1658 1242
rect 1614 358 1618 362
rect 1510 288 1514 292
rect 1518 268 1522 272
rect 882 103 886 107
rect 889 103 890 107
rect 890 103 893 107
rect 382 68 386 72
rect 454 68 458 72
rect 1806 1458 1810 1462
rect 1766 1338 1770 1342
rect 1750 1148 1754 1152
rect 1718 1028 1722 1032
rect 1718 748 1722 752
rect 1686 678 1690 682
rect 1710 668 1714 672
rect 1638 368 1642 372
rect 1678 368 1682 372
rect 1662 268 1666 272
rect 1758 848 1762 852
rect 1774 768 1778 772
rect 1766 668 1770 672
rect 1822 1158 1826 1162
rect 1838 1148 1842 1152
rect 1914 1703 1918 1707
rect 1921 1703 1922 1707
rect 1922 1703 1925 1707
rect 1870 1658 1874 1662
rect 1862 1338 1866 1342
rect 1990 1548 1994 1552
rect 1914 1503 1918 1507
rect 1921 1503 1922 1507
rect 1922 1503 1925 1507
rect 1914 1303 1918 1307
rect 1921 1303 1922 1307
rect 1922 1303 1925 1307
rect 1910 1248 1914 1252
rect 1870 948 1874 952
rect 1914 1103 1918 1107
rect 1921 1103 1922 1107
rect 1922 1103 1925 1107
rect 1914 903 1918 907
rect 1921 903 1922 907
rect 1922 903 1925 907
rect 1982 948 1986 952
rect 1914 703 1918 707
rect 1921 703 1922 707
rect 1922 703 1925 707
rect 1914 503 1918 507
rect 1921 503 1922 507
rect 1922 503 1925 507
rect 1998 928 2002 932
rect 2054 948 2058 952
rect 1914 303 1918 307
rect 1921 303 1922 307
rect 1922 303 1925 307
rect 2142 1548 2146 1552
rect 2046 278 2050 282
rect 1914 103 1918 107
rect 1921 103 1922 107
rect 1922 103 1925 107
rect 2214 1548 2218 1552
rect 2294 848 2298 852
rect 2294 768 2298 772
rect 378 3 382 7
rect 385 3 386 7
rect 386 3 389 7
rect 1394 3 1398 7
rect 1401 3 1402 7
rect 1402 3 1405 7
<< metal5 >>
rect 886 2103 889 2107
rect 885 2102 890 2103
rect 895 2102 896 2107
rect 1918 2103 1921 2107
rect 1917 2102 1922 2103
rect 1927 2102 1928 2107
rect 290 2058 326 2061
rect 306 2048 582 2051
rect 586 2048 758 2051
rect 382 2003 385 2007
rect 381 2002 386 2003
rect 391 2002 392 2007
rect 1398 2003 1401 2007
rect 1397 2002 1402 2003
rect 1407 2002 1408 2007
rect 186 1918 590 1921
rect 886 1903 889 1907
rect 885 1902 890 1903
rect 895 1902 896 1907
rect 1918 1903 1921 1907
rect 1917 1902 1922 1903
rect 1927 1902 1928 1907
rect 1762 1878 1782 1881
rect 602 1838 950 1841
rect 954 1838 1550 1841
rect 382 1803 385 1807
rect 381 1802 386 1803
rect 391 1802 392 1807
rect 1398 1803 1401 1807
rect 1397 1802 1402 1803
rect 1407 1802 1408 1807
rect 714 1738 1302 1741
rect 1306 1738 1526 1741
rect 886 1703 889 1707
rect 885 1702 890 1703
rect 895 1702 896 1707
rect 1918 1703 1921 1707
rect 1917 1702 1922 1703
rect 1927 1702 1928 1707
rect 682 1658 1558 1661
rect 1018 1648 1262 1651
rect 1870 1651 1873 1658
rect 1794 1648 1873 1651
rect 382 1603 385 1607
rect 381 1602 386 1603
rect 391 1602 392 1607
rect 1398 1603 1401 1607
rect 1397 1602 1402 1603
rect 1407 1602 1408 1607
rect 1482 1548 1990 1551
rect 2146 1548 2214 1551
rect 1186 1538 1814 1541
rect 886 1503 889 1507
rect 885 1502 890 1503
rect 895 1502 896 1507
rect 1918 1503 1921 1507
rect 1917 1502 1922 1503
rect 1927 1502 1928 1507
rect 874 1478 1286 1481
rect 314 1468 790 1471
rect 458 1458 1302 1461
rect 1354 1458 1422 1461
rect 1506 1458 1806 1461
rect 1026 1448 1494 1451
rect 1250 1418 1534 1421
rect 382 1403 385 1407
rect 381 1402 386 1403
rect 391 1402 392 1407
rect 1398 1403 1401 1407
rect 1397 1402 1402 1403
rect 1407 1402 1408 1407
rect 626 1358 1406 1361
rect 810 1348 918 1351
rect 1106 1348 1369 1351
rect 1394 1348 1454 1351
rect 1366 1342 1369 1348
rect 1770 1338 1862 1341
rect 886 1303 889 1307
rect 885 1302 890 1303
rect 895 1302 896 1307
rect 1918 1303 1921 1307
rect 1917 1302 1922 1303
rect 1927 1302 1928 1307
rect 1142 1271 1145 1278
rect 1142 1268 1438 1271
rect 146 1258 670 1261
rect 1114 1258 1206 1261
rect 1042 1248 1166 1251
rect 1714 1248 1910 1251
rect 1138 1238 1654 1241
rect 382 1203 385 1207
rect 381 1202 386 1203
rect 391 1202 392 1207
rect 1398 1203 1401 1207
rect 1397 1202 1402 1203
rect 1407 1202 1408 1207
rect 1106 1168 1558 1171
rect 866 1158 1278 1161
rect 1610 1158 1822 1161
rect 482 1148 702 1151
rect 706 1148 846 1151
rect 850 1148 1030 1151
rect 1034 1148 1198 1151
rect 1754 1148 1838 1151
rect 782 1138 1166 1141
rect 782 1132 785 1138
rect 1026 1128 1294 1131
rect 886 1103 889 1107
rect 885 1102 890 1103
rect 895 1102 896 1107
rect 1918 1103 1921 1107
rect 1917 1102 1922 1103
rect 1927 1102 1928 1107
rect 202 1068 246 1071
rect 1218 1058 1582 1061
rect 1370 1048 1566 1051
rect 1002 1038 1462 1041
rect 1018 1028 1718 1031
rect 382 1003 385 1007
rect 381 1002 386 1003
rect 391 1002 392 1007
rect 1398 1003 1401 1007
rect 1397 1002 1402 1003
rect 1407 1002 1408 1007
rect 1058 978 1086 981
rect 1526 951 1529 958
rect 778 948 1529 951
rect 1546 948 1870 951
rect 1986 948 2054 951
rect 1578 938 2001 941
rect 1998 932 2001 938
rect 634 928 1262 931
rect 886 903 889 907
rect 885 902 890 903
rect 895 902 896 907
rect 1918 903 1921 907
rect 1917 902 1922 903
rect 1927 902 1928 907
rect 762 888 1534 891
rect 530 878 1566 881
rect 1530 868 1590 871
rect 1762 848 2294 851
rect 382 803 385 807
rect 381 802 386 803
rect 391 802 392 807
rect 1398 803 1401 807
rect 1397 802 1402 803
rect 1407 802 1408 807
rect 1778 768 2294 771
rect 1154 748 1718 751
rect 650 738 1190 741
rect 658 728 1062 731
rect 1026 708 1166 711
rect 886 703 889 707
rect 885 702 890 703
rect 895 702 896 707
rect 1918 703 1921 707
rect 1917 702 1922 703
rect 1927 702 1928 707
rect 1486 691 1489 698
rect 1486 688 1590 691
rect 998 681 1001 688
rect 1126 681 1129 688
rect 998 678 1129 681
rect 1546 678 1686 681
rect 762 668 1550 671
rect 1714 668 1766 671
rect 382 603 385 607
rect 381 602 386 603
rect 391 602 392 607
rect 1398 603 1401 607
rect 1397 602 1402 603
rect 1407 602 1408 607
rect 1202 568 1238 571
rect 886 503 889 507
rect 885 502 890 503
rect 895 502 896 507
rect 1918 503 1921 507
rect 1917 502 1922 503
rect 1927 502 1928 507
rect 290 458 334 461
rect 994 418 1430 421
rect 382 403 385 407
rect 381 402 386 403
rect 391 402 392 407
rect 1398 403 1401 407
rect 1397 402 1402 403
rect 1407 402 1408 407
rect 746 368 1174 371
rect 1642 368 1678 371
rect 498 358 1614 361
rect 338 348 910 351
rect 578 338 1038 341
rect 754 328 1174 331
rect 886 303 889 307
rect 885 302 890 303
rect 895 302 896 307
rect 1918 303 1921 307
rect 1917 302 1922 303
rect 1927 302 1928 307
rect 1018 288 1510 291
rect 1130 278 2046 281
rect 1522 268 1662 271
rect 382 203 385 207
rect 381 202 386 203
rect 391 202 392 207
rect 1398 203 1401 207
rect 1397 202 1402 203
rect 1407 202 1408 207
rect 442 148 1150 151
rect 886 103 889 107
rect 885 102 890 103
rect 895 102 896 107
rect 1918 103 1921 107
rect 1917 102 1922 103
rect 1927 102 1928 107
rect 386 68 454 71
rect 382 3 385 7
rect 381 2 386 3
rect 391 2 392 7
rect 1398 3 1401 7
rect 1397 2 1402 3
rect 1407 2 1408 7
<< m6contact >>
rect 880 2103 882 2107
rect 882 2103 885 2107
rect 890 2103 893 2107
rect 893 2103 895 2107
rect 880 2102 885 2103
rect 890 2102 895 2103
rect 1912 2103 1914 2107
rect 1914 2103 1917 2107
rect 1922 2103 1925 2107
rect 1925 2103 1927 2107
rect 1912 2102 1917 2103
rect 1922 2102 1927 2103
rect 376 2003 378 2007
rect 378 2003 381 2007
rect 386 2003 389 2007
rect 389 2003 391 2007
rect 376 2002 381 2003
rect 386 2002 391 2003
rect 1392 2003 1394 2007
rect 1394 2003 1397 2007
rect 1402 2003 1405 2007
rect 1405 2003 1407 2007
rect 1392 2002 1397 2003
rect 1402 2002 1407 2003
rect 880 1903 882 1907
rect 882 1903 885 1907
rect 890 1903 893 1907
rect 893 1903 895 1907
rect 880 1902 885 1903
rect 890 1902 895 1903
rect 1912 1903 1914 1907
rect 1914 1903 1917 1907
rect 1922 1903 1925 1907
rect 1925 1903 1927 1907
rect 1912 1902 1917 1903
rect 1922 1902 1927 1903
rect 376 1803 378 1807
rect 378 1803 381 1807
rect 386 1803 389 1807
rect 389 1803 391 1807
rect 376 1802 381 1803
rect 386 1802 391 1803
rect 1392 1803 1394 1807
rect 1394 1803 1397 1807
rect 1402 1803 1405 1807
rect 1405 1803 1407 1807
rect 1392 1802 1397 1803
rect 1402 1802 1407 1803
rect 880 1703 882 1707
rect 882 1703 885 1707
rect 890 1703 893 1707
rect 893 1703 895 1707
rect 880 1702 885 1703
rect 890 1702 895 1703
rect 1912 1703 1914 1707
rect 1914 1703 1917 1707
rect 1922 1703 1925 1707
rect 1925 1703 1927 1707
rect 1912 1702 1917 1703
rect 1922 1702 1927 1703
rect 376 1603 378 1607
rect 378 1603 381 1607
rect 386 1603 389 1607
rect 389 1603 391 1607
rect 376 1602 381 1603
rect 386 1602 391 1603
rect 1392 1603 1394 1607
rect 1394 1603 1397 1607
rect 1402 1603 1405 1607
rect 1405 1603 1407 1607
rect 1392 1602 1397 1603
rect 1402 1602 1407 1603
rect 880 1503 882 1507
rect 882 1503 885 1507
rect 890 1503 893 1507
rect 893 1503 895 1507
rect 880 1502 885 1503
rect 890 1502 895 1503
rect 1912 1503 1914 1507
rect 1914 1503 1917 1507
rect 1922 1503 1925 1507
rect 1925 1503 1927 1507
rect 1912 1502 1917 1503
rect 1922 1502 1927 1503
rect 376 1403 378 1407
rect 378 1403 381 1407
rect 386 1403 389 1407
rect 389 1403 391 1407
rect 376 1402 381 1403
rect 386 1402 391 1403
rect 1392 1403 1394 1407
rect 1394 1403 1397 1407
rect 1402 1403 1405 1407
rect 1405 1403 1407 1407
rect 1392 1402 1397 1403
rect 1402 1402 1407 1403
rect 880 1303 882 1307
rect 882 1303 885 1307
rect 890 1303 893 1307
rect 893 1303 895 1307
rect 880 1302 885 1303
rect 890 1302 895 1303
rect 1912 1303 1914 1307
rect 1914 1303 1917 1307
rect 1922 1303 1925 1307
rect 1925 1303 1927 1307
rect 1912 1302 1917 1303
rect 1922 1302 1927 1303
rect 376 1203 378 1207
rect 378 1203 381 1207
rect 386 1203 389 1207
rect 389 1203 391 1207
rect 376 1202 381 1203
rect 386 1202 391 1203
rect 1392 1203 1394 1207
rect 1394 1203 1397 1207
rect 1402 1203 1405 1207
rect 1405 1203 1407 1207
rect 1392 1202 1397 1203
rect 1402 1202 1407 1203
rect 880 1103 882 1107
rect 882 1103 885 1107
rect 890 1103 893 1107
rect 893 1103 895 1107
rect 880 1102 885 1103
rect 890 1102 895 1103
rect 1912 1103 1914 1107
rect 1914 1103 1917 1107
rect 1922 1103 1925 1107
rect 1925 1103 1927 1107
rect 1912 1102 1917 1103
rect 1922 1102 1927 1103
rect 376 1003 378 1007
rect 378 1003 381 1007
rect 386 1003 389 1007
rect 389 1003 391 1007
rect 376 1002 381 1003
rect 386 1002 391 1003
rect 1392 1003 1394 1007
rect 1394 1003 1397 1007
rect 1402 1003 1405 1007
rect 1405 1003 1407 1007
rect 1392 1002 1397 1003
rect 1402 1002 1407 1003
rect 880 903 882 907
rect 882 903 885 907
rect 890 903 893 907
rect 893 903 895 907
rect 880 902 885 903
rect 890 902 895 903
rect 1912 903 1914 907
rect 1914 903 1917 907
rect 1922 903 1925 907
rect 1925 903 1927 907
rect 1912 902 1917 903
rect 1922 902 1927 903
rect 376 803 378 807
rect 378 803 381 807
rect 386 803 389 807
rect 389 803 391 807
rect 376 802 381 803
rect 386 802 391 803
rect 1392 803 1394 807
rect 1394 803 1397 807
rect 1402 803 1405 807
rect 1405 803 1407 807
rect 1392 802 1397 803
rect 1402 802 1407 803
rect 880 703 882 707
rect 882 703 885 707
rect 890 703 893 707
rect 893 703 895 707
rect 880 702 885 703
rect 890 702 895 703
rect 1912 703 1914 707
rect 1914 703 1917 707
rect 1922 703 1925 707
rect 1925 703 1927 707
rect 1912 702 1917 703
rect 1922 702 1927 703
rect 376 603 378 607
rect 378 603 381 607
rect 386 603 389 607
rect 389 603 391 607
rect 376 602 381 603
rect 386 602 391 603
rect 1392 603 1394 607
rect 1394 603 1397 607
rect 1402 603 1405 607
rect 1405 603 1407 607
rect 1392 602 1397 603
rect 1402 602 1407 603
rect 880 503 882 507
rect 882 503 885 507
rect 890 503 893 507
rect 893 503 895 507
rect 880 502 885 503
rect 890 502 895 503
rect 1912 503 1914 507
rect 1914 503 1917 507
rect 1922 503 1925 507
rect 1925 503 1927 507
rect 1912 502 1917 503
rect 1922 502 1927 503
rect 376 403 378 407
rect 378 403 381 407
rect 386 403 389 407
rect 389 403 391 407
rect 376 402 381 403
rect 386 402 391 403
rect 1392 403 1394 407
rect 1394 403 1397 407
rect 1402 403 1405 407
rect 1405 403 1407 407
rect 1392 402 1397 403
rect 1402 402 1407 403
rect 880 303 882 307
rect 882 303 885 307
rect 890 303 893 307
rect 893 303 895 307
rect 880 302 885 303
rect 890 302 895 303
rect 1912 303 1914 307
rect 1914 303 1917 307
rect 1922 303 1925 307
rect 1925 303 1927 307
rect 1912 302 1917 303
rect 1922 302 1927 303
rect 376 203 378 207
rect 378 203 381 207
rect 386 203 389 207
rect 389 203 391 207
rect 376 202 381 203
rect 386 202 391 203
rect 1392 203 1394 207
rect 1394 203 1397 207
rect 1402 203 1405 207
rect 1405 203 1407 207
rect 1392 202 1397 203
rect 1402 202 1407 203
rect 880 103 882 107
rect 882 103 885 107
rect 890 103 893 107
rect 893 103 895 107
rect 880 102 885 103
rect 890 102 895 103
rect 1912 103 1914 107
rect 1914 103 1917 107
rect 1922 103 1925 107
rect 1925 103 1927 107
rect 1912 102 1917 103
rect 1922 102 1927 103
rect 376 3 378 7
rect 378 3 381 7
rect 386 3 389 7
rect 389 3 391 7
rect 376 2 381 3
rect 386 2 391 3
rect 1392 3 1394 7
rect 1394 3 1397 7
rect 1402 3 1405 7
rect 1405 3 1407 7
rect 1392 2 1397 3
rect 1402 2 1407 3
<< metal6 >>
rect 376 2007 392 2130
rect 381 2002 386 2007
rect 391 2002 392 2007
rect 376 1807 392 2002
rect 381 1802 386 1807
rect 391 1802 392 1807
rect 376 1607 392 1802
rect 381 1602 386 1607
rect 391 1602 392 1607
rect 376 1407 392 1602
rect 381 1402 386 1407
rect 391 1402 392 1407
rect 376 1207 392 1402
rect 381 1202 386 1207
rect 391 1202 392 1207
rect 376 1007 392 1202
rect 381 1002 386 1007
rect 391 1002 392 1007
rect 376 807 392 1002
rect 381 802 386 807
rect 391 802 392 807
rect 376 607 392 802
rect 381 602 386 607
rect 391 602 392 607
rect 376 407 392 602
rect 381 402 386 407
rect 391 402 392 407
rect 376 207 392 402
rect 381 202 386 207
rect 391 202 392 207
rect 376 7 392 202
rect 381 2 386 7
rect 391 2 392 7
rect 376 -30 392 2
rect 880 2107 896 2130
rect 885 2102 890 2107
rect 895 2102 896 2107
rect 880 1907 896 2102
rect 885 1902 890 1907
rect 895 1902 896 1907
rect 880 1707 896 1902
rect 885 1702 890 1707
rect 895 1702 896 1707
rect 880 1507 896 1702
rect 885 1502 890 1507
rect 895 1502 896 1507
rect 880 1307 896 1502
rect 885 1302 890 1307
rect 895 1302 896 1307
rect 880 1107 896 1302
rect 885 1102 890 1107
rect 895 1102 896 1107
rect 880 907 896 1102
rect 885 902 890 907
rect 895 902 896 907
rect 880 707 896 902
rect 885 702 890 707
rect 895 702 896 707
rect 880 507 896 702
rect 885 502 890 507
rect 895 502 896 507
rect 880 307 896 502
rect 885 302 890 307
rect 895 302 896 307
rect 880 107 896 302
rect 885 102 890 107
rect 895 102 896 107
rect 880 -30 896 102
rect 1392 2007 1408 2130
rect 1397 2002 1402 2007
rect 1407 2002 1408 2007
rect 1392 1807 1408 2002
rect 1397 1802 1402 1807
rect 1407 1802 1408 1807
rect 1392 1607 1408 1802
rect 1397 1602 1402 1607
rect 1407 1602 1408 1607
rect 1392 1407 1408 1602
rect 1397 1402 1402 1407
rect 1407 1402 1408 1407
rect 1392 1207 1408 1402
rect 1397 1202 1402 1207
rect 1407 1202 1408 1207
rect 1392 1007 1408 1202
rect 1397 1002 1402 1007
rect 1407 1002 1408 1007
rect 1392 807 1408 1002
rect 1397 802 1402 807
rect 1407 802 1408 807
rect 1392 607 1408 802
rect 1397 602 1402 607
rect 1407 602 1408 607
rect 1392 407 1408 602
rect 1397 402 1402 407
rect 1407 402 1408 407
rect 1392 207 1408 402
rect 1397 202 1402 207
rect 1407 202 1408 207
rect 1392 7 1408 202
rect 1397 2 1402 7
rect 1407 2 1408 7
rect 1392 -30 1408 2
rect 1912 2107 1928 2130
rect 1917 2102 1922 2107
rect 1927 2102 1928 2107
rect 1912 1907 1928 2102
rect 1917 1902 1922 1907
rect 1927 1902 1928 1907
rect 1912 1707 1928 1902
rect 1917 1702 1922 1707
rect 1927 1702 1928 1707
rect 1912 1507 1928 1702
rect 1917 1502 1922 1507
rect 1927 1502 1928 1507
rect 1912 1307 1928 1502
rect 1917 1302 1922 1307
rect 1927 1302 1928 1307
rect 1912 1107 1928 1302
rect 1917 1102 1922 1107
rect 1927 1102 1928 1107
rect 1912 907 1928 1102
rect 1917 902 1922 907
rect 1927 902 1928 907
rect 1912 707 1928 902
rect 1917 702 1922 707
rect 1927 702 1928 707
rect 1912 507 1928 702
rect 1917 502 1922 507
rect 1927 502 1928 507
rect 1912 307 1928 502
rect 1917 302 1922 307
rect 1927 302 1928 307
rect 1912 107 1928 302
rect 1917 102 1922 107
rect 1927 102 1928 107
rect 1912 -30 1928 102
use OAI21X1  OAI21X1_217
timestamp 1732943601
transform -1 0 36 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_174
timestamp 1732943601
transform -1 0 60 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_43
timestamp 1732943601
transform -1 0 92 0 -1 105
box -2 -3 34 103
use INVX8  INVX8_10
timestamp 1732943601
transform 1 0 92 0 -1 105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1732943601
transform 1 0 4 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_212
timestamp 1732943601
transform 1 0 100 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1732943601
transform -1 0 156 0 -1 105
box -2 -3 26 103
use INVX8  INVX8_5
timestamp 1732943601
transform 1 0 156 0 -1 105
box -2 -3 42 103
use BUFX4  BUFX4_2
timestamp 1732943601
transform 1 0 196 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1732943601
transform 1 0 132 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_6
timestamp 1732943601
transform 1 0 228 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1732943601
transform 1 0 300 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_22
timestamp 1732943601
transform 1 0 228 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1732943601
transform 1 0 244 0 1 105
box -2 -3 98 103
use FILL  FILL_0_0_0
timestamp 1732943601
transform -1 0 404 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1732943601
transform -1 0 412 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_16
timestamp 1732943601
transform -1 0 372 0 1 105
box -2 -3 34 103
use FILL  FILL_1_0_0
timestamp 1732943601
transform -1 0 380 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1732943601
transform -1 0 388 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_72
timestamp 1732943601
transform -1 0 436 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_15
timestamp 1732943601
transform -1 0 436 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_165
timestamp 1732943601
transform 1 0 436 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_209
timestamp 1732943601
transform -1 0 492 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1732943601
transform -1 0 588 0 -1 105
box -2 -3 98 103
use BUFX4  BUFX4_41
timestamp 1732943601
transform 1 0 436 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1732943601
transform 1 0 468 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1732943601
transform 1 0 588 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_80
timestamp 1732943601
transform 1 0 564 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1732943601
transform -1 0 620 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1732943601
transform 1 0 684 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_49
timestamp 1732943601
transform 1 0 620 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_262
timestamp 1732943601
transform 1 0 636 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_204
timestamp 1732943601
transform -1 0 692 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1732943601
transform 1 0 692 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_2
timestamp 1732943601
transform -1 0 812 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1732943601
transform 1 0 788 0 1 105
box -2 -3 18 103
use INVX2  INVX2_1
timestamp 1732943601
transform 1 0 804 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_74
timestamp 1732943601
transform -1 0 876 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_75
timestamp 1732943601
transform 1 0 820 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1732943601
transform -1 0 868 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1732943601
transform 1 0 812 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1_1
timestamp 1732943601
transform 1 0 884 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_0
timestamp 1732943601
transform 1 0 876 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_11
timestamp 1732943601
transform 1 0 908 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_1
timestamp 1732943601
transform 1 0 900 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_0
timestamp 1732943601
transform 1 0 892 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_4
timestamp 1732943601
transform 1 0 868 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1732943601
transform 1 0 892 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_10
timestamp 1732943601
transform -1 0 964 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1732943601
transform 1 0 964 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_18
timestamp 1732943601
transform 1 0 988 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1732943601
transform 1 0 1004 0 1 105
box -2 -3 98 103
use INVX8  INVX8_7
timestamp 1732943601
transform -1 0 1100 0 -1 105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1732943601
transform 1 0 1100 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_61
timestamp 1732943601
transform 1 0 1100 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1732943601
transform 1 0 1196 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_60
timestamp 1732943601
transform -1 0 1156 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_19
timestamp 1732943601
transform 1 0 1156 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_51
timestamp 1732943601
transform 1 0 1204 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_204
timestamp 1732943601
transform -1 0 1324 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_50
timestamp 1732943601
transform -1 0 1260 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_55
timestamp 1732943601
transform 1 0 1260 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1732943601
transform 1 0 1292 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_20
timestamp 1732943601
transform -1 0 1364 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1732943601
transform -1 0 1420 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_58
timestamp 1732943601
transform 1 0 1364 0 1 105
box -2 -3 26 103
use FILL  FILL_1_2_0
timestamp 1732943601
transform -1 0 1396 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1732943601
transform -1 0 1404 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_59
timestamp 1732943601
transform -1 0 1436 0 1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1732943601
transform -1 0 1428 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1732943601
transform -1 0 1436 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1732943601
transform -1 0 1532 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_38
timestamp 1732943601
transform -1 0 1484 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1732943601
transform 1 0 1484 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_162
timestamp 1732943601
transform 1 0 1532 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_206
timestamp 1732943601
transform -1 0 1588 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1732943601
transform 1 0 1588 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1732943601
transform 1 0 1580 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_12
timestamp 1732943601
transform -1 0 1644 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1732943601
transform -1 0 1740 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_61
timestamp 1732943601
transform 1 0 1676 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_62
timestamp 1732943601
transform -1 0 1732 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1732943601
transform 1 0 1740 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1732943601
transform 1 0 1764 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_155
timestamp 1732943601
transform -1 0 1812 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_1
timestamp 1732943601
transform 1 0 1812 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1732943601
transform 1 0 1732 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_3
timestamp 1732943601
transform 1 0 1844 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1732943601
transform 1 0 1868 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1732943601
transform 1 0 1900 0 -1 105
box -2 -3 26 103
use INVX4  INVX4_5
timestamp 1732943601
transform -1 0 1852 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_11
timestamp 1732943601
transform 1 0 1852 0 1 105
box -2 -3 26 103
use INVX4  INVX4_6
timestamp 1732943601
transform -1 0 1900 0 1 105
box -2 -3 26 103
use FILL  FILL_1_3_0
timestamp 1732943601
transform -1 0 1908 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1732943601
transform -1 0 1916 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1732943601
transform -1 0 2012 0 1 105
box -2 -3 98 103
use FILL  FILL_0_3_0
timestamp 1732943601
transform 1 0 1924 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1732943601
transform 1 0 1932 0 -1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_5
timestamp 1732943601
transform 1 0 1940 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1732943601
transform 1 0 1972 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1732943601
transform 1 0 1996 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_50
timestamp 1732943601
transform 1 0 2012 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1732943601
transform -1 0 2188 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_163
timestamp 1732943601
transform 1 0 2060 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_207
timestamp 1732943601
transform -1 0 2116 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1732943601
transform 1 0 2116 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1732943601
transform -1 0 2212 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1732943601
transform -1 0 2308 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_13
timestamp 1732943601
transform -1 0 2172 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_2
timestamp 1732943601
transform 1 0 2172 0 1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_21
timestamp 1732943601
transform 1 0 2244 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_22
timestamp 1732943601
transform -1 0 2300 0 1 105
box -2 -3 34 103
use FILL  FILL_2_1
timestamp 1732943601
transform 1 0 2300 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_40
timestamp 1732943601
transform -1 0 36 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1732943601
transform -1 0 132 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1732943601
transform -1 0 228 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_56
timestamp 1732943601
transform 1 0 228 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_34
timestamp 1732943601
transform 1 0 244 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_35
timestamp 1732943601
transform -1 0 300 0 -1 305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_14
timestamp 1732943601
transform -1 0 372 0 -1 305
box -2 -3 74 103
use FILL  FILL_2_0_0
timestamp 1732943601
transform -1 0 380 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1732943601
transform -1 0 388 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1732943601
transform -1 0 484 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_32
timestamp 1732943601
transform 1 0 484 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1732943601
transform 1 0 516 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_209
timestamp 1732943601
transform 1 0 540 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_267
timestamp 1732943601
transform -1 0 596 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1732943601
transform 1 0 596 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1732943601
transform -1 0 788 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_59
timestamp 1732943601
transform 1 0 788 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_60
timestamp 1732943601
transform -1 0 844 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1732943601
transform -1 0 852 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1732943601
transform -1 0 860 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1732943601
transform -1 0 956 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_166
timestamp 1732943601
transform 1 0 956 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_185
timestamp 1732943601
transform 1 0 980 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_157
timestamp 1732943601
transform -1 0 1028 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_77
timestamp 1732943601
transform 1 0 1028 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1732943601
transform 1 0 1060 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1732943601
transform -1 0 1252 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_110
timestamp 1732943601
transform -1 0 1276 0 -1 305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_7
timestamp 1732943601
transform 1 0 1276 0 -1 305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_9
timestamp 1732943601
transform 1 0 1348 0 -1 305
box -2 -3 74 103
use FILL  FILL_2_2_0
timestamp 1732943601
transform 1 0 1420 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1732943601
transform 1 0 1428 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_52
timestamp 1732943601
transform 1 0 1436 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_53
timestamp 1732943601
transform -1 0 1492 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1732943601
transform -1 0 1588 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_214
timestamp 1732943601
transform 1 0 1588 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_246
timestamp 1732943601
transform 1 0 1620 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_188
timestamp 1732943601
transform -1 0 1676 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1732943601
transform -1 0 1772 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1732943601
transform -1 0 1868 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_3_0
timestamp 1732943601
transform 1 0 1868 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1732943601
transform 1 0 1876 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1732943601
transform 1 0 1884 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_53
timestamp 1732943601
transform -1 0 2004 0 -1 305
box -2 -3 26 103
use BUFX4  BUFX4_21
timestamp 1732943601
transform 1 0 2004 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1732943601
transform 1 0 2036 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1732943601
transform -1 0 2092 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1732943601
transform -1 0 2188 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_205
timestamp 1732943601
transform -1 0 2212 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1732943601
transform -1 0 2308 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_39
timestamp 1732943601
transform -1 0 28 0 1 305
box -2 -3 26 103
use INVX1  INVX1_51
timestamp 1732943601
transform 1 0 28 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_226
timestamp 1732943601
transform 1 0 44 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_182
timestamp 1732943601
transform -1 0 100 0 1 305
box -2 -3 26 103
use INVX1  INVX1_52
timestamp 1732943601
transform 1 0 100 0 1 305
box -2 -3 18 103
use OAI22X1  OAI22X1_12
timestamp 1732943601
transform -1 0 156 0 1 305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1732943601
transform 1 0 156 0 1 305
box -2 -3 98 103
use INVX1  INVX1_20
timestamp 1732943601
transform 1 0 252 0 1 305
box -2 -3 18 103
use OAI22X1  OAI22X1_14
timestamp 1732943601
transform -1 0 308 0 1 305
box -2 -3 42 103
use INVX1  INVX1_55
timestamp 1732943601
transform -1 0 324 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1732943601
transform 1 0 324 0 1 305
box -2 -3 98 103
use FILL  FILL_3_0_0
timestamp 1732943601
transform -1 0 428 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1732943601
transform -1 0 436 0 1 305
box -2 -3 10 103
use INVX1  INVX1_30
timestamp 1732943601
transform -1 0 452 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_170
timestamp 1732943601
transform 1 0 452 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_213
timestamp 1732943601
transform -1 0 508 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1732943601
transform 1 0 508 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_76
timestamp 1732943601
transform -1 0 588 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_201
timestamp 1732943601
transform 1 0 588 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_52
timestamp 1732943601
transform 1 0 612 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1732943601
transform -1 0 668 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_29
timestamp 1732943601
transform -1 0 716 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_194
timestamp 1732943601
transform 1 0 716 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_149
timestamp 1732943601
transform 1 0 748 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_254
timestamp 1732943601
transform 1 0 772 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_196
timestamp 1732943601
transform -1 0 828 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_23
timestamp 1732943601
transform -1 0 876 0 1 305
box -2 -3 50 103
use FILL  FILL_3_1_0
timestamp 1732943601
transform -1 0 884 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1732943601
transform -1 0 892 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1732943601
transform -1 0 988 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_36
timestamp 1732943601
transform 1 0 988 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1732943601
transform -1 0 1044 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_76
timestamp 1732943601
transform -1 0 1068 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_22
timestamp 1732943601
transform 1 0 1068 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_18
timestamp 1732943601
transform 1 0 1116 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_19
timestamp 1732943601
transform -1 0 1172 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_156
timestamp 1732943601
transform 1 0 1172 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_21
timestamp 1732943601
transform -1 0 1252 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_39
timestamp 1732943601
transform 1 0 1252 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_40
timestamp 1732943601
transform 1 0 1300 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_2
timestamp 1732943601
transform 1 0 1348 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_3
timestamp 1732943601
transform -1 0 1404 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1732943601
transform -1 0 1412 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1732943601
transform -1 0 1420 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1732943601
transform -1 0 1516 0 1 305
box -2 -3 98 103
use OAI22X1  OAI22X1_11
timestamp 1732943601
transform 1 0 1516 0 1 305
box -2 -3 42 103
use MUX2X1  MUX2X1_37
timestamp 1732943601
transform -1 0 1604 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_171
timestamp 1732943601
transform 1 0 1604 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_179
timestamp 1732943601
transform 1 0 1628 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_223
timestamp 1732943601
transform 1 0 1652 0 1 305
box -2 -3 34 103
use INVX1  INVX1_44
timestamp 1732943601
transform -1 0 1700 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_16
timestamp 1732943601
transform -1 0 1732 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_172
timestamp 1732943601
transform 1 0 1732 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_215
timestamp 1732943601
transform -1 0 1788 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_51
timestamp 1732943601
transform 1 0 1788 0 1 305
box -2 -3 50 103
use INVX1  INVX1_43
timestamp 1732943601
transform -1 0 1852 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1732943601
transform -1 0 1948 0 1 305
box -2 -3 98 103
use FILL  FILL_3_3_0
timestamp 1732943601
transform 1 0 1948 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1732943601
transform 1 0 1956 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_54
timestamp 1732943601
transform 1 0 1964 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1732943601
transform 1 0 1996 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1732943601
transform -1 0 2052 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1732943601
transform -1 0 2148 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_20
timestamp 1732943601
transform 1 0 2148 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1732943601
transform -1 0 2204 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1732943601
transform -1 0 2300 0 1 305
box -2 -3 98 103
use FILL  FILL_4_1
timestamp 1732943601
transform 1 0 2300 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1732943601
transform 1 0 4 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_66
timestamp 1732943601
transform 1 0 100 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1732943601
transform -1 0 156 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1732943601
transform 1 0 156 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1732943601
transform 1 0 180 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_42
timestamp 1732943601
transform 1 0 276 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1732943601
transform -1 0 332 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_115
timestamp 1732943601
transform 1 0 332 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1732943601
transform 1 0 356 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1732943601
transform 1 0 364 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1732943601
transform 1 0 372 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_72
timestamp 1732943601
transform 1 0 468 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_71
timestamp 1732943601
transform -1 0 524 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1732943601
transform -1 0 620 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_259
timestamp 1732943601
transform -1 0 652 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1732943601
transform 1 0 652 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_64
timestamp 1732943601
transform -1 0 780 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_251
timestamp 1732943601
transform 1 0 780 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_193
timestamp 1732943601
transform -1 0 836 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1732943601
transform -1 0 932 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_1_0
timestamp 1732943601
transform 1 0 932 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1732943601
transform 1 0 940 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_76
timestamp 1732943601
transform 1 0 948 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1732943601
transform -1 0 1004 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1732943601
transform 1 0 1004 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_33
timestamp 1732943601
transform 1 0 1100 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_24
timestamp 1732943601
transform -1 0 1164 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_44
timestamp 1732943601
transform 1 0 1164 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_112
timestamp 1732943601
transform -1 0 1236 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1732943601
transform -1 0 1260 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1732943601
transform -1 0 1356 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_190
timestamp 1732943601
transform 1 0 1356 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_248
timestamp 1732943601
transform -1 0 1412 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1732943601
transform 1 0 1412 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1732943601
transform 1 0 1420 0 -1 505
box -2 -3 10 103
use INVX4  INVX4_4
timestamp 1732943601
transform 1 0 1428 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_129
timestamp 1732943601
transform -1 0 1476 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1732943601
transform 1 0 1476 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1732943601
transform 1 0 1508 0 -1 505
box -2 -3 98 103
use BUFX2  BUFX2_8
timestamp 1732943601
transform 1 0 1604 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1732943601
transform 1 0 1628 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1732943601
transform -1 0 1684 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1732943601
transform -1 0 1780 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_18
timestamp 1732943601
transform -1 0 1812 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_52
timestamp 1732943601
transform 1 0 1812 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1732943601
transform -1 0 1956 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_3_0
timestamp 1732943601
transform 1 0 1956 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1732943601
transform 1 0 1964 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_15
timestamp 1732943601
transform 1 0 1972 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_17
timestamp 1732943601
transform -1 0 2036 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_31
timestamp 1732943601
transform -1 0 2084 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_197
timestamp 1732943601
transform 1 0 2084 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_255
timestamp 1732943601
transform -1 0 2140 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_77
timestamp 1732943601
transform 1 0 2140 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_263
timestamp 1732943601
transform 1 0 2164 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1732943601
transform -1 0 2292 0 -1 505
box -2 -3 98 103
use FILL  FILL_5_1
timestamp 1732943601
transform -1 0 2300 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1732943601
transform -1 0 2308 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_30
timestamp 1732943601
transform 1 0 4 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1732943601
transform 1 0 36 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_177
timestamp 1732943601
transform 1 0 132 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1732943601
transform 1 0 156 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1732943601
transform -1 0 212 0 1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_1
timestamp 1732943601
transform 1 0 212 0 1 505
box -2 -3 74 103
use NAND2X1  NAND2X1_124
timestamp 1732943601
transform 1 0 284 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_161
timestamp 1732943601
transform 1 0 308 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1732943601
transform 1 0 340 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1732943601
transform 1 0 348 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1732943601
transform 1 0 356 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_270
timestamp 1732943601
transform 1 0 452 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_212
timestamp 1732943601
transform -1 0 508 0 1 505
box -2 -3 26 103
use INVX1  INVX1_50
timestamp 1732943601
transform 1 0 508 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_198
timestamp 1732943601
transform 1 0 524 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_197
timestamp 1732943601
transform 1 0 556 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_271
timestamp 1732943601
transform 1 0 588 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1732943601
transform 1 0 620 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_28
timestamp 1732943601
transform 1 0 716 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_63
timestamp 1732943601
transform 1 0 748 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_73
timestamp 1732943601
transform 1 0 772 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_74
timestamp 1732943601
transform -1 0 868 0 1 505
box -2 -3 50 103
use FILL  FILL_5_1_0
timestamp 1732943601
transform 1 0 868 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1732943601
transform 1 0 876 0 1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_30
timestamp 1732943601
transform 1 0 884 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1732943601
transform 1 0 932 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_28
timestamp 1732943601
transform -1 0 1052 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_126
timestamp 1732943601
transform -1 0 1076 0 1 505
box -2 -3 26 103
use INVX1  INVX1_26
timestamp 1732943601
transform 1 0 1076 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_173
timestamp 1732943601
transform -1 0 1124 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1732943601
transform 1 0 1124 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_46
timestamp 1732943601
transform 1 0 1156 0 1 505
box -2 -3 50 103
use NAND3X1  NAND3X1_13
timestamp 1732943601
transform -1 0 1236 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1732943601
transform -1 0 1260 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_56
timestamp 1732943601
transform 1 0 1260 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1732943601
transform 1 0 1292 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_132
timestamp 1732943601
transform 1 0 1324 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_49
timestamp 1732943601
transform 1 0 1348 0 1 505
box -2 -3 50 103
use FILL  FILL_5_2_0
timestamp 1732943601
transform -1 0 1404 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1732943601
transform -1 0 1412 0 1 505
box -2 -3 10 103
use INVX1  INVX1_34
timestamp 1732943601
transform -1 0 1428 0 1 505
box -2 -3 18 103
use OR2X2  OR2X2_2
timestamp 1732943601
transform -1 0 1460 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1732943601
transform -1 0 1492 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1732943601
transform -1 0 1516 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1732943601
transform 1 0 1516 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_68
timestamp 1732943601
transform 1 0 1612 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1732943601
transform -1 0 1668 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1732943601
transform 1 0 1668 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1732943601
transform 1 0 1716 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_22
timestamp 1732943601
transform -1 0 1844 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_5
timestamp 1732943601
transform 1 0 1844 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_194
timestamp 1732943601
transform 1 0 1892 0 1 505
box -2 -3 26 103
use FILL  FILL_5_3_0
timestamp 1732943601
transform -1 0 1924 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1732943601
transform -1 0 1932 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_252
timestamp 1732943601
transform -1 0 1964 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1732943601
transform 1 0 1964 0 1 505
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1732943601
transform -1 0 2012 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_33
timestamp 1732943601
transform 1 0 2012 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_32
timestamp 1732943601
transform 1 0 2060 0 1 505
box -2 -3 50 103
use BUFX4  BUFX4_69
timestamp 1732943601
transform -1 0 2140 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_78
timestamp 1732943601
transform 1 0 2140 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1732943601
transform -1 0 2268 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_70
timestamp 1732943601
transform 1 0 2268 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1732943601
transform 1 0 2300 0 1 505
box -2 -3 10 103
use INVX8  INVX8_6
timestamp 1732943601
transform 1 0 4 0 -1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1732943601
transform 1 0 44 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_221
timestamp 1732943601
transform -1 0 172 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1732943601
transform 1 0 172 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_159
timestamp 1732943601
transform 1 0 188 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1732943601
transform 1 0 220 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_160
timestamp 1732943601
transform 1 0 316 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1732943601
transform -1 0 380 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1732943601
transform -1 0 388 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1732943601
transform -1 0 396 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_170
timestamp 1732943601
transform -1 0 428 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1732943601
transform 1 0 428 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_116
timestamp 1732943601
transform 1 0 460 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_108
timestamp 1732943601
transform 1 0 484 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1732943601
transform 1 0 508 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_213
timestamp 1732943601
transform -1 0 628 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_153
timestamp 1732943601
transform 1 0 628 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_117
timestamp 1732943601
transform 1 0 652 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_45
timestamp 1732943601
transform 1 0 676 0 -1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_205
timestamp 1732943601
transform 1 0 724 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1732943601
transform -1 0 780 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1732943601
transform 1 0 780 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_1_0
timestamp 1732943601
transform -1 0 884 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1732943601
transform -1 0 892 0 -1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_28
timestamp 1732943601
transform -1 0 940 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_150
timestamp 1732943601
transform -1 0 964 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_195
timestamp 1732943601
transform -1 0 996 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_25
timestamp 1732943601
transform 1 0 996 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1732943601
transform -1 0 1060 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_196
timestamp 1732943601
transform 1 0 1060 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1732943601
transform -1 0 1116 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_119
timestamp 1732943601
transform 1 0 1116 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_189
timestamp 1732943601
transform 1 0 1140 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_247
timestamp 1732943601
transform -1 0 1196 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1732943601
transform 1 0 1196 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1732943601
transform 1 0 1228 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_158
timestamp 1732943601
transform 1 0 1260 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1732943601
transform -1 0 1388 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_2_0
timestamp 1732943601
transform 1 0 1388 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1732943601
transform 1 0 1396 0 -1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_18
timestamp 1732943601
transform 1 0 1404 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1732943601
transform 1 0 1436 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_177
timestamp 1732943601
transform 1 0 1468 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_48
timestamp 1732943601
transform 1 0 1500 0 -1 705
box -2 -3 50 103
use AOI21X1  AOI21X1_26
timestamp 1732943601
transform 1 0 1548 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1732943601
transform 1 0 1580 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1732943601
transform 1 0 1612 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_200
timestamp 1732943601
transform -1 0 1676 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1732943601
transform 1 0 1676 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_163
timestamp 1732943601
transform -1 0 1740 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1732943601
transform 1 0 1740 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_136
timestamp 1732943601
transform -1 0 1860 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_121
timestamp 1732943601
transform 1 0 1860 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_19
timestamp 1732943601
transform 1 0 1884 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_3_0
timestamp 1732943601
transform -1 0 1924 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1732943601
transform -1 0 1932 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1732943601
transform -1 0 2028 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_260
timestamp 1732943601
transform 1 0 2028 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_202
timestamp 1732943601
transform 1 0 2060 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_6
timestamp 1732943601
transform -1 0 2116 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1732943601
transform -1 0 2212 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1732943601
transform 1 0 2212 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1732943601
transform 1 0 4 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_28
timestamp 1732943601
transform 1 0 100 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1732943601
transform -1 0 156 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_219
timestamp 1732943601
transform 1 0 156 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1732943601
transform -1 0 212 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1732943601
transform 1 0 212 0 1 705
box -2 -3 98 103
use OAI22X1  OAI22X1_5
timestamp 1732943601
transform -1 0 348 0 1 705
box -2 -3 42 103
use INVX1  INVX1_21
timestamp 1732943601
transform -1 0 364 0 1 705
box -2 -3 18 103
use INVX1  INVX1_31
timestamp 1732943601
transform 1 0 364 0 1 705
box -2 -3 18 103
use FILL  FILL_7_0_0
timestamp 1732943601
transform -1 0 388 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1732943601
transform -1 0 396 0 1 705
box -2 -3 10 103
use OAI22X1  OAI22X1_8
timestamp 1732943601
transform -1 0 436 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_171
timestamp 1732943601
transform 1 0 436 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1732943601
transform 1 0 468 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1732943601
transform 1 0 500 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_133
timestamp 1732943601
transform -1 0 564 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_86
timestamp 1732943601
transform -1 0 588 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_155
timestamp 1732943601
transform 1 0 588 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_199
timestamp 1732943601
transform -1 0 652 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_272
timestamp 1732943601
transform 1 0 652 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_214
timestamp 1732943601
transform -1 0 708 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1732943601
transform -1 0 804 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_9
timestamp 1732943601
transform 1 0 804 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_12
timestamp 1732943601
transform 1 0 828 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1732943601
transform -1 0 884 0 1 705
box -2 -3 26 103
use FILL  FILL_7_1_0
timestamp 1732943601
transform -1 0 892 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1732943601
transform -1 0 900 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1732943601
transform -1 0 996 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_77
timestamp 1732943601
transform 1 0 996 0 1 705
box -2 -3 50 103
use NAND3X1  NAND3X1_21
timestamp 1732943601
transform 1 0 1044 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_151
timestamp 1732943601
transform -1 0 1100 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_165
timestamp 1732943601
transform 1 0 1100 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1732943601
transform 1 0 1132 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_53
timestamp 1732943601
transform -1 0 1196 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_109
timestamp 1732943601
transform 1 0 1196 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_54
timestamp 1732943601
transform -1 0 1252 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1732943601
transform 1 0 1252 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_256
timestamp 1732943601
transform 1 0 1348 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_198
timestamp 1732943601
transform -1 0 1404 0 1 705
box -2 -3 26 103
use FILL  FILL_7_2_0
timestamp 1732943601
transform 1 0 1404 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1732943601
transform 1 0 1412 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_264
timestamp 1732943601
transform 1 0 1420 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_206
timestamp 1732943601
transform -1 0 1476 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1732943601
transform 1 0 1476 0 1 705
box -2 -3 98 103
use INVX8  INVX8_11
timestamp 1732943601
transform -1 0 1612 0 1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1732943601
transform 1 0 1612 0 1 705
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1732943601
transform 1 0 1708 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_180
timestamp 1732943601
transform -1 0 1764 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1732943601
transform 1 0 1764 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1732943601
transform -1 0 1828 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_137
timestamp 1732943601
transform 1 0 1828 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_6
timestamp 1732943601
transform 1 0 1852 0 1 705
box -2 -3 50 103
use FILL  FILL_7_3_0
timestamp 1732943601
transform -1 0 1908 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1732943601
transform -1 0 1916 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_179
timestamp 1732943601
transform -1 0 1948 0 1 705
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1732943601
transform -1 0 1964 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_55
timestamp 1732943601
transform -1 0 2012 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_53
timestamp 1732943601
transform -1 0 2060 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1732943601
transform -1 0 2156 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_87
timestamp 1732943601
transform 1 0 2156 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1732943601
transform -1 0 2212 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_11
timestamp 1732943601
transform 1 0 2212 0 1 705
box -2 -3 74 103
use BUFX2  BUFX2_3
timestamp 1732943601
transform 1 0 2284 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1732943601
transform 1 0 4 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_122
timestamp 1732943601
transform -1 0 132 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1732943601
transform -1 0 164 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1732943601
transform 1 0 164 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1732943601
transform -1 0 228 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1732943601
transform 1 0 228 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_113
timestamp 1732943601
transform 1 0 260 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1732943601
transform 1 0 292 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_0_0
timestamp 1732943601
transform 1 0 388 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1732943601
transform 1 0 396 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_125
timestamp 1732943601
transform 1 0 404 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1732943601
transform 1 0 428 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_131
timestamp 1732943601
transform 1 0 524 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1732943601
transform -1 0 580 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1732943601
transform 1 0 580 0 -1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_13
timestamp 1732943601
transform 1 0 596 0 -1 905
box -2 -3 42 103
use INVX1  INVX1_53
timestamp 1732943601
transform -1 0 652 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_164
timestamp 1732943601
transform 1 0 652 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_5
timestamp 1732943601
transform -1 0 756 0 -1 905
box -2 -3 74 103
use NAND3X1  NAND3X1_22
timestamp 1732943601
transform 1 0 756 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1732943601
transform -1 0 884 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_1_0
timestamp 1732943601
transform 1 0 884 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1732943601
transform 1 0 892 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_56
timestamp 1732943601
transform 1 0 900 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1732943601
transform 1 0 932 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_24
timestamp 1732943601
transform 1 0 956 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1732943601
transform 1 0 988 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_166
timestamp 1732943601
transform 1 0 1084 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1732943601
transform 1 0 1116 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_167
timestamp 1732943601
transform 1 0 1148 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1732943601
transform 1 0 1180 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1732943601
transform 1 0 1212 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1732943601
transform -1 0 1404 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_2_0
timestamp 1732943601
transform 1 0 1404 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1732943601
transform 1 0 1412 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_72
timestamp 1732943601
transform 1 0 1420 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_73
timestamp 1732943601
transform -1 0 1476 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_191
timestamp 1732943601
transform -1 0 1500 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_135
timestamp 1732943601
transform -1 0 1524 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_7
timestamp 1732943601
transform 1 0 1524 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_16
timestamp 1732943601
transform 1 0 1556 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_17
timestamp 1732943601
transform 1 0 1588 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_8
timestamp 1732943601
transform 1 0 1620 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1732943601
transform -1 0 1684 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1732943601
transform -1 0 1716 0 -1 905
box -2 -3 34 103
use BUFX2  BUFX2_4
timestamp 1732943601
transform 1 0 1716 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_181
timestamp 1732943601
transform -1 0 1772 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_20
timestamp 1732943601
transform -1 0 1804 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_182
timestamp 1732943601
transform 1 0 1804 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_134
timestamp 1732943601
transform -1 0 1860 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_4
timestamp 1732943601
transform -1 0 1908 0 -1 905
box -2 -3 50 103
use FILL  FILL_8_3_0
timestamp 1732943601
transform 1 0 1908 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1732943601
transform 1 0 1916 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_17
timestamp 1732943601
transform 1 0 1924 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1732943601
transform -1 0 1980 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1732943601
transform -1 0 2076 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_54
timestamp 1732943601
transform 1 0 2076 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1732943601
transform -1 0 2220 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_207
timestamp 1732943601
transform 1 0 2220 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_265
timestamp 1732943601
transform -1 0 2276 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1732943601
transform 1 0 2276 0 -1 905
box -2 -3 26 103
use FILL  FILL_9_1
timestamp 1732943601
transform -1 0 2308 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1732943601
transform -1 0 100 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_178
timestamp 1732943601
transform 1 0 100 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_222
timestamp 1732943601
transform -1 0 156 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1732943601
transform 1 0 156 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_64
timestamp 1732943601
transform -1 0 212 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1732943601
transform 1 0 212 0 1 905
box -2 -3 98 103
use INVX1  INVX1_35
timestamp 1732943601
transform 1 0 308 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_96
timestamp 1732943601
transform 1 0 324 0 1 905
box -2 -3 26 103
use INVX1  INVX1_3
timestamp 1732943601
transform 1 0 348 0 1 905
box -2 -3 18 103
use FILL  FILL_9_0_0
timestamp 1732943601
transform 1 0 364 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1732943601
transform 1 0 372 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_141
timestamp 1732943601
transform 1 0 380 0 1 905
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1732943601
transform 1 0 412 0 1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_1
timestamp 1732943601
transform 1 0 428 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_142
timestamp 1732943601
transform 1 0 468 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_98
timestamp 1732943601
transform 1 0 500 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_128
timestamp 1732943601
transform -1 0 548 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_175
timestamp 1732943601
transform 1 0 548 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1732943601
transform 1 0 580 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_47
timestamp 1732943601
transform 1 0 676 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_48
timestamp 1732943601
transform -1 0 732 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1732943601
transform -1 0 764 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_128
timestamp 1732943601
transform 1 0 764 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1732943601
transform -1 0 892 0 1 905
box -2 -3 98 103
use FILL  FILL_9_1_0
timestamp 1732943601
transform 1 0 892 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1732943601
transform 1 0 900 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_55
timestamp 1732943601
transform 1 0 908 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_18
timestamp 1732943601
transform -1 0 964 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_183
timestamp 1732943601
transform -1 0 988 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_148
timestamp 1732943601
transform 1 0 988 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_218
timestamp 1732943601
transform -1 0 1044 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1732943601
transform -1 0 1068 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_152
timestamp 1732943601
transform -1 0 1092 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_75
timestamp 1732943601
transform -1 0 1140 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_122
timestamp 1732943601
transform -1 0 1164 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_10
timestamp 1732943601
transform -1 0 1196 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_34
timestamp 1732943601
transform -1 0 1228 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1732943601
transform -1 0 1252 0 1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_1
timestamp 1732943601
transform -1 0 1292 0 1 905
box -2 -3 42 103
use INVX1  INVX1_2
timestamp 1732943601
transform -1 0 1308 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_127
timestamp 1732943601
transform -1 0 1332 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_174
timestamp 1732943601
transform -1 0 1364 0 1 905
box -2 -3 34 103
use FILL  FILL_9_2_0
timestamp 1732943601
transform 1 0 1364 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1732943601
transform 1 0 1372 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1732943601
transform 1 0 1380 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_249
timestamp 1732943601
transform -1 0 1508 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_185
timestamp 1732943601
transform -1 0 1540 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1732943601
transform -1 0 1572 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1732943601
transform 1 0 1572 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1732943601
transform 1 0 1604 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1732943601
transform 1 0 1700 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_1
timestamp 1732943601
transform 1 0 1796 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1732943601
transform -1 0 1852 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_12
timestamp 1732943601
transform -1 0 1884 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_133
timestamp 1732943601
transform 1 0 1884 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1732943601
transform 1 0 1908 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1732943601
transform 1 0 1916 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_22
timestamp 1732943601
transform 1 0 1924 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_186
timestamp 1732943601
transform -1 0 1988 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_19
timestamp 1732943601
transform 1 0 1988 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1732943601
transform -1 0 2052 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1732943601
transform 1 0 2052 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1732943601
transform 1 0 2148 0 1 905
box -2 -3 98 103
use BUFX2  BUFX2_5
timestamp 1732943601
transform 1 0 2244 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1732943601
transform 1 0 2268 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1732943601
transform 1 0 2292 0 1 905
box -2 -3 10 103
use FILL  FILL_10_2
timestamp 1732943601
transform 1 0 2300 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_67
timestamp 1732943601
transform -1 0 28 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1732943601
transform 1 0 28 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_123
timestamp 1732943601
transform 1 0 44 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_168
timestamp 1732943601
transform -1 0 100 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1732943601
transform 1 0 100 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_33
timestamp 1732943601
transform 1 0 196 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1732943601
transform -1 0 252 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_169
timestamp 1732943601
transform 1 0 252 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1732943601
transform -1 0 316 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1732943601
transform 1 0 316 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_0_0
timestamp 1732943601
transform 1 0 332 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1732943601
transform 1 0 340 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1732943601
transform 1 0 348 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_42
timestamp 1732943601
transform 1 0 444 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1732943601
transform 1 0 476 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_54
timestamp 1732943601
transform 1 0 572 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_217
timestamp 1732943601
transform 1 0 588 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_275
timestamp 1732943601
transform -1 0 644 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1732943601
transform 1 0 644 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_7
timestamp 1732943601
transform 1 0 740 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_127
timestamp 1732943601
transform 1 0 772 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_123
timestamp 1732943601
transform 1 0 804 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1732943601
transform -1 0 868 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1732943601
transform 1 0 868 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1732943601
transform 1 0 876 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1732943601
transform 1 0 884 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_8
timestamp 1732943601
transform 1 0 980 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1732943601
transform -1 0 1036 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1732943601
transform 1 0 1036 0 -1 1105
box -2 -3 98 103
use INVX4  INVX4_10
timestamp 1732943601
transform 1 0 1132 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1732943601
transform -1 0 1180 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_33
timestamp 1732943601
transform -1 0 1212 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_11
timestamp 1732943601
transform 1 0 1212 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_138
timestamp 1732943601
transform -1 0 1276 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1732943601
transform 1 0 1276 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_70
timestamp 1732943601
transform 1 0 1372 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_2_0
timestamp 1732943601
transform -1 0 1412 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1732943601
transform -1 0 1420 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_69
timestamp 1732943601
transform -1 0 1444 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_38
timestamp 1732943601
transform 1 0 1444 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_183
timestamp 1732943601
transform -1 0 1492 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_184
timestamp 1732943601
transform 1 0 1492 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1732943601
transform 1 0 1524 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1732943601
transform -1 0 1572 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_139
timestamp 1732943601
transform -1 0 1604 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1732943601
transform 1 0 1604 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1732943601
transform -1 0 1668 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1732943601
transform -1 0 1684 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1732943601
transform -1 0 1780 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_82
timestamp 1732943601
transform 1 0 1780 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_129
timestamp 1732943601
transform -1 0 1836 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1732943601
transform 1 0 1836 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_273
timestamp 1732943601
transform 1 0 1860 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_215
timestamp 1732943601
transform -1 0 1916 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_3_0
timestamp 1732943601
transform -1 0 1924 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1732943601
transform -1 0 1932 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1732943601
transform -1 0 2028 0 -1 1105
box -2 -3 98 103
use INVX8  INVX8_1
timestamp 1732943601
transform 1 0 2028 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_258
timestamp 1732943601
transform 1 0 2068 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1732943601
transform -1 0 2196 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1732943601
transform 1 0 2196 0 -1 1105
box -2 -3 98 103
use FILL  FILL_11_1
timestamp 1732943601
transform -1 0 2300 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1732943601
transform -1 0 2308 0 -1 1105
box -2 -3 10 103
use INVX8  INVX8_2
timestamp 1732943601
transform 1 0 4 0 1 1105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1732943601
transform 1 0 44 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_120
timestamp 1732943601
transform 1 0 140 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1732943601
transform -1 0 204 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_29
timestamp 1732943601
transform 1 0 204 0 1 1105
box -2 -3 18 103
use OAI22X1  OAI22X1_7
timestamp 1732943601
transform -1 0 260 0 1 1105
box -2 -3 42 103
use OAI22X1  OAI22X1_6
timestamp 1732943601
transform -1 0 300 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_24
timestamp 1732943601
transform -1 0 316 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_46
timestamp 1732943601
transform -1 0 348 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_301
timestamp 1732943601
transform 1 0 348 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1732943601
transform 1 0 380 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1732943601
transform 1 0 388 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_300
timestamp 1732943601
transform 1 0 396 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_1
timestamp 1732943601
transform 1 0 428 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_306
timestamp 1732943601
transform 1 0 460 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_307
timestamp 1732943601
transform -1 0 524 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1732943601
transform -1 0 620 0 1 1105
box -2 -3 98 103
use OR2X2  OR2X2_1
timestamp 1732943601
transform -1 0 652 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1732943601
transform 1 0 652 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_116
timestamp 1732943601
transform 1 0 684 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1732943601
transform -1 0 748 0 1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1732943601
transform 1 0 748 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_41
timestamp 1732943601
transform -1 0 804 0 1 1105
box -2 -3 18 103
use INVX4  INVX4_9
timestamp 1732943601
transform 1 0 804 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1732943601
transform -1 0 924 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_1_0
timestamp 1732943601
transform 1 0 924 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1732943601
transform 1 0 932 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_45
timestamp 1732943601
transform 1 0 940 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_46
timestamp 1732943601
transform -1 0 996 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1732943601
transform 1 0 996 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_90
timestamp 1732943601
transform -1 0 1044 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_34
timestamp 1732943601
transform 1 0 1044 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_33
timestamp 1732943601
transform -1 0 1100 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_12
timestamp 1732943601
transform -1 0 1116 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_113
timestamp 1732943601
transform -1 0 1140 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_16
timestamp 1732943601
transform -1 0 1164 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1732943601
transform -1 0 1196 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1732943601
transform 1 0 1196 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1732943601
transform 1 0 1220 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_130
timestamp 1732943601
transform -1 0 1276 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_38
timestamp 1732943601
transform 1 0 1276 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1732943601
transform -1 0 1404 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_2_0
timestamp 1732943601
transform 1 0 1404 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1732943601
transform 1 0 1412 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_37
timestamp 1732943601
transform 1 0 1420 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_38
timestamp 1732943601
transform -1 0 1476 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1732943601
transform 1 0 1476 0 1 1105
box -2 -3 18 103
use OAI22X1  OAI22X1_9
timestamp 1732943601
transform 1 0 1492 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_138
timestamp 1732943601
transform -1 0 1556 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_137
timestamp 1732943601
transform -1 0 1588 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_91
timestamp 1732943601
transform 1 0 1588 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_156
timestamp 1732943601
transform 1 0 1612 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_10
timestamp 1732943601
transform 1 0 1636 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_21
timestamp 1732943601
transform 1 0 1668 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_71
timestamp 1732943601
transform -1 0 1732 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1732943601
transform -1 0 1764 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_9
timestamp 1732943601
transform -1 0 1796 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_148
timestamp 1732943601
transform 1 0 1796 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_100
timestamp 1732943601
transform -1 0 1852 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1732943601
transform 1 0 1852 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1732943601
transform -1 0 1916 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_3_0
timestamp 1732943601
transform 1 0 1916 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1732943601
transform 1 0 1924 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1732943601
transform 1 0 1932 0 1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_70
timestamp 1732943601
transform -1 0 2076 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_200
timestamp 1732943601
transform 1 0 2076 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1732943601
transform -1 0 2196 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1732943601
transform 1 0 2196 0 1 1105
box -2 -3 98 103
use FILL  FILL_12_1
timestamp 1732943601
transform 1 0 2292 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1732943601
transform 1 0 2300 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_68
timestamp 1732943601
transform -1 0 36 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1732943601
transform -1 0 132 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_28
timestamp 1732943601
transform 1 0 132 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1732943601
transform 1 0 148 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_23
timestamp 1732943601
transform 1 0 244 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_297
timestamp 1732943601
transform 1 0 260 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_296
timestamp 1732943601
transform -1 0 324 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1732943601
transform 1 0 324 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_0_0
timestamp 1732943601
transform -1 0 428 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1732943601
transform -1 0 436 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_32
timestamp 1732943601
transform -1 0 452 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1732943601
transform -1 0 484 0 -1 1305
box -2 -3 34 103
use INVX4  INVX4_8
timestamp 1732943601
transform -1 0 508 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_136
timestamp 1732943601
transform 1 0 508 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1732943601
transform -1 0 564 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_48
timestamp 1732943601
transform 1 0 564 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_193
timestamp 1732943601
transform 1 0 580 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1732943601
transform -1 0 636 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_25
timestamp 1732943601
transform 1 0 636 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1732943601
transform 1 0 652 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_42
timestamp 1732943601
transform 1 0 748 0 -1 1305
box -2 -3 18 103
use INVX1  INVX1_13
timestamp 1732943601
transform 1 0 764 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_268
timestamp 1732943601
transform 1 0 780 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_210
timestamp 1732943601
transform -1 0 836 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1732943601
transform 1 0 836 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_1_0
timestamp 1732943601
transform -1 0 940 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1732943601
transform -1 0 948 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_186
timestamp 1732943601
transform -1 0 972 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_18
timestamp 1732943601
transform -1 0 996 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_31
timestamp 1732943601
transform -1 0 1028 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1732943601
transform -1 0 1060 0 -1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1732943601
transform 1 0 1060 0 -1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_9
timestamp 1732943601
transform -1 0 1132 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_3
timestamp 1732943601
transform -1 0 1164 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1732943601
transform 1 0 1164 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_4
timestamp 1732943601
transform 1 0 1188 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_64
timestamp 1732943601
transform -1 0 1252 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1732943601
transform 1 0 1252 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_66
timestamp 1732943601
transform -1 0 1380 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_105
timestamp 1732943601
transform 1 0 1380 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_2_0
timestamp 1732943601
transform -1 0 1412 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1732943601
transform -1 0 1420 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_151
timestamp 1732943601
transform -1 0 1452 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_107
timestamp 1732943601
transform 1 0 1452 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_150
timestamp 1732943601
transform -1 0 1508 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1732943601
transform -1 0 1524 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1732943601
transform -1 0 1620 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_26
timestamp 1732943601
transform -1 0 1652 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1732943601
transform -1 0 1684 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_146
timestamp 1732943601
transform 1 0 1684 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_72
timestamp 1732943601
transform -1 0 1740 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_220
timestamp 1732943601
transform 1 0 1740 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_176
timestamp 1732943601
transform -1 0 1796 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1732943601
transform -1 0 1892 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_147
timestamp 1732943601
transform -1 0 1924 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1732943601
transform 1 0 1924 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1732943601
transform 1 0 1932 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_13
timestamp 1732943601
transform 1 0 1940 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_71
timestamp 1732943601
transform 1 0 1972 0 -1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_24
timestamp 1732943601
transform 1 0 2020 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_192
timestamp 1732943601
transform -1 0 2084 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_69
timestamp 1732943601
transform 1 0 2084 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_6
timestamp 1732943601
transform 1 0 2132 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1732943601
transform -1 0 2188 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1732943601
transform -1 0 2284 0 -1 1305
box -2 -3 98 103
use BUFX2  BUFX2_2
timestamp 1732943601
transform 1 0 2284 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1732943601
transform 1 0 4 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_35
timestamp 1732943601
transform 1 0 100 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_36
timestamp 1732943601
transform -1 0 156 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1732943601
transform 1 0 156 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_293
timestamp 1732943601
transform 1 0 252 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1732943601
transform 1 0 284 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_0_0
timestamp 1732943601
transform 1 0 380 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1732943601
transform 1 0 388 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_299
timestamp 1732943601
transform 1 0 396 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_298
timestamp 1732943601
transform -1 0 460 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1732943601
transform -1 0 484 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_45
timestamp 1732943601
transform -1 0 516 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1732943601
transform 1 0 516 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_106
timestamp 1732943601
transform 1 0 612 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1732943601
transform 1 0 636 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_303
timestamp 1732943601
transform -1 0 764 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_219
timestamp 1732943601
transform -1 0 788 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_30
timestamp 1732943601
transform 1 0 788 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1732943601
transform 1 0 820 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1732943601
transform 1 0 852 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1732943601
transform 1 0 860 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1732943601
transform 1 0 868 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_20
timestamp 1732943601
transform 1 0 964 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_61
timestamp 1732943601
transform -1 0 1020 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1732943601
transform 1 0 1020 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1732943601
transform 1 0 1052 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_62
timestamp 1732943601
transform -1 0 1116 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_29
timestamp 1732943601
transform -1 0 1148 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1732943601
transform 1 0 1148 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1732943601
transform 1 0 1180 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1732943601
transform -1 0 1244 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1732943601
transform -1 0 1276 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1732943601
transform 1 0 1276 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_63
timestamp 1732943601
transform -1 0 1332 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1732943601
transform 1 0 1332 0 1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1732943601
transform 1 0 1356 0 1 1305
box -2 -3 42 103
use FILL  FILL_13_2_0
timestamp 1732943601
transform -1 0 1404 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1732943601
transform -1 0 1412 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_152
timestamp 1732943601
transform -1 0 1444 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1732943601
transform 1 0 1444 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1732943601
transform -1 0 1492 0 1 1305
box -2 -3 18 103
use INVX8  INVX8_3
timestamp 1732943601
transform -1 0 1532 0 1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_15
timestamp 1732943601
transform -1 0 1556 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_227
timestamp 1732943601
transform -1 0 1588 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1732943601
transform 1 0 1588 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_145
timestamp 1732943601
transform 1 0 1612 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_20
timestamp 1732943601
transform 1 0 1636 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_191
timestamp 1732943601
transform -1 0 1700 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_190
timestamp 1732943601
transform 1 0 1700 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_245
timestamp 1732943601
transform 1 0 1732 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1732943601
transform -1 0 1788 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_78
timestamp 1732943601
transform 1 0 1788 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_79
timestamp 1732943601
transform -1 0 1844 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_101
timestamp 1732943601
transform -1 0 1868 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_3_0
timestamp 1732943601
transform -1 0 1876 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1732943601
transform -1 0 1884 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1732943601
transform -1 0 1980 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_146
timestamp 1732943601
transform -1 0 2012 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1732943601
transform -1 0 2028 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_73
timestamp 1732943601
transform 1 0 2028 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_74
timestamp 1732943601
transform -1 0 2084 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1732943601
transform -1 0 2180 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1732943601
transform 1 0 2180 0 1 1305
box -2 -3 98 103
use BUFX2  BUFX2_7
timestamp 1732943601
transform 1 0 2276 0 1 1305
box -2 -3 26 103
use FILL  FILL_14_1
timestamp 1732943601
transform 1 0 2300 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1732943601
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_41
timestamp 1732943601
transform 1 0 100 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_40
timestamp 1732943601
transform -1 0 156 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_97
timestamp 1732943601
transform 1 0 156 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_26
timestamp 1732943601
transform -1 0 204 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_143
timestamp 1732943601
transform 1 0 204 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1732943601
transform 1 0 236 0 -1 1505
box -2 -3 18 103
use INVX1  INVX1_8
timestamp 1732943601
transform 1 0 252 0 -1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_2
timestamp 1732943601
transform 1 0 268 0 -1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_292
timestamp 1732943601
transform -1 0 340 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1732943601
transform 1 0 340 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_0_0
timestamp 1732943601
transform 1 0 372 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1732943601
transform 1 0 380 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_144
timestamp 1732943601
transform 1 0 388 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_295
timestamp 1732943601
transform -1 0 452 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_294
timestamp 1732943601
transform -1 0 484 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_65
timestamp 1732943601
transform -1 0 516 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_66
timestamp 1732943601
transform 1 0 516 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1732943601
transform 1 0 548 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_305
timestamp 1732943601
transform 1 0 644 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_304
timestamp 1732943601
transform -1 0 708 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_302
timestamp 1732943601
transform 1 0 708 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_59
timestamp 1732943601
transform 1 0 740 0 -1 1505
box -2 -3 50 103
use INVX4  INVX4_7
timestamp 1732943601
transform 1 0 788 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1732943601
transform 1 0 812 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_201
timestamp 1732943601
transform -1 0 876 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_1_0
timestamp 1732943601
transform -1 0 884 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1732943601
transform -1 0 892 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_1
timestamp 1732943601
transform -1 0 924 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1732943601
transform 1 0 924 0 -1 1505
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1732943601
transform 1 0 956 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_6
timestamp 1732943601
transform 1 0 980 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1732943601
transform -1 0 1036 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_7
timestamp 1732943601
transform 1 0 1036 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1732943601
transform -1 0 1100 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_19
timestamp 1732943601
transform 1 0 1100 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1732943601
transform -1 0 1148 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_4
timestamp 1732943601
transform -1 0 1180 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_47
timestamp 1732943601
transform 1 0 1180 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1732943601
transform -1 0 1236 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_218
timestamp 1732943601
transform -1 0 1260 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_141
timestamp 1732943601
transform -1 0 1284 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_188
timestamp 1732943601
transform 1 0 1284 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1732943601
transform 1 0 1316 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_39
timestamp 1732943601
transform -1 0 1364 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1732943601
transform -1 0 1388 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_2_0
timestamp 1732943601
transform 1 0 1388 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1732943601
transform 1 0 1396 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_250
timestamp 1732943601
transform 1 0 1404 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_192
timestamp 1732943601
transform -1 0 1460 0 -1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_2
timestamp 1732943601
transform 1 0 1460 0 -1 1505
box -2 -3 42 103
use NAND3X1  NAND3X1_19
timestamp 1732943601
transform 1 0 1500 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1732943601
transform -1 0 1548 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_66
timestamp 1732943601
transform -1 0 1596 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_68
timestamp 1732943601
transform -1 0 1644 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1732943601
transform -1 0 1740 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_224
timestamp 1732943601
transform 1 0 1740 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_180
timestamp 1732943601
transform -1 0 1796 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1732943601
transform -1 0 1892 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_18
timestamp 1732943601
transform 1 0 1892 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1732943601
transform -1 0 1932 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1732943601
transform -1 0 1940 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_17
timestamp 1732943601
transform -1 0 1964 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1732943601
transform 1 0 1964 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_9
timestamp 1732943601
transform -1 0 2076 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1732943601
transform 1 0 2076 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_2
timestamp 1732943601
transform 1 0 2172 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1732943601
transform 1 0 2204 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1732943601
transform -1 0 2308 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_25
timestamp 1732943601
transform -1 0 36 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1732943601
transform -1 0 60 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_37
timestamp 1732943601
transform 1 0 60 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1732943601
transform 1 0 92 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1732943601
transform 1 0 4 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_6
timestamp 1732943601
transform 1 0 100 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1732943601
transform 1 0 124 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_167
timestamp 1732943601
transform 1 0 116 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1732943601
transform -1 0 172 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1732943601
transform 1 0 172 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1732943601
transform 1 0 204 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1732943601
transform 1 0 220 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_85
timestamp 1732943601
transform 1 0 300 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1732943601
transform 1 0 316 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_132
timestamp 1732943601
transform -1 0 356 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_0_0
timestamp 1732943601
transform 1 0 356 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1732943601
transform 1 0 364 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1732943601
transform 1 0 372 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_0_0
timestamp 1732943601
transform 1 0 412 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1732943601
transform 1 0 420 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_126
timestamp 1732943601
transform 1 0 428 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1732943601
transform -1 0 492 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_27
timestamp 1732943601
transform -1 0 540 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_25
timestamp 1732943601
transform -1 0 516 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1732943601
transform 1 0 540 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_233
timestamp 1732943601
transform 1 0 516 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_232
timestamp 1732943601
transform -1 0 580 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_68
timestamp 1732943601
transform 1 0 580 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_71
timestamp 1732943601
transform 1 0 636 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1732943601
transform -1 0 692 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_46
timestamp 1732943601
transform 1 0 692 0 1 1505
box -2 -3 18 103
use BUFX4  BUFX4_8
timestamp 1732943601
transform -1 0 740 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_80
timestamp 1732943601
transform 1 0 612 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_78
timestamp 1732943601
transform 1 0 660 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_242
timestamp 1732943601
transform 1 0 708 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1732943601
transform 1 0 740 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_243
timestamp 1732943601
transform -1 0 772 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1732943601
transform 1 0 772 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_231
timestamp 1732943601
transform 1 0 836 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_1_0
timestamp 1732943601
transform 1 0 868 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1732943601
transform 1 0 876 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1732943601
transform 1 0 884 0 1 1505
box -2 -3 98 103
use BUFX4  BUFX4_67
timestamp 1732943601
transform 1 0 868 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_1_0
timestamp 1732943601
transform -1 0 908 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1732943601
transform -1 0 916 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_184
timestamp 1732943601
transform -1 0 1004 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_285
timestamp 1732943601
transform -1 0 1036 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1732943601
transform -1 0 948 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_16
timestamp 1732943601
transform 1 0 948 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_284
timestamp 1732943601
transform 1 0 996 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_95
timestamp 1732943601
transform -1 0 1060 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1732943601
transform 1 0 1060 0 1 1505
box -2 -3 98 103
use BUFX4  BUFX4_6
timestamp 1732943601
transform 1 0 1028 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1732943601
transform 1 0 1060 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1732943601
transform 1 0 1156 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_41
timestamp 1732943601
transform 1 0 1156 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_43
timestamp 1732943601
transform -1 0 1252 0 -1 1705
box -2 -3 50 103
use BUFX4  BUFX4_27
timestamp 1732943601
transform -1 0 1284 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1732943601
transform -1 0 1308 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1732943601
transform 1 0 1308 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_18
timestamp 1732943601
transform -1 0 1300 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_63
timestamp 1732943601
transform -1 0 1348 0 -1 1705
box -2 -3 50 103
use FILL  FILL_15_2_0
timestamp 1732943601
transform 1 0 1404 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1732943601
transform 1 0 1412 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_65
timestamp 1732943601
transform -1 0 1396 0 -1 1705
box -2 -3 50 103
use FILL  FILL_16_2_0
timestamp 1732943601
transform 1 0 1396 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1732943601
transform 1 0 1404 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1732943601
transform 1 0 1412 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_45
timestamp 1732943601
transform 1 0 1420 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_144
timestamp 1732943601
transform -1 0 1460 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_187
timestamp 1732943601
transform 1 0 1460 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_23
timestamp 1732943601
transform 1 0 1492 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1732943601
transform -1 0 1524 0 -1 1705
box -2 -3 18 103
use BUFX4  BUFX4_57
timestamp 1732943601
transform -1 0 1556 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_140
timestamp 1732943601
transform 1 0 1556 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_30
timestamp 1732943601
transform 1 0 1580 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1732943601
transform -1 0 1700 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_189
timestamp 1732943601
transform -1 0 1556 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_142
timestamp 1732943601
transform 1 0 1556 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1732943601
transform 1 0 1580 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_31
timestamp 1732943601
transform -1 0 1732 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_88
timestamp 1732943601
transform 1 0 1676 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_135
timestamp 1732943601
transform -1 0 1732 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_67
timestamp 1732943601
transform 1 0 1732 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_143
timestamp 1732943601
transform 1 0 1780 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_274
timestamp 1732943601
transform 1 0 1804 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1732943601
transform -1 0 1764 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1732943601
transform 1 0 1764 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_26
timestamp 1732943601
transform 1 0 1788 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1732943601
transform 1 0 1820 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_216
timestamp 1732943601
transform -1 0 1860 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1732943601
transform -1 0 1956 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1732943601
transform 1 0 1852 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_3_0
timestamp 1732943601
transform 1 0 1956 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1732943601
transform 1 0 1964 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_99
timestamp 1732943601
transform 1 0 1972 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_13
timestamp 1732943601
transform 1 0 1996 0 1 1505
box -2 -3 50 103
use FILL  FILL_16_3_0
timestamp 1732943601
transform 1 0 1948 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1732943601
transform 1 0 1956 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_15
timestamp 1732943601
transform 1 0 1964 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_14
timestamp 1732943601
transform 1 0 2012 0 -1 1705
box -2 -3 50 103
use BUFX4  BUFX4_60
timestamp 1732943601
transform -1 0 2076 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1732943601
transform 1 0 2076 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1732943601
transform -1 0 2132 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1732943601
transform -1 0 2156 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_130
timestamp 1732943601
transform -1 0 2164 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1732943601
transform -1 0 2260 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_203
timestamp 1732943601
transform 1 0 2156 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_261
timestamp 1732943601
transform -1 0 2212 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1732943601
transform 1 0 2212 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_23
timestamp 1732943601
transform -1 0 2292 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1
timestamp 1732943601
transform 1 0 2292 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1732943601
transform 1 0 2300 0 1 1505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_10
timestamp 1732943601
transform 1 0 2236 0 -1 1705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_3
timestamp 1732943601
transform 1 0 4 0 1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1732943601
transform -1 0 172 0 1 1705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_8
timestamp 1732943601
transform 1 0 172 0 1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1732943601
transform 1 0 244 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_86
timestamp 1732943601
transform -1 0 372 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_0_0
timestamp 1732943601
transform -1 0 380 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1732943601
transform -1 0 388 0 1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_26
timestamp 1732943601
transform -1 0 436 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1732943601
transform 1 0 436 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_235
timestamp 1732943601
transform 1 0 532 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_234
timestamp 1732943601
transform -1 0 596 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_34
timestamp 1732943601
transform 1 0 596 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_8
timestamp 1732943601
transform -1 0 692 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_9
timestamp 1732943601
transform 1 0 692 0 1 1705
box -2 -3 50 103
use BUFX4  BUFX4_36
timestamp 1732943601
transform 1 0 740 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1732943601
transform 1 0 772 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_279
timestamp 1732943601
transform 1 0 868 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_1_0
timestamp 1732943601
transform -1 0 908 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1732943601
transform -1 0 916 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_278
timestamp 1732943601
transform -1 0 948 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_12
timestamp 1732943601
transform -1 0 988 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_81
timestamp 1732943601
transform 1 0 988 0 1 1705
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1732943601
transform 1 0 1012 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_240
timestamp 1732943601
transform 1 0 1036 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_241
timestamp 1732943601
transform -1 0 1100 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1732943601
transform 1 0 1100 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1732943601
transform 1 0 1132 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1732943601
transform 1 0 1164 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_42
timestamp 1732943601
transform -1 0 1308 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_80
timestamp 1732943601
transform -1 0 1332 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_17
timestamp 1732943601
transform -1 0 1380 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_84
timestamp 1732943601
transform 1 0 1380 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_2_0
timestamp 1732943601
transform -1 0 1420 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1732943601
transform -1 0 1428 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1732943601
transform -1 0 1524 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_58
timestamp 1732943601
transform 1 0 1524 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1732943601
transform -1 0 1580 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_50
timestamp 1732943601
transform 1 0 1580 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_49
timestamp 1732943601
transform -1 0 1636 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1732943601
transform 1 0 1636 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_11
timestamp 1732943601
transform 1 0 1732 0 1 1705
box -2 -3 50 103
use BUFX4  BUFX4_24
timestamp 1732943601
transform 1 0 1780 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1732943601
transform 1 0 1812 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_93
timestamp 1732943601
transform 1 0 1836 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_14
timestamp 1732943601
transform -1 0 1884 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_60
timestamp 1732943601
transform 1 0 1884 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_3_0
timestamp 1732943601
transform -1 0 1940 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1732943601
transform -1 0 1948 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_211
timestamp 1732943601
transform -1 0 1972 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_269
timestamp 1732943601
transform -1 0 2004 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1732943601
transform -1 0 2100 0 1 1705
box -2 -3 98 103
use BUFX4  BUFX4_58
timestamp 1732943601
transform 1 0 2100 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_83
timestamp 1732943601
transform 1 0 2132 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1732943601
transform -1 0 2252 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_164
timestamp 1732943601
transform 1 0 2252 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1732943601
transform -1 0 2308 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1732943601
transform 1 0 4 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_102
timestamp 1732943601
transform -1 0 132 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1732943601
transform -1 0 164 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1732943601
transform 1 0 164 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_82
timestamp 1732943601
transform 1 0 260 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1732943601
transform -1 0 324 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_85
timestamp 1732943601
transform 1 0 324 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_0_0
timestamp 1732943601
transform -1 0 364 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1732943601
transform -1 0 372 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_79
timestamp 1732943601
transform -1 0 420 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1732943601
transform 1 0 420 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_281
timestamp 1732943601
transform 1 0 516 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_280
timestamp 1732943601
transform -1 0 580 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1732943601
transform -1 0 612 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_36
timestamp 1732943601
transform 1 0 612 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_290
timestamp 1732943601
transform -1 0 692 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_51
timestamp 1732943601
transform 1 0 692 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_7
timestamp 1732943601
transform -1 0 772 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1732943601
transform -1 0 868 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_276
timestamp 1732943601
transform -1 0 900 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_1_0
timestamp 1732943601
transform -1 0 908 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1732943601
transform -1 0 916 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_277
timestamp 1732943601
transform -1 0 948 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_57
timestamp 1732943601
transform 1 0 948 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_58
timestamp 1732943601
transform 1 0 996 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_56
timestamp 1732943601
transform -1 0 1092 0 -1 1905
box -2 -3 50 103
use BUFX4  BUFX4_52
timestamp 1732943601
transform -1 0 1124 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1732943601
transform 1 0 1124 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_286
timestamp 1732943601
transform 1 0 1156 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_287
timestamp 1732943601
transform -1 0 1220 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1732943601
transform -1 0 1316 0 -1 1905
box -2 -3 98 103
use INVX4  INVX4_1
timestamp 1732943601
transform 1 0 1316 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_64
timestamp 1732943601
transform -1 0 1388 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_2_0
timestamp 1732943601
transform 1 0 1388 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1732943601
transform 1 0 1396 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_83
timestamp 1732943601
transform 1 0 1404 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_288
timestamp 1732943601
transform 1 0 1436 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_289
timestamp 1732943601
transform 1 0 1468 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1732943601
transform 1 0 1500 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_168
timestamp 1732943601
transform 1 0 1596 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_211
timestamp 1732943601
transform -1 0 1652 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1732943601
transform -1 0 1668 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1732943601
transform -1 0 1764 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_173
timestamp 1732943601
transform 1 0 1764 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_216
timestamp 1732943601
transform -1 0 1820 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_2
timestamp 1732943601
transform 1 0 1820 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_62
timestamp 1732943601
transform 1 0 1868 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_3_0
timestamp 1732943601
transform 1 0 1916 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1732943601
transform 1 0 1924 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_3
timestamp 1732943601
transform 1 0 1932 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_12
timestamp 1732943601
transform 1 0 1980 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_10
timestamp 1732943601
transform 1 0 2028 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1732943601
transform -1 0 2172 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_9
timestamp 1732943601
transform 1 0 2172 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_10
timestamp 1732943601
transform -1 0 2228 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1732943601
transform 1 0 2228 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_203
timestamp 1732943601
transform -1 0 2284 0 -1 1905
box -2 -3 34 103
use FILL  FILL_19_1
timestamp 1732943601
transform -1 0 2292 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_2
timestamp 1732943601
transform -1 0 2300 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_3
timestamp 1732943601
transform -1 0 2308 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1732943601
transform -1 0 100 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_112
timestamp 1732943601
transform -1 0 132 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1732943601
transform -1 0 164 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1732943601
transform -1 0 196 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1732943601
transform -1 0 228 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1732943601
transform 1 0 228 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1732943601
transform -1 0 292 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1732943601
transform 1 0 292 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_0_0
timestamp 1732943601
transform 1 0 388 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1732943601
transform 1 0 396 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1732943601
transform 1 0 404 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_283
timestamp 1732943601
transform -1 0 532 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_35
timestamp 1732943601
transform -1 0 580 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_291
timestamp 1732943601
transform 1 0 580 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1732943601
transform 1 0 612 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_228
timestamp 1732943601
transform 1 0 708 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_92
timestamp 1732943601
transform 1 0 740 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1732943601
transform -1 0 804 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1732943601
transform -1 0 836 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_239
timestamp 1732943601
transform 1 0 836 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_238
timestamp 1732943601
transform 1 0 868 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_1_0
timestamp 1732943601
transform 1 0 900 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1732943601
transform 1 0 908 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1732943601
transform 1 0 916 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_237
timestamp 1732943601
transform 1 0 1012 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_236
timestamp 1732943601
transform 1 0 1044 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1732943601
transform 1 0 1076 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1732943601
transform 1 0 1172 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_90
timestamp 1732943601
transform 1 0 1268 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1732943601
transform -1 0 1332 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1732943601
transform 1 0 1332 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1732943601
transform -1 0 1396 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1732943601
transform -1 0 1404 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1732943601
transform -1 0 1412 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1732943601
transform -1 0 1508 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1732943601
transform -1 0 1604 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_225
timestamp 1732943601
transform 1 0 1604 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1732943601
transform -1 0 1660 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1732943601
transform -1 0 1756 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_57
timestamp 1732943601
transform 1 0 1756 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1732943601
transform -1 0 1812 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_61
timestamp 1732943601
transform -1 0 1860 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_63
timestamp 1732943601
transform 1 0 1860 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1732943601
transform -1 0 1916 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_3_0
timestamp 1732943601
transform -1 0 1924 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1732943601
transform -1 0 1932 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1732943601
transform -1 0 2028 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_9
timestamp 1732943601
transform 1 0 2028 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1732943601
transform -1 0 2084 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1732943601
transform -1 0 2180 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_266
timestamp 1732943601
transform 1 0 2180 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1732943601
transform -1 0 2308 0 1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_12
timestamp 1732943601
transform 1 0 4 0 -1 2105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_4
timestamp 1732943601
transform 1 0 76 0 -1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1732943601
transform 1 0 148 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_97
timestamp 1732943601
transform 1 0 244 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_98
timestamp 1732943601
transform -1 0 308 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1732943601
transform 1 0 308 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_0_0
timestamp 1732943601
transform -1 0 412 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1732943601
transform -1 0 420 0 -1 2105
box -2 -3 10 103
use BUFX4  BUFX4_49
timestamp 1732943601
transform -1 0 452 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1732943601
transform 1 0 452 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_104
timestamp 1732943601
transform 1 0 548 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1732943601
transform -1 0 612 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_50
timestamp 1732943601
transform -1 0 644 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1732943601
transform 1 0 644 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1732943601
transform -1 0 836 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_107
timestamp 1732943601
transform 1 0 836 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_108
timestamp 1732943601
transform -1 0 900 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_1_0
timestamp 1732943601
transform 1 0 900 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1732943601
transform 1 0 908 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1732943601
transform 1 0 916 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1732943601
transform 1 0 1012 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_110
timestamp 1732943601
transform 1 0 1108 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1732943601
transform -1 0 1172 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_100
timestamp 1732943601
transform 1 0 1172 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1732943601
transform 1 0 1204 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1732943601
transform 1 0 1236 0 -1 2105
box -2 -3 98 103
use BUFX4  BUFX4_25
timestamp 1732943601
transform -1 0 1364 0 -1 2105
box -2 -3 34 103
use INVX8  INVX8_9
timestamp 1732943601
transform 1 0 1364 0 -1 2105
box -2 -3 42 103
use FILL  FILL_20_2_0
timestamp 1732943601
transform 1 0 1404 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1732943601
transform 1 0 1412 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1732943601
transform 1 0 1420 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_55
timestamp 1732943601
transform 1 0 1516 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1732943601
transform -1 0 1572 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_59
timestamp 1732943601
transform 1 0 1572 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1732943601
transform -1 0 1700 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_49
timestamp 1732943601
transform 1 0 1700 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1732943601
transform -1 0 1756 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1732943601
transform 1 0 1756 0 -1 2105
box -2 -3 98 103
use INVX8  INVX8_4
timestamp 1732943601
transform -1 0 1892 0 -1 2105
box -2 -3 42 103
use FILL  FILL_20_3_0
timestamp 1732943601
transform -1 0 1900 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1732943601
transform -1 0 1908 0 -1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_13
timestamp 1732943601
transform -1 0 1980 0 -1 2105
box -2 -3 74 103
use MUX2X1  MUX2X1_1
timestamp 1732943601
transform -1 0 2028 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_202
timestamp 1732943601
transform 1 0 2028 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_158
timestamp 1732943601
transform -1 0 2084 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_5
timestamp 1732943601
transform 1 0 2084 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1732943601
transform -1 0 2204 0 -1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_208
timestamp 1732943601
transform -1 0 2228 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_257
timestamp 1732943601
transform 1 0 2228 0 -1 2105
box -2 -3 34 103
use INVX8  INVX8_8
timestamp 1732943601
transform -1 0 2300 0 -1 2105
box -2 -3 42 103
use FILL  FILL_21_1
timestamp 1732943601
transform -1 0 2308 0 -1 2105
box -2 -3 10 103
<< labels >>
flabel metal6 s 376 -30 392 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 880 -30 896 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1750 -22 1754 -18 7 FreeSans 24 270 0 0 en
port 2 nsew
flabel metal3 s 2334 1068 2338 1072 3 FreeSans 24 0 0 0 rw
port 3 nsew
flabel metal3 s -26 2048 -22 2052 7 FreeSans 24 90 0 0 clk
port 4 nsew
flabel metal2 s 814 -22 818 -18 7 FreeSans 24 270 0 0 ras
port 5 nsew
flabel metal2 s 1814 -22 1818 -18 7 FreeSans 24 270 0 0 cas
port 6 nsew
flabel metal2 s 1798 -22 1802 -18 7 FreeSans 24 270 0 0 vas
port 7 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 datain[0]
port 8 nsew
flabel metal2 s 1870 2128 1874 2132 3 FreeSans 24 90 0 0 datain[1]
port 9 nsew
flabel metal2 s 174 -22 178 -18 7 FreeSans 24 270 0 0 datain[2]
port 10 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 datain[3]
port 11 nsew
flabel metal2 s 1078 -22 1082 -18 7 FreeSans 24 270 0 0 datain[4]
port 12 nsew
flabel metal3 s 2334 2048 2338 2052 3 FreeSans 24 90 0 0 datain[5]
port 13 nsew
flabel metal2 s 1382 2128 1386 2132 3 FreeSans 24 90 0 0 datain[6]
port 14 nsew
flabel metal2 s 110 -22 114 -18 7 FreeSans 24 270 0 0 datain[7]
port 15 nsew
flabel metal2 s 1854 -22 1858 -18 7 FreeSans 24 270 0 0 address[0]
port 16 nsew
flabel metal2 s 902 -22 906 -18 7 FreeSans 24 270 0 0 address[1]
port 17 nsew
flabel metal2 s 854 -22 858 -18 7 FreeSans 24 270 0 0 address[2]
port 18 nsew
flabel metal2 s 1934 -22 1938 -18 7 FreeSans 24 270 0 0 address[3]
port 19 nsew
flabel metal2 s 1982 -22 1986 -18 7 FreeSans 24 270 0 0 address[4]
port 20 nsew
flabel metal3 s 2334 768 2338 772 3 FreeSans 24 0 0 0 dataout[0]
port 21 nsew
flabel metal3 s 2334 1248 2338 1252 3 FreeSans 24 0 0 0 dataout[1]
port 22 nsew
flabel metal3 s 2334 748 2338 752 3 FreeSans 24 0 0 0 dataout[2]
port 23 nsew
flabel metal3 s 2334 848 2338 852 3 FreeSans 24 0 0 0 dataout[3]
port 24 nsew
flabel metal3 s 2334 948 2338 952 3 FreeSans 24 0 0 0 dataout[4]
port 25 nsew
flabel metal3 s 2334 968 2338 972 3 FreeSans 24 0 0 0 dataout[5]
port 26 nsew
flabel metal3 s 2334 1348 2338 1352 3 FreeSans 24 0 0 0 dataout[6]
port 27 nsew
flabel metal2 s 1614 -22 1618 -18 7 FreeSans 24 270 0 0 dataout[7]
port 28 nsew
<< end >>
