magic
tech scmos
timestamp 1732942936
<< metal1 >>
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 493 2403 496 2407
rect 1496 2403 1498 2407
rect 1502 2403 1505 2407
rect 1509 2403 1512 2407
rect 114 2368 121 2371
rect 554 2368 561 2371
rect 694 2368 702 2371
rect 741 2368 742 2372
rect 1254 2368 1262 2371
rect 1618 2368 1625 2371
rect 2030 2368 2054 2371
rect 54 2348 65 2351
rect 86 2351 89 2361
rect 86 2348 105 2351
rect 254 2351 258 2352
rect 238 2348 258 2351
rect 310 2351 313 2361
rect 310 2348 329 2351
rect 62 2342 65 2348
rect 570 2348 585 2351
rect 726 2351 729 2361
rect 710 2348 729 2351
rect 1030 2348 1046 2351
rect 1286 2351 1289 2361
rect 1270 2348 1289 2351
rect 1342 2351 1345 2361
rect 1342 2348 1361 2351
rect 1406 2348 1422 2351
rect 1590 2351 1593 2361
rect 1922 2358 1926 2362
rect 1570 2348 1577 2351
rect 1590 2348 1609 2351
rect 1974 2348 1990 2351
rect 2078 2351 2081 2361
rect 2062 2348 2081 2351
rect 2486 2351 2489 2361
rect 2486 2348 2505 2351
rect 86 2338 94 2341
rect 206 2338 214 2341
rect 310 2338 318 2341
rect 974 2338 982 2341
rect 1282 2338 1289 2341
rect 1310 2338 1318 2341
rect 1590 2338 1598 2341
rect 1806 2338 1818 2341
rect 14 2328 33 2331
rect 1494 2328 1529 2331
rect 2213 2318 2214 2322
rect 984 2303 986 2307
rect 990 2303 993 2307
rect 997 2303 1000 2307
rect 2016 2303 2018 2307
rect 2022 2303 2025 2307
rect 2029 2303 2032 2307
rect 2050 2288 2051 2292
rect 1166 2278 1185 2281
rect 1622 2278 1641 2281
rect 1893 2278 1894 2282
rect 1006 2272 1009 2278
rect 370 2268 377 2271
rect 398 2268 406 2271
rect 1006 2268 1010 2272
rect 1242 2268 1249 2271
rect 1718 2268 1730 2271
rect 1962 2268 1969 2271
rect 2278 2268 2286 2271
rect 2310 2271 2314 2274
rect 2302 2268 2314 2271
rect 50 2258 65 2261
rect 198 2258 217 2261
rect 398 2258 417 2261
rect 574 2258 582 2261
rect 670 2258 678 2261
rect 874 2258 889 2261
rect 894 2258 910 2261
rect 1086 2258 1094 2261
rect 1142 2258 1150 2261
rect 1230 2261 1233 2268
rect 1230 2258 1249 2261
rect 1478 2258 1486 2261
rect 1554 2258 1561 2261
rect 1854 2258 1862 2261
rect 1990 2258 2009 2261
rect 2302 2262 2305 2268
rect 2210 2258 2217 2261
rect 2278 2258 2297 2261
rect 198 2248 201 2258
rect 398 2248 401 2258
rect 858 2248 865 2251
rect 1094 2248 1113 2251
rect 1394 2248 1398 2252
rect 1406 2248 1425 2251
rect 1990 2248 1993 2258
rect 2278 2248 2281 2258
rect 933 2218 934 2222
rect 1141 2218 1142 2222
rect 1938 2218 1939 2222
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 493 2203 496 2207
rect 1496 2203 1498 2207
rect 1502 2203 1505 2207
rect 1509 2203 1512 2207
rect 2397 2188 2398 2192
rect 378 2168 381 2172
rect 701 2168 702 2172
rect 1198 2168 1209 2171
rect 1822 2168 1833 2171
rect 1198 2166 1202 2168
rect 1822 2166 1826 2168
rect 126 2151 129 2161
rect 922 2158 926 2162
rect 934 2158 953 2161
rect 1026 2158 1033 2161
rect 126 2148 145 2151
rect 258 2148 265 2151
rect 390 2148 398 2151
rect 494 2151 498 2153
rect 470 2148 498 2151
rect 970 2148 977 2151
rect 1006 2148 1014 2151
rect 1238 2148 1246 2151
rect 1326 2151 1329 2161
rect 1326 2148 1345 2151
rect 310 2138 329 2141
rect 786 2138 793 2141
rect 1062 2138 1065 2148
rect 1590 2151 1593 2161
rect 1590 2148 1609 2151
rect 1646 2151 1649 2161
rect 1646 2148 1665 2151
rect 1882 2148 1889 2151
rect 2070 2151 2073 2161
rect 2182 2158 2201 2161
rect 2210 2158 2214 2162
rect 2070 2148 2089 2151
rect 1326 2138 1334 2141
rect 1646 2138 1654 2141
rect 2046 2141 2049 2148
rect 2382 2151 2385 2161
rect 2366 2148 2385 2151
rect 2014 2138 2049 2141
rect 2070 2138 2078 2141
rect 326 2128 329 2138
rect 277 2118 278 2122
rect 984 2103 986 2107
rect 990 2103 993 2107
rect 997 2103 1000 2107
rect 2016 2103 2018 2107
rect 2022 2103 2025 2107
rect 2029 2103 2032 2107
rect 2026 2088 2041 2091
rect 278 2074 282 2078
rect 750 2072 753 2081
rect 1390 2078 1409 2081
rect 1950 2072 1953 2081
rect 2454 2078 2462 2081
rect 542 2068 550 2071
rect 1506 2068 1514 2071
rect 1678 2068 1686 2071
rect 1822 2068 1838 2071
rect 1982 2068 1990 2071
rect 2298 2068 2305 2071
rect 2462 2068 2478 2071
rect 126 2058 145 2061
rect 182 2058 201 2061
rect 246 2058 266 2061
rect 366 2058 385 2061
rect 398 2058 406 2061
rect 534 2058 553 2061
rect 586 2058 593 2061
rect 926 2058 942 2061
rect 1082 2058 1089 2061
rect 1202 2058 1209 2061
rect 1678 2058 1697 2061
rect 1890 2058 1897 2061
rect 1982 2058 1985 2068
rect 2090 2058 2097 2061
rect 2370 2058 2385 2061
rect 2462 2058 2465 2068
rect 126 2048 129 2058
rect 182 2048 185 2058
rect 262 2057 266 2058
rect 382 2048 385 2058
rect 670 2052 674 2057
rect 514 2048 529 2051
rect 1678 2048 1681 2058
rect 605 2018 606 2022
rect 1861 2018 1862 2022
rect 2002 2018 2003 2022
rect 2274 2018 2275 2022
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 493 2003 496 2007
rect 1496 2003 1498 2007
rect 1502 2003 1505 2007
rect 1509 2003 1512 2007
rect 634 1988 635 1992
rect 797 1988 798 1992
rect 1837 1988 1838 1992
rect 1733 1978 1734 1982
rect 395 1968 398 1972
rect 834 1968 837 1972
rect 1618 1968 1621 1972
rect 2210 1968 2217 1971
rect 294 1951 297 1961
rect 306 1958 310 1962
rect 50 1948 65 1951
rect 278 1948 297 1951
rect 590 1951 593 1961
rect 982 1958 990 1961
rect 574 1948 593 1951
rect 650 1948 657 1951
rect 698 1948 705 1951
rect 746 1948 753 1951
rect 94 1938 106 1941
rect 486 1938 510 1941
rect 562 1938 569 1941
rect 658 1938 665 1941
rect 710 1938 718 1941
rect 774 1941 777 1948
rect 974 1948 998 1951
rect 1718 1951 1721 1961
rect 2138 1958 2142 1962
rect 1702 1948 1721 1951
rect 1838 1948 1865 1951
rect 2182 1951 2185 1961
rect 2182 1948 2201 1951
rect 2394 1948 2401 1951
rect 766 1938 777 1941
rect 994 1938 1017 1941
rect 1022 1938 1034 1941
rect 1030 1936 1034 1938
rect 1062 1932 1065 1942
rect 1262 1938 1270 1941
rect 1322 1938 1329 1941
rect 1390 1938 1417 1941
rect 1478 1938 1486 1941
rect 1962 1938 1977 1941
rect 2182 1938 2190 1941
rect 1149 1928 1150 1932
rect 1293 1918 1294 1922
rect 1389 1918 1390 1922
rect 1938 1918 1939 1922
rect 984 1903 986 1907
rect 990 1903 993 1907
rect 997 1903 1000 1907
rect 2016 1903 2018 1907
rect 2022 1903 2025 1907
rect 2029 1903 2032 1907
rect 730 1888 731 1892
rect 1874 1888 1875 1892
rect 2005 1888 2006 1892
rect 2034 1888 2041 1891
rect 414 1878 433 1881
rect 1422 1878 1441 1881
rect 342 1876 346 1878
rect 1102 1872 1106 1877
rect 54 1868 62 1871
rect 110 1868 118 1871
rect 722 1868 729 1871
rect 1118 1871 1122 1874
rect 1118 1868 1129 1871
rect 1146 1868 1153 1871
rect 1178 1868 1185 1871
rect 1566 1868 1585 1871
rect 1830 1868 1838 1871
rect 1854 1868 1862 1871
rect 2014 1868 2030 1871
rect 2070 1868 2073 1878
rect 2202 1868 2217 1871
rect 2278 1868 2286 1871
rect 1582 1862 1585 1868
rect 14 1858 33 1861
rect 86 1858 105 1861
rect 114 1858 129 1861
rect 702 1858 710 1861
rect 790 1858 798 1861
rect 862 1858 881 1861
rect 918 1858 937 1861
rect 970 1858 977 1861
rect 1006 1858 1014 1861
rect 1134 1858 1153 1861
rect 1166 1858 1182 1861
rect 1198 1858 1206 1861
rect 1266 1858 1273 1861
rect 1622 1858 1641 1861
rect 1706 1858 1721 1861
rect 1830 1858 1849 1861
rect 2082 1858 2097 1861
rect 2190 1858 2206 1861
rect 2278 1858 2297 1861
rect 30 1848 33 1858
rect 86 1848 89 1858
rect 878 1848 881 1858
rect 934 1848 937 1858
rect 1150 1848 1153 1858
rect 1622 1848 1625 1858
rect 1830 1848 1833 1858
rect 2278 1848 2281 1858
rect 1622 1842 1626 1844
rect 1682 1838 1685 1842
rect 1922 1838 1925 1842
rect 690 1828 691 1832
rect 1778 1828 1779 1832
rect 594 1818 595 1822
rect 2178 1818 2179 1822
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 493 1803 496 1807
rect 1496 1803 1498 1807
rect 1502 1803 1505 1807
rect 1509 1803 1512 1807
rect 1413 1788 1414 1792
rect 2002 1788 2003 1792
rect 1741 1768 1742 1772
rect 1778 1768 1781 1772
rect 134 1751 137 1758
rect 118 1748 137 1751
rect 206 1751 209 1761
rect 206 1748 225 1751
rect 290 1748 297 1751
rect 510 1748 518 1751
rect 614 1751 617 1761
rect 626 1758 630 1762
rect 598 1748 617 1751
rect 746 1748 753 1751
rect 878 1751 882 1753
rect 878 1748 897 1751
rect 1166 1751 1169 1761
rect 1150 1748 1169 1751
rect 1246 1748 1254 1751
rect 1526 1751 1529 1761
rect 1538 1758 1542 1762
rect 1494 1748 1529 1751
rect 1726 1751 1729 1761
rect 2490 1758 2494 1762
rect 1710 1748 1729 1751
rect 1810 1748 1817 1751
rect 1918 1748 1926 1751
rect 2162 1748 2177 1751
rect 2294 1748 2302 1751
rect 2414 1748 2422 1751
rect 138 1738 145 1741
rect 206 1738 214 1741
rect 510 1738 526 1741
rect 554 1738 561 1741
rect 890 1738 897 1741
rect 986 1738 1009 1741
rect 1085 1738 1086 1742
rect 1162 1738 1169 1741
rect 1438 1741 1441 1748
rect 1326 1738 1353 1741
rect 1438 1738 1449 1741
rect 1658 1738 1665 1741
rect 2218 1738 2225 1741
rect 2314 1738 2321 1741
rect 1277 1728 1278 1732
rect 2282 1728 2283 1732
rect 2058 1718 2059 1722
rect 2370 1718 2371 1722
rect 984 1703 986 1707
rect 990 1703 993 1707
rect 997 1703 1000 1707
rect 2016 1703 2018 1707
rect 2022 1703 2025 1707
rect 2029 1703 2032 1707
rect 706 1688 707 1692
rect 1221 1688 1222 1692
rect 1309 1688 1310 1692
rect 1778 1688 1779 1692
rect 1813 1688 1814 1692
rect 453 1678 454 1682
rect 2066 1678 2067 1682
rect 70 1668 82 1671
rect 406 1662 409 1671
rect 806 1668 814 1671
rect 830 1668 838 1671
rect 1194 1668 1201 1671
rect 1598 1668 1625 1671
rect 1742 1668 1750 1671
rect 2090 1668 2097 1671
rect 2374 1668 2377 1678
rect 238 1658 254 1661
rect 310 1658 329 1661
rect 362 1658 369 1661
rect 482 1658 497 1661
rect 654 1658 673 1661
rect 718 1658 726 1661
rect 738 1658 745 1661
rect 806 1658 825 1661
rect 982 1658 1017 1661
rect 1146 1658 1153 1661
rect 1198 1661 1201 1668
rect 1166 1658 1185 1661
rect 1198 1658 1209 1661
rect 1254 1658 1273 1661
rect 1426 1658 1433 1661
rect 1506 1658 1513 1661
rect 1658 1658 1665 1661
rect 1678 1658 1697 1661
rect 1790 1658 1798 1661
rect 1874 1658 1889 1661
rect 1950 1658 1969 1661
rect 2078 1658 2097 1661
rect 2126 1658 2145 1661
rect 2218 1658 2233 1661
rect 326 1648 329 1658
rect 642 1648 646 1652
rect 654 1648 657 1658
rect 806 1648 809 1658
rect 1014 1648 1017 1658
rect 1166 1648 1169 1658
rect 1270 1648 1273 1658
rect 1282 1648 1286 1652
rect 1678 1648 1681 1658
rect 1950 1648 1953 1658
rect 2094 1652 2097 1658
rect 2142 1648 2145 1658
rect 189 1638 190 1642
rect 381 1638 382 1642
rect 1115 1638 1118 1642
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 493 1603 496 1607
rect 1496 1603 1498 1607
rect 1502 1603 1505 1607
rect 1509 1603 1512 1607
rect 365 1588 366 1592
rect 389 1588 390 1592
rect 445 1588 446 1592
rect 517 1588 518 1592
rect 1314 1588 1315 1592
rect 1525 1588 1526 1592
rect 1802 1588 1803 1592
rect 94 1568 102 1571
rect 1230 1568 1238 1571
rect 1602 1568 1609 1571
rect 2074 1568 2077 1572
rect 2370 1568 2377 1571
rect 38 1548 46 1551
rect 126 1551 129 1561
rect 110 1548 129 1551
rect 162 1548 169 1551
rect 230 1551 233 1561
rect 230 1548 249 1551
rect 306 1548 321 1551
rect 378 1548 385 1551
rect 426 1548 433 1551
rect 498 1548 513 1551
rect 654 1551 657 1561
rect 782 1558 801 1561
rect 638 1548 657 1551
rect 774 1548 782 1551
rect 1262 1551 1265 1561
rect 1246 1548 1265 1551
rect 1374 1548 1382 1551
rect 1482 1548 1513 1551
rect 1574 1551 1577 1561
rect 1574 1548 1593 1551
rect 1750 1551 1753 1561
rect 1750 1548 1769 1551
rect 1814 1548 1822 1551
rect 1950 1551 1953 1561
rect 2006 1558 2014 1561
rect 1934 1548 1953 1551
rect 1998 1548 2022 1551
rect 2106 1548 2113 1551
rect 2342 1551 2345 1561
rect 2510 1558 2518 1561
rect 2342 1548 2361 1551
rect 478 1538 510 1541
rect 1258 1538 1265 1541
rect 1574 1538 1582 1541
rect 1974 1538 1982 1541
rect 2018 1538 2041 1541
rect 2342 1538 2350 1541
rect 2490 1538 2497 1541
rect 550 1533 554 1538
rect 398 1528 409 1531
rect 958 1528 977 1531
rect 982 1528 998 1531
rect 1030 1528 1049 1531
rect 1086 1528 1105 1531
rect 181 1518 182 1522
rect 2506 1518 2507 1522
rect 984 1503 986 1507
rect 990 1503 993 1507
rect 997 1503 1000 1507
rect 2016 1503 2018 1507
rect 2022 1503 2025 1507
rect 2029 1503 2032 1507
rect 338 1488 339 1492
rect 542 1472 545 1481
rect 570 1478 577 1481
rect 2058 1478 2059 1482
rect 122 1468 129 1471
rect 366 1468 377 1471
rect 446 1468 454 1471
rect 598 1468 609 1471
rect 58 1458 65 1461
rect 110 1458 129 1461
rect 190 1458 198 1461
rect 278 1458 297 1461
rect 318 1458 329 1461
rect 518 1461 521 1468
rect 518 1458 529 1461
rect 766 1458 785 1461
rect 1206 1458 1214 1461
rect 1486 1462 1489 1471
rect 1590 1468 1598 1471
rect 1789 1468 1790 1472
rect 1962 1468 1969 1471
rect 1990 1468 1998 1471
rect 2014 1468 2022 1471
rect 1562 1458 1577 1461
rect 1590 1458 1609 1461
rect 2230 1462 2233 1471
rect 1802 1458 1809 1461
rect 1990 1458 2009 1461
rect 2238 1458 2257 1461
rect 2270 1458 2278 1461
rect 126 1448 129 1458
rect 278 1448 281 1458
rect 326 1452 329 1458
rect 346 1448 353 1451
rect 1486 1448 1505 1451
rect 1590 1448 1593 1458
rect 1990 1448 1993 1458
rect 2254 1448 2257 1458
rect 2266 1448 2270 1452
rect 94 1438 102 1441
rect 413 1418 414 1422
rect 533 1418 534 1422
rect 1194 1418 1195 1422
rect 1938 1418 1939 1422
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 493 1403 496 1407
rect 1496 1403 1498 1407
rect 1502 1403 1505 1407
rect 1509 1403 1512 1407
rect 397 1388 398 1392
rect 698 1388 699 1392
rect 837 1388 838 1392
rect 1110 1368 1118 1371
rect 1462 1368 1470 1371
rect 2018 1368 2025 1371
rect 2194 1368 2197 1372
rect 166 1351 169 1361
rect 166 1348 185 1351
rect 218 1348 225 1351
rect 378 1348 385 1351
rect 654 1348 662 1351
rect 714 1348 721 1351
rect 822 1351 825 1361
rect 806 1348 825 1351
rect 878 1351 881 1361
rect 878 1348 897 1351
rect 286 1338 294 1341
rect 510 1338 518 1341
rect 790 1341 793 1348
rect 962 1348 969 1351
rect 1142 1351 1145 1361
rect 1126 1348 1145 1351
rect 1246 1351 1249 1361
rect 1230 1348 1249 1351
rect 1406 1348 1422 1351
rect 1490 1348 1521 1351
rect 1726 1351 1729 1361
rect 1690 1348 1697 1351
rect 1710 1348 1729 1351
rect 1974 1351 1977 1361
rect 1974 1348 1993 1351
rect 2142 1351 2145 1361
rect 2126 1348 2145 1351
rect 658 1338 665 1341
rect 670 1338 689 1341
rect 790 1338 801 1341
rect 878 1338 886 1341
rect 1138 1338 1145 1341
rect 1694 1341 1697 1348
rect 1694 1338 1705 1341
rect 1722 1338 1729 1341
rect 1790 1338 1817 1341
rect 1898 1338 1913 1341
rect 1974 1338 1982 1341
rect 1998 1338 2014 1341
rect 2390 1338 2409 1341
rect 642 1328 646 1332
rect 770 1318 771 1322
rect 1482 1318 1483 1322
rect 1533 1318 1534 1322
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 2016 1303 2018 1307
rect 2022 1303 2025 1307
rect 2029 1303 2032 1307
rect 490 1288 505 1291
rect 1026 1288 1027 1292
rect 1914 1288 1915 1292
rect 2370 1288 2371 1292
rect 781 1278 782 1282
rect 846 1278 854 1282
rect 2178 1278 2179 1282
rect 846 1272 849 1278
rect 366 1268 374 1271
rect 414 1268 430 1271
rect 670 1268 678 1271
rect 898 1268 913 1271
rect 982 1268 1006 1271
rect 1046 1268 1065 1271
rect 1106 1268 1113 1271
rect 1174 1268 1182 1271
rect 1341 1268 1342 1272
rect 1446 1268 1454 1271
rect 1541 1268 1542 1272
rect 1618 1268 1625 1271
rect 1886 1268 1897 1271
rect 1934 1268 1953 1271
rect 2122 1268 2129 1271
rect 2453 1268 2454 1272
rect 38 1258 54 1261
rect 290 1258 297 1261
rect 414 1258 422 1261
rect 478 1258 494 1261
rect 606 1258 625 1261
rect 906 1258 913 1261
rect 1046 1258 1049 1268
rect 1058 1258 1065 1261
rect 1154 1258 1161 1261
rect 1174 1258 1193 1261
rect 1406 1258 1425 1261
rect 1606 1258 1625 1261
rect 1726 1258 1745 1261
rect 1894 1262 1897 1268
rect 1934 1258 1937 1268
rect 2110 1258 2129 1261
rect 2406 1258 2409 1268
rect 2458 1258 2473 1261
rect 110 1248 129 1251
rect 622 1248 625 1258
rect 1174 1248 1177 1258
rect 1422 1248 1425 1258
rect 1622 1248 1625 1258
rect 1726 1248 1729 1258
rect 2126 1248 2129 1258
rect 2214 1248 2233 1251
rect 2242 1248 2246 1252
rect 2026 1238 2029 1242
rect 1674 1218 1675 1222
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 1496 1203 1498 1207
rect 1502 1203 1505 1207
rect 1509 1203 1512 1207
rect 773 1188 774 1192
rect 1786 1188 1787 1192
rect 1722 1168 1723 1172
rect 102 1151 105 1161
rect 282 1158 289 1161
rect 586 1158 590 1162
rect 86 1148 105 1151
rect 118 1148 126 1151
rect 262 1148 281 1151
rect 298 1148 313 1151
rect 366 1148 374 1151
rect 434 1148 441 1151
rect 598 1151 601 1161
rect 598 1148 617 1151
rect 630 1148 641 1151
rect 754 1148 761 1151
rect 822 1151 825 1161
rect 966 1158 974 1161
rect 822 1148 841 1151
rect 1014 1151 1017 1161
rect 982 1148 1017 1151
rect 1038 1148 1046 1151
rect 1070 1151 1073 1161
rect 1054 1148 1073 1151
rect 1146 1148 1161 1151
rect 1438 1151 1441 1161
rect 1402 1148 1417 1151
rect 1422 1148 1441 1151
rect 1454 1148 1462 1151
rect 278 1142 281 1148
rect 454 1138 462 1141
rect 630 1141 633 1148
rect 626 1138 633 1141
rect 970 1138 977 1141
rect 1038 1138 1041 1148
rect 1286 1138 1294 1141
rect 1398 1138 1406 1141
rect 1414 1138 1417 1148
rect 1734 1151 1737 1161
rect 1878 1158 1897 1161
rect 1734 1148 1753 1151
rect 1798 1148 1814 1151
rect 1950 1151 1953 1161
rect 2202 1158 2206 1162
rect 1950 1148 1969 1151
rect 2042 1148 2057 1151
rect 1462 1138 1470 1141
rect 1922 1138 1929 1141
rect 1974 1138 2002 1141
rect 2222 1141 2225 1148
rect 2222 1138 2233 1141
rect 1998 1136 2002 1138
rect 1010 1128 1017 1131
rect 2322 1128 2323 1132
rect 2274 1118 2275 1122
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 2016 1103 2018 1107
rect 2022 1103 2025 1107
rect 2029 1103 2032 1107
rect 1010 1088 1017 1091
rect 1346 1088 1347 1092
rect 94 1071 98 1074
rect 558 1072 562 1077
rect 94 1068 102 1071
rect 230 1062 233 1071
rect 250 1068 257 1071
rect 470 1068 478 1071
rect 686 1068 694 1071
rect 718 1068 726 1071
rect 750 1071 754 1074
rect 742 1068 754 1071
rect 838 1068 850 1071
rect 990 1068 998 1071
rect 1030 1068 1038 1071
rect 1226 1068 1233 1071
rect 1326 1068 1334 1071
rect 1446 1068 1457 1071
rect 1538 1068 1545 1071
rect 1598 1068 1625 1071
rect 238 1058 257 1061
rect 330 1058 345 1061
rect 526 1058 546 1061
rect 718 1058 737 1061
rect 802 1058 809 1061
rect 1046 1058 1057 1061
rect 1238 1058 1257 1061
rect 1546 1058 1553 1061
rect 1678 1061 1681 1071
rect 1702 1068 1710 1071
rect 2026 1068 2057 1071
rect 1662 1058 1681 1061
rect 1734 1058 1753 1061
rect 1818 1058 1825 1061
rect 1946 1058 1953 1061
rect 2022 1058 2030 1061
rect 2238 1062 2241 1071
rect 2390 1062 2393 1071
rect 2398 1058 2417 1061
rect 254 1048 257 1058
rect 542 1057 546 1058
rect 646 1048 665 1051
rect 718 1048 721 1058
rect 1054 1052 1057 1058
rect 994 1048 1017 1051
rect 1082 1048 1089 1051
rect 1114 1048 1121 1051
rect 1222 1048 1230 1051
rect 1254 1048 1257 1058
rect 1782 1052 1786 1057
rect 2414 1048 2417 1058
rect 1330 1038 1345 1041
rect 1758 1041 1762 1044
rect 1758 1038 1769 1041
rect 2195 1038 2198 1042
rect 514 1018 515 1022
rect 954 1018 955 1022
rect 1877 1018 1878 1022
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 1496 1003 1498 1007
rect 1502 1003 1505 1007
rect 1509 1003 1512 1007
rect 21 988 22 992
rect 2114 988 2115 992
rect 2490 988 2491 992
rect 138 948 145 951
rect 206 951 209 961
rect 190 948 209 951
rect 262 951 265 961
rect 246 948 265 951
rect 182 938 185 948
rect 486 948 510 951
rect 686 951 689 961
rect 974 958 1009 961
rect 1018 958 1022 962
rect 1350 952 1353 961
rect 670 948 689 951
rect 714 948 729 951
rect 878 948 894 951
rect 1022 948 1030 951
rect 1142 948 1158 951
rect 1446 948 1454 951
rect 1538 948 1545 951
rect 1650 948 1665 951
rect 1918 951 1921 961
rect 1902 948 1921 951
rect 2050 948 2073 951
rect 2278 948 2286 951
rect 2318 951 2321 961
rect 2318 948 2337 951
rect 202 938 209 941
rect 286 938 294 941
rect 382 932 385 942
rect 658 938 665 941
rect 958 938 966 941
rect 982 938 998 941
rect 1154 938 1161 941
rect 1490 938 1497 941
rect 1694 938 1706 941
rect 1914 938 1921 941
rect 2262 938 2265 948
rect 2502 948 2510 951
rect 2286 938 2294 941
rect 157 928 158 932
rect 1606 931 1610 933
rect 1602 928 1610 931
rect 949 918 950 922
rect 1170 918 1171 922
rect 1205 918 1206 922
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 2016 903 2018 907
rect 2022 903 2025 907
rect 2029 903 2032 907
rect 426 888 427 892
rect 829 888 830 892
rect 906 888 907 892
rect 1962 888 1963 892
rect 1662 878 1681 881
rect 398 868 406 871
rect 598 868 606 871
rect 838 868 846 871
rect 886 868 894 871
rect 934 868 942 871
rect 982 868 1006 871
rect 1514 868 1521 871
rect 1538 868 1545 871
rect 1566 868 1577 871
rect 1682 868 1689 871
rect 2142 868 2153 871
rect 2254 868 2262 871
rect 134 858 142 861
rect 154 858 161 861
rect 414 861 417 868
rect 398 858 417 861
rect 498 858 513 861
rect 574 858 593 861
rect 706 858 713 861
rect 878 858 889 861
rect 430 848 438 851
rect 574 848 577 858
rect 886 852 889 858
rect 910 858 918 861
rect 1086 858 1102 861
rect 1174 858 1193 861
rect 1238 858 1246 861
rect 1278 858 1297 861
rect 1354 858 1369 861
rect 1574 862 1577 868
rect 1526 858 1545 861
rect 1610 858 1617 861
rect 1810 858 1817 861
rect 1950 861 1953 868
rect 2142 862 2145 868
rect 1934 858 1953 861
rect 1982 858 2001 861
rect 2014 858 2030 861
rect 2254 861 2257 868
rect 2246 858 2257 861
rect 2270 858 2289 861
rect 2430 858 2438 861
rect 910 848 913 858
rect 1174 848 1177 858
rect 1278 848 1281 858
rect 1542 848 1545 858
rect 1998 848 2001 858
rect 2010 848 2014 852
rect 2286 848 2289 858
rect 2298 848 2302 852
rect 910 842 914 844
rect 674 838 677 842
rect 317 818 318 822
rect 629 818 630 822
rect 1226 818 1227 822
rect 1629 818 1630 822
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 1496 803 1498 807
rect 1502 803 1505 807
rect 1509 803 1512 807
rect 586 768 589 772
rect 1954 768 1955 772
rect 1574 766 1578 768
rect 206 751 209 761
rect 206 748 225 751
rect 318 751 321 761
rect 318 748 337 751
rect 478 748 494 751
rect 690 748 697 751
rect 750 751 753 761
rect 750 748 769 751
rect 1006 751 1009 761
rect 974 748 1009 751
rect 1114 748 1121 751
rect 1198 748 1217 751
rect 1222 748 1230 751
rect 1242 748 1249 751
rect 1318 742 1321 751
rect 1358 748 1366 751
rect 1510 748 1518 751
rect 1582 748 1601 751
rect 1666 748 1673 751
rect 1686 751 1689 761
rect 1686 748 1705 751
rect 1878 748 1886 751
rect 1966 751 1969 761
rect 2154 758 2161 761
rect 1946 748 1953 751
rect 1966 748 1985 751
rect 2110 748 2118 751
rect 2166 751 2169 758
rect 2166 748 2185 751
rect 2202 748 2217 751
rect 2298 748 2313 751
rect 2494 748 2518 751
rect 318 738 326 741
rect 710 738 729 741
rect 1090 738 1105 741
rect 1446 738 1470 741
rect 1566 738 1574 741
rect 1938 738 1945 741
rect 2026 738 2049 741
rect 2210 738 2217 741
rect 150 728 169 731
rect 262 728 281 731
rect 498 728 513 731
rect 518 728 537 731
rect 1110 728 1118 731
rect 2430 728 2449 731
rect 930 718 931 722
rect 1298 718 1299 722
rect 1418 718 1419 722
rect 1914 718 1915 722
rect 2098 718 2099 722
rect 2138 718 2139 722
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 2016 703 2018 707
rect 2022 703 2025 707
rect 2029 703 2032 707
rect 942 688 961 691
rect 1114 688 1115 692
rect 958 682 961 688
rect 778 678 782 682
rect 1162 678 1166 682
rect 1366 678 1385 681
rect 1722 678 1723 682
rect 1893 678 1894 682
rect 2034 678 2038 682
rect 382 668 398 671
rect 598 668 617 671
rect 14 658 33 661
rect 66 658 73 661
rect 238 658 254 661
rect 334 658 342 661
rect 438 658 446 661
rect 486 658 502 661
rect 642 658 649 661
rect 686 658 697 661
rect 702 658 710 661
rect 822 661 825 671
rect 1098 668 1105 671
rect 1598 671 1602 674
rect 2358 672 2361 678
rect 1598 668 1609 671
rect 1654 668 1662 671
rect 2026 668 2033 671
rect 2058 668 2073 671
rect 822 658 841 661
rect 1010 658 1025 661
rect 1130 658 1137 661
rect 1294 658 1313 661
rect 1334 661 1337 668
rect 1334 658 1345 661
rect 2150 662 2153 671
rect 2258 668 2265 671
rect 2358 668 2362 672
rect 2414 668 2426 671
rect 1450 658 1457 661
rect 1542 658 1558 661
rect 1614 658 1633 661
rect 1658 658 1665 661
rect 1782 658 1790 661
rect 1962 658 1969 661
rect 2010 658 2025 661
rect 2086 658 2094 661
rect 2210 658 2217 661
rect 30 648 33 658
rect 686 652 689 658
rect 702 648 705 658
rect 1310 648 1313 658
rect 1630 648 1633 658
rect 626 618 627 622
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 1496 603 1498 607
rect 1502 603 1505 607
rect 1509 603 1512 607
rect 429 588 430 592
rect 474 588 475 592
rect 898 588 899 592
rect 1949 588 1950 592
rect 246 568 254 571
rect 30 551 33 561
rect 14 548 33 551
rect 278 551 281 561
rect 262 548 281 551
rect 654 551 657 561
rect 654 548 673 551
rect 958 548 966 551
rect 1110 551 1113 561
rect 1182 561 1185 568
rect 1182 558 1193 561
rect 1262 558 1281 561
rect 1094 548 1113 551
rect 1158 548 1177 551
rect 1282 548 1289 551
rect 1466 548 1473 551
rect 1550 551 1553 561
rect 1550 548 1569 551
rect 1806 548 1822 551
rect 654 538 662 541
rect 1106 538 1113 541
rect 1466 538 1473 541
rect 1902 541 1905 551
rect 1922 548 1937 551
rect 2022 548 2030 551
rect 2042 548 2049 551
rect 1890 538 1905 541
rect 2250 538 2257 541
rect 590 528 598 531
rect 1430 528 1449 531
rect 1982 528 2001 531
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 2016 503 2018 507
rect 2022 503 2025 507
rect 2029 503 2032 507
rect 277 488 278 492
rect 461 488 462 492
rect 1486 488 1494 491
rect 2282 488 2283 492
rect 1126 476 1130 478
rect 446 468 454 471
rect 470 468 494 471
rect 854 471 858 474
rect 854 468 865 471
rect 882 468 889 471
rect 1018 468 1033 471
rect 1050 468 1057 471
rect 1214 468 1222 471
rect 1394 468 1402 471
rect 2014 468 2030 471
rect 2202 468 2209 471
rect 2302 468 2321 471
rect 2382 468 2390 471
rect 110 458 129 461
rect 258 458 265 461
rect 310 458 329 461
rect 734 458 753 461
rect 870 458 889 461
rect 1038 458 1057 461
rect 1214 458 1233 461
rect 1450 458 1457 461
rect 1566 458 1585 461
rect 1670 458 1678 461
rect 1706 458 1713 461
rect 2190 458 2209 461
rect 2302 461 2305 468
rect 2294 458 2305 461
rect 2314 458 2321 461
rect 2382 458 2401 461
rect 126 448 129 458
rect 138 448 142 452
rect 326 448 329 458
rect 734 448 737 458
rect 886 448 889 458
rect 1054 448 1057 458
rect 1214 448 1217 458
rect 1582 448 1585 458
rect 2206 448 2209 458
rect 2382 448 2385 458
rect 454 442 458 444
rect 510 442 514 444
rect 514 438 521 441
rect 1242 438 1249 441
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 1496 403 1498 407
rect 1502 403 1505 407
rect 1509 403 1512 407
rect 125 388 126 392
rect 373 388 374 392
rect 933 388 934 392
rect 1226 388 1227 392
rect 1714 388 1715 392
rect 1994 388 1995 392
rect 1179 368 1182 372
rect 94 351 98 353
rect 94 348 113 351
rect 174 351 177 361
rect 174 348 193 351
rect 422 351 425 361
rect 406 348 425 351
rect 526 351 529 361
rect 510 348 529 351
rect 542 348 550 351
rect 590 348 601 351
rect 1078 351 1081 361
rect 1078 348 1097 351
rect 174 338 182 341
rect 446 338 465 341
rect 598 341 601 348
rect 1162 348 1169 351
rect 1630 348 1638 351
rect 1726 348 1734 351
rect 1846 351 1849 361
rect 1858 358 1862 362
rect 1806 348 1817 351
rect 1830 348 1849 351
rect 1910 348 1918 351
rect 2090 348 2097 351
rect 2190 348 2198 351
rect 2230 351 2233 361
rect 2230 348 2249 351
rect 2262 348 2273 351
rect 2390 351 2393 361
rect 2390 348 2409 351
rect 598 338 617 341
rect 878 338 897 341
rect 1654 338 1670 341
rect 1686 338 1689 348
rect 1814 341 1817 348
rect 2262 342 2265 348
rect 1814 338 1822 341
rect 2254 338 2262 341
rect 2358 341 2361 348
rect 2358 338 2369 341
rect 2390 338 2398 341
rect 78 332 82 336
rect 878 328 881 338
rect 2318 328 2337 331
rect 1410 318 1411 322
rect 1677 318 1678 322
rect 2034 318 2041 321
rect 2141 318 2142 322
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 2016 303 2018 307
rect 2022 303 2025 307
rect 2029 303 2032 307
rect 1474 288 1475 292
rect 1538 288 1539 292
rect 1986 288 1987 292
rect 2290 288 2291 292
rect 170 268 171 272
rect 786 268 793 271
rect 818 268 825 271
rect 942 268 958 271
rect 1082 268 1089 271
rect 1294 268 1302 271
rect 1590 268 1601 271
rect 2058 268 2065 271
rect 2110 268 2118 271
rect 2154 268 2161 271
rect 14 258 33 261
rect 70 258 89 261
rect 266 258 273 261
rect 590 258 609 261
rect 774 258 793 261
rect 906 258 913 261
rect 1070 258 1089 261
rect 1114 258 1126 261
rect 1142 258 1161 261
rect 1226 258 1233 261
rect 1294 258 1313 261
rect 1590 262 1593 268
rect 1562 258 1569 261
rect 1606 258 1625 261
rect 1682 258 1689 261
rect 1822 258 1841 261
rect 2070 258 2089 261
rect 2134 258 2150 261
rect 2214 258 2222 261
rect 2430 258 2438 261
rect 30 248 33 258
rect 86 248 89 258
rect 98 248 102 252
rect 590 248 593 258
rect 790 248 793 258
rect 1086 248 1089 258
rect 1142 248 1145 258
rect 1294 248 1297 258
rect 1622 248 1625 258
rect 1686 248 1689 258
rect 1838 248 1841 258
rect 1850 248 1854 252
rect 2086 248 2089 258
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 1496 203 1498 207
rect 1502 203 1505 207
rect 1509 203 1512 207
rect 469 188 470 192
rect 2122 188 2123 192
rect 1589 178 1590 182
rect 779 168 782 172
rect 798 168 806 171
rect 1162 168 1165 172
rect 2258 168 2265 171
rect 126 151 129 161
rect 110 148 129 151
rect 178 148 185 151
rect 206 142 209 151
rect 450 148 457 151
rect 630 151 633 161
rect 614 148 633 151
rect 658 148 673 151
rect 830 151 833 161
rect 814 148 833 151
rect 1042 148 1049 151
rect 1110 151 1113 161
rect 1094 148 1113 151
rect 1270 148 1278 151
rect 1406 151 1409 161
rect 1390 148 1409 151
rect 1574 151 1577 161
rect 1710 158 1729 161
rect 1558 148 1577 151
rect 1810 148 1817 151
rect 1878 151 1881 161
rect 1878 148 1897 151
rect 1998 151 2002 153
rect 1998 148 2033 151
rect 2174 151 2177 161
rect 2174 148 2193 151
rect 2230 151 2233 161
rect 2230 148 2249 151
rect 826 138 833 141
rect 854 138 862 141
rect 1325 138 1326 142
rect 1402 138 1409 141
rect 1498 138 1513 141
rect 2018 138 2033 141
rect 2074 138 2081 141
rect 2230 138 2238 141
rect 206 128 225 131
rect 1013 128 1014 132
rect 165 118 166 122
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 2016 103 2018 107
rect 2022 103 2025 107
rect 2029 103 2032 107
rect 498 88 505 91
rect 302 71 305 81
rect 786 78 802 81
rect 1210 78 1226 81
rect 798 74 802 78
rect 1222 74 1226 78
rect 286 68 305 71
rect 454 68 462 71
rect 482 68 494 71
rect 814 71 818 74
rect 814 68 825 71
rect 842 68 849 71
rect 1010 68 1025 71
rect 1042 68 1049 71
rect 1202 68 1203 72
rect 1238 71 1242 74
rect 1238 68 1249 71
rect 1266 68 1273 71
rect 1422 68 1430 71
rect 142 58 150 61
rect 454 58 473 61
rect 642 58 657 61
rect 830 58 849 61
rect 1030 58 1049 61
rect 1254 58 1273 61
rect 1470 61 1473 68
rect 1670 62 1673 71
rect 1974 68 1982 71
rect 1998 68 2006 71
rect 2238 68 2246 71
rect 2270 71 2274 74
rect 2262 68 2274 71
rect 2470 68 2478 71
rect 2518 71 2521 78
rect 2510 68 2521 71
rect 1446 58 1473 61
rect 1974 58 1993 61
rect 2150 58 2166 61
rect 2238 58 2257 61
rect 454 48 457 58
rect 846 48 849 58
rect 1046 48 1049 58
rect 1270 48 1273 58
rect 1454 48 1462 51
rect 1670 48 1689 51
rect 1806 48 1825 51
rect 1834 48 1838 52
rect 1974 48 1977 58
rect 2238 48 2241 58
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
rect 1496 3 1498 7
rect 1502 3 1505 7
rect 1509 3 1512 7
<< m2contact >>
rect 482 2403 486 2407
rect 489 2403 493 2407
rect 1498 2403 1502 2407
rect 1505 2403 1509 2407
rect 886 2388 890 2392
rect 1542 2388 1546 2392
rect 1134 2378 1138 2382
rect 110 2368 114 2372
rect 550 2368 554 2372
rect 702 2368 706 2372
rect 742 2368 746 2372
rect 1262 2368 1266 2372
rect 1614 2368 1618 2372
rect 2054 2368 2058 2372
rect 22 2348 26 2352
rect 70 2348 74 2352
rect 94 2358 98 2362
rect 174 2348 178 2352
rect 294 2348 298 2352
rect 318 2358 322 2362
rect 566 2358 570 2362
rect 574 2358 578 2362
rect 718 2358 722 2362
rect 366 2347 370 2351
rect 518 2347 522 2351
rect 566 2348 570 2352
rect 590 2348 594 2352
rect 638 2348 642 2352
rect 1118 2358 1122 2362
rect 1278 2358 1282 2362
rect 742 2348 746 2352
rect 822 2347 826 2351
rect 854 2348 858 2352
rect 902 2348 906 2352
rect 1046 2348 1050 2352
rect 1102 2348 1106 2352
rect 1110 2348 1114 2352
rect 1198 2348 1202 2352
rect 1302 2348 1306 2352
rect 1326 2348 1330 2352
rect 1350 2358 1354 2362
rect 1422 2348 1426 2352
rect 1470 2348 1474 2352
rect 1518 2348 1522 2352
rect 1558 2348 1562 2352
rect 1566 2348 1570 2352
rect 1598 2358 1602 2362
rect 1918 2358 1922 2362
rect 1934 2358 1938 2362
rect 2070 2358 2074 2362
rect 1678 2348 1682 2352
rect 1782 2347 1786 2351
rect 1846 2348 1850 2352
rect 1918 2348 1922 2352
rect 1990 2348 1994 2352
rect 2206 2358 2210 2362
rect 2086 2348 2090 2352
rect 2094 2348 2098 2352
rect 2134 2347 2138 2351
rect 2262 2348 2266 2352
rect 2358 2348 2362 2352
rect 2470 2348 2474 2352
rect 2494 2358 2498 2362
rect 46 2338 50 2342
rect 62 2338 66 2342
rect 94 2338 98 2342
rect 110 2338 114 2342
rect 214 2338 218 2342
rect 222 2338 226 2342
rect 246 2338 250 2342
rect 286 2338 290 2342
rect 318 2338 322 2342
rect 334 2338 338 2342
rect 374 2338 378 2342
rect 534 2338 538 2342
rect 550 2338 554 2342
rect 598 2338 602 2342
rect 702 2338 706 2342
rect 750 2338 754 2342
rect 838 2338 842 2342
rect 910 2338 914 2342
rect 982 2338 986 2342
rect 1006 2338 1010 2342
rect 1094 2338 1098 2342
rect 1158 2338 1162 2342
rect 1174 2338 1178 2342
rect 1262 2338 1266 2342
rect 1278 2338 1282 2342
rect 1318 2338 1322 2342
rect 1366 2338 1370 2342
rect 1406 2338 1410 2342
rect 1478 2338 1482 2342
rect 1566 2338 1570 2342
rect 1598 2338 1602 2342
rect 1614 2338 1618 2342
rect 1702 2338 1706 2342
rect 1854 2338 1858 2342
rect 1910 2338 1914 2342
rect 1982 2338 1986 2342
rect 2054 2338 2058 2342
rect 2102 2338 2106 2342
rect 2142 2338 2146 2342
rect 2222 2338 2226 2342
rect 2238 2338 2242 2342
rect 2334 2338 2338 2342
rect 2454 2338 2458 2342
rect 2462 2338 2466 2342
rect 2510 2338 2514 2342
rect 6 2328 10 2332
rect 630 2328 634 2332
rect 1534 2328 1538 2332
rect 38 2318 42 2322
rect 270 2318 274 2322
rect 430 2318 434 2322
rect 454 2318 458 2322
rect 758 2318 762 2322
rect 870 2318 874 2322
rect 1086 2318 1090 2322
rect 1134 2318 1138 2322
rect 1342 2318 1346 2322
rect 1462 2318 1466 2322
rect 1486 2318 1490 2322
rect 1718 2318 1722 2322
rect 1902 2318 1906 2322
rect 2198 2318 2202 2322
rect 2214 2318 2218 2322
rect 2318 2318 2322 2322
rect 2414 2318 2418 2322
rect 2446 2318 2450 2322
rect 2486 2318 2490 2322
rect 986 2303 990 2307
rect 993 2303 997 2307
rect 2018 2303 2022 2307
rect 2025 2303 2029 2307
rect 6 2288 10 2292
rect 318 2288 322 2292
rect 518 2288 522 2292
rect 758 2288 762 2292
rect 974 2288 978 2292
rect 1190 2288 1194 2292
rect 1214 2288 1218 2292
rect 1286 2288 1290 2292
rect 1502 2288 1506 2292
rect 1814 2288 1818 2292
rect 1990 2288 1994 2292
rect 2046 2288 2050 2292
rect 1006 2278 1010 2282
rect 1158 2278 1162 2282
rect 1614 2278 1618 2282
rect 1646 2278 1650 2282
rect 1894 2278 1898 2282
rect 86 2268 90 2272
rect 166 2268 170 2272
rect 174 2268 178 2272
rect 198 2268 202 2272
rect 222 2268 226 2272
rect 366 2268 370 2272
rect 406 2268 410 2272
rect 422 2268 426 2272
rect 438 2268 442 2272
rect 574 2268 578 2272
rect 686 2268 690 2272
rect 838 2268 842 2272
rect 854 2268 858 2272
rect 902 2268 906 2272
rect 1038 2268 1042 2272
rect 1070 2268 1074 2272
rect 1102 2268 1106 2272
rect 1150 2268 1154 2272
rect 1198 2268 1202 2272
rect 1230 2268 1234 2272
rect 1238 2268 1242 2272
rect 1366 2268 1370 2272
rect 1382 2268 1386 2272
rect 1414 2268 1418 2272
rect 1582 2268 1586 2272
rect 1606 2268 1610 2272
rect 1758 2268 1762 2272
rect 1958 2268 1962 2272
rect 2014 2268 2018 2272
rect 2038 2268 2042 2272
rect 2102 2268 2106 2272
rect 2214 2268 2218 2272
rect 2254 2268 2258 2272
rect 2286 2268 2290 2272
rect 2390 2268 2394 2272
rect 46 2258 50 2262
rect 182 2258 186 2262
rect 254 2259 258 2263
rect 286 2258 290 2262
rect 326 2258 330 2262
rect 334 2258 338 2262
rect 350 2258 354 2262
rect 358 2258 362 2262
rect 382 2258 386 2262
rect 454 2259 458 2263
rect 542 2258 546 2262
rect 550 2258 554 2262
rect 582 2258 586 2262
rect 590 2258 594 2262
rect 598 2258 602 2262
rect 622 2258 626 2262
rect 638 2258 642 2262
rect 646 2258 650 2262
rect 678 2258 682 2262
rect 750 2258 754 2262
rect 790 2258 794 2262
rect 822 2259 826 2263
rect 870 2258 874 2262
rect 910 2258 914 2262
rect 918 2258 922 2262
rect 942 2258 946 2262
rect 950 2258 954 2262
rect 1030 2258 1034 2262
rect 1078 2258 1082 2262
rect 1094 2258 1098 2262
rect 1150 2258 1154 2262
rect 1174 2258 1178 2262
rect 1206 2258 1210 2262
rect 1270 2258 1274 2262
rect 1278 2258 1282 2262
rect 1350 2259 1354 2263
rect 1390 2258 1394 2262
rect 1446 2258 1450 2262
rect 1470 2258 1474 2262
rect 1486 2258 1490 2262
rect 1550 2258 1554 2262
rect 1598 2258 1602 2262
rect 1630 2258 1634 2262
rect 1750 2259 1754 2263
rect 1822 2258 1826 2262
rect 1830 2258 1834 2262
rect 1862 2258 1866 2262
rect 1878 2258 1882 2262
rect 1902 2258 1906 2262
rect 1910 2258 1914 2262
rect 1918 2258 1922 2262
rect 1926 2258 1930 2262
rect 1950 2258 1954 2262
rect 1974 2258 1978 2262
rect 2086 2259 2090 2263
rect 2158 2258 2162 2262
rect 2166 2258 2170 2262
rect 2190 2258 2194 2262
rect 2206 2258 2210 2262
rect 2238 2258 2242 2262
rect 2246 2258 2250 2262
rect 2262 2258 2266 2262
rect 2302 2258 2306 2262
rect 2366 2258 2370 2262
rect 2438 2258 2442 2262
rect 2470 2259 2474 2263
rect 206 2248 210 2252
rect 406 2248 410 2252
rect 854 2248 858 2252
rect 870 2248 874 2252
rect 878 2248 882 2252
rect 1118 2248 1122 2252
rect 1126 2248 1130 2252
rect 1214 2248 1218 2252
rect 1390 2248 1394 2252
rect 1430 2248 1434 2252
rect 1998 2248 2002 2252
rect 2054 2248 2058 2252
rect 2286 2248 2290 2252
rect 6 2218 10 2222
rect 110 2218 114 2222
rect 614 2218 618 2222
rect 662 2218 666 2222
rect 934 2218 938 2222
rect 1142 2218 1146 2222
rect 1454 2218 1458 2222
rect 1662 2218 1666 2222
rect 1846 2218 1850 2222
rect 1934 2218 1938 2222
rect 2150 2218 2154 2222
rect 2182 2218 2186 2222
rect 2406 2218 2410 2222
rect 482 2203 486 2207
rect 489 2203 493 2207
rect 1498 2203 1502 2207
rect 1505 2203 1509 2207
rect 6 2188 10 2192
rect 454 2188 458 2192
rect 1070 2188 1074 2192
rect 1206 2188 1210 2192
rect 1782 2188 1786 2192
rect 1830 2188 1834 2192
rect 2158 2188 2162 2192
rect 2398 2188 2402 2192
rect 1982 2178 1986 2182
rect 358 2168 362 2172
rect 374 2168 378 2172
rect 702 2168 706 2172
rect 1086 2168 1090 2172
rect 70 2147 74 2151
rect 110 2148 114 2152
rect 118 2148 122 2152
rect 134 2158 138 2162
rect 686 2158 690 2162
rect 918 2158 922 2162
rect 958 2158 962 2162
rect 1022 2158 1026 2162
rect 1078 2158 1082 2162
rect 182 2147 186 2151
rect 254 2148 258 2152
rect 286 2148 290 2152
rect 294 2148 298 2152
rect 302 2148 306 2152
rect 350 2148 354 2152
rect 398 2148 402 2152
rect 414 2148 418 2152
rect 526 2148 530 2152
rect 558 2147 562 2151
rect 622 2148 626 2152
rect 654 2147 658 2151
rect 702 2148 706 2152
rect 718 2148 722 2152
rect 750 2148 754 2152
rect 806 2148 810 2152
rect 846 2148 850 2152
rect 918 2148 922 2152
rect 966 2148 970 2152
rect 998 2148 1002 2152
rect 1014 2148 1018 2152
rect 1046 2148 1050 2152
rect 1062 2148 1066 2152
rect 1142 2148 1146 2152
rect 1246 2148 1250 2152
rect 1262 2148 1266 2152
rect 1310 2148 1314 2152
rect 1334 2158 1338 2162
rect 86 2138 90 2142
rect 102 2138 106 2142
rect 150 2138 154 2142
rect 166 2138 170 2142
rect 342 2138 346 2142
rect 438 2138 442 2142
rect 670 2138 674 2142
rect 710 2138 714 2142
rect 726 2138 730 2142
rect 766 2138 770 2142
rect 782 2138 786 2142
rect 838 2138 842 2142
rect 910 2138 914 2142
rect 942 2138 946 2142
rect 1054 2138 1058 2142
rect 1382 2147 1386 2151
rect 1510 2148 1514 2152
rect 1574 2148 1578 2152
rect 1598 2158 1602 2162
rect 1630 2148 1634 2152
rect 1654 2158 1658 2162
rect 1702 2147 1706 2151
rect 1798 2148 1802 2152
rect 1878 2148 1882 2152
rect 1998 2148 2002 2152
rect 2046 2148 2050 2152
rect 2054 2148 2058 2152
rect 2078 2158 2082 2162
rect 2174 2158 2178 2162
rect 2214 2158 2218 2162
rect 2326 2158 2330 2162
rect 2374 2158 2378 2162
rect 2214 2148 2218 2152
rect 1118 2138 1122 2142
rect 1166 2138 1170 2142
rect 1182 2138 1186 2142
rect 1302 2138 1306 2142
rect 1334 2138 1338 2142
rect 1350 2138 1354 2142
rect 1366 2138 1370 2142
rect 1534 2138 1538 2142
rect 1566 2138 1570 2142
rect 1614 2138 1618 2142
rect 1622 2138 1626 2142
rect 1654 2138 1658 2142
rect 1670 2138 1674 2142
rect 1686 2138 1690 2142
rect 1806 2138 1810 2142
rect 1886 2138 1890 2142
rect 1926 2138 1930 2142
rect 2254 2147 2258 2151
rect 2342 2148 2346 2152
rect 2398 2148 2402 2152
rect 2446 2148 2450 2152
rect 2478 2147 2482 2151
rect 2078 2138 2082 2142
rect 2094 2138 2098 2142
rect 2102 2138 2106 2142
rect 2190 2138 2194 2142
rect 2222 2138 2226 2142
rect 2238 2138 2242 2142
rect 2334 2138 2338 2142
rect 2350 2138 2354 2142
rect 2358 2138 2362 2142
rect 2406 2138 2410 2142
rect 2494 2138 2498 2142
rect 318 2128 322 2132
rect 742 2128 746 2132
rect 246 2118 250 2122
rect 278 2118 282 2122
rect 334 2118 338 2122
rect 494 2118 498 2122
rect 590 2118 594 2122
rect 734 2118 738 2122
rect 902 2118 906 2122
rect 982 2118 986 2122
rect 1030 2118 1034 2122
rect 1198 2118 1202 2122
rect 1446 2118 1450 2122
rect 1454 2118 1458 2122
rect 1590 2118 1594 2122
rect 1766 2118 1770 2122
rect 1822 2118 1826 2122
rect 2318 2118 2322 2122
rect 2414 2118 2418 2122
rect 986 2103 990 2107
rect 993 2103 997 2107
rect 2018 2103 2022 2107
rect 2025 2103 2029 2107
rect 6 2088 10 2092
rect 182 2088 186 2092
rect 566 2088 570 2092
rect 646 2088 650 2092
rect 654 2088 658 2092
rect 758 2088 762 2092
rect 886 2088 890 2092
rect 1022 2088 1026 2092
rect 1030 2088 1034 2092
rect 1190 2088 1194 2092
rect 1222 2088 1226 2092
rect 1286 2088 1290 2092
rect 1414 2088 1418 2092
rect 1446 2088 1450 2092
rect 1470 2088 1474 2092
rect 1598 2088 1602 2092
rect 1798 2088 1802 2092
rect 1814 2088 1818 2092
rect 1942 2088 1946 2092
rect 2022 2088 2026 2092
rect 2318 2088 2322 2092
rect 2326 2088 2330 2092
rect 2486 2088 2490 2092
rect 278 2078 282 2082
rect 574 2078 578 2082
rect 1230 2078 1234 2082
rect 1382 2078 1386 2082
rect 1454 2078 1458 2082
rect 1462 2078 1466 2082
rect 1806 2078 1810 2082
rect 1958 2078 1962 2082
rect 2390 2078 2394 2082
rect 2446 2078 2450 2082
rect 2462 2078 2466 2082
rect 2494 2078 2498 2082
rect 86 2068 90 2072
rect 102 2068 106 2072
rect 150 2068 154 2072
rect 158 2068 162 2072
rect 206 2068 210 2072
rect 358 2068 362 2072
rect 406 2068 410 2072
rect 438 2068 442 2072
rect 550 2068 554 2072
rect 558 2068 562 2072
rect 630 2068 634 2072
rect 750 2068 754 2072
rect 774 2068 778 2072
rect 830 2068 834 2072
rect 1006 2068 1010 2072
rect 1110 2068 1114 2072
rect 1214 2068 1218 2072
rect 1366 2068 1370 2072
rect 1422 2068 1426 2072
rect 1478 2068 1482 2072
rect 1502 2068 1506 2072
rect 1654 2068 1658 2072
rect 1686 2068 1690 2072
rect 1702 2068 1706 2072
rect 1718 2068 1722 2072
rect 1838 2068 1842 2072
rect 1894 2068 1898 2072
rect 1950 2068 1954 2072
rect 1974 2068 1978 2072
rect 1990 2068 1994 2072
rect 2094 2068 2098 2072
rect 2118 2068 2122 2072
rect 2134 2068 2138 2072
rect 2198 2068 2202 2072
rect 2294 2068 2298 2072
rect 2422 2068 2426 2072
rect 2478 2068 2482 2072
rect 70 2059 74 2063
rect 110 2058 114 2062
rect 118 2058 122 2062
rect 166 2058 170 2062
rect 214 2058 218 2062
rect 222 2058 226 2062
rect 294 2058 298 2062
rect 326 2059 330 2063
rect 390 2058 394 2062
rect 406 2058 410 2062
rect 446 2058 450 2062
rect 582 2058 586 2062
rect 614 2058 618 2062
rect 622 2058 626 2062
rect 686 2058 690 2062
rect 718 2059 722 2063
rect 766 2058 770 2062
rect 822 2059 826 2063
rect 894 2058 898 2062
rect 902 2058 906 2062
rect 942 2058 946 2062
rect 950 2058 954 2062
rect 974 2058 978 2062
rect 982 2058 986 2062
rect 1078 2058 1082 2062
rect 1126 2058 1130 2062
rect 1134 2058 1138 2062
rect 1158 2058 1162 2062
rect 1174 2058 1178 2062
rect 1198 2058 1202 2062
rect 1238 2058 1242 2062
rect 1246 2058 1250 2062
rect 1270 2058 1274 2062
rect 1350 2059 1354 2063
rect 1398 2058 1402 2062
rect 1430 2058 1434 2062
rect 1438 2058 1442 2062
rect 1486 2058 1490 2062
rect 1542 2058 1546 2062
rect 1566 2058 1570 2062
rect 1606 2058 1610 2062
rect 1614 2058 1618 2062
rect 1638 2058 1642 2062
rect 1662 2058 1666 2062
rect 1734 2059 1738 2063
rect 1830 2058 1834 2062
rect 1846 2058 1850 2062
rect 1870 2058 1874 2062
rect 1878 2058 1882 2062
rect 1886 2058 1890 2062
rect 1918 2058 1922 2062
rect 1926 2058 1930 2062
rect 1934 2058 1938 2062
rect 1966 2058 1970 2062
rect 1998 2058 2002 2062
rect 2086 2058 2090 2062
rect 2214 2058 2218 2062
rect 2238 2058 2242 2062
rect 2246 2058 2250 2062
rect 2254 2058 2258 2062
rect 2262 2058 2266 2062
rect 2286 2058 2290 2062
rect 2366 2058 2370 2062
rect 2470 2058 2474 2062
rect 134 2048 138 2052
rect 190 2048 194 2052
rect 374 2048 378 2052
rect 510 2048 514 2052
rect 646 2048 650 2052
rect 670 2048 674 2052
rect 790 2048 794 2052
rect 1022 2048 1026 2052
rect 1686 2048 1690 2052
rect 2014 2048 2018 2052
rect 2318 2048 2322 2052
rect 2438 2048 2442 2052
rect 238 2018 242 2022
rect 502 2018 506 2022
rect 606 2018 610 2022
rect 782 2018 786 2022
rect 918 2018 922 2022
rect 958 2018 962 2022
rect 1150 2018 1154 2022
rect 1262 2018 1266 2022
rect 1630 2018 1634 2022
rect 1862 2018 1866 2022
rect 1998 2018 2002 2022
rect 2222 2018 2226 2022
rect 2270 2018 2274 2022
rect 2430 2018 2434 2022
rect 482 2003 486 2007
rect 489 2003 493 2007
rect 1498 2003 1502 2007
rect 1505 2003 1509 2007
rect 630 1988 634 1992
rect 798 1988 802 1992
rect 1030 1988 1034 1992
rect 1758 1988 1762 1992
rect 1838 1988 1842 1992
rect 2486 1988 2490 1992
rect 1734 1978 1738 1982
rect 398 1968 402 1972
rect 414 1968 418 1972
rect 830 1968 834 1972
rect 1598 1968 1602 1972
rect 1614 1968 1618 1972
rect 2206 1968 2210 1972
rect 286 1958 290 1962
rect 46 1948 50 1952
rect 310 1958 314 1962
rect 582 1958 586 1962
rect 126 1947 130 1951
rect 310 1948 314 1952
rect 350 1947 354 1951
rect 446 1948 450 1952
rect 454 1948 458 1952
rect 462 1948 466 1952
rect 486 1948 490 1952
rect 518 1948 522 1952
rect 526 1948 530 1952
rect 550 1948 554 1952
rect 646 1958 650 1962
rect 678 1958 682 1962
rect 694 1958 698 1962
rect 782 1958 786 1962
rect 990 1958 994 1962
rect 1006 1958 1010 1962
rect 1478 1958 1482 1962
rect 1710 1958 1714 1962
rect 606 1948 610 1952
rect 630 1948 634 1952
rect 646 1948 650 1952
rect 686 1948 690 1952
rect 694 1948 698 1952
rect 742 1948 746 1952
rect 774 1948 778 1952
rect 798 1948 802 1952
rect 142 1938 146 1942
rect 262 1938 266 1942
rect 270 1938 274 1942
rect 318 1938 322 1942
rect 334 1938 338 1942
rect 510 1938 514 1942
rect 558 1938 562 1942
rect 590 1938 594 1942
rect 614 1938 618 1942
rect 622 1938 626 1942
rect 654 1938 658 1942
rect 678 1938 682 1942
rect 718 1938 722 1942
rect 878 1947 882 1951
rect 918 1948 922 1952
rect 942 1948 946 1952
rect 950 1948 954 1952
rect 966 1948 970 1952
rect 998 1948 1002 1952
rect 1086 1948 1090 1952
rect 1134 1948 1138 1952
rect 1158 1948 1162 1952
rect 1166 1948 1170 1952
rect 1206 1948 1210 1952
rect 1238 1947 1242 1951
rect 1278 1948 1282 1952
rect 1302 1948 1306 1952
rect 1310 1948 1314 1952
rect 1326 1948 1330 1952
rect 1350 1948 1354 1952
rect 1358 1948 1362 1952
rect 1366 1948 1370 1952
rect 1398 1948 1402 1952
rect 1414 1948 1418 1952
rect 1438 1948 1442 1952
rect 1446 1948 1450 1952
rect 1462 1948 1466 1952
rect 1822 1958 1826 1962
rect 1854 1958 1858 1962
rect 1886 1958 1890 1962
rect 2134 1958 2138 1962
rect 2150 1958 2154 1962
rect 1526 1947 1530 1951
rect 1662 1947 1666 1951
rect 1734 1948 1738 1952
rect 1878 1948 1882 1952
rect 1910 1948 1914 1952
rect 1918 1948 1922 1952
rect 1926 1948 1930 1952
rect 1950 1948 1954 1952
rect 1974 1948 1978 1952
rect 1998 1948 2002 1952
rect 2006 1948 2010 1952
rect 2086 1948 2090 1952
rect 2134 1948 2138 1952
rect 2166 1948 2170 1952
rect 2190 1958 2194 1962
rect 2334 1958 2338 1962
rect 2438 1958 2442 1962
rect 2246 1948 2250 1952
rect 2270 1948 2274 1952
rect 2318 1948 2322 1952
rect 2390 1948 2394 1952
rect 2454 1948 2458 1952
rect 2470 1948 2474 1952
rect 806 1938 810 1942
rect 894 1938 898 1942
rect 958 1938 962 1942
rect 990 1938 994 1942
rect 1110 1938 1114 1942
rect 1270 1938 1274 1942
rect 1318 1938 1322 1942
rect 1374 1938 1378 1942
rect 1454 1938 1458 1942
rect 1486 1938 1490 1942
rect 1534 1938 1538 1942
rect 1558 1938 1562 1942
rect 1678 1938 1682 1942
rect 1694 1938 1698 1942
rect 1742 1938 1746 1942
rect 1814 1938 1818 1942
rect 1846 1938 1850 1942
rect 1870 1938 1874 1942
rect 1886 1938 1890 1942
rect 1902 1938 1906 1942
rect 1958 1938 1962 1942
rect 2094 1938 2098 1942
rect 2126 1938 2130 1942
rect 2158 1938 2162 1942
rect 2190 1938 2194 1942
rect 2206 1938 2210 1942
rect 2294 1938 2298 1942
rect 2310 1938 2314 1942
rect 2334 1938 2338 1942
rect 2462 1938 2466 1942
rect 726 1928 730 1932
rect 1062 1928 1066 1932
rect 1150 1928 1154 1932
rect 2406 1928 2410 1932
rect 6 1918 10 1922
rect 190 1918 194 1922
rect 206 1918 210 1922
rect 430 1918 434 1922
rect 542 1918 546 1922
rect 814 1918 818 1922
rect 926 1918 930 1922
rect 1174 1918 1178 1922
rect 1294 1918 1298 1922
rect 1390 1918 1394 1922
rect 1590 1918 1594 1922
rect 1934 1918 1938 1922
rect 2030 1918 2034 1922
rect 2342 1918 2346 1922
rect 2438 1918 2442 1922
rect 986 1903 990 1907
rect 993 1903 997 1907
rect 2018 1903 2022 1907
rect 2025 1903 2029 1907
rect 86 1888 90 1892
rect 478 1888 482 1892
rect 726 1888 730 1892
rect 846 1888 850 1892
rect 934 1888 938 1892
rect 1334 1888 1338 1892
rect 1446 1888 1450 1892
rect 1470 1888 1474 1892
rect 1526 1888 1530 1892
rect 1582 1888 1586 1892
rect 1662 1888 1666 1892
rect 1870 1888 1874 1892
rect 1902 1888 1906 1892
rect 2006 1888 2010 1892
rect 2030 1888 2034 1892
rect 2150 1888 2154 1892
rect 342 1878 346 1882
rect 406 1878 410 1882
rect 1414 1878 1418 1882
rect 2070 1878 2074 1882
rect 2334 1878 2338 1882
rect 6 1868 10 1872
rect 38 1868 42 1872
rect 62 1868 66 1872
rect 118 1868 122 1872
rect 230 1868 234 1872
rect 398 1868 402 1872
rect 446 1868 450 1872
rect 718 1868 722 1872
rect 742 1868 746 1872
rect 790 1868 794 1872
rect 854 1868 858 1872
rect 878 1868 882 1872
rect 902 1868 906 1872
rect 910 1868 914 1872
rect 958 1868 962 1872
rect 1038 1868 1042 1872
rect 1102 1868 1106 1872
rect 1142 1868 1146 1872
rect 1174 1868 1178 1872
rect 1270 1868 1274 1872
rect 1310 1868 1314 1872
rect 1406 1868 1410 1872
rect 1454 1868 1458 1872
rect 1486 1868 1490 1872
rect 1518 1868 1522 1872
rect 1534 1868 1538 1872
rect 1598 1868 1602 1872
rect 1606 1868 1610 1872
rect 1630 1868 1634 1872
rect 1654 1868 1658 1872
rect 1718 1868 1722 1872
rect 1742 1868 1746 1872
rect 1806 1868 1810 1872
rect 1838 1868 1842 1872
rect 1862 1868 1866 1872
rect 1870 1868 1874 1872
rect 1886 1868 1890 1872
rect 1982 1868 1986 1872
rect 2030 1868 2034 1872
rect 2118 1868 2122 1872
rect 2134 1868 2138 1872
rect 2198 1868 2202 1872
rect 2254 1868 2258 1872
rect 2286 1868 2290 1872
rect 2302 1868 2306 1872
rect 2406 1868 2410 1872
rect 2470 1868 2474 1872
rect 46 1858 50 1862
rect 70 1858 74 1862
rect 110 1858 114 1862
rect 150 1858 154 1862
rect 158 1858 162 1862
rect 246 1858 250 1862
rect 270 1858 274 1862
rect 278 1858 282 1862
rect 294 1858 298 1862
rect 318 1858 322 1862
rect 326 1858 330 1862
rect 422 1858 426 1862
rect 438 1858 442 1862
rect 454 1858 458 1862
rect 510 1858 514 1862
rect 534 1858 538 1862
rect 574 1858 578 1862
rect 582 1858 586 1862
rect 606 1858 610 1862
rect 630 1858 634 1862
rect 638 1858 642 1862
rect 654 1858 658 1862
rect 662 1858 666 1862
rect 670 1858 674 1862
rect 678 1858 682 1862
rect 710 1858 714 1862
rect 718 1858 722 1862
rect 750 1858 754 1862
rect 798 1858 802 1862
rect 894 1858 898 1862
rect 950 1858 954 1862
rect 966 1858 970 1862
rect 998 1858 1002 1862
rect 1014 1858 1018 1862
rect 1062 1858 1066 1862
rect 1182 1858 1186 1862
rect 1190 1858 1194 1862
rect 1206 1858 1210 1862
rect 1262 1858 1266 1862
rect 1318 1858 1322 1862
rect 1430 1858 1434 1862
rect 1462 1858 1466 1862
rect 1510 1858 1514 1862
rect 1542 1858 1546 1862
rect 1550 1858 1554 1862
rect 1582 1858 1586 1862
rect 1702 1858 1706 1862
rect 1758 1858 1762 1862
rect 1766 1858 1770 1862
rect 1790 1858 1794 1862
rect 1814 1858 1818 1862
rect 1862 1858 1866 1862
rect 1894 1858 1898 1862
rect 1958 1858 1962 1862
rect 2078 1858 2082 1862
rect 2158 1858 2162 1862
rect 2166 1858 2170 1862
rect 2206 1858 2210 1862
rect 2214 1858 2218 1862
rect 2238 1858 2242 1862
rect 2246 1858 2250 1862
rect 2262 1858 2266 1862
rect 2334 1859 2338 1863
rect 2502 1858 2506 1862
rect 22 1848 26 1852
rect 94 1848 98 1852
rect 134 1848 138 1852
rect 870 1848 874 1852
rect 926 1848 930 1852
rect 1142 1848 1146 1852
rect 1206 1848 1210 1852
rect 1334 1848 1338 1852
rect 1470 1848 1474 1852
rect 1582 1848 1586 1852
rect 1614 1848 1618 1852
rect 1654 1848 1658 1852
rect 1838 1848 1842 1852
rect 1998 1848 2002 1852
rect 2150 1848 2154 1852
rect 2286 1848 2290 1852
rect 1622 1838 1626 1842
rect 1678 1838 1682 1842
rect 1918 1838 1922 1842
rect 686 1828 690 1832
rect 1774 1828 1778 1832
rect 2398 1828 2402 1832
rect 174 1818 178 1822
rect 254 1818 258 1822
rect 302 1818 306 1822
rect 590 1818 594 1822
rect 982 1818 986 1822
rect 1214 1818 1218 1822
rect 1350 1818 1354 1822
rect 1566 1818 1570 1822
rect 2174 1818 2178 1822
rect 2486 1818 2490 1822
rect 482 1803 486 1807
rect 489 1803 493 1807
rect 1498 1803 1502 1807
rect 1505 1803 1509 1807
rect 534 1788 538 1792
rect 1206 1788 1210 1792
rect 1414 1788 1418 1792
rect 1998 1788 2002 1792
rect 6 1778 10 1782
rect 646 1778 650 1782
rect 326 1768 330 1772
rect 1046 1768 1050 1772
rect 1558 1768 1562 1772
rect 1742 1768 1746 1772
rect 1758 1768 1762 1772
rect 1774 1768 1778 1772
rect 102 1758 106 1762
rect 134 1758 138 1762
rect 174 1758 178 1762
rect 70 1747 74 1751
rect 110 1748 114 1752
rect 190 1748 194 1752
rect 214 1758 218 1762
rect 430 1758 434 1762
rect 526 1758 530 1762
rect 606 1758 610 1762
rect 262 1747 266 1751
rect 286 1748 290 1752
rect 366 1748 370 1752
rect 398 1747 402 1751
rect 438 1748 442 1752
rect 446 1748 450 1752
rect 478 1748 482 1752
rect 486 1748 490 1752
rect 518 1748 522 1752
rect 550 1748 554 1752
rect 582 1748 586 1752
rect 630 1758 634 1762
rect 1158 1758 1162 1762
rect 630 1748 634 1752
rect 702 1748 706 1752
rect 742 1748 746 1752
rect 774 1748 778 1752
rect 782 1748 786 1752
rect 814 1747 818 1751
rect 918 1748 922 1752
rect 926 1748 930 1752
rect 942 1748 946 1752
rect 966 1748 970 1752
rect 974 1748 978 1752
rect 1006 1748 1010 1752
rect 1030 1748 1034 1752
rect 1038 1748 1042 1752
rect 1198 1758 1202 1762
rect 1502 1758 1506 1762
rect 1110 1747 1114 1751
rect 1182 1748 1186 1752
rect 1254 1748 1258 1752
rect 1262 1748 1266 1752
rect 1286 1748 1290 1752
rect 1294 1748 1298 1752
rect 1302 1748 1306 1752
rect 1334 1748 1338 1752
rect 1350 1748 1354 1752
rect 1374 1748 1378 1752
rect 1382 1748 1386 1752
rect 1398 1748 1402 1752
rect 1422 1748 1426 1752
rect 1430 1748 1434 1752
rect 1438 1748 1442 1752
rect 1446 1748 1450 1752
rect 1470 1748 1474 1752
rect 1478 1748 1482 1752
rect 1542 1758 1546 1762
rect 1718 1758 1722 1762
rect 1542 1748 1546 1752
rect 1590 1748 1594 1752
rect 1614 1748 1618 1752
rect 1662 1748 1666 1752
rect 1686 1748 1690 1752
rect 1694 1748 1698 1752
rect 2110 1758 2114 1762
rect 2374 1758 2378 1762
rect 2486 1758 2490 1762
rect 2502 1758 2506 1762
rect 1742 1748 1746 1752
rect 1806 1748 1810 1752
rect 1854 1748 1858 1752
rect 1926 1748 1930 1752
rect 1982 1748 1986 1752
rect 1990 1748 1994 1752
rect 2014 1748 2018 1752
rect 2046 1748 2050 1752
rect 2078 1748 2082 1752
rect 2094 1748 2098 1752
rect 2102 1748 2106 1752
rect 2158 1748 2162 1752
rect 2222 1748 2226 1752
rect 2246 1748 2250 1752
rect 2254 1748 2258 1752
rect 2262 1748 2266 1752
rect 2270 1748 2274 1752
rect 2302 1748 2306 1752
rect 2318 1748 2322 1752
rect 2342 1748 2346 1752
rect 2350 1748 2354 1752
rect 2422 1748 2426 1752
rect 86 1738 90 1742
rect 126 1738 130 1742
rect 134 1738 138 1742
rect 150 1738 154 1742
rect 158 1738 162 1742
rect 182 1738 186 1742
rect 214 1738 218 1742
rect 230 1738 234 1742
rect 246 1738 250 1742
rect 414 1738 418 1742
rect 454 1738 458 1742
rect 526 1738 530 1742
rect 542 1738 546 1742
rect 550 1738 554 1742
rect 566 1738 570 1742
rect 574 1738 578 1742
rect 590 1738 594 1742
rect 638 1738 642 1742
rect 750 1738 754 1742
rect 798 1738 802 1742
rect 886 1738 890 1742
rect 982 1738 986 1742
rect 1086 1738 1090 1742
rect 1126 1738 1130 1742
rect 1142 1738 1146 1742
rect 1158 1738 1162 1742
rect 1190 1738 1194 1742
rect 1214 1738 1218 1742
rect 1310 1738 1314 1742
rect 2446 1747 2450 1751
rect 2486 1748 2490 1752
rect 1486 1738 1490 1742
rect 1550 1738 1554 1742
rect 1654 1738 1658 1742
rect 1702 1738 1706 1742
rect 1750 1738 1754 1742
rect 1838 1738 1842 1742
rect 1918 1738 1922 1742
rect 2054 1738 2058 1742
rect 2070 1738 2074 1742
rect 2086 1738 2090 1742
rect 2214 1738 2218 1742
rect 2310 1738 2314 1742
rect 2358 1738 2362 1742
rect 2478 1738 2482 1742
rect 710 1728 714 1732
rect 1278 1728 1282 1732
rect 2182 1728 2186 1732
rect 2278 1728 2282 1732
rect 174 1718 178 1722
rect 334 1718 338 1722
rect 878 1718 882 1722
rect 950 1718 954 1722
rect 1230 1718 1234 1722
rect 1318 1718 1322 1722
rect 1870 1718 1874 1722
rect 1974 1718 1978 1722
rect 2054 1718 2058 1722
rect 2118 1718 2122 1722
rect 2366 1718 2370 1722
rect 2382 1718 2386 1722
rect 986 1703 990 1707
rect 993 1703 997 1707
rect 2018 1703 2022 1707
rect 2025 1703 2029 1707
rect 166 1688 170 1692
rect 294 1688 298 1692
rect 422 1688 426 1692
rect 510 1688 514 1692
rect 622 1688 626 1692
rect 702 1688 706 1692
rect 878 1688 882 1692
rect 1134 1688 1138 1692
rect 1222 1688 1226 1692
rect 1310 1688 1314 1692
rect 1326 1688 1330 1692
rect 1774 1688 1778 1692
rect 1814 1688 1818 1692
rect 1830 1688 1834 1692
rect 1950 1688 1954 1692
rect 2006 1688 2010 1692
rect 2110 1688 2114 1692
rect 2342 1688 2346 1692
rect 230 1678 234 1682
rect 454 1678 458 1682
rect 558 1678 562 1682
rect 1518 1678 1522 1682
rect 2062 1678 2066 1682
rect 2142 1678 2146 1682
rect 2374 1678 2378 1682
rect 2470 1678 2474 1682
rect 118 1668 122 1672
rect 198 1668 202 1672
rect 302 1668 306 1672
rect 326 1668 330 1672
rect 350 1668 354 1672
rect 502 1668 506 1672
rect 518 1668 522 1672
rect 630 1668 634 1672
rect 678 1668 682 1672
rect 742 1668 746 1672
rect 782 1668 786 1672
rect 814 1668 818 1672
rect 838 1668 842 1672
rect 846 1668 850 1672
rect 862 1668 866 1672
rect 958 1668 962 1672
rect 974 1668 978 1672
rect 1014 1668 1018 1672
rect 1038 1668 1042 1672
rect 1086 1668 1090 1672
rect 1142 1668 1146 1672
rect 1190 1668 1194 1672
rect 1246 1668 1250 1672
rect 1294 1668 1298 1672
rect 1318 1668 1322 1672
rect 1374 1668 1378 1672
rect 1422 1668 1426 1672
rect 1446 1668 1450 1672
rect 1638 1668 1642 1672
rect 1654 1668 1658 1672
rect 1678 1668 1682 1672
rect 1702 1668 1706 1672
rect 1750 1668 1754 1672
rect 1822 1668 1826 1672
rect 1894 1668 1898 1672
rect 1926 1668 1930 1672
rect 1974 1668 1978 1672
rect 2086 1668 2090 1672
rect 2118 1668 2122 1672
rect 2166 1668 2170 1672
rect 2254 1668 2258 1672
rect 2334 1668 2338 1672
rect 2422 1668 2426 1672
rect 2494 1668 2498 1672
rect 110 1658 114 1662
rect 190 1658 194 1662
rect 254 1658 258 1662
rect 342 1658 346 1662
rect 358 1658 362 1662
rect 390 1658 394 1662
rect 398 1658 402 1662
rect 406 1658 410 1662
rect 438 1658 442 1662
rect 462 1658 466 1662
rect 470 1658 474 1662
rect 478 1658 482 1662
rect 526 1658 530 1662
rect 566 1658 570 1662
rect 638 1658 642 1662
rect 686 1658 690 1662
rect 694 1658 698 1662
rect 726 1658 730 1662
rect 734 1658 738 1662
rect 766 1658 770 1662
rect 774 1658 778 1662
rect 790 1658 794 1662
rect 838 1658 842 1662
rect 870 1658 874 1662
rect 942 1659 946 1663
rect 1030 1658 1034 1662
rect 1078 1658 1082 1662
rect 1142 1658 1146 1662
rect 1158 1658 1162 1662
rect 1230 1658 1234 1662
rect 1238 1658 1242 1662
rect 1286 1658 1290 1662
rect 1382 1658 1386 1662
rect 1422 1658 1426 1662
rect 1502 1658 1506 1662
rect 1566 1658 1570 1662
rect 1574 1658 1578 1662
rect 1598 1658 1602 1662
rect 1614 1658 1618 1662
rect 1646 1658 1650 1662
rect 1654 1658 1658 1662
rect 1710 1658 1714 1662
rect 1718 1658 1722 1662
rect 1742 1658 1746 1662
rect 1758 1658 1762 1662
rect 1766 1658 1770 1662
rect 1798 1658 1802 1662
rect 1870 1658 1874 1662
rect 1934 1658 1938 1662
rect 1982 1658 1986 1662
rect 1990 1658 1994 1662
rect 2014 1658 2018 1662
rect 2046 1658 2050 1662
rect 2054 1658 2058 1662
rect 2158 1658 2162 1662
rect 2214 1658 2218 1662
rect 2406 1659 2410 1663
rect 2462 1658 2466 1662
rect 2486 1658 2490 1662
rect 174 1648 178 1652
rect 318 1648 322 1652
rect 422 1648 426 1652
rect 638 1648 642 1652
rect 662 1648 666 1652
rect 814 1648 818 1652
rect 990 1648 994 1652
rect 1174 1648 1178 1652
rect 1262 1648 1266 1652
rect 1286 1648 1290 1652
rect 1302 1648 1306 1652
rect 1446 1648 1450 1652
rect 1686 1648 1690 1652
rect 1806 1648 1810 1652
rect 1958 1648 1962 1652
rect 2094 1648 2098 1652
rect 2110 1648 2114 1652
rect 2134 1648 2138 1652
rect 2470 1648 2474 1652
rect 190 1638 194 1642
rect 382 1638 386 1642
rect 1118 1638 1122 1642
rect 1622 1638 1626 1642
rect 2174 1638 2178 1642
rect 846 1628 850 1632
rect 14 1618 18 1622
rect 166 1618 170 1622
rect 1454 1618 1458 1622
rect 2278 1618 2282 1622
rect 2446 1618 2450 1622
rect 482 1603 486 1607
rect 489 1603 493 1607
rect 1498 1603 1502 1607
rect 1505 1603 1509 1607
rect 366 1588 370 1592
rect 390 1588 394 1592
rect 446 1588 450 1592
rect 518 1588 522 1592
rect 742 1588 746 1592
rect 926 1588 930 1592
rect 1126 1588 1130 1592
rect 1310 1588 1314 1592
rect 1446 1588 1450 1592
rect 1526 1588 1530 1592
rect 1798 1588 1802 1592
rect 2150 1588 2154 1592
rect 102 1568 106 1572
rect 262 1568 266 1572
rect 534 1568 538 1572
rect 814 1568 818 1572
rect 1238 1568 1242 1572
rect 1430 1568 1434 1572
rect 1598 1568 1602 1572
rect 1830 1568 1834 1572
rect 2054 1568 2058 1572
rect 2070 1568 2074 1572
rect 2366 1568 2370 1572
rect 118 1558 122 1562
rect 46 1548 50 1552
rect 134 1548 138 1552
rect 142 1548 146 1552
rect 158 1548 162 1552
rect 190 1548 194 1552
rect 198 1548 202 1552
rect 214 1548 218 1552
rect 238 1558 242 1562
rect 646 1558 650 1562
rect 302 1548 306 1552
rect 358 1548 362 1552
rect 374 1548 378 1552
rect 422 1548 426 1552
rect 454 1548 458 1552
rect 462 1548 466 1552
rect 470 1548 474 1552
rect 494 1548 498 1552
rect 566 1548 570 1552
rect 806 1558 810 1562
rect 1254 1558 1258 1562
rect 598 1547 602 1551
rect 662 1548 666 1552
rect 670 1548 674 1552
rect 766 1548 770 1552
rect 782 1548 786 1552
rect 846 1548 850 1552
rect 870 1548 874 1552
rect 910 1548 914 1552
rect 934 1548 938 1552
rect 966 1548 970 1552
rect 1006 1548 1010 1552
rect 1038 1548 1042 1552
rect 1062 1548 1066 1552
rect 1094 1548 1098 1552
rect 1174 1548 1178 1552
rect 1438 1558 1442 1562
rect 1478 1558 1482 1562
rect 1278 1548 1282 1552
rect 1294 1548 1298 1552
rect 1302 1548 1306 1552
rect 1326 1548 1330 1552
rect 1382 1548 1386 1552
rect 1398 1548 1402 1552
rect 1478 1548 1482 1552
rect 1534 1548 1538 1552
rect 1542 1548 1546 1552
rect 1558 1548 1562 1552
rect 1582 1558 1586 1562
rect 1718 1558 1722 1562
rect 1662 1548 1666 1552
rect 1734 1548 1738 1552
rect 1758 1558 1762 1562
rect 1942 1558 1946 1562
rect 1782 1548 1786 1552
rect 1790 1548 1794 1552
rect 1822 1548 1826 1552
rect 1886 1548 1890 1552
rect 2014 1558 2018 1562
rect 2030 1558 2034 1562
rect 1958 1548 1962 1552
rect 1966 1548 1970 1552
rect 1990 1548 1994 1552
rect 2022 1548 2026 1552
rect 2102 1548 2106 1552
rect 2206 1548 2210 1552
rect 2326 1548 2330 1552
rect 2350 1558 2354 1562
rect 2518 1558 2522 1562
rect 2430 1548 2434 1552
rect 2486 1548 2490 1552
rect 14 1538 18 1542
rect 102 1538 106 1542
rect 150 1538 154 1542
rect 206 1538 210 1542
rect 254 1538 258 1542
rect 342 1538 346 1542
rect 414 1538 418 1542
rect 510 1538 514 1542
rect 550 1538 554 1542
rect 630 1538 634 1542
rect 678 1538 682 1542
rect 686 1538 690 1542
rect 758 1538 762 1542
rect 790 1538 794 1542
rect 894 1538 898 1542
rect 942 1538 946 1542
rect 1014 1538 1018 1542
rect 1070 1538 1074 1542
rect 1134 1538 1138 1542
rect 1150 1538 1154 1542
rect 1238 1538 1242 1542
rect 1254 1538 1258 1542
rect 1286 1538 1290 1542
rect 1374 1538 1378 1542
rect 1454 1538 1458 1542
rect 1462 1538 1466 1542
rect 1550 1538 1554 1542
rect 1582 1538 1586 1542
rect 1598 1538 1602 1542
rect 1686 1538 1690 1542
rect 1702 1538 1706 1542
rect 1726 1538 1730 1542
rect 1750 1538 1754 1542
rect 1774 1538 1778 1542
rect 1894 1538 1898 1542
rect 1926 1538 1930 1542
rect 1982 1538 1986 1542
rect 2014 1538 2018 1542
rect 2046 1538 2050 1542
rect 2134 1538 2138 1542
rect 2230 1538 2234 1542
rect 2246 1538 2250 1542
rect 2318 1538 2322 1542
rect 2350 1538 2354 1542
rect 2366 1538 2370 1542
rect 2454 1538 2458 1542
rect 2486 1538 2490 1542
rect 230 1528 234 1532
rect 374 1528 378 1532
rect 486 1528 490 1532
rect 526 1528 530 1532
rect 998 1528 1002 1532
rect 1054 1528 1058 1532
rect 1110 1528 1114 1532
rect 2470 1528 2474 1532
rect 182 1518 186 1522
rect 366 1518 370 1522
rect 390 1518 394 1522
rect 406 1518 410 1522
rect 950 1518 954 1522
rect 1022 1518 1026 1522
rect 1078 1518 1082 1522
rect 1478 1518 1482 1522
rect 1718 1518 1722 1522
rect 2302 1518 2306 1522
rect 2478 1518 2482 1522
rect 2502 1518 2506 1522
rect 986 1503 990 1507
rect 993 1503 997 1507
rect 2018 1503 2022 1507
rect 2025 1503 2029 1507
rect 334 1488 338 1492
rect 350 1488 354 1492
rect 558 1488 562 1492
rect 798 1488 802 1492
rect 1070 1488 1074 1492
rect 1166 1488 1170 1492
rect 1310 1488 1314 1492
rect 1366 1488 1370 1492
rect 1534 1488 1538 1492
rect 1710 1488 1714 1492
rect 1750 1488 1754 1492
rect 2086 1488 2090 1492
rect 2198 1488 2202 1492
rect 2286 1488 2290 1492
rect 2502 1488 2506 1492
rect 310 1478 314 1482
rect 382 1478 386 1482
rect 502 1478 506 1482
rect 550 1478 554 1482
rect 566 1478 570 1482
rect 742 1478 746 1482
rect 2054 1478 2058 1482
rect 14 1468 18 1472
rect 102 1468 106 1472
rect 118 1468 122 1472
rect 150 1468 154 1472
rect 166 1468 170 1472
rect 254 1468 258 1472
rect 302 1468 306 1472
rect 326 1468 330 1472
rect 438 1468 442 1472
rect 454 1468 458 1472
rect 462 1468 466 1472
rect 518 1468 522 1472
rect 542 1468 546 1472
rect 582 1468 586 1472
rect 686 1468 690 1472
rect 758 1468 762 1472
rect 790 1468 794 1472
rect 862 1468 866 1472
rect 894 1468 898 1472
rect 990 1468 994 1472
rect 1086 1468 1090 1472
rect 1230 1468 1234 1472
rect 1462 1468 1466 1472
rect 38 1458 42 1462
rect 54 1458 58 1462
rect 142 1458 146 1462
rect 198 1458 202 1462
rect 262 1458 266 1462
rect 270 1458 274 1462
rect 374 1458 378 1462
rect 398 1458 402 1462
rect 422 1458 426 1462
rect 430 1458 434 1462
rect 470 1458 474 1462
rect 566 1458 570 1462
rect 678 1458 682 1462
rect 750 1458 754 1462
rect 854 1458 858 1462
rect 958 1458 962 1462
rect 1006 1459 1010 1463
rect 1102 1459 1106 1463
rect 1174 1458 1178 1462
rect 1182 1458 1186 1462
rect 1214 1458 1218 1462
rect 1246 1459 1250 1463
rect 1326 1458 1330 1462
rect 1350 1458 1354 1462
rect 1358 1458 1362 1462
rect 1398 1458 1402 1462
rect 1430 1459 1434 1463
rect 1494 1468 1498 1472
rect 1558 1468 1562 1472
rect 1566 1468 1570 1472
rect 1598 1468 1602 1472
rect 1614 1468 1618 1472
rect 1630 1468 1634 1472
rect 1742 1468 1746 1472
rect 1790 1468 1794 1472
rect 1830 1468 1834 1472
rect 1910 1468 1914 1472
rect 1958 1468 1962 1472
rect 1998 1468 2002 1472
rect 2022 1468 2026 1472
rect 2166 1468 2170 1472
rect 1470 1458 1474 1462
rect 1486 1458 1490 1462
rect 1550 1458 1554 1462
rect 1558 1458 1562 1462
rect 1646 1459 1650 1463
rect 2278 1468 2282 1472
rect 2318 1468 2322 1472
rect 2382 1468 2386 1472
rect 2406 1468 2410 1472
rect 2438 1468 2442 1472
rect 1678 1458 1682 1462
rect 1726 1458 1730 1462
rect 1734 1458 1738 1462
rect 1798 1458 1802 1462
rect 1918 1458 1922 1462
rect 1926 1458 1930 1462
rect 1950 1458 1954 1462
rect 1974 1458 1978 1462
rect 2038 1458 2042 1462
rect 2046 1458 2050 1462
rect 2070 1458 2074 1462
rect 2142 1458 2146 1462
rect 2190 1458 2194 1462
rect 2214 1458 2218 1462
rect 2222 1458 2226 1462
rect 2230 1458 2234 1462
rect 2278 1458 2282 1462
rect 2342 1458 2346 1462
rect 2390 1458 2394 1462
rect 2446 1458 2450 1462
rect 118 1448 122 1452
rect 286 1448 290 1452
rect 326 1448 330 1452
rect 342 1448 346 1452
rect 454 1448 458 1452
rect 478 1448 482 1452
rect 774 1448 778 1452
rect 1510 1448 1514 1452
rect 1534 1448 1538 1452
rect 1598 1448 1602 1452
rect 1718 1448 1722 1452
rect 1998 1448 2002 1452
rect 2246 1448 2250 1452
rect 2270 1448 2274 1452
rect 2406 1448 2410 1452
rect 102 1438 106 1442
rect 246 1418 250 1422
rect 414 1418 418 1422
rect 518 1418 522 1422
rect 534 1418 538 1422
rect 630 1418 634 1422
rect 734 1418 738 1422
rect 1190 1418 1194 1422
rect 1334 1418 1338 1422
rect 1854 1418 1858 1422
rect 1934 1418 1938 1422
rect 482 1403 486 1407
rect 489 1403 493 1407
rect 1498 1403 1502 1407
rect 1505 1403 1509 1407
rect 30 1388 34 1392
rect 358 1388 362 1392
rect 398 1388 402 1392
rect 446 1388 450 1392
rect 694 1388 698 1392
rect 838 1388 842 1392
rect 2406 1388 2410 1392
rect 2438 1388 2442 1392
rect 246 1368 250 1372
rect 1118 1368 1122 1372
rect 1470 1368 1474 1372
rect 1646 1368 1650 1372
rect 2014 1368 2018 1372
rect 2174 1368 2178 1372
rect 2190 1368 2194 1372
rect 78 1348 82 1352
rect 150 1348 154 1352
rect 158 1348 162 1352
rect 174 1358 178 1362
rect 198 1358 202 1362
rect 678 1358 682 1362
rect 710 1358 714 1362
rect 734 1358 738 1362
rect 814 1358 818 1362
rect 214 1348 218 1352
rect 230 1348 234 1352
rect 254 1348 258 1352
rect 270 1348 274 1352
rect 374 1348 378 1352
rect 406 1348 410 1352
rect 414 1348 418 1352
rect 422 1348 426 1352
rect 454 1348 458 1352
rect 478 1348 482 1352
rect 486 1348 490 1352
rect 510 1348 514 1352
rect 582 1348 586 1352
rect 622 1348 626 1352
rect 662 1348 666 1352
rect 694 1348 698 1352
rect 710 1348 714 1352
rect 750 1348 754 1352
rect 758 1348 762 1352
rect 782 1348 786 1352
rect 790 1348 794 1352
rect 838 1348 842 1352
rect 862 1348 866 1352
rect 886 1358 890 1362
rect 1134 1358 1138 1362
rect 6 1338 10 1342
rect 54 1338 58 1342
rect 142 1338 146 1342
rect 190 1338 194 1342
rect 214 1338 218 1342
rect 294 1338 298 1342
rect 302 1338 306 1342
rect 430 1338 434 1342
rect 446 1338 450 1342
rect 518 1338 522 1342
rect 606 1338 610 1342
rect 630 1338 634 1342
rect 646 1338 650 1342
rect 654 1338 658 1342
rect 934 1347 938 1351
rect 958 1348 962 1352
rect 1054 1348 1058 1352
rect 1238 1358 1242 1362
rect 1158 1348 1162 1352
rect 1182 1348 1186 1352
rect 1206 1348 1210 1352
rect 1214 1348 1218 1352
rect 1486 1358 1490 1362
rect 1678 1358 1682 1362
rect 1718 1358 1722 1362
rect 1262 1348 1266 1352
rect 1334 1348 1338 1352
rect 1422 1348 1426 1352
rect 1486 1348 1490 1352
rect 1542 1348 1546 1352
rect 1550 1348 1554 1352
rect 1590 1348 1594 1352
rect 1654 1348 1658 1352
rect 1662 1348 1666 1352
rect 1686 1348 1690 1352
rect 1846 1358 1850 1362
rect 1742 1348 1746 1352
rect 1758 1348 1762 1352
rect 1766 1348 1770 1352
rect 1790 1348 1794 1352
rect 1806 1348 1810 1352
rect 1822 1348 1826 1352
rect 1838 1348 1842 1352
rect 1870 1348 1874 1352
rect 1910 1348 1914 1352
rect 1934 1348 1938 1352
rect 1942 1348 1946 1352
rect 1958 1348 1962 1352
rect 1982 1358 1986 1362
rect 2134 1358 2138 1362
rect 2078 1348 2082 1352
rect 2366 1358 2370 1362
rect 2150 1348 2154 1352
rect 2158 1348 2162 1352
rect 2230 1348 2234 1352
rect 2302 1348 2306 1352
rect 846 1338 850 1342
rect 854 1338 858 1342
rect 886 1338 890 1342
rect 902 1338 906 1342
rect 1046 1338 1050 1342
rect 1118 1338 1122 1342
rect 1134 1338 1138 1342
rect 1166 1338 1170 1342
rect 1222 1338 1226 1342
rect 1270 1338 1274 1342
rect 1382 1338 1386 1342
rect 1470 1338 1474 1342
rect 1566 1338 1570 1342
rect 2334 1347 2338 1351
rect 2374 1348 2378 1352
rect 2382 1348 2386 1352
rect 2422 1348 2426 1352
rect 1718 1338 1722 1342
rect 1750 1338 1754 1342
rect 1830 1338 1834 1342
rect 1862 1338 1866 1342
rect 1886 1338 1890 1342
rect 1894 1338 1898 1342
rect 1950 1338 1954 1342
rect 1982 1338 1986 1342
rect 2014 1338 2018 1342
rect 2070 1338 2074 1342
rect 2102 1338 2106 1342
rect 2118 1338 2122 1342
rect 2166 1338 2170 1342
rect 2254 1338 2258 1342
rect 2494 1338 2498 1342
rect 646 1328 650 1332
rect 1342 1328 1346 1332
rect 134 1318 138 1322
rect 198 1318 202 1322
rect 526 1318 530 1322
rect 766 1318 770 1322
rect 998 1318 1002 1322
rect 1190 1318 1194 1322
rect 1246 1318 1250 1322
rect 1278 1318 1282 1322
rect 1478 1318 1482 1322
rect 1534 1318 1538 1322
rect 1846 1318 1850 1322
rect 2270 1318 2274 1322
rect 2438 1318 2442 1322
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 2018 1303 2022 1307
rect 2025 1303 2029 1307
rect 94 1288 98 1292
rect 278 1288 282 1292
rect 486 1288 490 1292
rect 622 1288 626 1292
rect 742 1288 746 1292
rect 886 1288 890 1292
rect 1022 1288 1026 1292
rect 1294 1288 1298 1292
rect 1502 1288 1506 1292
rect 1846 1288 1850 1292
rect 1910 1288 1914 1292
rect 2006 1288 2010 1292
rect 2366 1288 2370 1292
rect 2414 1288 2418 1292
rect 438 1278 442 1282
rect 446 1278 450 1282
rect 454 1278 458 1282
rect 782 1278 786 1282
rect 1230 1278 1234 1282
rect 1782 1278 1786 1282
rect 2070 1278 2074 1282
rect 2174 1278 2178 1282
rect 2406 1278 2410 1282
rect 14 1268 18 1272
rect 118 1268 122 1272
rect 126 1268 130 1272
rect 150 1268 154 1272
rect 158 1268 162 1272
rect 182 1268 186 1272
rect 214 1268 218 1272
rect 374 1268 378 1272
rect 430 1268 434 1272
rect 470 1268 474 1272
rect 582 1268 586 1272
rect 598 1268 602 1272
rect 646 1268 650 1272
rect 678 1268 682 1272
rect 686 1268 690 1272
rect 814 1268 818 1272
rect 830 1268 834 1272
rect 846 1268 850 1272
rect 862 1268 866 1272
rect 894 1268 898 1272
rect 1006 1268 1010 1272
rect 1022 1268 1026 1272
rect 1038 1268 1042 1272
rect 1102 1268 1106 1272
rect 1150 1268 1154 1272
rect 1182 1268 1186 1272
rect 1198 1268 1202 1272
rect 1342 1268 1346 1272
rect 1382 1268 1386 1272
rect 1398 1268 1402 1272
rect 1422 1268 1426 1272
rect 1454 1268 1458 1272
rect 1470 1268 1474 1272
rect 1542 1268 1546 1272
rect 1582 1268 1586 1272
rect 1598 1268 1602 1272
rect 1614 1268 1618 1272
rect 1646 1268 1650 1272
rect 1702 1268 1706 1272
rect 1726 1268 1730 1272
rect 1750 1268 1754 1272
rect 1910 1268 1914 1272
rect 1926 1268 1930 1272
rect 2086 1268 2090 1272
rect 2102 1268 2106 1272
rect 2118 1268 2122 1272
rect 2150 1268 2154 1272
rect 2222 1268 2226 1272
rect 2254 1268 2258 1272
rect 2342 1268 2346 1272
rect 2358 1268 2362 1272
rect 2390 1268 2394 1272
rect 2406 1268 2410 1272
rect 2454 1268 2458 1272
rect 2494 1268 2498 1272
rect 54 1258 58 1262
rect 142 1258 146 1262
rect 166 1258 170 1262
rect 222 1258 226 1262
rect 286 1258 290 1262
rect 302 1258 306 1262
rect 318 1258 322 1262
rect 326 1258 330 1262
rect 334 1258 338 1262
rect 342 1258 346 1262
rect 366 1258 370 1262
rect 382 1258 386 1262
rect 390 1258 394 1262
rect 422 1258 426 1262
rect 430 1258 434 1262
rect 462 1258 466 1262
rect 494 1258 498 1262
rect 558 1258 562 1262
rect 638 1258 642 1262
rect 654 1258 658 1262
rect 766 1258 770 1262
rect 790 1258 794 1262
rect 798 1258 802 1262
rect 806 1258 810 1262
rect 838 1258 842 1262
rect 870 1258 874 1262
rect 902 1258 906 1262
rect 934 1258 938 1262
rect 942 1258 946 1262
rect 950 1258 954 1262
rect 958 1258 962 1262
rect 982 1258 986 1262
rect 1014 1258 1018 1262
rect 1054 1258 1058 1262
rect 1086 1258 1090 1262
rect 1094 1258 1098 1262
rect 1110 1258 1114 1262
rect 1134 1258 1138 1262
rect 1142 1258 1146 1262
rect 1150 1258 1154 1262
rect 1238 1258 1242 1262
rect 1366 1259 1370 1263
rect 1438 1258 1442 1262
rect 1462 1258 1466 1262
rect 1566 1259 1570 1263
rect 1638 1258 1642 1262
rect 1654 1258 1658 1262
rect 1662 1258 1666 1262
rect 1686 1258 1690 1262
rect 1710 1258 1714 1262
rect 1782 1259 1786 1263
rect 1814 1258 1818 1262
rect 1854 1258 1858 1262
rect 1862 1258 1866 1262
rect 1886 1258 1890 1262
rect 1894 1258 1898 1262
rect 1902 1258 1906 1262
rect 1950 1258 1954 1262
rect 1974 1258 1978 1262
rect 1982 1258 1986 1262
rect 2070 1259 2074 1263
rect 2142 1258 2146 1262
rect 2158 1258 2162 1262
rect 2166 1258 2170 1262
rect 2190 1258 2194 1262
rect 2246 1258 2250 1262
rect 2318 1258 2322 1262
rect 2382 1258 2386 1262
rect 2454 1258 2458 1262
rect 102 1248 106 1252
rect 182 1248 186 1252
rect 614 1248 618 1252
rect 830 1248 834 1252
rect 846 1248 850 1252
rect 1182 1248 1186 1252
rect 1414 1248 1418 1252
rect 1478 1248 1482 1252
rect 1614 1248 1618 1252
rect 1734 1248 1738 1252
rect 2118 1248 2122 1252
rect 2206 1248 2210 1252
rect 2246 1248 2250 1252
rect 2374 1248 2378 1252
rect 2022 1238 2026 1242
rect 2262 1238 2266 1242
rect 742 1218 746 1222
rect 886 1218 890 1222
rect 1302 1218 1306 1222
rect 1670 1218 1674 1222
rect 2414 1218 2418 1222
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 1498 1203 1502 1207
rect 1505 1203 1509 1207
rect 14 1188 18 1192
rect 254 1188 258 1192
rect 702 1188 706 1192
rect 774 1188 778 1192
rect 1102 1188 1106 1192
rect 1350 1188 1354 1192
rect 1782 1188 1786 1192
rect 2390 1178 2394 1182
rect 2494 1178 2498 1182
rect 222 1168 226 1172
rect 478 1168 482 1172
rect 942 1168 946 1172
rect 1718 1168 1722 1172
rect 94 1158 98 1162
rect 278 1158 282 1162
rect 294 1158 298 1162
rect 326 1158 330 1162
rect 430 1158 434 1162
rect 582 1158 586 1162
rect 110 1148 114 1152
rect 126 1148 130 1152
rect 158 1147 162 1151
rect 230 1148 234 1152
rect 238 1148 242 1152
rect 294 1148 298 1152
rect 374 1148 378 1152
rect 430 1148 434 1152
rect 446 1148 450 1152
rect 534 1148 538 1152
rect 582 1148 586 1152
rect 606 1158 610 1162
rect 646 1158 650 1162
rect 742 1158 746 1162
rect 662 1148 666 1152
rect 670 1148 674 1152
rect 678 1148 682 1152
rect 686 1148 690 1152
rect 710 1148 714 1152
rect 750 1148 754 1152
rect 782 1148 786 1152
rect 790 1148 794 1152
rect 806 1148 810 1152
rect 830 1158 834 1162
rect 974 1158 978 1162
rect 990 1158 994 1162
rect 886 1148 890 1152
rect 910 1148 914 1152
rect 1062 1158 1066 1162
rect 1030 1148 1034 1152
rect 1046 1148 1050 1152
rect 1430 1158 1434 1162
rect 1078 1148 1082 1152
rect 1086 1148 1090 1152
rect 1142 1148 1146 1152
rect 1254 1148 1258 1152
rect 1366 1148 1370 1152
rect 1374 1148 1378 1152
rect 1398 1148 1402 1152
rect 1582 1158 1586 1162
rect 1462 1148 1466 1152
rect 1518 1148 1522 1152
rect 70 1138 74 1142
rect 78 1138 82 1142
rect 126 1138 130 1142
rect 174 1138 178 1142
rect 278 1138 282 1142
rect 302 1138 306 1142
rect 342 1138 346 1142
rect 390 1138 394 1142
rect 462 1138 466 1142
rect 542 1138 546 1142
rect 574 1138 578 1142
rect 622 1138 626 1142
rect 726 1138 730 1142
rect 798 1138 802 1142
rect 846 1138 850 1142
rect 950 1138 954 1142
rect 966 1138 970 1142
rect 1046 1138 1050 1142
rect 1094 1138 1098 1142
rect 1182 1138 1186 1142
rect 1230 1138 1234 1142
rect 1294 1138 1298 1142
rect 1406 1138 1410 1142
rect 1550 1147 1554 1151
rect 1598 1148 1602 1152
rect 1646 1148 1650 1152
rect 1718 1148 1722 1152
rect 1742 1158 1746 1162
rect 1862 1158 1866 1162
rect 1870 1158 1874 1162
rect 1766 1148 1770 1152
rect 1774 1148 1778 1152
rect 1814 1148 1818 1152
rect 1838 1148 1842 1152
rect 1910 1148 1914 1152
rect 1934 1148 1938 1152
rect 1958 1158 1962 1162
rect 2198 1158 2202 1162
rect 2214 1158 2218 1162
rect 2398 1158 2402 1162
rect 2038 1148 2042 1152
rect 2126 1148 2130 1152
rect 2198 1148 2202 1152
rect 2222 1148 2226 1152
rect 2246 1148 2250 1152
rect 2254 1148 2258 1152
rect 2262 1148 2266 1152
rect 2286 1148 2290 1152
rect 2302 1148 2306 1152
rect 2310 1148 2314 1152
rect 2334 1148 2338 1152
rect 2350 1148 2354 1152
rect 1470 1138 1474 1142
rect 1566 1138 1570 1142
rect 1606 1138 1610 1142
rect 1622 1138 1626 1142
rect 1710 1138 1714 1142
rect 1758 1138 1762 1142
rect 1822 1138 1826 1142
rect 1846 1138 1850 1142
rect 1886 1138 1890 1142
rect 1918 1138 1922 1142
rect 1950 1138 1954 1142
rect 2062 1138 2066 1142
rect 2102 1138 2106 1142
rect 2150 1138 2154 1142
rect 2190 1138 2194 1142
rect 2430 1147 2434 1151
rect 2382 1138 2386 1142
rect 2414 1138 2418 1142
rect 878 1128 882 1132
rect 1006 1128 1010 1132
rect 2318 1128 2322 1132
rect 14 1118 18 1122
rect 326 1118 330 1122
rect 422 1118 426 1122
rect 742 1118 746 1122
rect 822 1118 826 1122
rect 966 1118 970 1122
rect 1198 1118 1202 1122
rect 1438 1118 1442 1122
rect 1486 1118 1490 1122
rect 1582 1118 1586 1122
rect 1702 1118 1706 1122
rect 1862 1118 1866 1122
rect 1894 1118 1898 1122
rect 1998 1118 2002 1122
rect 2182 1118 2186 1122
rect 2270 1118 2274 1122
rect 2366 1118 2370 1122
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 2018 1103 2022 1107
rect 2025 1103 2029 1107
rect 110 1088 114 1092
rect 134 1088 138 1092
rect 286 1088 290 1092
rect 390 1088 394 1092
rect 454 1088 458 1092
rect 750 1088 754 1092
rect 934 1088 938 1092
rect 1006 1088 1010 1092
rect 1078 1088 1082 1092
rect 1086 1088 1090 1092
rect 1190 1088 1194 1092
rect 1254 1088 1258 1092
rect 1310 1088 1314 1092
rect 1342 1088 1346 1092
rect 1358 1088 1362 1092
rect 1894 1088 1898 1092
rect 2222 1088 2226 1092
rect 2374 1088 2378 1092
rect 2414 1088 2418 1092
rect 2502 1088 2506 1092
rect 814 1078 818 1082
rect 1422 1078 1426 1082
rect 1710 1078 1714 1082
rect 2150 1078 2154 1082
rect 14 1068 18 1072
rect 102 1068 106 1072
rect 182 1068 186 1072
rect 30 1059 34 1063
rect 126 1058 130 1062
rect 198 1059 202 1063
rect 246 1068 250 1072
rect 278 1068 282 1072
rect 342 1068 346 1072
rect 446 1068 450 1072
rect 478 1068 482 1072
rect 558 1068 562 1072
rect 590 1068 594 1072
rect 654 1068 658 1072
rect 662 1068 666 1072
rect 694 1068 698 1072
rect 726 1068 730 1072
rect 942 1068 946 1072
rect 998 1068 1002 1072
rect 1038 1068 1042 1072
rect 1054 1068 1058 1072
rect 1062 1068 1066 1072
rect 1102 1068 1106 1072
rect 1110 1068 1114 1072
rect 1134 1068 1138 1072
rect 1206 1068 1210 1072
rect 1222 1068 1226 1072
rect 1278 1068 1282 1072
rect 1286 1068 1290 1072
rect 1334 1068 1338 1072
rect 1534 1068 1538 1072
rect 1638 1068 1642 1072
rect 1670 1068 1674 1072
rect 230 1058 234 1062
rect 270 1058 274 1062
rect 326 1058 330 1062
rect 494 1058 498 1062
rect 502 1058 506 1062
rect 606 1059 610 1063
rect 678 1058 682 1062
rect 702 1058 706 1062
rect 798 1058 802 1062
rect 870 1059 874 1063
rect 950 1058 954 1062
rect 1270 1058 1274 1062
rect 1422 1059 1426 1063
rect 1518 1058 1522 1062
rect 1542 1058 1546 1062
rect 1566 1058 1570 1062
rect 1574 1058 1578 1062
rect 1598 1058 1602 1062
rect 1614 1058 1618 1062
rect 1646 1058 1650 1062
rect 1710 1068 1714 1072
rect 1726 1068 1730 1072
rect 1742 1068 1746 1072
rect 1822 1068 1826 1072
rect 1886 1068 1890 1072
rect 1974 1068 1978 1072
rect 1998 1068 2002 1072
rect 2014 1068 2018 1072
rect 2022 1068 2026 1072
rect 2094 1068 2098 1072
rect 2118 1068 2122 1072
rect 1686 1058 1690 1062
rect 1814 1058 1818 1062
rect 1878 1058 1882 1062
rect 1942 1058 1946 1062
rect 1990 1058 1994 1062
rect 2006 1058 2010 1062
rect 2030 1058 2034 1062
rect 2054 1058 2058 1062
rect 2078 1058 2082 1062
rect 2086 1058 2090 1062
rect 2102 1058 2106 1062
rect 2150 1059 2154 1063
rect 2318 1068 2322 1072
rect 2438 1068 2442 1072
rect 2446 1068 2450 1072
rect 2238 1058 2242 1062
rect 2246 1058 2250 1062
rect 2254 1058 2258 1062
rect 2278 1058 2282 1062
rect 2294 1058 2298 1062
rect 2390 1058 2394 1062
rect 2430 1058 2434 1062
rect 246 1048 250 1052
rect 454 1048 458 1052
rect 638 1048 642 1052
rect 726 1048 730 1052
rect 966 1048 970 1052
rect 974 1048 978 1052
rect 990 1048 994 1052
rect 1038 1048 1042 1052
rect 1054 1048 1058 1052
rect 1078 1048 1082 1052
rect 1110 1048 1114 1052
rect 1126 1048 1130 1052
rect 1230 1048 1234 1052
rect 1246 1048 1250 1052
rect 1302 1048 1306 1052
rect 1310 1048 1314 1052
rect 1350 1048 1354 1052
rect 1558 1048 1562 1052
rect 1654 1048 1658 1052
rect 1702 1048 1706 1052
rect 1782 1048 1786 1052
rect 1862 1048 1866 1052
rect 2118 1048 2122 1052
rect 2222 1048 2226 1052
rect 2270 1048 2274 1052
rect 2406 1048 2410 1052
rect 1326 1038 1330 1042
rect 1622 1038 1626 1042
rect 2198 1038 2202 1042
rect 2310 1038 2314 1042
rect 1710 1028 1714 1032
rect 94 1018 98 1022
rect 110 1018 114 1022
rect 134 1018 138 1022
rect 510 1018 514 1022
rect 950 1018 954 1022
rect 982 1018 986 1022
rect 1094 1018 1098 1022
rect 1214 1018 1218 1022
rect 1294 1018 1298 1022
rect 1318 1018 1322 1022
rect 1878 1018 1882 1022
rect 2214 1018 2218 1022
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 1498 1003 1502 1007
rect 1505 1003 1509 1007
rect 22 988 26 992
rect 478 988 482 992
rect 838 988 842 992
rect 934 988 938 992
rect 950 988 954 992
rect 1166 988 1170 992
rect 1342 988 1346 992
rect 1366 988 1370 992
rect 1398 988 1402 992
rect 1470 988 1474 992
rect 1550 988 1554 992
rect 1790 988 1794 992
rect 2110 988 2114 992
rect 2150 988 2154 992
rect 2486 988 2490 992
rect 126 968 130 972
rect 606 968 610 972
rect 1126 968 1130 972
rect 6 958 10 962
rect 198 958 202 962
rect 22 948 26 952
rect 70 948 74 952
rect 134 948 138 952
rect 166 948 170 952
rect 174 948 178 952
rect 182 948 186 952
rect 254 958 258 962
rect 222 948 226 952
rect 318 958 322 962
rect 422 958 426 962
rect 678 958 682 962
rect 278 948 282 952
rect 302 948 306 952
rect 30 938 34 942
rect 350 947 354 951
rect 438 948 442 952
rect 454 948 458 952
rect 462 948 466 952
rect 510 948 514 952
rect 550 948 554 952
rect 614 948 618 952
rect 622 948 626 952
rect 646 948 650 952
rect 742 958 746 962
rect 942 958 946 962
rect 966 958 970 962
rect 1022 958 1026 962
rect 1150 958 1154 962
rect 1174 958 1178 962
rect 1910 958 1914 962
rect 702 948 706 952
rect 710 948 714 952
rect 734 948 738 952
rect 774 947 778 951
rect 894 948 898 952
rect 1030 948 1034 952
rect 1062 947 1066 951
rect 1158 948 1162 952
rect 1190 948 1194 952
rect 1214 948 1218 952
rect 1222 948 1226 952
rect 1350 948 1354 952
rect 1382 948 1386 952
rect 1414 948 1418 952
rect 1454 948 1458 952
rect 1510 948 1514 952
rect 1534 948 1538 952
rect 1566 948 1570 952
rect 1574 948 1578 952
rect 1582 948 1586 952
rect 1646 948 1650 952
rect 1734 948 1738 952
rect 1758 948 1762 952
rect 1830 948 1834 952
rect 2062 958 2066 962
rect 2142 958 2146 962
rect 2262 958 2266 962
rect 1862 947 1866 951
rect 1934 948 1938 952
rect 1982 948 1986 952
rect 2014 947 2018 951
rect 2046 948 2050 952
rect 2078 948 2082 952
rect 2094 948 2098 952
rect 2102 948 2106 952
rect 2126 948 2130 952
rect 2198 948 2202 952
rect 2230 947 2234 951
rect 2262 948 2266 952
rect 2286 948 2290 952
rect 2302 948 2306 952
rect 2326 958 2330 962
rect 2446 958 2450 962
rect 198 938 202 942
rect 230 938 234 942
rect 238 938 242 942
rect 294 938 298 942
rect 318 938 322 942
rect 430 938 434 942
rect 446 938 450 942
rect 526 938 530 942
rect 654 938 658 942
rect 686 938 690 942
rect 710 938 714 942
rect 718 938 722 942
rect 758 938 762 942
rect 878 938 882 942
rect 966 938 970 942
rect 998 938 1002 942
rect 1030 938 1034 942
rect 1134 938 1138 942
rect 1150 938 1154 942
rect 1246 940 1250 944
rect 1254 938 1258 942
rect 1262 938 1266 942
rect 1334 938 1338 942
rect 1486 938 1490 942
rect 1894 938 1898 942
rect 1910 938 1914 942
rect 1942 938 1946 942
rect 2086 938 2090 942
rect 2158 938 2162 942
rect 2374 947 2378 951
rect 2470 948 2474 952
rect 2478 948 2482 952
rect 2510 948 2514 952
rect 2294 938 2298 942
rect 2318 938 2322 942
rect 2342 938 2346 942
rect 2358 938 2362 942
rect 2462 938 2466 942
rect 62 928 66 932
rect 158 928 162 932
rect 350 928 354 932
rect 382 928 386 932
rect 1062 928 1066 932
rect 1398 928 1402 932
rect 1598 928 1602 932
rect 262 918 266 922
rect 414 918 418 922
rect 638 918 642 922
rect 950 918 954 922
rect 1166 918 1170 922
rect 1206 918 1210 922
rect 1230 918 1234 922
rect 1318 918 1322 922
rect 1366 918 1370 922
rect 1430 918 1434 922
rect 1470 918 1474 922
rect 1590 918 1594 922
rect 1798 918 1802 922
rect 1950 918 1954 922
rect 2166 918 2170 922
rect 2438 918 2442 922
rect 2446 918 2450 922
rect 986 903 990 907
rect 993 903 997 907
rect 2018 903 2022 907
rect 2025 903 2029 907
rect 62 888 66 892
rect 78 888 82 892
rect 198 888 202 892
rect 342 888 346 892
rect 422 888 426 892
rect 454 888 458 892
rect 654 888 658 892
rect 830 888 834 892
rect 846 888 850 892
rect 902 888 906 892
rect 958 888 962 892
rect 966 888 970 892
rect 1022 888 1026 892
rect 1046 888 1050 892
rect 1142 888 1146 892
rect 1310 888 1314 892
rect 1406 888 1410 892
rect 1590 888 1594 892
rect 1710 888 1714 892
rect 1958 888 1962 892
rect 2046 888 2050 892
rect 2206 888 2210 892
rect 2406 888 2410 892
rect 2454 888 2458 892
rect 1078 878 1082 882
rect 1598 878 1602 882
rect 1654 878 1658 882
rect 6 868 10 872
rect 94 868 98 872
rect 110 868 114 872
rect 358 868 362 872
rect 406 868 410 872
rect 414 868 418 872
rect 534 868 538 872
rect 550 868 554 872
rect 574 868 578 872
rect 606 868 610 872
rect 734 868 738 872
rect 750 868 754 872
rect 814 868 818 872
rect 846 868 850 872
rect 862 868 866 872
rect 894 868 898 872
rect 942 868 946 872
rect 1006 868 1010 872
rect 1030 868 1034 872
rect 1150 868 1154 872
rect 1198 868 1202 872
rect 1254 868 1258 872
rect 1302 868 1306 872
rect 1486 868 1490 872
rect 1510 868 1514 872
rect 1534 868 1538 872
rect 1582 868 1586 872
rect 1678 868 1682 872
rect 1694 868 1698 872
rect 1758 868 1762 872
rect 1950 868 1954 872
rect 1974 868 1978 872
rect 2022 868 2026 872
rect 2126 868 2130 872
rect 2190 868 2194 872
rect 2262 868 2266 872
rect 2310 868 2314 872
rect 2326 868 2330 872
rect 2414 868 2418 872
rect 2510 868 2514 872
rect 142 858 146 862
rect 150 858 154 862
rect 230 858 234 862
rect 262 859 266 863
rect 302 858 306 862
rect 326 858 330 862
rect 334 858 338 862
rect 366 858 370 862
rect 374 858 378 862
rect 494 858 498 862
rect 558 858 562 862
rect 614 858 618 862
rect 638 858 642 862
rect 646 858 650 862
rect 702 858 706 862
rect 78 848 82 852
rect 342 848 346 852
rect 438 848 442 852
rect 918 858 922 862
rect 1102 858 1106 862
rect 1158 858 1162 862
rect 1166 858 1170 862
rect 1206 858 1210 862
rect 1214 858 1218 862
rect 1246 858 1250 862
rect 1262 858 1266 862
rect 1270 858 1274 862
rect 1342 858 1346 862
rect 1350 858 1354 862
rect 1470 859 1474 863
rect 1558 858 1562 862
rect 1574 858 1578 862
rect 1606 858 1610 862
rect 1638 858 1642 862
rect 1646 858 1650 862
rect 1670 858 1674 862
rect 1702 858 1706 862
rect 1766 858 1770 862
rect 1806 858 1810 862
rect 1822 858 1826 862
rect 1838 858 1842 862
rect 1846 858 1850 862
rect 1854 858 1858 862
rect 1862 858 1866 862
rect 1886 858 1890 862
rect 1902 858 1906 862
rect 1910 858 1914 862
rect 2030 858 2034 862
rect 2102 858 2106 862
rect 2142 858 2146 862
rect 2150 858 2154 862
rect 2174 858 2178 862
rect 2182 858 2186 862
rect 2214 858 2218 862
rect 2222 858 2226 862
rect 2302 858 2306 862
rect 2342 859 2346 863
rect 2422 858 2426 862
rect 2438 858 2442 862
rect 582 848 586 852
rect 822 848 826 852
rect 846 848 850 852
rect 870 848 874 852
rect 886 848 890 852
rect 918 848 922 852
rect 958 848 962 852
rect 966 848 970 852
rect 1022 848 1026 852
rect 1046 848 1050 852
rect 1182 848 1186 852
rect 1286 848 1290 852
rect 1534 848 1538 852
rect 1966 848 1970 852
rect 1990 848 1994 852
rect 2014 848 2018 852
rect 2206 848 2210 852
rect 2278 848 2282 852
rect 2302 848 2306 852
rect 2438 848 2442 852
rect 190 838 194 842
rect 670 838 674 842
rect 910 838 914 842
rect 318 818 322 822
rect 630 818 634 822
rect 830 818 834 822
rect 926 818 930 822
rect 974 818 978 822
rect 1014 818 1018 822
rect 1038 818 1042 822
rect 1222 818 1226 822
rect 1630 818 1634 822
rect 1878 818 1882 822
rect 1926 818 1930 822
rect 2238 818 2242 822
rect 482 803 486 807
rect 489 803 493 807
rect 1498 803 1502 807
rect 1505 803 1509 807
rect 710 788 714 792
rect 950 788 954 792
rect 1078 788 1082 792
rect 1398 788 1402 792
rect 1414 788 1418 792
rect 1638 788 1642 792
rect 2006 788 2010 792
rect 102 768 106 772
rect 438 768 442 772
rect 566 768 570 772
rect 582 768 586 772
rect 1478 768 1482 772
rect 1574 768 1578 772
rect 1950 768 1954 772
rect 2254 768 2258 772
rect 30 747 34 751
rect 62 748 66 752
rect 118 748 122 752
rect 126 748 130 752
rect 158 748 162 752
rect 190 748 194 752
rect 198 748 202 752
rect 214 758 218 762
rect 238 748 242 752
rect 270 748 274 752
rect 302 748 306 752
rect 326 758 330 762
rect 374 747 378 751
rect 446 748 450 752
rect 454 748 458 752
rect 494 748 498 752
rect 526 748 530 752
rect 542 748 546 752
rect 558 748 562 752
rect 622 748 626 752
rect 686 748 690 752
rect 734 748 738 752
rect 742 748 746 752
rect 758 758 762 762
rect 934 758 938 762
rect 942 758 946 762
rect 982 758 986 762
rect 814 748 818 752
rect 878 748 882 752
rect 910 748 914 752
rect 1086 758 1090 762
rect 1126 758 1130 762
rect 1206 758 1210 762
rect 1422 758 1426 762
rect 1022 748 1026 752
rect 1046 748 1050 752
rect 1094 748 1098 752
rect 1110 748 1114 752
rect 1150 748 1154 752
rect 1174 748 1178 752
rect 1182 748 1186 752
rect 1230 748 1234 752
rect 1238 748 1242 752
rect 1270 748 1274 752
rect 1278 748 1282 752
rect 1286 748 1290 752
rect 1326 748 1330 752
rect 1334 748 1338 752
rect 1350 748 1354 752
rect 1366 748 1370 752
rect 1382 748 1386 752
rect 1430 748 1434 752
rect 1518 748 1522 752
rect 1542 747 1546 751
rect 1614 748 1618 752
rect 1654 748 1658 752
rect 1662 748 1666 752
rect 1678 748 1682 752
rect 1694 758 1698 762
rect 1814 758 1818 762
rect 1742 747 1746 751
rect 1830 748 1834 752
rect 1846 748 1850 752
rect 1854 748 1858 752
rect 1886 748 1890 752
rect 1894 748 1898 752
rect 1902 748 1906 752
rect 1926 748 1930 752
rect 1942 748 1946 752
rect 1974 758 1978 762
rect 2014 758 2018 762
rect 2046 758 2050 762
rect 2142 758 2146 762
rect 2150 758 2154 762
rect 2166 758 2170 762
rect 2198 758 2202 762
rect 2478 758 2482 762
rect 2038 748 2042 752
rect 2070 748 2074 752
rect 2078 748 2082 752
rect 2086 748 2090 752
rect 2118 748 2122 752
rect 2198 748 2202 752
rect 2238 748 2242 752
rect 2246 748 2250 752
rect 2294 748 2298 752
rect 2438 748 2442 752
rect 2470 748 2474 752
rect 2518 748 2522 752
rect 134 738 138 742
rect 182 738 186 742
rect 230 738 234 742
rect 246 738 250 742
rect 294 738 298 742
rect 326 738 330 742
rect 342 738 346 742
rect 358 738 362 742
rect 478 738 482 742
rect 550 738 554 742
rect 646 738 650 742
rect 774 738 778 742
rect 806 738 810 742
rect 886 738 890 742
rect 902 738 906 742
rect 918 738 922 742
rect 958 738 962 742
rect 966 738 970 742
rect 1030 738 1034 742
rect 1038 738 1042 742
rect 1070 738 1074 742
rect 1086 738 1090 742
rect 1190 738 1194 742
rect 1246 738 1250 742
rect 1294 738 1298 742
rect 1310 738 1314 742
rect 1318 738 1322 742
rect 1374 738 1378 742
rect 1406 738 1410 742
rect 1470 738 1474 742
rect 1574 738 1578 742
rect 1590 738 1594 742
rect 1606 738 1610 742
rect 1662 738 1666 742
rect 1710 738 1714 742
rect 1726 738 1730 742
rect 1838 738 1842 742
rect 1878 738 1882 742
rect 1934 738 1938 742
rect 1990 738 1994 742
rect 1998 738 2002 742
rect 2022 738 2026 742
rect 2062 738 2066 742
rect 2126 738 2130 742
rect 2150 738 2154 742
rect 2174 738 2178 742
rect 2198 738 2202 742
rect 2206 738 2210 742
rect 2350 738 2354 742
rect 2462 738 2466 742
rect 2502 738 2506 742
rect 174 728 178 732
rect 286 728 290 732
rect 494 728 498 732
rect 1118 728 1122 732
rect 1134 728 1138 732
rect 1230 728 1234 732
rect 1622 728 1626 732
rect 1814 728 1818 732
rect 2318 728 2322 732
rect 2422 728 2426 732
rect 94 718 98 722
rect 142 718 146 722
rect 254 718 258 722
rect 670 718 674 722
rect 870 718 874 722
rect 894 718 898 722
rect 926 718 930 722
rect 1006 718 1010 722
rect 1062 718 1066 722
rect 1086 718 1090 722
rect 1158 718 1162 722
rect 1294 718 1298 722
rect 1414 718 1418 722
rect 1806 718 1810 722
rect 1910 718 1914 722
rect 2094 718 2098 722
rect 2134 718 2138 722
rect 2406 718 2410 722
rect 2454 718 2458 722
rect 2478 718 2482 722
rect 986 703 990 707
rect 993 703 997 707
rect 2018 703 2022 707
rect 2025 703 2029 707
rect 30 688 34 692
rect 198 688 202 692
rect 966 688 970 692
rect 1094 688 1098 692
rect 1110 688 1114 692
rect 1190 688 1194 692
rect 1598 688 1602 692
rect 1838 688 1842 692
rect 1846 688 1850 692
rect 1934 688 1938 692
rect 1974 688 1978 692
rect 2110 688 2114 692
rect 2158 688 2162 692
rect 2326 688 2330 692
rect 2510 688 2514 692
rect 662 678 666 682
rect 782 678 786 682
rect 958 678 962 682
rect 1062 678 1066 682
rect 1158 678 1162 682
rect 1390 678 1394 682
rect 1718 678 1722 682
rect 1774 678 1778 682
rect 1894 678 1898 682
rect 2030 678 2034 682
rect 2358 678 2362 682
rect 6 668 10 672
rect 54 668 58 672
rect 118 668 122 672
rect 150 668 154 672
rect 214 668 218 672
rect 334 668 338 672
rect 398 668 402 672
rect 518 668 522 672
rect 534 668 538 672
rect 558 668 562 672
rect 574 668 578 672
rect 590 668 594 672
rect 654 668 658 672
rect 670 668 674 672
rect 686 668 690 672
rect 766 668 770 672
rect 782 668 786 672
rect 46 658 50 662
rect 62 658 66 662
rect 78 658 82 662
rect 94 658 98 662
rect 102 658 106 662
rect 142 658 146 662
rect 254 658 258 662
rect 262 658 266 662
rect 302 658 306 662
rect 310 658 314 662
rect 342 658 346 662
rect 350 658 354 662
rect 358 658 362 662
rect 382 658 386 662
rect 406 658 410 662
rect 414 658 418 662
rect 430 658 434 662
rect 446 658 450 662
rect 454 658 458 662
rect 462 658 466 662
rect 478 658 482 662
rect 502 658 506 662
rect 510 658 514 662
rect 542 658 546 662
rect 550 658 554 662
rect 582 658 586 662
rect 622 658 626 662
rect 638 658 642 662
rect 678 658 682 662
rect 710 658 714 662
rect 718 658 722 662
rect 742 658 746 662
rect 750 658 754 662
rect 758 658 762 662
rect 790 658 794 662
rect 806 658 810 662
rect 814 658 818 662
rect 830 668 834 672
rect 854 668 858 672
rect 894 668 898 672
rect 910 668 914 672
rect 926 668 930 672
rect 1046 668 1050 672
rect 1078 668 1082 672
rect 1094 668 1098 672
rect 1142 668 1146 672
rect 1158 668 1162 672
rect 1174 668 1178 672
rect 1286 668 1290 672
rect 1310 668 1314 672
rect 1334 668 1338 672
rect 1350 668 1354 672
rect 1518 668 1522 672
rect 1630 668 1634 672
rect 1662 668 1666 672
rect 1670 668 1674 672
rect 1686 668 1690 672
rect 1862 668 1866 672
rect 1926 668 1930 672
rect 1942 668 1946 672
rect 2022 668 2026 672
rect 2046 668 2050 672
rect 2054 668 2058 672
rect 2126 668 2130 672
rect 862 658 866 662
rect 886 658 890 662
rect 902 658 906 662
rect 918 658 922 662
rect 1006 658 1010 662
rect 1070 658 1074 662
rect 1126 658 1130 662
rect 1150 658 1154 662
rect 1182 658 1186 662
rect 1222 658 1226 662
rect 1254 659 1258 663
rect 1326 658 1330 662
rect 1366 658 1370 662
rect 1374 658 1378 662
rect 1422 659 1426 663
rect 2238 668 2242 672
rect 2254 668 2258 672
rect 2302 668 2306 672
rect 2406 668 2410 672
rect 1446 658 1450 662
rect 1558 658 1562 662
rect 1646 658 1650 662
rect 1654 658 1658 662
rect 1678 658 1682 662
rect 1694 658 1698 662
rect 1702 658 1706 662
rect 1710 658 1714 662
rect 1734 658 1738 662
rect 1790 658 1794 662
rect 1878 658 1882 662
rect 1902 658 1906 662
rect 1910 658 1914 662
rect 1918 658 1922 662
rect 1950 658 1954 662
rect 1958 658 1962 662
rect 1990 658 1994 662
rect 1998 658 2002 662
rect 2006 658 2010 662
rect 2054 658 2058 662
rect 2094 658 2098 662
rect 2134 658 2138 662
rect 2150 658 2154 662
rect 2206 658 2210 662
rect 2262 658 2266 662
rect 2286 658 2290 662
rect 2294 658 2298 662
rect 2390 659 2394 663
rect 2454 658 2458 662
rect 22 648 26 652
rect 606 648 610 652
rect 638 648 642 652
rect 686 648 690 652
rect 798 648 802 652
rect 846 648 850 652
rect 942 648 946 652
rect 1094 648 1098 652
rect 1118 648 1122 652
rect 1126 648 1130 652
rect 1302 648 1306 652
rect 1622 648 1626 652
rect 1846 648 1850 652
rect 2150 648 2154 652
rect 2318 648 2322 652
rect 294 638 298 642
rect 518 638 522 642
rect 574 638 578 642
rect 622 618 626 622
rect 726 618 730 622
rect 878 618 882 622
rect 966 618 970 622
rect 1486 618 1490 622
rect 2310 618 2314 622
rect 482 603 486 607
rect 489 603 493 607
rect 1498 603 1502 607
rect 1505 603 1509 607
rect 430 588 434 592
rect 470 588 474 592
rect 542 588 546 592
rect 846 588 850 592
rect 894 588 898 592
rect 1158 588 1162 592
rect 1230 588 1234 592
rect 1398 588 1402 592
rect 1950 588 1954 592
rect 2062 588 2066 592
rect 2278 588 2282 592
rect 2406 588 2410 592
rect 150 578 154 582
rect 254 568 258 572
rect 774 568 778 572
rect 990 568 994 572
rect 1182 568 1186 572
rect 22 558 26 562
rect 270 558 274 562
rect 38 548 42 552
rect 46 548 50 552
rect 86 547 90 551
rect 190 548 194 552
rect 294 548 298 552
rect 366 548 370 552
rect 414 548 418 552
rect 438 548 442 552
rect 446 548 450 552
rect 454 548 458 552
rect 462 548 466 552
rect 486 548 490 552
rect 518 548 522 552
rect 526 548 530 552
rect 550 548 554 552
rect 566 548 570 552
rect 622 548 626 552
rect 638 548 642 552
rect 662 558 666 562
rect 1102 558 1106 562
rect 710 547 714 551
rect 790 548 794 552
rect 798 548 802 552
rect 814 548 818 552
rect 822 548 826 552
rect 838 548 842 552
rect 862 548 866 552
rect 870 548 874 552
rect 878 548 882 552
rect 886 548 890 552
rect 910 548 914 552
rect 926 548 930 552
rect 934 548 938 552
rect 950 548 954 552
rect 966 548 970 552
rect 1166 558 1170 562
rect 1254 558 1258 562
rect 1054 547 1058 551
rect 1126 548 1130 552
rect 1206 548 1210 552
rect 1214 548 1218 552
rect 1238 548 1242 552
rect 1278 548 1282 552
rect 1294 548 1298 552
rect 1334 547 1338 551
rect 1406 548 1410 552
rect 1438 548 1442 552
rect 1462 548 1466 552
rect 1494 548 1498 552
rect 1502 548 1506 552
rect 1534 548 1538 552
rect 1558 558 1562 562
rect 2374 558 2378 562
rect 1606 547 1610 551
rect 1734 548 1738 552
rect 1822 548 1826 552
rect 1870 548 1874 552
rect 1894 548 1898 552
rect 6 538 10 542
rect 54 538 58 542
rect 70 538 74 542
rect 166 538 170 542
rect 254 538 258 542
rect 278 538 282 542
rect 302 538 306 542
rect 390 538 394 542
rect 574 538 578 542
rect 614 538 618 542
rect 630 538 634 542
rect 662 538 666 542
rect 678 538 682 542
rect 694 538 698 542
rect 1070 538 1074 542
rect 1086 538 1090 542
rect 1102 538 1106 542
rect 1134 538 1138 542
rect 1182 538 1186 542
rect 1270 538 1274 542
rect 1302 538 1306 542
rect 1414 538 1418 542
rect 1462 538 1466 542
rect 1526 538 1530 542
rect 1550 538 1554 542
rect 1574 538 1578 542
rect 1590 538 1594 542
rect 1742 538 1746 542
rect 1806 538 1810 542
rect 1886 538 1890 542
rect 1918 548 1922 552
rect 1958 548 1962 552
rect 1966 548 1970 552
rect 1990 548 1994 552
rect 2030 548 2034 552
rect 2038 548 2042 552
rect 2142 548 2146 552
rect 2182 548 2186 552
rect 2214 547 2218 551
rect 2270 548 2274 552
rect 2310 548 2314 552
rect 2342 547 2346 551
rect 2382 548 2386 552
rect 2390 548 2394 552
rect 2470 547 2474 551
rect 1910 538 1914 542
rect 2014 538 2018 542
rect 2078 538 2082 542
rect 2246 538 2250 542
rect 2262 538 2266 542
rect 2398 538 2402 542
rect 2462 538 2466 542
rect 598 528 602 532
rect 1142 528 1146 532
rect 1198 528 1202 532
rect 1334 528 1338 532
rect 1454 528 1458 532
rect 1870 528 1874 532
rect 1918 528 1922 532
rect 1974 528 1978 532
rect 2246 528 2250 532
rect 310 518 314 522
rect 582 518 586 522
rect 606 518 610 522
rect 1422 518 1426 522
rect 1670 518 1674 522
rect 1678 518 1682 522
rect 1862 518 1866 522
rect 2006 518 2010 522
rect 2150 518 2154 522
rect 986 503 990 507
rect 993 503 997 507
rect 2018 503 2022 507
rect 2025 503 2029 507
rect 38 488 42 492
rect 246 488 250 492
rect 278 488 282 492
rect 326 488 330 492
rect 462 488 466 492
rect 510 488 514 492
rect 702 488 706 492
rect 854 488 858 492
rect 918 488 922 492
rect 1094 488 1098 492
rect 1358 488 1362 492
rect 1494 488 1498 492
rect 1526 488 1530 492
rect 1582 488 1586 492
rect 1622 488 1626 492
rect 1686 488 1690 492
rect 1758 488 1762 492
rect 1902 488 1906 492
rect 1926 488 1930 492
rect 2054 488 2058 492
rect 2086 488 2090 492
rect 2246 488 2250 492
rect 2278 488 2282 492
rect 2502 488 2506 492
rect 1126 478 1130 482
rect 1382 478 1386 482
rect 2238 478 2242 482
rect 94 468 98 472
rect 102 468 106 472
rect 150 468 154 472
rect 166 468 170 472
rect 302 468 306 472
rect 350 468 354 472
rect 454 468 458 472
rect 494 468 498 472
rect 598 468 602 472
rect 622 468 626 472
rect 710 468 714 472
rect 726 468 730 472
rect 758 468 762 472
rect 774 468 778 472
rect 878 468 882 472
rect 910 468 914 472
rect 998 468 1002 472
rect 1014 468 1018 472
rect 1046 468 1050 472
rect 1078 468 1082 472
rect 1182 468 1186 472
rect 1190 468 1194 472
rect 1222 468 1226 472
rect 1238 468 1242 472
rect 1326 468 1330 472
rect 1374 468 1378 472
rect 1390 468 1394 472
rect 1558 468 1562 472
rect 1606 468 1610 472
rect 1806 468 1810 472
rect 2030 468 2034 472
rect 2182 468 2186 472
rect 2198 468 2202 472
rect 2230 468 2234 472
rect 2358 468 2362 472
rect 2390 468 2394 472
rect 2406 468 2410 472
rect 2422 468 2426 472
rect 22 458 26 462
rect 142 458 146 462
rect 182 459 186 463
rect 254 458 258 462
rect 286 458 290 462
rect 294 458 298 462
rect 342 458 346 462
rect 390 458 394 462
rect 422 459 426 463
rect 582 459 586 463
rect 646 458 650 462
rect 718 458 722 462
rect 798 458 802 462
rect 902 458 906 462
rect 982 459 986 463
rect 1070 458 1074 462
rect 1110 458 1114 462
rect 1198 458 1202 462
rect 1278 458 1282 462
rect 1302 458 1306 462
rect 1342 458 1346 462
rect 1422 459 1426 463
rect 1446 458 1450 462
rect 1518 458 1522 462
rect 1542 458 1546 462
rect 1550 458 1554 462
rect 1598 458 1602 462
rect 1638 458 1642 462
rect 1678 458 1682 462
rect 1702 458 1706 462
rect 1742 458 1746 462
rect 1798 458 1802 462
rect 1878 458 1882 462
rect 1886 458 1890 462
rect 1910 458 1914 462
rect 1958 458 1962 462
rect 1990 459 1994 463
rect 2046 458 2050 462
rect 2070 458 2074 462
rect 2078 458 2082 462
rect 2118 458 2122 462
rect 2150 459 2154 463
rect 2222 458 2226 462
rect 2254 458 2258 462
rect 2262 458 2266 462
rect 2270 458 2274 462
rect 2310 458 2314 462
rect 2342 458 2346 462
rect 2350 458 2354 462
rect 2366 458 2370 462
rect 2438 459 2442 463
rect 118 448 122 452
rect 142 448 146 452
rect 318 448 322 452
rect 742 448 746 452
rect 878 448 882 452
rect 1046 448 1050 452
rect 1222 448 1226 452
rect 1390 448 1394 452
rect 1574 448 1578 452
rect 2198 448 2202 452
rect 2390 448 2394 452
rect 6 438 10 442
rect 358 438 362 442
rect 454 438 458 442
rect 510 438 514 442
rect 1238 438 1242 442
rect 38 418 42 422
rect 1654 418 1658 422
rect 1726 418 1730 422
rect 1782 418 1786 422
rect 1862 418 1866 422
rect 482 403 486 407
rect 489 403 493 407
rect 1498 403 1502 407
rect 1505 403 1509 407
rect 126 388 130 392
rect 326 388 330 392
rect 374 388 378 392
rect 462 388 466 392
rect 582 388 586 392
rect 670 388 674 392
rect 710 388 714 392
rect 934 388 938 392
rect 1022 388 1026 392
rect 1222 388 1226 392
rect 1430 388 1434 392
rect 1462 388 1466 392
rect 1614 388 1618 392
rect 1710 388 1714 392
rect 1798 388 1802 392
rect 1990 388 1994 392
rect 294 368 298 372
rect 822 368 826 372
rect 1182 368 1186 372
rect 1198 368 1202 372
rect 1302 368 1306 372
rect 1878 368 1882 372
rect 2510 368 2514 372
rect 30 347 34 351
rect 134 348 138 352
rect 142 348 146 352
rect 158 348 162 352
rect 182 358 186 362
rect 414 358 418 362
rect 230 347 234 351
rect 302 348 306 352
rect 310 348 314 352
rect 334 348 338 352
rect 358 348 362 352
rect 382 348 386 352
rect 390 348 394 352
rect 518 358 522 362
rect 438 348 442 352
rect 478 348 482 352
rect 846 358 850 362
rect 550 348 554 352
rect 558 348 562 352
rect 566 348 570 352
rect 614 348 618 352
rect 638 348 642 352
rect 646 348 650 352
rect 662 348 666 352
rect 686 348 690 352
rect 694 348 698 352
rect 726 348 730 352
rect 766 348 770 352
rect 854 348 858 352
rect 902 348 906 352
rect 918 348 922 352
rect 942 348 946 352
rect 950 348 954 352
rect 982 348 986 352
rect 1014 348 1018 352
rect 1038 348 1042 352
rect 1046 348 1050 352
rect 1062 348 1066 352
rect 1086 358 1090 362
rect 1414 358 1418 362
rect 1670 358 1674 362
rect 1838 358 1842 362
rect 38 338 42 342
rect 150 338 154 342
rect 182 338 186 342
rect 198 338 202 342
rect 214 338 218 342
rect 398 338 402 342
rect 502 338 506 342
rect 550 338 554 342
rect 1134 347 1138 351
rect 1158 348 1162 352
rect 1206 348 1210 352
rect 1214 348 1218 352
rect 1238 348 1242 352
rect 1262 348 1266 352
rect 1286 348 1290 352
rect 1294 348 1298 352
rect 1366 347 1370 351
rect 1454 348 1458 352
rect 1478 348 1482 352
rect 1486 348 1490 352
rect 1574 347 1578 351
rect 1638 348 1642 352
rect 1686 348 1690 352
rect 1694 348 1698 352
rect 1702 348 1706 352
rect 1734 348 1738 352
rect 1742 348 1746 352
rect 1774 348 1778 352
rect 1782 348 1786 352
rect 1862 358 1866 362
rect 2134 358 2138 362
rect 1862 348 1866 352
rect 1918 348 1922 352
rect 1934 348 1938 352
rect 1974 348 1978 352
rect 1982 348 1986 352
rect 2006 348 2010 352
rect 2070 348 2074 352
rect 2086 348 2090 352
rect 2158 348 2162 352
rect 2166 348 2170 352
rect 2198 348 2202 352
rect 2214 348 2218 352
rect 2238 358 2242 362
rect 2294 348 2298 352
rect 2302 348 2306 352
rect 2326 348 2330 352
rect 2358 348 2362 352
rect 2374 348 2378 352
rect 2398 358 2402 362
rect 774 338 778 342
rect 830 338 834 342
rect 862 338 866 342
rect 870 338 874 342
rect 1054 338 1058 342
rect 1078 338 1082 342
rect 1102 338 1106 342
rect 1382 338 1386 342
rect 1398 338 1402 342
rect 1422 338 1426 342
rect 1566 338 1570 342
rect 1670 338 1674 342
rect 1822 338 1826 342
rect 1870 338 1874 342
rect 2150 338 2154 342
rect 2190 338 2194 342
rect 2206 338 2210 342
rect 2262 338 2266 342
rect 2270 338 2274 342
rect 2350 338 2354 342
rect 2446 347 2450 351
rect 2398 338 2402 342
rect 2414 338 2418 342
rect 2430 338 2434 342
rect 78 328 82 332
rect 526 328 530 332
rect 886 328 890 332
rect 966 328 970 332
rect 1366 328 1370 332
rect 1574 328 1578 332
rect 2310 328 2314 332
rect 422 318 426 322
rect 846 318 850 322
rect 1270 318 1274 322
rect 1406 318 1410 322
rect 1510 318 1514 322
rect 1614 318 1618 322
rect 1678 318 1682 322
rect 1758 318 1762 322
rect 2030 318 2034 322
rect 2142 318 2146 322
rect 2230 318 2234 322
rect 2342 318 2346 322
rect 986 303 990 307
rect 993 303 997 307
rect 2018 303 2022 307
rect 2025 303 2029 307
rect 30 288 34 292
rect 206 288 210 292
rect 302 288 306 292
rect 310 288 314 292
rect 542 288 546 292
rect 710 288 714 292
rect 734 288 738 292
rect 854 288 858 292
rect 966 288 970 292
rect 1414 288 1418 292
rect 1422 288 1426 292
rect 1470 288 1474 292
rect 1534 288 1538 292
rect 1582 288 1586 292
rect 1622 288 1626 292
rect 1670 288 1674 292
rect 1718 288 1722 292
rect 1870 288 1874 292
rect 1982 288 1986 292
rect 2046 288 2050 292
rect 2086 288 2090 292
rect 2182 288 2186 292
rect 2286 288 2290 292
rect 2302 288 2306 292
rect 2398 288 2402 292
rect 2518 288 2522 292
rect 374 278 378 282
rect 1142 278 1146 282
rect 2462 278 2466 282
rect 6 268 10 272
rect 54 268 58 272
rect 62 268 66 272
rect 110 268 114 272
rect 166 268 170 272
rect 390 268 394 272
rect 486 268 490 272
rect 566 268 570 272
rect 582 268 586 272
rect 614 268 618 272
rect 662 268 666 272
rect 766 268 770 272
rect 782 268 786 272
rect 814 268 818 272
rect 958 268 962 272
rect 1062 268 1066 272
rect 1078 268 1082 272
rect 1110 268 1114 272
rect 1118 268 1122 272
rect 1166 268 1170 272
rect 1270 268 1274 272
rect 1302 268 1306 272
rect 1318 268 1322 272
rect 1334 268 1338 272
rect 1446 268 1450 272
rect 1646 268 1650 272
rect 1694 268 1698 272
rect 1710 268 1714 272
rect 1766 268 1770 272
rect 1814 268 1818 272
rect 1862 268 1866 272
rect 1950 268 1954 272
rect 2054 268 2058 272
rect 2118 268 2122 272
rect 2150 268 2154 272
rect 2278 268 2282 272
rect 2366 268 2370 272
rect 2494 268 2498 272
rect 46 258 50 262
rect 102 258 106 262
rect 142 259 146 263
rect 174 258 178 262
rect 246 258 250 262
rect 262 258 266 262
rect 374 259 378 263
rect 470 259 474 263
rect 518 258 522 262
rect 526 258 530 262
rect 550 258 554 262
rect 574 258 578 262
rect 654 258 658 262
rect 726 258 730 262
rect 750 258 754 262
rect 758 258 762 262
rect 806 258 810 262
rect 830 258 834 262
rect 838 258 842 262
rect 902 258 906 262
rect 998 258 1002 262
rect 1030 259 1034 263
rect 1102 258 1106 262
rect 1110 258 1114 262
rect 1126 258 1130 262
rect 1198 259 1202 263
rect 1222 258 1226 262
rect 1278 258 1282 262
rect 1350 259 1354 263
rect 1438 258 1442 262
rect 1454 258 1458 262
rect 1462 258 1466 262
rect 1486 258 1490 262
rect 1518 258 1522 262
rect 1526 258 1530 262
rect 1550 258 1554 262
rect 1558 258 1562 262
rect 1590 258 1594 262
rect 1638 258 1642 262
rect 1654 258 1658 262
rect 1678 258 1682 262
rect 1702 258 1706 262
rect 1774 258 1778 262
rect 1854 258 1858 262
rect 1902 258 1906 262
rect 1926 258 1930 262
rect 1966 258 1970 262
rect 1974 258 1978 262
rect 1998 258 2002 262
rect 2030 258 2034 262
rect 2102 258 2106 262
rect 2126 258 2130 262
rect 2150 258 2154 262
rect 2174 258 2178 262
rect 2222 258 2226 262
rect 2238 258 2242 262
rect 2358 258 2362 262
rect 2438 258 2442 262
rect 2454 258 2458 262
rect 2502 258 2506 262
rect 22 248 26 252
rect 78 248 82 252
rect 102 248 106 252
rect 598 248 602 252
rect 782 248 786 252
rect 846 248 850 252
rect 1078 248 1082 252
rect 1150 248 1154 252
rect 1302 248 1306 252
rect 1422 248 1426 252
rect 1614 248 1618 252
rect 1830 248 1834 252
rect 1854 248 1858 252
rect 2078 248 2082 252
rect 2142 248 2146 252
rect 2294 248 2298 252
rect 2518 248 2522 252
rect 1262 238 1266 242
rect 406 228 410 232
rect 1582 218 1586 222
rect 2046 218 2050 222
rect 482 203 486 207
rect 489 203 493 207
rect 1498 203 1502 207
rect 1505 203 1509 207
rect 390 188 394 192
rect 430 188 434 192
rect 470 188 474 192
rect 678 188 682 192
rect 886 188 890 192
rect 958 188 962 192
rect 1262 188 1266 192
rect 1758 188 1762 192
rect 2118 188 2122 192
rect 2366 188 2370 192
rect 2438 188 2442 192
rect 2510 188 2514 192
rect 1590 178 1594 182
rect 6 168 10 172
rect 782 168 786 172
rect 806 168 810 172
rect 1142 168 1146 172
rect 1158 168 1162 172
rect 1286 168 1290 172
rect 1694 168 1698 172
rect 1998 168 2002 172
rect 2254 168 2258 172
rect 118 158 122 162
rect 158 158 162 162
rect 622 158 626 162
rect 70 147 74 151
rect 142 148 146 152
rect 174 148 178 152
rect 214 148 218 152
rect 262 147 266 151
rect 446 148 450 152
rect 478 148 482 152
rect 486 148 490 152
rect 510 148 514 152
rect 822 158 826 162
rect 646 148 650 152
rect 654 148 658 152
rect 694 148 698 152
rect 702 148 706 152
rect 742 148 746 152
rect 1102 158 1106 162
rect 846 148 850 152
rect 998 148 1002 152
rect 1022 148 1026 152
rect 1030 148 1034 152
rect 1038 148 1042 152
rect 1070 148 1074 152
rect 1078 148 1082 152
rect 1398 158 1402 162
rect 1118 148 1122 152
rect 1126 148 1130 152
rect 1198 148 1202 152
rect 1238 148 1242 152
rect 1246 148 1250 152
rect 1278 148 1282 152
rect 1342 148 1346 152
rect 1438 158 1442 162
rect 1462 158 1466 162
rect 1566 158 1570 162
rect 1422 148 1426 152
rect 1510 148 1514 152
rect 1534 148 1538 152
rect 1542 148 1546 152
rect 1702 158 1706 162
rect 1590 148 1594 152
rect 1630 147 1634 151
rect 1734 148 1738 152
rect 1742 148 1746 152
rect 1806 148 1810 152
rect 1862 148 1866 152
rect 1886 158 1890 162
rect 1942 148 1946 152
rect 2054 148 2058 152
rect 2062 148 2066 152
rect 2094 148 2098 152
rect 2102 148 2106 152
rect 2110 148 2114 152
rect 2134 148 2138 152
rect 2158 148 2162 152
rect 2182 158 2186 162
rect 2214 148 2218 152
rect 2238 158 2242 162
rect 2502 158 2506 162
rect 2318 148 2322 152
rect 102 138 106 142
rect 126 138 130 142
rect 150 138 154 142
rect 174 138 178 142
rect 190 138 194 142
rect 206 138 210 142
rect 246 138 250 142
rect 334 138 338 142
rect 438 138 442 142
rect 534 138 538 142
rect 598 138 602 142
rect 606 138 610 142
rect 638 138 642 142
rect 654 138 658 142
rect 718 138 722 142
rect 806 138 810 142
rect 822 138 826 142
rect 862 138 866 142
rect 894 138 898 142
rect 902 138 906 142
rect 1046 138 1050 142
rect 1086 138 1090 142
rect 1134 138 1138 142
rect 1222 138 1226 142
rect 1326 138 1330 142
rect 1366 138 1370 142
rect 1382 138 1386 142
rect 1398 138 1402 142
rect 1430 138 1434 142
rect 1454 138 1458 142
rect 1478 138 1482 142
rect 1494 138 1498 142
rect 1550 138 1554 142
rect 1598 138 1602 142
rect 1614 138 1618 142
rect 1718 138 1722 142
rect 1750 138 1754 142
rect 1838 138 1842 142
rect 1854 138 1858 142
rect 1902 138 1906 142
rect 1918 138 1922 142
rect 2014 138 2018 142
rect 2070 138 2074 142
rect 2150 138 2154 142
rect 2166 138 2170 142
rect 2198 138 2202 142
rect 2206 138 2210 142
rect 2238 138 2242 142
rect 2254 138 2258 142
rect 2342 138 2346 142
rect 2358 138 2362 142
rect 2422 138 2426 142
rect 2430 138 2434 142
rect 2494 138 2498 142
rect 2518 138 2522 142
rect 70 128 74 132
rect 230 128 234 132
rect 1014 128 1018 132
rect 1878 128 1882 132
rect 166 118 170 122
rect 326 118 330 122
rect 430 118 434 122
rect 526 118 530 122
rect 958 118 962 122
rect 1438 118 1442 122
rect 1462 118 1466 122
rect 986 103 990 107
rect 993 103 997 107
rect 2018 103 2022 107
rect 2025 103 2029 107
rect 270 88 274 92
rect 422 88 426 92
rect 494 88 498 92
rect 598 88 602 92
rect 710 88 714 92
rect 894 88 898 92
rect 910 88 914 92
rect 1390 88 1394 92
rect 1478 88 1482 92
rect 1702 88 1706 92
rect 1942 88 1946 92
rect 2110 88 2114 92
rect 2206 88 2210 92
rect 2270 88 2274 92
rect 2446 88 2450 92
rect 2486 88 2490 92
rect 294 78 298 82
rect 6 68 10 72
rect 70 68 74 72
rect 78 68 82 72
rect 150 68 154 72
rect 190 68 194 72
rect 662 78 666 82
rect 782 78 786 82
rect 1206 78 1210 82
rect 1326 78 1330 82
rect 1766 78 1770 82
rect 2518 78 2522 82
rect 318 68 322 72
rect 342 68 346 72
rect 430 68 434 72
rect 462 68 466 72
rect 478 68 482 72
rect 494 68 498 72
rect 534 68 538 72
rect 582 68 586 72
rect 678 68 682 72
rect 734 68 738 72
rect 838 68 842 72
rect 870 68 874 72
rect 958 68 962 72
rect 1006 68 1010 72
rect 1038 68 1042 72
rect 1070 68 1074 72
rect 1078 68 1082 72
rect 1142 68 1146 72
rect 1158 68 1162 72
rect 1198 68 1202 72
rect 1262 68 1266 72
rect 1294 68 1298 72
rect 1398 68 1402 72
rect 1430 68 1434 72
rect 1470 68 1474 72
rect 1558 68 1562 72
rect 1574 68 1578 72
rect 1638 68 1642 72
rect 1646 68 1650 72
rect 150 58 154 62
rect 158 58 162 62
rect 166 58 170 62
rect 206 59 210 63
rect 278 58 282 62
rect 310 58 314 62
rect 326 58 330 62
rect 358 59 362 63
rect 438 58 442 62
rect 558 58 562 62
rect 638 58 642 62
rect 694 58 698 62
rect 758 58 762 62
rect 862 58 866 62
rect 878 58 882 62
rect 974 59 978 63
rect 1062 58 1066 62
rect 1182 58 1186 62
rect 1286 58 1290 62
rect 1334 58 1338 62
rect 1414 58 1418 62
rect 1438 58 1442 62
rect 1678 68 1682 72
rect 1782 68 1786 72
rect 1814 68 1818 72
rect 1846 68 1850 72
rect 1894 68 1898 72
rect 1950 68 1954 72
rect 1982 68 1986 72
rect 2006 68 2010 72
rect 2062 68 2066 72
rect 2158 68 2162 72
rect 2214 68 2218 72
rect 2246 68 2250 72
rect 2350 68 2354 72
rect 2366 68 2370 72
rect 2430 68 2434 72
rect 2478 68 2482 72
rect 1534 58 1538 62
rect 1654 58 1658 62
rect 1670 58 1674 62
rect 1758 58 1762 62
rect 1838 58 1842 62
rect 1878 59 1882 63
rect 1958 58 1962 62
rect 2046 59 2050 63
rect 2166 58 2170 62
rect 2222 58 2226 62
rect 2326 58 2330 62
rect 174 48 178 52
rect 462 48 466 52
rect 838 48 842 52
rect 1038 48 1042 52
rect 1262 48 1266 52
rect 1398 48 1402 52
rect 1462 48 1466 52
rect 1694 48 1698 52
rect 1798 48 1802 52
rect 1838 48 1842 52
rect 1982 48 1986 52
rect 2246 48 2250 52
rect 482 3 486 7
rect 489 3 493 7
rect 1498 3 1502 7
rect 1505 3 1509 7
<< metal2 >>
rect 262 2428 266 2432
rect 462 2428 466 2432
rect 894 2431 898 2432
rect 886 2428 898 2431
rect 918 2428 922 2432
rect 1142 2428 1146 2432
rect 1550 2431 1554 2432
rect 1542 2428 1554 2431
rect 1806 2428 1810 2432
rect 262 2402 265 2428
rect 90 2358 94 2361
rect 70 2352 73 2358
rect 22 2342 25 2348
rect 50 2338 54 2341
rect 62 2332 65 2338
rect 6 2292 9 2328
rect 42 2318 49 2321
rect 46 2262 49 2318
rect 10 2218 14 2221
rect 70 2212 73 2348
rect 94 2342 97 2348
rect 110 2342 113 2368
rect 170 2348 174 2351
rect 246 2342 249 2398
rect 314 2358 318 2361
rect 294 2352 297 2358
rect 290 2348 294 2351
rect 366 2351 369 2358
rect 318 2342 321 2348
rect 282 2338 286 2341
rect 110 2272 113 2338
rect 174 2272 177 2328
rect 86 2242 89 2268
rect 166 2242 169 2268
rect 186 2258 190 2261
rect 198 2252 201 2268
rect 206 2252 209 2258
rect 10 2188 14 2191
rect 110 2172 113 2218
rect 70 2151 73 2158
rect 86 2142 89 2168
rect 134 2162 137 2228
rect 118 2152 121 2158
rect 134 2152 137 2158
rect 106 2148 110 2151
rect 102 2112 105 2138
rect 10 2088 14 2091
rect 86 2072 89 2078
rect 102 2072 105 2108
rect 66 2059 70 2061
rect 66 2058 73 2059
rect 102 1972 105 2068
rect 122 2058 126 2061
rect 110 2052 113 2058
rect 134 2042 137 2048
rect 6 1872 9 1918
rect 10 1868 14 1871
rect 46 1871 49 1948
rect 42 1868 49 1871
rect 62 1872 65 1968
rect 86 1892 89 1948
rect 126 1942 129 1947
rect 142 1942 145 2168
rect 150 2142 153 2188
rect 166 2142 169 2168
rect 150 2072 153 2078
rect 158 2072 161 2108
rect 182 2092 185 2147
rect 190 2062 193 2208
rect 206 2152 209 2248
rect 214 2132 217 2338
rect 222 2332 225 2338
rect 286 2332 289 2338
rect 334 2322 337 2338
rect 222 2272 225 2288
rect 254 2252 257 2259
rect 254 2152 257 2218
rect 242 2118 246 2121
rect 206 2072 209 2118
rect 246 2102 249 2118
rect 222 2062 225 2068
rect 170 2058 174 2061
rect 190 2052 193 2058
rect 190 1992 193 2048
rect 214 1922 217 2058
rect 110 1862 113 1868
rect 118 1862 121 1868
rect 190 1862 193 1918
rect 206 1872 209 1918
rect 226 1868 230 1871
rect 74 1858 78 1861
rect 146 1858 150 1861
rect 46 1852 49 1858
rect 94 1852 97 1858
rect 26 1848 30 1851
rect 10 1778 14 1781
rect 46 1652 49 1848
rect 94 1802 97 1848
rect 134 1842 137 1848
rect 158 1842 161 1858
rect 70 1751 73 1758
rect 86 1742 89 1768
rect 138 1758 142 1761
rect 102 1742 105 1758
rect 114 1748 118 1751
rect 150 1742 153 1778
rect 174 1772 177 1818
rect 178 1758 182 1761
rect 186 1748 190 1751
rect 138 1738 142 1741
rect 126 1732 129 1738
rect 158 1691 161 1738
rect 182 1732 185 1738
rect 158 1688 166 1691
rect 118 1672 121 1688
rect 114 1658 118 1661
rect 14 1542 17 1618
rect 50 1548 54 1551
rect 102 1542 105 1568
rect 114 1558 118 1561
rect 142 1552 145 1558
rect 130 1548 134 1551
rect 150 1542 153 1668
rect 174 1652 177 1718
rect 206 1692 209 1868
rect 238 1862 241 2018
rect 270 1992 273 2318
rect 314 2288 318 2291
rect 334 2262 337 2288
rect 366 2272 369 2328
rect 358 2262 361 2268
rect 286 2242 289 2258
rect 326 2222 329 2258
rect 350 2252 353 2258
rect 374 2242 377 2338
rect 454 2322 457 2338
rect 426 2318 430 2321
rect 422 2272 425 2288
rect 406 2262 409 2268
rect 382 2252 385 2258
rect 410 2248 414 2251
rect 374 2172 377 2238
rect 286 2152 289 2158
rect 278 2092 281 2118
rect 278 2072 281 2078
rect 294 2072 297 2148
rect 302 2142 305 2148
rect 318 2132 321 2158
rect 350 2152 353 2168
rect 358 2162 361 2168
rect 438 2162 441 2268
rect 454 2252 457 2259
rect 462 2241 465 2428
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 493 2403 496 2407
rect 886 2392 889 2428
rect 918 2402 921 2428
rect 1142 2402 1145 2428
rect 1496 2403 1498 2407
rect 1502 2403 1505 2407
rect 1509 2403 1512 2407
rect 1130 2378 1134 2381
rect 742 2372 745 2378
rect 554 2368 558 2371
rect 574 2362 577 2368
rect 562 2358 566 2361
rect 590 2352 593 2358
rect 638 2352 641 2368
rect 514 2348 518 2351
rect 562 2348 566 2351
rect 598 2342 601 2348
rect 702 2342 705 2368
rect 718 2352 721 2358
rect 854 2352 857 2378
rect 1046 2352 1049 2368
rect 1102 2352 1105 2358
rect 1110 2352 1113 2368
rect 1122 2358 1126 2361
rect 746 2348 750 2351
rect 554 2338 558 2341
rect 754 2338 758 2341
rect 534 2332 537 2338
rect 514 2288 518 2291
rect 550 2262 553 2288
rect 570 2268 574 2271
rect 582 2262 585 2338
rect 622 2262 625 2268
rect 630 2262 633 2328
rect 702 2322 705 2338
rect 646 2262 649 2318
rect 758 2312 761 2318
rect 758 2282 761 2288
rect 678 2262 681 2278
rect 454 2238 465 2241
rect 454 2192 457 2238
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 493 2203 496 2207
rect 330 2118 334 2121
rect 270 1942 273 1968
rect 246 1782 249 1858
rect 254 1792 257 1818
rect 262 1812 265 1938
rect 278 1862 281 2058
rect 286 1952 289 1958
rect 294 1872 297 2058
rect 326 2052 329 2059
rect 342 2022 345 2138
rect 358 2072 361 2078
rect 374 2052 377 2058
rect 390 2052 393 2058
rect 314 1958 318 1961
rect 350 1951 353 1958
rect 214 1752 217 1758
rect 230 1742 233 1758
rect 246 1742 249 1768
rect 270 1762 273 1858
rect 262 1742 265 1747
rect 218 1738 222 1741
rect 230 1682 233 1688
rect 194 1668 198 1671
rect 194 1658 198 1661
rect 190 1632 193 1638
rect 166 1552 169 1618
rect 238 1562 241 1708
rect 246 1682 249 1738
rect 254 1662 257 1668
rect 278 1592 281 1858
rect 294 1852 297 1858
rect 302 1792 305 1818
rect 310 1772 313 1948
rect 318 1932 321 1938
rect 334 1872 337 1938
rect 342 1882 345 1888
rect 330 1858 334 1861
rect 318 1852 321 1858
rect 326 1762 329 1768
rect 290 1748 294 1751
rect 366 1742 369 1748
rect 294 1681 297 1688
rect 294 1678 302 1681
rect 302 1672 305 1678
rect 334 1672 337 1718
rect 350 1692 353 1728
rect 374 1712 377 2048
rect 398 1972 401 2148
rect 406 2112 409 2138
rect 414 2122 417 2148
rect 438 2142 441 2158
rect 526 2132 529 2148
rect 406 2072 409 2108
rect 438 2072 441 2128
rect 406 2052 409 2058
rect 410 1968 414 1971
rect 430 1922 433 1938
rect 406 1882 409 1888
rect 394 1868 398 1871
rect 430 1862 433 1918
rect 438 1882 441 2068
rect 494 2062 497 2118
rect 542 2112 545 2258
rect 590 2242 593 2258
rect 598 2252 601 2258
rect 638 2222 641 2258
rect 614 2202 617 2218
rect 662 2202 665 2218
rect 686 2212 689 2268
rect 746 2258 750 2261
rect 622 2152 625 2158
rect 558 2111 561 2147
rect 558 2108 569 2111
rect 566 2092 569 2108
rect 446 2052 449 2058
rect 510 2052 513 2058
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 493 2003 496 2007
rect 446 1952 449 1988
rect 502 1982 505 2018
rect 462 1952 465 1968
rect 454 1942 457 1948
rect 486 1892 489 1948
rect 510 1942 513 1958
rect 526 1952 529 1958
rect 542 1951 545 2088
rect 574 2082 577 2088
rect 550 1962 553 2068
rect 558 2042 561 2068
rect 582 2062 585 2098
rect 590 2062 593 2118
rect 622 2062 625 2068
rect 630 2062 633 2068
rect 610 2058 614 2061
rect 542 1948 550 1951
rect 518 1942 521 1948
rect 558 1942 561 1978
rect 582 1952 585 1958
rect 590 1942 593 2048
rect 606 2012 609 2018
rect 630 1992 633 2038
rect 626 1948 630 1951
rect 638 1951 641 2198
rect 646 2092 649 2158
rect 654 2151 657 2168
rect 670 2142 673 2208
rect 702 2172 705 2178
rect 690 2158 694 2161
rect 766 2152 769 2338
rect 790 2262 793 2268
rect 806 2152 809 2308
rect 822 2302 825 2347
rect 838 2332 841 2338
rect 854 2312 857 2348
rect 870 2292 873 2318
rect 902 2282 905 2348
rect 1102 2342 1105 2348
rect 1158 2342 1161 2398
rect 1542 2392 1545 2428
rect 1806 2402 1809 2428
rect 1198 2342 1201 2348
rect 978 2338 982 2341
rect 854 2272 857 2278
rect 910 2272 913 2338
rect 1006 2332 1009 2338
rect 818 2259 822 2261
rect 818 2258 825 2259
rect 722 2148 726 2151
rect 654 2082 657 2088
rect 646 2022 649 2048
rect 650 1958 654 1961
rect 638 1948 646 1951
rect 606 1942 609 1948
rect 650 1938 654 1941
rect 542 1892 545 1918
rect 474 1888 478 1891
rect 558 1882 561 1938
rect 614 1932 617 1938
rect 422 1822 425 1858
rect 438 1852 441 1858
rect 446 1822 449 1868
rect 454 1862 457 1868
rect 510 1862 513 1878
rect 606 1862 609 1868
rect 398 1751 401 1758
rect 350 1672 353 1688
rect 414 1682 417 1738
rect 430 1721 433 1758
rect 446 1752 449 1798
rect 438 1742 441 1748
rect 422 1718 433 1721
rect 422 1692 425 1718
rect 322 1668 326 1671
rect 358 1662 361 1678
rect 390 1662 393 1668
rect 406 1662 409 1668
rect 342 1652 345 1658
rect 198 1552 201 1558
rect 238 1552 241 1558
rect 186 1548 190 1551
rect 218 1548 222 1551
rect 158 1542 161 1548
rect 206 1542 209 1548
rect 106 1538 110 1541
rect 14 1472 17 1538
rect 150 1472 153 1538
rect 226 1528 230 1531
rect 178 1518 182 1521
rect 122 1468 126 1471
rect 146 1468 150 1471
rect 38 1462 41 1468
rect 54 1442 57 1458
rect 102 1442 105 1468
rect 146 1458 150 1461
rect 118 1452 121 1458
rect 166 1442 169 1468
rect 202 1458 206 1461
rect 34 1388 38 1391
rect 6 1342 9 1348
rect 54 1342 57 1438
rect 102 1402 105 1438
rect 150 1352 153 1378
rect 174 1362 177 1378
rect 198 1352 201 1358
rect 214 1352 217 1428
rect 230 1352 233 1398
rect 82 1348 86 1351
rect 162 1348 166 1351
rect 146 1338 150 1341
rect 134 1322 137 1328
rect 94 1282 97 1288
rect 118 1272 121 1278
rect 14 1192 17 1268
rect 54 1262 57 1268
rect 126 1262 129 1268
rect 142 1262 145 1318
rect 158 1272 161 1338
rect 190 1332 193 1338
rect 214 1332 217 1338
rect 190 1292 193 1328
rect 178 1268 182 1271
rect 142 1252 145 1258
rect 106 1248 110 1251
rect 150 1241 153 1268
rect 170 1258 174 1261
rect 182 1252 185 1258
rect 198 1252 201 1318
rect 238 1272 241 1548
rect 262 1542 265 1568
rect 258 1538 262 1541
rect 302 1532 305 1548
rect 254 1431 257 1468
rect 274 1458 278 1461
rect 262 1442 265 1458
rect 286 1442 289 1448
rect 254 1428 265 1431
rect 250 1418 254 1421
rect 246 1362 249 1368
rect 254 1332 257 1348
rect 262 1342 265 1428
rect 302 1422 305 1468
rect 310 1452 313 1478
rect 270 1362 273 1388
rect 270 1352 273 1358
rect 290 1338 294 1341
rect 278 1292 281 1328
rect 302 1282 305 1338
rect 318 1322 321 1648
rect 378 1638 382 1641
rect 366 1592 369 1628
rect 390 1592 393 1618
rect 398 1612 401 1658
rect 426 1648 430 1651
rect 438 1642 441 1658
rect 446 1652 449 1748
rect 454 1742 457 1858
rect 534 1852 537 1858
rect 574 1852 577 1858
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 493 1803 496 1807
rect 534 1792 537 1838
rect 486 1752 489 1778
rect 474 1748 478 1751
rect 454 1692 457 1738
rect 510 1692 513 1758
rect 518 1752 521 1788
rect 526 1762 529 1768
rect 546 1748 550 1751
rect 526 1742 529 1748
rect 574 1742 577 1828
rect 582 1781 585 1858
rect 622 1842 625 1938
rect 630 1862 633 1878
rect 654 1862 657 1878
rect 662 1862 665 2108
rect 670 2062 673 2138
rect 690 2058 694 2061
rect 670 1872 673 2048
rect 702 2022 705 2148
rect 714 2138 718 2141
rect 726 2112 729 2138
rect 750 2132 753 2148
rect 766 2142 769 2148
rect 838 2142 841 2268
rect 866 2258 870 2261
rect 878 2252 881 2258
rect 858 2248 862 2251
rect 870 2232 873 2248
rect 870 2202 873 2228
rect 846 2152 849 2158
rect 778 2138 782 2141
rect 742 2122 745 2128
rect 734 2062 737 2118
rect 758 2092 761 2118
rect 750 2072 753 2078
rect 766 2062 769 2108
rect 774 2072 777 2078
rect 718 2052 721 2059
rect 766 2002 769 2058
rect 790 2052 793 2108
rect 886 2082 889 2088
rect 678 1962 681 1968
rect 690 1958 694 1961
rect 698 1948 702 1951
rect 686 1942 689 1948
rect 678 1922 681 1938
rect 678 1862 681 1868
rect 710 1862 713 1958
rect 742 1952 745 1988
rect 782 1962 785 2018
rect 790 1951 793 2048
rect 822 2042 825 2059
rect 798 1992 801 2038
rect 830 1972 833 2068
rect 894 2062 897 2218
rect 902 2152 905 2268
rect 918 2262 921 2318
rect 1086 2312 1089 2318
rect 984 2303 986 2307
rect 990 2303 993 2307
rect 997 2303 1000 2307
rect 1094 2292 1097 2338
rect 1174 2332 1177 2338
rect 974 2282 977 2288
rect 942 2262 945 2278
rect 1006 2272 1009 2278
rect 1102 2272 1105 2278
rect 1074 2268 1078 2271
rect 1030 2262 1033 2268
rect 954 2258 958 2261
rect 910 2202 913 2258
rect 918 2162 921 2168
rect 922 2148 926 2151
rect 910 2142 913 2148
rect 906 2118 910 2121
rect 902 2062 905 2078
rect 894 2042 897 2058
rect 918 1952 921 2018
rect 790 1948 798 1951
rect 802 1948 806 1951
rect 774 1942 777 1948
rect 934 1951 937 2218
rect 958 2152 961 2158
rect 966 2152 969 2188
rect 998 2152 1001 2178
rect 1014 2152 1017 2258
rect 1038 2212 1041 2268
rect 942 2122 945 2138
rect 986 2118 990 2121
rect 942 2062 945 2118
rect 984 2103 986 2107
rect 990 2103 993 2107
rect 997 2103 1000 2107
rect 974 2062 977 2078
rect 1006 2072 1009 2078
rect 1014 2062 1017 2148
rect 1022 2092 1025 2158
rect 1054 2152 1057 2268
rect 1090 2258 1094 2261
rect 1078 2252 1081 2258
rect 1114 2248 1118 2251
rect 1126 2242 1129 2248
rect 1070 2192 1073 2238
rect 1062 2152 1065 2178
rect 1030 2102 1033 2118
rect 1030 2082 1033 2088
rect 1046 2062 1049 2148
rect 1054 2142 1057 2148
rect 1062 2142 1065 2148
rect 1078 2132 1081 2158
rect 1086 2142 1089 2168
rect 1078 2062 1081 2098
rect 1118 2091 1121 2138
rect 1134 2112 1137 2318
rect 1190 2292 1193 2318
rect 1214 2292 1217 2358
rect 1262 2342 1265 2368
rect 1282 2358 1286 2361
rect 1346 2358 1350 2361
rect 1278 2352 1281 2358
rect 1302 2352 1305 2358
rect 1326 2352 1329 2358
rect 1598 2352 1601 2358
rect 1514 2348 1518 2351
rect 1570 2348 1574 2351
rect 1282 2338 1286 2341
rect 1150 2272 1153 2288
rect 1142 2152 1145 2218
rect 1150 2132 1153 2258
rect 1158 2222 1161 2278
rect 1198 2262 1201 2268
rect 1206 2262 1209 2288
rect 1230 2272 1233 2308
rect 1178 2258 1182 2261
rect 1166 2212 1169 2238
rect 1166 2142 1169 2208
rect 1206 2192 1209 2228
rect 1214 2222 1217 2248
rect 1182 2132 1185 2138
rect 1110 2088 1121 2091
rect 1110 2072 1113 2088
rect 950 2032 953 2058
rect 982 2052 985 2058
rect 1022 2052 1025 2058
rect 958 1962 961 2018
rect 1010 1958 1014 1961
rect 966 1952 969 1958
rect 934 1948 942 1951
rect 954 1948 958 1951
rect 802 1938 806 1941
rect 718 1921 721 1938
rect 726 1932 729 1938
rect 718 1918 729 1921
rect 726 1892 729 1918
rect 806 1902 809 1938
rect 718 1872 721 1888
rect 814 1882 817 1918
rect 878 1892 881 1947
rect 894 1932 897 1938
rect 930 1918 934 1921
rect 958 1902 961 1938
rect 966 1932 969 1948
rect 990 1942 993 1958
rect 1002 1948 1006 1951
rect 984 1903 986 1907
rect 990 1903 993 1907
rect 997 1903 1000 1907
rect 846 1872 849 1888
rect 902 1872 905 1898
rect 930 1888 934 1891
rect 958 1882 961 1898
rect 910 1872 913 1878
rect 958 1872 961 1878
rect 738 1868 742 1871
rect 858 1868 862 1871
rect 638 1852 641 1858
rect 662 1842 665 1858
rect 670 1852 673 1858
rect 718 1852 721 1858
rect 690 1828 694 1831
rect 590 1792 593 1818
rect 582 1778 590 1781
rect 642 1778 646 1781
rect 542 1732 545 1738
rect 550 1721 553 1738
rect 566 1732 569 1738
rect 542 1718 553 1721
rect 454 1672 457 1678
rect 498 1668 502 1671
rect 462 1642 465 1658
rect 470 1652 473 1658
rect 446 1592 449 1638
rect 478 1622 481 1658
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 493 1603 496 1607
rect 454 1552 457 1568
rect 370 1548 374 1551
rect 474 1548 478 1551
rect 490 1548 494 1551
rect 342 1532 345 1538
rect 330 1488 334 1491
rect 326 1472 329 1478
rect 342 1472 345 1528
rect 350 1492 353 1508
rect 358 1492 361 1548
rect 422 1542 425 1548
rect 462 1542 465 1548
rect 326 1452 329 1458
rect 342 1452 345 1458
rect 358 1392 361 1468
rect 366 1412 369 1518
rect 374 1502 377 1528
rect 374 1492 377 1498
rect 378 1478 382 1481
rect 382 1472 385 1478
rect 374 1462 377 1468
rect 374 1352 377 1418
rect 390 1322 393 1518
rect 406 1482 409 1518
rect 414 1492 417 1538
rect 422 1462 425 1518
rect 470 1512 473 1548
rect 510 1542 513 1638
rect 518 1632 521 1668
rect 526 1662 529 1698
rect 542 1622 545 1718
rect 558 1682 561 1688
rect 566 1652 569 1658
rect 582 1642 585 1748
rect 590 1742 593 1778
rect 630 1762 633 1768
rect 606 1722 609 1758
rect 702 1752 705 1758
rect 630 1722 633 1748
rect 638 1742 641 1748
rect 626 1688 630 1691
rect 638 1682 641 1738
rect 638 1671 641 1678
rect 634 1668 641 1671
rect 678 1672 681 1688
rect 686 1662 689 1718
rect 702 1692 705 1698
rect 710 1662 713 1728
rect 726 1662 729 1758
rect 734 1662 737 1688
rect 742 1672 745 1748
rect 750 1742 753 1858
rect 790 1851 793 1868
rect 878 1862 881 1868
rect 966 1862 969 1868
rect 998 1862 1001 1868
rect 802 1858 806 1861
rect 894 1852 897 1858
rect 790 1848 801 1851
rect 874 1848 878 1851
rect 798 1832 801 1848
rect 774 1732 777 1748
rect 782 1742 785 1748
rect 798 1742 801 1828
rect 642 1658 646 1661
rect 698 1658 702 1661
rect 662 1652 665 1658
rect 638 1642 641 1648
rect 518 1592 521 1618
rect 662 1612 665 1648
rect 686 1582 689 1658
rect 530 1568 534 1571
rect 598 1551 601 1568
rect 650 1558 654 1561
rect 662 1552 665 1568
rect 670 1552 673 1558
rect 546 1538 550 1541
rect 486 1482 489 1528
rect 502 1482 505 1488
rect 434 1468 438 1471
rect 450 1468 454 1471
rect 434 1458 438 1461
rect 398 1392 401 1458
rect 450 1448 454 1451
rect 462 1451 465 1468
rect 474 1458 478 1461
rect 458 1448 465 1451
rect 474 1448 478 1451
rect 414 1361 417 1418
rect 510 1412 513 1538
rect 566 1532 569 1548
rect 630 1542 633 1548
rect 526 1492 529 1528
rect 558 1492 561 1508
rect 670 1492 673 1548
rect 678 1542 681 1558
rect 686 1532 689 1538
rect 550 1482 553 1488
rect 542 1472 545 1478
rect 566 1472 569 1478
rect 582 1472 585 1478
rect 686 1472 689 1528
rect 518 1462 521 1468
rect 566 1462 569 1468
rect 678 1452 681 1458
rect 414 1358 425 1361
rect 422 1352 425 1358
rect 430 1352 433 1408
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 493 1403 496 1407
rect 518 1402 521 1418
rect 450 1388 454 1391
rect 486 1352 489 1368
rect 474 1348 478 1351
rect 406 1342 409 1348
rect 142 1238 153 1241
rect 94 1162 97 1168
rect 78 1142 81 1158
rect 70 1132 73 1138
rect 14 1092 17 1118
rect 14 1072 17 1088
rect 102 1072 105 1238
rect 126 1172 129 1218
rect 126 1152 129 1168
rect 114 1148 118 1151
rect 142 1142 145 1238
rect 214 1192 217 1268
rect 222 1262 225 1268
rect 286 1262 289 1278
rect 254 1192 257 1208
rect 162 1148 166 1151
rect 122 1138 126 1141
rect 110 1092 113 1138
rect 174 1132 177 1138
rect 182 1092 185 1188
rect 226 1168 230 1171
rect 134 1072 137 1088
rect 182 1072 185 1088
rect 126 1062 129 1068
rect 30 1021 33 1059
rect 194 1059 198 1062
rect 22 1018 33 1021
rect 22 992 25 1018
rect 6 932 9 958
rect 22 952 25 978
rect 74 948 78 951
rect 10 868 14 871
rect 22 852 25 948
rect 30 942 33 948
rect 62 892 65 928
rect 78 892 81 928
rect 62 882 65 888
rect 94 872 97 1018
rect 110 942 113 1018
rect 126 942 129 968
rect 134 952 137 1018
rect 202 958 206 961
rect 166 942 169 948
rect 154 928 158 931
rect 110 872 113 878
rect 82 848 86 851
rect 142 772 145 858
rect 102 752 105 768
rect 118 752 121 758
rect 30 692 33 747
rect 54 681 57 738
rect 50 678 57 681
rect 62 681 65 748
rect 126 742 129 748
rect 134 742 137 748
rect 62 678 73 681
rect 54 672 57 678
rect 10 668 14 671
rect 62 662 65 668
rect 50 658 54 661
rect 22 652 25 658
rect 6 542 9 578
rect 22 562 25 568
rect 46 552 49 558
rect 38 542 41 548
rect 70 542 73 678
rect 94 672 97 718
rect 102 662 105 688
rect 78 652 81 658
rect 94 582 97 658
rect 86 551 89 558
rect 50 538 54 541
rect 70 532 73 538
rect 38 492 41 528
rect 118 502 121 668
rect 142 662 145 718
rect 150 672 153 858
rect 174 832 177 948
rect 182 942 185 948
rect 198 942 201 948
rect 202 888 206 891
rect 194 838 198 841
rect 190 752 193 758
rect 198 752 201 768
rect 214 762 217 1168
rect 222 1162 225 1168
rect 238 1152 241 1168
rect 294 1162 297 1268
rect 326 1262 329 1298
rect 374 1272 377 1308
rect 390 1262 393 1288
rect 362 1258 366 1261
rect 302 1252 305 1258
rect 318 1242 321 1258
rect 334 1252 337 1258
rect 342 1212 345 1258
rect 382 1252 385 1258
rect 282 1158 286 1161
rect 322 1158 326 1161
rect 294 1152 297 1158
rect 378 1148 382 1151
rect 230 1092 233 1148
rect 278 1091 281 1138
rect 278 1088 286 1091
rect 274 1068 278 1071
rect 230 1062 233 1068
rect 246 1062 249 1068
rect 246 1042 249 1048
rect 270 1042 273 1058
rect 222 962 225 1028
rect 278 972 281 1068
rect 222 952 225 958
rect 230 942 233 968
rect 294 962 297 1148
rect 302 1142 305 1148
rect 302 1072 305 1138
rect 342 1132 345 1138
rect 326 1062 329 1118
rect 342 1072 345 1128
rect 390 1092 393 1138
rect 258 958 262 961
rect 278 952 281 958
rect 302 952 305 968
rect 318 952 321 958
rect 242 938 246 941
rect 238 892 241 938
rect 230 862 233 878
rect 262 863 265 918
rect 262 858 265 859
rect 214 752 217 758
rect 162 748 166 751
rect 230 742 233 838
rect 278 822 281 948
rect 314 938 318 941
rect 294 872 297 938
rect 302 862 305 938
rect 334 911 337 958
rect 350 942 353 947
rect 334 908 345 911
rect 342 892 345 908
rect 350 882 353 928
rect 326 842 329 858
rect 334 852 337 858
rect 342 852 345 858
rect 302 752 305 758
rect 242 748 246 751
rect 238 742 241 748
rect 270 742 273 748
rect 294 742 297 748
rect 186 738 190 741
rect 250 738 254 741
rect 174 702 177 728
rect 198 692 201 698
rect 214 672 217 678
rect 254 662 257 718
rect 146 578 150 581
rect 254 552 257 568
rect 190 542 193 548
rect 254 542 257 548
rect 94 472 97 498
rect 102 472 105 488
rect 150 472 153 478
rect 166 472 169 538
rect 242 488 246 491
rect 146 458 150 461
rect 6 442 9 448
rect 22 442 25 458
rect 118 452 121 458
rect 146 448 150 451
rect 10 268 14 271
rect 22 252 25 298
rect 30 292 33 347
rect 38 342 41 418
rect 126 392 129 428
rect 38 332 41 338
rect 46 262 49 298
rect 54 272 57 368
rect 62 272 65 288
rect 78 272 81 328
rect 102 262 105 358
rect 130 348 134 351
rect 142 342 145 348
rect 150 342 153 368
rect 158 352 161 388
rect 110 272 113 278
rect 78 252 81 258
rect 142 252 145 259
rect 106 248 110 251
rect 6 152 9 168
rect 150 162 153 338
rect 166 272 169 468
rect 182 452 185 459
rect 182 362 185 388
rect 254 352 257 458
rect 198 342 201 348
rect 230 342 233 347
rect 178 338 182 341
rect 214 332 217 338
rect 206 292 209 308
rect 202 288 206 291
rect 246 262 249 328
rect 262 262 265 658
rect 286 641 289 728
rect 294 692 297 738
rect 318 682 321 818
rect 350 771 353 878
rect 358 862 361 868
rect 366 862 369 1088
rect 414 1022 417 1348
rect 430 1342 433 1348
rect 430 1272 433 1328
rect 446 1312 449 1338
rect 454 1322 457 1348
rect 510 1332 513 1348
rect 518 1342 521 1348
rect 526 1322 529 1338
rect 526 1312 529 1318
rect 534 1302 537 1418
rect 630 1382 633 1418
rect 626 1348 630 1351
rect 438 1282 441 1288
rect 454 1282 457 1288
rect 422 1262 425 1268
rect 446 1262 449 1278
rect 430 1242 433 1258
rect 462 1252 465 1258
rect 470 1242 473 1268
rect 486 1262 489 1288
rect 494 1262 497 1268
rect 494 1232 497 1258
rect 434 1158 438 1161
rect 434 1148 438 1151
rect 446 1132 449 1148
rect 422 1072 425 1118
rect 454 1092 457 1158
rect 462 1142 465 1228
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 482 1168 486 1171
rect 534 1152 537 1158
rect 542 1142 545 1328
rect 582 1292 585 1348
rect 646 1342 649 1368
rect 662 1352 665 1408
rect 678 1362 681 1388
rect 634 1338 638 1341
rect 606 1332 609 1338
rect 654 1331 657 1338
rect 650 1328 657 1331
rect 598 1272 601 1308
rect 622 1282 625 1288
rect 650 1268 654 1271
rect 582 1262 585 1268
rect 558 1252 561 1258
rect 638 1252 641 1258
rect 654 1252 657 1258
rect 618 1248 622 1251
rect 638 1202 641 1248
rect 662 1202 665 1348
rect 686 1272 689 1468
rect 694 1392 697 1468
rect 694 1282 697 1348
rect 674 1268 678 1271
rect 686 1262 689 1268
rect 586 1158 590 1161
rect 606 1152 609 1158
rect 586 1148 590 1151
rect 574 1142 577 1148
rect 446 1072 449 1078
rect 382 932 385 938
rect 410 918 414 921
rect 382 862 385 918
rect 422 892 425 958
rect 438 952 441 1058
rect 462 1051 465 1128
rect 482 1068 486 1071
rect 494 1062 497 1108
rect 542 1092 545 1138
rect 606 1092 609 1148
rect 622 1142 625 1168
rect 646 1162 649 1168
rect 686 1152 689 1158
rect 662 1122 665 1148
rect 670 1112 673 1148
rect 678 1142 681 1148
rect 590 1072 593 1088
rect 694 1072 697 1268
rect 702 1192 705 1368
rect 718 1361 721 1598
rect 742 1592 745 1658
rect 758 1562 761 1678
rect 782 1672 785 1678
rect 798 1662 801 1738
rect 814 1672 817 1747
rect 886 1732 889 1738
rect 874 1718 878 1721
rect 838 1672 841 1718
rect 846 1672 849 1708
rect 858 1668 862 1671
rect 870 1662 873 1698
rect 878 1682 881 1688
rect 766 1592 769 1658
rect 758 1542 761 1558
rect 774 1552 777 1658
rect 790 1652 793 1658
rect 838 1652 841 1658
rect 782 1552 785 1558
rect 790 1552 793 1588
rect 814 1582 817 1648
rect 894 1642 897 1848
rect 926 1822 929 1848
rect 950 1822 953 1858
rect 918 1752 921 1778
rect 982 1762 985 1818
rect 1014 1762 1017 1858
rect 962 1748 966 1751
rect 926 1672 929 1748
rect 942 1732 945 1748
rect 974 1742 977 1748
rect 974 1722 977 1738
rect 982 1732 985 1738
rect 950 1702 953 1718
rect 984 1703 986 1707
rect 990 1703 993 1707
rect 997 1703 1000 1707
rect 958 1672 961 1688
rect 1006 1682 1009 1748
rect 1022 1702 1025 2048
rect 1046 2042 1049 2058
rect 1030 1992 1033 2028
rect 1110 1952 1113 2068
rect 1158 2062 1161 2078
rect 1174 2062 1177 2108
rect 1126 2052 1129 2058
rect 1134 2041 1137 2058
rect 1126 2038 1137 2041
rect 1126 2012 1129 2038
rect 1134 1952 1137 2028
rect 1150 2012 1153 2018
rect 1082 1948 1086 1951
rect 1110 1942 1113 1948
rect 1062 1932 1065 1938
rect 1150 1932 1153 1938
rect 1158 1922 1161 1948
rect 1166 1872 1169 1948
rect 1174 1932 1177 2058
rect 1182 1972 1185 2128
rect 1190 2092 1193 2138
rect 1198 2062 1201 2118
rect 1222 2092 1225 2148
rect 1230 2082 1233 2088
rect 1238 2082 1241 2268
rect 1246 2182 1249 2328
rect 1262 2312 1265 2338
rect 1302 2322 1305 2348
rect 1318 2292 1321 2338
rect 1286 2282 1289 2288
rect 1270 2262 1273 2278
rect 1278 2232 1281 2258
rect 1326 2252 1329 2348
rect 1342 2302 1345 2318
rect 1366 2302 1369 2338
rect 1382 2272 1385 2288
rect 1350 2252 1353 2259
rect 1366 2242 1369 2268
rect 1386 2258 1390 2261
rect 1406 2252 1409 2338
rect 1422 2282 1425 2348
rect 1470 2342 1473 2348
rect 1478 2342 1481 2348
rect 1414 2272 1417 2278
rect 1446 2262 1449 2308
rect 1462 2262 1465 2318
rect 1470 2262 1473 2298
rect 1478 2272 1481 2338
rect 1486 2312 1489 2318
rect 1502 2292 1505 2298
rect 1534 2292 1537 2328
rect 1550 2262 1553 2268
rect 1430 2252 1433 2258
rect 1394 2248 1398 2251
rect 1246 2152 1249 2178
rect 1334 2152 1337 2158
rect 1258 2148 1262 2151
rect 1306 2148 1310 2151
rect 1366 2142 1369 2178
rect 1382 2142 1385 2147
rect 1454 2142 1457 2218
rect 1486 2182 1489 2258
rect 1558 2232 1561 2348
rect 1614 2342 1617 2368
rect 1918 2362 1921 2368
rect 1846 2352 1849 2358
rect 1934 2352 1937 2358
rect 1990 2352 1993 2358
rect 1678 2342 1681 2348
rect 1702 2342 1705 2348
rect 1914 2348 1918 2351
rect 1594 2338 1598 2341
rect 1566 2222 1569 2338
rect 1614 2302 1617 2338
rect 1782 2332 1785 2347
rect 1986 2338 1990 2341
rect 1718 2282 1721 2318
rect 1618 2278 1622 2281
rect 1582 2252 1585 2268
rect 1598 2222 1601 2258
rect 1606 2242 1609 2268
rect 1646 2262 1649 2278
rect 1750 2263 1753 2308
rect 1818 2288 1822 2291
rect 1750 2258 1753 2259
rect 1630 2242 1633 2258
rect 1758 2252 1761 2268
rect 1830 2262 1833 2268
rect 1822 2252 1825 2258
rect 1496 2203 1498 2207
rect 1502 2203 1505 2207
rect 1509 2203 1512 2207
rect 1598 2162 1601 2188
rect 1594 2158 1598 2161
rect 1574 2152 1577 2158
rect 1630 2152 1633 2168
rect 1654 2162 1657 2168
rect 1662 2152 1665 2218
rect 1506 2148 1510 2151
rect 1306 2138 1310 2141
rect 1330 2138 1334 2141
rect 1214 2052 1217 2068
rect 1238 2062 1241 2068
rect 1246 2062 1249 2118
rect 1310 2112 1313 2138
rect 1350 2122 1353 2138
rect 1442 2118 1446 2121
rect 1458 2118 1462 2121
rect 1286 2062 1289 2088
rect 1350 2063 1353 2098
rect 1414 2092 1417 2098
rect 1366 2072 1369 2078
rect 1274 2058 1278 2061
rect 1382 2062 1385 2078
rect 1422 2062 1425 2068
rect 1430 2062 1433 2108
rect 1470 2092 1473 2148
rect 1534 2142 1537 2148
rect 1686 2142 1689 2148
rect 1702 2142 1705 2147
rect 1650 2138 1654 2141
rect 1450 2088 1465 2091
rect 1462 2082 1465 2088
rect 1450 2078 1454 2081
rect 1262 1982 1265 2018
rect 1270 1982 1273 1998
rect 1206 1952 1209 1958
rect 1326 1952 1329 1998
rect 1178 1918 1182 1921
rect 1238 1902 1241 1947
rect 1278 1942 1281 1948
rect 1302 1942 1305 1948
rect 1254 1882 1257 1928
rect 1174 1872 1177 1878
rect 1106 1868 1110 1871
rect 1038 1832 1041 1868
rect 1142 1862 1145 1868
rect 1066 1858 1070 1861
rect 1202 1858 1206 1861
rect 1182 1852 1185 1858
rect 1146 1848 1150 1851
rect 1190 1851 1193 1858
rect 1190 1848 1201 1851
rect 1050 1768 1054 1771
rect 1030 1752 1033 1768
rect 1038 1742 1041 1748
rect 1106 1747 1110 1750
rect 1126 1742 1129 1788
rect 1142 1742 1145 1768
rect 1182 1762 1185 1848
rect 1198 1772 1201 1848
rect 1206 1792 1209 1848
rect 1214 1782 1217 1818
rect 1198 1762 1201 1768
rect 1162 1758 1166 1761
rect 1182 1752 1185 1758
rect 1158 1742 1161 1748
rect 974 1672 977 1678
rect 1038 1672 1041 1708
rect 1086 1692 1089 1738
rect 1086 1672 1089 1688
rect 1134 1682 1137 1688
rect 1142 1672 1145 1708
rect 938 1659 942 1661
rect 1014 1662 1017 1668
rect 938 1658 945 1659
rect 1082 1658 1086 1661
rect 1162 1658 1166 1661
rect 846 1632 849 1638
rect 766 1522 769 1548
rect 774 1511 777 1548
rect 790 1542 793 1548
rect 766 1508 777 1511
rect 738 1478 742 1481
rect 754 1468 758 1471
rect 754 1458 758 1461
rect 766 1422 769 1508
rect 790 1502 793 1528
rect 806 1522 809 1558
rect 814 1552 817 1568
rect 870 1552 873 1558
rect 846 1542 849 1548
rect 774 1452 777 1488
rect 790 1472 793 1498
rect 798 1482 801 1488
rect 734 1402 737 1418
rect 714 1358 721 1361
rect 734 1362 737 1368
rect 710 1292 713 1348
rect 710 1252 713 1288
rect 710 1152 713 1228
rect 554 1068 558 1071
rect 650 1068 654 1071
rect 502 1062 505 1068
rect 458 1048 465 1051
rect 606 1052 609 1059
rect 638 1052 641 1058
rect 662 1052 665 1068
rect 682 1058 686 1061
rect 454 972 457 1048
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 474 988 478 991
rect 510 952 513 1018
rect 550 952 553 968
rect 430 922 433 938
rect 414 872 417 888
rect 406 862 409 868
rect 378 858 382 861
rect 366 792 369 858
rect 438 852 441 948
rect 446 872 449 938
rect 454 912 457 948
rect 462 932 465 948
rect 526 942 529 948
rect 454 882 457 888
rect 494 862 497 918
rect 558 882 561 1038
rect 606 962 609 968
rect 614 952 617 1018
rect 678 972 681 1028
rect 678 962 681 968
rect 622 952 625 958
rect 610 948 614 951
rect 550 872 553 878
rect 350 768 361 771
rect 434 768 438 771
rect 330 758 334 761
rect 326 742 329 748
rect 342 742 345 768
rect 358 742 361 768
rect 446 752 449 838
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 534 802 537 868
rect 454 752 457 768
rect 494 752 497 768
rect 538 748 542 751
rect 550 751 553 868
rect 558 862 561 878
rect 574 852 577 868
rect 582 852 585 878
rect 606 872 609 888
rect 638 862 641 918
rect 646 892 649 948
rect 654 942 657 958
rect 686 942 689 958
rect 694 952 697 1068
rect 702 1052 705 1058
rect 702 952 705 968
rect 710 952 713 1138
rect 718 1102 721 1358
rect 750 1352 753 1418
rect 758 1352 761 1398
rect 782 1352 785 1398
rect 750 1331 753 1348
rect 758 1342 761 1348
rect 790 1342 793 1348
rect 806 1342 809 1518
rect 862 1462 865 1468
rect 850 1458 854 1461
rect 838 1392 841 1448
rect 854 1362 857 1388
rect 878 1362 881 1608
rect 926 1592 929 1658
rect 990 1642 993 1648
rect 1030 1642 1033 1658
rect 1002 1548 1006 1551
rect 894 1482 897 1538
rect 910 1492 913 1548
rect 894 1472 897 1478
rect 882 1358 886 1361
rect 814 1352 817 1358
rect 842 1348 846 1351
rect 854 1342 857 1358
rect 862 1352 865 1358
rect 886 1342 889 1348
rect 846 1332 849 1338
rect 750 1328 761 1331
rect 742 1292 745 1328
rect 742 1182 745 1218
rect 746 1158 750 1161
rect 742 1142 745 1158
rect 726 1122 729 1138
rect 726 1062 729 1068
rect 730 1048 734 1051
rect 742 962 745 1118
rect 750 1092 753 1148
rect 758 1022 761 1328
rect 766 1262 769 1318
rect 782 1272 785 1278
rect 798 1262 801 1308
rect 886 1292 889 1328
rect 894 1292 897 1468
rect 934 1422 937 1548
rect 966 1542 969 1548
rect 1018 1538 1022 1541
rect 934 1392 937 1418
rect 942 1412 945 1538
rect 998 1522 1001 1528
rect 950 1472 953 1518
rect 984 1503 986 1507
rect 990 1503 993 1507
rect 997 1503 1000 1507
rect 990 1462 993 1468
rect 1006 1463 1009 1468
rect 1022 1462 1025 1518
rect 934 1351 937 1358
rect 902 1322 905 1338
rect 846 1272 849 1278
rect 862 1272 865 1278
rect 826 1268 830 1271
rect 786 1258 790 1261
rect 774 1192 777 1258
rect 806 1202 809 1258
rect 814 1252 817 1268
rect 870 1262 873 1288
rect 834 1258 838 1261
rect 834 1248 846 1251
rect 894 1232 897 1268
rect 790 1152 793 1188
rect 782 1142 785 1148
rect 798 1142 801 1168
rect 794 1058 798 1061
rect 738 948 742 951
rect 718 942 721 948
rect 778 948 782 951
rect 650 888 654 891
rect 710 872 713 938
rect 758 932 761 938
rect 806 922 809 1148
rect 814 1082 817 1178
rect 886 1172 889 1218
rect 902 1202 905 1258
rect 830 1152 833 1158
rect 822 1102 825 1118
rect 846 1092 849 1138
rect 886 1132 889 1148
rect 830 892 833 1088
rect 870 1063 873 1098
rect 838 992 841 998
rect 846 892 849 918
rect 814 872 817 888
rect 858 868 862 871
rect 610 858 614 861
rect 650 858 654 861
rect 702 852 705 858
rect 582 772 585 798
rect 630 782 633 818
rect 562 768 566 771
rect 670 752 673 838
rect 550 748 558 751
rect 618 748 622 751
rect 374 742 377 747
rect 446 742 449 748
rect 330 668 334 671
rect 342 662 345 698
rect 350 662 353 668
rect 358 662 361 678
rect 398 672 401 678
rect 446 662 449 718
rect 454 662 457 668
rect 462 662 465 668
rect 478 662 481 738
rect 494 732 497 748
rect 526 742 529 748
rect 646 742 649 748
rect 546 738 550 741
rect 518 672 521 678
rect 510 662 513 668
rect 298 658 302 661
rect 378 658 382 661
rect 402 658 406 661
rect 310 652 313 658
rect 414 652 417 658
rect 294 642 297 648
rect 286 638 294 641
rect 270 562 273 588
rect 270 392 273 558
rect 294 552 297 588
rect 282 538 286 541
rect 278 492 281 528
rect 286 462 289 498
rect 302 482 305 538
rect 310 502 313 518
rect 310 471 313 498
rect 326 492 329 538
rect 306 468 313 471
rect 294 462 297 468
rect 342 462 345 628
rect 430 592 433 658
rect 446 651 449 658
rect 446 648 457 651
rect 454 562 457 648
rect 470 592 473 658
rect 502 612 505 658
rect 518 642 521 648
rect 526 622 529 738
rect 534 672 537 708
rect 558 672 561 678
rect 578 668 582 671
rect 630 671 633 738
rect 686 722 689 748
rect 670 692 673 718
rect 666 678 689 681
rect 686 672 689 678
rect 702 672 705 838
rect 710 792 713 868
rect 734 862 737 868
rect 750 862 753 868
rect 742 752 745 768
rect 758 752 761 758
rect 730 748 734 751
rect 630 668 641 671
rect 650 668 654 671
rect 674 668 678 671
rect 550 662 553 668
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 518 582 521 598
rect 542 592 545 658
rect 582 652 585 658
rect 574 642 577 648
rect 590 642 593 668
rect 638 662 641 668
rect 710 662 713 698
rect 718 662 721 728
rect 766 682 769 758
rect 774 732 777 738
rect 778 678 782 681
rect 766 672 769 678
rect 750 662 753 668
rect 626 658 630 661
rect 670 658 678 661
rect 738 658 742 661
rect 762 658 766 661
rect 606 642 609 648
rect 638 642 641 648
rect 446 552 449 558
rect 454 552 457 558
rect 518 552 521 578
rect 550 552 553 568
rect 622 562 625 618
rect 662 562 665 608
rect 410 548 414 551
rect 466 548 470 551
rect 366 542 369 548
rect 354 468 358 471
rect 298 458 305 461
rect 294 352 297 368
rect 302 352 305 458
rect 318 452 321 458
rect 326 392 329 448
rect 350 372 353 468
rect 362 438 366 441
rect 374 392 377 498
rect 390 462 393 538
rect 422 463 425 518
rect 438 492 441 548
rect 462 492 465 538
rect 486 502 489 548
rect 454 472 457 488
rect 494 472 497 498
rect 510 492 513 548
rect 390 372 393 458
rect 454 442 457 448
rect 462 392 465 468
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 310 312 313 348
rect 334 322 337 348
rect 302 292 305 298
rect 310 292 313 298
rect 174 222 177 258
rect 262 172 265 258
rect 158 162 161 168
rect 70 151 73 158
rect 118 152 121 158
rect 102 142 105 148
rect 126 142 129 158
rect 146 148 150 151
rect 146 138 150 141
rect 6 72 9 78
rect 70 72 73 128
rect 74 68 78 71
rect 146 68 150 71
rect 158 62 161 158
rect 174 152 177 158
rect 262 151 265 158
rect 206 142 209 148
rect 214 142 217 148
rect 334 142 337 168
rect 194 138 198 141
rect 166 71 169 118
rect 174 102 177 138
rect 214 82 217 138
rect 246 132 249 138
rect 230 122 233 128
rect 322 118 326 121
rect 270 92 273 98
rect 294 82 297 88
rect 166 68 177 71
rect 146 58 150 61
rect 166 52 169 58
rect 174 52 177 68
rect 190 62 193 68
rect 278 62 281 78
rect 318 72 321 78
rect 342 72 345 128
rect 358 122 361 348
rect 374 282 377 368
rect 414 352 417 358
rect 478 352 481 358
rect 394 348 398 351
rect 442 348 446 351
rect 382 342 385 348
rect 402 338 406 341
rect 382 302 385 338
rect 370 259 374 262
rect 390 192 393 268
rect 422 262 425 318
rect 502 292 505 338
rect 486 272 489 278
rect 470 263 473 268
rect 502 262 505 288
rect 410 228 414 231
rect 470 192 473 218
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 434 188 438 191
rect 486 152 489 178
rect 510 152 513 438
rect 526 432 529 548
rect 566 542 569 548
rect 574 542 577 558
rect 638 552 641 558
rect 618 548 622 551
rect 662 542 665 548
rect 618 538 622 541
rect 634 538 638 541
rect 602 528 606 531
rect 582 522 585 528
rect 606 502 609 518
rect 518 362 521 368
rect 518 262 521 348
rect 526 332 529 338
rect 526 252 529 258
rect 534 172 537 468
rect 582 463 585 498
rect 598 452 601 468
rect 622 462 625 468
rect 646 462 649 468
rect 550 372 553 418
rect 582 392 585 438
rect 670 392 673 658
rect 686 652 689 658
rect 726 572 729 618
rect 782 592 785 668
rect 790 662 793 828
rect 806 742 809 858
rect 846 852 849 868
rect 850 848 854 851
rect 822 832 825 848
rect 862 842 865 868
rect 870 852 873 988
rect 878 942 881 1128
rect 894 952 897 1008
rect 902 1002 905 1198
rect 910 1152 913 1288
rect 934 1262 937 1288
rect 942 1262 945 1268
rect 950 1262 953 1438
rect 958 1352 961 1458
rect 1030 1342 1033 1568
rect 1118 1552 1121 1638
rect 1142 1612 1145 1658
rect 1182 1652 1185 1748
rect 1190 1712 1193 1738
rect 1190 1672 1193 1688
rect 1174 1612 1177 1648
rect 1126 1592 1129 1598
rect 1182 1582 1185 1648
rect 1058 1548 1062 1551
rect 1178 1548 1182 1551
rect 1038 1542 1041 1548
rect 1094 1542 1097 1548
rect 1150 1542 1153 1548
rect 1074 1538 1078 1541
rect 1134 1532 1137 1538
rect 1054 1502 1057 1528
rect 1082 1518 1086 1521
rect 1070 1492 1073 1518
rect 1110 1512 1113 1528
rect 1166 1492 1169 1498
rect 1086 1472 1089 1478
rect 1102 1463 1105 1468
rect 1182 1462 1185 1498
rect 1174 1432 1177 1458
rect 1058 1348 1062 1351
rect 1046 1342 1049 1348
rect 994 1318 998 1321
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 1014 1288 1022 1291
rect 1014 1282 1017 1288
rect 1022 1272 1025 1278
rect 1006 1262 1009 1268
rect 1014 1262 1017 1268
rect 978 1258 982 1261
rect 926 1092 929 1248
rect 942 1192 945 1258
rect 950 1232 953 1258
rect 934 1121 937 1168
rect 942 1152 945 1168
rect 950 1142 953 1198
rect 958 1152 961 1258
rect 1014 1202 1017 1258
rect 1030 1232 1033 1338
rect 966 1142 969 1148
rect 934 1118 945 1121
rect 930 1088 934 1091
rect 942 1072 945 1118
rect 950 1062 953 1068
rect 878 932 881 938
rect 878 892 881 928
rect 902 892 905 958
rect 902 882 905 888
rect 886 852 889 858
rect 894 852 897 868
rect 918 862 921 1058
rect 966 1052 969 1118
rect 974 1072 977 1158
rect 990 1152 993 1158
rect 1030 1152 1033 1228
rect 1038 1222 1041 1268
rect 1050 1258 1054 1261
rect 1026 1148 1030 1151
rect 1002 1128 1006 1131
rect 1038 1122 1041 1218
rect 1046 1152 1049 1168
rect 1054 1141 1057 1218
rect 1070 1162 1073 1388
rect 1118 1372 1121 1398
rect 1086 1262 1089 1268
rect 1094 1262 1097 1368
rect 1118 1342 1121 1368
rect 1138 1358 1142 1361
rect 1158 1352 1161 1358
rect 1134 1342 1137 1348
rect 1102 1262 1105 1268
rect 1134 1262 1137 1318
rect 1158 1302 1161 1348
rect 1166 1342 1169 1418
rect 1190 1351 1193 1418
rect 1198 1362 1201 1758
rect 1214 1742 1217 1778
rect 1254 1752 1257 1878
rect 1270 1872 1273 1938
rect 1294 1912 1297 1918
rect 1310 1892 1313 1948
rect 1318 1942 1321 1948
rect 1334 1892 1337 2048
rect 1350 1952 1353 1968
rect 1366 1952 1369 2008
rect 1398 1982 1401 2058
rect 1438 2022 1441 2058
rect 1446 2002 1449 2078
rect 1478 2062 1481 2068
rect 1486 2062 1489 2108
rect 1498 2068 1502 2071
rect 1478 2022 1481 2058
rect 1496 2003 1498 2007
rect 1502 2003 1505 2007
rect 1509 2003 1512 2007
rect 1414 1952 1417 1978
rect 1402 1948 1406 1951
rect 1434 1948 1438 1951
rect 1466 1948 1470 1951
rect 1262 1862 1265 1868
rect 1310 1862 1313 1868
rect 1318 1862 1321 1888
rect 1330 1848 1334 1851
rect 1350 1792 1353 1818
rect 1262 1752 1265 1758
rect 1294 1752 1297 1758
rect 1350 1752 1353 1758
rect 1278 1732 1281 1738
rect 1230 1712 1233 1718
rect 1222 1692 1225 1698
rect 1246 1672 1249 1688
rect 1286 1682 1289 1748
rect 1302 1742 1305 1748
rect 1314 1738 1318 1741
rect 1294 1672 1297 1708
rect 1310 1692 1313 1718
rect 1238 1662 1241 1668
rect 1246 1662 1249 1668
rect 1226 1658 1230 1661
rect 1282 1658 1286 1661
rect 1238 1622 1241 1658
rect 1262 1652 1265 1658
rect 1262 1572 1265 1648
rect 1286 1642 1289 1648
rect 1294 1601 1297 1668
rect 1302 1632 1305 1648
rect 1286 1598 1297 1601
rect 1238 1552 1241 1568
rect 1250 1558 1254 1561
rect 1278 1552 1281 1558
rect 1238 1542 1241 1548
rect 1286 1542 1289 1598
rect 1310 1592 1313 1678
rect 1318 1672 1321 1718
rect 1326 1692 1329 1698
rect 1334 1592 1337 1748
rect 1358 1592 1361 1948
rect 1446 1942 1449 1948
rect 1458 1938 1465 1941
rect 1374 1932 1377 1938
rect 1390 1842 1393 1918
rect 1414 1882 1417 1918
rect 1446 1892 1449 1898
rect 1402 1868 1406 1871
rect 1450 1868 1454 1871
rect 1430 1862 1433 1868
rect 1462 1862 1465 1938
rect 1478 1932 1481 1958
rect 1526 1942 1529 1947
rect 1534 1942 1537 2138
rect 1566 2112 1569 2138
rect 1590 2072 1593 2118
rect 1598 2082 1601 2088
rect 1542 2062 1545 2068
rect 1606 2062 1609 2098
rect 1614 2082 1617 2138
rect 1622 2112 1625 2138
rect 1670 2122 1673 2138
rect 1614 2062 1617 2078
rect 1654 2072 1657 2108
rect 1670 2072 1673 2118
rect 1702 2072 1705 2078
rect 1682 2068 1686 2071
rect 1638 2062 1641 2068
rect 1566 2012 1569 2058
rect 1606 1992 1609 2058
rect 1662 2042 1665 2058
rect 1686 2042 1689 2048
rect 1614 1972 1617 2008
rect 1630 1982 1633 2018
rect 1602 1968 1606 1971
rect 1662 1951 1665 1978
rect 1490 1938 1494 1941
rect 1474 1888 1478 1891
rect 1522 1888 1526 1891
rect 1486 1872 1489 1888
rect 1534 1872 1537 1908
rect 1522 1868 1526 1871
rect 1542 1862 1545 1868
rect 1550 1862 1553 1878
rect 1506 1858 1510 1861
rect 1382 1752 1385 1798
rect 1414 1792 1417 1858
rect 1430 1812 1433 1858
rect 1462 1852 1465 1858
rect 1470 1842 1473 1848
rect 1478 1761 1481 1838
rect 1496 1803 1498 1807
rect 1502 1803 1505 1807
rect 1509 1803 1512 1807
rect 1558 1792 1561 1938
rect 1574 1852 1577 1948
rect 1694 1942 1697 1968
rect 1710 1952 1713 1958
rect 1582 1892 1585 1928
rect 1594 1918 1601 1921
rect 1598 1872 1601 1918
rect 1658 1888 1662 1891
rect 1606 1872 1609 1888
rect 1626 1868 1630 1871
rect 1582 1862 1585 1868
rect 1578 1848 1582 1851
rect 1566 1822 1569 1848
rect 1470 1758 1481 1761
rect 1498 1758 1502 1761
rect 1470 1752 1473 1758
rect 1450 1748 1454 1751
rect 1374 1742 1377 1748
rect 1398 1722 1401 1748
rect 1422 1732 1425 1748
rect 1422 1672 1425 1678
rect 1294 1552 1297 1588
rect 1302 1552 1305 1558
rect 1330 1548 1334 1551
rect 1258 1538 1262 1541
rect 1214 1462 1217 1498
rect 1230 1472 1233 1478
rect 1186 1348 1193 1351
rect 1206 1352 1209 1378
rect 1214 1352 1217 1448
rect 1190 1282 1193 1318
rect 1198 1272 1201 1288
rect 1146 1268 1150 1271
rect 1182 1262 1185 1268
rect 1110 1252 1113 1258
rect 1102 1192 1105 1218
rect 1142 1192 1145 1258
rect 1150 1252 1153 1258
rect 1178 1248 1182 1251
rect 1066 1158 1070 1161
rect 1086 1152 1089 1158
rect 1050 1138 1057 1141
rect 1078 1142 1081 1148
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 1006 1092 1009 1118
rect 1038 1072 1041 1108
rect 986 1048 990 1051
rect 950 1012 953 1018
rect 934 992 937 998
rect 950 992 953 998
rect 962 958 966 961
rect 942 892 945 958
rect 942 872 945 888
rect 814 752 817 768
rect 830 712 833 818
rect 870 731 873 848
rect 886 822 889 848
rect 878 752 881 778
rect 886 742 889 778
rect 894 742 897 848
rect 910 782 913 838
rect 910 752 913 768
rect 918 762 921 848
rect 926 812 929 818
rect 942 772 945 858
rect 950 822 953 918
rect 958 892 961 948
rect 966 942 969 948
rect 966 922 969 938
rect 966 892 969 898
rect 974 892 977 1048
rect 982 982 985 1018
rect 998 992 1001 1068
rect 1038 1062 1041 1068
rect 1034 1048 1038 1051
rect 982 942 985 978
rect 998 942 1001 968
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 958 871 961 888
rect 1006 872 1009 1048
rect 1014 952 1017 1038
rect 1022 952 1025 958
rect 1030 952 1033 958
rect 1026 938 1030 941
rect 1022 892 1025 908
rect 1046 892 1049 1128
rect 1054 1102 1057 1118
rect 1054 1072 1057 1098
rect 1078 1092 1081 1118
rect 1086 1092 1089 1148
rect 1094 1142 1097 1178
rect 1138 1148 1142 1151
rect 1150 1132 1153 1248
rect 1158 1212 1161 1218
rect 1214 1212 1217 1348
rect 1222 1322 1225 1338
rect 1230 1282 1233 1468
rect 1246 1463 1249 1518
rect 1294 1472 1297 1548
rect 1374 1542 1377 1668
rect 1382 1652 1385 1658
rect 1422 1652 1425 1658
rect 1422 1562 1425 1648
rect 1430 1632 1433 1748
rect 1438 1742 1441 1748
rect 1478 1712 1481 1748
rect 1486 1742 1489 1748
rect 1518 1682 1521 1788
rect 1546 1758 1550 1761
rect 1538 1748 1542 1751
rect 1550 1742 1553 1748
rect 1558 1742 1561 1768
rect 1566 1752 1569 1818
rect 1590 1752 1593 1788
rect 1598 1762 1601 1868
rect 1606 1842 1609 1868
rect 1654 1862 1657 1868
rect 1614 1852 1617 1858
rect 1650 1848 1654 1851
rect 1678 1842 1681 1938
rect 1698 1858 1702 1861
rect 1622 1822 1625 1838
rect 1662 1752 1665 1758
rect 1686 1752 1689 1758
rect 1610 1748 1614 1751
rect 1654 1732 1657 1738
rect 1694 1732 1697 1748
rect 1702 1742 1705 1748
rect 1710 1742 1713 1948
rect 1718 1872 1721 2068
rect 1734 2063 1737 2068
rect 1726 1952 1729 2008
rect 1758 1992 1761 2248
rect 1854 2242 1857 2338
rect 1862 2262 1865 2288
rect 1878 2262 1881 2298
rect 1782 2192 1785 2218
rect 1830 2192 1833 2228
rect 1802 2148 1806 2151
rect 1806 2132 1809 2138
rect 1766 2112 1769 2118
rect 1814 2092 1817 2138
rect 1798 2082 1801 2088
rect 1734 1972 1737 1978
rect 1730 1948 1734 1951
rect 1742 1882 1745 1938
rect 1742 1812 1745 1868
rect 1766 1862 1769 2078
rect 1806 2052 1809 2078
rect 1822 2061 1825 2118
rect 1822 2058 1830 2061
rect 1838 1992 1841 2068
rect 1846 2062 1849 2218
rect 1878 2142 1881 2148
rect 1886 2142 1889 2338
rect 1902 2292 1905 2318
rect 1910 2312 1913 2338
rect 1894 2262 1897 2278
rect 1902 2262 1905 2278
rect 1958 2272 1961 2308
rect 1990 2292 1993 2328
rect 2016 2303 2018 2307
rect 2022 2303 2025 2307
rect 2029 2303 2032 2307
rect 2046 2292 2049 2348
rect 2054 2342 2057 2368
rect 2210 2358 2214 2361
rect 2070 2352 2073 2358
rect 2086 2352 2089 2358
rect 2094 2352 2097 2358
rect 2266 2348 2270 2351
rect 2362 2348 2366 2351
rect 2054 2322 2057 2338
rect 2102 2332 2105 2338
rect 2014 2272 2017 2278
rect 2038 2272 2041 2278
rect 1926 2262 1929 2268
rect 1950 2262 1953 2268
rect 1910 2102 1913 2258
rect 1918 2182 1921 2258
rect 1958 2222 1961 2268
rect 1970 2258 1974 2261
rect 1998 2252 2001 2258
rect 2050 2248 2054 2251
rect 1926 2132 1929 2138
rect 1934 2092 1937 2218
rect 1974 2182 1977 2238
rect 1978 2178 1982 2181
rect 1946 2088 1950 2091
rect 1870 2062 1873 2068
rect 1886 2062 1889 2078
rect 1898 2068 1902 2071
rect 1878 2032 1881 2058
rect 1862 1982 1865 2018
rect 1818 1958 1822 1961
rect 1858 1958 1886 1961
rect 1910 1952 1913 2088
rect 1958 2082 1961 2088
rect 1950 2072 1953 2078
rect 1990 2072 1993 2218
rect 1998 2152 2001 2238
rect 2054 2152 2057 2158
rect 2078 2152 2081 2158
rect 2046 2142 2049 2148
rect 2016 2103 2018 2107
rect 2022 2103 2025 2107
rect 2029 2103 2032 2107
rect 2022 2082 2025 2088
rect 1918 2062 1921 2068
rect 1974 2062 1977 2068
rect 1938 2058 1942 2061
rect 1994 2058 1998 2061
rect 1926 2052 1929 2058
rect 1966 2052 1969 2058
rect 1950 1952 1953 1998
rect 1998 1962 2001 2018
rect 1930 1948 1934 1951
rect 1818 1938 1822 1941
rect 1790 1862 1793 1888
rect 1802 1868 1806 1871
rect 1834 1868 1838 1871
rect 1718 1772 1721 1788
rect 1758 1782 1761 1858
rect 1814 1842 1817 1858
rect 1838 1842 1841 1848
rect 1778 1828 1782 1831
rect 1846 1812 1849 1938
rect 1870 1892 1873 1938
rect 1878 1922 1881 1948
rect 1886 1922 1889 1938
rect 1902 1912 1905 1938
rect 1898 1888 1902 1891
rect 1862 1872 1865 1888
rect 1870 1872 1873 1878
rect 1886 1862 1889 1868
rect 1742 1772 1745 1778
rect 1774 1772 1777 1808
rect 1718 1762 1721 1768
rect 1758 1762 1761 1768
rect 1718 1752 1721 1758
rect 1806 1752 1809 1768
rect 1738 1748 1742 1751
rect 1750 1742 1753 1748
rect 1446 1662 1449 1668
rect 1498 1658 1502 1661
rect 1562 1658 1566 1661
rect 1602 1658 1606 1661
rect 1446 1592 1449 1648
rect 1310 1492 1313 1498
rect 1326 1462 1329 1488
rect 1350 1462 1353 1478
rect 1358 1462 1361 1508
rect 1382 1492 1385 1548
rect 1398 1512 1401 1548
rect 1430 1542 1433 1568
rect 1442 1558 1446 1561
rect 1454 1552 1457 1618
rect 1496 1603 1498 1607
rect 1502 1603 1505 1607
rect 1509 1603 1512 1607
rect 1526 1592 1529 1608
rect 1482 1558 1486 1561
rect 1542 1552 1545 1618
rect 1574 1612 1577 1658
rect 1614 1652 1617 1658
rect 1622 1642 1625 1648
rect 1598 1572 1601 1618
rect 1586 1558 1590 1561
rect 1558 1552 1561 1558
rect 1454 1542 1457 1548
rect 1478 1542 1481 1548
rect 1466 1538 1470 1541
rect 1534 1532 1537 1548
rect 1366 1482 1369 1488
rect 1430 1463 1433 1468
rect 1246 1458 1249 1459
rect 1238 1352 1241 1358
rect 1258 1348 1262 1351
rect 1270 1342 1273 1408
rect 1334 1382 1337 1418
rect 1358 1362 1361 1458
rect 1266 1338 1270 1341
rect 1274 1318 1278 1321
rect 1246 1312 1249 1318
rect 1290 1288 1294 1291
rect 1110 1072 1113 1108
rect 1134 1072 1137 1078
rect 1054 1052 1057 1058
rect 1062 1042 1065 1068
rect 1102 1052 1105 1068
rect 1074 1048 1078 1051
rect 1114 1048 1118 1051
rect 1078 1022 1081 1048
rect 1066 947 1070 950
rect 1030 872 1033 888
rect 958 868 966 871
rect 958 852 961 858
rect 1018 848 1022 851
rect 966 842 969 848
rect 950 792 953 798
rect 942 762 945 768
rect 930 758 934 761
rect 922 738 926 741
rect 954 738 958 741
rect 870 728 881 731
rect 830 672 833 678
rect 854 672 857 728
rect 866 718 870 721
rect 878 682 881 728
rect 902 722 905 738
rect 894 702 897 718
rect 926 702 929 718
rect 910 672 913 688
rect 898 668 902 671
rect 918 662 921 678
rect 930 668 934 671
rect 818 658 822 661
rect 890 658 897 661
rect 906 658 910 661
rect 790 652 793 658
rect 798 652 801 658
rect 806 582 809 658
rect 846 652 849 658
rect 862 652 865 658
rect 878 622 881 628
rect 850 588 854 591
rect 774 562 777 568
rect 678 542 681 558
rect 814 552 817 568
rect 870 552 873 558
rect 878 552 881 598
rect 894 592 897 658
rect 942 652 945 738
rect 966 692 969 738
rect 958 682 961 688
rect 938 648 942 651
rect 942 592 945 648
rect 966 552 969 618
rect 714 547 718 550
rect 802 548 806 551
rect 834 548 838 551
rect 914 548 918 551
rect 954 548 958 551
rect 694 492 697 538
rect 790 492 793 548
rect 706 488 710 491
rect 710 472 713 478
rect 758 472 761 488
rect 730 468 734 471
rect 710 392 713 468
rect 722 458 726 461
rect 742 452 745 458
rect 774 452 777 468
rect 798 462 801 468
rect 550 352 553 368
rect 558 352 561 358
rect 726 352 729 378
rect 666 348 670 351
rect 698 348 702 351
rect 566 342 569 348
rect 542 292 545 338
rect 550 332 553 338
rect 566 272 569 328
rect 614 302 617 348
rect 638 322 641 348
rect 586 268 590 271
rect 550 242 553 258
rect 430 92 433 118
rect 418 88 422 91
rect 438 82 441 138
rect 446 102 449 148
rect 326 62 329 68
rect 206 52 209 59
rect 310 52 313 58
rect 358 52 361 59
rect 422 -18 425 78
rect 478 72 481 148
rect 534 142 537 168
rect 526 101 529 118
rect 518 98 529 101
rect 494 72 497 88
rect 434 68 438 71
rect 458 68 462 71
rect 434 58 438 61
rect 462 52 465 58
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
rect 518 -18 521 98
rect 534 72 537 138
rect 566 122 569 268
rect 578 258 582 261
rect 602 248 606 251
rect 598 142 601 148
rect 606 142 609 238
rect 614 232 617 268
rect 646 232 649 348
rect 662 272 665 278
rect 654 262 657 268
rect 614 152 617 228
rect 646 182 649 228
rect 622 162 625 168
rect 646 152 649 168
rect 654 152 657 158
rect 606 91 609 138
rect 602 88 609 91
rect 582 72 585 78
rect 558 62 561 68
rect 638 62 641 138
rect 654 122 657 138
rect 662 82 665 268
rect 678 192 681 348
rect 686 312 689 348
rect 766 342 769 348
rect 774 342 777 448
rect 822 442 825 548
rect 862 542 865 548
rect 854 492 857 528
rect 822 352 825 368
rect 846 362 849 448
rect 834 338 841 341
rect 734 292 737 308
rect 710 262 713 288
rect 758 262 761 278
rect 766 262 769 268
rect 730 258 734 261
rect 702 152 705 208
rect 694 132 697 148
rect 718 142 721 148
rect 742 142 745 148
rect 750 122 753 258
rect 774 241 777 338
rect 786 268 790 271
rect 806 262 809 268
rect 782 252 785 258
rect 774 238 785 241
rect 782 172 785 238
rect 806 162 809 168
rect 806 142 809 158
rect 710 92 713 118
rect 678 62 681 68
rect 694 62 697 88
rect 782 82 785 128
rect 814 92 817 268
rect 822 162 825 288
rect 830 262 833 328
rect 838 292 841 338
rect 846 332 849 358
rect 854 352 857 368
rect 838 262 841 268
rect 846 252 849 318
rect 854 311 857 348
rect 862 342 865 408
rect 870 362 873 548
rect 886 542 889 548
rect 926 542 929 548
rect 926 512 929 538
rect 934 532 937 548
rect 922 488 926 491
rect 882 468 886 471
rect 914 468 921 471
rect 906 458 910 461
rect 878 452 881 458
rect 902 352 905 408
rect 918 372 921 468
rect 926 352 929 488
rect 934 392 937 448
rect 950 352 953 428
rect 974 422 977 818
rect 982 762 985 778
rect 982 752 985 758
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 1006 662 1009 718
rect 1014 642 1017 818
rect 1022 792 1025 848
rect 1022 752 1025 778
rect 1030 762 1033 868
rect 1046 842 1049 848
rect 1038 772 1041 818
rect 1046 752 1049 758
rect 1030 748 1038 751
rect 1030 742 1033 748
rect 1062 742 1065 928
rect 1078 882 1081 928
rect 1078 792 1081 848
rect 1094 762 1097 1018
rect 1110 1002 1113 1048
rect 1126 1022 1129 1048
rect 1142 1012 1145 1108
rect 1150 1092 1153 1128
rect 1122 968 1126 971
rect 1134 942 1137 988
rect 1150 962 1153 1018
rect 1150 942 1153 958
rect 1158 952 1161 1208
rect 1230 1152 1233 1278
rect 1238 1262 1241 1268
rect 1302 1162 1305 1218
rect 1182 1142 1185 1148
rect 1198 1112 1201 1118
rect 1190 1092 1193 1098
rect 1166 992 1169 998
rect 1102 852 1105 858
rect 1086 742 1089 758
rect 1074 738 1078 741
rect 994 568 998 571
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 998 472 1001 478
rect 1014 472 1017 488
rect 982 463 985 468
rect 938 348 942 351
rect 870 332 873 338
rect 886 332 889 348
rect 918 332 921 348
rect 890 328 894 331
rect 854 308 865 311
rect 854 292 857 298
rect 822 152 825 158
rect 842 148 846 151
rect 862 142 865 308
rect 898 258 902 261
rect 950 212 953 348
rect 966 342 969 368
rect 974 352 977 418
rect 1022 392 1025 718
rect 1030 532 1033 738
rect 1038 732 1041 738
rect 1046 682 1049 738
rect 1062 702 1065 718
rect 1066 678 1070 681
rect 1046 672 1049 678
rect 1070 652 1073 658
rect 1078 652 1081 668
rect 1086 582 1089 718
rect 1094 692 1097 748
rect 1094 662 1097 668
rect 1094 652 1097 658
rect 1102 572 1105 768
rect 1126 762 1129 938
rect 1134 802 1137 938
rect 1142 872 1145 888
rect 1150 872 1153 878
rect 1158 862 1161 948
rect 1174 932 1177 958
rect 1190 952 1193 968
rect 1198 952 1201 1108
rect 1206 1072 1209 1128
rect 1222 1072 1225 1108
rect 1230 1102 1233 1138
rect 1254 1092 1257 1148
rect 1294 1122 1297 1138
rect 1242 1048 1246 1051
rect 1214 992 1217 1018
rect 1222 952 1225 1018
rect 1210 948 1214 951
rect 1166 892 1169 918
rect 1174 902 1177 928
rect 1222 922 1225 948
rect 1230 941 1233 1048
rect 1230 940 1238 941
rect 1242 940 1246 943
rect 1262 942 1265 1078
rect 1286 1072 1289 1098
rect 1310 1092 1313 1298
rect 1270 1052 1273 1058
rect 1270 982 1273 1048
rect 1278 971 1281 1068
rect 1318 1052 1321 1318
rect 1334 1312 1337 1348
rect 1342 1272 1345 1328
rect 1382 1312 1385 1338
rect 1350 1192 1353 1308
rect 1398 1292 1401 1458
rect 1382 1272 1385 1288
rect 1422 1282 1425 1348
rect 1418 1268 1422 1271
rect 1366 1263 1369 1268
rect 1366 1258 1369 1259
rect 1374 1152 1377 1158
rect 1366 1142 1369 1148
rect 1334 1072 1337 1098
rect 1342 1092 1345 1128
rect 1314 1048 1318 1051
rect 1270 968 1281 971
rect 1294 1022 1297 1028
rect 1230 938 1241 940
rect 1206 902 1209 918
rect 1230 892 1233 918
rect 1166 852 1169 858
rect 1182 852 1185 858
rect 1198 852 1201 868
rect 1206 862 1209 868
rect 1214 852 1217 858
rect 1174 752 1177 758
rect 1182 752 1185 808
rect 1206 762 1209 828
rect 1154 748 1158 751
rect 1110 692 1113 748
rect 1118 722 1121 728
rect 1134 722 1137 728
rect 1122 658 1126 661
rect 1134 661 1137 718
rect 1142 672 1145 678
rect 1150 662 1153 728
rect 1158 712 1161 718
rect 1162 678 1166 681
rect 1174 672 1177 738
rect 1182 692 1185 748
rect 1194 738 1198 741
rect 1194 688 1198 691
rect 1134 658 1145 661
rect 1130 648 1134 651
rect 1054 551 1057 558
rect 1086 542 1089 568
rect 1102 562 1105 568
rect 1118 562 1121 648
rect 1126 552 1129 568
rect 1102 542 1105 548
rect 1070 472 1073 538
rect 1078 472 1081 508
rect 1094 492 1097 528
rect 1134 512 1137 538
rect 1142 532 1145 658
rect 1158 642 1161 668
rect 1182 652 1185 658
rect 1206 612 1209 758
rect 1222 752 1225 818
rect 1238 761 1241 938
rect 1254 932 1257 938
rect 1254 872 1257 878
rect 1246 862 1249 868
rect 1262 862 1265 918
rect 1270 882 1273 968
rect 1258 858 1262 861
rect 1270 852 1273 858
rect 1230 758 1241 761
rect 1278 762 1281 898
rect 1294 882 1297 1018
rect 1302 1012 1305 1048
rect 1318 932 1321 1018
rect 1310 872 1313 888
rect 1298 868 1302 871
rect 1318 862 1321 918
rect 1326 912 1329 1038
rect 1334 942 1337 1068
rect 1342 992 1345 1068
rect 1350 1052 1353 1098
rect 1358 1092 1361 1108
rect 1390 1101 1393 1208
rect 1398 1162 1401 1268
rect 1414 1222 1417 1248
rect 1430 1162 1433 1418
rect 1462 1412 1465 1468
rect 1470 1452 1473 1458
rect 1478 1452 1481 1518
rect 1530 1488 1534 1491
rect 1494 1472 1497 1478
rect 1486 1462 1489 1468
rect 1510 1452 1513 1458
rect 1530 1448 1534 1451
rect 1542 1411 1545 1548
rect 1598 1542 1601 1568
rect 1638 1562 1641 1668
rect 1646 1662 1649 1688
rect 1654 1672 1657 1698
rect 1682 1668 1686 1671
rect 1702 1662 1705 1668
rect 1710 1662 1713 1668
rect 1654 1652 1657 1658
rect 1682 1648 1686 1651
rect 1578 1538 1582 1541
rect 1550 1481 1553 1538
rect 1550 1478 1558 1481
rect 1558 1472 1561 1478
rect 1594 1468 1598 1471
rect 1550 1422 1553 1458
rect 1558 1452 1561 1458
rect 1542 1408 1553 1411
rect 1496 1403 1498 1407
rect 1502 1403 1505 1407
rect 1509 1403 1512 1407
rect 1550 1382 1553 1408
rect 1558 1392 1561 1448
rect 1454 1272 1457 1298
rect 1438 1262 1441 1268
rect 1462 1262 1465 1358
rect 1470 1342 1473 1368
rect 1482 1358 1486 1361
rect 1550 1352 1553 1378
rect 1566 1352 1569 1468
rect 1594 1448 1598 1451
rect 1538 1348 1542 1351
rect 1486 1342 1489 1348
rect 1474 1338 1478 1341
rect 1470 1272 1473 1278
rect 1438 1222 1441 1258
rect 1462 1172 1465 1258
rect 1478 1252 1481 1318
rect 1502 1292 1505 1348
rect 1550 1342 1553 1348
rect 1502 1282 1505 1288
rect 1496 1203 1498 1207
rect 1502 1203 1505 1207
rect 1509 1203 1512 1207
rect 1434 1158 1438 1161
rect 1462 1152 1465 1158
rect 1518 1152 1521 1308
rect 1534 1242 1537 1318
rect 1566 1312 1569 1338
rect 1542 1272 1545 1288
rect 1582 1272 1585 1418
rect 1590 1342 1593 1348
rect 1598 1272 1601 1278
rect 1562 1259 1566 1262
rect 1606 1252 1609 1558
rect 1614 1472 1617 1488
rect 1630 1472 1633 1508
rect 1646 1463 1649 1468
rect 1646 1352 1649 1368
rect 1654 1362 1657 1648
rect 1718 1622 1721 1658
rect 1662 1542 1665 1548
rect 1718 1542 1721 1558
rect 1726 1542 1729 1698
rect 1814 1692 1817 1808
rect 1854 1752 1857 1858
rect 1862 1842 1865 1858
rect 1894 1842 1897 1858
rect 1838 1742 1841 1748
rect 1778 1688 1782 1691
rect 1742 1662 1745 1678
rect 1822 1672 1825 1688
rect 1830 1682 1833 1688
rect 1750 1662 1753 1668
rect 1738 1658 1742 1661
rect 1770 1658 1774 1661
rect 1758 1652 1761 1658
rect 1798 1592 1801 1658
rect 1806 1642 1809 1648
rect 1734 1552 1737 1568
rect 1758 1562 1761 1568
rect 1750 1542 1753 1558
rect 1822 1552 1825 1558
rect 1778 1548 1782 1551
rect 1790 1542 1793 1548
rect 1830 1542 1833 1568
rect 1778 1538 1782 1541
rect 1686 1502 1689 1538
rect 1702 1532 1705 1538
rect 1706 1488 1710 1491
rect 1662 1352 1665 1488
rect 1678 1462 1681 1468
rect 1718 1452 1721 1518
rect 1726 1482 1729 1538
rect 1734 1462 1737 1538
rect 1750 1492 1753 1528
rect 1742 1472 1745 1478
rect 1726 1452 1729 1458
rect 1678 1362 1681 1368
rect 1718 1352 1721 1358
rect 1690 1348 1694 1351
rect 1646 1272 1649 1298
rect 1654 1292 1657 1348
rect 1722 1338 1726 1341
rect 1614 1262 1617 1268
rect 1638 1252 1641 1258
rect 1610 1248 1614 1251
rect 1582 1162 1585 1168
rect 1398 1112 1401 1148
rect 1390 1098 1401 1101
rect 1350 1042 1353 1048
rect 1366 992 1369 1048
rect 1398 992 1401 1098
rect 1406 1042 1409 1138
rect 1422 1082 1425 1118
rect 1422 1052 1425 1059
rect 1438 1052 1441 1118
rect 1350 952 1353 958
rect 1386 948 1390 951
rect 1418 948 1422 951
rect 1338 938 1342 941
rect 1286 852 1289 858
rect 1230 752 1233 758
rect 1290 748 1294 751
rect 1230 722 1233 728
rect 1238 692 1241 748
rect 1246 732 1249 738
rect 1222 662 1225 668
rect 1254 663 1257 668
rect 1254 658 1257 659
rect 1154 588 1158 591
rect 1142 502 1145 528
rect 1126 482 1129 488
rect 1038 468 1046 471
rect 1038 462 1041 468
rect 1074 458 1078 461
rect 1046 452 1049 458
rect 1110 442 1113 458
rect 1110 382 1113 438
rect 982 352 985 378
rect 1058 348 1062 351
rect 966 332 969 338
rect 1014 322 1017 348
rect 1038 331 1041 348
rect 1046 342 1049 348
rect 1078 342 1081 358
rect 1086 352 1089 358
rect 1102 342 1105 368
rect 1134 351 1137 358
rect 1054 332 1057 338
rect 1038 328 1049 331
rect 966 292 969 318
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 970 288 974 291
rect 958 262 961 268
rect 998 262 1001 268
rect 1030 263 1033 268
rect 886 192 889 198
rect 958 192 961 258
rect 902 142 905 178
rect 998 152 1001 158
rect 1030 152 1033 158
rect 1022 142 1025 148
rect 826 138 830 141
rect 894 101 897 138
rect 1010 128 1014 131
rect 1038 122 1041 148
rect 1046 142 1049 328
rect 1062 272 1065 288
rect 1110 272 1113 278
rect 1118 272 1121 328
rect 1142 282 1145 288
rect 1082 268 1086 271
rect 1102 262 1105 268
rect 1078 252 1081 258
rect 1070 152 1073 178
rect 1078 152 1081 228
rect 1086 152 1089 168
rect 1098 158 1102 161
rect 1086 142 1089 148
rect 886 98 897 101
rect 734 72 737 78
rect 870 72 873 88
rect 842 68 846 71
rect 758 62 761 68
rect 862 62 865 68
rect 874 58 878 61
rect 862 52 865 58
rect 842 48 846 51
rect 422 -22 426 -18
rect 518 -22 522 -18
rect 878 -19 882 -18
rect 886 -19 889 98
rect 910 92 913 118
rect 894 82 897 88
rect 958 82 961 118
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 958 72 961 78
rect 1006 72 1009 118
rect 1070 72 1073 88
rect 1078 72 1081 78
rect 1110 72 1113 258
rect 1118 192 1121 268
rect 1150 262 1153 578
rect 1182 562 1185 568
rect 1170 558 1174 561
rect 1206 552 1209 568
rect 1182 532 1185 538
rect 1202 528 1206 531
rect 1214 521 1217 548
rect 1206 518 1217 521
rect 1190 472 1193 508
rect 1182 372 1185 468
rect 1198 462 1201 518
rect 1206 452 1209 518
rect 1222 482 1225 658
rect 1270 642 1273 748
rect 1278 722 1281 748
rect 1310 742 1313 768
rect 1326 752 1329 898
rect 1342 862 1345 868
rect 1350 852 1353 858
rect 1334 752 1337 758
rect 1346 748 1350 751
rect 1318 742 1321 748
rect 1294 732 1297 738
rect 1294 712 1297 718
rect 1286 672 1289 688
rect 1306 668 1310 671
rect 1326 662 1329 708
rect 1334 672 1337 678
rect 1358 672 1361 888
rect 1366 782 1369 918
rect 1366 752 1369 758
rect 1374 742 1377 788
rect 1390 752 1393 938
rect 1398 932 1401 938
rect 1406 872 1409 888
rect 1398 838 1406 841
rect 1398 792 1401 838
rect 1414 792 1417 938
rect 1430 922 1433 928
rect 1430 902 1433 918
rect 1422 762 1425 798
rect 1386 748 1390 751
rect 1406 742 1409 748
rect 1414 712 1417 718
rect 1422 712 1425 758
rect 1430 752 1433 758
rect 1438 702 1441 778
rect 1354 668 1358 671
rect 1374 662 1377 668
rect 1362 658 1366 661
rect 1302 652 1305 658
rect 1230 592 1233 638
rect 1254 562 1257 598
rect 1238 532 1241 548
rect 1270 542 1273 638
rect 1294 602 1297 628
rect 1294 552 1297 598
rect 1374 592 1377 658
rect 1390 612 1393 678
rect 1426 659 1430 661
rect 1422 658 1430 659
rect 1398 592 1401 638
rect 1282 548 1286 551
rect 1334 551 1337 558
rect 1218 468 1222 471
rect 1222 452 1225 458
rect 1238 442 1241 468
rect 1278 462 1281 478
rect 1194 368 1198 371
rect 1206 352 1209 418
rect 1222 392 1225 398
rect 1214 352 1217 368
rect 1238 352 1241 438
rect 1286 352 1289 368
rect 1294 352 1297 538
rect 1302 512 1305 538
rect 1334 511 1337 528
rect 1406 512 1409 548
rect 1418 538 1422 541
rect 1326 508 1337 511
rect 1326 472 1329 508
rect 1358 492 1361 508
rect 1382 482 1385 498
rect 1378 468 1382 471
rect 1302 462 1305 468
rect 1390 461 1393 468
rect 1382 458 1393 461
rect 1422 463 1425 518
rect 1342 442 1345 458
rect 1342 382 1345 438
rect 1306 368 1310 371
rect 1298 348 1302 351
rect 1130 258 1134 261
rect 1150 252 1153 258
rect 1158 172 1161 348
rect 1262 292 1265 348
rect 1366 342 1369 347
rect 1382 342 1385 458
rect 1390 442 1393 448
rect 1398 342 1401 368
rect 1414 362 1417 388
rect 1422 342 1425 448
rect 1430 392 1433 638
rect 1438 552 1441 698
rect 1446 672 1449 858
rect 1454 762 1457 948
rect 1462 922 1465 1148
rect 1474 1138 1478 1141
rect 1490 1118 1494 1121
rect 1470 992 1473 1028
rect 1486 942 1489 1108
rect 1534 1072 1537 1118
rect 1496 1003 1498 1007
rect 1502 1003 1505 1007
rect 1509 1003 1512 1007
rect 1506 948 1510 951
rect 1462 902 1465 918
rect 1470 912 1473 918
rect 1518 882 1521 1058
rect 1534 952 1537 1068
rect 1542 1062 1545 1158
rect 1646 1152 1649 1168
rect 1590 1148 1598 1151
rect 1550 1122 1553 1147
rect 1566 1142 1569 1148
rect 1578 1118 1582 1121
rect 1550 992 1553 1008
rect 1558 942 1561 1048
rect 1566 1032 1569 1058
rect 1574 1042 1577 1058
rect 1590 1052 1593 1148
rect 1622 1142 1625 1148
rect 1602 1138 1606 1141
rect 1614 1062 1617 1118
rect 1638 1072 1641 1098
rect 1646 1062 1649 1118
rect 1654 1112 1657 1258
rect 1662 1242 1665 1258
rect 1686 1242 1689 1258
rect 1670 1122 1673 1218
rect 1566 972 1569 1028
rect 1598 1012 1601 1058
rect 1574 952 1577 958
rect 1486 872 1489 878
rect 1506 868 1510 871
rect 1466 859 1470 862
rect 1496 803 1498 807
rect 1502 803 1505 807
rect 1509 803 1512 807
rect 1482 768 1486 771
rect 1518 752 1521 878
rect 1534 862 1537 868
rect 1558 852 1561 858
rect 1530 848 1534 851
rect 1566 802 1569 948
rect 1582 892 1585 948
rect 1590 912 1593 918
rect 1598 911 1601 928
rect 1598 908 1609 911
rect 1594 888 1598 891
rect 1582 872 1585 888
rect 1594 878 1598 881
rect 1606 862 1609 908
rect 1578 858 1582 861
rect 1614 852 1617 1058
rect 1622 1042 1625 1048
rect 1654 1042 1657 1048
rect 1670 1042 1673 1068
rect 1694 1061 1697 1308
rect 1734 1272 1737 1458
rect 1766 1352 1769 1358
rect 1742 1282 1745 1348
rect 1758 1342 1761 1348
rect 1750 1302 1753 1338
rect 1750 1272 1753 1288
rect 1782 1282 1785 1498
rect 1838 1491 1841 1738
rect 1862 1512 1865 1838
rect 1870 1702 1873 1718
rect 1870 1682 1873 1698
rect 1870 1652 1873 1658
rect 1894 1582 1897 1668
rect 1882 1548 1886 1551
rect 1894 1542 1897 1578
rect 1910 1542 1913 1938
rect 1918 1932 1921 1948
rect 1958 1942 1961 1948
rect 1974 1922 1977 1948
rect 1938 1918 1942 1921
rect 1998 1892 2001 1948
rect 2006 1942 2009 1948
rect 2014 1931 2017 2048
rect 2054 2042 2057 2148
rect 2086 2141 2089 2259
rect 2082 2138 2089 2141
rect 2094 2142 2097 2218
rect 2102 2182 2105 2268
rect 2134 2212 2137 2347
rect 2238 2342 2241 2348
rect 2334 2342 2337 2348
rect 2454 2342 2457 2358
rect 2494 2352 2497 2358
rect 2466 2348 2470 2351
rect 2218 2338 2222 2341
rect 2142 2252 2145 2338
rect 2462 2332 2465 2338
rect 2190 2262 2193 2278
rect 2154 2258 2158 2261
rect 2146 2218 2150 2221
rect 2158 2202 2161 2248
rect 2166 2222 2169 2258
rect 2158 2192 2161 2198
rect 2102 2142 2105 2178
rect 2174 2162 2177 2168
rect 2174 2152 2177 2158
rect 2086 2052 2089 2058
rect 2094 1972 2097 2068
rect 2118 2062 2121 2068
rect 2134 2062 2137 2068
rect 2006 1928 2017 1931
rect 2006 1892 2009 1928
rect 2034 1918 2038 1921
rect 2016 1903 2018 1907
rect 2022 1903 2025 1907
rect 2029 1903 2032 1907
rect 2030 1872 2033 1888
rect 2070 1872 2073 1878
rect 1958 1862 1961 1868
rect 1982 1862 1985 1868
rect 2078 1862 2081 1958
rect 2086 1952 2089 1958
rect 2094 1942 2097 1968
rect 2138 1958 2142 1961
rect 2138 1948 2145 1951
rect 2130 1938 2134 1941
rect 1998 1852 2001 1858
rect 1918 1752 1921 1838
rect 1990 1752 1993 1808
rect 1998 1792 2001 1838
rect 2006 1748 2014 1751
rect 2042 1748 2046 1751
rect 2062 1751 2065 1758
rect 2054 1748 2065 1751
rect 1918 1742 1921 1748
rect 1926 1702 1929 1748
rect 1982 1742 1985 1748
rect 1950 1692 1953 1698
rect 1926 1672 1929 1678
rect 1974 1672 1977 1718
rect 2006 1692 2009 1748
rect 2054 1742 2057 1748
rect 2066 1738 2070 1741
rect 2016 1703 2018 1707
rect 2022 1703 2025 1707
rect 2029 1703 2032 1707
rect 1978 1668 1993 1671
rect 1990 1662 1993 1668
rect 1930 1658 1934 1661
rect 1958 1652 1961 1658
rect 1982 1612 1985 1658
rect 1926 1542 1929 1558
rect 1942 1552 1945 1558
rect 1958 1552 1961 1558
rect 1830 1488 1841 1491
rect 1830 1472 1833 1488
rect 1794 1468 1798 1471
rect 1794 1458 1798 1461
rect 1850 1418 1854 1421
rect 1822 1352 1825 1358
rect 1838 1352 1841 1408
rect 1846 1362 1849 1368
rect 1794 1348 1798 1351
rect 1806 1322 1809 1348
rect 1830 1332 1833 1338
rect 1846 1312 1849 1318
rect 1862 1312 1865 1338
rect 1842 1288 1846 1291
rect 1702 1142 1705 1268
rect 1710 1232 1713 1258
rect 1726 1252 1729 1268
rect 1862 1262 1865 1288
rect 1782 1252 1785 1259
rect 1734 1232 1737 1248
rect 1782 1192 1785 1238
rect 1814 1222 1817 1258
rect 1854 1252 1857 1258
rect 1722 1168 1726 1171
rect 1718 1152 1721 1158
rect 1714 1138 1718 1141
rect 1706 1118 1710 1121
rect 1710 1082 1713 1098
rect 1690 1058 1697 1061
rect 1710 1052 1713 1068
rect 1726 1052 1729 1068
rect 1698 1048 1702 1051
rect 1702 1002 1705 1048
rect 1714 1028 1718 1031
rect 1734 992 1737 1168
rect 1746 1158 1750 1161
rect 1774 1152 1777 1158
rect 1758 1142 1761 1148
rect 1758 1122 1761 1138
rect 1742 1072 1745 1108
rect 1734 952 1737 958
rect 1646 892 1649 948
rect 1654 882 1657 888
rect 1654 872 1657 878
rect 1638 862 1641 868
rect 1630 812 1633 818
rect 1638 792 1641 828
rect 1578 768 1582 771
rect 1538 747 1542 750
rect 1590 742 1593 788
rect 1646 772 1649 858
rect 1662 772 1665 898
rect 1706 888 1710 891
rect 1682 868 1686 871
rect 1706 868 1713 871
rect 1670 852 1673 858
rect 1694 852 1697 868
rect 1710 862 1713 868
rect 1670 782 1673 848
rect 1702 782 1705 858
rect 1742 792 1745 1068
rect 1766 1022 1769 1148
rect 1814 1122 1817 1148
rect 1822 1142 1825 1148
rect 1822 1072 1825 1108
rect 1778 1048 1782 1051
rect 1814 1032 1817 1058
rect 1794 988 1798 991
rect 1754 948 1758 951
rect 1758 872 1761 948
rect 1798 922 1801 928
rect 1762 858 1766 861
rect 1654 752 1657 758
rect 1662 752 1665 768
rect 1694 762 1697 768
rect 1678 752 1681 758
rect 1610 748 1614 751
rect 1610 738 1614 741
rect 1446 662 1449 668
rect 1438 542 1441 548
rect 1446 462 1449 658
rect 1462 552 1465 608
rect 1454 532 1457 538
rect 1462 532 1465 538
rect 1462 392 1465 408
rect 1274 318 1278 321
rect 1166 242 1169 268
rect 1198 263 1201 278
rect 1318 272 1321 288
rect 1298 268 1302 271
rect 1138 168 1142 171
rect 1126 152 1129 158
rect 1194 148 1198 151
rect 1118 142 1121 148
rect 1222 142 1225 258
rect 1258 238 1262 241
rect 1262 192 1265 218
rect 1238 142 1241 148
rect 1130 138 1134 141
rect 1222 122 1225 138
rect 1246 132 1249 148
rect 1198 72 1201 108
rect 1206 82 1209 118
rect 1270 92 1273 268
rect 1278 262 1281 268
rect 1302 252 1305 258
rect 1286 172 1289 178
rect 1290 168 1294 171
rect 1278 132 1281 148
rect 1326 122 1329 138
rect 1266 68 1270 71
rect 970 59 974 62
rect 1038 62 1041 68
rect 1066 58 1070 61
rect 1062 52 1065 58
rect 1042 48 1046 51
rect 1110 32 1113 68
rect 1142 62 1145 68
rect 1158 62 1161 68
rect 1182 62 1185 68
rect 1286 62 1289 98
rect 1294 72 1297 88
rect 1326 82 1329 118
rect 1334 112 1337 268
rect 1350 263 1353 268
rect 1342 142 1345 148
rect 1366 142 1369 328
rect 1414 321 1417 338
rect 1422 331 1425 338
rect 1422 328 1430 331
rect 1414 318 1425 321
rect 1406 302 1409 318
rect 1422 292 1425 318
rect 1410 288 1414 291
rect 1422 252 1425 268
rect 1438 262 1441 388
rect 1470 362 1473 738
rect 1574 722 1577 738
rect 1518 672 1521 678
rect 1558 662 1561 668
rect 1486 612 1489 618
rect 1534 612 1537 648
rect 1496 603 1498 607
rect 1502 603 1505 607
rect 1509 603 1512 607
rect 1534 572 1537 608
rect 1590 582 1593 738
rect 1622 732 1625 748
rect 1654 732 1657 748
rect 1702 742 1705 778
rect 1742 751 1745 758
rect 1710 742 1713 748
rect 1666 738 1670 741
rect 1622 721 1625 728
rect 1614 718 1625 721
rect 1598 692 1601 698
rect 1614 642 1617 718
rect 1626 668 1630 671
rect 1654 662 1657 708
rect 1662 672 1665 738
rect 1670 672 1673 708
rect 1726 692 1729 738
rect 1774 722 1777 908
rect 1806 862 1809 868
rect 1682 678 1689 681
rect 1686 672 1689 678
rect 1722 678 1726 681
rect 1694 662 1697 678
rect 1702 662 1705 668
rect 1734 662 1737 668
rect 1646 652 1649 658
rect 1678 652 1681 658
rect 1626 648 1630 651
rect 1534 552 1537 568
rect 1558 562 1561 568
rect 1606 551 1609 558
rect 1494 542 1497 548
rect 1502 542 1505 548
rect 1526 542 1529 548
rect 1550 542 1553 548
rect 1494 492 1497 538
rect 1526 492 1529 518
rect 1518 462 1521 478
rect 1558 472 1561 498
rect 1542 462 1545 468
rect 1558 462 1561 468
rect 1550 422 1553 458
rect 1496 403 1498 407
rect 1502 403 1505 407
rect 1509 403 1512 407
rect 1486 352 1489 358
rect 1454 342 1457 348
rect 1382 142 1385 168
rect 1398 162 1401 248
rect 1438 242 1441 258
rect 1394 158 1398 161
rect 1434 158 1438 161
rect 1398 152 1401 158
rect 1402 138 1406 141
rect 1366 112 1369 138
rect 1390 92 1393 98
rect 1402 68 1406 71
rect 1334 62 1337 68
rect 1414 62 1417 158
rect 1426 148 1430 151
rect 1446 142 1449 268
rect 1454 262 1457 318
rect 1470 292 1473 338
rect 1478 312 1481 348
rect 1510 272 1513 318
rect 1462 262 1465 268
rect 1518 262 1521 298
rect 1534 292 1537 308
rect 1550 262 1553 268
rect 1558 262 1561 378
rect 1566 342 1569 488
rect 1574 482 1577 538
rect 1582 492 1585 518
rect 1590 492 1593 538
rect 1602 468 1606 471
rect 1574 452 1577 458
rect 1574 342 1577 347
rect 1462 162 1465 188
rect 1486 141 1489 258
rect 1496 203 1498 207
rect 1502 203 1505 207
rect 1509 203 1512 207
rect 1514 148 1518 151
rect 1482 138 1489 141
rect 1430 92 1433 138
rect 1442 118 1446 121
rect 1454 102 1457 138
rect 1430 72 1433 78
rect 1438 62 1441 68
rect 1262 52 1265 58
rect 1398 52 1401 58
rect 1414 52 1417 58
rect 1462 52 1465 118
rect 1478 92 1481 138
rect 1494 132 1497 138
rect 1526 102 1529 258
rect 1542 152 1545 228
rect 1566 202 1569 258
rect 1566 162 1569 198
rect 1566 152 1569 158
rect 1534 92 1537 148
rect 1550 142 1553 148
rect 1574 72 1577 328
rect 1590 292 1593 468
rect 1602 458 1606 461
rect 1614 392 1617 598
rect 1626 488 1630 491
rect 1670 482 1673 518
rect 1678 502 1681 518
rect 1686 492 1689 508
rect 1642 458 1646 461
rect 1682 458 1686 461
rect 1638 352 1641 458
rect 1702 452 1705 458
rect 1654 422 1657 438
rect 1654 352 1657 418
rect 1666 358 1670 361
rect 1614 302 1617 318
rect 1622 292 1625 338
rect 1586 288 1590 291
rect 1646 272 1649 288
rect 1590 262 1593 268
rect 1638 262 1641 268
rect 1662 262 1665 358
rect 1694 352 1697 428
rect 1710 392 1713 658
rect 1734 522 1737 548
rect 1742 542 1745 688
rect 1774 682 1777 718
rect 1790 662 1793 768
rect 1814 762 1817 998
rect 1830 952 1833 1218
rect 1870 1202 1873 1348
rect 1894 1342 1897 1348
rect 1886 1332 1889 1338
rect 1886 1302 1889 1328
rect 1894 1262 1897 1268
rect 1902 1262 1905 1508
rect 1910 1472 1913 1538
rect 1926 1462 1929 1478
rect 1950 1462 1953 1488
rect 1914 1458 1918 1461
rect 1958 1451 1961 1468
rect 1950 1448 1961 1451
rect 1934 1412 1937 1418
rect 1910 1352 1913 1368
rect 1910 1292 1913 1308
rect 1910 1272 1913 1278
rect 1926 1272 1929 1398
rect 1942 1352 1945 1378
rect 1934 1292 1937 1348
rect 1950 1342 1953 1448
rect 1958 1352 1961 1358
rect 1946 1338 1950 1341
rect 1838 1152 1841 1198
rect 1870 1162 1873 1168
rect 1858 1158 1862 1161
rect 1846 992 1849 1138
rect 1862 1052 1865 1118
rect 1878 1092 1881 1158
rect 1886 1142 1889 1258
rect 1902 1182 1905 1258
rect 1886 1091 1889 1138
rect 1894 1102 1897 1118
rect 1886 1088 1894 1091
rect 1878 1062 1881 1088
rect 1886 1022 1889 1068
rect 1878 962 1881 1018
rect 1862 942 1865 947
rect 1894 932 1897 938
rect 1838 862 1841 928
rect 1854 862 1857 918
rect 1886 862 1889 878
rect 1902 872 1905 1178
rect 1910 1172 1913 1258
rect 1910 1152 1913 1168
rect 1914 1138 1918 1141
rect 1910 962 1913 978
rect 1910 942 1913 948
rect 1898 858 1902 861
rect 1822 852 1825 858
rect 1830 752 1833 788
rect 1846 762 1849 858
rect 1862 852 1865 858
rect 1910 852 1913 858
rect 1878 762 1881 818
rect 1894 752 1897 838
rect 1842 748 1846 751
rect 1842 738 1849 741
rect 1806 722 1809 738
rect 1814 722 1817 728
rect 1838 692 1841 718
rect 1846 692 1849 738
rect 1854 702 1857 748
rect 1878 742 1881 748
rect 1886 742 1889 748
rect 1902 742 1905 748
rect 1910 712 1913 718
rect 1862 672 1865 688
rect 1890 678 1894 681
rect 1918 662 1921 868
rect 1926 852 1929 1268
rect 1950 1262 1953 1268
rect 1958 1172 1961 1348
rect 1958 1152 1961 1158
rect 1966 1151 1969 1548
rect 1982 1542 1985 1598
rect 2014 1592 2017 1658
rect 1990 1522 1993 1548
rect 2014 1542 2017 1558
rect 2022 1552 2025 1558
rect 2030 1522 2033 1558
rect 2016 1503 2018 1507
rect 2022 1503 2025 1507
rect 2029 1503 2032 1507
rect 1994 1468 1998 1471
rect 2026 1468 2030 1471
rect 2038 1462 2041 1738
rect 2078 1732 2081 1748
rect 2086 1742 2089 1938
rect 2118 1872 2121 1898
rect 2134 1872 2137 1918
rect 2118 1792 2121 1868
rect 2142 1832 2145 1948
rect 2150 1892 2153 1958
rect 2158 1942 2161 2138
rect 2182 1982 2185 2218
rect 2190 2122 2193 2138
rect 2190 2062 2193 2118
rect 2198 2102 2201 2318
rect 2206 2262 2209 2318
rect 2214 2282 2217 2318
rect 2254 2272 2257 2328
rect 2322 2318 2326 2321
rect 2410 2318 2414 2321
rect 2450 2318 2454 2321
rect 2218 2268 2222 2271
rect 2238 2262 2241 2268
rect 2246 2232 2249 2258
rect 2254 2222 2257 2268
rect 2286 2262 2289 2268
rect 2302 2262 2305 2268
rect 2390 2262 2393 2268
rect 2438 2262 2441 2268
rect 2362 2258 2366 2261
rect 2442 2258 2449 2261
rect 2262 2252 2265 2258
rect 2282 2248 2286 2251
rect 2214 2162 2217 2168
rect 2210 2148 2214 2151
rect 2238 2142 2241 2198
rect 2254 2151 2257 2158
rect 2218 2138 2222 2141
rect 2314 2118 2318 2121
rect 2326 2111 2329 2158
rect 2342 2152 2345 2188
rect 2350 2152 2353 2218
rect 2370 2158 2374 2161
rect 2318 2108 2329 2111
rect 2186 1958 2190 1961
rect 2166 1952 2169 1958
rect 2190 1942 2193 1948
rect 2198 1902 2201 2068
rect 2238 2062 2241 2068
rect 2254 2062 2257 2088
rect 2262 2062 2265 2098
rect 2318 2092 2321 2108
rect 2286 2062 2289 2088
rect 2326 2072 2329 2088
rect 2298 2068 2302 2071
rect 2334 2062 2337 2138
rect 2210 2058 2214 2061
rect 2222 2002 2225 2018
rect 2246 1992 2249 2058
rect 2342 2052 2345 2148
rect 2350 2142 2353 2148
rect 2358 2102 2361 2138
rect 2390 2082 2393 2258
rect 2410 2218 2414 2221
rect 2398 2192 2401 2208
rect 2398 2152 2401 2158
rect 2406 2142 2409 2148
rect 2410 2138 2414 2141
rect 2410 2118 2414 2121
rect 2406 2092 2409 2118
rect 2422 2082 2425 2218
rect 2446 2152 2449 2258
rect 2470 2252 2473 2259
rect 2486 2192 2489 2318
rect 2446 2082 2449 2118
rect 2422 2072 2425 2078
rect 2362 2058 2366 2061
rect 2314 2048 2318 2051
rect 2206 1942 2209 1968
rect 2154 1858 2158 1861
rect 2170 1858 2174 1861
rect 2150 1832 2153 1848
rect 2174 1812 2177 1818
rect 2198 1762 2201 1868
rect 2206 1862 2209 1938
rect 2214 1862 2217 1978
rect 2094 1722 2097 1748
rect 2102 1742 2105 1748
rect 2054 1692 2057 1718
rect 2066 1678 2070 1681
rect 2086 1672 2089 1708
rect 2110 1692 2113 1758
rect 2222 1752 2225 1958
rect 2246 1952 2249 1968
rect 2270 1962 2273 2018
rect 2266 1948 2270 1951
rect 2310 1942 2313 1978
rect 2430 1972 2433 2018
rect 2438 2012 2441 2048
rect 2330 1958 2334 1961
rect 2442 1958 2446 1961
rect 2454 1952 2457 2158
rect 2462 2082 2465 2088
rect 2470 2062 2473 2138
rect 2478 2111 2481 2147
rect 2478 2108 2489 2111
rect 2486 2092 2489 2108
rect 2494 2102 2497 2138
rect 2490 2078 2494 2081
rect 2470 2052 2473 2058
rect 2470 1952 2473 2028
rect 2386 1948 2390 1951
rect 2254 1872 2257 1938
rect 2294 1882 2297 1938
rect 2318 1912 2321 1948
rect 2334 1942 2337 1948
rect 2338 1918 2342 1921
rect 2334 1882 2337 1888
rect 2406 1872 2409 1928
rect 2286 1862 2289 1868
rect 2238 1812 2241 1858
rect 2246 1852 2249 1858
rect 2262 1852 2265 1858
rect 2282 1848 2286 1851
rect 2262 1802 2265 1848
rect 2302 1832 2305 1868
rect 2334 1863 2337 1868
rect 2394 1828 2398 1831
rect 2254 1752 2257 1758
rect 2302 1752 2305 1828
rect 2154 1748 2158 1751
rect 2214 1732 2217 1738
rect 2246 1732 2249 1748
rect 2262 1742 2265 1748
rect 2118 1712 2121 1718
rect 2146 1678 2150 1681
rect 2086 1662 2089 1668
rect 2118 1662 2121 1668
rect 2058 1658 2062 1661
rect 2046 1642 2049 1658
rect 2094 1652 2097 1658
rect 2158 1652 2161 1658
rect 2110 1642 2113 1648
rect 2046 1542 2049 1588
rect 2134 1582 2137 1648
rect 2166 1602 2169 1668
rect 2182 1662 2185 1728
rect 2270 1722 2273 1748
rect 2310 1742 2313 1808
rect 2282 1728 2286 1731
rect 2318 1692 2321 1748
rect 2214 1662 2217 1678
rect 2254 1662 2257 1668
rect 2174 1642 2177 1658
rect 2146 1588 2150 1591
rect 2070 1572 2073 1578
rect 2166 1572 2169 1598
rect 2058 1568 2062 1571
rect 2206 1552 2209 1558
rect 2278 1552 2281 1618
rect 2098 1548 2102 1551
rect 2134 1542 2137 1548
rect 2230 1542 2233 1548
rect 2318 1542 2321 1568
rect 2326 1562 2329 1818
rect 2406 1792 2409 1868
rect 2334 1672 2337 1788
rect 2374 1762 2377 1768
rect 2342 1752 2345 1758
rect 2350 1742 2353 1748
rect 2358 1692 2361 1738
rect 2366 1712 2369 1718
rect 2374 1702 2377 1758
rect 2386 1718 2390 1721
rect 2346 1688 2350 1691
rect 2374 1672 2377 1678
rect 2406 1663 2409 1678
rect 2422 1672 2425 1748
rect 2366 1572 2369 1618
rect 2346 1558 2350 1561
rect 2326 1552 2329 1558
rect 2250 1538 2254 1541
rect 2202 1488 2206 1491
rect 2282 1488 2286 1491
rect 2058 1478 2062 1481
rect 2086 1472 2089 1488
rect 2070 1462 2073 1468
rect 2138 1458 2142 1461
rect 1974 1452 1977 1458
rect 1994 1448 1998 1451
rect 1974 1392 1977 1448
rect 2014 1372 2017 1458
rect 2038 1432 2041 1458
rect 2046 1452 2049 1458
rect 2166 1452 2169 1468
rect 2190 1462 2193 1478
rect 2230 1472 2233 1488
rect 2282 1468 2286 1471
rect 2214 1462 2217 1468
rect 2230 1462 2233 1468
rect 2302 1462 2305 1518
rect 2318 1462 2321 1468
rect 2282 1458 2286 1461
rect 2222 1452 2225 1458
rect 2246 1452 2249 1458
rect 2274 1448 2278 1451
rect 1978 1358 1982 1361
rect 1982 1342 1985 1348
rect 2014 1342 2017 1368
rect 2016 1303 2018 1307
rect 2022 1303 2025 1307
rect 2029 1303 2032 1307
rect 2010 1288 2014 1291
rect 1974 1262 1977 1278
rect 1982 1212 1985 1258
rect 2022 1222 2025 1238
rect 2038 1212 2041 1428
rect 2074 1348 2078 1351
rect 2102 1342 2105 1358
rect 2118 1342 2121 1368
rect 2134 1362 2137 1408
rect 2158 1352 2161 1408
rect 2190 1372 2193 1448
rect 2170 1368 2174 1371
rect 2302 1362 2305 1458
rect 2302 1352 2305 1358
rect 2146 1348 2150 1351
rect 2226 1348 2230 1351
rect 2170 1338 2174 1341
rect 1962 1148 1969 1151
rect 1934 1132 1937 1148
rect 2038 1142 2041 1148
rect 2062 1142 2065 1308
rect 2070 1282 2073 1338
rect 2150 1292 2153 1338
rect 2254 1312 2257 1338
rect 2270 1302 2273 1318
rect 2102 1272 2105 1288
rect 2150 1272 2153 1288
rect 2070 1263 2073 1268
rect 2086 1172 2089 1268
rect 2118 1262 2121 1268
rect 2166 1262 2169 1298
rect 2178 1278 2182 1281
rect 2254 1272 2257 1288
rect 2258 1268 2262 1271
rect 2222 1262 2225 1268
rect 2246 1262 2249 1268
rect 2194 1258 2198 1261
rect 2142 1252 2145 1258
rect 2122 1248 2126 1251
rect 2158 1242 2161 1258
rect 2202 1248 2206 1251
rect 2246 1242 2249 1248
rect 2262 1242 2265 1258
rect 2318 1252 2321 1258
rect 2102 1142 2105 1168
rect 2198 1162 2201 1168
rect 2126 1152 2129 1158
rect 2202 1148 2206 1151
rect 1954 1138 1958 1141
rect 2194 1138 2198 1141
rect 1974 1112 1977 1128
rect 1994 1118 1998 1121
rect 1942 1062 1945 1098
rect 1974 1072 1977 1108
rect 2016 1103 2018 1107
rect 2022 1103 2025 1107
rect 2029 1103 2032 1107
rect 2006 1078 2025 1081
rect 2006 1071 2009 1078
rect 2022 1072 2025 1078
rect 2002 1068 2009 1071
rect 2014 1062 2017 1068
rect 2030 1062 2033 1088
rect 2094 1072 2097 1108
rect 2150 1082 2153 1138
rect 2182 1072 2185 1118
rect 2190 1112 2193 1138
rect 2214 1131 2217 1158
rect 2246 1152 2249 1198
rect 2254 1152 2257 1168
rect 2302 1152 2305 1208
rect 2310 1152 2313 1158
rect 2326 1152 2329 1548
rect 2350 1542 2353 1548
rect 2366 1542 2369 1568
rect 2342 1452 2345 1458
rect 2382 1432 2385 1468
rect 2390 1462 2393 1468
rect 2406 1462 2409 1468
rect 2402 1448 2406 1451
rect 2334 1342 2337 1347
rect 2342 1272 2345 1308
rect 2358 1272 2361 1298
rect 2366 1292 2369 1358
rect 2382 1352 2385 1358
rect 2374 1342 2377 1348
rect 2382 1271 2385 1348
rect 2374 1268 2385 1271
rect 2374 1252 2377 1268
rect 2382 1252 2385 1258
rect 2390 1252 2393 1268
rect 2350 1152 2353 1198
rect 2390 1192 2393 1248
rect 2398 1181 2401 1438
rect 2406 1392 2409 1428
rect 2422 1421 2425 1668
rect 2430 1542 2433 1548
rect 2438 1492 2441 1918
rect 2454 1822 2457 1948
rect 2462 1932 2465 1938
rect 2470 1882 2473 1948
rect 2466 1868 2470 1871
rect 2478 1822 2481 2068
rect 2486 1992 2489 2058
rect 2486 1982 2489 1988
rect 2502 1862 2505 1878
rect 2486 1781 2489 1818
rect 2486 1778 2497 1781
rect 2486 1762 2489 1768
rect 2446 1751 2449 1758
rect 2482 1748 2486 1751
rect 2478 1732 2481 1738
rect 2494 1732 2497 1778
rect 2502 1752 2505 1758
rect 2462 1671 2465 1708
rect 2470 1682 2473 1688
rect 2462 1668 2473 1671
rect 2446 1612 2449 1618
rect 2462 1582 2465 1658
rect 2470 1652 2473 1668
rect 2486 1662 2489 1698
rect 2494 1672 2497 1728
rect 2494 1572 2497 1668
rect 2482 1548 2486 1551
rect 2422 1418 2433 1421
rect 2414 1292 2417 1298
rect 2410 1278 2417 1281
rect 2406 1262 2409 1268
rect 2394 1178 2401 1181
rect 2382 1162 2385 1178
rect 2398 1162 2401 1168
rect 2338 1148 2342 1151
rect 2222 1142 2225 1148
rect 2214 1128 2225 1131
rect 2222 1092 2225 1128
rect 1994 1058 1998 1061
rect 1934 952 1937 978
rect 1942 872 1945 938
rect 1950 872 1953 918
rect 1958 892 1961 938
rect 1982 912 1985 948
rect 1966 852 1969 888
rect 1974 862 1977 868
rect 1926 752 1929 818
rect 1990 812 1993 848
rect 1934 742 1937 778
rect 1942 752 1945 808
rect 1950 762 1953 768
rect 1974 762 1977 808
rect 1998 751 2001 1058
rect 2006 1042 2009 1058
rect 2054 1032 2057 1058
rect 2078 1052 2081 1058
rect 2086 1042 2089 1058
rect 2094 1022 2097 1068
rect 2102 1062 2105 1068
rect 2118 1062 2121 1068
rect 2150 1063 2153 1068
rect 2238 1062 2241 1068
rect 2254 1062 2257 1068
rect 2046 952 2049 958
rect 2010 948 2014 951
rect 2016 903 2018 907
rect 2022 903 2025 907
rect 2029 903 2032 907
rect 2026 868 2030 871
rect 2018 848 2022 851
rect 2030 812 2033 858
rect 2010 788 2014 791
rect 2018 758 2022 761
rect 2038 752 2041 918
rect 2046 862 2049 888
rect 2054 881 2057 968
rect 2062 942 2065 958
rect 2078 952 2081 1008
rect 2102 1002 2105 1058
rect 2114 1048 2118 1051
rect 2110 992 2113 1028
rect 2102 952 2105 988
rect 2142 962 2145 998
rect 2150 992 2153 1048
rect 2198 1042 2201 1058
rect 2158 952 2161 1018
rect 2198 952 2201 1038
rect 2210 1018 2214 1021
rect 2130 948 2134 951
rect 2078 892 2081 948
rect 2086 912 2089 938
rect 2054 878 2065 881
rect 2046 752 2049 758
rect 1998 748 2009 751
rect 1934 692 1937 728
rect 1974 692 1977 748
rect 1990 722 1993 738
rect 1998 732 2001 738
rect 1926 672 1929 678
rect 1938 668 1942 671
rect 1990 662 1993 668
rect 2006 662 2009 748
rect 2018 738 2022 741
rect 2016 703 2018 707
rect 2022 703 2025 707
rect 2029 703 2032 707
rect 2022 672 2025 688
rect 2034 678 2038 681
rect 2046 672 2049 738
rect 2054 672 2057 868
rect 2062 742 2065 878
rect 2086 872 2089 908
rect 2094 842 2097 948
rect 2158 942 2161 948
rect 2126 872 2129 878
rect 2166 871 2169 918
rect 2206 892 2209 958
rect 2166 868 2174 871
rect 2194 868 2198 871
rect 2142 862 2145 868
rect 2174 862 2177 868
rect 2214 862 2217 1008
rect 2222 952 2225 1048
rect 2246 1042 2249 1058
rect 2262 1032 2265 1148
rect 2286 1142 2289 1148
rect 2270 1092 2273 1118
rect 2278 1062 2281 1068
rect 2270 1042 2273 1048
rect 2266 958 2270 961
rect 2286 952 2289 1088
rect 2294 1052 2297 1058
rect 2302 1012 2305 1148
rect 2318 1132 2321 1138
rect 2318 1062 2321 1068
rect 2310 1042 2313 1048
rect 2326 962 2329 1148
rect 2382 1142 2385 1158
rect 2414 1152 2417 1218
rect 2422 1202 2425 1348
rect 2430 1232 2433 1418
rect 2438 1392 2441 1468
rect 2446 1462 2449 1468
rect 2438 1312 2441 1318
rect 2454 1272 2457 1538
rect 2470 1292 2473 1528
rect 2478 1502 2481 1518
rect 2486 1322 2489 1538
rect 2502 1512 2505 1518
rect 2502 1482 2505 1488
rect 2494 1272 2497 1338
rect 2450 1258 2454 1261
rect 2430 1151 2433 1158
rect 2374 1132 2377 1138
rect 2414 1132 2417 1138
rect 2366 1092 2369 1118
rect 2374 1092 2377 1128
rect 2414 1092 2417 1108
rect 2438 1072 2441 1088
rect 2446 1072 2449 1078
rect 2390 1062 2393 1068
rect 2434 1058 2438 1061
rect 2306 948 2310 951
rect 2230 942 2233 947
rect 2262 942 2265 948
rect 2222 862 2225 918
rect 2262 872 2265 888
rect 2186 858 2190 861
rect 2102 852 2105 858
rect 2070 752 2073 758
rect 1874 658 1878 661
rect 1946 658 1950 661
rect 1842 648 1846 651
rect 1902 592 1905 658
rect 1910 652 1913 658
rect 1958 651 1961 658
rect 1950 648 1961 651
rect 1998 652 2001 658
rect 1950 592 1953 648
rect 1758 542 1761 578
rect 1822 542 1825 548
rect 1870 542 1873 548
rect 1886 542 1889 588
rect 2030 562 2033 668
rect 2046 561 2049 588
rect 2054 572 2057 658
rect 2062 592 2065 658
rect 2078 582 2081 748
rect 2086 722 2089 748
rect 2094 702 2097 718
rect 2094 662 2097 678
rect 2046 558 2057 561
rect 1894 552 1897 558
rect 2030 552 2033 558
rect 1986 548 1990 551
rect 1906 538 1910 541
rect 1758 492 1761 538
rect 1798 462 1801 478
rect 1806 472 1809 538
rect 1878 531 1881 538
rect 1918 532 1921 548
rect 1958 542 1961 548
rect 1874 528 1881 531
rect 1866 518 1870 521
rect 1902 492 1905 528
rect 1918 522 1921 528
rect 1926 492 1929 538
rect 1966 522 1969 548
rect 2014 542 2017 548
rect 1974 532 1977 538
rect 1966 512 1969 518
rect 1810 468 1814 471
rect 1958 462 1961 468
rect 1990 463 1993 468
rect 1794 458 1798 461
rect 1874 458 1878 461
rect 2006 462 2009 518
rect 2016 503 2018 507
rect 2022 503 2025 507
rect 2029 503 2032 507
rect 2038 482 2041 548
rect 2030 462 2033 468
rect 1670 342 1673 348
rect 1686 342 1689 348
rect 1670 322 1673 338
rect 1694 332 1697 348
rect 1702 342 1705 348
rect 1670 292 1673 298
rect 1670 282 1673 288
rect 1678 262 1681 318
rect 1694 272 1697 278
rect 1710 272 1713 318
rect 1718 292 1721 338
rect 1634 258 1638 261
rect 1650 258 1654 261
rect 1698 258 1702 261
rect 1614 252 1617 258
rect 1582 172 1585 218
rect 1594 178 1598 181
rect 1586 148 1590 151
rect 1598 142 1601 168
rect 1630 151 1633 178
rect 1598 82 1601 138
rect 1614 72 1617 138
rect 1638 72 1641 108
rect 1646 72 1649 168
rect 1470 62 1473 68
rect 1558 62 1561 68
rect 1574 62 1577 68
rect 1654 62 1657 238
rect 1694 142 1697 168
rect 1702 162 1705 208
rect 1710 142 1713 268
rect 1726 232 1729 418
rect 1742 352 1745 458
rect 1886 452 1889 458
rect 1782 422 1785 428
rect 1798 392 1801 448
rect 1862 392 1865 418
rect 1874 368 1878 371
rect 1770 348 1774 351
rect 1718 142 1721 188
rect 1726 182 1729 228
rect 1734 192 1737 348
rect 1774 342 1777 348
rect 1758 312 1761 318
rect 1782 292 1785 348
rect 1822 342 1825 368
rect 1866 358 1870 361
rect 1838 352 1841 358
rect 1858 348 1862 351
rect 1742 152 1745 208
rect 1754 188 1758 191
rect 1730 148 1734 151
rect 1746 138 1750 141
rect 1698 88 1702 91
rect 1678 72 1681 88
rect 1766 82 1769 268
rect 1774 262 1777 278
rect 1814 272 1817 288
rect 1830 252 1833 258
rect 1826 248 1830 251
rect 1838 222 1841 348
rect 1862 338 1870 341
rect 1862 322 1865 338
rect 1862 282 1865 318
rect 1874 288 1878 291
rect 1862 272 1865 278
rect 1850 258 1854 261
rect 1858 248 1862 251
rect 1902 221 1905 258
rect 1910 232 1913 458
rect 1918 352 1921 388
rect 1934 352 1937 358
rect 1894 218 1905 221
rect 1882 158 1886 161
rect 1862 152 1865 158
rect 1802 148 1806 151
rect 1838 142 1841 148
rect 1858 138 1862 141
rect 1854 91 1857 138
rect 1878 122 1881 128
rect 1846 88 1857 91
rect 1782 72 1785 78
rect 1814 72 1817 88
rect 1846 72 1849 88
rect 1894 82 1897 218
rect 1902 142 1905 168
rect 1918 152 1921 348
rect 1958 311 1961 458
rect 1990 392 1993 448
rect 1974 352 1977 378
rect 1950 308 1961 311
rect 1950 272 1953 308
rect 1966 262 1969 308
rect 1982 292 1985 348
rect 2006 291 2009 348
rect 2026 318 2030 321
rect 2016 303 2018 307
rect 2022 303 2025 307
rect 2029 303 2032 307
rect 2006 288 2017 291
rect 2002 258 2006 261
rect 1926 252 1929 258
rect 1918 142 1921 148
rect 1934 92 1937 258
rect 1974 252 1977 258
rect 1994 168 1998 171
rect 1942 132 1945 148
rect 2014 142 2017 288
rect 2038 261 2041 478
rect 2046 462 2049 508
rect 2054 492 2057 558
rect 2070 462 2073 488
rect 2078 472 2081 538
rect 2090 488 2094 491
rect 2078 442 2081 458
rect 2070 352 2073 388
rect 2046 292 2049 328
rect 2034 258 2041 261
rect 2054 272 2057 318
rect 2086 292 2089 348
rect 2102 272 2105 838
rect 2110 722 2113 778
rect 2118 742 2121 748
rect 2126 742 2129 798
rect 2142 762 2145 808
rect 2150 782 2153 858
rect 2202 848 2206 851
rect 2198 822 2201 848
rect 2166 762 2169 768
rect 2154 758 2158 761
rect 2194 758 2198 761
rect 2110 692 2113 718
rect 2126 702 2129 738
rect 2134 672 2137 718
rect 2122 668 2126 671
rect 2134 632 2137 658
rect 2142 631 2145 758
rect 2190 748 2198 751
rect 2150 742 2153 748
rect 2174 722 2177 738
rect 2158 692 2161 698
rect 2150 662 2153 668
rect 2150 642 2153 648
rect 2138 628 2145 631
rect 2138 548 2142 551
rect 2182 542 2185 548
rect 2150 512 2153 518
rect 2182 472 2185 488
rect 2118 462 2121 468
rect 2146 459 2150 462
rect 2134 362 2137 368
rect 2118 272 2121 278
rect 2122 268 2126 271
rect 2054 262 2057 268
rect 1938 88 1942 91
rect 1894 72 1897 78
rect 1950 72 1953 138
rect 2006 72 2009 128
rect 2038 112 2041 258
rect 2078 252 2081 268
rect 2102 262 2105 268
rect 2134 261 2137 358
rect 2170 348 2174 351
rect 2178 348 2185 351
rect 2150 342 2153 348
rect 2158 342 2161 348
rect 2130 258 2137 261
rect 2046 152 2049 218
rect 2062 152 2065 178
rect 2094 152 2097 258
rect 2142 252 2145 318
rect 2182 292 2185 348
rect 2190 342 2193 748
rect 2198 732 2201 738
rect 2206 692 2209 738
rect 2206 662 2209 668
rect 2214 602 2217 858
rect 2278 852 2281 858
rect 2286 852 2289 948
rect 2318 942 2321 958
rect 2326 952 2329 958
rect 2358 942 2361 1058
rect 2406 1052 2409 1058
rect 2374 951 2377 958
rect 2294 912 2297 938
rect 2342 922 2345 938
rect 2302 862 2305 898
rect 2310 872 2313 908
rect 2326 872 2329 878
rect 2302 842 2305 848
rect 2326 841 2329 868
rect 2342 852 2345 859
rect 2318 838 2329 841
rect 2238 752 2241 818
rect 2246 752 2249 828
rect 2254 752 2257 768
rect 2294 742 2297 748
rect 2238 672 2241 678
rect 2254 672 2257 678
rect 2262 662 2265 688
rect 2286 678 2294 681
rect 2286 662 2289 678
rect 2302 672 2305 778
rect 2318 732 2321 838
rect 2358 741 2361 938
rect 2406 902 2409 1048
rect 2446 962 2449 1058
rect 2442 958 2446 961
rect 2402 888 2406 891
rect 2414 872 2417 878
rect 2354 738 2361 741
rect 2422 862 2425 958
rect 2434 918 2438 921
rect 2434 858 2438 861
rect 2422 742 2425 858
rect 2446 851 2449 918
rect 2454 892 2457 1228
rect 2490 1178 2494 1181
rect 2498 1088 2502 1091
rect 2486 992 2489 1028
rect 2510 952 2513 2338
rect 2518 1562 2521 2008
rect 2466 948 2470 951
rect 2478 942 2481 948
rect 2466 938 2470 941
rect 2510 892 2513 948
rect 2442 848 2449 851
rect 2470 752 2473 878
rect 2506 868 2510 871
rect 2482 758 2486 761
rect 2518 752 2521 1558
rect 2442 748 2446 751
rect 2462 742 2465 748
rect 2470 742 2473 748
rect 2498 738 2502 741
rect 2318 682 2321 728
rect 2330 688 2334 691
rect 2358 672 2361 678
rect 2214 542 2217 547
rect 2262 542 2265 618
rect 2278 592 2281 598
rect 2286 592 2289 658
rect 2294 652 2297 658
rect 2270 542 2273 548
rect 2250 538 2254 541
rect 2238 482 2241 508
rect 2246 492 2249 528
rect 2198 462 2201 468
rect 2198 442 2201 448
rect 2154 268 2158 271
rect 2170 258 2174 261
rect 2150 252 2153 258
rect 2118 192 2121 228
rect 2102 152 2105 158
rect 2134 152 2137 158
rect 2182 152 2185 158
rect 2154 148 2158 151
rect 2054 132 2057 148
rect 2074 138 2078 141
rect 2016 103 2018 107
rect 2022 103 2025 107
rect 2029 103 2032 107
rect 2054 102 2057 128
rect 2094 92 2097 148
rect 2110 132 2113 148
rect 2198 142 2201 348
rect 2206 342 2209 478
rect 2230 472 2233 478
rect 2262 471 2265 538
rect 2270 482 2273 538
rect 2278 492 2281 568
rect 2254 468 2265 471
rect 2254 462 2257 468
rect 2222 442 2225 458
rect 2262 452 2265 458
rect 2238 362 2241 368
rect 2214 352 2217 358
rect 2270 342 2273 458
rect 2230 272 2233 318
rect 2262 292 2265 338
rect 2278 272 2281 468
rect 2286 292 2289 578
rect 2294 381 2297 648
rect 2302 602 2305 668
rect 2390 663 2393 678
rect 2406 672 2409 718
rect 2422 692 2425 728
rect 2454 682 2457 718
rect 2454 662 2457 668
rect 2310 562 2313 618
rect 2318 612 2321 648
rect 2462 622 2465 738
rect 2314 548 2318 551
rect 2294 378 2305 381
rect 2294 352 2297 368
rect 2302 352 2305 378
rect 2310 332 2313 458
rect 2326 352 2329 568
rect 2374 562 2377 568
rect 2390 552 2393 608
rect 2402 588 2406 591
rect 2478 591 2481 718
rect 2510 692 2513 698
rect 2470 588 2481 591
rect 2338 548 2342 551
rect 2378 548 2382 551
rect 2470 551 2473 588
rect 2402 538 2406 541
rect 2342 471 2345 518
rect 2358 472 2361 538
rect 2406 472 2409 488
rect 2342 468 2353 471
rect 2350 462 2353 468
rect 2386 468 2390 471
rect 2338 458 2342 461
rect 2358 352 2361 468
rect 2370 458 2374 461
rect 2390 452 2393 458
rect 2422 421 2425 468
rect 2438 463 2441 468
rect 2422 418 2433 421
rect 2402 358 2406 361
rect 2374 352 2377 358
rect 2326 342 2329 348
rect 2398 342 2401 348
rect 2346 338 2350 341
rect 2310 292 2313 328
rect 2298 288 2302 291
rect 2342 262 2345 318
rect 2366 272 2369 338
rect 2394 288 2398 291
rect 2358 262 2361 268
rect 2214 152 2217 198
rect 2146 138 2150 141
rect 2210 138 2214 141
rect 2110 92 2113 98
rect 2062 72 2065 78
rect 2158 72 2161 78
rect 1978 68 1982 71
rect 1670 62 1673 68
rect 1758 62 1761 68
rect 1530 58 1534 61
rect 1694 52 1697 58
rect 1806 52 1809 68
rect 1838 62 1841 68
rect 2046 63 2049 68
rect 1878 52 1881 59
rect 2166 62 2169 138
rect 2198 91 2201 138
rect 2198 88 2206 91
rect 2214 72 2217 138
rect 2222 82 2225 258
rect 2238 252 2241 258
rect 2294 242 2297 248
rect 2238 162 2241 198
rect 2366 192 2369 268
rect 2254 162 2257 168
rect 2406 162 2409 358
rect 2414 342 2417 368
rect 2430 342 2433 418
rect 2446 351 2449 358
rect 2430 332 2433 338
rect 2462 282 2465 538
rect 2498 488 2502 491
rect 2518 442 2521 748
rect 2506 368 2510 371
rect 2494 272 2497 278
rect 2502 262 2505 298
rect 2450 258 2454 261
rect 2438 192 2441 258
rect 2510 192 2513 358
rect 2518 302 2521 438
rect 2518 282 2521 288
rect 2518 252 2521 258
rect 2498 158 2502 161
rect 2238 142 2241 148
rect 2254 142 2257 158
rect 2314 148 2318 151
rect 2342 142 2345 148
rect 2358 142 2361 148
rect 2518 142 2521 238
rect 2426 138 2430 141
rect 2490 138 2494 141
rect 2270 92 2273 128
rect 2350 72 2353 78
rect 2366 72 2369 138
rect 2422 72 2425 138
rect 2442 88 2446 91
rect 2482 88 2486 91
rect 2518 72 2521 78
rect 2242 68 2246 71
rect 2434 68 2438 71
rect 2326 62 2329 68
rect 2218 58 2222 61
rect 1802 48 1806 51
rect 1838 42 1841 48
rect 1958 32 1961 58
rect 2246 52 2249 58
rect 2478 52 2481 68
rect 1982 32 1985 48
rect 878 -22 889 -19
rect 1422 -18 1425 8
rect 1496 3 1498 7
rect 1502 3 1505 7
rect 1509 3 1512 7
rect 1654 -18 1657 8
rect 2038 -18 2041 8
rect 1422 -22 1426 -18
rect 1654 -22 1658 -18
rect 2038 -22 2042 -18
<< m3contact >>
rect 246 2398 250 2402
rect 262 2398 266 2402
rect 70 2358 74 2362
rect 86 2358 90 2362
rect 94 2348 98 2352
rect 22 2338 26 2342
rect 54 2338 58 2342
rect 62 2328 66 2332
rect 14 2218 18 2222
rect 166 2348 170 2352
rect 294 2358 298 2362
rect 310 2358 314 2362
rect 366 2358 370 2362
rect 286 2348 290 2352
rect 318 2348 322 2352
rect 278 2338 282 2342
rect 454 2338 458 2342
rect 174 2328 178 2332
rect 110 2268 114 2272
rect 190 2258 194 2262
rect 206 2258 210 2262
rect 198 2248 202 2252
rect 86 2238 90 2242
rect 166 2238 170 2242
rect 134 2228 138 2232
rect 70 2208 74 2212
rect 14 2188 18 2192
rect 86 2168 90 2172
rect 110 2168 114 2172
rect 70 2158 74 2162
rect 190 2208 194 2212
rect 150 2188 154 2192
rect 142 2168 146 2172
rect 118 2158 122 2162
rect 102 2148 106 2152
rect 134 2148 138 2152
rect 102 2108 106 2112
rect 14 2088 18 2092
rect 86 2078 90 2082
rect 62 2058 66 2062
rect 126 2058 130 2062
rect 110 2048 114 2052
rect 134 2038 138 2042
rect 62 1968 66 1972
rect 102 1968 106 1972
rect 14 1868 18 1872
rect 86 1948 90 1952
rect 166 2168 170 2172
rect 158 2108 162 2112
rect 150 2078 154 2082
rect 206 2148 210 2152
rect 222 2328 226 2332
rect 286 2328 290 2332
rect 366 2328 370 2332
rect 334 2318 338 2322
rect 222 2288 226 2292
rect 254 2248 258 2252
rect 254 2218 258 2222
rect 214 2128 218 2132
rect 206 2118 210 2122
rect 238 2118 242 2122
rect 246 2098 250 2102
rect 222 2068 226 2072
rect 174 2058 178 2062
rect 190 2058 194 2062
rect 190 1988 194 1992
rect 126 1938 130 1942
rect 214 1918 218 1922
rect 110 1868 114 1872
rect 206 1868 210 1872
rect 222 1868 226 1872
rect 78 1858 82 1862
rect 94 1858 98 1862
rect 118 1858 122 1862
rect 142 1858 146 1862
rect 190 1858 194 1862
rect 30 1848 34 1852
rect 46 1848 50 1852
rect 14 1778 18 1782
rect 134 1838 138 1842
rect 158 1838 162 1842
rect 94 1798 98 1802
rect 150 1778 154 1782
rect 86 1768 90 1772
rect 70 1758 74 1762
rect 142 1758 146 1762
rect 118 1748 122 1752
rect 174 1768 178 1772
rect 182 1758 186 1762
rect 182 1748 186 1752
rect 102 1738 106 1742
rect 142 1738 146 1742
rect 126 1728 130 1732
rect 118 1688 122 1692
rect 182 1728 186 1732
rect 150 1668 154 1672
rect 118 1658 122 1662
rect 46 1648 50 1652
rect 54 1548 58 1552
rect 110 1558 114 1562
rect 142 1558 146 1562
rect 126 1548 130 1552
rect 310 2288 314 2292
rect 334 2288 338 2292
rect 358 2268 362 2272
rect 286 2238 290 2242
rect 350 2248 354 2252
rect 422 2318 426 2322
rect 422 2288 426 2292
rect 406 2258 410 2262
rect 382 2248 386 2252
rect 414 2248 418 2252
rect 374 2238 378 2242
rect 326 2218 330 2222
rect 350 2168 354 2172
rect 286 2158 290 2162
rect 318 2158 322 2162
rect 278 2088 282 2092
rect 302 2138 306 2142
rect 454 2248 458 2252
rect 482 2403 486 2407
rect 489 2403 493 2407
rect 1498 2403 1502 2407
rect 1505 2403 1509 2407
rect 918 2398 922 2402
rect 1142 2398 1146 2402
rect 1158 2398 1162 2402
rect 742 2378 746 2382
rect 854 2378 858 2382
rect 1126 2378 1130 2382
rect 558 2368 562 2372
rect 574 2368 578 2372
rect 638 2368 642 2372
rect 558 2358 562 2362
rect 590 2358 594 2362
rect 510 2348 514 2352
rect 558 2348 562 2352
rect 598 2348 602 2352
rect 1046 2368 1050 2372
rect 1110 2368 1114 2372
rect 1102 2358 1106 2362
rect 1126 2358 1130 2362
rect 718 2348 722 2352
rect 750 2348 754 2352
rect 558 2338 562 2342
rect 582 2338 586 2342
rect 758 2338 762 2342
rect 766 2338 770 2342
rect 534 2328 538 2332
rect 510 2288 514 2292
rect 550 2288 554 2292
rect 566 2268 570 2272
rect 630 2328 634 2332
rect 622 2268 626 2272
rect 646 2318 650 2322
rect 702 2318 706 2322
rect 758 2308 762 2312
rect 678 2278 682 2282
rect 758 2278 762 2282
rect 630 2258 634 2262
rect 482 2203 486 2207
rect 489 2203 493 2207
rect 358 2158 362 2162
rect 438 2158 442 2162
rect 342 2138 346 2142
rect 326 2118 330 2122
rect 278 2068 282 2072
rect 294 2068 298 2072
rect 278 2058 282 2062
rect 270 1988 274 1992
rect 270 1968 274 1972
rect 238 1858 242 1862
rect 286 1948 290 1952
rect 326 2048 330 2052
rect 358 2078 362 2082
rect 374 2058 378 2062
rect 390 2048 394 2052
rect 342 2018 346 2022
rect 318 1958 322 1962
rect 350 1958 354 1962
rect 310 1948 314 1952
rect 294 1868 298 1872
rect 262 1808 266 1812
rect 254 1788 258 1792
rect 246 1778 250 1782
rect 246 1768 250 1772
rect 230 1758 234 1762
rect 214 1748 218 1752
rect 270 1758 274 1762
rect 222 1738 226 1742
rect 262 1738 266 1742
rect 238 1708 242 1712
rect 206 1688 210 1692
rect 230 1688 234 1692
rect 190 1668 194 1672
rect 198 1658 202 1662
rect 190 1628 194 1632
rect 246 1678 250 1682
rect 254 1668 258 1672
rect 294 1848 298 1852
rect 302 1788 306 1792
rect 318 1928 322 1932
rect 342 1888 346 1892
rect 334 1868 338 1872
rect 334 1858 338 1862
rect 318 1848 322 1852
rect 310 1768 314 1772
rect 326 1758 330 1762
rect 294 1748 298 1752
rect 366 1738 370 1742
rect 350 1728 354 1732
rect 302 1678 306 1682
rect 406 2138 410 2142
rect 438 2128 442 2132
rect 526 2128 530 2132
rect 414 2118 418 2122
rect 406 2108 410 2112
rect 406 2048 410 2052
rect 406 1968 410 1972
rect 430 1938 434 1942
rect 406 1888 410 1892
rect 390 1868 394 1872
rect 598 2248 602 2252
rect 590 2238 594 2242
rect 638 2218 642 2222
rect 742 2258 746 2262
rect 670 2208 674 2212
rect 686 2208 690 2212
rect 614 2198 618 2202
rect 638 2198 642 2202
rect 662 2198 666 2202
rect 622 2158 626 2162
rect 542 2108 546 2112
rect 582 2098 586 2102
rect 542 2088 546 2092
rect 574 2088 578 2092
rect 494 2058 498 2062
rect 510 2058 514 2062
rect 446 2048 450 2052
rect 482 2003 486 2007
rect 489 2003 493 2007
rect 446 1988 450 1992
rect 502 1978 506 1982
rect 462 1968 466 1972
rect 510 1958 514 1962
rect 526 1958 530 1962
rect 454 1938 458 1942
rect 622 2068 626 2072
rect 590 2058 594 2062
rect 606 2058 610 2062
rect 630 2058 634 2062
rect 590 2048 594 2052
rect 558 2038 562 2042
rect 558 1978 562 1982
rect 550 1958 554 1962
rect 582 1948 586 1952
rect 630 2038 634 2042
rect 606 2008 610 2012
rect 622 1948 626 1952
rect 654 2168 658 2172
rect 646 2158 650 2162
rect 702 2178 706 2182
rect 694 2158 698 2162
rect 806 2308 810 2312
rect 790 2268 794 2272
rect 838 2328 842 2332
rect 854 2308 858 2312
rect 822 2298 826 2302
rect 870 2288 874 2292
rect 1806 2398 1810 2402
rect 1918 2368 1922 2372
rect 1214 2358 1218 2362
rect 910 2338 914 2342
rect 974 2338 978 2342
rect 1102 2338 1106 2342
rect 1198 2338 1202 2342
rect 854 2278 858 2282
rect 902 2278 906 2282
rect 1006 2328 1010 2332
rect 918 2318 922 2322
rect 910 2268 914 2272
rect 814 2258 818 2262
rect 702 2148 706 2152
rect 726 2148 730 2152
rect 766 2148 770 2152
rect 662 2108 666 2112
rect 654 2078 658 2082
rect 646 2018 650 2022
rect 654 1958 658 1962
rect 518 1938 522 1942
rect 606 1938 610 1942
rect 646 1938 650 1942
rect 470 1888 474 1892
rect 486 1888 490 1892
rect 542 1888 546 1892
rect 614 1928 618 1932
rect 438 1878 442 1882
rect 510 1878 514 1882
rect 558 1878 562 1882
rect 454 1868 458 1872
rect 430 1858 434 1862
rect 438 1848 442 1852
rect 606 1868 610 1872
rect 422 1818 426 1822
rect 446 1818 450 1822
rect 446 1798 450 1802
rect 398 1758 402 1762
rect 374 1708 378 1712
rect 350 1688 354 1692
rect 438 1738 442 1742
rect 358 1678 362 1682
rect 414 1678 418 1682
rect 318 1668 322 1672
rect 334 1668 338 1672
rect 390 1668 394 1672
rect 406 1668 410 1672
rect 318 1648 322 1652
rect 342 1648 346 1652
rect 278 1588 282 1592
rect 198 1558 202 1562
rect 166 1548 170 1552
rect 182 1548 186 1552
rect 206 1548 210 1552
rect 222 1548 226 1552
rect 238 1548 242 1552
rect 110 1538 114 1542
rect 158 1538 162 1542
rect 222 1528 226 1532
rect 174 1518 178 1522
rect 38 1468 42 1472
rect 126 1468 130 1472
rect 142 1468 146 1472
rect 118 1458 122 1462
rect 150 1458 154 1462
rect 206 1458 210 1462
rect 54 1438 58 1442
rect 166 1438 170 1442
rect 38 1388 42 1392
rect 6 1348 10 1352
rect 214 1428 218 1432
rect 102 1398 106 1402
rect 150 1378 154 1382
rect 174 1378 178 1382
rect 230 1398 234 1402
rect 86 1348 90 1352
rect 166 1348 170 1352
rect 198 1348 202 1352
rect 150 1338 154 1342
rect 158 1338 162 1342
rect 134 1328 138 1332
rect 142 1318 146 1322
rect 94 1278 98 1282
rect 118 1278 122 1282
rect 54 1268 58 1272
rect 190 1328 194 1332
rect 214 1328 218 1332
rect 190 1288 194 1292
rect 174 1268 178 1272
rect 126 1258 130 1262
rect 110 1248 114 1252
rect 142 1248 146 1252
rect 102 1238 106 1242
rect 174 1258 178 1262
rect 182 1258 186 1262
rect 262 1538 266 1542
rect 302 1528 306 1532
rect 254 1468 258 1472
rect 278 1458 282 1462
rect 262 1438 266 1442
rect 286 1438 290 1442
rect 254 1418 258 1422
rect 246 1358 250 1362
rect 310 1448 314 1452
rect 302 1418 306 1422
rect 270 1388 274 1392
rect 270 1358 274 1362
rect 262 1338 266 1342
rect 286 1338 290 1342
rect 254 1328 258 1332
rect 278 1328 282 1332
rect 374 1638 378 1642
rect 366 1628 370 1632
rect 390 1618 394 1622
rect 430 1648 434 1652
rect 534 1848 538 1852
rect 574 1848 578 1852
rect 534 1838 538 1842
rect 482 1803 486 1807
rect 489 1803 493 1807
rect 574 1828 578 1832
rect 518 1788 522 1792
rect 486 1778 490 1782
rect 510 1758 514 1762
rect 470 1748 474 1752
rect 526 1768 530 1772
rect 526 1748 530 1752
rect 542 1748 546 1752
rect 630 1878 634 1882
rect 654 1878 658 1882
rect 670 2058 674 2062
rect 694 2058 698 2062
rect 718 2138 722 2142
rect 862 2258 866 2262
rect 878 2258 882 2262
rect 862 2248 866 2252
rect 870 2228 874 2232
rect 894 2218 898 2222
rect 870 2198 874 2202
rect 846 2158 850 2162
rect 774 2138 778 2142
rect 750 2128 754 2132
rect 742 2118 746 2122
rect 758 2118 762 2122
rect 726 2108 730 2112
rect 766 2108 770 2112
rect 790 2108 794 2112
rect 750 2078 754 2082
rect 774 2078 778 2082
rect 734 2058 738 2062
rect 718 2048 722 2052
rect 702 2018 706 2022
rect 886 2078 890 2082
rect 766 1998 770 2002
rect 742 1988 746 1992
rect 678 1968 682 1972
rect 686 1958 690 1962
rect 710 1958 714 1962
rect 702 1948 706 1952
rect 686 1938 690 1942
rect 678 1918 682 1922
rect 670 1868 674 1872
rect 678 1868 682 1872
rect 798 2038 802 2042
rect 822 2038 826 2042
rect 1086 2308 1090 2312
rect 986 2303 990 2307
rect 993 2303 997 2307
rect 1174 2328 1178 2332
rect 1190 2318 1194 2322
rect 1094 2288 1098 2292
rect 942 2278 946 2282
rect 974 2278 978 2282
rect 1102 2278 1106 2282
rect 1006 2268 1010 2272
rect 1030 2268 1034 2272
rect 1054 2268 1058 2272
rect 1078 2268 1082 2272
rect 958 2258 962 2262
rect 1014 2258 1018 2262
rect 910 2198 914 2202
rect 918 2168 922 2172
rect 902 2148 906 2152
rect 910 2148 914 2152
rect 926 2148 930 2152
rect 910 2138 914 2142
rect 910 2118 914 2122
rect 902 2078 906 2082
rect 894 2038 898 2042
rect 806 1948 810 1952
rect 966 2188 970 2192
rect 998 2178 1002 2182
rect 1038 2208 1042 2212
rect 958 2148 962 2152
rect 942 2118 946 2122
rect 990 2118 994 2122
rect 986 2103 990 2107
rect 993 2103 997 2107
rect 974 2078 978 2082
rect 1006 2078 1010 2082
rect 1086 2258 1090 2262
rect 1078 2248 1082 2252
rect 1110 2248 1114 2252
rect 1070 2238 1074 2242
rect 1126 2238 1130 2242
rect 1062 2178 1066 2182
rect 1054 2148 1058 2152
rect 1030 2098 1034 2102
rect 1030 2078 1034 2082
rect 1062 2138 1066 2142
rect 1086 2138 1090 2142
rect 1078 2128 1082 2132
rect 1078 2098 1082 2102
rect 1286 2358 1290 2362
rect 1302 2358 1306 2362
rect 1326 2358 1330 2362
rect 1342 2358 1346 2362
rect 1278 2348 1282 2352
rect 1478 2348 1482 2352
rect 1510 2348 1514 2352
rect 1574 2348 1578 2352
rect 1598 2348 1602 2352
rect 1286 2338 1290 2342
rect 1246 2328 1250 2332
rect 1230 2308 1234 2312
rect 1150 2288 1154 2292
rect 1206 2288 1210 2292
rect 1182 2258 1186 2262
rect 1198 2258 1202 2262
rect 1166 2238 1170 2242
rect 1158 2218 1162 2222
rect 1206 2228 1210 2232
rect 1166 2208 1170 2212
rect 1214 2218 1218 2222
rect 1222 2148 1226 2152
rect 1190 2138 1194 2142
rect 1150 2128 1154 2132
rect 1182 2128 1186 2132
rect 1134 2108 1138 2112
rect 1174 2108 1178 2112
rect 1158 2078 1162 2082
rect 1014 2058 1018 2062
rect 1022 2058 1026 2062
rect 1046 2058 1050 2062
rect 982 2048 986 2052
rect 950 2028 954 2032
rect 958 1958 962 1962
rect 966 1958 970 1962
rect 1014 1958 1018 1962
rect 958 1948 962 1952
rect 726 1938 730 1942
rect 774 1938 778 1942
rect 798 1938 802 1942
rect 806 1898 810 1902
rect 718 1888 722 1892
rect 894 1928 898 1932
rect 934 1918 938 1922
rect 1006 1948 1010 1952
rect 966 1928 970 1932
rect 986 1903 990 1907
rect 993 1903 997 1907
rect 902 1898 906 1902
rect 958 1898 962 1902
rect 878 1888 882 1892
rect 814 1878 818 1882
rect 926 1888 930 1892
rect 910 1878 914 1882
rect 958 1878 962 1882
rect 734 1868 738 1872
rect 846 1868 850 1872
rect 862 1868 866 1872
rect 966 1868 970 1872
rect 998 1868 1002 1872
rect 638 1848 642 1852
rect 670 1848 674 1852
rect 718 1848 722 1852
rect 622 1838 626 1842
rect 662 1838 666 1842
rect 694 1828 698 1832
rect 590 1788 594 1792
rect 590 1778 594 1782
rect 638 1778 642 1782
rect 542 1728 546 1732
rect 566 1728 570 1732
rect 526 1698 530 1702
rect 454 1688 458 1692
rect 454 1668 458 1672
rect 494 1668 498 1672
rect 518 1668 522 1672
rect 446 1648 450 1652
rect 470 1648 474 1652
rect 438 1638 442 1642
rect 446 1638 450 1642
rect 462 1638 466 1642
rect 398 1608 402 1612
rect 510 1638 514 1642
rect 478 1618 482 1622
rect 482 1603 486 1607
rect 489 1603 493 1607
rect 454 1568 458 1572
rect 358 1548 362 1552
rect 366 1548 370 1552
rect 478 1548 482 1552
rect 486 1548 490 1552
rect 342 1528 346 1532
rect 326 1488 330 1492
rect 326 1478 330 1482
rect 350 1508 354 1512
rect 422 1538 426 1542
rect 462 1538 466 1542
rect 358 1488 362 1492
rect 342 1468 346 1472
rect 358 1468 362 1472
rect 326 1458 330 1462
rect 342 1458 346 1462
rect 374 1498 378 1502
rect 374 1488 378 1492
rect 374 1478 378 1482
rect 374 1468 378 1472
rect 382 1468 386 1472
rect 374 1418 378 1422
rect 366 1408 370 1412
rect 422 1518 426 1522
rect 414 1488 418 1492
rect 406 1478 410 1482
rect 518 1628 522 1632
rect 558 1688 562 1692
rect 566 1648 570 1652
rect 630 1768 634 1772
rect 702 1758 706 1762
rect 726 1758 730 1762
rect 638 1748 642 1752
rect 606 1718 610 1722
rect 630 1718 634 1722
rect 630 1688 634 1692
rect 686 1718 690 1722
rect 678 1688 682 1692
rect 638 1678 642 1682
rect 702 1698 706 1702
rect 734 1688 738 1692
rect 806 1858 810 1862
rect 878 1858 882 1862
rect 878 1848 882 1852
rect 894 1848 898 1852
rect 798 1828 802 1832
rect 782 1738 786 1742
rect 774 1728 778 1732
rect 758 1678 762 1682
rect 782 1678 786 1682
rect 646 1658 650 1662
rect 662 1658 666 1662
rect 702 1658 706 1662
rect 710 1658 714 1662
rect 742 1658 746 1662
rect 582 1638 586 1642
rect 638 1638 642 1642
rect 518 1618 522 1622
rect 542 1618 546 1622
rect 662 1608 666 1612
rect 718 1598 722 1602
rect 686 1578 690 1582
rect 526 1568 530 1572
rect 598 1568 602 1572
rect 662 1568 666 1572
rect 654 1558 658 1562
rect 670 1558 674 1562
rect 678 1558 682 1562
rect 542 1538 546 1542
rect 470 1508 474 1512
rect 502 1488 506 1492
rect 486 1478 490 1482
rect 430 1468 434 1472
rect 446 1468 450 1472
rect 438 1458 442 1462
rect 446 1448 450 1452
rect 478 1458 482 1462
rect 470 1448 474 1452
rect 630 1548 634 1552
rect 566 1528 570 1532
rect 558 1508 562 1512
rect 686 1538 690 1542
rect 686 1528 690 1532
rect 526 1488 530 1492
rect 550 1488 554 1492
rect 670 1488 674 1492
rect 542 1478 546 1482
rect 582 1478 586 1482
rect 566 1468 570 1472
rect 694 1468 698 1472
rect 518 1458 522 1462
rect 678 1448 682 1452
rect 430 1408 434 1412
rect 510 1408 514 1412
rect 482 1403 486 1407
rect 489 1403 493 1407
rect 518 1398 522 1402
rect 454 1388 458 1392
rect 486 1368 490 1372
rect 414 1348 418 1352
rect 430 1348 434 1352
rect 470 1348 474 1352
rect 518 1348 522 1352
rect 406 1338 410 1342
rect 318 1318 322 1322
rect 390 1318 394 1322
rect 374 1308 378 1312
rect 326 1298 330 1302
rect 286 1278 290 1282
rect 302 1278 306 1282
rect 222 1268 226 1272
rect 238 1268 242 1272
rect 198 1248 202 1252
rect 94 1168 98 1172
rect 78 1158 82 1162
rect 70 1128 74 1132
rect 14 1088 18 1092
rect 126 1218 130 1222
rect 126 1168 130 1172
rect 118 1148 122 1152
rect 294 1268 298 1272
rect 254 1208 258 1212
rect 182 1188 186 1192
rect 214 1188 218 1192
rect 166 1148 170 1152
rect 110 1138 114 1142
rect 118 1138 122 1142
rect 142 1138 146 1142
rect 174 1128 178 1132
rect 214 1168 218 1172
rect 230 1168 234 1172
rect 238 1168 242 1172
rect 182 1088 186 1092
rect 126 1068 130 1072
rect 134 1068 138 1072
rect 190 1059 194 1063
rect 22 978 26 982
rect 30 948 34 952
rect 78 948 82 952
rect 6 928 10 932
rect 14 868 18 872
rect 78 928 82 932
rect 62 878 66 882
rect 206 958 210 962
rect 198 948 202 952
rect 110 938 114 942
rect 126 938 130 942
rect 166 938 170 942
rect 150 928 154 932
rect 110 878 114 882
rect 22 848 26 852
rect 86 848 90 852
rect 142 768 146 772
rect 118 758 122 762
rect 102 748 106 752
rect 134 748 138 752
rect 54 738 58 742
rect 46 678 50 682
rect 126 738 130 742
rect 14 668 18 672
rect 62 668 66 672
rect 22 658 26 662
rect 54 658 58 662
rect 6 578 10 582
rect 22 568 26 572
rect 46 558 50 562
rect 102 688 106 692
rect 94 668 98 672
rect 78 648 82 652
rect 94 578 98 582
rect 86 558 90 562
rect 38 538 42 542
rect 46 538 50 542
rect 38 528 42 532
rect 70 528 74 532
rect 182 938 186 942
rect 206 888 210 892
rect 198 838 202 842
rect 174 828 178 832
rect 198 768 202 772
rect 190 758 194 762
rect 222 1158 226 1162
rect 390 1288 394 1292
rect 358 1258 362 1262
rect 302 1248 306 1252
rect 334 1248 338 1252
rect 318 1238 322 1242
rect 382 1248 386 1252
rect 342 1208 346 1212
rect 286 1158 290 1162
rect 318 1158 322 1162
rect 302 1148 306 1152
rect 382 1148 386 1152
rect 230 1088 234 1092
rect 230 1068 234 1072
rect 270 1068 274 1072
rect 246 1058 250 1062
rect 246 1038 250 1042
rect 270 1038 274 1042
rect 222 1028 226 1032
rect 230 968 234 972
rect 278 968 282 972
rect 222 958 226 962
rect 342 1128 346 1132
rect 302 1068 306 1072
rect 366 1088 370 1092
rect 302 968 306 972
rect 262 958 266 962
rect 278 958 282 962
rect 294 958 298 962
rect 334 958 338 962
rect 318 948 322 952
rect 246 938 250 942
rect 238 888 242 892
rect 230 878 234 882
rect 230 838 234 842
rect 166 748 170 752
rect 214 748 218 752
rect 302 938 306 942
rect 310 938 314 942
rect 294 868 298 872
rect 350 938 354 942
rect 350 878 354 882
rect 342 858 346 862
rect 334 848 338 852
rect 326 838 330 842
rect 278 818 282 822
rect 302 758 306 762
rect 246 748 250 752
rect 294 748 298 752
rect 190 738 194 742
rect 238 738 242 742
rect 254 738 258 742
rect 270 738 274 742
rect 174 698 178 702
rect 198 698 202 702
rect 214 678 218 682
rect 150 668 154 672
rect 142 578 146 582
rect 254 548 258 552
rect 190 538 194 542
rect 94 498 98 502
rect 118 498 122 502
rect 102 488 106 492
rect 150 478 154 482
rect 238 488 242 492
rect 118 458 122 462
rect 150 458 154 462
rect 6 448 10 452
rect 150 448 154 452
rect 22 438 26 442
rect 126 428 130 432
rect 22 298 26 302
rect 14 268 18 272
rect 158 388 162 392
rect 54 368 58 372
rect 150 368 154 372
rect 38 328 42 332
rect 46 298 50 302
rect 102 358 106 362
rect 62 288 66 292
rect 78 268 82 272
rect 126 348 130 352
rect 142 338 146 342
rect 110 278 114 282
rect 78 258 82 262
rect 102 258 106 262
rect 110 248 114 252
rect 142 248 146 252
rect 182 448 186 452
rect 182 388 186 392
rect 198 348 202 352
rect 254 348 258 352
rect 174 338 178 342
rect 230 338 234 342
rect 214 328 218 332
rect 246 328 250 332
rect 206 308 210 312
rect 198 288 202 292
rect 294 688 298 692
rect 342 768 346 772
rect 430 1328 434 1332
rect 526 1338 530 1342
rect 510 1328 514 1332
rect 454 1318 458 1322
rect 446 1308 450 1312
rect 526 1308 530 1312
rect 662 1408 666 1412
rect 630 1378 634 1382
rect 646 1368 650 1372
rect 630 1348 634 1352
rect 542 1328 546 1332
rect 534 1298 538 1302
rect 438 1288 442 1292
rect 454 1288 458 1292
rect 422 1268 426 1272
rect 446 1258 450 1262
rect 462 1248 466 1252
rect 494 1268 498 1272
rect 486 1258 490 1262
rect 430 1238 434 1242
rect 470 1238 474 1242
rect 462 1228 466 1232
rect 494 1228 498 1232
rect 438 1158 442 1162
rect 454 1158 458 1162
rect 438 1148 442 1152
rect 446 1128 450 1132
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 486 1168 490 1172
rect 534 1158 538 1162
rect 678 1388 682 1392
rect 638 1338 642 1342
rect 606 1328 610 1332
rect 598 1308 602 1312
rect 582 1288 586 1292
rect 622 1278 626 1282
rect 654 1268 658 1272
rect 582 1258 586 1262
rect 558 1248 562 1252
rect 622 1248 626 1252
rect 638 1248 642 1252
rect 654 1248 658 1252
rect 702 1368 706 1372
rect 694 1278 698 1282
rect 670 1268 674 1272
rect 694 1268 698 1272
rect 686 1258 690 1262
rect 638 1198 642 1202
rect 662 1198 666 1202
rect 622 1168 626 1172
rect 646 1168 650 1172
rect 590 1158 594 1162
rect 574 1148 578 1152
rect 590 1148 594 1152
rect 606 1148 610 1152
rect 462 1138 466 1142
rect 462 1128 466 1132
rect 446 1078 450 1082
rect 422 1068 426 1072
rect 438 1058 442 1062
rect 414 1018 418 1022
rect 382 938 386 942
rect 382 918 386 922
rect 406 918 410 922
rect 494 1108 498 1112
rect 486 1068 490 1072
rect 686 1158 690 1162
rect 662 1118 666 1122
rect 678 1138 682 1142
rect 670 1108 674 1112
rect 542 1088 546 1092
rect 590 1088 594 1092
rect 606 1088 610 1092
rect 886 1728 890 1732
rect 838 1718 842 1722
rect 870 1718 874 1722
rect 846 1708 850 1712
rect 870 1698 874 1702
rect 854 1668 858 1672
rect 878 1678 882 1682
rect 798 1658 802 1662
rect 766 1588 770 1592
rect 758 1558 762 1562
rect 790 1648 794 1652
rect 814 1648 818 1652
rect 838 1648 842 1652
rect 790 1588 794 1592
rect 782 1558 786 1562
rect 926 1818 930 1822
rect 950 1818 954 1822
rect 918 1778 922 1782
rect 982 1758 986 1762
rect 1014 1758 1018 1762
rect 958 1748 962 1752
rect 974 1738 978 1742
rect 942 1728 946 1732
rect 982 1728 986 1732
rect 974 1718 978 1722
rect 986 1703 990 1707
rect 993 1703 997 1707
rect 950 1698 954 1702
rect 958 1688 962 1692
rect 1046 2038 1050 2042
rect 1030 2028 1034 2032
rect 1126 2048 1130 2052
rect 1134 2028 1138 2032
rect 1126 2008 1130 2012
rect 1150 2008 1154 2012
rect 1078 1948 1082 1952
rect 1110 1948 1114 1952
rect 1062 1938 1066 1942
rect 1150 1938 1154 1942
rect 1158 1918 1162 1922
rect 1230 2088 1234 2092
rect 1302 2318 1306 2322
rect 1262 2308 1266 2312
rect 1318 2288 1322 2292
rect 1270 2278 1274 2282
rect 1286 2278 1290 2282
rect 1342 2298 1346 2302
rect 1366 2298 1370 2302
rect 1382 2288 1386 2292
rect 1326 2248 1330 2252
rect 1350 2248 1354 2252
rect 1382 2258 1386 2262
rect 1470 2338 1474 2342
rect 1446 2308 1450 2312
rect 1414 2278 1418 2282
rect 1422 2278 1426 2282
rect 1470 2298 1474 2302
rect 1486 2308 1490 2312
rect 1502 2298 1506 2302
rect 1534 2288 1538 2292
rect 1478 2268 1482 2272
rect 1550 2268 1554 2272
rect 1430 2258 1434 2262
rect 1462 2258 1466 2262
rect 1398 2248 1402 2252
rect 1406 2248 1410 2252
rect 1366 2238 1370 2242
rect 1278 2228 1282 2232
rect 1246 2178 1250 2182
rect 1366 2178 1370 2182
rect 1254 2148 1258 2152
rect 1302 2148 1306 2152
rect 1334 2148 1338 2152
rect 1846 2358 1850 2362
rect 1990 2358 1994 2362
rect 1702 2348 1706 2352
rect 1910 2348 1914 2352
rect 1934 2348 1938 2352
rect 2046 2348 2050 2352
rect 1566 2338 1570 2342
rect 1590 2338 1594 2342
rect 1678 2338 1682 2342
rect 1558 2228 1562 2232
rect 1886 2338 1890 2342
rect 1990 2338 1994 2342
rect 1782 2328 1786 2332
rect 1614 2298 1618 2302
rect 1750 2308 1754 2312
rect 1622 2278 1626 2282
rect 1718 2278 1722 2282
rect 1582 2248 1586 2252
rect 1822 2288 1826 2292
rect 1830 2268 1834 2272
rect 1646 2258 1650 2262
rect 1758 2248 1762 2252
rect 1822 2248 1826 2252
rect 1606 2238 1610 2242
rect 1630 2238 1634 2242
rect 1566 2218 1570 2222
rect 1598 2218 1602 2222
rect 1498 2203 1502 2207
rect 1505 2203 1509 2207
rect 1598 2188 1602 2192
rect 1486 2178 1490 2182
rect 1630 2168 1634 2172
rect 1654 2168 1658 2172
rect 1574 2158 1578 2162
rect 1590 2158 1594 2162
rect 1470 2148 1474 2152
rect 1502 2148 1506 2152
rect 1534 2148 1538 2152
rect 1662 2148 1666 2152
rect 1686 2148 1690 2152
rect 1310 2138 1314 2142
rect 1326 2138 1330 2142
rect 1382 2138 1386 2142
rect 1454 2138 1458 2142
rect 1246 2118 1250 2122
rect 1238 2078 1242 2082
rect 1238 2068 1242 2072
rect 1350 2118 1354 2122
rect 1438 2118 1442 2122
rect 1462 2118 1466 2122
rect 1310 2108 1314 2112
rect 1430 2108 1434 2112
rect 1350 2098 1354 2102
rect 1414 2098 1418 2102
rect 1366 2078 1370 2082
rect 1278 2058 1282 2062
rect 1286 2058 1290 2062
rect 1646 2138 1650 2142
rect 1702 2138 1706 2142
rect 1486 2108 1490 2112
rect 1446 2078 1450 2082
rect 1382 2058 1386 2062
rect 1398 2058 1402 2062
rect 1422 2058 1426 2062
rect 1214 2048 1218 2052
rect 1334 2048 1338 2052
rect 1270 1998 1274 2002
rect 1326 1998 1330 2002
rect 1262 1978 1266 1982
rect 1270 1978 1274 1982
rect 1182 1968 1186 1972
rect 1206 1958 1210 1962
rect 1318 1948 1322 1952
rect 1174 1928 1178 1932
rect 1182 1918 1186 1922
rect 1278 1938 1282 1942
rect 1302 1938 1306 1942
rect 1254 1928 1258 1932
rect 1238 1898 1242 1902
rect 1174 1878 1178 1882
rect 1254 1878 1258 1882
rect 1110 1868 1114 1872
rect 1166 1868 1170 1872
rect 1070 1858 1074 1862
rect 1142 1858 1146 1862
rect 1198 1858 1202 1862
rect 1150 1848 1154 1852
rect 1182 1848 1186 1852
rect 1038 1828 1042 1832
rect 1126 1788 1130 1792
rect 1030 1768 1034 1772
rect 1054 1768 1058 1772
rect 1102 1747 1106 1751
rect 1142 1768 1146 1772
rect 1214 1778 1218 1782
rect 1198 1768 1202 1772
rect 1166 1758 1170 1762
rect 1182 1758 1186 1762
rect 1158 1748 1162 1752
rect 1038 1738 1042 1742
rect 1038 1708 1042 1712
rect 1022 1698 1026 1702
rect 974 1678 978 1682
rect 1006 1678 1010 1682
rect 1142 1708 1146 1712
rect 1086 1688 1090 1692
rect 1134 1678 1138 1682
rect 926 1668 930 1672
rect 926 1658 930 1662
rect 934 1658 938 1662
rect 1014 1658 1018 1662
rect 1086 1658 1090 1662
rect 1166 1658 1170 1662
rect 846 1638 850 1642
rect 894 1638 898 1642
rect 878 1608 882 1612
rect 814 1578 818 1582
rect 774 1548 778 1552
rect 790 1548 794 1552
rect 766 1518 770 1522
rect 790 1528 794 1532
rect 734 1478 738 1482
rect 750 1468 754 1472
rect 758 1458 762 1462
rect 870 1558 874 1562
rect 814 1548 818 1552
rect 846 1538 850 1542
rect 806 1518 810 1522
rect 790 1498 794 1502
rect 774 1488 778 1492
rect 798 1478 802 1482
rect 750 1418 754 1422
rect 766 1418 770 1422
rect 734 1398 738 1402
rect 734 1368 738 1372
rect 710 1288 714 1292
rect 710 1248 714 1252
rect 710 1228 714 1232
rect 710 1138 714 1142
rect 502 1068 506 1072
rect 550 1068 554 1072
rect 646 1068 650 1072
rect 638 1058 642 1062
rect 686 1058 690 1062
rect 606 1048 610 1052
rect 662 1048 666 1052
rect 558 1038 562 1042
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 470 988 474 992
rect 454 968 458 972
rect 550 968 554 972
rect 526 948 530 952
rect 430 918 434 922
rect 414 888 418 892
rect 358 858 362 862
rect 382 858 386 862
rect 406 858 410 862
rect 462 928 466 932
rect 494 918 498 922
rect 454 908 458 912
rect 454 878 458 882
rect 446 868 450 872
rect 678 1028 682 1032
rect 614 1018 618 1022
rect 606 958 610 962
rect 678 968 682 972
rect 622 958 626 962
rect 654 958 658 962
rect 686 958 690 962
rect 606 948 610 952
rect 606 888 610 892
rect 550 878 554 882
rect 558 878 562 882
rect 582 878 586 882
rect 446 838 450 842
rect 366 788 370 792
rect 430 768 434 772
rect 334 758 338 762
rect 326 748 330 752
rect 482 803 486 807
rect 489 803 493 807
rect 534 798 538 802
rect 454 768 458 772
rect 494 768 498 772
rect 534 748 538 752
rect 702 1048 706 1052
rect 702 968 706 972
rect 758 1398 762 1402
rect 782 1398 786 1402
rect 742 1328 746 1332
rect 846 1458 850 1462
rect 862 1458 866 1462
rect 838 1448 842 1452
rect 854 1388 858 1392
rect 990 1638 994 1642
rect 1030 1638 1034 1642
rect 1030 1568 1034 1572
rect 934 1548 938 1552
rect 998 1548 1002 1552
rect 910 1488 914 1492
rect 894 1478 898 1482
rect 854 1358 858 1362
rect 862 1358 866 1362
rect 878 1358 882 1362
rect 814 1348 818 1352
rect 846 1348 850 1352
rect 886 1348 890 1352
rect 758 1338 762 1342
rect 790 1338 794 1342
rect 806 1338 810 1342
rect 846 1328 850 1332
rect 886 1328 890 1332
rect 742 1178 746 1182
rect 750 1158 754 1162
rect 742 1138 746 1142
rect 726 1118 730 1122
rect 718 1098 722 1102
rect 726 1058 730 1062
rect 734 1048 738 1052
rect 798 1308 802 1312
rect 782 1268 786 1272
rect 942 1538 946 1542
rect 966 1538 970 1542
rect 1022 1538 1026 1542
rect 934 1418 938 1422
rect 998 1518 1002 1522
rect 986 1503 990 1507
rect 993 1503 997 1507
rect 950 1468 954 1472
rect 1006 1468 1010 1472
rect 958 1458 962 1462
rect 990 1458 994 1462
rect 1022 1458 1026 1462
rect 950 1438 954 1442
rect 942 1408 946 1412
rect 934 1388 938 1392
rect 934 1358 938 1362
rect 902 1318 906 1322
rect 870 1288 874 1292
rect 894 1288 898 1292
rect 910 1288 914 1292
rect 934 1288 938 1292
rect 846 1278 850 1282
rect 862 1278 866 1282
rect 822 1268 826 1272
rect 774 1258 778 1262
rect 782 1258 786 1262
rect 830 1258 834 1262
rect 814 1248 818 1252
rect 894 1228 898 1232
rect 806 1198 810 1202
rect 790 1188 794 1192
rect 814 1178 818 1182
rect 798 1168 802 1172
rect 806 1148 810 1152
rect 782 1138 786 1142
rect 790 1058 794 1062
rect 758 1018 762 1022
rect 694 948 698 952
rect 718 948 722 952
rect 742 948 746 952
rect 782 948 786 952
rect 646 888 650 892
rect 758 928 762 932
rect 902 1198 906 1202
rect 886 1168 890 1172
rect 830 1148 834 1152
rect 822 1098 826 1102
rect 886 1128 890 1132
rect 870 1098 874 1102
rect 830 1088 834 1092
rect 846 1088 850 1092
rect 806 918 810 922
rect 838 998 842 1002
rect 870 988 874 992
rect 846 918 850 922
rect 814 888 818 892
rect 710 868 714 872
rect 854 868 858 872
rect 606 858 610 862
rect 654 858 658 862
rect 574 848 578 852
rect 702 848 706 852
rect 702 838 706 842
rect 582 798 586 802
rect 630 778 634 782
rect 558 768 562 772
rect 614 748 618 752
rect 646 748 650 752
rect 670 748 674 752
rect 374 738 378 742
rect 446 738 450 742
rect 446 718 450 722
rect 342 698 346 702
rect 318 678 322 682
rect 326 668 330 672
rect 358 678 362 682
rect 398 678 402 682
rect 350 668 354 672
rect 454 668 458 672
rect 462 668 466 672
rect 526 738 530 742
rect 542 738 546 742
rect 630 738 634 742
rect 518 678 522 682
rect 510 668 514 672
rect 294 658 298 662
rect 374 658 378 662
rect 398 658 402 662
rect 470 658 474 662
rect 294 648 298 652
rect 310 648 314 652
rect 414 648 418 652
rect 342 628 346 632
rect 270 588 274 592
rect 294 588 298 592
rect 286 538 290 542
rect 326 538 330 542
rect 278 528 282 532
rect 286 498 290 502
rect 310 498 314 502
rect 302 478 306 482
rect 294 468 298 472
rect 518 648 522 652
rect 534 708 538 712
rect 558 678 562 682
rect 550 668 554 672
rect 582 668 586 672
rect 686 718 690 722
rect 670 688 674 692
rect 734 858 738 862
rect 750 858 754 862
rect 806 858 810 862
rect 790 828 794 832
rect 742 768 746 772
rect 766 758 770 762
rect 726 748 730 752
rect 758 748 762 752
rect 718 728 722 732
rect 710 698 714 702
rect 646 668 650 672
rect 678 668 682 672
rect 702 668 706 672
rect 526 618 530 622
rect 502 608 506 612
rect 482 603 486 607
rect 489 603 493 607
rect 518 598 522 602
rect 574 648 578 652
rect 582 648 586 652
rect 774 728 778 732
rect 766 678 770 682
rect 774 678 778 682
rect 750 668 754 672
rect 630 658 634 662
rect 686 658 690 662
rect 734 658 738 662
rect 766 658 770 662
rect 590 638 594 642
rect 606 638 610 642
rect 638 638 642 642
rect 518 578 522 582
rect 446 558 450 562
rect 454 558 458 562
rect 550 568 554 572
rect 662 608 666 612
rect 574 558 578 562
rect 622 558 626 562
rect 638 558 642 562
rect 662 558 666 562
rect 406 548 410 552
rect 470 548 474 552
rect 510 548 514 552
rect 366 538 370 542
rect 374 498 378 502
rect 358 468 362 472
rect 270 388 274 392
rect 318 458 322 462
rect 342 458 346 462
rect 326 448 330 452
rect 366 438 370 442
rect 422 518 426 522
rect 462 538 466 542
rect 486 498 490 502
rect 494 498 498 502
rect 438 488 442 492
rect 454 488 458 492
rect 462 468 466 472
rect 454 448 458 452
rect 482 403 486 407
rect 489 403 493 407
rect 350 368 354 372
rect 374 368 378 372
rect 390 368 394 372
rect 294 348 298 352
rect 334 318 338 322
rect 310 308 314 312
rect 302 298 306 302
rect 310 298 314 302
rect 174 218 178 222
rect 158 168 162 172
rect 262 168 266 172
rect 334 168 338 172
rect 70 158 74 162
rect 126 158 130 162
rect 150 158 154 162
rect 174 158 178 162
rect 262 158 266 162
rect 6 148 10 152
rect 102 148 106 152
rect 118 148 122 152
rect 150 148 154 152
rect 142 138 146 142
rect 70 128 74 132
rect 6 78 10 82
rect 142 68 146 72
rect 206 148 210 152
rect 198 138 202 142
rect 214 138 218 142
rect 174 98 178 102
rect 246 128 250 132
rect 342 128 346 132
rect 230 118 234 122
rect 318 118 322 122
rect 270 98 274 102
rect 294 88 298 92
rect 214 78 218 82
rect 278 78 282 82
rect 318 78 322 82
rect 142 58 146 62
rect 190 58 194 62
rect 414 358 418 362
rect 478 358 482 362
rect 398 348 402 352
rect 414 348 418 352
rect 446 348 450 352
rect 382 338 386 342
rect 406 338 410 342
rect 382 298 386 302
rect 366 259 370 263
rect 502 288 506 292
rect 486 278 490 282
rect 470 268 474 272
rect 422 258 426 262
rect 502 258 506 262
rect 414 228 418 232
rect 470 218 474 222
rect 482 203 486 207
rect 489 203 493 207
rect 438 188 442 192
rect 486 178 490 182
rect 614 548 618 552
rect 662 548 666 552
rect 566 538 570 542
rect 622 538 626 542
rect 638 538 642 542
rect 582 528 586 532
rect 606 528 610 532
rect 582 498 586 502
rect 606 498 610 502
rect 534 468 538 472
rect 526 428 530 432
rect 518 368 522 372
rect 518 348 522 352
rect 526 338 530 342
rect 526 248 530 252
rect 646 468 650 472
rect 622 458 626 462
rect 598 448 602 452
rect 582 438 586 442
rect 550 418 554 422
rect 854 848 858 852
rect 894 1008 898 1012
rect 942 1268 946 1272
rect 958 1348 962 1352
rect 1190 1708 1194 1712
rect 1190 1688 1194 1692
rect 1182 1648 1186 1652
rect 1142 1608 1146 1612
rect 1174 1608 1178 1612
rect 1126 1598 1130 1602
rect 1182 1578 1186 1582
rect 1054 1548 1058 1552
rect 1118 1548 1122 1552
rect 1150 1548 1154 1552
rect 1182 1548 1186 1552
rect 1038 1538 1042 1542
rect 1078 1538 1082 1542
rect 1094 1538 1098 1542
rect 1134 1528 1138 1532
rect 1070 1518 1074 1522
rect 1086 1518 1090 1522
rect 1054 1498 1058 1502
rect 1110 1508 1114 1512
rect 1166 1498 1170 1502
rect 1182 1498 1186 1502
rect 1070 1488 1074 1492
rect 1086 1478 1090 1482
rect 1102 1468 1106 1472
rect 1174 1428 1178 1432
rect 1166 1418 1170 1422
rect 1118 1398 1122 1402
rect 1070 1388 1074 1392
rect 1046 1348 1050 1352
rect 1062 1348 1066 1352
rect 1030 1338 1034 1342
rect 990 1318 994 1322
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 1014 1278 1018 1282
rect 1022 1278 1026 1282
rect 1014 1268 1018 1272
rect 974 1258 978 1262
rect 1006 1258 1010 1262
rect 926 1248 930 1252
rect 950 1228 954 1232
rect 950 1198 954 1202
rect 942 1188 946 1192
rect 934 1168 938 1172
rect 942 1148 946 1152
rect 1030 1228 1034 1232
rect 1014 1198 1018 1202
rect 974 1158 978 1162
rect 958 1148 962 1152
rect 966 1148 970 1152
rect 926 1088 930 1092
rect 950 1068 954 1072
rect 918 1058 922 1062
rect 902 998 906 1002
rect 902 958 906 962
rect 878 928 882 932
rect 878 888 882 892
rect 902 878 906 882
rect 886 858 890 862
rect 1046 1258 1050 1262
rect 1038 1218 1042 1222
rect 1054 1218 1058 1222
rect 990 1148 994 1152
rect 1022 1148 1026 1152
rect 998 1128 1002 1132
rect 1046 1168 1050 1172
rect 1046 1138 1050 1142
rect 1094 1368 1098 1372
rect 1086 1268 1090 1272
rect 1142 1358 1146 1362
rect 1158 1358 1162 1362
rect 1134 1348 1138 1352
rect 1134 1318 1138 1322
rect 1294 1908 1298 1912
rect 1366 2008 1370 2012
rect 1350 1968 1354 1972
rect 1438 2018 1442 2022
rect 1494 2068 1498 2072
rect 1478 2058 1482 2062
rect 1478 2018 1482 2022
rect 1498 2003 1502 2007
rect 1505 2003 1509 2007
rect 1446 1998 1450 2002
rect 1398 1978 1402 1982
rect 1414 1978 1418 1982
rect 1406 1948 1410 1952
rect 1430 1948 1434 1952
rect 1470 1948 1474 1952
rect 1310 1888 1314 1892
rect 1318 1888 1322 1892
rect 1262 1868 1266 1872
rect 1270 1868 1274 1872
rect 1310 1858 1314 1862
rect 1326 1848 1330 1852
rect 1350 1788 1354 1792
rect 1262 1758 1266 1762
rect 1294 1758 1298 1762
rect 1350 1758 1354 1762
rect 1278 1738 1282 1742
rect 1230 1708 1234 1712
rect 1222 1698 1226 1702
rect 1246 1688 1250 1692
rect 1302 1738 1306 1742
rect 1318 1738 1322 1742
rect 1310 1718 1314 1722
rect 1294 1708 1298 1712
rect 1286 1678 1290 1682
rect 1310 1678 1314 1682
rect 1238 1668 1242 1672
rect 1294 1668 1298 1672
rect 1222 1658 1226 1662
rect 1246 1658 1250 1662
rect 1262 1658 1266 1662
rect 1278 1658 1282 1662
rect 1238 1618 1242 1622
rect 1286 1638 1290 1642
rect 1302 1628 1306 1632
rect 1262 1568 1266 1572
rect 1246 1558 1250 1562
rect 1278 1558 1282 1562
rect 1238 1548 1242 1552
rect 1326 1698 1330 1702
rect 1446 1938 1450 1942
rect 1374 1928 1378 1932
rect 1414 1918 1418 1922
rect 1446 1898 1450 1902
rect 1398 1868 1402 1872
rect 1430 1868 1434 1872
rect 1446 1868 1450 1872
rect 1566 2108 1570 2112
rect 1606 2098 1610 2102
rect 1598 2078 1602 2082
rect 1542 2068 1546 2072
rect 1590 2068 1594 2072
rect 1670 2118 1674 2122
rect 1622 2108 1626 2112
rect 1654 2108 1658 2112
rect 1614 2078 1618 2082
rect 1702 2078 1706 2082
rect 1638 2068 1642 2072
rect 1670 2068 1674 2072
rect 1678 2068 1682 2072
rect 1734 2068 1738 2072
rect 1566 2008 1570 2012
rect 1662 2038 1666 2042
rect 1686 2038 1690 2042
rect 1614 2008 1618 2012
rect 1606 1988 1610 1992
rect 1630 1978 1634 1982
rect 1662 1978 1666 1982
rect 1606 1968 1610 1972
rect 1574 1948 1578 1952
rect 1694 1968 1698 1972
rect 1494 1938 1498 1942
rect 1526 1938 1530 1942
rect 1478 1928 1482 1932
rect 1534 1908 1538 1912
rect 1478 1888 1482 1892
rect 1486 1888 1490 1892
rect 1518 1888 1522 1892
rect 1550 1878 1554 1882
rect 1526 1868 1530 1872
rect 1542 1868 1546 1872
rect 1414 1858 1418 1862
rect 1502 1858 1506 1862
rect 1390 1838 1394 1842
rect 1382 1798 1386 1802
rect 1462 1848 1466 1852
rect 1470 1838 1474 1842
rect 1478 1838 1482 1842
rect 1430 1808 1434 1812
rect 1498 1803 1502 1807
rect 1505 1803 1509 1807
rect 1710 1948 1714 1952
rect 1582 1928 1586 1932
rect 1606 1888 1610 1892
rect 1654 1888 1658 1892
rect 1582 1868 1586 1872
rect 1622 1868 1626 1872
rect 1566 1848 1570 1852
rect 1574 1848 1578 1852
rect 1518 1788 1522 1792
rect 1558 1788 1562 1792
rect 1494 1758 1498 1762
rect 1454 1748 1458 1752
rect 1486 1748 1490 1752
rect 1374 1738 1378 1742
rect 1422 1728 1426 1732
rect 1398 1718 1402 1722
rect 1422 1678 1426 1682
rect 1294 1588 1298 1592
rect 1334 1588 1338 1592
rect 1358 1588 1362 1592
rect 1302 1558 1306 1562
rect 1334 1548 1338 1552
rect 1262 1538 1266 1542
rect 1246 1518 1250 1522
rect 1214 1498 1218 1502
rect 1230 1478 1234 1482
rect 1214 1448 1218 1452
rect 1206 1378 1210 1382
rect 1198 1358 1202 1362
rect 1166 1338 1170 1342
rect 1158 1298 1162 1302
rect 1198 1288 1202 1292
rect 1190 1278 1194 1282
rect 1142 1268 1146 1272
rect 1102 1258 1106 1262
rect 1182 1258 1186 1262
rect 1110 1248 1114 1252
rect 1102 1218 1106 1222
rect 1150 1248 1154 1252
rect 1174 1248 1178 1252
rect 1142 1188 1146 1192
rect 1094 1178 1098 1182
rect 1070 1158 1074 1162
rect 1086 1158 1090 1162
rect 1078 1138 1082 1142
rect 1046 1128 1050 1132
rect 1006 1118 1010 1122
rect 1038 1118 1042 1122
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 1038 1108 1042 1112
rect 974 1068 978 1072
rect 974 1048 978 1052
rect 982 1048 986 1052
rect 950 1008 954 1012
rect 934 998 938 1002
rect 950 998 954 1002
rect 958 958 962 962
rect 958 948 962 952
rect 966 948 970 952
rect 942 888 946 892
rect 942 858 946 862
rect 894 848 898 852
rect 918 848 922 852
rect 862 838 866 842
rect 822 828 826 832
rect 814 768 818 772
rect 854 728 858 732
rect 886 818 890 822
rect 878 778 882 782
rect 886 778 890 782
rect 910 778 914 782
rect 910 768 914 772
rect 926 808 930 812
rect 966 918 970 922
rect 966 898 970 902
rect 1038 1058 1042 1062
rect 1006 1048 1010 1052
rect 1030 1048 1034 1052
rect 998 988 1002 992
rect 982 978 986 982
rect 998 968 1002 972
rect 982 938 986 942
rect 986 903 990 907
rect 993 903 997 907
rect 974 888 978 892
rect 1014 1038 1018 1042
rect 1030 958 1034 962
rect 1014 948 1018 952
rect 1022 948 1026 952
rect 1022 938 1026 942
rect 1022 908 1026 912
rect 1054 1118 1058 1122
rect 1078 1118 1082 1122
rect 1054 1098 1058 1102
rect 1134 1148 1138 1152
rect 1158 1218 1162 1222
rect 1222 1318 1226 1322
rect 1382 1648 1386 1652
rect 1422 1648 1426 1652
rect 1438 1738 1442 1742
rect 1486 1738 1490 1742
rect 1478 1708 1482 1712
rect 1550 1758 1554 1762
rect 1534 1748 1538 1752
rect 1550 1748 1554 1752
rect 1590 1788 1594 1792
rect 1614 1858 1618 1862
rect 1654 1858 1658 1862
rect 1646 1848 1650 1852
rect 1694 1858 1698 1862
rect 1606 1838 1610 1842
rect 1622 1818 1626 1822
rect 1598 1758 1602 1762
rect 1662 1758 1666 1762
rect 1686 1758 1690 1762
rect 1566 1748 1570 1752
rect 1606 1748 1610 1752
rect 1702 1748 1706 1752
rect 1558 1738 1562 1742
rect 1726 2008 1730 2012
rect 1878 2298 1882 2302
rect 1862 2288 1866 2292
rect 1854 2238 1858 2242
rect 1830 2228 1834 2232
rect 1782 2218 1786 2222
rect 1806 2148 1810 2152
rect 1814 2138 1818 2142
rect 1806 2128 1810 2132
rect 1766 2108 1770 2112
rect 1766 2078 1770 2082
rect 1798 2078 1802 2082
rect 1734 1968 1738 1972
rect 1726 1948 1730 1952
rect 1742 1878 1746 1882
rect 1806 2048 1810 2052
rect 1990 2328 1994 2332
rect 1910 2308 1914 2312
rect 1958 2308 1962 2312
rect 1902 2288 1906 2292
rect 1902 2278 1906 2282
rect 2018 2303 2022 2307
rect 2025 2303 2029 2307
rect 2086 2358 2090 2362
rect 2094 2358 2098 2362
rect 2214 2358 2218 2362
rect 2454 2358 2458 2362
rect 2070 2348 2074 2352
rect 2094 2348 2098 2352
rect 2238 2348 2242 2352
rect 2270 2348 2274 2352
rect 2334 2348 2338 2352
rect 2366 2348 2370 2352
rect 2102 2328 2106 2332
rect 2054 2318 2058 2322
rect 2014 2278 2018 2282
rect 2038 2278 2042 2282
rect 1926 2268 1930 2272
rect 1950 2268 1954 2272
rect 1894 2258 1898 2262
rect 1878 2138 1882 2142
rect 1966 2258 1970 2262
rect 1998 2258 2002 2262
rect 2046 2248 2050 2252
rect 1974 2238 1978 2242
rect 1998 2238 2002 2242
rect 1958 2218 1962 2222
rect 1918 2178 1922 2182
rect 1926 2128 1930 2132
rect 1910 2098 1914 2102
rect 1990 2218 1994 2222
rect 1974 2178 1978 2182
rect 1910 2088 1914 2092
rect 1934 2088 1938 2092
rect 1950 2088 1954 2092
rect 1958 2088 1962 2092
rect 1886 2078 1890 2082
rect 1870 2068 1874 2072
rect 1902 2068 1906 2072
rect 1878 2028 1882 2032
rect 1862 1978 1866 1982
rect 1814 1958 1818 1962
rect 1950 2078 1954 2082
rect 2054 2158 2058 2162
rect 1998 2148 2002 2152
rect 2078 2148 2082 2152
rect 2046 2138 2050 2142
rect 2018 2103 2022 2107
rect 2025 2103 2029 2107
rect 2022 2078 2026 2082
rect 1918 2068 1922 2072
rect 1942 2058 1946 2062
rect 1974 2058 1978 2062
rect 1990 2058 1994 2062
rect 1926 2048 1930 2052
rect 1966 2048 1970 2052
rect 1950 1998 1954 2002
rect 1998 1958 2002 1962
rect 1934 1948 1938 1952
rect 1958 1948 1962 1952
rect 1822 1938 1826 1942
rect 1790 1888 1794 1892
rect 1798 1868 1802 1872
rect 1830 1868 1834 1872
rect 1742 1808 1746 1812
rect 1718 1788 1722 1792
rect 1814 1838 1818 1842
rect 1838 1838 1842 1842
rect 1782 1828 1786 1832
rect 1910 1938 1914 1942
rect 1878 1918 1882 1922
rect 1886 1918 1890 1922
rect 1902 1908 1906 1912
rect 1862 1888 1866 1892
rect 1894 1888 1898 1892
rect 1870 1878 1874 1882
rect 1854 1858 1858 1862
rect 1886 1858 1890 1862
rect 1774 1808 1778 1812
rect 1814 1808 1818 1812
rect 1846 1808 1850 1812
rect 1742 1778 1746 1782
rect 1758 1778 1762 1782
rect 1718 1768 1722 1772
rect 1806 1768 1810 1772
rect 1758 1758 1762 1762
rect 1718 1748 1722 1752
rect 1734 1748 1738 1752
rect 1750 1748 1754 1752
rect 1710 1738 1714 1742
rect 1654 1728 1658 1732
rect 1694 1728 1698 1732
rect 1654 1698 1658 1702
rect 1726 1698 1730 1702
rect 1646 1688 1650 1692
rect 1446 1658 1450 1662
rect 1494 1658 1498 1662
rect 1558 1658 1562 1662
rect 1606 1658 1610 1662
rect 1430 1628 1434 1632
rect 1542 1618 1546 1622
rect 1422 1558 1426 1562
rect 1358 1508 1362 1512
rect 1310 1498 1314 1502
rect 1326 1488 1330 1492
rect 1294 1468 1298 1472
rect 1350 1478 1354 1482
rect 1446 1558 1450 1562
rect 1526 1608 1530 1612
rect 1498 1603 1502 1607
rect 1505 1603 1509 1607
rect 1486 1558 1490 1562
rect 1614 1648 1618 1652
rect 1622 1648 1626 1652
rect 1598 1618 1602 1622
rect 1574 1608 1578 1612
rect 1558 1558 1562 1562
rect 1590 1558 1594 1562
rect 1454 1548 1458 1552
rect 1430 1538 1434 1542
rect 1470 1538 1474 1542
rect 1478 1538 1482 1542
rect 1534 1528 1538 1532
rect 1398 1508 1402 1512
rect 1382 1488 1386 1492
rect 1366 1478 1370 1482
rect 1430 1468 1434 1472
rect 1270 1408 1274 1412
rect 1238 1348 1242 1352
rect 1254 1348 1258 1352
rect 1334 1378 1338 1382
rect 1358 1358 1362 1362
rect 1262 1338 1266 1342
rect 1270 1318 1274 1322
rect 1318 1318 1322 1322
rect 1246 1308 1250 1312
rect 1310 1298 1314 1302
rect 1286 1288 1290 1292
rect 1158 1208 1162 1212
rect 1214 1208 1218 1212
rect 1150 1128 1154 1132
rect 1110 1108 1114 1112
rect 1142 1108 1146 1112
rect 1134 1078 1138 1082
rect 1054 1058 1058 1062
rect 1070 1048 1074 1052
rect 1102 1048 1106 1052
rect 1118 1048 1122 1052
rect 1062 1038 1066 1042
rect 1078 1018 1082 1022
rect 1070 947 1074 951
rect 1078 928 1082 932
rect 1030 888 1034 892
rect 966 868 970 872
rect 958 858 962 862
rect 1014 848 1018 852
rect 966 838 970 842
rect 950 818 954 822
rect 950 798 954 802
rect 942 768 946 772
rect 918 758 922 762
rect 926 758 930 762
rect 894 738 898 742
rect 926 738 930 742
rect 942 738 946 742
rect 950 738 954 742
rect 830 708 834 712
rect 830 678 834 682
rect 862 718 866 722
rect 902 718 906 722
rect 894 698 898 702
rect 926 698 930 702
rect 910 688 914 692
rect 878 678 882 682
rect 918 678 922 682
rect 902 668 906 672
rect 934 668 938 672
rect 798 658 802 662
rect 822 658 826 662
rect 846 658 850 662
rect 910 658 914 662
rect 790 648 794 652
rect 782 588 786 592
rect 862 648 866 652
rect 878 628 882 632
rect 878 598 882 602
rect 854 588 858 592
rect 806 578 810 582
rect 726 568 730 572
rect 814 568 818 572
rect 678 558 682 562
rect 774 558 778 562
rect 870 558 874 562
rect 958 688 962 692
rect 934 648 938 652
rect 942 588 946 592
rect 718 547 722 551
rect 806 548 810 552
rect 830 548 834 552
rect 918 548 922 552
rect 958 548 962 552
rect 694 488 698 492
rect 710 488 714 492
rect 758 488 762 492
rect 790 488 794 492
rect 710 478 714 482
rect 734 468 738 472
rect 798 468 802 472
rect 726 458 730 462
rect 742 458 746 462
rect 774 448 778 452
rect 726 378 730 382
rect 550 368 554 372
rect 558 358 562 362
rect 670 348 674 352
rect 678 348 682 352
rect 702 348 706 352
rect 542 338 546 342
rect 566 338 570 342
rect 550 328 554 332
rect 566 328 570 332
rect 638 318 642 322
rect 614 298 618 302
rect 590 268 594 272
rect 550 238 554 242
rect 534 168 538 172
rect 358 118 362 122
rect 414 88 418 92
rect 430 88 434 92
rect 446 98 450 102
rect 422 78 426 82
rect 438 78 442 82
rect 326 68 330 72
rect 166 48 170 52
rect 206 48 210 52
rect 310 48 314 52
rect 358 48 362 52
rect 438 68 442 72
rect 454 68 458 72
rect 430 58 434 62
rect 462 58 466 62
rect 482 3 486 7
rect 489 3 493 7
rect 582 258 586 262
rect 606 248 610 252
rect 606 238 610 242
rect 598 148 602 152
rect 662 278 666 282
rect 654 268 658 272
rect 614 228 618 232
rect 646 228 650 232
rect 646 178 650 182
rect 622 168 626 172
rect 646 168 650 172
rect 654 158 658 162
rect 614 148 618 152
rect 566 118 570 122
rect 582 78 586 82
rect 558 68 562 72
rect 654 118 658 122
rect 862 538 866 542
rect 854 528 858 532
rect 846 448 850 452
rect 822 438 826 442
rect 862 408 866 412
rect 854 368 858 372
rect 822 348 826 352
rect 766 338 770 342
rect 686 308 690 312
rect 734 308 738 312
rect 758 278 762 282
rect 710 258 714 262
rect 734 258 738 262
rect 766 258 770 262
rect 702 208 706 212
rect 718 148 722 152
rect 742 138 746 142
rect 694 128 698 132
rect 830 328 834 332
rect 822 288 826 292
rect 790 268 794 272
rect 806 268 810 272
rect 782 258 786 262
rect 806 158 810 162
rect 782 128 786 132
rect 710 118 714 122
rect 750 118 754 122
rect 694 88 698 92
rect 710 88 714 92
rect 846 328 850 332
rect 838 288 842 292
rect 838 268 842 272
rect 886 538 890 542
rect 926 538 930 542
rect 934 528 938 532
rect 926 508 930 512
rect 926 488 930 492
rect 886 468 890 472
rect 878 458 882 462
rect 910 458 914 462
rect 902 408 906 412
rect 870 358 874 362
rect 918 368 922 372
rect 934 448 938 452
rect 950 428 954 432
rect 982 778 986 782
rect 982 748 986 752
rect 986 703 990 707
rect 993 703 997 707
rect 1022 788 1026 792
rect 1022 778 1026 782
rect 1046 838 1050 842
rect 1038 768 1042 772
rect 1030 758 1034 762
rect 1046 758 1050 762
rect 1038 748 1042 752
rect 1078 848 1082 852
rect 1126 1018 1130 1022
rect 1150 1088 1154 1092
rect 1150 1018 1154 1022
rect 1142 1008 1146 1012
rect 1110 998 1114 1002
rect 1134 988 1138 992
rect 1118 968 1122 972
rect 1238 1268 1242 1272
rect 1302 1158 1306 1162
rect 1182 1148 1186 1152
rect 1230 1148 1234 1152
rect 1206 1128 1210 1132
rect 1198 1108 1202 1112
rect 1190 1098 1194 1102
rect 1166 998 1170 1002
rect 1190 968 1194 972
rect 1126 938 1130 942
rect 1150 938 1154 942
rect 1102 848 1106 852
rect 1102 768 1106 772
rect 1086 758 1090 762
rect 1094 758 1098 762
rect 1046 738 1050 742
rect 1062 738 1066 742
rect 1078 738 1082 742
rect 1022 718 1026 722
rect 1014 638 1018 642
rect 998 568 1002 572
rect 986 503 990 507
rect 993 503 997 507
rect 1014 488 1018 492
rect 998 478 1002 482
rect 982 468 986 472
rect 974 418 978 422
rect 966 368 970 372
rect 886 348 890 352
rect 926 348 930 352
rect 934 348 938 352
rect 870 328 874 332
rect 894 328 898 332
rect 918 328 922 332
rect 854 298 858 302
rect 822 148 826 152
rect 838 148 842 152
rect 894 258 898 262
rect 1038 728 1042 732
rect 1062 698 1066 702
rect 1046 678 1050 682
rect 1070 678 1074 682
rect 1070 648 1074 652
rect 1078 648 1082 652
rect 1094 658 1098 662
rect 1086 578 1090 582
rect 1150 878 1154 882
rect 1142 868 1146 872
rect 1222 1108 1226 1112
rect 1230 1098 1234 1102
rect 1294 1118 1298 1122
rect 1286 1098 1290 1102
rect 1262 1078 1266 1082
rect 1238 1048 1242 1052
rect 1222 1018 1226 1022
rect 1214 988 1218 992
rect 1198 948 1202 952
rect 1206 948 1210 952
rect 1174 928 1178 932
rect 1238 940 1242 944
rect 1270 1048 1274 1052
rect 1270 978 1274 982
rect 1334 1308 1338 1312
rect 1350 1308 1354 1312
rect 1382 1308 1386 1312
rect 1430 1418 1434 1422
rect 1382 1288 1386 1292
rect 1398 1288 1402 1292
rect 1422 1278 1426 1282
rect 1366 1268 1370 1272
rect 1414 1268 1418 1272
rect 1390 1208 1394 1212
rect 1374 1158 1378 1162
rect 1366 1138 1370 1142
rect 1342 1128 1346 1132
rect 1334 1098 1338 1102
rect 1358 1108 1362 1112
rect 1350 1098 1354 1102
rect 1342 1068 1346 1072
rect 1318 1048 1322 1052
rect 1294 1028 1298 1032
rect 1222 918 1226 922
rect 1174 898 1178 902
rect 1206 898 1210 902
rect 1166 888 1170 892
rect 1230 888 1234 892
rect 1198 868 1202 872
rect 1206 868 1210 872
rect 1158 858 1162 862
rect 1182 858 1186 862
rect 1166 848 1170 852
rect 1198 848 1202 852
rect 1214 848 1218 852
rect 1206 828 1210 832
rect 1182 808 1186 812
rect 1134 798 1138 802
rect 1174 758 1178 762
rect 1158 748 1162 752
rect 1174 738 1178 742
rect 1150 728 1154 732
rect 1118 718 1122 722
rect 1134 718 1138 722
rect 1118 658 1122 662
rect 1142 678 1146 682
rect 1158 708 1162 712
rect 1166 678 1170 682
rect 1198 738 1202 742
rect 1182 688 1186 692
rect 1198 688 1202 692
rect 1134 648 1138 652
rect 1086 568 1090 572
rect 1102 568 1106 572
rect 1054 558 1058 562
rect 1126 568 1130 572
rect 1118 558 1122 562
rect 1102 548 1106 552
rect 1030 528 1034 532
rect 1094 528 1098 532
rect 1078 508 1082 512
rect 1182 648 1186 652
rect 1158 638 1162 642
rect 1254 928 1258 932
rect 1262 918 1266 922
rect 1254 878 1258 882
rect 1246 868 1250 872
rect 1278 898 1282 902
rect 1270 878 1274 882
rect 1254 858 1258 862
rect 1270 848 1274 852
rect 1302 1008 1306 1012
rect 1318 928 1322 932
rect 1294 878 1298 882
rect 1294 868 1298 872
rect 1310 868 1314 872
rect 1414 1218 1418 1222
rect 1526 1488 1530 1492
rect 1494 1478 1498 1482
rect 1486 1468 1490 1472
rect 1510 1458 1514 1462
rect 1470 1448 1474 1452
rect 1478 1448 1482 1452
rect 1526 1448 1530 1452
rect 1462 1408 1466 1412
rect 1686 1668 1690 1672
rect 1710 1668 1714 1672
rect 1702 1658 1706 1662
rect 1654 1648 1658 1652
rect 1678 1648 1682 1652
rect 1606 1558 1610 1562
rect 1638 1558 1642 1562
rect 1574 1538 1578 1542
rect 1558 1478 1562 1482
rect 1590 1468 1594 1472
rect 1558 1448 1562 1452
rect 1550 1418 1554 1422
rect 1498 1403 1502 1407
rect 1505 1403 1509 1407
rect 1558 1388 1562 1392
rect 1550 1378 1554 1382
rect 1462 1358 1466 1362
rect 1454 1298 1458 1302
rect 1438 1268 1442 1272
rect 1478 1358 1482 1362
rect 1590 1448 1594 1452
rect 1582 1418 1586 1422
rect 1502 1348 1506 1352
rect 1534 1348 1538 1352
rect 1566 1348 1570 1352
rect 1478 1338 1482 1342
rect 1486 1338 1490 1342
rect 1470 1278 1474 1282
rect 1438 1218 1442 1222
rect 1550 1338 1554 1342
rect 1518 1308 1522 1312
rect 1502 1278 1506 1282
rect 1498 1203 1502 1207
rect 1505 1203 1509 1207
rect 1462 1168 1466 1172
rect 1398 1158 1402 1162
rect 1438 1158 1442 1162
rect 1462 1158 1466 1162
rect 1566 1308 1570 1312
rect 1542 1288 1546 1292
rect 1590 1338 1594 1342
rect 1598 1278 1602 1282
rect 1558 1259 1562 1263
rect 1630 1508 1634 1512
rect 1614 1488 1618 1492
rect 1646 1468 1650 1472
rect 1718 1618 1722 1622
rect 1862 1838 1866 1842
rect 1894 1838 1898 1842
rect 1838 1748 1842 1752
rect 1782 1688 1786 1692
rect 1822 1688 1826 1692
rect 1742 1678 1746 1682
rect 1830 1678 1834 1682
rect 1734 1658 1738 1662
rect 1750 1658 1754 1662
rect 1774 1658 1778 1662
rect 1758 1648 1762 1652
rect 1806 1638 1810 1642
rect 1734 1568 1738 1572
rect 1758 1568 1762 1572
rect 1750 1558 1754 1562
rect 1822 1558 1826 1562
rect 1774 1548 1778 1552
rect 1662 1538 1666 1542
rect 1718 1538 1722 1542
rect 1734 1538 1738 1542
rect 1782 1538 1786 1542
rect 1790 1538 1794 1542
rect 1830 1538 1834 1542
rect 1702 1528 1706 1532
rect 1686 1498 1690 1502
rect 1662 1488 1666 1492
rect 1702 1488 1706 1492
rect 1654 1358 1658 1362
rect 1678 1468 1682 1472
rect 1726 1478 1730 1482
rect 1750 1528 1754 1532
rect 1782 1498 1786 1502
rect 1742 1478 1746 1482
rect 1726 1448 1730 1452
rect 1678 1368 1682 1372
rect 1646 1348 1650 1352
rect 1694 1348 1698 1352
rect 1718 1348 1722 1352
rect 1646 1298 1650 1302
rect 1726 1338 1730 1342
rect 1694 1308 1698 1312
rect 1654 1288 1658 1292
rect 1614 1258 1618 1262
rect 1654 1258 1658 1262
rect 1606 1248 1610 1252
rect 1638 1248 1642 1252
rect 1534 1238 1538 1242
rect 1582 1168 1586 1172
rect 1646 1168 1650 1172
rect 1542 1158 1546 1162
rect 1398 1108 1402 1112
rect 1366 1048 1370 1052
rect 1350 1038 1354 1042
rect 1422 1118 1426 1122
rect 1422 1048 1426 1052
rect 1438 1048 1442 1052
rect 1406 1038 1410 1042
rect 1350 958 1354 962
rect 1390 948 1394 952
rect 1422 948 1426 952
rect 1454 948 1458 952
rect 1342 938 1346 942
rect 1390 938 1394 942
rect 1398 938 1402 942
rect 1414 938 1418 942
rect 1326 908 1330 912
rect 1326 898 1330 902
rect 1286 858 1290 862
rect 1318 858 1322 862
rect 1310 768 1314 772
rect 1278 758 1282 762
rect 1222 748 1226 752
rect 1294 748 1298 752
rect 1230 718 1234 722
rect 1246 728 1250 732
rect 1238 688 1242 692
rect 1222 668 1226 672
rect 1254 668 1258 672
rect 1206 608 1210 612
rect 1150 588 1154 592
rect 1150 578 1154 582
rect 1134 508 1138 512
rect 1142 498 1146 502
rect 1126 488 1130 492
rect 1070 468 1074 472
rect 1038 458 1042 462
rect 1046 458 1050 462
rect 1078 458 1082 462
rect 1110 438 1114 442
rect 982 378 986 382
rect 1110 378 1114 382
rect 1102 368 1106 372
rect 1078 358 1082 362
rect 974 348 978 352
rect 1054 348 1058 352
rect 966 338 970 342
rect 1086 348 1090 352
rect 1134 358 1138 362
rect 1046 338 1050 342
rect 1054 328 1058 332
rect 1118 328 1122 332
rect 966 318 970 322
rect 1014 318 1018 322
rect 986 303 990 307
rect 993 303 997 307
rect 974 288 978 292
rect 998 268 1002 272
rect 1030 268 1034 272
rect 958 258 962 262
rect 950 208 954 212
rect 886 198 890 202
rect 902 178 906 182
rect 998 158 1002 162
rect 1030 158 1034 162
rect 830 138 834 142
rect 1022 138 1026 142
rect 1006 128 1010 132
rect 1062 288 1066 292
rect 1110 278 1114 282
rect 1142 288 1146 292
rect 1086 268 1090 272
rect 1102 268 1106 272
rect 1078 258 1082 262
rect 1102 258 1106 262
rect 1078 228 1082 232
rect 1070 178 1074 182
rect 1086 168 1090 172
rect 1094 158 1098 162
rect 1086 148 1090 152
rect 910 118 914 122
rect 1006 118 1010 122
rect 1038 118 1042 122
rect 814 88 818 92
rect 870 88 874 92
rect 734 78 738 82
rect 758 68 762 72
rect 846 68 850 72
rect 862 68 866 72
rect 678 58 682 62
rect 694 58 698 62
rect 870 58 874 62
rect 846 48 850 52
rect 862 48 866 52
rect 986 103 990 107
rect 993 103 997 107
rect 894 78 898 82
rect 958 78 962 82
rect 1070 88 1074 92
rect 1078 78 1082 82
rect 1206 568 1210 572
rect 1174 558 1178 562
rect 1182 558 1186 562
rect 1182 528 1186 532
rect 1206 528 1210 532
rect 1198 518 1202 522
rect 1190 508 1194 512
rect 1182 468 1186 472
rect 1198 458 1202 462
rect 1358 888 1362 892
rect 1342 868 1346 872
rect 1350 848 1354 852
rect 1334 758 1338 762
rect 1318 748 1322 752
rect 1342 748 1346 752
rect 1294 728 1298 732
rect 1278 718 1282 722
rect 1294 708 1298 712
rect 1326 708 1330 712
rect 1286 688 1290 692
rect 1302 668 1306 672
rect 1334 678 1338 682
rect 1374 788 1378 792
rect 1366 778 1370 782
rect 1366 758 1370 762
rect 1406 868 1410 872
rect 1406 838 1410 842
rect 1430 928 1434 932
rect 1430 898 1434 902
rect 1446 858 1450 862
rect 1422 798 1426 802
rect 1438 778 1442 782
rect 1430 758 1434 762
rect 1390 748 1394 752
rect 1406 748 1410 752
rect 1414 708 1418 712
rect 1422 708 1426 712
rect 1438 698 1442 702
rect 1358 668 1362 672
rect 1374 668 1378 672
rect 1302 658 1306 662
rect 1326 658 1330 662
rect 1358 658 1362 662
rect 1230 638 1234 642
rect 1270 638 1274 642
rect 1254 598 1258 602
rect 1294 628 1298 632
rect 1294 598 1298 602
rect 1430 658 1434 662
rect 1398 638 1402 642
rect 1430 638 1434 642
rect 1390 608 1394 612
rect 1374 588 1378 592
rect 1334 558 1338 562
rect 1286 548 1290 552
rect 1406 548 1410 552
rect 1294 538 1298 542
rect 1238 528 1242 532
rect 1222 478 1226 482
rect 1278 478 1282 482
rect 1214 468 1218 472
rect 1222 458 1226 462
rect 1206 448 1210 452
rect 1206 418 1210 422
rect 1190 368 1194 372
rect 1222 398 1226 402
rect 1214 368 1218 372
rect 1286 368 1290 372
rect 1302 508 1306 512
rect 1422 538 1426 542
rect 1358 508 1362 512
rect 1406 508 1410 512
rect 1382 498 1386 502
rect 1302 468 1306 472
rect 1382 468 1386 472
rect 1342 438 1346 442
rect 1342 378 1346 382
rect 1310 368 1314 372
rect 1302 348 1306 352
rect 1134 258 1138 262
rect 1150 258 1154 262
rect 1118 188 1122 192
rect 1422 448 1426 452
rect 1390 438 1394 442
rect 1414 388 1418 392
rect 1398 368 1402 372
rect 1478 1138 1482 1142
rect 1494 1118 1498 1122
rect 1534 1118 1538 1122
rect 1486 1108 1490 1112
rect 1470 1028 1474 1032
rect 1498 1003 1502 1007
rect 1505 1003 1509 1007
rect 1502 948 1506 952
rect 1462 918 1466 922
rect 1470 908 1474 912
rect 1462 898 1466 902
rect 1566 1148 1570 1152
rect 1622 1148 1626 1152
rect 1550 1118 1554 1122
rect 1574 1118 1578 1122
rect 1558 1048 1562 1052
rect 1550 1008 1554 1012
rect 1598 1138 1602 1142
rect 1614 1118 1618 1122
rect 1646 1118 1650 1122
rect 1638 1098 1642 1102
rect 1662 1238 1666 1242
rect 1686 1238 1690 1242
rect 1670 1118 1674 1122
rect 1654 1108 1658 1112
rect 1590 1048 1594 1052
rect 1574 1038 1578 1042
rect 1566 1028 1570 1032
rect 1598 1008 1602 1012
rect 1566 968 1570 972
rect 1574 958 1578 962
rect 1558 938 1562 942
rect 1486 878 1490 882
rect 1518 878 1522 882
rect 1502 868 1506 872
rect 1462 859 1466 863
rect 1498 803 1502 807
rect 1505 803 1509 807
rect 1486 768 1490 772
rect 1454 758 1458 762
rect 1534 858 1538 862
rect 1526 848 1530 852
rect 1558 848 1562 852
rect 1590 908 1594 912
rect 1582 888 1586 892
rect 1598 888 1602 892
rect 1590 878 1594 882
rect 1582 858 1586 862
rect 1622 1048 1626 1052
rect 1766 1358 1770 1362
rect 1742 1348 1746 1352
rect 1758 1338 1762 1342
rect 1750 1298 1754 1302
rect 1750 1288 1754 1292
rect 1742 1278 1746 1282
rect 1870 1698 1874 1702
rect 1870 1678 1874 1682
rect 1870 1648 1874 1652
rect 1894 1578 1898 1582
rect 1878 1548 1882 1552
rect 1918 1928 1922 1932
rect 1942 1918 1946 1922
rect 1974 1918 1978 1922
rect 2006 1938 2010 1942
rect 2094 2218 2098 2222
rect 2462 2348 2466 2352
rect 2494 2348 2498 2352
rect 2142 2338 2146 2342
rect 2214 2338 2218 2342
rect 2254 2328 2258 2332
rect 2462 2328 2466 2332
rect 2206 2318 2210 2322
rect 2190 2278 2194 2282
rect 2150 2258 2154 2262
rect 2142 2248 2146 2252
rect 2158 2248 2162 2252
rect 2142 2218 2146 2222
rect 2134 2208 2138 2212
rect 2166 2218 2170 2222
rect 2158 2198 2162 2202
rect 2102 2178 2106 2182
rect 2174 2168 2178 2172
rect 2174 2148 2178 2152
rect 2158 2138 2162 2142
rect 2086 2048 2090 2052
rect 2054 2038 2058 2042
rect 2118 2058 2122 2062
rect 2134 2058 2138 2062
rect 2094 1968 2098 1972
rect 2078 1958 2082 1962
rect 2086 1958 2090 1962
rect 2038 1918 2042 1922
rect 2018 1903 2022 1907
rect 2025 1903 2029 1907
rect 1998 1888 2002 1892
rect 2030 1888 2034 1892
rect 1958 1868 1962 1872
rect 2070 1868 2074 1872
rect 2142 1958 2146 1962
rect 2086 1938 2090 1942
rect 2134 1938 2138 1942
rect 1982 1858 1986 1862
rect 1998 1858 2002 1862
rect 1998 1838 2002 1842
rect 1990 1808 1994 1812
rect 2062 1758 2066 1762
rect 1918 1748 1922 1752
rect 2038 1748 2042 1752
rect 1982 1738 1986 1742
rect 1926 1698 1930 1702
rect 1950 1698 1954 1702
rect 1926 1678 1930 1682
rect 2038 1738 2042 1742
rect 2062 1738 2066 1742
rect 2018 1703 2022 1707
rect 2025 1703 2029 1707
rect 1926 1658 1930 1662
rect 1958 1658 1962 1662
rect 1982 1608 1986 1612
rect 1982 1598 1986 1602
rect 1926 1558 1930 1562
rect 1958 1558 1962 1562
rect 1942 1548 1946 1552
rect 1966 1548 1970 1552
rect 1910 1538 1914 1542
rect 1862 1508 1866 1512
rect 1902 1508 1906 1512
rect 1798 1468 1802 1472
rect 1790 1458 1794 1462
rect 1846 1418 1850 1422
rect 1838 1408 1842 1412
rect 1822 1358 1826 1362
rect 1846 1368 1850 1372
rect 1798 1348 1802 1352
rect 1894 1348 1898 1352
rect 1830 1328 1834 1332
rect 1806 1318 1810 1322
rect 1846 1308 1850 1312
rect 1862 1308 1866 1312
rect 1838 1288 1842 1292
rect 1862 1288 1866 1292
rect 1734 1268 1738 1272
rect 1726 1248 1730 1252
rect 1782 1248 1786 1252
rect 1782 1238 1786 1242
rect 1710 1228 1714 1232
rect 1734 1228 1738 1232
rect 1854 1248 1858 1252
rect 1814 1218 1818 1222
rect 1830 1218 1834 1222
rect 1726 1168 1730 1172
rect 1734 1168 1738 1172
rect 1718 1158 1722 1162
rect 1702 1138 1706 1142
rect 1718 1138 1722 1142
rect 1710 1118 1714 1122
rect 1710 1098 1714 1102
rect 1694 1048 1698 1052
rect 1710 1048 1714 1052
rect 1726 1048 1730 1052
rect 1654 1038 1658 1042
rect 1670 1038 1674 1042
rect 1718 1028 1722 1032
rect 1702 998 1706 1002
rect 1750 1158 1754 1162
rect 1774 1158 1778 1162
rect 1758 1148 1762 1152
rect 1822 1148 1826 1152
rect 1758 1118 1762 1122
rect 1742 1108 1746 1112
rect 1734 988 1738 992
rect 1734 958 1738 962
rect 1662 898 1666 902
rect 1646 888 1650 892
rect 1654 888 1658 892
rect 1638 868 1642 872
rect 1654 868 1658 872
rect 1614 848 1618 852
rect 1638 828 1642 832
rect 1630 808 1634 812
rect 1566 798 1570 802
rect 1590 788 1594 792
rect 1582 768 1586 772
rect 1534 747 1538 751
rect 1702 888 1706 892
rect 1686 868 1690 872
rect 1702 868 1706 872
rect 1702 858 1706 862
rect 1710 858 1714 862
rect 1670 848 1674 852
rect 1694 848 1698 852
rect 1814 1118 1818 1122
rect 1822 1108 1826 1112
rect 1774 1048 1778 1052
rect 1814 1028 1818 1032
rect 1766 1018 1770 1022
rect 1814 998 1818 1002
rect 1798 988 1802 992
rect 1750 948 1754 952
rect 1798 928 1802 932
rect 1774 908 1778 912
rect 1758 858 1762 862
rect 1742 788 1746 792
rect 1670 778 1674 782
rect 1702 778 1706 782
rect 1646 768 1650 772
rect 1662 768 1666 772
rect 1694 768 1698 772
rect 1654 758 1658 762
rect 1678 758 1682 762
rect 1606 748 1610 752
rect 1622 748 1626 752
rect 1614 738 1618 742
rect 1446 668 1450 672
rect 1438 538 1442 542
rect 1462 608 1466 612
rect 1454 538 1458 542
rect 1462 528 1466 532
rect 1462 408 1466 412
rect 1438 388 1442 392
rect 1366 338 1370 342
rect 1414 338 1418 342
rect 1278 318 1282 322
rect 1262 288 1266 292
rect 1318 288 1322 292
rect 1198 278 1202 282
rect 1270 268 1274 272
rect 1278 268 1282 272
rect 1294 268 1298 272
rect 1350 268 1354 272
rect 1166 238 1170 242
rect 1134 168 1138 172
rect 1126 158 1130 162
rect 1190 148 1194 152
rect 1254 238 1258 242
rect 1262 218 1266 222
rect 1118 138 1122 142
rect 1126 138 1130 142
rect 1238 138 1242 142
rect 1246 128 1250 132
rect 1206 118 1210 122
rect 1222 118 1226 122
rect 1198 108 1202 112
rect 1302 258 1306 262
rect 1286 178 1290 182
rect 1294 168 1298 172
rect 1278 128 1282 132
rect 1326 118 1330 122
rect 1286 98 1290 102
rect 1270 88 1274 92
rect 1110 68 1114 72
rect 1182 68 1186 72
rect 1270 68 1274 72
rect 966 59 970 63
rect 1038 58 1042 62
rect 1070 58 1074 62
rect 1046 48 1050 52
rect 1062 48 1066 52
rect 1294 88 1298 92
rect 1430 328 1434 332
rect 1406 298 1410 302
rect 1406 288 1410 292
rect 1422 268 1426 272
rect 1574 718 1578 722
rect 1518 678 1522 682
rect 1558 668 1562 672
rect 1534 648 1538 652
rect 1486 608 1490 612
rect 1534 608 1538 612
rect 1498 603 1502 607
rect 1505 603 1509 607
rect 1742 758 1746 762
rect 1710 748 1714 752
rect 1670 738 1674 742
rect 1702 738 1706 742
rect 1654 728 1658 732
rect 1598 698 1602 702
rect 1654 708 1658 712
rect 1622 668 1626 672
rect 1670 708 1674 712
rect 1806 868 1810 872
rect 1790 768 1794 772
rect 1774 718 1778 722
rect 1726 688 1730 692
rect 1742 688 1746 692
rect 1678 678 1682 682
rect 1694 678 1698 682
rect 1726 678 1730 682
rect 1702 668 1706 672
rect 1734 668 1738 672
rect 1630 648 1634 652
rect 1646 648 1650 652
rect 1678 648 1682 652
rect 1614 638 1618 642
rect 1614 598 1618 602
rect 1590 578 1594 582
rect 1534 568 1538 572
rect 1558 568 1562 572
rect 1606 558 1610 562
rect 1526 548 1530 552
rect 1550 548 1554 552
rect 1494 538 1498 542
rect 1502 538 1506 542
rect 1526 518 1530 522
rect 1558 498 1562 502
rect 1518 478 1522 482
rect 1566 488 1570 492
rect 1542 468 1546 472
rect 1558 458 1562 462
rect 1550 418 1554 422
rect 1498 403 1502 407
rect 1505 403 1509 407
rect 1558 378 1562 382
rect 1470 358 1474 362
rect 1486 358 1490 362
rect 1454 338 1458 342
rect 1470 338 1474 342
rect 1454 318 1458 322
rect 1398 248 1402 252
rect 1382 168 1386 172
rect 1438 238 1442 242
rect 1390 158 1394 162
rect 1414 158 1418 162
rect 1430 158 1434 162
rect 1398 148 1402 152
rect 1342 138 1346 142
rect 1406 138 1410 142
rect 1334 108 1338 112
rect 1366 108 1370 112
rect 1390 98 1394 102
rect 1334 68 1338 72
rect 1406 68 1410 72
rect 1430 148 1434 152
rect 1478 308 1482 312
rect 1534 308 1538 312
rect 1518 298 1522 302
rect 1462 268 1466 272
rect 1510 268 1514 272
rect 1550 268 1554 272
rect 1582 518 1586 522
rect 1590 488 1594 492
rect 1574 478 1578 482
rect 1590 468 1594 472
rect 1598 468 1602 472
rect 1574 458 1578 462
rect 1574 338 1578 342
rect 1566 258 1570 262
rect 1462 188 1466 192
rect 1462 158 1466 162
rect 1430 138 1434 142
rect 1446 138 1450 142
rect 1498 203 1502 207
rect 1505 203 1509 207
rect 1518 148 1522 152
rect 1446 118 1450 122
rect 1454 98 1458 102
rect 1430 88 1434 92
rect 1430 78 1434 82
rect 1438 68 1442 72
rect 1142 58 1146 62
rect 1158 58 1162 62
rect 1262 58 1266 62
rect 1286 58 1290 62
rect 1398 58 1402 62
rect 1494 128 1498 132
rect 1542 228 1546 232
rect 1566 198 1570 202
rect 1550 148 1554 152
rect 1566 148 1570 152
rect 1526 98 1530 102
rect 1550 138 1554 142
rect 1534 88 1538 92
rect 1606 458 1610 462
rect 1630 488 1634 492
rect 1686 508 1690 512
rect 1678 498 1682 502
rect 1670 478 1674 482
rect 1646 458 1650 462
rect 1686 458 1690 462
rect 1702 448 1706 452
rect 1654 438 1658 442
rect 1694 428 1698 432
rect 1662 358 1666 362
rect 1654 348 1658 352
rect 1622 338 1626 342
rect 1614 298 1618 302
rect 1590 288 1594 292
rect 1646 288 1650 292
rect 1590 268 1594 272
rect 1638 268 1642 272
rect 1886 1328 1890 1332
rect 1886 1298 1890 1302
rect 1894 1268 1898 1272
rect 1950 1488 1954 1492
rect 1926 1478 1930 1482
rect 1910 1458 1914 1462
rect 1934 1408 1938 1412
rect 1926 1398 1930 1402
rect 1910 1368 1914 1372
rect 1910 1308 1914 1312
rect 1910 1278 1914 1282
rect 1942 1378 1946 1382
rect 1958 1358 1962 1362
rect 1942 1338 1946 1342
rect 1934 1288 1938 1292
rect 1950 1268 1954 1272
rect 1910 1258 1914 1262
rect 1838 1198 1842 1202
rect 1870 1198 1874 1202
rect 1870 1168 1874 1172
rect 1854 1158 1858 1162
rect 1878 1158 1882 1162
rect 1902 1178 1906 1182
rect 1878 1088 1882 1092
rect 1894 1098 1898 1102
rect 1886 1018 1890 1022
rect 1846 988 1850 992
rect 1878 958 1882 962
rect 1830 948 1834 952
rect 1862 938 1866 942
rect 1838 928 1842 932
rect 1894 928 1898 932
rect 1854 918 1858 922
rect 1886 878 1890 882
rect 1910 1168 1914 1172
rect 1910 1138 1914 1142
rect 1910 978 1914 982
rect 1910 948 1914 952
rect 1902 868 1906 872
rect 1918 868 1922 872
rect 1894 858 1898 862
rect 1822 848 1826 852
rect 1830 788 1834 792
rect 1862 848 1866 852
rect 1910 848 1914 852
rect 1894 838 1898 842
rect 1846 758 1850 762
rect 1878 758 1882 762
rect 1838 748 1842 752
rect 1878 748 1882 752
rect 1806 738 1810 742
rect 1814 718 1818 722
rect 1838 718 1842 722
rect 1886 738 1890 742
rect 1902 738 1906 742
rect 1910 708 1914 712
rect 1854 698 1858 702
rect 1862 688 1866 692
rect 1886 678 1890 682
rect 1958 1168 1962 1172
rect 1934 1148 1938 1152
rect 1958 1148 1962 1152
rect 2014 1588 2018 1592
rect 2022 1558 2026 1562
rect 1990 1518 1994 1522
rect 2030 1518 2034 1522
rect 2018 1503 2022 1507
rect 2025 1503 2029 1507
rect 1990 1468 1994 1472
rect 2030 1468 2034 1472
rect 2134 1918 2138 1922
rect 2118 1898 2122 1902
rect 2190 2118 2194 2122
rect 2214 2278 2218 2282
rect 2326 2318 2330 2322
rect 2406 2318 2410 2322
rect 2454 2318 2458 2322
rect 2222 2268 2226 2272
rect 2238 2268 2242 2272
rect 2302 2268 2306 2272
rect 2438 2268 2442 2272
rect 2246 2228 2250 2232
rect 2286 2258 2290 2262
rect 2358 2258 2362 2262
rect 2390 2258 2394 2262
rect 2262 2248 2266 2252
rect 2278 2248 2282 2252
rect 2254 2218 2258 2222
rect 2350 2218 2354 2222
rect 2238 2198 2242 2202
rect 2214 2168 2218 2172
rect 2206 2148 2210 2152
rect 2342 2188 2346 2192
rect 2254 2158 2258 2162
rect 2214 2138 2218 2142
rect 2310 2118 2314 2122
rect 2366 2158 2370 2162
rect 2350 2148 2354 2152
rect 2198 2098 2202 2102
rect 2262 2098 2266 2102
rect 2254 2088 2258 2092
rect 2238 2068 2242 2072
rect 2190 2058 2194 2062
rect 2182 1978 2186 1982
rect 2166 1958 2170 1962
rect 2182 1958 2186 1962
rect 2190 1948 2194 1952
rect 2158 1938 2162 1942
rect 2286 2088 2290 2092
rect 2302 2068 2306 2072
rect 2326 2068 2330 2072
rect 2206 2058 2210 2062
rect 2334 2058 2338 2062
rect 2222 1998 2226 2002
rect 2358 2098 2362 2102
rect 2414 2218 2418 2222
rect 2422 2218 2426 2222
rect 2398 2208 2402 2212
rect 2398 2158 2402 2162
rect 2406 2148 2410 2152
rect 2414 2138 2418 2142
rect 2406 2118 2410 2122
rect 2406 2088 2410 2092
rect 2470 2248 2474 2252
rect 2486 2188 2490 2192
rect 2454 2158 2458 2162
rect 2446 2118 2450 2122
rect 2422 2078 2426 2082
rect 2358 2058 2362 2062
rect 2310 2048 2314 2052
rect 2342 2048 2346 2052
rect 2246 1988 2250 1992
rect 2214 1978 2218 1982
rect 2198 1898 2202 1902
rect 2150 1858 2154 1862
rect 2174 1858 2178 1862
rect 2142 1828 2146 1832
rect 2150 1828 2154 1832
rect 2174 1808 2178 1812
rect 2118 1788 2122 1792
rect 2246 1968 2250 1972
rect 2222 1958 2226 1962
rect 2198 1758 2202 1762
rect 2078 1728 2082 1732
rect 2102 1738 2106 1742
rect 2094 1718 2098 1722
rect 2086 1708 2090 1712
rect 2054 1688 2058 1692
rect 2070 1678 2074 1682
rect 2310 1978 2314 1982
rect 2270 1958 2274 1962
rect 2262 1948 2266 1952
rect 2438 2008 2442 2012
rect 2430 1968 2434 1972
rect 2326 1958 2330 1962
rect 2446 1958 2450 1962
rect 2470 2138 2474 2142
rect 2462 2088 2466 2092
rect 2494 2098 2498 2102
rect 2486 2078 2490 2082
rect 2470 2048 2474 2052
rect 2470 2028 2474 2032
rect 2334 1948 2338 1952
rect 2382 1948 2386 1952
rect 2254 1938 2258 1942
rect 2334 1918 2338 1922
rect 2318 1908 2322 1912
rect 2334 1888 2338 1892
rect 2294 1878 2298 1882
rect 2334 1868 2338 1872
rect 2286 1858 2290 1862
rect 2246 1848 2250 1852
rect 2262 1848 2266 1852
rect 2278 1848 2282 1852
rect 2238 1808 2242 1812
rect 2302 1828 2306 1832
rect 2390 1828 2394 1832
rect 2262 1798 2266 1802
rect 2254 1758 2258 1762
rect 2326 1818 2330 1822
rect 2310 1808 2314 1812
rect 2150 1748 2154 1752
rect 2262 1738 2266 1742
rect 2214 1728 2218 1732
rect 2246 1728 2250 1732
rect 2118 1708 2122 1712
rect 2150 1678 2154 1682
rect 2062 1658 2066 1662
rect 2086 1658 2090 1662
rect 2094 1658 2098 1662
rect 2118 1658 2122 1662
rect 2134 1648 2138 1652
rect 2158 1648 2162 1652
rect 2046 1638 2050 1642
rect 2110 1638 2114 1642
rect 2046 1588 2050 1592
rect 2286 1728 2290 1732
rect 2270 1718 2274 1722
rect 2318 1688 2322 1692
rect 2214 1678 2218 1682
rect 2174 1658 2178 1662
rect 2182 1658 2186 1662
rect 2254 1658 2258 1662
rect 2166 1598 2170 1602
rect 2142 1588 2146 1592
rect 2070 1578 2074 1582
rect 2134 1578 2138 1582
rect 2062 1568 2066 1572
rect 2166 1568 2170 1572
rect 2206 1558 2210 1562
rect 2318 1568 2322 1572
rect 2094 1548 2098 1552
rect 2134 1548 2138 1552
rect 2230 1548 2234 1552
rect 2278 1548 2282 1552
rect 2334 1788 2338 1792
rect 2406 1788 2410 1792
rect 2374 1768 2378 1772
rect 2342 1758 2346 1762
rect 2350 1738 2354 1742
rect 2366 1708 2370 1712
rect 2390 1718 2394 1722
rect 2374 1698 2378 1702
rect 2350 1688 2354 1692
rect 2358 1688 2362 1692
rect 2406 1678 2410 1682
rect 2374 1668 2378 1672
rect 2366 1618 2370 1622
rect 2326 1558 2330 1562
rect 2342 1558 2346 1562
rect 2350 1548 2354 1552
rect 2254 1538 2258 1542
rect 2206 1488 2210 1492
rect 2230 1488 2234 1492
rect 2278 1488 2282 1492
rect 2062 1478 2066 1482
rect 2190 1478 2194 1482
rect 2070 1468 2074 1472
rect 2086 1468 2090 1472
rect 2014 1458 2018 1462
rect 2134 1458 2138 1462
rect 1974 1448 1978 1452
rect 1990 1448 1994 1452
rect 1974 1388 1978 1392
rect 2214 1468 2218 1472
rect 2230 1468 2234 1472
rect 2286 1468 2290 1472
rect 2246 1458 2250 1462
rect 2286 1458 2290 1462
rect 2302 1458 2306 1462
rect 2318 1458 2322 1462
rect 2046 1448 2050 1452
rect 2166 1448 2170 1452
rect 2190 1448 2194 1452
rect 2222 1448 2226 1452
rect 2278 1448 2282 1452
rect 2038 1428 2042 1432
rect 1974 1358 1978 1362
rect 1982 1348 1986 1352
rect 2018 1303 2022 1307
rect 2025 1303 2029 1307
rect 2014 1288 2018 1292
rect 1974 1278 1978 1282
rect 2022 1218 2026 1222
rect 2134 1408 2138 1412
rect 2158 1408 2162 1412
rect 2118 1368 2122 1372
rect 2102 1358 2106 1362
rect 2070 1348 2074 1352
rect 2166 1368 2170 1372
rect 2302 1358 2306 1362
rect 2142 1348 2146 1352
rect 2222 1348 2226 1352
rect 2150 1338 2154 1342
rect 2174 1338 2178 1342
rect 2062 1308 2066 1312
rect 1982 1208 1986 1212
rect 2038 1208 2042 1212
rect 2254 1308 2258 1312
rect 2166 1298 2170 1302
rect 2270 1298 2274 1302
rect 2102 1288 2106 1292
rect 2150 1288 2154 1292
rect 2070 1268 2074 1272
rect 2254 1288 2258 1292
rect 2182 1278 2186 1282
rect 2246 1268 2250 1272
rect 2262 1268 2266 1272
rect 2118 1258 2122 1262
rect 2198 1258 2202 1262
rect 2222 1258 2226 1262
rect 2262 1258 2266 1262
rect 2126 1248 2130 1252
rect 2142 1248 2146 1252
rect 2198 1248 2202 1252
rect 2318 1248 2322 1252
rect 2158 1238 2162 1242
rect 2246 1238 2250 1242
rect 2302 1208 2306 1212
rect 2246 1198 2250 1202
rect 2086 1168 2090 1172
rect 2102 1168 2106 1172
rect 2198 1168 2202 1172
rect 2126 1158 2130 1162
rect 2206 1148 2210 1152
rect 1958 1138 1962 1142
rect 2038 1138 2042 1142
rect 2198 1138 2202 1142
rect 1934 1128 1938 1132
rect 1974 1128 1978 1132
rect 1990 1118 1994 1122
rect 1974 1108 1978 1112
rect 2094 1108 2098 1112
rect 1942 1098 1946 1102
rect 2018 1103 2022 1107
rect 2025 1103 2029 1107
rect 2030 1088 2034 1092
rect 2254 1168 2258 1172
rect 2310 1158 2314 1162
rect 2382 1468 2386 1472
rect 2390 1468 2394 1472
rect 2342 1448 2346 1452
rect 2406 1458 2410 1462
rect 2398 1448 2402 1452
rect 2398 1438 2402 1442
rect 2382 1428 2386 1432
rect 2382 1358 2386 1362
rect 2334 1338 2338 1342
rect 2342 1308 2346 1312
rect 2358 1298 2362 1302
rect 2374 1338 2378 1342
rect 2382 1248 2386 1252
rect 2390 1248 2394 1252
rect 2350 1198 2354 1202
rect 2390 1188 2394 1192
rect 2382 1178 2386 1182
rect 2406 1428 2410 1432
rect 2430 1538 2434 1542
rect 2462 1928 2466 1932
rect 2470 1878 2474 1882
rect 2462 1868 2466 1872
rect 2486 2058 2490 2062
rect 2486 1978 2490 1982
rect 2502 1878 2506 1882
rect 2454 1818 2458 1822
rect 2478 1818 2482 1822
rect 2486 1768 2490 1772
rect 2446 1758 2450 1762
rect 2478 1748 2482 1752
rect 2502 1748 2506 1752
rect 2478 1728 2482 1732
rect 2494 1728 2498 1732
rect 2462 1708 2466 1712
rect 2486 1698 2490 1702
rect 2470 1688 2474 1692
rect 2446 1608 2450 1612
rect 2462 1578 2466 1582
rect 2494 1568 2498 1572
rect 2478 1548 2482 1552
rect 2438 1488 2442 1492
rect 2446 1468 2450 1472
rect 2414 1298 2418 1302
rect 2406 1278 2410 1282
rect 2406 1258 2410 1262
rect 2398 1168 2402 1172
rect 2382 1158 2386 1162
rect 2326 1148 2330 1152
rect 2342 1148 2346 1152
rect 2222 1138 2226 1142
rect 2190 1108 2194 1112
rect 2102 1068 2106 1072
rect 2150 1068 2154 1072
rect 2182 1068 2186 1072
rect 2238 1068 2242 1072
rect 2254 1068 2258 1072
rect 1998 1058 2002 1062
rect 2014 1058 2018 1062
rect 1934 978 1938 982
rect 1958 938 1962 942
rect 1982 908 1986 912
rect 1966 888 1970 892
rect 1942 868 1946 872
rect 1974 858 1978 862
rect 1926 848 1930 852
rect 1942 808 1946 812
rect 1974 808 1978 812
rect 1990 808 1994 812
rect 1934 778 1938 782
rect 1950 758 1954 762
rect 1974 748 1978 752
rect 2006 1038 2010 1042
rect 2078 1048 2082 1052
rect 2086 1038 2090 1042
rect 2054 1028 2058 1032
rect 2118 1058 2122 1062
rect 2198 1058 2202 1062
rect 2094 1018 2098 1022
rect 2078 1008 2082 1012
rect 2054 968 2058 972
rect 2046 958 2050 962
rect 2006 948 2010 952
rect 2038 918 2042 922
rect 2018 903 2022 907
rect 2025 903 2029 907
rect 2030 868 2034 872
rect 2022 848 2026 852
rect 2030 808 2034 812
rect 2014 788 2018 792
rect 2022 758 2026 762
rect 2110 1048 2114 1052
rect 2150 1048 2154 1052
rect 2110 1028 2114 1032
rect 2102 998 2106 1002
rect 2142 998 2146 1002
rect 2102 988 2106 992
rect 2158 1018 2162 1022
rect 2206 1018 2210 1022
rect 2214 1008 2218 1012
rect 2206 958 2210 962
rect 2134 948 2138 952
rect 2158 948 2162 952
rect 2062 938 2066 942
rect 2086 908 2090 912
rect 2078 888 2082 892
rect 2054 868 2058 872
rect 2046 858 2050 862
rect 2046 748 2050 752
rect 1934 728 1938 732
rect 1998 728 2002 732
rect 1990 718 1994 722
rect 1926 678 1930 682
rect 1934 668 1938 672
rect 1990 668 1994 672
rect 2014 738 2018 742
rect 2046 738 2050 742
rect 2018 703 2022 707
rect 2025 703 2029 707
rect 2022 688 2026 692
rect 2038 678 2042 682
rect 2086 868 2090 872
rect 2126 878 2130 882
rect 2142 868 2146 872
rect 2174 868 2178 872
rect 2198 868 2202 872
rect 2246 1038 2250 1042
rect 2286 1138 2290 1142
rect 2270 1088 2274 1092
rect 2286 1088 2290 1092
rect 2278 1068 2282 1072
rect 2270 1038 2274 1042
rect 2262 1028 2266 1032
rect 2270 958 2274 962
rect 2294 1048 2298 1052
rect 2318 1138 2322 1142
rect 2318 1058 2322 1062
rect 2310 1048 2314 1052
rect 2302 1008 2306 1012
rect 2438 1308 2442 1312
rect 2478 1498 2482 1502
rect 2502 1508 2506 1512
rect 2502 1478 2506 1482
rect 2486 1318 2490 1322
rect 2470 1288 2474 1292
rect 2454 1268 2458 1272
rect 2446 1258 2450 1262
rect 2430 1228 2434 1232
rect 2454 1228 2458 1232
rect 2422 1198 2426 1202
rect 2430 1158 2434 1162
rect 2414 1148 2418 1152
rect 2374 1138 2378 1142
rect 2374 1128 2378 1132
rect 2414 1128 2418 1132
rect 2414 1108 2418 1112
rect 2366 1088 2370 1092
rect 2438 1088 2442 1092
rect 2446 1078 2450 1082
rect 2390 1068 2394 1072
rect 2358 1058 2362 1062
rect 2406 1058 2410 1062
rect 2438 1058 2442 1062
rect 2446 1058 2450 1062
rect 2318 958 2322 962
rect 2222 948 2226 952
rect 2310 948 2314 952
rect 2230 938 2234 942
rect 2262 938 2266 942
rect 2222 918 2226 922
rect 2262 888 2266 892
rect 2190 858 2194 862
rect 2214 858 2218 862
rect 2278 858 2282 862
rect 2102 848 2106 852
rect 2094 838 2098 842
rect 2102 838 2106 842
rect 2070 758 2074 762
rect 2030 668 2034 672
rect 1870 658 1874 662
rect 1942 658 1946 662
rect 1838 648 1842 652
rect 1910 648 1914 652
rect 1998 648 2002 652
rect 1886 588 1890 592
rect 1902 588 1906 592
rect 1758 578 1762 582
rect 2062 658 2066 662
rect 2046 588 2050 592
rect 1894 558 1898 562
rect 2030 558 2034 562
rect 2086 718 2090 722
rect 2094 698 2098 702
rect 2094 678 2098 682
rect 2078 578 2082 582
rect 2054 568 2058 572
rect 1982 548 1986 552
rect 2014 548 2018 552
rect 1758 538 1762 542
rect 1822 538 1826 542
rect 1870 538 1874 542
rect 1878 538 1882 542
rect 1902 538 1906 542
rect 1734 518 1738 522
rect 1798 478 1802 482
rect 1926 538 1930 542
rect 1958 538 1962 542
rect 1902 528 1906 532
rect 1870 518 1874 522
rect 1918 518 1922 522
rect 1974 538 1978 542
rect 1966 518 1970 522
rect 1966 508 1970 512
rect 1814 468 1818 472
rect 1958 468 1962 472
rect 1990 468 1994 472
rect 1742 458 1746 462
rect 1790 458 1794 462
rect 1870 458 1874 462
rect 2018 503 2022 507
rect 2025 503 2029 507
rect 2046 508 2050 512
rect 2038 478 2042 482
rect 2006 458 2010 462
rect 2030 458 2034 462
rect 1670 348 1674 352
rect 1686 338 1690 342
rect 1702 338 1706 342
rect 1718 338 1722 342
rect 1694 328 1698 332
rect 1670 318 1674 322
rect 1710 318 1714 322
rect 1670 298 1674 302
rect 1670 278 1674 282
rect 1694 278 1698 282
rect 1614 258 1618 262
rect 1630 258 1634 262
rect 1646 258 1650 262
rect 1662 258 1666 262
rect 1694 258 1698 262
rect 1654 238 1658 242
rect 1598 178 1602 182
rect 1630 178 1634 182
rect 1582 168 1586 172
rect 1598 168 1602 172
rect 1582 148 1586 152
rect 1646 168 1650 172
rect 1598 78 1602 82
rect 1638 108 1642 112
rect 1614 68 1618 72
rect 1702 208 1706 212
rect 1798 448 1802 452
rect 1886 448 1890 452
rect 1782 428 1786 432
rect 1862 388 1866 392
rect 1822 368 1826 372
rect 1870 368 1874 372
rect 1766 348 1770 352
rect 1726 228 1730 232
rect 1718 188 1722 192
rect 1774 338 1778 342
rect 1758 308 1762 312
rect 1870 358 1874 362
rect 1838 348 1842 352
rect 1854 348 1858 352
rect 1782 288 1786 292
rect 1814 288 1818 292
rect 1774 278 1778 282
rect 1742 208 1746 212
rect 1734 188 1738 192
rect 1726 178 1730 182
rect 1750 188 1754 192
rect 1726 148 1730 152
rect 1694 138 1698 142
rect 1710 138 1714 142
rect 1742 138 1746 142
rect 1678 88 1682 92
rect 1694 88 1698 92
rect 1830 258 1834 262
rect 1822 248 1826 252
rect 1862 318 1866 322
rect 1878 288 1882 292
rect 1862 278 1866 282
rect 1846 258 1850 262
rect 1862 248 1866 252
rect 1838 218 1842 222
rect 1918 388 1922 392
rect 1934 358 1938 362
rect 1910 228 1914 232
rect 1862 158 1866 162
rect 1878 158 1882 162
rect 1798 148 1802 152
rect 1838 148 1842 152
rect 1862 138 1866 142
rect 1814 88 1818 92
rect 1878 118 1882 122
rect 1782 78 1786 82
rect 1902 168 1906 172
rect 1990 448 1994 452
rect 1974 378 1978 382
rect 1966 308 1970 312
rect 2022 318 2026 322
rect 2018 303 2022 307
rect 2025 303 2029 307
rect 1934 258 1938 262
rect 2006 258 2010 262
rect 1926 248 1930 252
rect 1918 148 1922 152
rect 1974 248 1978 252
rect 1990 168 1994 172
rect 2070 488 2074 492
rect 2094 488 2098 492
rect 2078 468 2082 472
rect 2078 438 2082 442
rect 2070 388 2074 392
rect 2046 328 2050 332
rect 2054 318 2058 322
rect 2142 808 2146 812
rect 2126 798 2130 802
rect 2110 778 2114 782
rect 2198 848 2202 852
rect 2198 818 2202 822
rect 2150 778 2154 782
rect 2166 768 2170 772
rect 2158 758 2162 762
rect 2190 758 2194 762
rect 2118 738 2122 742
rect 2110 718 2114 722
rect 2126 698 2130 702
rect 2118 668 2122 672
rect 2134 668 2138 672
rect 2134 628 2138 632
rect 2150 748 2154 752
rect 2174 718 2178 722
rect 2158 698 2162 702
rect 2150 668 2154 672
rect 2150 638 2154 642
rect 2134 548 2138 552
rect 2182 538 2186 542
rect 2150 508 2154 512
rect 2182 488 2186 492
rect 2118 468 2122 472
rect 2142 459 2146 463
rect 2134 368 2138 372
rect 2118 278 2122 282
rect 2078 268 2082 272
rect 2102 268 2106 272
rect 2126 268 2130 272
rect 2054 258 2058 262
rect 1950 138 1954 142
rect 1942 128 1946 132
rect 1934 88 1938 92
rect 1894 78 1898 82
rect 2006 128 2010 132
rect 2094 258 2098 262
rect 2150 348 2154 352
rect 2174 348 2178 352
rect 2158 338 2162 342
rect 2062 178 2066 182
rect 2198 728 2202 732
rect 2206 688 2210 692
rect 2206 668 2210 672
rect 2326 948 2330 952
rect 2374 958 2378 962
rect 2342 918 2346 922
rect 2294 908 2298 912
rect 2310 908 2314 912
rect 2302 898 2306 902
rect 2326 878 2330 882
rect 2302 858 2306 862
rect 2286 848 2290 852
rect 2302 838 2306 842
rect 2342 848 2346 852
rect 2246 828 2250 832
rect 2302 778 2306 782
rect 2254 748 2258 752
rect 2294 738 2298 742
rect 2262 688 2266 692
rect 2238 678 2242 682
rect 2254 678 2258 682
rect 2294 678 2298 682
rect 2422 958 2426 962
rect 2438 958 2442 962
rect 2406 898 2410 902
rect 2398 888 2402 892
rect 2414 878 2418 882
rect 2430 918 2434 922
rect 2430 858 2434 862
rect 2486 1178 2490 1182
rect 2494 1088 2498 1092
rect 2486 1028 2490 1032
rect 2518 2008 2522 2012
rect 2462 948 2466 952
rect 2470 938 2474 942
rect 2478 938 2482 942
rect 2510 888 2514 892
rect 2470 878 2474 882
rect 2502 868 2506 872
rect 2486 758 2490 762
rect 2446 748 2450 752
rect 2462 748 2466 752
rect 2422 738 2426 742
rect 2470 738 2474 742
rect 2494 738 2498 742
rect 2334 688 2338 692
rect 2318 678 2322 682
rect 2390 678 2394 682
rect 2358 668 2362 672
rect 2262 618 2266 622
rect 2214 598 2218 602
rect 2278 598 2282 602
rect 2294 648 2298 652
rect 2286 588 2290 592
rect 2286 578 2290 582
rect 2278 568 2282 572
rect 2214 538 2218 542
rect 2254 538 2258 542
rect 2270 538 2274 542
rect 2238 508 2242 512
rect 2206 478 2210 482
rect 2230 478 2234 482
rect 2198 458 2202 462
rect 2198 438 2202 442
rect 2158 268 2162 272
rect 2166 258 2170 262
rect 2150 248 2154 252
rect 2118 228 2122 232
rect 2102 158 2106 162
rect 2134 158 2138 162
rect 2046 148 2050 152
rect 2150 148 2154 152
rect 2182 148 2186 152
rect 2078 138 2082 142
rect 2054 128 2058 132
rect 2038 108 2042 112
rect 2018 103 2022 107
rect 2025 103 2029 107
rect 2054 98 2058 102
rect 2270 478 2274 482
rect 2278 468 2282 472
rect 2262 448 2266 452
rect 2222 438 2226 442
rect 2238 368 2242 372
rect 2214 358 2218 362
rect 2262 288 2266 292
rect 2422 688 2426 692
rect 2454 678 2458 682
rect 2454 668 2458 672
rect 2302 598 2306 602
rect 2462 618 2466 622
rect 2318 608 2322 612
rect 2390 608 2394 612
rect 2326 568 2330 572
rect 2374 568 2378 572
rect 2310 558 2314 562
rect 2318 548 2322 552
rect 2294 368 2298 372
rect 2398 588 2402 592
rect 2510 698 2514 702
rect 2334 548 2338 552
rect 2374 548 2378 552
rect 2358 538 2362 542
rect 2406 538 2410 542
rect 2342 518 2346 522
rect 2406 488 2410 492
rect 2382 468 2386 472
rect 2438 468 2442 472
rect 2334 458 2338 462
rect 2374 458 2378 462
rect 2390 458 2394 462
rect 2414 368 2418 372
rect 2374 358 2378 362
rect 2406 358 2410 362
rect 2398 348 2402 352
rect 2326 338 2330 342
rect 2342 338 2346 342
rect 2366 338 2370 342
rect 2294 288 2298 292
rect 2310 288 2314 292
rect 2230 268 2234 272
rect 2390 288 2394 292
rect 2358 268 2362 272
rect 2342 258 2346 262
rect 2214 198 2218 202
rect 2142 138 2146 142
rect 2214 138 2218 142
rect 2110 128 2114 132
rect 2110 98 2114 102
rect 2094 88 2098 92
rect 2062 78 2066 82
rect 2158 78 2162 82
rect 1670 68 1674 72
rect 1758 68 1762 72
rect 1806 68 1810 72
rect 1838 68 1842 72
rect 1974 68 1978 72
rect 2046 68 2050 72
rect 1470 58 1474 62
rect 1526 58 1530 62
rect 1558 58 1562 62
rect 1574 58 1578 62
rect 1654 58 1658 62
rect 1694 58 1698 62
rect 2238 248 2242 252
rect 2294 238 2298 242
rect 2238 198 2242 202
rect 2446 358 2450 362
rect 2430 328 2434 332
rect 2494 488 2498 492
rect 2518 438 2522 442
rect 2502 368 2506 372
rect 2510 358 2514 362
rect 2502 298 2506 302
rect 2494 278 2498 282
rect 2446 258 2450 262
rect 2518 298 2522 302
rect 2518 278 2522 282
rect 2518 258 2522 262
rect 2518 238 2522 242
rect 2254 158 2258 162
rect 2406 158 2410 162
rect 2494 158 2498 162
rect 2238 148 2242 152
rect 2310 148 2314 152
rect 2342 148 2346 152
rect 2358 148 2362 152
rect 2366 138 2370 142
rect 2486 138 2490 142
rect 2270 128 2274 132
rect 2222 78 2226 82
rect 2350 78 2354 82
rect 2438 88 2442 92
rect 2478 88 2482 92
rect 2238 68 2242 72
rect 2326 68 2330 72
rect 2422 68 2426 72
rect 2438 68 2442 72
rect 2518 68 2522 72
rect 2214 58 2218 62
rect 2246 58 2250 62
rect 1414 48 1418 52
rect 1806 48 1810 52
rect 1878 48 1882 52
rect 1838 38 1842 42
rect 2478 48 2482 52
rect 1110 28 1114 32
rect 1958 28 1962 32
rect 1982 28 1986 32
rect 1422 8 1426 12
rect 1654 8 1658 12
rect 2038 8 2042 12
rect 1498 3 1502 7
rect 1505 3 1509 7
<< metal3 >>
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 494 2403 496 2407
rect 1496 2403 1498 2407
rect 1502 2403 1505 2407
rect 1510 2403 1512 2407
rect 250 2398 262 2401
rect 922 2398 926 2401
rect 1146 2398 1158 2401
rect 1806 2392 1809 2398
rect 858 2378 1126 2381
rect 562 2368 574 2371
rect 742 2371 745 2378
rect 642 2368 745 2371
rect 1050 2368 1110 2371
rect 74 2358 86 2361
rect 298 2358 310 2361
rect 562 2358 590 2361
rect 594 2358 1102 2361
rect 1130 2358 1214 2361
rect 1290 2358 1302 2361
rect 1330 2358 1342 2361
rect 1918 2361 1921 2368
rect 1850 2358 1921 2361
rect 1994 2358 2086 2361
rect 2098 2358 2214 2361
rect 2218 2358 2382 2361
rect 2458 2358 2553 2361
rect 98 2348 166 2351
rect 194 2348 286 2351
rect 366 2351 369 2358
rect 2550 2352 2553 2358
rect 322 2348 369 2351
rect 514 2348 558 2351
rect 722 2348 750 2351
rect 754 2348 1278 2351
rect 1482 2348 1510 2351
rect 1570 2348 1574 2351
rect 1578 2348 1598 2351
rect 1834 2348 1910 2351
rect 1938 2348 2046 2351
rect 2074 2348 2094 2351
rect 2274 2348 2310 2351
rect 2362 2348 2366 2351
rect 2418 2348 2462 2351
rect 2466 2348 2494 2351
rect 2550 2348 2554 2352
rect 26 2338 46 2341
rect 50 2338 54 2341
rect 222 2338 278 2341
rect 458 2338 558 2341
rect 562 2338 582 2341
rect 598 2341 601 2348
rect 598 2338 758 2341
rect 762 2338 766 2341
rect 838 2338 910 2341
rect 978 2338 1009 2341
rect 1106 2338 1190 2341
rect 1202 2338 1286 2341
rect 1474 2338 1566 2341
rect 1594 2338 1678 2341
rect 1702 2341 1705 2348
rect 2238 2342 2241 2348
rect 1702 2338 1886 2341
rect 1890 2338 1990 2341
rect 1994 2338 2142 2341
rect 2210 2338 2214 2341
rect 2334 2341 2337 2348
rect 2306 2338 2337 2341
rect 222 2332 225 2338
rect 838 2332 841 2338
rect 1006 2332 1009 2338
rect 2462 2332 2465 2338
rect 66 2328 174 2331
rect 178 2328 222 2331
rect 290 2328 342 2331
rect 346 2328 366 2331
rect 538 2328 630 2331
rect 1010 2328 1174 2331
rect 1178 2328 1246 2331
rect 1786 2328 1990 2331
rect 2106 2328 2254 2331
rect 338 2318 422 2321
rect 426 2318 646 2321
rect 706 2318 918 2321
rect 978 2318 1190 2321
rect 1306 2318 1761 2321
rect 2058 2318 2206 2321
rect 2330 2318 2334 2321
rect 2394 2318 2406 2321
rect 2450 2318 2454 2321
rect 762 2308 766 2311
rect 810 2308 854 2311
rect 1090 2308 1230 2311
rect 1266 2308 1446 2311
rect 1490 2308 1750 2311
rect 1758 2311 1761 2318
rect 1758 2308 1814 2311
rect 1914 2308 1958 2311
rect 984 2303 986 2307
rect 990 2303 993 2307
rect 998 2303 1000 2307
rect 2016 2303 2018 2307
rect 2022 2303 2025 2307
rect 2030 2303 2032 2307
rect 826 2298 974 2301
rect 1346 2298 1358 2301
rect 1370 2298 1470 2301
rect 1474 2298 1502 2301
rect 1618 2298 1878 2301
rect 226 2288 310 2291
rect 314 2288 334 2291
rect 426 2288 510 2291
rect 514 2288 550 2291
rect 874 2288 1094 2291
rect 1098 2288 1150 2291
rect 1154 2288 1206 2291
rect 1210 2288 1318 2291
rect 1322 2288 1382 2291
rect 1538 2288 1822 2291
rect 1826 2288 1862 2291
rect 1906 2288 2041 2291
rect 2038 2282 2041 2288
rect 682 2278 758 2281
rect 762 2278 854 2281
rect 906 2278 910 2281
rect 946 2278 974 2281
rect 978 2278 1102 2281
rect 1274 2278 1286 2281
rect 1290 2278 1414 2281
rect 1426 2278 1622 2281
rect 1722 2278 1902 2281
rect 1906 2278 2014 2281
rect 2042 2278 2190 2281
rect 2218 2278 2358 2281
rect 114 2268 358 2271
rect 570 2268 622 2271
rect 914 2268 1006 2271
rect 1058 2268 1078 2271
rect 1198 2268 1222 2271
rect 1226 2268 1478 2271
rect 1546 2268 1550 2271
rect 1954 2268 2222 2271
rect 2242 2268 2302 2271
rect 194 2258 206 2261
rect 350 2258 390 2261
rect 410 2258 457 2261
rect 350 2252 353 2258
rect 454 2252 457 2258
rect 634 2258 742 2261
rect 790 2261 793 2268
rect 746 2258 793 2261
rect 818 2258 862 2261
rect 962 2258 1014 2261
rect 1030 2261 1033 2268
rect 1198 2262 1201 2268
rect 1030 2258 1086 2261
rect 1186 2258 1198 2261
rect 1250 2258 1382 2261
rect 1386 2258 1430 2261
rect 1434 2258 1446 2261
rect 1466 2258 1646 2261
rect 1830 2261 1833 2268
rect 1650 2258 1833 2261
rect 1926 2261 1929 2268
rect 1898 2258 1929 2261
rect 1970 2258 1974 2261
rect 1978 2258 1998 2261
rect 2154 2258 2158 2261
rect 2290 2258 2358 2261
rect 2438 2261 2441 2268
rect 2394 2258 2441 2261
rect 598 2252 601 2258
rect 202 2248 254 2251
rect 386 2248 414 2251
rect 418 2248 438 2251
rect 878 2251 881 2258
rect 2262 2252 2265 2258
rect 2470 2252 2473 2258
rect 866 2248 881 2251
rect 1082 2248 1102 2251
rect 1106 2248 1110 2251
rect 1114 2248 1326 2251
rect 1354 2248 1398 2251
rect 1410 2248 1582 2251
rect 1586 2248 1758 2251
rect 1834 2248 2046 2251
rect 2146 2248 2158 2251
rect 2266 2248 2278 2251
rect 2282 2248 2286 2251
rect 90 2238 166 2241
rect 170 2238 286 2241
rect 290 2238 374 2241
rect 594 2238 1054 2241
rect 1074 2238 1126 2241
rect 1170 2238 1366 2241
rect 1406 2241 1409 2248
rect 1822 2242 1825 2248
rect 1370 2238 1409 2241
rect 1490 2238 1606 2241
rect 1610 2238 1630 2241
rect 1858 2238 1974 2241
rect 2002 2238 2446 2241
rect 138 2228 870 2231
rect 906 2228 1206 2231
rect 1282 2228 1342 2231
rect 1562 2228 1830 2231
rect 2250 2228 2350 2231
rect 18 2218 254 2221
rect 330 2218 574 2221
rect 642 2218 894 2221
rect 1154 2218 1158 2221
rect 1194 2218 1214 2221
rect 1570 2218 1598 2221
rect 1602 2218 1782 2221
rect 1786 2218 1958 2221
rect 1962 2218 1990 2221
rect 2098 2218 2142 2221
rect 2146 2218 2166 2221
rect 2258 2218 2350 2221
rect 2418 2218 2422 2221
rect 74 2208 190 2211
rect 674 2208 686 2211
rect 1042 2208 1166 2211
rect 2138 2208 2398 2211
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 494 2203 496 2207
rect 1496 2203 1498 2207
rect 1502 2203 1505 2207
rect 1510 2203 1512 2207
rect 618 2198 638 2201
rect 666 2198 694 2201
rect 874 2198 910 2201
rect 914 2198 1062 2201
rect 2162 2198 2238 2201
rect 18 2188 150 2191
rect 154 2188 966 2191
rect 1602 2188 2118 2191
rect 2122 2188 2342 2191
rect 2458 2188 2486 2191
rect 1002 2178 1062 2181
rect 1250 2178 1366 2181
rect 1490 2178 1822 2181
rect 1906 2178 1918 2181
rect 1978 2178 2102 2181
rect 90 2168 110 2171
rect 114 2168 142 2171
rect 146 2168 166 2171
rect 346 2168 350 2171
rect 702 2171 705 2178
rect 658 2168 705 2171
rect 1010 2168 1630 2171
rect 1634 2168 1654 2171
rect 1658 2168 2126 2171
rect 2130 2168 2174 2171
rect 74 2158 118 2161
rect 290 2158 318 2161
rect 322 2158 358 2161
rect 442 2158 622 2161
rect 650 2158 694 2161
rect 918 2161 921 2168
rect 850 2158 921 2161
rect 946 2158 1574 2161
rect 1578 2158 1590 2161
rect 2214 2161 2217 2168
rect 2058 2158 2081 2161
rect 2214 2158 2254 2161
rect 2370 2158 2374 2161
rect 2378 2158 2398 2161
rect 2402 2158 2454 2161
rect 2078 2152 2081 2158
rect 106 2148 110 2151
rect 114 2148 134 2151
rect 210 2148 702 2151
rect 730 2148 766 2151
rect 770 2148 902 2151
rect 906 2148 910 2151
rect 930 2148 958 2151
rect 962 2148 1006 2151
rect 1226 2148 1254 2151
rect 1306 2148 1310 2151
rect 1314 2148 1334 2151
rect 1474 2148 1502 2151
rect 1538 2148 1662 2151
rect 1666 2148 1686 2151
rect 1810 2148 1854 2151
rect 1858 2148 1998 2151
rect 2178 2148 2206 2151
rect 2354 2148 2406 2151
rect 306 2138 342 2141
rect 410 2138 718 2141
rect 722 2138 774 2141
rect 1054 2141 1057 2148
rect 914 2138 1057 2141
rect 1066 2138 1086 2141
rect 1194 2138 1310 2141
rect 1330 2138 1382 2141
rect 1442 2138 1454 2141
rect 1650 2138 1702 2141
rect 1818 2138 1878 2141
rect 1922 2138 1929 2141
rect 2050 2138 2158 2141
rect 2162 2138 2214 2141
rect 2418 2138 2470 2141
rect 1926 2132 1929 2138
rect 218 2128 438 2131
rect 442 2128 526 2131
rect 746 2128 750 2131
rect 1082 2128 1150 2131
rect 1186 2128 1742 2131
rect 1746 2128 1806 2131
rect 1078 2122 1081 2128
rect 210 2118 238 2121
rect 330 2118 414 2121
rect 746 2118 758 2121
rect 914 2118 942 2121
rect 970 2118 990 2121
rect 1250 2118 1350 2121
rect 1354 2118 1438 2121
rect 1458 2118 1462 2121
rect 1674 2118 1769 2121
rect 2194 2118 2310 2121
rect 2410 2118 2446 2121
rect 1766 2112 1769 2118
rect 106 2108 158 2111
rect 162 2108 406 2111
rect 546 2108 662 2111
rect 730 2108 766 2111
rect 794 2108 942 2111
rect 1138 2108 1174 2111
rect 1314 2108 1430 2111
rect 1434 2108 1486 2111
rect 1490 2108 1566 2111
rect 1570 2108 1622 2111
rect 1626 2108 1654 2111
rect 984 2103 986 2107
rect 990 2103 993 2107
rect 998 2103 1000 2107
rect 2016 2103 2018 2107
rect 2022 2103 2025 2107
rect 2030 2103 2032 2107
rect 250 2098 582 2101
rect 1034 2098 1078 2101
rect 1354 2098 1414 2101
rect 1610 2098 1910 2101
rect 1914 2098 2009 2101
rect 2202 2098 2262 2101
rect 2266 2098 2358 2101
rect 18 2088 153 2091
rect 282 2088 542 2091
rect 578 2088 734 2091
rect 738 2088 1230 2091
rect 1234 2088 1694 2091
rect 1914 2088 1934 2091
rect 1942 2088 1950 2091
rect 1954 2088 1958 2091
rect 2006 2091 2009 2098
rect 2494 2092 2497 2098
rect 2006 2088 2254 2091
rect 2290 2088 2406 2091
rect 150 2082 153 2088
rect 278 2078 358 2081
rect 658 2078 750 2081
rect 778 2078 886 2081
rect 890 2078 902 2081
rect 978 2078 1006 2081
rect 1010 2078 1030 2081
rect 1162 2078 1238 2081
rect 1450 2078 1454 2081
rect 1602 2078 1614 2081
rect 1706 2078 1766 2081
rect 1770 2078 1798 2081
rect 1890 2078 1950 2081
rect 1954 2078 2022 2081
rect 2030 2078 2422 2081
rect 2462 2081 2465 2088
rect 2462 2078 2486 2081
rect 86 2072 89 2078
rect 150 2071 153 2078
rect 278 2072 281 2078
rect 150 2068 222 2071
rect 298 2068 622 2071
rect 626 2068 1238 2071
rect 1366 2071 1369 2078
rect 1366 2068 1494 2071
rect 1546 2068 1590 2071
rect 1642 2068 1670 2071
rect 1682 2068 1734 2071
rect 1874 2068 1902 2071
rect 2030 2071 2033 2078
rect 1922 2068 2033 2071
rect 2118 2068 2137 2071
rect 2242 2068 2302 2071
rect 2306 2068 2326 2071
rect 66 2058 126 2061
rect 178 2058 190 2061
rect 294 2061 297 2068
rect 2118 2062 2121 2068
rect 2134 2062 2137 2068
rect 282 2058 297 2061
rect 378 2058 409 2061
rect 498 2058 510 2061
rect 594 2058 606 2061
rect 610 2058 630 2061
rect 674 2058 694 2061
rect 718 2058 734 2061
rect 978 2058 1014 2061
rect 1026 2058 1046 2061
rect 1058 2058 1126 2061
rect 1282 2058 1286 2061
rect 1290 2058 1382 2061
rect 1402 2058 1422 2061
rect 1482 2058 1942 2061
rect 1946 2058 1974 2061
rect 1994 2058 1998 2061
rect 2194 2058 2206 2061
rect 2338 2058 2358 2061
rect 2470 2058 2486 2061
rect 406 2052 409 2058
rect 718 2052 721 2058
rect 982 2052 985 2058
rect 1126 2052 1129 2058
rect 2470 2052 2473 2058
rect 114 2048 134 2051
rect 330 2048 390 2051
rect 450 2048 590 2051
rect 1218 2048 1334 2051
rect 1698 2048 1806 2051
rect 1930 2048 1934 2051
rect 1970 2048 2086 2051
rect 2314 2048 2342 2051
rect 134 2042 137 2048
rect 562 2038 630 2041
rect 802 2038 822 2041
rect 898 2038 1022 2041
rect 1050 2038 1662 2041
rect 1666 2038 1686 2041
rect 1690 2038 2054 2041
rect 954 2028 1030 2031
rect 1138 2028 1158 2031
rect 1306 2028 1878 2031
rect 2450 2028 2470 2031
rect 346 2018 502 2021
rect 594 2018 646 2021
rect 650 2018 702 2021
rect 1130 2018 1438 2021
rect 1442 2018 1478 2021
rect 610 2008 1126 2011
rect 1154 2008 1366 2011
rect 1570 2008 1614 2011
rect 1730 2008 2438 2011
rect 2442 2008 2518 2011
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 494 2003 496 2007
rect 1496 2003 1498 2007
rect 1502 2003 1505 2007
rect 1510 2003 1512 2007
rect 770 1998 1270 2001
rect 1330 1998 1446 2001
rect 1954 1998 2222 2001
rect 194 1988 230 1991
rect 274 1988 446 1991
rect 450 1988 742 1991
rect 746 1988 750 1991
rect 978 1988 1606 1991
rect 2226 1988 2246 1991
rect 506 1978 558 1981
rect 1274 1978 1398 1981
rect 1402 1978 1406 1981
rect 1418 1978 1630 1981
rect 1666 1978 1737 1981
rect 1262 1972 1265 1978
rect 1734 1972 1737 1978
rect 2186 1978 2214 1981
rect 2314 1978 2366 1981
rect 2370 1978 2486 1981
rect 1862 1972 1865 1978
rect 66 1968 102 1971
rect 274 1968 406 1971
rect 410 1968 462 1971
rect 1178 1968 1182 1971
rect 1354 1968 1606 1971
rect 1610 1968 1694 1971
rect 2098 1968 2246 1971
rect 2434 1968 2518 1971
rect 310 1958 318 1961
rect 322 1958 350 1961
rect 514 1958 526 1961
rect 554 1958 566 1961
rect 650 1958 654 1961
rect 678 1961 681 1968
rect 678 1958 686 1961
rect 714 1958 958 1961
rect 970 1958 1014 1961
rect 1330 1958 1654 1961
rect 1658 1958 1814 1961
rect 2002 1958 2078 1961
rect 2090 1958 2142 1961
rect 2170 1958 2182 1961
rect 2186 1958 2198 1961
rect 2226 1958 2270 1961
rect 2426 1958 2446 1961
rect 90 1948 129 1951
rect 290 1948 310 1951
rect 418 1948 457 1951
rect 126 1942 129 1948
rect 454 1942 457 1948
rect 586 1948 606 1951
rect 626 1948 630 1951
rect 802 1948 806 1951
rect 954 1948 958 1951
rect 1010 1948 1078 1951
rect 1206 1951 1209 1958
rect 2326 1952 2329 1958
rect 1114 1948 1209 1951
rect 1302 1948 1318 1951
rect 1434 1948 1438 1951
rect 1474 1948 1574 1951
rect 1714 1948 1726 1951
rect 1938 1948 1958 1951
rect 2010 1948 2158 1951
rect 2194 1948 2262 1951
rect 2338 1948 2382 1951
rect 518 1942 521 1948
rect 606 1942 609 1948
rect 686 1942 689 1948
rect 702 1942 705 1948
rect 1302 1942 1305 1948
rect 1406 1942 1409 1948
rect 2006 1942 2009 1948
rect 318 1938 430 1941
rect 650 1938 654 1941
rect 778 1938 798 1941
rect 894 1938 1062 1941
rect 1154 1938 1278 1941
rect 1410 1938 1438 1941
rect 1498 1938 1526 1941
rect 1826 1938 1910 1941
rect 1914 1938 1918 1941
rect 2090 1938 2134 1941
rect 2138 1938 2158 1941
rect 2162 1938 2254 1941
rect 2450 1938 2462 1941
rect 318 1932 321 1938
rect 618 1928 638 1931
rect 726 1931 729 1938
rect 642 1928 729 1931
rect 894 1932 897 1938
rect 1374 1932 1377 1938
rect 1446 1932 1449 1938
rect 2462 1932 2465 1938
rect 954 1928 966 1931
rect 1178 1928 1254 1931
rect 1482 1928 1582 1931
rect 1914 1928 1918 1931
rect 682 1918 934 1921
rect 1162 1918 1182 1921
rect 1186 1918 1414 1921
rect 1442 1918 1878 1921
rect 1890 1918 1942 1921
rect 1978 1918 2038 1921
rect 2042 1918 2134 1921
rect 2186 1918 2334 1921
rect 214 1912 217 1918
rect 1298 1908 1534 1911
rect 1874 1908 1902 1911
rect 2106 1908 2318 1911
rect 984 1903 986 1907
rect 990 1903 993 1907
rect 998 1903 1000 1907
rect 2016 1903 2018 1907
rect 2022 1903 2025 1907
rect 2030 1903 2032 1907
rect 810 1898 902 1901
rect 906 1898 958 1901
rect 1242 1898 1446 1901
rect 2122 1898 2198 1901
rect 410 1888 470 1891
rect 474 1888 486 1891
rect 546 1888 718 1891
rect 882 1888 926 1891
rect 1306 1888 1310 1891
rect 1322 1888 1478 1891
rect 1490 1888 1518 1891
rect 1522 1888 1529 1891
rect 1610 1888 1654 1891
rect 1794 1888 1862 1891
rect 1866 1888 1894 1891
rect 2002 1888 2030 1891
rect 342 1881 345 1888
rect 342 1878 438 1881
rect 442 1878 510 1881
rect 562 1878 630 1881
rect 658 1878 814 1881
rect 818 1878 910 1881
rect 962 1878 1174 1881
rect 1258 1878 1550 1881
rect 1866 1878 1870 1881
rect 2334 1881 2337 1888
rect 2298 1878 2337 1881
rect 2474 1878 2502 1881
rect 18 1868 110 1871
rect 210 1868 222 1871
rect 226 1868 294 1871
rect 298 1868 334 1871
rect 338 1868 390 1871
rect 610 1868 670 1871
rect 738 1868 742 1871
rect 850 1868 862 1871
rect 866 1868 966 1871
rect 1002 1868 1110 1871
rect 1170 1868 1174 1871
rect 1274 1868 1398 1871
rect 1434 1868 1446 1871
rect 1450 1868 1486 1871
rect 1498 1868 1526 1871
rect 1586 1868 1622 1871
rect 1742 1871 1745 1878
rect 1626 1868 1750 1871
rect 1754 1868 1798 1871
rect 1834 1868 1958 1871
rect 1982 1868 2070 1871
rect 2346 1868 2462 1871
rect 82 1858 94 1861
rect 122 1858 142 1861
rect 146 1858 190 1861
rect 242 1858 321 1861
rect 338 1858 350 1861
rect 454 1861 457 1868
rect 434 1858 457 1861
rect 474 1858 574 1861
rect 678 1861 681 1868
rect 638 1858 681 1861
rect 810 1858 878 1861
rect 1074 1858 1142 1861
rect 1262 1861 1265 1868
rect 1542 1862 1545 1868
rect 1982 1862 1985 1868
rect 1202 1858 1265 1861
rect 1418 1858 1502 1861
rect 1658 1858 1694 1861
rect 1850 1858 1854 1861
rect 1882 1858 1886 1861
rect 2098 1858 2150 1861
rect 2178 1858 2182 1861
rect 2334 1861 2337 1868
rect 2290 1858 2337 1861
rect 318 1852 321 1858
rect 574 1852 577 1858
rect 638 1852 641 1858
rect 718 1852 721 1858
rect 1310 1852 1313 1858
rect 34 1848 46 1851
rect 134 1848 294 1851
rect 442 1848 534 1851
rect 666 1848 670 1851
rect 882 1848 894 1851
rect 1154 1848 1182 1851
rect 1466 1848 1566 1851
rect 1578 1848 1582 1851
rect 1614 1851 1617 1858
rect 1614 1848 1646 1851
rect 1998 1851 2001 1858
rect 1714 1848 2001 1851
rect 2186 1848 2246 1851
rect 2266 1848 2278 1851
rect 2282 1848 2414 1851
rect 134 1842 137 1848
rect 1326 1842 1329 1848
rect 162 1838 382 1841
rect 538 1838 622 1841
rect 666 1838 1070 1841
rect 1394 1838 1470 1841
rect 1482 1838 1606 1841
rect 1818 1838 1830 1841
rect 1834 1838 1838 1841
rect 1858 1838 1862 1841
rect 1898 1838 1998 1841
rect 578 1828 694 1831
rect 802 1828 1038 1831
rect 1482 1828 1782 1831
rect 1818 1828 2142 1831
rect 2146 1828 2150 1831
rect 2306 1828 2390 1831
rect 426 1818 446 1821
rect 450 1818 854 1821
rect 874 1818 926 1821
rect 930 1818 950 1821
rect 954 1818 1622 1821
rect 1626 1818 2326 1821
rect 2402 1818 2454 1821
rect 2482 1818 2486 1821
rect 266 1808 302 1811
rect 506 1808 1054 1811
rect 1058 1808 1430 1811
rect 1746 1808 1774 1811
rect 1818 1808 1846 1811
rect 1994 1808 2174 1811
rect 2242 1808 2310 1811
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 494 1803 496 1807
rect 1496 1803 1498 1807
rect 1502 1803 1505 1807
rect 1510 1803 1512 1807
rect 98 1798 446 1801
rect 666 1798 1382 1801
rect 1554 1798 2230 1801
rect 2234 1798 2262 1801
rect 258 1788 297 1791
rect 306 1788 510 1791
rect 522 1788 590 1791
rect 1130 1788 1350 1791
rect 1522 1788 1558 1791
rect 1562 1788 1590 1791
rect 1722 1788 2102 1791
rect 2122 1788 2334 1791
rect 2338 1788 2406 1791
rect 18 1778 150 1781
rect 154 1778 246 1781
rect 294 1781 297 1788
rect 294 1778 486 1781
rect 594 1778 638 1781
rect 922 1778 1214 1781
rect 1762 1778 1822 1781
rect 1826 1778 1854 1781
rect 90 1768 174 1771
rect 178 1768 246 1771
rect 314 1768 318 1771
rect 1034 1768 1054 1771
rect 1058 1768 1142 1771
rect 1202 1768 1718 1771
rect 1742 1771 1745 1778
rect 1742 1768 1806 1771
rect 2106 1768 2374 1771
rect 146 1758 166 1761
rect 186 1758 190 1761
rect 234 1758 270 1761
rect 274 1758 326 1761
rect 526 1761 529 1768
rect 514 1758 529 1761
rect 630 1761 633 1768
rect 630 1758 702 1761
rect 730 1758 982 1761
rect 1170 1758 1182 1761
rect 1354 1758 1478 1761
rect 1498 1758 1502 1761
rect 1542 1758 1550 1761
rect 1554 1758 1593 1761
rect 1602 1758 1662 1761
rect 1690 1758 1758 1761
rect 2066 1758 2198 1761
rect 2346 1758 2374 1761
rect 2486 1761 2489 1768
rect 2450 1758 2489 1761
rect 2502 1758 2510 1761
rect 70 1751 73 1758
rect 70 1748 118 1751
rect 146 1748 182 1751
rect 186 1748 214 1751
rect 398 1751 401 1758
rect 1014 1752 1017 1758
rect 1262 1752 1265 1758
rect 298 1748 369 1751
rect 398 1748 441 1751
rect 466 1748 470 1751
rect 530 1748 542 1751
rect 782 1748 862 1751
rect 962 1748 966 1751
rect 366 1742 369 1748
rect 438 1742 441 1748
rect 638 1742 641 1748
rect 782 1742 785 1748
rect 1106 1748 1158 1751
rect 1294 1751 1297 1758
rect 1294 1748 1334 1751
rect 1458 1748 1486 1751
rect 1502 1751 1505 1758
rect 1502 1748 1534 1751
rect 1554 1748 1566 1751
rect 1590 1751 1593 1758
rect 1590 1748 1606 1751
rect 1686 1751 1689 1758
rect 2254 1752 2257 1758
rect 2502 1752 2505 1758
rect 1686 1748 1702 1751
rect 1722 1748 1734 1751
rect 1754 1748 1758 1751
rect 1842 1748 1918 1751
rect 1970 1748 2038 1751
rect 2102 1748 2150 1751
rect 2170 1748 2254 1751
rect 2102 1742 2105 1748
rect 2350 1742 2353 1748
rect 2478 1742 2481 1748
rect 106 1738 142 1741
rect 214 1738 222 1741
rect 226 1738 262 1741
rect 542 1738 569 1741
rect 794 1738 974 1741
rect 1026 1738 1038 1741
rect 1042 1738 1230 1741
rect 1282 1738 1302 1741
rect 1378 1738 1438 1741
rect 1490 1738 1558 1741
rect 1706 1738 1710 1741
rect 1962 1738 1982 1741
rect 2010 1738 2038 1741
rect 2050 1738 2062 1741
rect 2114 1738 2262 1741
rect 542 1732 545 1738
rect 566 1732 569 1738
rect 1318 1732 1321 1738
rect 130 1728 182 1731
rect 186 1728 206 1731
rect 210 1728 350 1731
rect 778 1728 886 1731
rect 946 1728 982 1731
rect 1426 1728 1654 1731
rect 1674 1728 1694 1731
rect 2082 1728 2214 1731
rect 2250 1728 2286 1731
rect 2482 1728 2494 1731
rect 1310 1722 1313 1728
rect 602 1718 606 1721
rect 610 1718 630 1721
rect 690 1718 790 1721
rect 842 1718 870 1721
rect 978 1718 1238 1721
rect 1334 1718 1398 1721
rect 2098 1718 2110 1721
rect 2274 1718 2390 1721
rect 2394 1718 2406 1721
rect 242 1708 374 1711
rect 514 1708 846 1711
rect 1042 1708 1142 1711
rect 1146 1708 1190 1711
rect 1194 1708 1230 1711
rect 1234 1708 1294 1711
rect 1334 1711 1337 1718
rect 1318 1708 1337 1711
rect 1346 1708 1478 1711
rect 1482 1708 1926 1711
rect 2090 1708 2118 1711
rect 2370 1708 2462 1711
rect 984 1703 986 1707
rect 990 1703 993 1707
rect 998 1703 1000 1707
rect 530 1698 702 1701
rect 874 1698 950 1701
rect 1026 1698 1038 1701
rect 1318 1701 1321 1708
rect 2016 1703 2018 1707
rect 2022 1703 2025 1707
rect 2030 1703 2032 1707
rect 1226 1698 1321 1701
rect 1658 1698 1726 1701
rect 1730 1698 1870 1701
rect 1930 1698 1950 1701
rect 2378 1698 2438 1701
rect 2442 1698 2486 1701
rect 122 1688 206 1691
rect 354 1688 454 1691
rect 634 1688 678 1691
rect 682 1688 734 1691
rect 962 1688 1086 1691
rect 1134 1688 1190 1691
rect 1326 1691 1329 1698
rect 1250 1688 1329 1691
rect 1650 1688 1782 1691
rect 1826 1688 2054 1691
rect 2322 1688 2350 1691
rect 2354 1688 2358 1691
rect 230 1681 233 1688
rect 230 1678 246 1681
rect 306 1678 358 1681
rect 558 1681 561 1688
rect 1134 1682 1137 1688
rect 418 1678 561 1681
rect 642 1678 758 1681
rect 762 1678 782 1681
rect 882 1678 974 1681
rect 978 1678 1006 1681
rect 1290 1678 1310 1681
rect 1746 1678 1830 1681
rect 1874 1678 1926 1681
rect 1938 1678 2070 1681
rect 2154 1678 2214 1681
rect 2470 1681 2473 1688
rect 2410 1678 2473 1681
rect 154 1668 190 1671
rect 258 1668 318 1671
rect 338 1668 390 1671
rect 394 1668 406 1671
rect 458 1668 494 1671
rect 522 1668 854 1671
rect 930 1668 942 1671
rect 946 1668 1238 1671
rect 1422 1671 1425 1678
rect 1298 1668 1425 1671
rect 1682 1668 1686 1671
rect 1714 1668 2222 1671
rect 2254 1668 2374 1671
rect 2254 1662 2257 1668
rect 122 1658 174 1661
rect 194 1658 198 1661
rect 354 1658 473 1661
rect 650 1658 662 1661
rect 698 1658 702 1661
rect 714 1658 742 1661
rect 746 1658 798 1661
rect 922 1658 926 1661
rect 938 1658 1014 1661
rect 1090 1658 1166 1661
rect 1226 1658 1246 1661
rect 1266 1658 1278 1661
rect 1450 1658 1494 1661
rect 1602 1658 1606 1661
rect 1706 1658 1734 1661
rect 1738 1658 1745 1661
rect 1754 1658 1774 1661
rect 1802 1658 1926 1661
rect 1930 1658 1958 1661
rect 2066 1658 2086 1661
rect 2098 1658 2118 1661
rect 2122 1658 2174 1661
rect 2186 1658 2254 1661
rect 470 1652 473 1658
rect 1558 1652 1561 1658
rect 50 1648 318 1651
rect 322 1648 342 1651
rect 426 1648 430 1651
rect 434 1648 446 1651
rect 570 1648 641 1651
rect 794 1648 814 1651
rect 842 1648 846 1651
rect 962 1648 1182 1651
rect 1286 1648 1382 1651
rect 1426 1648 1550 1651
rect 1610 1648 1614 1651
rect 1658 1648 1678 1651
rect 1754 1648 1758 1651
rect 1770 1648 1870 1651
rect 2138 1648 2158 1651
rect 638 1642 641 1648
rect 1286 1642 1289 1648
rect 186 1638 193 1641
rect 378 1638 438 1641
rect 450 1638 462 1641
rect 514 1638 582 1641
rect 882 1638 894 1641
rect 898 1638 990 1641
rect 994 1638 1030 1641
rect 1034 1638 1166 1641
rect 1622 1641 1625 1648
rect 2110 1642 2113 1648
rect 1622 1638 1806 1641
rect 1850 1638 2046 1641
rect 190 1632 193 1638
rect 370 1628 518 1631
rect 846 1631 849 1638
rect 846 1628 1302 1631
rect 1314 1628 1430 1631
rect 1434 1628 1958 1631
rect 394 1618 478 1621
rect 522 1618 542 1621
rect 546 1618 582 1621
rect 1242 1618 1542 1621
rect 1602 1618 1718 1621
rect 2370 1618 2374 1621
rect 666 1608 878 1611
rect 882 1608 1142 1611
rect 1146 1608 1174 1611
rect 1530 1608 1574 1611
rect 1730 1608 1982 1611
rect 2426 1608 2446 1611
rect 398 1602 401 1608
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 494 1603 496 1607
rect 1496 1603 1498 1607
rect 1502 1603 1505 1607
rect 1510 1603 1512 1607
rect 650 1598 718 1601
rect 722 1598 1126 1601
rect 1130 1598 1326 1601
rect 1986 1598 2166 1601
rect 770 1588 790 1591
rect 1178 1588 1294 1591
rect 1330 1588 1334 1591
rect 1362 1588 1846 1591
rect 2018 1588 2046 1591
rect 2050 1588 2142 1591
rect 278 1582 281 1588
rect 434 1578 686 1581
rect 1186 1578 1545 1581
rect 1898 1578 2070 1581
rect 2098 1578 2134 1581
rect 2170 1578 2462 1581
rect 814 1572 817 1578
rect 458 1568 526 1571
rect 602 1568 662 1571
rect 1034 1568 1262 1571
rect 1542 1571 1545 1578
rect 1542 1568 1718 1571
rect 1722 1568 1734 1571
rect 1738 1568 1758 1571
rect 1926 1568 2062 1571
rect 2170 1568 2318 1571
rect 2322 1568 2494 1571
rect 1926 1562 1929 1568
rect 106 1558 110 1561
rect 114 1558 142 1561
rect 202 1558 294 1561
rect 298 1558 641 1561
rect 658 1558 670 1561
rect 682 1558 758 1561
rect 786 1558 870 1561
rect 1146 1558 1246 1561
rect 1250 1558 1278 1561
rect 1426 1558 1438 1561
rect 1442 1558 1446 1561
rect 1482 1558 1486 1561
rect 1562 1558 1590 1561
rect 1594 1558 1606 1561
rect 1754 1558 1817 1561
rect 1826 1558 1926 1561
rect 1962 1558 1977 1561
rect 2026 1558 2206 1561
rect 2330 1558 2342 1561
rect -26 1551 -22 1552
rect -26 1548 6 1551
rect 58 1548 126 1551
rect 170 1548 182 1551
rect 226 1548 238 1551
rect 362 1548 366 1551
rect 386 1548 465 1551
rect 482 1548 486 1551
rect 638 1551 641 1558
rect 638 1548 774 1551
rect 794 1548 814 1551
rect 938 1548 998 1551
rect 1002 1548 1054 1551
rect 1122 1548 1150 1551
rect 1186 1548 1233 1551
rect 1302 1551 1305 1558
rect 1638 1552 1641 1558
rect 1242 1548 1305 1551
rect 1338 1548 1454 1551
rect 1674 1548 1774 1551
rect 1814 1551 1817 1558
rect 1814 1548 1878 1551
rect 1946 1548 1966 1551
rect 1974 1551 1977 1558
rect 1974 1548 2094 1551
rect 2138 1548 2230 1551
rect 2234 1548 2278 1551
rect 2354 1548 2433 1551
rect 2482 1548 2486 1551
rect 206 1542 209 1548
rect 462 1542 465 1548
rect 114 1538 158 1541
rect 266 1538 422 1541
rect 630 1541 633 1548
rect 546 1538 633 1541
rect 690 1538 846 1541
rect 858 1538 942 1541
rect 946 1538 966 1541
rect 1026 1538 1038 1541
rect 1042 1538 1054 1541
rect 1082 1538 1094 1541
rect 1098 1538 1222 1541
rect 1230 1541 1233 1548
rect 2430 1542 2433 1548
rect 1230 1538 1262 1541
rect 1434 1538 1470 1541
rect 1474 1538 1478 1541
rect 1578 1538 1662 1541
rect 1722 1538 1734 1541
rect 1774 1538 1782 1541
rect 1786 1538 1790 1541
rect 1794 1538 1830 1541
rect 1914 1538 2246 1541
rect 2250 1538 2254 1541
rect 2258 1538 2342 1541
rect 226 1528 302 1531
rect 346 1528 566 1531
rect 570 1528 686 1531
rect 794 1528 1134 1531
rect 1138 1528 1182 1531
rect 1538 1528 1702 1531
rect 1706 1528 1750 1531
rect 178 1518 422 1521
rect 770 1518 806 1521
rect 1002 1518 1070 1521
rect 1090 1518 1246 1521
rect 1986 1518 1990 1521
rect 1994 1518 2030 1521
rect 354 1508 470 1511
rect 562 1508 742 1511
rect 1114 1508 1217 1511
rect 1234 1508 1358 1511
rect 1402 1508 1630 1511
rect 1866 1508 1902 1511
rect 984 1503 986 1507
rect 990 1503 993 1507
rect 998 1503 1000 1507
rect 1214 1502 1217 1508
rect 2016 1503 2018 1507
rect 2022 1503 2025 1507
rect 2030 1503 2032 1507
rect 2502 1502 2505 1508
rect 10 1498 374 1501
rect 570 1498 574 1501
rect 578 1498 790 1501
rect 1058 1498 1166 1501
rect 1170 1498 1182 1501
rect 1218 1498 1310 1501
rect 1690 1498 1782 1501
rect 2418 1498 2478 1501
rect 330 1488 358 1491
rect 378 1488 414 1491
rect 418 1488 502 1491
rect 506 1488 526 1491
rect 530 1488 550 1491
rect 674 1488 678 1491
rect 778 1488 910 1491
rect 1074 1488 1326 1491
rect 1386 1488 1526 1491
rect 1618 1488 1662 1491
rect 1666 1488 1702 1491
rect 1954 1488 2206 1491
rect 2234 1488 2278 1491
rect 2434 1488 2438 1491
rect 734 1482 737 1488
rect 798 1482 801 1488
rect 34 1478 326 1481
rect 330 1478 374 1481
rect 410 1478 486 1481
rect 490 1478 542 1481
rect 546 1478 582 1481
rect 898 1478 1086 1481
rect 1090 1478 1230 1481
rect 1354 1478 1366 1481
rect 1370 1478 1494 1481
rect 1562 1478 1726 1481
rect 1730 1478 1742 1481
rect 1930 1478 2062 1481
rect 2194 1478 2214 1481
rect 2218 1478 2502 1481
rect -26 1471 -22 1472
rect -26 1468 6 1471
rect 42 1468 126 1471
rect 146 1468 254 1471
rect 346 1468 358 1471
rect 386 1468 430 1471
rect 450 1468 566 1471
rect 698 1468 750 1471
rect 954 1468 1006 1471
rect 1298 1468 1358 1471
rect 1434 1468 1486 1471
rect 1594 1468 1646 1471
rect 1682 1468 1798 1471
rect 1994 1468 2022 1471
rect 2034 1468 2070 1471
rect 2074 1468 2086 1471
rect 2218 1468 2230 1471
rect 2290 1468 2382 1471
rect 374 1462 377 1468
rect -26 1458 30 1461
rect 122 1458 142 1461
rect 146 1458 150 1461
rect 210 1458 278 1461
rect 330 1458 342 1461
rect 434 1458 438 1461
rect 482 1458 518 1461
rect 750 1458 758 1461
rect 762 1458 846 1461
rect 866 1458 958 1461
rect 962 1458 990 1461
rect 1102 1461 1105 1468
rect 1026 1458 1105 1461
rect 1258 1458 1510 1461
rect 1514 1458 1702 1461
rect 1726 1458 1790 1461
rect 1842 1458 1902 1461
rect 1906 1458 1910 1461
rect 2018 1458 2049 1461
rect 2138 1458 2142 1461
rect 2250 1458 2286 1461
rect 2290 1458 2294 1461
rect 2306 1458 2318 1461
rect 2390 1461 2393 1468
rect 2386 1458 2393 1461
rect 2446 1461 2449 1468
rect 2410 1458 2449 1461
rect -26 1452 -23 1458
rect 1470 1452 1473 1458
rect 1726 1452 1729 1458
rect 2046 1452 2049 1458
rect 2222 1452 2225 1458
rect -26 1448 -22 1452
rect 10 1448 310 1451
rect 314 1448 446 1451
rect 474 1448 478 1451
rect 682 1448 838 1451
rect 1218 1448 1302 1451
rect 1482 1448 1526 1451
rect 1562 1448 1590 1451
rect 1594 1448 1710 1451
rect 1978 1448 1990 1451
rect 2170 1448 2190 1451
rect 2270 1448 2278 1451
rect 2282 1448 2342 1451
rect 2362 1448 2398 1451
rect 58 1438 166 1441
rect 266 1438 286 1441
rect 290 1438 878 1441
rect 954 1438 974 1441
rect 2394 1438 2398 1441
rect 218 1428 1014 1431
rect 1018 1428 1174 1431
rect 1178 1428 2038 1431
rect 2386 1428 2390 1431
rect 2394 1428 2406 1431
rect 258 1418 302 1421
rect 306 1418 374 1421
rect 754 1418 766 1421
rect 938 1418 1166 1421
rect 1434 1418 1478 1421
rect 1482 1418 1550 1421
rect 1586 1418 1846 1421
rect 370 1408 430 1411
rect 514 1408 662 1411
rect 890 1408 942 1411
rect 1274 1408 1462 1411
rect 1842 1408 1934 1411
rect 2130 1408 2134 1411
rect 2138 1408 2158 1411
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 494 1403 496 1407
rect 1496 1403 1498 1407
rect 1502 1403 1505 1407
rect 1510 1403 1512 1407
rect 106 1398 230 1401
rect 522 1398 654 1401
rect 658 1398 726 1401
rect 738 1398 758 1401
rect 786 1398 1118 1401
rect 1882 1398 1926 1401
rect 42 1388 126 1391
rect 130 1388 270 1391
rect 446 1388 454 1391
rect 458 1388 678 1391
rect 858 1388 934 1391
rect 1074 1388 1110 1391
rect 1114 1388 1558 1391
rect 1570 1388 1974 1391
rect 154 1378 174 1381
rect 178 1378 598 1381
rect 634 1378 718 1381
rect 722 1378 1014 1381
rect 1210 1378 1334 1381
rect 1554 1378 1942 1381
rect 246 1368 486 1371
rect 650 1368 702 1371
rect 866 1368 1094 1371
rect 1098 1368 1310 1371
rect 1914 1368 2118 1371
rect 2122 1368 2166 1371
rect 246 1362 249 1368
rect 170 1358 201 1361
rect 274 1358 646 1361
rect 734 1361 737 1368
rect 734 1358 854 1361
rect 866 1358 878 1361
rect 882 1358 894 1361
rect 1010 1358 1142 1361
rect 1146 1358 1158 1361
rect 1202 1358 1238 1361
rect 1362 1358 1390 1361
rect 1466 1358 1478 1361
rect 1482 1358 1654 1361
rect 1678 1361 1681 1368
rect 1678 1358 1766 1361
rect 1846 1361 1849 1368
rect 1826 1358 1849 1361
rect 1962 1358 1974 1361
rect 2106 1358 2302 1361
rect 2322 1358 2382 1361
rect 198 1352 201 1358
rect -26 1351 -22 1352
rect -26 1348 6 1351
rect 90 1348 166 1351
rect 410 1348 414 1351
rect 434 1348 454 1351
rect 466 1348 470 1351
rect 522 1348 630 1351
rect 802 1348 814 1351
rect 818 1348 846 1351
rect 850 1348 854 1351
rect 934 1351 937 1358
rect 1238 1352 1241 1358
rect 890 1348 937 1351
rect 962 1348 1046 1351
rect 1066 1348 1134 1351
rect 1242 1348 1254 1351
rect 1506 1348 1534 1351
rect 1570 1348 1574 1351
rect 1650 1348 1694 1351
rect 1722 1348 1742 1351
rect 1802 1348 1894 1351
rect 1986 1348 2070 1351
rect 2146 1348 2222 1351
rect 2334 1348 2377 1351
rect 2334 1342 2337 1348
rect 2374 1342 2377 1348
rect 154 1338 158 1341
rect 162 1338 262 1341
rect 266 1338 286 1341
rect 410 1338 526 1341
rect 586 1338 638 1341
rect 762 1338 790 1341
rect 810 1338 1030 1341
rect 1170 1338 1262 1341
rect 1482 1338 1486 1341
rect 1522 1338 1550 1341
rect 1594 1338 1726 1341
rect 1762 1338 1878 1341
rect 1886 1338 1942 1341
rect 2154 1338 2174 1341
rect 1886 1332 1889 1338
rect 138 1328 190 1331
rect 218 1328 254 1331
rect 258 1328 278 1331
rect 434 1328 510 1331
rect 546 1328 606 1331
rect 610 1328 742 1331
rect 850 1328 886 1331
rect 1306 1328 1374 1331
rect 1378 1328 1830 1331
rect 1834 1328 1870 1331
rect 146 1318 318 1321
rect 394 1318 454 1321
rect 458 1318 838 1321
rect 906 1318 974 1321
rect 978 1318 990 1321
rect 1138 1318 1222 1321
rect 1226 1318 1270 1321
rect 1322 1318 1406 1321
rect 1410 1318 1806 1321
rect 1810 1318 1862 1321
rect 2290 1318 2486 1321
rect 378 1308 446 1311
rect 530 1308 598 1311
rect 802 1308 822 1311
rect 1250 1308 1334 1311
rect 1354 1308 1382 1311
rect 1386 1308 1518 1311
rect 1522 1308 1566 1311
rect 1698 1308 1846 1311
rect 1866 1308 1910 1311
rect 2066 1308 2254 1311
rect 2258 1308 2342 1311
rect 2346 1308 2438 1311
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 2016 1303 2018 1307
rect 2022 1303 2025 1307
rect 2030 1303 2032 1307
rect 330 1298 470 1301
rect 538 1298 686 1301
rect 690 1298 822 1301
rect 1162 1298 1310 1301
rect 1458 1298 1574 1301
rect 1578 1298 1646 1301
rect 1650 1298 1750 1301
rect 1754 1298 1886 1301
rect 2170 1298 2270 1301
rect 2274 1298 2358 1301
rect 194 1288 390 1291
rect 586 1288 625 1291
rect 714 1288 870 1291
rect 898 1288 910 1291
rect 938 1288 1198 1291
rect 1202 1288 1286 1291
rect 1386 1288 1398 1291
rect 1402 1288 1542 1291
rect 1658 1288 1670 1291
rect 1754 1288 1838 1291
rect 1842 1288 1862 1291
rect 1938 1288 2014 1291
rect 2018 1288 2102 1291
rect 2154 1288 2254 1291
rect 2414 1291 2417 1298
rect 2414 1288 2470 1291
rect 98 1278 118 1281
rect 122 1278 286 1281
rect 438 1281 441 1288
rect 454 1281 457 1288
rect 438 1278 457 1281
rect 622 1282 625 1288
rect 698 1278 846 1281
rect 866 1278 1014 1281
rect 1026 1278 1190 1281
rect 1426 1278 1470 1281
rect 1506 1278 1598 1281
rect 1746 1278 1814 1281
rect 1914 1278 1950 1281
rect 1978 1278 2182 1281
rect 2410 1278 2414 1281
rect 302 1272 305 1278
rect 58 1268 129 1271
rect 178 1268 222 1271
rect 242 1268 294 1271
rect 498 1268 654 1271
rect 658 1268 670 1271
rect 674 1268 694 1271
rect 786 1268 822 1271
rect 1018 1268 1022 1271
rect 1146 1268 1150 1271
rect 1370 1268 1414 1271
rect 1442 1268 1614 1271
rect 1618 1268 1734 1271
rect 1898 1268 1950 1271
rect 2210 1268 2246 1271
rect 2266 1268 2390 1271
rect 2458 1268 2470 1271
rect 126 1262 129 1268
rect 170 1258 174 1261
rect 302 1258 358 1261
rect 422 1261 425 1268
rect 942 1262 945 1268
rect 974 1262 977 1268
rect 422 1258 446 1261
rect 450 1258 486 1261
rect 586 1258 686 1261
rect 778 1258 782 1261
rect 826 1258 830 1261
rect 834 1258 926 1261
rect 1010 1258 1046 1261
rect 1086 1261 1089 1268
rect 1086 1258 1102 1261
rect 1238 1261 1241 1268
rect 1186 1258 1241 1261
rect 1562 1259 1614 1261
rect 1558 1258 1614 1259
rect 1658 1258 1758 1261
rect 1914 1258 1990 1261
rect 2070 1261 2073 1268
rect 2070 1258 2118 1261
rect 2202 1258 2222 1261
rect 2226 1258 2262 1261
rect 2382 1258 2390 1261
rect 2410 1258 2446 1261
rect 50 1248 110 1251
rect 114 1248 142 1251
rect 182 1251 185 1258
rect 302 1252 305 1258
rect 382 1252 385 1258
rect 1854 1252 1857 1258
rect 2382 1252 2385 1258
rect 182 1248 198 1251
rect 338 1248 350 1251
rect 466 1248 558 1251
rect 626 1248 638 1251
rect 650 1248 654 1251
rect 658 1248 710 1251
rect 730 1248 814 1251
rect 818 1248 862 1251
rect 930 1248 1110 1251
rect 1154 1248 1174 1251
rect 1282 1248 1606 1251
rect 1610 1248 1638 1251
rect 1642 1248 1662 1251
rect 1730 1248 1782 1251
rect 2122 1248 2126 1251
rect 2130 1248 2142 1251
rect 2202 1248 2206 1251
rect 2246 1248 2318 1251
rect 2394 1248 2486 1251
rect 2246 1242 2249 1248
rect 106 1238 318 1241
rect 362 1238 430 1241
rect 434 1238 470 1241
rect 474 1238 1398 1241
rect 1538 1238 1662 1241
rect 1690 1238 1782 1241
rect 1930 1238 2150 1241
rect 2154 1238 2158 1241
rect 466 1228 494 1231
rect 714 1228 894 1231
rect 954 1228 1006 1231
rect 1034 1228 1710 1231
rect 1714 1228 1734 1231
rect 1738 1228 1798 1231
rect 2434 1228 2454 1231
rect 130 1218 134 1221
rect 138 1218 670 1221
rect 746 1218 878 1221
rect 882 1218 1038 1221
rect 1058 1218 1102 1221
rect 1162 1218 1414 1221
rect 1418 1218 1438 1221
rect 1818 1218 1830 1221
rect 1834 1218 2022 1221
rect 258 1208 342 1211
rect 674 1208 1158 1211
rect 1218 1208 1390 1211
rect 1922 1208 1958 1211
rect 1962 1208 1982 1211
rect 2042 1208 2302 1211
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 1496 1203 1498 1207
rect 1502 1203 1505 1207
rect 1510 1203 1512 1207
rect 666 1198 718 1201
rect 802 1198 806 1201
rect 906 1198 950 1201
rect 1018 1198 1158 1201
rect 1842 1198 1870 1201
rect 1874 1198 2246 1201
rect 2250 1198 2350 1201
rect 2354 1198 2422 1201
rect 2426 1198 2462 1201
rect 638 1192 641 1198
rect 186 1188 214 1191
rect 698 1188 790 1191
rect 794 1188 942 1191
rect 1074 1188 1142 1191
rect 1402 1188 2326 1191
rect 2330 1188 2390 1191
rect 746 1178 814 1181
rect 1046 1178 1094 1181
rect 1098 1178 1150 1181
rect 1162 1178 1902 1181
rect 2386 1178 2486 1181
rect 1046 1172 1049 1178
rect 2254 1172 2257 1178
rect 98 1168 126 1171
rect 130 1168 214 1171
rect 234 1168 238 1171
rect 490 1168 622 1171
rect 802 1168 886 1171
rect 890 1168 934 1171
rect 938 1168 1046 1171
rect 1066 1168 1150 1171
rect 1154 1168 1462 1171
rect 1650 1168 1726 1171
rect 1738 1168 1870 1171
rect 1874 1168 1910 1171
rect 2090 1168 2102 1171
rect 82 1158 222 1161
rect 290 1158 318 1161
rect 442 1158 454 1161
rect 538 1158 590 1161
rect 646 1161 649 1168
rect 646 1158 686 1161
rect 754 1158 870 1161
rect 954 1158 974 1161
rect 1074 1158 1086 1161
rect 1306 1158 1374 1161
rect 1378 1158 1398 1161
rect 1442 1158 1462 1161
rect 1582 1161 1585 1168
rect 1958 1162 1961 1168
rect 1546 1158 1585 1161
rect 1722 1158 1750 1161
rect 1754 1158 1758 1161
rect 1858 1158 1878 1161
rect 2198 1161 2201 1168
rect 2398 1162 2401 1168
rect 2130 1158 2201 1161
rect 2314 1158 2382 1161
rect 1718 1152 1721 1158
rect 122 1148 166 1151
rect 386 1148 438 1151
rect 594 1148 606 1151
rect 674 1148 681 1151
rect 114 1138 118 1141
rect 122 1138 142 1141
rect 302 1141 305 1148
rect 146 1138 305 1141
rect 574 1141 577 1148
rect 466 1138 577 1141
rect 678 1142 681 1148
rect 810 1148 814 1151
rect 818 1148 830 1151
rect 946 1148 958 1151
rect 962 1148 966 1151
rect 994 1148 1022 1151
rect 1026 1148 1046 1151
rect 1078 1148 1134 1151
rect 1186 1148 1230 1151
rect 1570 1148 1622 1151
rect 1774 1151 1777 1158
rect 2430 1152 2433 1158
rect 1762 1148 1777 1151
rect 1938 1148 1958 1151
rect 1962 1148 1974 1151
rect 2210 1148 2326 1151
rect 2346 1148 2414 1151
rect 782 1142 785 1148
rect 1078 1142 1081 1148
rect 714 1138 742 1141
rect 970 1138 1046 1141
rect 1362 1138 1366 1141
rect 1482 1138 1598 1141
rect 1602 1138 1702 1141
rect 1706 1138 1718 1141
rect 1822 1141 1825 1148
rect 1722 1138 1910 1141
rect 1962 1138 2038 1141
rect 2202 1138 2222 1141
rect 2290 1138 2318 1141
rect 2378 1138 2417 1141
rect 2414 1132 2417 1138
rect 74 1128 174 1131
rect 178 1128 342 1131
rect 442 1128 446 1131
rect 450 1128 462 1131
rect 466 1128 833 1131
rect 890 1128 998 1131
rect 1042 1128 1046 1131
rect 1050 1128 1150 1131
rect 1186 1128 1206 1131
rect 1346 1128 1934 1131
rect 1978 1128 2302 1131
rect 2306 1128 2374 1131
rect 666 1118 726 1121
rect 730 1118 822 1121
rect 830 1121 833 1128
rect 830 1118 1006 1121
rect 1042 1118 1054 1121
rect 1082 1118 1278 1121
rect 1298 1118 1422 1121
rect 1498 1118 1534 1121
rect 1554 1118 1574 1121
rect 1610 1118 1614 1121
rect 1650 1118 1670 1121
rect 1714 1118 1758 1121
rect 1818 1118 1990 1121
rect 2414 1112 2417 1118
rect 402 1108 494 1111
rect 498 1108 670 1111
rect 674 1108 710 1111
rect 1042 1108 1110 1111
rect 1114 1108 1142 1111
rect 1202 1108 1222 1111
rect 1362 1108 1398 1111
rect 1490 1108 1654 1111
rect 1658 1108 1702 1111
rect 1746 1108 1750 1111
rect 1826 1108 1974 1111
rect 2098 1108 2190 1111
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 2016 1103 2018 1107
rect 2022 1103 2025 1107
rect 2030 1103 2032 1107
rect 722 1098 790 1101
rect 826 1098 870 1101
rect 1058 1098 1078 1101
rect 1082 1098 1182 1101
rect 1194 1098 1230 1101
rect 1290 1098 1334 1101
rect 1354 1098 1638 1101
rect 1642 1098 1686 1101
rect 1698 1098 1710 1101
rect 1898 1098 1942 1101
rect 2494 1092 2497 1098
rect 18 1088 182 1091
rect 234 1088 278 1091
rect 282 1088 366 1091
rect 546 1088 590 1091
rect 610 1088 830 1091
rect 850 1088 926 1091
rect 1154 1088 1878 1091
rect 1882 1088 1982 1091
rect 2034 1088 2270 1091
rect 2290 1088 2294 1091
rect 2370 1088 2414 1091
rect 2418 1088 2438 1091
rect 2442 1088 2446 1091
rect 10 1078 302 1081
rect 306 1078 446 1081
rect 450 1078 902 1081
rect 906 1078 1134 1081
rect 1138 1078 1262 1081
rect 1266 1078 2246 1081
rect 2250 1078 2446 1081
rect 138 1068 230 1071
rect 274 1068 302 1071
rect 426 1068 486 1071
rect 490 1068 502 1071
rect 554 1068 646 1071
rect 850 1068 950 1071
rect 954 1068 974 1071
rect 978 1068 1342 1071
rect 1346 1068 1830 1071
rect 1834 1068 2102 1071
rect 2186 1068 2238 1071
rect 2242 1068 2254 1071
rect 2282 1068 2374 1071
rect 2378 1068 2390 1071
rect 126 1062 129 1068
rect 194 1059 246 1061
rect 190 1058 246 1059
rect 442 1058 638 1061
rect 642 1058 678 1061
rect 682 1058 686 1061
rect 730 1058 790 1061
rect 866 1058 918 1061
rect 922 1058 1038 1061
rect 1058 1058 1086 1061
rect 1090 1058 1238 1061
rect 1330 1058 1966 1061
rect 1970 1058 1998 1061
rect 2010 1058 2014 1061
rect 2150 1061 2153 1068
rect 2438 1062 2441 1068
rect 2122 1058 2153 1061
rect 2202 1058 2318 1061
rect 2322 1058 2358 1061
rect 2410 1058 2438 1061
rect 2450 1058 2478 1061
rect 2078 1052 2081 1058
rect 610 1048 662 1051
rect 706 1048 726 1051
rect 730 1048 734 1051
rect 978 1048 982 1051
rect 1010 1048 1030 1051
rect 1034 1048 1070 1051
rect 1098 1048 1102 1051
rect 1122 1048 1238 1051
rect 1242 1048 1270 1051
rect 1314 1048 1318 1051
rect 1338 1048 1366 1051
rect 1426 1048 1438 1051
rect 1562 1048 1590 1051
rect 1658 1048 1694 1051
rect 1714 1048 1726 1051
rect 1778 1048 1910 1051
rect 2114 1048 2150 1051
rect 2162 1048 2273 1051
rect 2298 1048 2302 1051
rect 2550 1051 2554 1052
rect 2314 1048 2554 1051
rect 234 1038 246 1041
rect 250 1038 270 1041
rect 274 1038 558 1041
rect 1018 1038 1062 1041
rect 1066 1038 1206 1041
rect 1346 1038 1350 1041
rect 1410 1038 1574 1041
rect 1622 1041 1625 1048
rect 2270 1042 2273 1048
rect 1622 1038 1654 1041
rect 1674 1038 2006 1041
rect 2082 1038 2086 1041
rect 2090 1038 2182 1041
rect 2202 1038 2222 1041
rect 2226 1038 2246 1041
rect 2306 1038 2318 1041
rect 226 1028 590 1031
rect 594 1028 678 1031
rect 898 1028 1182 1031
rect 1194 1028 1294 1031
rect 1474 1028 1558 1031
rect 1562 1028 1566 1031
rect 1710 1028 1718 1031
rect 1722 1028 1814 1031
rect 2058 1028 2110 1031
rect 2266 1028 2486 1031
rect 394 1018 414 1021
rect 418 1018 614 1021
rect 762 1018 1062 1021
rect 1082 1018 1126 1021
rect 1130 1018 1150 1021
rect 1226 1018 1766 1021
rect 1770 1018 1846 1021
rect 1890 1018 2094 1021
rect 2098 1018 2126 1021
rect 2162 1018 2206 1021
rect 898 1008 950 1011
rect 1146 1008 1302 1011
rect 1554 1008 1598 1011
rect 2082 1008 2094 1011
rect 2218 1008 2302 1011
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 1496 1003 1498 1007
rect 1502 1003 1505 1007
rect 1510 1003 1512 1007
rect 826 998 838 1001
rect 906 998 934 1001
rect 954 998 958 1001
rect 970 998 1110 1001
rect 1170 998 1254 1001
rect 1706 998 1814 1001
rect 2106 998 2142 1001
rect 2146 998 2158 1001
rect 474 988 806 991
rect 842 988 870 991
rect 874 988 998 991
rect 1002 988 1134 991
rect 1186 988 1214 991
rect 1218 988 1382 991
rect 1386 988 1734 991
rect 1802 988 1846 991
rect 1850 988 2102 991
rect 26 978 422 981
rect 426 978 982 981
rect 1274 978 1910 981
rect 1914 978 1934 981
rect 1938 978 1958 981
rect 234 968 278 971
rect 306 968 342 971
rect 346 968 454 971
rect 554 968 665 971
rect 682 968 702 971
rect 706 968 966 971
rect 1002 968 1118 971
rect 1122 968 1190 971
rect 1570 968 1782 971
rect 1874 968 2054 971
rect 210 958 222 961
rect 266 958 278 961
rect 282 958 294 961
rect 318 958 334 961
rect 610 958 622 961
rect 626 958 654 961
rect 662 961 665 968
rect 662 958 686 961
rect 906 958 958 961
rect 962 958 1030 961
rect 1034 958 1118 961
rect 1178 958 1326 961
rect 1330 958 1350 961
rect 1578 958 1726 961
rect 1738 958 1878 961
rect 2210 958 2270 961
rect 2322 958 2374 961
rect 2426 958 2430 961
rect 2434 958 2438 961
rect 318 952 321 958
rect 1574 952 1577 958
rect 82 948 198 951
rect 610 948 678 951
rect 698 948 718 951
rect 746 948 782 951
rect 858 948 958 951
rect 970 948 1014 951
rect 1026 948 1070 951
rect 30 941 33 948
rect 30 938 110 941
rect 130 938 166 941
rect 170 938 182 941
rect 250 938 302 941
rect 314 938 350 941
rect 526 941 529 948
rect 1202 948 1206 951
rect 1394 948 1422 951
rect 1426 948 1454 951
rect 1458 948 1502 951
rect 1754 948 1830 951
rect 1862 948 1910 951
rect 2046 951 2049 958
rect 2010 948 2049 951
rect 2138 948 2158 951
rect 2226 948 2310 951
rect 2314 948 2326 951
rect 2354 948 2430 951
rect 2434 948 2462 951
rect 386 938 761 941
rect 986 938 1014 941
rect 1026 938 1030 941
rect 1130 938 1150 941
rect 1862 942 1865 948
rect 1242 940 1342 941
rect 1238 938 1342 940
rect 1346 938 1390 941
rect 1418 938 1558 941
rect 1562 938 1750 941
rect 1962 938 2062 941
rect 2234 938 2262 941
rect 2338 938 2470 941
rect 2474 938 2478 941
rect 758 932 761 938
rect 10 928 78 931
rect 154 928 462 931
rect 882 928 1078 931
rect 1178 928 1254 931
rect 1290 928 1318 931
rect 1398 931 1401 938
rect 1378 928 1401 931
rect 1434 928 1745 931
rect 1802 928 1838 931
rect 1842 928 1894 931
rect 386 918 406 921
rect 434 918 494 921
rect 810 918 846 921
rect 938 918 966 921
rect 1066 918 1222 921
rect 1266 918 1462 921
rect 1742 921 1745 928
rect 1742 918 1838 921
rect 1842 918 1854 921
rect 1866 918 2038 921
rect 2226 918 2342 921
rect 2346 918 2430 921
rect 458 908 646 911
rect 1026 908 1142 911
rect 1170 908 1326 911
rect 1338 908 1470 911
rect 1594 908 1598 911
rect 1778 908 1982 911
rect 2090 908 2294 911
rect 2298 908 2310 911
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 2016 903 2018 907
rect 2022 903 2025 907
rect 2030 903 2032 907
rect 874 898 966 901
rect 1162 898 1174 901
rect 1210 898 1278 901
rect 1298 898 1326 901
rect 1330 898 1430 901
rect 1466 898 1662 901
rect 2306 898 2406 901
rect 210 888 238 891
rect 418 888 457 891
rect 610 888 646 891
rect 818 888 878 891
rect 946 888 974 891
rect 978 888 1030 891
rect 1114 888 1166 891
rect 1226 888 1230 891
rect 1234 888 1358 891
rect 1362 888 1582 891
rect 1602 888 1646 891
rect 1658 888 1702 891
rect 1754 888 1966 891
rect 1970 888 2078 891
rect 2266 888 2398 891
rect 454 882 457 888
rect 2510 882 2513 888
rect 66 878 110 881
rect 114 878 230 881
rect 234 878 350 881
rect 562 878 582 881
rect 586 878 902 881
rect 1034 878 1150 881
rect 1154 878 1254 881
rect 1258 878 1270 881
rect 1274 878 1278 881
rect 1298 878 1414 881
rect 1490 878 1518 881
rect 1594 878 1598 881
rect 1890 878 2097 881
rect 2130 878 2326 881
rect 2418 878 2470 881
rect -26 871 -22 872
rect -26 868 6 871
rect 10 868 14 871
rect 298 868 446 871
rect 550 871 553 878
rect 450 868 710 871
rect 734 868 753 871
rect 858 868 878 871
rect 962 868 966 871
rect 1146 868 1198 871
rect 1250 868 1294 871
rect 1298 868 1310 871
rect 1410 868 1502 871
rect 1506 868 1598 871
rect 1642 868 1654 871
rect 1690 868 1702 871
rect 1714 868 1806 871
rect 1906 868 1918 871
rect 1946 868 2030 871
rect 2034 868 2054 871
rect 2058 868 2086 871
rect 2094 871 2097 878
rect 2414 872 2417 878
rect 2094 868 2142 871
rect 2178 868 2198 871
rect 2474 868 2502 871
rect 734 862 737 868
rect 750 862 753 868
rect 362 858 382 861
rect 410 858 606 861
rect 650 858 654 861
rect 754 858 806 861
rect 890 858 910 861
rect 930 858 942 861
rect 946 858 958 861
rect 1162 858 1182 861
rect 1206 861 1209 868
rect 1206 858 1238 861
rect 1258 858 1286 861
rect 1342 861 1345 868
rect 1322 858 1446 861
rect 1466 859 1534 861
rect 1462 858 1534 859
rect 1586 858 1702 861
rect 1714 858 1758 861
rect 1822 858 1865 861
rect 1890 858 1894 861
rect 1910 858 1974 861
rect 1978 858 2046 861
rect 2194 858 2214 861
rect 2282 858 2302 861
rect 2314 858 2430 861
rect 334 852 337 858
rect 342 852 345 858
rect 1254 852 1257 858
rect 1822 852 1825 858
rect 1862 852 1865 858
rect 1910 852 1913 858
rect 26 848 86 851
rect 578 848 702 851
rect 858 848 894 851
rect 922 848 1014 851
rect 1050 848 1078 851
rect 1106 848 1166 851
rect 1202 848 1214 851
rect 1274 848 1350 851
rect 1506 848 1526 851
rect 1530 848 1558 851
rect 1562 848 1566 851
rect 1618 848 1622 851
rect 1674 848 1694 851
rect 2014 848 2022 851
rect 2026 848 2102 851
rect 2202 848 2286 851
rect 2302 848 2342 851
rect 1926 842 1929 848
rect 2302 842 2305 848
rect 202 838 230 841
rect 234 838 326 841
rect 450 838 694 841
rect 706 838 862 841
rect 970 838 1046 841
rect 1050 838 1174 841
rect 1402 838 1406 841
rect 1786 838 1894 841
rect 2090 838 2094 841
rect 2106 838 2206 841
rect 178 828 382 831
rect 386 828 702 831
rect 722 828 790 831
rect 794 828 822 831
rect 966 831 969 838
rect 826 828 969 831
rect 1210 828 1638 831
rect 1642 828 2078 831
rect 2082 828 2246 831
rect 282 818 886 821
rect 914 818 950 821
rect 1602 818 2198 821
rect 514 808 598 811
rect 602 808 926 811
rect 1186 808 1334 811
rect 1634 808 1750 811
rect 1762 808 1942 811
rect 1946 808 1974 811
rect 1994 808 2030 811
rect 2034 808 2110 811
rect 2114 808 2142 811
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 1496 803 1498 807
rect 1502 803 1505 807
rect 1510 803 1512 807
rect 538 798 582 801
rect 730 798 798 801
rect 802 798 950 801
rect 1138 798 1422 801
rect 1570 798 2126 801
rect 370 788 526 791
rect 1026 788 1318 791
rect 1322 788 1374 791
rect 1594 788 1742 791
rect 1834 788 2014 791
rect 634 778 878 781
rect 890 778 910 781
rect 986 778 1022 781
rect 1026 778 1166 781
rect 1202 778 1366 781
rect 1442 778 1670 781
rect 1674 778 1678 781
rect 1706 778 1934 781
rect 1938 778 2110 781
rect 2154 778 2302 781
rect 146 768 198 771
rect 346 768 430 771
rect 434 768 454 771
rect 498 768 558 771
rect 746 768 814 771
rect 914 768 942 771
rect 1042 768 1102 771
rect 1306 768 1310 771
rect 1322 768 1486 771
rect 1490 768 1582 771
rect 1650 768 1654 771
rect 1666 768 1694 771
rect 1794 768 1953 771
rect 1978 768 2166 771
rect 1950 762 1953 768
rect 306 758 310 761
rect 314 758 326 761
rect 330 758 334 761
rect 770 758 918 761
rect 922 758 926 761
rect 1034 758 1046 761
rect 1050 758 1086 761
rect 1098 758 1102 761
rect 1282 758 1334 761
rect 1434 758 1454 761
rect 1458 758 1654 761
rect 1682 758 1742 761
rect 1842 758 1846 761
rect 1882 758 1942 761
rect 2026 758 2049 761
rect 118 752 121 758
rect -26 751 -22 752
rect -26 748 102 751
rect 138 748 158 751
rect 162 748 166 751
rect 190 751 193 758
rect 190 748 214 751
rect 250 748 294 751
rect 330 748 377 751
rect 538 748 614 751
rect 650 748 670 751
rect 730 748 758 751
rect 762 748 982 751
rect 1034 748 1038 751
rect 1162 748 1166 751
rect 1174 751 1177 758
rect 1366 752 1369 758
rect 2046 752 2049 758
rect 2162 758 2190 761
rect 2490 758 2494 761
rect 2070 752 2073 758
rect 1174 748 1222 751
rect 1298 748 1310 751
rect 1322 748 1342 751
rect 1346 748 1353 751
rect 1382 748 1390 751
rect 1394 748 1406 751
rect 374 742 377 748
rect 1078 742 1081 748
rect 1538 748 1606 751
rect 1610 748 1617 751
rect 1626 748 1694 751
rect 1842 748 1846 751
rect 1882 748 1905 751
rect 1954 748 1974 751
rect 2154 748 2254 751
rect 2450 748 2462 751
rect 58 738 126 741
rect 130 738 190 741
rect 194 738 238 741
rect 258 738 270 741
rect 274 738 310 741
rect 530 738 542 741
rect 634 738 857 741
rect 898 738 926 741
rect 930 738 942 741
rect 946 738 950 741
rect 1050 738 1062 741
rect 1082 738 1174 741
rect 1202 738 1518 741
rect 1610 738 1614 741
rect 1674 738 1702 741
rect 1710 741 1713 748
rect 1902 742 1905 748
rect 1710 738 1806 741
rect 1810 738 1886 741
rect 2010 738 2014 741
rect 2050 738 2054 741
rect 2150 741 2153 748
rect 2122 738 2153 741
rect 2198 738 2294 741
rect 2402 738 2422 741
rect 2474 738 2494 741
rect 446 732 449 738
rect 854 732 857 738
rect 1654 732 1657 738
rect 2198 732 2201 738
rect 722 728 774 731
rect 858 728 1038 731
rect 1042 728 1150 731
rect 1154 728 1158 731
rect 1170 728 1246 731
rect 1298 728 1302 731
rect 1698 728 1817 731
rect 1938 728 1998 731
rect 450 718 462 721
rect 506 718 686 721
rect 774 721 777 728
rect 1814 722 1817 728
rect 774 718 862 721
rect 906 718 1022 721
rect 1122 718 1134 721
rect 1138 718 1230 721
rect 1282 718 1390 721
rect 1394 718 1438 721
rect 1578 718 1774 721
rect 1842 718 1990 721
rect 1994 718 2086 721
rect 2114 718 2174 721
rect 458 708 534 711
rect 538 708 758 711
rect 834 708 974 711
rect 1010 708 1158 711
rect 1170 708 1294 711
rect 1330 708 1414 711
rect 1426 708 1622 711
rect 1626 708 1654 711
rect 1674 708 1910 711
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 2016 703 2018 707
rect 2022 703 2025 707
rect 2030 703 2032 707
rect 178 698 198 701
rect 202 698 342 701
rect 714 698 894 701
rect 902 698 926 701
rect 930 698 942 701
rect 1058 698 1062 701
rect 1066 698 1438 701
rect 1602 698 1854 701
rect 2042 698 2094 701
rect 2130 698 2158 701
rect 106 688 214 691
rect 298 688 630 691
rect 634 688 670 691
rect 902 691 905 698
rect 2510 692 2513 698
rect 690 688 905 691
rect 914 688 929 691
rect 962 688 1150 691
rect 1162 688 1182 691
rect 1202 688 1238 691
rect 1242 688 1286 691
rect 1518 688 1726 691
rect 1730 688 1742 691
rect 1866 688 1937 691
rect 2026 688 2206 691
rect 2266 688 2334 691
rect 2338 688 2422 691
rect 50 678 54 681
rect 322 678 358 681
rect 402 678 518 681
rect 562 678 582 681
rect 586 678 766 681
rect 778 678 830 681
rect 842 678 878 681
rect 882 678 918 681
rect 926 681 929 688
rect 1518 682 1521 688
rect 926 678 1006 681
rect 1066 678 1070 681
rect 1146 678 1166 681
rect 1282 678 1334 681
rect 1682 678 1686 681
rect 1698 678 1726 681
rect 1890 678 1926 681
rect 1934 681 1937 688
rect 1934 678 2038 681
rect 2098 678 2166 681
rect 2250 678 2254 681
rect 2290 678 2294 681
rect 2314 678 2318 681
rect 2394 678 2454 681
rect 18 668 62 671
rect 66 668 94 671
rect 214 671 217 678
rect 154 668 217 671
rect 330 668 334 671
rect 418 668 454 671
rect 466 668 486 671
rect 514 668 534 671
rect 650 668 654 671
rect 682 668 702 671
rect 762 668 902 671
rect 906 668 934 671
rect 938 668 942 671
rect 1046 671 1049 678
rect 1046 668 1222 671
rect 1258 668 1302 671
rect 1362 668 1374 671
rect 1518 671 1521 678
rect 1450 668 1521 671
rect 1562 668 1622 671
rect 1930 668 1934 671
rect 2034 668 2118 671
rect 2122 668 2126 671
rect 2138 668 2142 671
rect 2154 668 2206 671
rect 2238 671 2241 678
rect 2238 668 2358 671
rect 294 662 297 668
rect 350 662 353 668
rect 26 658 46 661
rect 50 658 54 661
rect 78 658 278 661
rect 378 658 382 661
rect 402 658 406 661
rect 414 658 454 661
rect 550 661 553 668
rect 474 658 553 661
rect 582 662 585 668
rect 750 662 753 668
rect 1702 662 1705 668
rect 1734 662 1737 668
rect 1990 662 1993 668
rect 2454 662 2457 668
rect 634 658 686 661
rect 738 658 742 661
rect 762 658 766 661
rect 794 658 798 661
rect 818 658 822 661
rect 850 658 910 661
rect 1070 658 1094 661
rect 1102 658 1118 661
rect 1146 658 1302 661
rect 1306 658 1326 661
rect 1362 658 1430 661
rect 1754 658 1870 661
rect 1946 658 1950 661
rect 2058 658 2062 661
rect 2066 658 2297 661
rect 78 652 81 658
rect 414 652 417 658
rect 1070 652 1073 658
rect 1102 652 1105 658
rect 1910 652 1913 658
rect 2294 652 2297 658
rect 298 648 310 651
rect 586 648 790 651
rect 866 648 934 651
rect 1138 648 1166 651
rect 1186 648 1206 651
rect 1418 648 1534 651
rect 1618 648 1630 651
rect 1634 648 1646 651
rect 1682 648 1838 651
rect 1914 648 1998 651
rect 2146 648 2153 651
rect 518 641 521 648
rect 518 638 558 641
rect 574 641 577 648
rect 1078 642 1081 648
rect 2150 642 2153 648
rect 574 638 590 641
rect 602 638 606 641
rect 642 638 790 641
rect 798 638 1014 641
rect 1162 638 1230 641
rect 1274 638 1398 641
rect 1434 638 1614 641
rect 798 631 801 638
rect 346 628 801 631
rect 1298 628 2134 631
rect 878 621 881 628
rect 530 618 886 621
rect 890 618 2262 621
rect 2266 618 2462 621
rect 506 608 590 611
rect 642 608 662 611
rect 666 608 910 611
rect 922 608 1206 611
rect 1394 608 1462 611
rect 1466 608 1486 611
rect 1538 608 2318 611
rect 2322 608 2382 611
rect 2386 608 2390 611
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 1496 603 1498 607
rect 1502 603 1505 607
rect 1510 603 1512 607
rect 522 598 878 601
rect 1018 598 1254 601
rect 1258 598 1294 601
rect 1618 598 2214 601
rect 2282 598 2302 601
rect 170 588 270 591
rect 274 588 294 591
rect 298 588 686 591
rect 786 588 854 591
rect 946 588 1150 591
rect 1378 588 1886 591
rect 1906 588 2046 591
rect 2290 588 2398 591
rect 10 578 94 581
rect 98 578 142 581
rect 434 578 518 581
rect 618 578 806 581
rect 1090 578 1150 581
rect 1402 578 1590 581
rect 1762 578 2078 581
rect 2290 578 2302 581
rect 2326 572 2329 578
rect 554 568 726 571
rect 818 568 998 571
rect 1002 568 1086 571
rect 1106 568 1126 571
rect 1146 568 1206 571
rect 1210 568 1374 571
rect 1538 568 1558 571
rect 2058 568 2278 571
rect 22 562 25 568
rect 446 562 449 568
rect 26 558 46 561
rect 458 558 462 561
rect 578 558 622 561
rect 642 558 662 561
rect 682 558 742 561
rect 746 558 774 561
rect 874 558 918 561
rect 1122 558 1174 561
rect 1178 558 1182 561
rect 1898 558 2030 561
rect 2374 561 2377 568
rect 2314 558 2377 561
rect 86 551 89 558
rect 38 548 89 551
rect 258 548 406 551
rect 466 548 470 551
rect 514 548 614 551
rect 666 548 718 551
rect 38 542 41 548
rect 798 548 806 551
rect 810 548 830 551
rect 882 548 889 551
rect 922 548 958 551
rect 1054 551 1057 558
rect 1054 548 1102 551
rect 1334 551 1337 558
rect 1290 548 1337 551
rect 1410 548 1526 551
rect 1606 551 1609 558
rect 1554 548 1609 551
rect 1682 548 1982 551
rect 1986 548 2014 551
rect 2138 548 2318 551
rect 2338 548 2374 551
rect 862 542 865 548
rect 886 542 889 548
rect 2182 542 2185 548
rect 50 538 54 541
rect 194 538 286 541
rect 330 538 366 541
rect 466 538 566 541
rect 618 538 622 541
rect 634 538 638 541
rect 930 538 1070 541
rect 1074 538 1294 541
rect 1426 538 1438 541
rect 1458 538 1494 541
rect 1506 538 1518 541
rect 1522 538 1758 541
rect 1826 538 1870 541
rect 1882 538 1902 541
rect 1906 538 1913 541
rect 1930 538 1958 541
rect 1962 538 1974 541
rect 2218 538 2254 541
rect 2274 538 2358 541
rect 2362 538 2406 541
rect 2410 538 2422 541
rect 42 528 70 531
rect 282 528 462 531
rect 610 528 734 531
rect 858 528 934 531
rect 1034 528 1094 531
rect 1186 528 1190 531
rect 1202 528 1206 531
rect 1242 528 1462 531
rect 1906 528 2006 531
rect 582 521 585 528
rect 426 518 585 521
rect 978 518 1198 521
rect 1370 518 1526 521
rect 1586 518 1734 521
rect 1874 518 1918 521
rect 1970 518 2342 521
rect 2346 518 2430 521
rect 154 508 926 511
rect 1082 508 1134 511
rect 1138 508 1190 511
rect 1194 508 1302 511
rect 1306 508 1358 511
rect 1362 508 1406 511
rect 1442 508 1686 511
rect 1690 508 1838 511
rect 1842 508 1966 511
rect 2050 508 2150 511
rect 2154 508 2238 511
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 2016 503 2018 507
rect 2022 503 2025 507
rect 2030 503 2032 507
rect 98 498 118 501
rect 290 498 310 501
rect 378 498 486 501
rect 498 498 574 501
rect 586 498 606 501
rect 1146 498 1382 501
rect 1562 498 1678 501
rect 106 488 238 491
rect 242 488 438 491
rect 458 488 694 491
rect 714 488 758 491
rect 762 488 790 491
rect 930 488 1014 491
rect 1570 488 1590 491
rect 1622 488 1630 491
rect 1634 488 1846 491
rect 2074 488 2094 491
rect 2098 488 2182 491
rect 2346 488 2406 491
rect 2410 488 2494 491
rect 122 478 150 481
rect 154 478 302 481
rect 306 478 710 481
rect 1126 481 1129 488
rect 1126 478 1222 481
rect 1226 478 1278 481
rect 1522 478 1574 481
rect 1578 478 1670 481
rect 1802 478 2038 481
rect 2210 478 2230 481
rect 2234 478 2270 481
rect 298 468 302 471
rect 362 468 462 471
rect 538 468 625 471
rect 650 468 734 471
rect 802 468 886 471
rect 998 471 1001 478
rect 998 468 1070 471
rect 1074 468 1182 471
rect 1218 468 1302 471
rect 1386 468 1398 471
rect 1594 468 1598 471
rect 1818 468 1958 471
rect 2082 468 2118 471
rect 2178 468 2278 471
rect 2386 468 2438 471
rect 622 462 625 468
rect 910 462 913 468
rect 122 458 142 461
rect 146 458 150 461
rect 154 458 318 461
rect 322 458 342 461
rect 730 458 742 461
rect 746 458 846 461
rect 882 458 910 461
rect 982 461 985 468
rect 982 458 1038 461
rect 1050 458 1078 461
rect 1082 458 1110 461
rect 1202 458 1222 461
rect 1542 461 1545 468
rect 1542 458 1558 461
rect 1578 458 1598 461
rect 1602 458 1606 461
rect 1650 458 1686 461
rect 1690 458 1742 461
rect 1746 458 1790 461
rect 1866 458 1870 461
rect 1874 458 1878 461
rect 1990 461 1993 468
rect 1990 458 2006 461
rect 2118 461 2121 468
rect 2034 458 2121 461
rect 2146 459 2198 461
rect 2142 458 2198 459
rect 2258 458 2265 461
rect 2338 458 2342 461
rect 2378 458 2390 461
rect 1702 452 1705 458
rect 2262 452 2265 458
rect 2390 452 2393 458
rect -26 451 -22 452
rect -26 448 6 451
rect 142 448 150 451
rect 154 448 182 451
rect 330 448 406 451
rect 602 448 774 451
rect 850 448 854 451
rect 938 448 1206 451
rect 1390 448 1422 451
rect 1802 448 1886 451
rect 1954 448 1990 451
rect 26 438 366 441
rect 454 441 457 448
rect 370 438 457 441
rect 582 442 585 448
rect 1390 442 1393 448
rect 610 438 822 441
rect 826 438 1030 441
rect 1114 438 1342 441
rect 1658 438 1854 441
rect 1858 438 2078 441
rect 2202 438 2222 441
rect 2226 438 2518 441
rect 130 428 526 431
rect 954 428 1182 431
rect 1186 428 1670 431
rect 1674 428 1694 431
rect 1786 428 1894 431
rect 554 418 974 421
rect 1210 418 1358 421
rect 1362 418 1550 421
rect 1782 421 1785 428
rect 1554 418 1785 421
rect 866 408 886 411
rect 890 408 902 411
rect 1210 408 1462 411
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 1496 403 1498 407
rect 1502 403 1505 407
rect 1510 403 1512 407
rect 866 398 1222 401
rect 162 388 182 391
rect 186 388 270 391
rect 962 388 1414 391
rect 1418 388 1438 391
rect 1866 388 1918 391
rect 1922 388 2070 391
rect 730 378 886 381
rect 890 378 982 381
rect 986 378 1110 381
rect 1346 378 1558 381
rect 1650 378 1918 381
rect 1922 378 1974 381
rect 58 368 150 371
rect 154 368 350 371
rect 378 368 390 371
rect 522 368 550 371
rect 858 368 918 371
rect 922 368 966 371
rect 1106 368 1190 371
rect 1194 368 1214 371
rect 1290 368 1310 371
rect 1314 368 1398 371
rect 1826 368 1870 371
rect 2298 368 2414 371
rect 2418 368 2502 371
rect 1662 362 1665 368
rect 106 358 414 361
rect 434 358 478 361
rect 482 358 502 361
rect 562 358 670 361
rect 674 358 870 361
rect 1082 358 1134 361
rect 1146 358 1470 361
rect 1474 358 1486 361
rect 1490 358 1646 361
rect 1862 358 1870 361
rect 1874 358 1934 361
rect 2134 361 2137 368
rect 1986 358 2137 361
rect 2218 358 2230 361
rect 2238 361 2241 368
rect 2234 358 2241 361
rect 2378 358 2398 361
rect 2402 358 2406 361
rect 2506 358 2510 361
rect 114 348 126 351
rect 142 348 150 351
rect 202 348 254 351
rect 258 348 294 351
rect 394 348 398 351
rect 418 348 446 351
rect 450 348 510 351
rect 522 348 526 351
rect 530 348 606 351
rect 674 348 678 351
rect 698 348 702 351
rect 826 348 886 351
rect 930 348 934 351
rect 978 348 1054 351
rect 1058 348 1086 351
rect 1306 348 1654 351
rect 1674 348 1766 351
rect 1818 348 1838 351
rect 1842 348 1854 351
rect 2154 348 2174 351
rect 2446 351 2449 358
rect 2402 348 2449 351
rect 142 342 145 348
rect 178 338 230 341
rect 386 338 406 341
rect 546 338 566 341
rect 770 338 873 341
rect 42 328 214 331
rect 526 331 529 338
rect 870 332 873 338
rect 1050 338 1078 341
rect 1082 338 1318 341
rect 1370 338 1414 341
rect 1458 338 1470 341
rect 1578 338 1622 341
rect 1690 338 1702 341
rect 1706 338 1718 341
rect 1778 338 2158 341
rect 2162 338 2198 341
rect 2330 338 2342 341
rect 2370 338 2433 341
rect 250 328 529 331
rect 554 328 566 331
rect 834 328 846 331
rect 886 328 894 331
rect 898 328 918 331
rect 966 331 969 338
rect 2430 332 2433 338
rect 966 328 1054 331
rect 1058 328 1118 331
rect 1426 328 1430 331
rect 1698 328 2046 331
rect 2050 328 2086 331
rect 330 318 334 321
rect 642 318 966 321
rect 1018 318 1278 321
rect 1286 318 1454 321
rect 1458 318 1670 321
rect 1714 318 1862 321
rect 2026 318 2054 321
rect 210 308 310 311
rect 690 308 734 311
rect 1286 311 1289 318
rect 1010 308 1289 311
rect 1482 308 1534 311
rect 1578 308 1758 311
rect 1762 308 1966 311
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 2016 303 2018 307
rect 2022 303 2025 307
rect 2030 303 2032 307
rect 26 298 46 301
rect 50 298 102 301
rect 314 298 382 301
rect 618 298 854 301
rect 1410 298 1414 301
rect 1522 298 1614 301
rect 1674 298 1862 301
rect 2506 298 2518 301
rect 66 288 198 291
rect 302 291 305 298
rect 302 288 502 291
rect 802 288 822 291
rect 854 291 857 298
rect 842 288 857 291
rect 978 288 1062 291
rect 1266 288 1318 291
rect 1322 288 1406 291
rect 1582 288 1590 291
rect 1594 288 1646 291
rect 1786 288 1814 291
rect 1818 288 1878 291
rect 2266 288 2294 291
rect 2314 288 2390 291
rect 2490 288 2521 291
rect 114 278 118 281
rect 490 278 662 281
rect 706 278 758 281
rect 762 278 1006 281
rect 1142 281 1145 288
rect 2518 282 2521 288
rect 1142 278 1198 281
rect 1322 278 1670 281
rect 1698 278 1774 281
rect 1866 278 2118 281
rect 1102 272 1105 278
rect 18 268 78 271
rect 474 268 590 271
rect 658 268 790 271
rect 1034 268 1086 271
rect 1110 271 1113 278
rect 1110 268 1270 271
rect 1282 268 1286 271
rect 1298 268 1350 271
rect 1418 268 1422 271
rect 1434 268 1462 271
rect 1514 268 1550 271
rect 1554 268 1590 271
rect 1642 268 2078 271
rect 2082 268 2102 271
rect 2130 268 2158 271
rect 2234 268 2358 271
rect 2494 271 2497 278
rect 2370 268 2497 271
rect 82 258 102 261
rect 806 262 809 268
rect 370 259 422 261
rect 366 258 422 259
rect 506 258 529 261
rect 586 258 601 261
rect 714 258 734 261
rect 738 258 766 261
rect 786 258 806 261
rect 838 261 841 268
rect 838 258 894 261
rect 998 261 1001 268
rect 962 258 1001 261
rect 1082 258 1102 261
rect 1138 258 1150 261
rect 1286 261 1289 268
rect 2166 262 2169 268
rect 1286 258 1302 261
rect 1306 258 1566 261
rect 1610 258 1614 261
rect 1618 258 1630 261
rect 1650 258 1654 261
rect 1666 258 1694 261
rect 1834 258 1846 261
rect 1938 258 1977 261
rect 2010 258 2054 261
rect 2098 258 2166 261
rect 2346 258 2446 261
rect 526 252 529 258
rect 598 252 601 258
rect 1974 252 1977 258
rect 2518 252 2521 258
rect 102 248 110 251
rect 114 248 142 251
rect 602 248 606 251
rect 1402 248 1822 251
rect 1854 248 1862 251
rect 1866 248 1926 251
rect 2154 248 2238 251
rect 554 238 606 241
rect 1170 238 1254 241
rect 1258 238 1430 241
rect 1442 238 1654 241
rect 1970 238 2294 241
rect 2410 238 2518 241
rect 418 228 614 231
rect 650 228 1078 231
rect 1082 228 1542 231
rect 1546 228 1726 231
rect 1914 228 2118 231
rect 474 218 878 221
rect 1266 218 1294 221
rect 1378 218 1838 221
rect 174 212 177 218
rect 706 208 710 211
rect 714 208 950 211
rect 1602 208 1702 211
rect 1706 208 1742 211
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 1496 203 1498 207
rect 1502 203 1505 207
rect 1510 203 1512 207
rect 1570 198 2214 201
rect 2218 198 2238 201
rect 886 192 889 198
rect 434 188 438 191
rect 1122 188 1126 191
rect 1386 188 1438 191
rect 1442 188 1462 191
rect 1722 188 1734 191
rect 1738 188 1750 191
rect 902 182 905 188
rect 490 178 646 181
rect 1074 178 1286 181
rect 1590 178 1598 181
rect 1602 178 1630 181
rect 1730 178 2062 181
rect 2066 178 2150 181
rect 106 168 158 171
rect 266 168 334 171
rect 338 168 534 171
rect 626 168 646 171
rect 650 168 974 171
rect 1090 168 1134 171
rect 1298 168 1382 171
rect 1586 168 1598 171
rect 1602 168 1646 171
rect 1906 168 1990 171
rect 74 158 126 161
rect 154 158 174 161
rect 810 158 998 161
rect 1034 158 1038 161
rect 1098 158 1102 161
rect 1106 158 1126 161
rect 1130 158 1390 161
rect 1418 158 1430 161
rect 1466 158 1862 161
rect 1866 158 1878 161
rect 2138 158 2254 161
rect 2410 158 2494 161
rect 10 148 102 151
rect 106 148 110 151
rect 122 148 150 151
rect 154 148 190 151
rect 262 151 265 158
rect 210 148 265 151
rect 654 151 657 158
rect 618 148 657 151
rect 826 148 838 151
rect 842 148 1014 151
rect 1022 148 1086 151
rect 1118 148 1190 151
rect 1238 148 1318 151
rect 1402 148 1430 151
rect 1522 148 1550 151
rect 1570 148 1582 151
rect 1730 148 1798 151
rect 1842 148 1918 151
rect 2102 151 2105 158
rect 2050 148 2105 151
rect 2154 148 2158 151
rect 2162 148 2182 151
rect 2242 148 2310 151
rect 146 138 150 141
rect 202 138 214 141
rect 598 141 601 148
rect 718 141 721 148
rect 1022 142 1025 148
rect 1118 142 1121 148
rect 1238 142 1241 148
rect 598 138 721 141
rect 746 138 830 141
rect 1130 138 1134 141
rect 1346 138 1406 141
rect 1434 138 1446 141
rect 1554 138 1694 141
rect 1714 138 1742 141
rect 1866 138 1950 141
rect 1954 138 2078 141
rect 2082 138 2142 141
rect 2146 138 2214 141
rect 2342 141 2345 148
rect 2358 141 2361 148
rect 2342 138 2361 141
rect 2370 138 2446 141
rect 2450 138 2486 141
rect 74 128 246 131
rect 250 128 342 131
rect 698 128 782 131
rect 1010 128 1246 131
rect 1282 128 1494 131
rect 1878 128 1942 131
rect 2010 128 2054 131
rect 2114 128 2270 131
rect 1878 122 1881 128
rect 234 118 318 121
rect 322 118 358 121
rect 570 118 654 121
rect 658 118 710 121
rect 754 118 910 121
rect 914 118 1006 121
rect 1042 118 1206 121
rect 1226 118 1326 121
rect 1402 118 1446 121
rect 1202 108 1334 111
rect 1370 108 1638 111
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect 2016 103 2018 107
rect 2022 103 2025 107
rect 2030 103 2032 107
rect 2038 102 2041 108
rect 178 98 270 101
rect 274 98 446 101
rect 1018 98 1286 101
rect 1290 98 1374 101
rect 1394 98 1454 101
rect 1458 98 1526 101
rect 2058 98 2110 101
rect 298 88 334 91
rect 338 88 414 91
rect 434 88 694 91
rect 714 88 814 91
rect 818 88 870 91
rect 894 88 1070 91
rect 1074 88 1270 91
rect 1274 88 1294 91
rect 1298 88 1430 91
rect 1538 88 1678 91
rect 1682 88 1694 91
rect 1818 88 1934 91
rect 2098 88 2438 91
rect 2466 88 2478 91
rect 894 82 897 88
rect 218 78 278 81
rect 282 78 318 81
rect 322 78 358 81
rect 426 78 438 81
rect 962 78 1078 81
rect 1434 78 1598 81
rect 1786 78 1894 81
rect 1898 78 2062 81
rect 2066 78 2158 81
rect 2162 78 2222 81
rect 2226 78 2350 81
rect 6 72 9 78
rect 122 68 142 71
rect 146 68 326 71
rect 330 68 438 71
rect 458 68 558 71
rect 582 71 585 78
rect 734 71 737 78
rect 582 68 737 71
rect 762 68 846 71
rect 866 68 1110 71
rect 1142 68 1161 71
rect 1186 68 1270 71
rect 1338 68 1406 71
rect 1558 68 1614 71
rect 1674 68 1758 71
rect 1810 68 1838 71
rect 1842 68 1966 71
rect 1978 68 2046 71
rect 2242 68 2326 71
rect 2350 71 2353 78
rect 2350 68 2422 71
rect 2442 68 2470 71
rect 2550 71 2554 72
rect 2522 68 2554 71
rect 146 58 174 61
rect 178 58 190 61
rect 202 58 430 61
rect 434 58 462 61
rect 682 58 686 61
rect 698 58 870 61
rect 1142 62 1145 68
rect 1158 62 1161 68
rect 1438 62 1441 68
rect 1558 62 1561 68
rect 1574 62 1577 68
rect 970 59 1038 61
rect 966 58 1038 59
rect 1074 58 1086 61
rect 1106 58 1142 61
rect 1266 58 1286 61
rect 1402 58 1406 61
rect 1474 58 1526 61
rect 1658 58 1694 61
rect 1698 58 2214 61
rect 2218 58 2246 61
rect 170 48 206 51
rect 314 48 358 51
rect 850 48 862 51
rect 1050 48 1062 51
rect 1066 48 1414 51
rect 1418 48 1806 51
rect 1838 48 1878 51
rect 2550 51 2554 52
rect 2482 48 2554 51
rect 1838 42 1841 48
rect 1114 28 1958 31
rect 1962 28 1982 31
rect 1422 12 1425 18
rect 1654 12 1657 18
rect 2038 12 2041 18
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
rect 1496 3 1498 7
rect 1502 3 1505 7
rect 1510 3 1512 7
<< m4contact >>
rect 482 2403 486 2407
rect 490 2403 493 2407
rect 493 2403 494 2407
rect 1498 2403 1502 2407
rect 1506 2403 1509 2407
rect 1509 2403 1510 2407
rect 926 2398 930 2402
rect 1806 2388 1810 2392
rect 2382 2358 2386 2362
rect 190 2348 194 2352
rect 1566 2348 1570 2352
rect 1830 2348 1834 2352
rect 2310 2348 2314 2352
rect 2358 2348 2362 2352
rect 2414 2348 2418 2352
rect 46 2338 50 2342
rect 1190 2338 1194 2342
rect 2206 2338 2210 2342
rect 2238 2338 2242 2342
rect 2302 2338 2306 2342
rect 2462 2338 2466 2342
rect 342 2328 346 2332
rect 974 2318 978 2322
rect 2334 2318 2338 2322
rect 2390 2318 2394 2322
rect 2446 2318 2450 2322
rect 766 2308 770 2312
rect 1814 2308 1818 2312
rect 986 2303 990 2307
rect 994 2303 997 2307
rect 997 2303 998 2307
rect 2018 2303 2022 2307
rect 2026 2303 2029 2307
rect 2029 2303 2030 2307
rect 974 2298 978 2302
rect 1358 2298 1362 2302
rect 910 2278 914 2282
rect 2358 2278 2362 2282
rect 1222 2268 1226 2272
rect 1542 2268 1546 2272
rect 390 2258 394 2262
rect 598 2258 602 2262
rect 1246 2258 1250 2262
rect 1446 2258 1450 2262
rect 1974 2258 1978 2262
rect 2158 2258 2162 2262
rect 2262 2258 2266 2262
rect 2470 2258 2474 2262
rect 438 2248 442 2252
rect 1102 2248 1106 2252
rect 1830 2248 1834 2252
rect 2286 2248 2290 2252
rect 86 2238 90 2242
rect 1054 2238 1058 2242
rect 1486 2238 1490 2242
rect 1822 2238 1826 2242
rect 2446 2238 2450 2242
rect 902 2228 906 2232
rect 1342 2228 1346 2232
rect 2350 2228 2354 2232
rect 574 2218 578 2222
rect 1150 2218 1154 2222
rect 1190 2218 1194 2222
rect 482 2203 486 2207
rect 490 2203 493 2207
rect 493 2203 494 2207
rect 1498 2203 1502 2207
rect 1506 2203 1509 2207
rect 1509 2203 1510 2207
rect 694 2198 698 2202
rect 1062 2198 1066 2202
rect 2118 2188 2122 2192
rect 2454 2188 2458 2192
rect 1822 2178 1826 2182
rect 1902 2178 1906 2182
rect 342 2168 346 2172
rect 1006 2168 1010 2172
rect 2126 2168 2130 2172
rect 942 2158 946 2162
rect 2374 2158 2378 2162
rect 110 2148 114 2152
rect 1006 2148 1010 2152
rect 1310 2148 1314 2152
rect 1854 2148 1858 2152
rect 1438 2138 1442 2142
rect 1918 2138 1922 2142
rect 742 2128 746 2132
rect 1742 2128 1746 2132
rect 1806 2128 1810 2132
rect 966 2118 970 2122
rect 1078 2118 1082 2122
rect 1454 2118 1458 2122
rect 942 2108 946 2112
rect 986 2103 990 2107
rect 994 2103 997 2107
rect 997 2103 998 2107
rect 2018 2103 2022 2107
rect 2026 2103 2029 2107
rect 2029 2103 2030 2107
rect 734 2088 738 2092
rect 1694 2088 1698 2092
rect 2494 2088 2498 2092
rect 1454 2078 1458 2082
rect 86 2068 90 2072
rect 974 2058 978 2062
rect 1054 2058 1058 2062
rect 1126 2058 1130 2062
rect 1998 2058 2002 2062
rect 134 2048 138 2052
rect 1694 2048 1698 2052
rect 1934 2048 1938 2052
rect 1022 2038 1026 2042
rect 1158 2028 1162 2032
rect 1302 2028 1306 2032
rect 2446 2028 2450 2032
rect 502 2018 506 2022
rect 590 2018 594 2022
rect 1126 2018 1130 2022
rect 482 2003 486 2007
rect 490 2003 493 2007
rect 493 2003 494 2007
rect 1498 2003 1502 2007
rect 1506 2003 1509 2007
rect 1509 2003 1510 2007
rect 230 1988 234 1992
rect 750 1988 754 1992
rect 974 1988 978 1992
rect 2222 1988 2226 1992
rect 1406 1978 1410 1982
rect 2366 1978 2370 1982
rect 1174 1968 1178 1972
rect 1262 1968 1266 1972
rect 1862 1968 1866 1972
rect 2518 1968 2522 1972
rect 566 1958 570 1962
rect 646 1958 650 1962
rect 1326 1958 1330 1962
rect 1654 1958 1658 1962
rect 2198 1958 2202 1962
rect 2422 1958 2426 1962
rect 414 1948 418 1952
rect 518 1948 522 1952
rect 606 1948 610 1952
rect 630 1948 634 1952
rect 686 1948 690 1952
rect 798 1948 802 1952
rect 950 1948 954 1952
rect 1438 1948 1442 1952
rect 2006 1948 2010 1952
rect 2158 1948 2162 1952
rect 2326 1948 2330 1952
rect 654 1938 658 1942
rect 702 1938 706 1942
rect 1374 1938 1378 1942
rect 1406 1938 1410 1942
rect 1438 1938 1442 1942
rect 1918 1938 1922 1942
rect 2446 1938 2450 1942
rect 2462 1938 2466 1942
rect 638 1928 642 1932
rect 950 1928 954 1932
rect 1446 1928 1450 1932
rect 1910 1928 1914 1932
rect 1438 1918 1442 1922
rect 2182 1918 2186 1922
rect 214 1908 218 1912
rect 1870 1908 1874 1912
rect 2102 1908 2106 1912
rect 2318 1908 2322 1912
rect 986 1903 990 1907
rect 994 1903 997 1907
rect 997 1903 998 1907
rect 2018 1903 2022 1907
rect 2026 1903 2029 1907
rect 2029 1903 2030 1907
rect 1302 1888 1306 1892
rect 1862 1878 1866 1882
rect 742 1868 746 1872
rect 1174 1868 1178 1872
rect 1486 1868 1490 1872
rect 1494 1868 1498 1872
rect 1750 1868 1754 1872
rect 2342 1868 2346 1872
rect 350 1858 354 1862
rect 470 1858 474 1862
rect 574 1858 578 1862
rect 718 1858 722 1862
rect 1542 1858 1546 1862
rect 1846 1858 1850 1862
rect 1878 1858 1882 1862
rect 1998 1858 2002 1862
rect 2094 1858 2098 1862
rect 2182 1858 2186 1862
rect 662 1848 666 1852
rect 1310 1848 1314 1852
rect 1582 1848 1586 1852
rect 1710 1848 1714 1852
rect 2182 1848 2186 1852
rect 2414 1848 2418 1852
rect 382 1838 386 1842
rect 1070 1838 1074 1842
rect 1326 1838 1330 1842
rect 1830 1838 1834 1842
rect 1854 1838 1858 1842
rect 1478 1828 1482 1832
rect 1814 1828 1818 1832
rect 854 1818 858 1822
rect 870 1818 874 1822
rect 2398 1818 2402 1822
rect 2486 1818 2490 1822
rect 302 1808 306 1812
rect 502 1808 506 1812
rect 1054 1808 1058 1812
rect 482 1803 486 1807
rect 490 1803 493 1807
rect 493 1803 494 1807
rect 1498 1803 1502 1807
rect 1506 1803 1509 1807
rect 1509 1803 1510 1807
rect 662 1798 666 1802
rect 1550 1798 1554 1802
rect 2230 1798 2234 1802
rect 510 1788 514 1792
rect 2102 1788 2106 1792
rect 1822 1778 1826 1782
rect 1854 1778 1858 1782
rect 318 1768 322 1772
rect 2102 1768 2106 1772
rect 166 1758 170 1762
rect 190 1758 194 1762
rect 1478 1758 1482 1762
rect 1502 1758 1506 1762
rect 2374 1758 2378 1762
rect 2510 1758 2514 1762
rect 142 1748 146 1752
rect 462 1748 466 1752
rect 862 1748 866 1752
rect 966 1748 970 1752
rect 1014 1748 1018 1752
rect 1262 1748 1266 1752
rect 1334 1748 1338 1752
rect 1758 1748 1762 1752
rect 1966 1748 1970 1752
rect 2166 1748 2170 1752
rect 2254 1748 2258 1752
rect 2350 1748 2354 1752
rect 638 1738 642 1742
rect 790 1738 794 1742
rect 1022 1738 1026 1742
rect 1230 1738 1234 1742
rect 1702 1738 1706 1742
rect 1958 1738 1962 1742
rect 2006 1738 2010 1742
rect 2046 1738 2050 1742
rect 2110 1738 2114 1742
rect 2478 1738 2482 1742
rect 206 1728 210 1732
rect 1310 1728 1314 1732
rect 1318 1728 1322 1732
rect 1670 1728 1674 1732
rect 598 1718 602 1722
rect 790 1718 794 1722
rect 1238 1718 1242 1722
rect 2110 1718 2114 1722
rect 2406 1718 2410 1722
rect 510 1708 514 1712
rect 1342 1708 1346 1712
rect 1926 1708 1930 1712
rect 986 1703 990 1707
rect 994 1703 997 1707
rect 997 1703 998 1707
rect 1038 1698 1042 1702
rect 2018 1703 2022 1707
rect 2026 1703 2029 1707
rect 2029 1703 2030 1707
rect 2438 1698 2442 1702
rect 1934 1678 1938 1682
rect 942 1668 946 1672
rect 1678 1668 1682 1672
rect 2222 1668 2226 1672
rect 174 1658 178 1662
rect 190 1658 194 1662
rect 350 1658 354 1662
rect 694 1658 698 1662
rect 918 1658 922 1662
rect 1598 1658 1602 1662
rect 1798 1658 1802 1662
rect 422 1648 426 1652
rect 846 1648 850 1652
rect 958 1648 962 1652
rect 1550 1648 1554 1652
rect 1558 1648 1562 1652
rect 1606 1648 1610 1652
rect 1750 1648 1754 1652
rect 1766 1648 1770 1652
rect 2110 1648 2114 1652
rect 182 1638 186 1642
rect 878 1638 882 1642
rect 1166 1638 1170 1642
rect 1846 1638 1850 1642
rect 1310 1628 1314 1632
rect 1958 1628 1962 1632
rect 582 1618 586 1622
rect 2374 1618 2378 1622
rect 1726 1608 1730 1612
rect 2422 1608 2426 1612
rect 482 1603 486 1607
rect 490 1603 493 1607
rect 493 1603 494 1607
rect 1498 1603 1502 1607
rect 1506 1603 1509 1607
rect 1509 1603 1510 1607
rect 398 1598 402 1602
rect 646 1598 650 1602
rect 1326 1598 1330 1602
rect 1174 1588 1178 1592
rect 1326 1588 1330 1592
rect 1846 1588 1850 1592
rect 278 1578 282 1582
rect 430 1578 434 1582
rect 2094 1578 2098 1582
rect 2166 1578 2170 1582
rect 814 1568 818 1572
rect 1718 1568 1722 1572
rect 102 1558 106 1562
rect 294 1558 298 1562
rect 1142 1558 1146 1562
rect 1438 1558 1442 1562
rect 1478 1558 1482 1562
rect 6 1548 10 1552
rect 382 1548 386 1552
rect 1638 1548 1642 1552
rect 1670 1548 1674 1552
rect 2486 1548 2490 1552
rect 206 1538 210 1542
rect 854 1538 858 1542
rect 1054 1538 1058 1542
rect 1222 1538 1226 1542
rect 2246 1538 2250 1542
rect 2342 1538 2346 1542
rect 1182 1528 1186 1532
rect 1982 1518 1986 1522
rect 742 1508 746 1512
rect 1230 1508 1234 1512
rect 986 1503 990 1507
rect 994 1503 997 1507
rect 997 1503 998 1507
rect 2018 1503 2022 1507
rect 2026 1503 2029 1507
rect 2029 1503 2030 1507
rect 6 1498 10 1502
rect 566 1498 570 1502
rect 574 1498 578 1502
rect 2414 1498 2418 1502
rect 2502 1498 2506 1502
rect 678 1488 682 1492
rect 734 1488 738 1492
rect 2430 1488 2434 1492
rect 30 1478 34 1482
rect 2214 1478 2218 1482
rect 6 1468 10 1472
rect 1358 1468 1362 1472
rect 2022 1468 2026 1472
rect 30 1458 34 1462
rect 142 1458 146 1462
rect 374 1458 378 1462
rect 430 1458 434 1462
rect 1254 1458 1258 1462
rect 1702 1458 1706 1462
rect 1838 1458 1842 1462
rect 1902 1458 1906 1462
rect 2142 1458 2146 1462
rect 2222 1458 2226 1462
rect 2294 1458 2298 1462
rect 2382 1458 2386 1462
rect 6 1448 10 1452
rect 478 1448 482 1452
rect 1302 1448 1306 1452
rect 1710 1448 1714 1452
rect 2358 1448 2362 1452
rect 878 1438 882 1442
rect 974 1438 978 1442
rect 2390 1438 2394 1442
rect 214 1428 218 1432
rect 1014 1428 1018 1432
rect 2390 1428 2394 1432
rect 1478 1418 1482 1422
rect 886 1408 890 1412
rect 2126 1408 2130 1412
rect 482 1403 486 1407
rect 490 1403 493 1407
rect 493 1403 494 1407
rect 1498 1403 1502 1407
rect 1506 1403 1509 1407
rect 1509 1403 1510 1407
rect 654 1398 658 1402
rect 726 1398 730 1402
rect 1878 1398 1882 1402
rect 126 1388 130 1392
rect 1110 1388 1114 1392
rect 1566 1388 1570 1392
rect 598 1378 602 1382
rect 718 1378 722 1382
rect 1014 1378 1018 1382
rect 862 1368 866 1372
rect 1310 1368 1314 1372
rect 166 1358 170 1362
rect 646 1358 650 1362
rect 894 1358 898 1362
rect 1006 1358 1010 1362
rect 1238 1358 1242 1362
rect 1390 1358 1394 1362
rect 1974 1358 1978 1362
rect 2318 1358 2322 1362
rect 406 1348 410 1352
rect 454 1348 458 1352
rect 462 1348 466 1352
rect 798 1348 802 1352
rect 854 1348 858 1352
rect 1574 1348 1578 1352
rect 582 1338 586 1342
rect 1518 1338 1522 1342
rect 1878 1338 1882 1342
rect 1302 1328 1306 1332
rect 1374 1328 1378 1332
rect 1870 1328 1874 1332
rect 838 1318 842 1322
rect 974 1318 978 1322
rect 1406 1318 1410 1322
rect 1862 1318 1866 1322
rect 2286 1318 2290 1322
rect 822 1308 826 1312
rect 986 1303 990 1307
rect 994 1303 997 1307
rect 997 1303 998 1307
rect 2018 1303 2022 1307
rect 2026 1303 2029 1307
rect 2029 1303 2030 1307
rect 470 1298 474 1302
rect 686 1298 690 1302
rect 822 1298 826 1302
rect 1574 1298 1578 1302
rect 1670 1288 1674 1292
rect 1814 1278 1818 1282
rect 1950 1278 1954 1282
rect 2414 1278 2418 1282
rect 302 1268 306 1272
rect 974 1268 978 1272
rect 1022 1268 1026 1272
rect 1150 1268 1154 1272
rect 1614 1268 1618 1272
rect 2206 1268 2210 1272
rect 2390 1268 2394 1272
rect 2470 1268 2474 1272
rect 166 1258 170 1262
rect 382 1258 386 1262
rect 822 1258 826 1262
rect 926 1258 930 1262
rect 942 1258 946 1262
rect 1758 1258 1762 1262
rect 1854 1258 1858 1262
rect 1990 1258 1994 1262
rect 2390 1258 2394 1262
rect 46 1248 50 1252
rect 350 1248 354 1252
rect 646 1248 650 1252
rect 726 1248 730 1252
rect 862 1248 866 1252
rect 1278 1248 1282 1252
rect 1662 1248 1666 1252
rect 2118 1248 2122 1252
rect 2206 1248 2210 1252
rect 2486 1248 2490 1252
rect 358 1238 362 1242
rect 1398 1238 1402 1242
rect 1926 1238 1930 1242
rect 2150 1238 2154 1242
rect 1006 1228 1010 1232
rect 1798 1228 1802 1232
rect 134 1218 138 1222
rect 670 1218 674 1222
rect 742 1218 746 1222
rect 878 1218 882 1222
rect 670 1208 674 1212
rect 1918 1208 1922 1212
rect 1958 1208 1962 1212
rect 482 1203 486 1207
rect 490 1203 493 1207
rect 493 1203 494 1207
rect 1498 1203 1502 1207
rect 1506 1203 1509 1207
rect 1509 1203 1510 1207
rect 718 1198 722 1202
rect 798 1198 802 1202
rect 1158 1198 1162 1202
rect 2462 1198 2466 1202
rect 638 1188 642 1192
rect 694 1188 698 1192
rect 1070 1188 1074 1192
rect 1398 1188 1402 1192
rect 2326 1188 2330 1192
rect 1150 1178 1154 1182
rect 1158 1178 1162 1182
rect 2254 1178 2258 1182
rect 1062 1168 1066 1172
rect 1150 1168 1154 1172
rect 870 1158 874 1162
rect 950 1158 954 1162
rect 1758 1158 1762 1162
rect 1958 1158 1962 1162
rect 2398 1158 2402 1162
rect 606 1148 610 1152
rect 670 1148 674 1152
rect 782 1148 786 1152
rect 814 1148 818 1152
rect 1046 1148 1050 1152
rect 1718 1148 1722 1152
rect 1974 1148 1978 1152
rect 2430 1148 2434 1152
rect 966 1138 970 1142
rect 1358 1138 1362 1142
rect 438 1128 442 1132
rect 1038 1128 1042 1132
rect 1182 1128 1186 1132
rect 2302 1128 2306 1132
rect 822 1118 826 1122
rect 1078 1118 1082 1122
rect 1278 1118 1282 1122
rect 1606 1118 1610 1122
rect 2414 1118 2418 1122
rect 398 1108 402 1112
rect 710 1108 714 1112
rect 1702 1108 1706 1112
rect 1750 1108 1754 1112
rect 986 1103 990 1107
rect 994 1103 997 1107
rect 997 1103 998 1107
rect 2018 1103 2022 1107
rect 2026 1103 2029 1107
rect 2029 1103 2030 1107
rect 790 1098 794 1102
rect 1078 1098 1082 1102
rect 1182 1098 1186 1102
rect 1638 1098 1642 1102
rect 1686 1098 1690 1102
rect 1694 1098 1698 1102
rect 2494 1098 2498 1102
rect 278 1088 282 1092
rect 1982 1088 1986 1092
rect 2294 1088 2298 1092
rect 2414 1088 2418 1092
rect 2446 1088 2450 1092
rect 6 1078 10 1082
rect 302 1078 306 1082
rect 902 1078 906 1082
rect 2246 1078 2250 1082
rect 2446 1078 2450 1082
rect 846 1068 850 1072
rect 1830 1068 1834 1072
rect 2374 1068 2378 1072
rect 2438 1068 2442 1072
rect 126 1058 130 1062
rect 678 1058 682 1062
rect 862 1058 866 1062
rect 1086 1058 1090 1062
rect 1238 1058 1242 1062
rect 1326 1058 1330 1062
rect 1966 1058 1970 1062
rect 2006 1058 2010 1062
rect 2078 1058 2082 1062
rect 2478 1058 2482 1062
rect 726 1048 730 1052
rect 1094 1048 1098 1052
rect 1310 1048 1314 1052
rect 1334 1048 1338 1052
rect 1654 1048 1658 1052
rect 1910 1048 1914 1052
rect 2158 1048 2162 1052
rect 2302 1048 2306 1052
rect 230 1038 234 1042
rect 1206 1038 1210 1042
rect 1342 1038 1346 1042
rect 2078 1038 2082 1042
rect 2182 1038 2186 1042
rect 2198 1038 2202 1042
rect 2222 1038 2226 1042
rect 2302 1038 2306 1042
rect 2318 1038 2322 1042
rect 590 1028 594 1032
rect 894 1028 898 1032
rect 1182 1028 1186 1032
rect 1190 1028 1194 1032
rect 1558 1028 1562 1032
rect 390 1018 394 1022
rect 1062 1018 1066 1022
rect 1846 1018 1850 1022
rect 2126 1018 2130 1022
rect 1302 1008 1306 1012
rect 2094 1008 2098 1012
rect 482 1003 486 1007
rect 490 1003 493 1007
rect 493 1003 494 1007
rect 1498 1003 1502 1007
rect 1506 1003 1509 1007
rect 1509 1003 1510 1007
rect 822 998 826 1002
rect 958 998 962 1002
rect 966 998 970 1002
rect 1254 998 1258 1002
rect 2158 998 2162 1002
rect 806 988 810 992
rect 838 988 842 992
rect 1182 988 1186 992
rect 1382 988 1386 992
rect 422 978 426 982
rect 1958 978 1962 982
rect 342 968 346 972
rect 966 968 970 972
rect 1782 968 1786 972
rect 1870 968 1874 972
rect 1118 958 1122 962
rect 1174 958 1178 962
rect 1326 958 1330 962
rect 1726 958 1730 962
rect 2430 958 2434 962
rect 678 948 682 952
rect 854 948 858 952
rect 1574 948 1578 952
rect 2350 948 2354 952
rect 2430 948 2434 952
rect 1014 938 1018 942
rect 1030 938 1034 942
rect 1750 938 1754 942
rect 2334 938 2338 942
rect 1286 928 1290 932
rect 1374 928 1378 932
rect 806 918 810 922
rect 934 918 938 922
rect 1062 918 1066 922
rect 1838 918 1842 922
rect 1862 918 1866 922
rect 646 908 650 912
rect 1142 908 1146 912
rect 1166 908 1170 912
rect 1334 908 1338 912
rect 1598 908 1602 912
rect 986 903 990 907
rect 994 903 997 907
rect 997 903 998 907
rect 2018 903 2022 907
rect 2026 903 2029 907
rect 2029 903 2030 907
rect 870 898 874 902
rect 1158 898 1162 902
rect 1294 898 1298 902
rect 1110 888 1114 892
rect 1222 888 1226 892
rect 1750 888 1754 892
rect 1030 878 1034 882
rect 1278 878 1282 882
rect 1414 878 1418 882
rect 1598 878 1602 882
rect 2510 878 2514 882
rect 6 868 10 872
rect 878 868 882 872
rect 958 868 962 872
rect 1598 868 1602 872
rect 1710 868 1714 872
rect 2414 868 2418 872
rect 2470 868 2474 872
rect 334 858 338 862
rect 646 858 650 862
rect 910 858 914 862
rect 926 858 930 862
rect 1238 858 1242 862
rect 1886 858 1890 862
rect 2310 858 2314 862
rect 22 848 26 852
rect 342 848 346 852
rect 1046 848 1050 852
rect 1254 848 1258 852
rect 1502 848 1506 852
rect 1566 848 1570 852
rect 1622 848 1626 852
rect 694 838 698 842
rect 1174 838 1178 842
rect 1398 838 1402 842
rect 1782 838 1786 842
rect 1926 838 1930 842
rect 2086 838 2090 842
rect 2206 838 2210 842
rect 382 828 386 832
rect 702 828 706 832
rect 718 828 722 832
rect 2078 828 2082 832
rect 910 818 914 822
rect 1598 818 1602 822
rect 510 808 514 812
rect 598 808 602 812
rect 1334 808 1338 812
rect 1750 808 1754 812
rect 1758 808 1762 812
rect 2110 808 2114 812
rect 482 803 486 807
rect 490 803 493 807
rect 493 803 494 807
rect 1498 803 1502 807
rect 1506 803 1509 807
rect 1509 803 1510 807
rect 726 798 730 802
rect 798 798 802 802
rect 526 788 530 792
rect 1318 788 1322 792
rect 1166 778 1170 782
rect 1198 778 1202 782
rect 1678 778 1682 782
rect 1302 768 1306 772
rect 1318 768 1322 772
rect 1654 768 1658 772
rect 1974 768 1978 772
rect 310 758 314 762
rect 326 758 330 762
rect 1102 758 1106 762
rect 1838 758 1842 762
rect 1942 758 1946 762
rect 118 748 122 752
rect 158 748 162 752
rect 1030 748 1034 752
rect 1078 748 1082 752
rect 1166 748 1170 752
rect 2494 758 2498 762
rect 1310 748 1314 752
rect 1366 748 1370 752
rect 1694 748 1698 752
rect 1846 748 1850 752
rect 1950 748 1954 752
rect 2070 748 2074 752
rect 310 738 314 742
rect 1518 738 1522 742
rect 1606 738 1610 742
rect 1654 738 1658 742
rect 2006 738 2010 742
rect 2054 738 2058 742
rect 2398 738 2402 742
rect 446 728 450 732
rect 1158 728 1162 732
rect 1166 728 1170 732
rect 1302 728 1306 732
rect 1694 728 1698 732
rect 462 718 466 722
rect 502 718 506 722
rect 1390 718 1394 722
rect 1438 718 1442 722
rect 454 708 458 712
rect 758 708 762 712
rect 974 708 978 712
rect 1006 708 1010 712
rect 1166 708 1170 712
rect 1622 708 1626 712
rect 986 703 990 707
rect 994 703 997 707
rect 997 703 998 707
rect 2018 703 2022 707
rect 2026 703 2029 707
rect 2029 703 2030 707
rect 942 698 946 702
rect 1054 698 1058 702
rect 2038 698 2042 702
rect 214 688 218 692
rect 630 688 634 692
rect 686 688 690 692
rect 1150 688 1154 692
rect 1158 688 1162 692
rect 2510 688 2514 692
rect 54 678 58 682
rect 582 678 586 682
rect 838 678 842 682
rect 1006 678 1010 682
rect 1062 678 1066 682
rect 1278 678 1282 682
rect 1686 678 1690 682
rect 2166 678 2170 682
rect 2238 678 2242 682
rect 2246 678 2250 682
rect 2286 678 2290 682
rect 2310 678 2314 682
rect 294 668 298 672
rect 334 668 338 672
rect 414 668 418 672
rect 486 668 490 672
rect 534 668 538 672
rect 654 668 658 672
rect 758 668 762 672
rect 942 668 946 672
rect 1926 668 1930 672
rect 2126 668 2130 672
rect 2142 668 2146 672
rect 46 658 50 662
rect 278 658 282 662
rect 350 658 354 662
rect 382 658 386 662
rect 406 658 410 662
rect 454 658 458 662
rect 582 658 586 662
rect 742 658 746 662
rect 750 658 754 662
rect 758 658 762 662
rect 790 658 794 662
rect 814 658 818 662
rect 1142 658 1146 662
rect 1702 658 1706 662
rect 1734 658 1738 662
rect 1750 658 1754 662
rect 1910 658 1914 662
rect 1950 658 1954 662
rect 1990 658 1994 662
rect 2054 658 2058 662
rect 2454 658 2458 662
rect 1102 648 1106 652
rect 1166 648 1170 652
rect 1206 648 1210 652
rect 1414 648 1418 652
rect 1614 648 1618 652
rect 2142 648 2146 652
rect 558 638 562 642
rect 598 638 602 642
rect 790 638 794 642
rect 1078 638 1082 642
rect 886 618 890 622
rect 590 608 594 612
rect 638 608 642 612
rect 910 608 914 612
rect 918 608 922 612
rect 2382 608 2386 612
rect 482 603 486 607
rect 490 603 493 607
rect 493 603 494 607
rect 1498 603 1502 607
rect 1506 603 1509 607
rect 1509 603 1510 607
rect 1014 598 1018 602
rect 166 588 170 592
rect 686 588 690 592
rect 430 578 434 582
rect 614 578 618 582
rect 1398 578 1402 582
rect 2302 578 2306 582
rect 2326 578 2330 582
rect 446 568 450 572
rect 1102 568 1106 572
rect 1142 568 1146 572
rect 1374 568 1378 572
rect 22 558 26 562
rect 462 558 466 562
rect 742 558 746 562
rect 918 558 922 562
rect 462 548 466 552
rect 862 548 866 552
rect 878 548 882 552
rect 1678 548 1682 552
rect 2318 548 2322 552
rect 54 538 58 542
rect 614 538 618 542
rect 630 538 634 542
rect 1070 538 1074 542
rect 1518 538 1522 542
rect 2422 538 2426 542
rect 462 528 466 532
rect 734 528 738 532
rect 1190 528 1194 532
rect 1198 528 1202 532
rect 2006 528 2010 532
rect 974 518 978 522
rect 1366 518 1370 522
rect 2430 518 2434 522
rect 150 508 154 512
rect 1438 508 1442 512
rect 1838 508 1842 512
rect 986 503 990 507
rect 994 503 997 507
rect 997 503 998 507
rect 2018 503 2022 507
rect 2026 503 2029 507
rect 2029 503 2030 507
rect 574 498 578 502
rect 1846 488 1850 492
rect 2342 488 2346 492
rect 118 478 122 482
rect 302 468 306 472
rect 910 468 914 472
rect 1398 468 1402 472
rect 2174 468 2178 472
rect 142 458 146 462
rect 846 458 850 462
rect 1110 458 1114 462
rect 1598 458 1602 462
rect 1862 458 1866 462
rect 1878 458 1882 462
rect 2254 458 2258 462
rect 2342 458 2346 462
rect 406 448 410 452
rect 582 448 586 452
rect 854 448 858 452
rect 1950 448 1954 452
rect 2390 448 2394 452
rect 606 438 610 442
rect 1030 438 1034 442
rect 1854 438 1858 442
rect 1182 428 1186 432
rect 1670 428 1674 432
rect 1894 428 1898 432
rect 1358 418 1362 422
rect 886 408 890 412
rect 1206 408 1210 412
rect 482 403 486 407
rect 490 403 493 407
rect 493 403 494 407
rect 1498 403 1502 407
rect 1506 403 1509 407
rect 1509 403 1510 407
rect 862 398 866 402
rect 958 388 962 392
rect 886 378 890 382
rect 1646 378 1650 382
rect 1918 378 1922 382
rect 1662 368 1666 372
rect 430 358 434 362
rect 502 358 506 362
rect 670 358 674 362
rect 1142 358 1146 362
rect 1646 358 1650 362
rect 1982 358 1986 362
rect 2230 358 2234 362
rect 2398 358 2402 362
rect 2502 358 2506 362
rect 110 348 114 352
rect 150 348 154 352
rect 390 348 394 352
rect 510 348 514 352
rect 526 348 530 352
rect 606 348 610 352
rect 694 348 698 352
rect 1814 348 1818 352
rect 1078 338 1082 342
rect 1318 338 1322 342
rect 2198 338 2202 342
rect 1422 328 1426 332
rect 2086 328 2090 332
rect 326 318 330 322
rect 1006 308 1010 312
rect 1574 308 1578 312
rect 986 303 990 307
rect 994 303 997 307
rect 997 303 998 307
rect 2018 303 2022 307
rect 2026 303 2029 307
rect 2029 303 2030 307
rect 102 298 106 302
rect 1414 298 1418 302
rect 1862 298 1866 302
rect 798 288 802 292
rect 2486 288 2490 292
rect 118 278 122 282
rect 702 278 706 282
rect 1006 278 1010 282
rect 1102 278 1106 282
rect 1318 278 1322 282
rect 1286 268 1290 272
rect 1414 268 1418 272
rect 1430 268 1434 272
rect 2166 268 2170 272
rect 2366 268 2370 272
rect 806 258 810 262
rect 1606 258 1610 262
rect 1654 258 1658 262
rect 598 248 602 252
rect 2518 248 2522 252
rect 1430 238 1434 242
rect 1966 238 1970 242
rect 2406 238 2410 242
rect 878 218 882 222
rect 1294 218 1298 222
rect 1374 218 1378 222
rect 174 208 178 212
rect 710 208 714 212
rect 1598 208 1602 212
rect 482 203 486 207
rect 490 203 493 207
rect 493 203 494 207
rect 1498 203 1502 207
rect 1506 203 1509 207
rect 1509 203 1510 207
rect 430 188 434 192
rect 886 188 890 192
rect 902 188 906 192
rect 1126 188 1130 192
rect 1382 188 1386 192
rect 1438 188 1442 192
rect 2150 178 2154 182
rect 102 168 106 172
rect 974 168 978 172
rect 150 158 154 162
rect 1038 158 1042 162
rect 1102 158 1106 162
rect 110 148 114 152
rect 190 148 194 152
rect 1014 148 1018 152
rect 1318 148 1322 152
rect 2158 148 2162 152
rect 150 138 154 142
rect 1134 138 1138 142
rect 2446 138 2450 142
rect 1398 118 1402 122
rect 986 103 990 107
rect 994 103 997 107
rect 997 103 998 107
rect 2018 103 2022 107
rect 2026 103 2029 107
rect 2029 103 2030 107
rect 1014 98 1018 102
rect 1374 98 1378 102
rect 2038 98 2042 102
rect 334 88 338 92
rect 2462 88 2466 92
rect 358 78 362 82
rect 6 68 10 72
rect 118 68 122 72
rect 1966 68 1970 72
rect 2470 68 2474 72
rect 174 58 178 62
rect 198 58 202 62
rect 686 58 690 62
rect 1086 58 1090 62
rect 1102 58 1106 62
rect 1406 58 1410 62
rect 1438 58 1442 62
rect 1422 18 1426 22
rect 1654 18 1658 22
rect 2038 18 2042 22
rect 482 3 486 7
rect 490 3 493 7
rect 493 3 494 7
rect 1498 3 1502 7
rect 1506 3 1509 7
rect 1509 3 1510 7
<< metal4 >>
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 494 2403 496 2407
rect 1496 2403 1498 2407
rect 1502 2403 1505 2407
rect 1510 2403 1512 2407
rect 918 2398 926 2401
rect 50 2338 54 2341
rect 86 2072 89 2238
rect 110 1561 113 2148
rect 106 1558 113 1561
rect 6 1502 9 1548
rect 6 1452 9 1468
rect 30 1462 33 1478
rect 6 872 9 1078
rect 6 72 9 868
rect 22 562 25 848
rect 46 662 49 1248
rect 46 652 49 658
rect 54 542 57 678
rect 102 302 105 1558
rect 126 1062 129 1388
rect 134 1222 137 2048
rect 190 1762 193 2348
rect 342 2172 345 2328
rect 758 2308 766 2311
rect 394 2258 398 2261
rect 594 2258 598 2261
rect 142 1462 145 1748
rect 122 748 126 751
rect 102 172 105 298
rect 110 152 113 348
rect 118 282 121 478
rect 142 462 145 1458
rect 166 1362 169 1758
rect 190 1672 193 1758
rect 190 1662 193 1668
rect 174 1651 177 1658
rect 174 1648 185 1651
rect 182 1642 185 1648
rect 166 1262 169 1358
rect 158 752 161 778
rect 166 592 169 1258
rect 150 352 153 508
rect 118 72 121 278
rect 150 142 153 158
rect 174 62 177 208
rect 190 152 193 1658
rect 206 1542 209 1728
rect 214 1432 217 1908
rect 214 692 217 1428
rect 230 1042 233 1988
rect 278 1092 281 1578
rect 294 672 297 1558
rect 302 1272 305 1808
rect 310 1768 318 1771
rect 302 1082 305 1268
rect 310 762 313 1768
rect 350 1662 353 1858
rect 350 1252 353 1658
rect 382 1552 385 1838
rect 374 1452 377 1458
rect 382 1262 385 1548
rect 334 842 337 858
rect 342 852 345 968
rect 330 758 334 761
rect 314 738 318 741
rect 350 692 353 1248
rect 338 668 342 671
rect 282 658 286 661
rect 294 471 297 668
rect 350 662 353 688
rect 294 468 302 471
rect 330 318 337 321
rect 194 148 201 151
rect 198 62 201 148
rect 334 92 337 318
rect 358 82 361 1238
rect 382 832 385 1258
rect 398 1112 401 1598
rect 414 1351 417 1948
rect 410 1348 417 1351
rect 378 658 382 661
rect 390 352 393 1018
rect 422 982 425 1648
rect 430 1462 433 1578
rect 410 668 414 671
rect 406 452 409 658
rect 430 582 433 1458
rect 438 1132 441 2248
rect 758 2242 761 2308
rect 902 2278 910 2281
rect 902 2232 905 2278
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 494 2203 496 2207
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 494 2003 496 2007
rect 462 1352 465 1748
rect 446 572 449 728
rect 454 712 457 1348
rect 462 722 465 1348
rect 470 1302 473 1858
rect 502 1812 505 2018
rect 518 1942 521 1948
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 494 1803 496 1807
rect 510 1712 513 1788
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 494 1603 496 1607
rect 566 1502 569 1958
rect 574 1862 577 2218
rect 578 1858 582 1861
rect 478 1452 481 1458
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 494 1403 496 1407
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 490 668 494 671
rect 458 658 462 661
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 458 558 462 561
rect 462 532 465 548
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 502 362 505 718
rect 430 192 433 358
rect 510 352 513 808
rect 526 352 529 788
rect 534 672 537 678
rect 562 638 566 641
rect 574 502 577 1498
rect 582 1342 585 1618
rect 582 682 585 1338
rect 590 1032 593 2018
rect 598 1722 601 2128
rect 634 1948 638 1951
rect 606 1772 609 1948
rect 598 1382 601 1718
rect 598 812 601 1378
rect 606 1152 609 1768
rect 638 1742 641 1928
rect 646 1602 649 1958
rect 654 1402 657 1938
rect 662 1802 665 1848
rect 646 1252 649 1358
rect 582 452 585 658
rect 602 638 606 641
rect 590 582 593 608
rect 614 542 617 578
rect 630 542 633 688
rect 638 612 641 1188
rect 662 1151 665 1798
rect 670 1488 678 1491
rect 670 1222 673 1488
rect 686 1302 689 1948
rect 694 1662 697 2198
rect 746 2128 753 2131
rect 702 1942 705 1948
rect 718 1382 721 1858
rect 734 1492 737 2088
rect 750 1992 753 2128
rect 742 1512 745 1868
rect 790 1722 793 1738
rect 726 1252 729 1398
rect 670 1212 673 1218
rect 662 1148 670 1151
rect 646 872 649 908
rect 646 862 649 868
rect 650 668 654 671
rect 606 352 609 438
rect 670 362 673 1148
rect 682 1058 686 1061
rect 678 942 681 948
rect 694 842 697 1188
rect 686 592 689 688
rect 694 352 697 358
rect 702 282 705 828
rect 598 242 601 248
rect 710 212 713 1108
rect 718 832 721 1198
rect 726 802 729 1048
rect 734 532 737 1488
rect 742 1222 745 1508
rect 798 1352 801 1948
rect 802 1198 809 1201
rect 786 1148 790 1151
rect 750 662 753 728
rect 758 672 761 708
rect 790 662 793 1098
rect 806 992 809 1198
rect 814 1152 817 1568
rect 822 1312 825 1958
rect 854 1822 857 2018
rect 838 1648 846 1651
rect 838 1322 841 1648
rect 854 1542 857 1818
rect 862 1372 865 1748
rect 822 1262 825 1298
rect 822 1002 825 1118
rect 838 992 841 1318
rect 762 658 766 661
rect 742 562 745 658
rect 790 642 793 658
rect 798 292 801 798
rect 806 262 809 918
rect 834 678 838 681
rect 818 658 822 661
rect 846 462 849 1068
rect 854 952 857 1348
rect 862 1062 865 1248
rect 870 1162 873 1818
rect 918 1662 921 2398
rect 974 2302 977 2318
rect 984 2303 986 2307
rect 990 2303 993 2307
rect 998 2303 1000 2307
rect 1106 2248 1113 2251
rect 942 2112 945 2158
rect 1006 2152 1009 2168
rect 950 1952 953 1958
rect 878 1442 881 1638
rect 870 902 873 1158
rect 878 872 881 1218
rect 886 622 889 1408
rect 894 1032 897 1358
rect 942 1262 945 1668
rect 846 451 849 458
rect 846 448 854 451
rect 862 402 865 548
rect 878 222 881 548
rect 886 412 889 618
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 886 192 889 378
rect 902 192 905 1078
rect 926 1052 929 1258
rect 950 1162 953 1928
rect 966 1752 969 2118
rect 984 2103 986 2107
rect 990 2103 993 2107
rect 998 2103 1000 2107
rect 974 1992 977 2058
rect 926 862 929 1048
rect 914 858 918 861
rect 910 612 913 818
rect 934 671 937 918
rect 942 702 945 1078
rect 958 1002 961 1648
rect 974 1442 977 1988
rect 984 1903 986 1907
rect 990 1903 993 1907
rect 998 1903 1000 1907
rect 984 1703 986 1707
rect 990 1703 993 1707
rect 998 1703 1000 1707
rect 984 1503 986 1507
rect 990 1503 993 1507
rect 998 1503 1000 1507
rect 1006 1362 1009 2148
rect 1054 2062 1057 2238
rect 1014 1432 1017 1748
rect 1022 1742 1025 2038
rect 974 1272 977 1318
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 1014 1271 1017 1378
rect 1014 1268 1022 1271
rect 966 1142 969 1148
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 966 972 969 998
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 934 668 942 671
rect 910 472 913 608
rect 918 562 921 608
rect 958 392 961 868
rect 1006 732 1009 1228
rect 1038 1132 1041 1698
rect 1054 1542 1057 1808
rect 974 522 977 708
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 1006 682 1009 708
rect 1014 602 1017 938
rect 1030 882 1033 938
rect 1030 752 1033 878
rect 1046 852 1049 1148
rect 1054 742 1057 1538
rect 1062 1172 1065 2198
rect 1070 1192 1073 1838
rect 1078 1662 1081 2118
rect 1062 922 1065 1018
rect 1054 702 1057 738
rect 1062 682 1065 918
rect 1070 542 1073 1188
rect 1078 1122 1081 1658
rect 1110 1392 1113 2248
rect 1150 2222 1153 2238
rect 1190 2222 1193 2338
rect 1222 2272 1225 2338
rect 1358 2272 1361 2298
rect 1546 2268 1550 2271
rect 1154 2218 1161 2221
rect 1130 2058 1134 2061
rect 1158 2032 1161 2218
rect 1122 2018 1126 2021
rect 1178 1968 1185 1971
rect 1174 1832 1177 1868
rect 1078 752 1081 1098
rect 974 172 977 518
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 1006 282 1009 308
rect 1030 162 1033 438
rect 1078 342 1081 638
rect 1034 158 1038 161
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect 1014 102 1017 148
rect 1086 62 1089 1058
rect 1098 1048 1102 1051
rect 1110 762 1113 888
rect 1118 852 1121 958
rect 1142 952 1145 1558
rect 1150 1182 1153 1268
rect 1158 1182 1161 1198
rect 1142 912 1145 948
rect 1094 758 1102 761
rect 1094 161 1097 758
rect 1102 652 1105 658
rect 1102 282 1105 568
rect 1110 462 1113 758
rect 1150 692 1153 1168
rect 1158 902 1161 1178
rect 1166 912 1169 1638
rect 1174 1592 1177 1828
rect 1182 1532 1185 1968
rect 1182 1102 1185 1128
rect 1190 1062 1193 2218
rect 1222 1542 1225 2268
rect 1246 2252 1249 2258
rect 1446 2252 1449 2258
rect 1310 2132 1313 2148
rect 1262 1752 1265 1968
rect 1302 1942 1305 2028
rect 1302 1892 1305 1938
rect 1190 1032 1193 1058
rect 1210 1038 1214 1041
rect 1182 992 1185 1028
rect 1158 732 1161 898
rect 1166 782 1169 908
rect 1174 842 1177 958
rect 1222 892 1225 1538
rect 1230 1512 1233 1738
rect 1238 1652 1241 1718
rect 1238 1062 1241 1358
rect 1254 1002 1257 1458
rect 1302 1452 1305 1888
rect 1310 1732 1313 1848
rect 1326 1842 1329 1958
rect 1342 1862 1345 2228
rect 1398 1978 1406 1981
rect 1310 1372 1313 1628
rect 1278 1122 1281 1248
rect 1302 1012 1305 1328
rect 1318 1062 1321 1728
rect 1326 1602 1329 1838
rect 1326 1062 1329 1588
rect 1310 1052 1313 1058
rect 1222 782 1225 888
rect 1166 732 1169 748
rect 1158 692 1161 698
rect 1142 652 1145 658
rect 1142 572 1145 578
rect 1150 372 1153 688
rect 1166 652 1169 708
rect 1198 562 1201 778
rect 1238 732 1241 858
rect 1254 852 1257 858
rect 1278 682 1281 878
rect 1198 532 1201 558
rect 1182 528 1190 531
rect 1182 432 1185 528
rect 1206 412 1209 648
rect 1142 352 1145 358
rect 1286 272 1289 928
rect 1294 872 1297 898
rect 1302 772 1305 1008
rect 1310 752 1313 1048
rect 1318 792 1321 1058
rect 1326 962 1329 1058
rect 1334 1052 1337 1748
rect 1342 1712 1345 1858
rect 1358 1142 1361 1468
rect 1374 1332 1377 1938
rect 1346 1038 1350 1041
rect 1358 942 1361 1138
rect 1334 812 1337 908
rect 1318 752 1321 768
rect 1294 728 1302 731
rect 1294 222 1297 728
rect 1358 422 1361 938
rect 1366 522 1369 748
rect 1374 662 1377 928
rect 1374 572 1377 658
rect 1318 282 1321 338
rect 1094 158 1102 161
rect 1126 141 1129 188
rect 1318 152 1321 278
rect 1382 242 1385 988
rect 1390 842 1393 1358
rect 1398 1242 1401 1978
rect 1438 1952 1441 2138
rect 1454 2082 1457 2118
rect 1406 1322 1409 1938
rect 1438 1922 1441 1938
rect 1446 1932 1449 1958
rect 1450 1928 1454 1931
rect 1486 1872 1489 2238
rect 1496 2203 1498 2207
rect 1502 2203 1505 2207
rect 1510 2203 1512 2207
rect 1496 2003 1498 2007
rect 1502 2003 1505 2007
rect 1510 2003 1512 2007
rect 1498 1868 1502 1871
rect 1542 1842 1545 1858
rect 1478 1762 1481 1828
rect 1496 1803 1498 1807
rect 1502 1803 1505 1807
rect 1510 1803 1512 1807
rect 1502 1762 1505 1768
rect 1550 1652 1553 1798
rect 1496 1603 1498 1607
rect 1502 1603 1505 1607
rect 1510 1603 1512 1607
rect 1398 1192 1401 1238
rect 1398 842 1401 1188
rect 1438 1082 1441 1558
rect 1478 1422 1481 1558
rect 1496 1403 1498 1407
rect 1502 1403 1505 1407
rect 1510 1403 1512 1407
rect 1496 1203 1498 1207
rect 1502 1203 1505 1207
rect 1510 1203 1512 1207
rect 1496 1003 1498 1007
rect 1502 1003 1505 1007
rect 1510 1003 1512 1007
rect 1390 722 1393 838
rect 1414 652 1417 878
rect 1498 848 1502 851
rect 1496 803 1498 807
rect 1502 803 1505 807
rect 1510 803 1512 807
rect 1518 742 1521 1338
rect 1558 1032 1561 1648
rect 1566 1392 1569 2348
rect 1806 2132 1809 2388
rect 2362 2348 2366 2351
rect 1694 2052 1697 2088
rect 1586 1848 1590 1851
rect 1598 1662 1601 1668
rect 1566 852 1569 1388
rect 1574 1302 1577 1348
rect 1606 1122 1609 1648
rect 1398 472 1401 578
rect 1438 512 1441 718
rect 1496 603 1498 607
rect 1502 603 1505 607
rect 1510 603 1512 607
rect 1518 542 1521 738
rect 1496 403 1498 407
rect 1502 403 1505 407
rect 1510 403 1512 407
rect 1414 272 1417 298
rect 1126 138 1134 141
rect 1374 102 1377 218
rect 1382 192 1385 238
rect 682 58 686 61
rect 1098 58 1102 61
rect 1398 61 1401 118
rect 1398 58 1406 61
rect 1422 22 1425 328
rect 1574 312 1577 948
rect 1598 882 1601 908
rect 1602 868 1606 871
rect 1598 462 1601 818
rect 1606 742 1609 748
rect 1614 652 1617 1268
rect 1638 1102 1641 1548
rect 1654 1052 1657 1958
rect 1670 1552 1673 1728
rect 1678 1662 1681 1668
rect 1670 1292 1673 1548
rect 1622 712 1625 848
rect 1646 768 1654 771
rect 1646 732 1649 768
rect 1430 242 1433 268
rect 1496 203 1498 207
rect 1502 203 1505 207
rect 1510 203 1512 207
rect 1438 62 1441 188
rect 1574 162 1577 308
rect 1598 212 1601 368
rect 1646 362 1649 378
rect 1654 262 1657 738
rect 1662 372 1665 1248
rect 1670 432 1673 1288
rect 1694 1102 1697 2048
rect 1702 1462 1705 1738
rect 1710 1452 1713 1848
rect 1718 1152 1721 1568
rect 1678 552 1681 778
rect 1686 682 1689 1098
rect 1694 752 1697 1098
rect 1694 732 1697 738
rect 1702 662 1705 1108
rect 1726 962 1729 1608
rect 1742 1111 1745 2128
rect 1750 1751 1753 1868
rect 1814 1832 1817 2308
rect 1830 2252 1833 2348
rect 2210 2338 2217 2341
rect 2016 2303 2018 2307
rect 2022 2303 2025 2307
rect 2030 2303 2032 2307
rect 1822 2182 1825 2238
rect 1750 1748 1758 1751
rect 1766 1652 1769 1658
rect 1754 1648 1761 1651
rect 1758 1262 1761 1648
rect 1798 1232 1801 1658
rect 1814 1282 1817 1828
rect 1822 1782 1825 2178
rect 1830 1842 1833 2248
rect 1854 1861 1857 2148
rect 1902 2062 1905 2178
rect 1862 1882 1865 1968
rect 1850 1858 1857 1861
rect 1850 1838 1854 1841
rect 1742 1108 1750 1111
rect 1750 892 1753 938
rect 1714 868 1718 871
rect 1758 812 1761 1158
rect 1782 842 1785 968
rect 1734 662 1737 668
rect 1750 662 1753 808
rect 1814 352 1817 1278
rect 1830 1072 1833 1838
rect 1854 1742 1857 1778
rect 1846 1592 1849 1638
rect 1838 922 1841 1458
rect 1846 1022 1849 1588
rect 1854 1262 1857 1738
rect 1870 1332 1873 1908
rect 1878 1862 1881 1868
rect 1878 1402 1881 1858
rect 1902 1462 1905 2058
rect 1918 1942 1921 2138
rect 1926 2048 1934 2051
rect 1914 1928 1921 1931
rect 1918 1392 1921 1928
rect 1926 1712 1929 2048
rect 1878 1342 1881 1388
rect 1838 512 1841 758
rect 1846 752 1849 1018
rect 1846 492 1849 748
rect 1854 442 1857 1258
rect 1862 922 1865 1318
rect 1870 972 1873 1328
rect 1878 462 1881 1338
rect 1926 1242 1929 1708
rect 1934 1672 1937 1678
rect 1958 1632 1961 1738
rect 1910 1042 1913 1048
rect 1890 858 1897 861
rect 1862 302 1865 458
rect 1894 432 1897 858
rect 1906 658 1910 661
rect 1918 382 1921 1208
rect 1926 672 1929 838
rect 1942 752 1945 758
rect 1950 752 1953 1278
rect 1958 1212 1961 1628
rect 1958 982 1961 1158
rect 1966 1062 1969 1748
rect 1974 1362 1977 2258
rect 2016 2103 2018 2107
rect 2022 2103 2025 2107
rect 2030 2103 2032 2107
rect 1998 1862 2001 2058
rect 2006 1742 2009 1948
rect 2016 1903 2018 1907
rect 2022 1903 2025 1907
rect 2030 1903 2032 1907
rect 2094 1832 2097 1858
rect 2102 1792 2105 1908
rect 2098 1768 2102 1771
rect 2106 1738 2110 1741
rect 2016 1703 2018 1707
rect 2022 1703 2025 1707
rect 2030 1703 2032 1707
rect 1986 1518 1993 1521
rect 1990 1262 1993 1518
rect 2016 1503 2018 1507
rect 2022 1503 2025 1507
rect 2030 1503 2032 1507
rect 2022 1462 2025 1468
rect 2016 1303 2018 1307
rect 2022 1303 2025 1307
rect 2030 1303 2032 1307
rect 1974 772 1977 1148
rect 2016 1103 2018 1107
rect 2022 1103 2025 1107
rect 2030 1103 2032 1107
rect 1950 452 1953 658
rect 1982 362 1985 1088
rect 2046 1062 2049 1738
rect 2110 1652 2113 1718
rect 2010 1058 2014 1061
rect 2082 1058 2086 1061
rect 2016 903 2018 907
rect 2022 903 2025 907
rect 2030 903 2032 907
rect 2046 741 2049 1058
rect 2078 832 2081 1038
rect 2094 1012 2097 1578
rect 2066 748 2070 751
rect 2046 738 2054 741
rect 1994 658 1998 661
rect 2006 532 2009 738
rect 2016 703 2018 707
rect 2022 703 2025 707
rect 2030 703 2032 707
rect 2038 672 2041 698
rect 2054 662 2057 728
rect 2016 503 2018 507
rect 2022 503 2025 507
rect 2030 503 2032 507
rect 2086 332 2089 838
rect 2110 812 2113 1648
rect 2118 1252 2121 2188
rect 2126 1412 2129 2168
rect 2158 1952 2161 2258
rect 2182 1862 2185 1918
rect 2174 1858 2182 1861
rect 2162 1748 2166 1751
rect 2138 1458 2142 1461
rect 2126 672 2129 1018
rect 2142 652 2145 668
rect 2016 303 2018 307
rect 2022 303 2025 307
rect 2030 303 2032 307
rect 1610 258 1614 261
rect 1654 22 1657 258
rect 1966 72 1969 238
rect 2150 182 2153 1238
rect 2158 1052 2161 1058
rect 2158 152 2161 998
rect 2166 682 2169 1578
rect 2166 272 2169 678
rect 2174 472 2177 1858
rect 2198 1852 2201 1958
rect 2182 1042 2185 1848
rect 2198 1271 2201 1848
rect 2214 1482 2217 2338
rect 2222 1672 2225 1988
rect 2222 1462 2225 1668
rect 2198 1268 2206 1271
rect 2206 1252 2209 1268
rect 2198 342 2201 1038
rect 2206 842 2209 1248
rect 2222 1042 2225 1458
rect 2230 362 2233 1798
rect 2238 682 2241 2338
rect 2262 2252 2265 2258
rect 2246 1082 2249 1538
rect 2254 1182 2257 1748
rect 2286 1461 2289 2248
rect 2286 1458 2294 1461
rect 2246 662 2249 678
rect 2254 462 2257 1178
rect 2286 682 2289 1318
rect 2294 1092 2297 1458
rect 2302 1132 2305 2338
rect 2298 1048 2302 1051
rect 2302 582 2305 1038
rect 2310 862 2313 2348
rect 2318 1362 2321 1908
rect 2326 1351 2329 1948
rect 2318 1348 2329 1351
rect 2318 1042 2321 1348
rect 2314 678 2321 681
rect 2318 552 2321 678
rect 2326 582 2329 1188
rect 2334 942 2337 2318
rect 2342 1542 2345 1868
rect 2350 1752 2353 2228
rect 2350 952 2353 1748
rect 2358 1452 2361 2278
rect 2374 2132 2377 2158
rect 2342 462 2345 488
rect 2366 272 2369 1978
rect 2374 1622 2377 1758
rect 2374 1072 2377 1608
rect 2382 1462 2385 2358
rect 2390 1612 2393 2318
rect 2414 1852 2417 2348
rect 2446 2242 2449 2318
rect 2446 2032 2449 2238
rect 2422 1841 2425 1958
rect 2414 1838 2425 1841
rect 2382 612 2385 1458
rect 2390 1442 2393 1598
rect 2390 1272 2393 1428
rect 2390 1262 2393 1268
rect 2398 1162 2401 1818
rect 2390 1158 2398 1161
rect 2390 452 2393 1158
rect 2398 362 2401 738
rect 2406 242 2409 1718
rect 2414 1602 2417 1838
rect 2414 1282 2417 1498
rect 2414 1122 2417 1268
rect 2414 872 2417 1088
rect 2422 542 2425 1608
rect 2430 1152 2433 1488
rect 2438 1072 2441 1698
rect 2446 1092 2449 1938
rect 2434 958 2441 961
rect 2438 952 2441 958
rect 2430 522 2433 948
rect 2446 142 2449 1078
rect 2454 662 2457 2188
rect 2462 1942 2465 2338
rect 2474 2258 2478 2261
rect 2016 103 2018 107
rect 2022 103 2025 107
rect 2030 103 2032 107
rect 2038 22 2041 98
rect 2462 92 2465 1198
rect 2470 872 2473 1268
rect 2478 1062 2481 1738
rect 2486 1552 2489 1818
rect 2486 1252 2489 1548
rect 2470 72 2473 868
rect 2486 292 2489 1238
rect 2494 1102 2497 2088
rect 2502 1071 2505 1498
rect 2494 1068 2505 1071
rect 2494 762 2497 1068
rect 2510 1061 2513 1758
rect 2502 1058 2513 1061
rect 2502 362 2505 1058
rect 2510 692 2513 878
rect 2518 252 2521 1968
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
rect 1496 3 1498 7
rect 1502 3 1505 7
rect 1510 3 1512 7
<< m5contact >>
rect 482 2403 486 2407
rect 489 2403 490 2407
rect 490 2403 493 2407
rect 1498 2403 1502 2407
rect 1505 2403 1506 2407
rect 1506 2403 1509 2407
rect 54 2338 58 2342
rect 46 648 50 652
rect 398 2258 402 2262
rect 590 2258 594 2262
rect 438 2248 442 2252
rect 126 748 130 752
rect 190 1668 194 1672
rect 158 778 162 782
rect 374 1448 378 1452
rect 334 838 338 842
rect 334 758 338 762
rect 318 738 322 742
rect 350 688 354 692
rect 342 668 346 672
rect 286 658 290 662
rect 374 658 378 662
rect 406 668 410 672
rect 758 2238 762 2242
rect 482 2203 486 2207
rect 489 2203 490 2207
rect 490 2203 493 2207
rect 482 2003 486 2007
rect 489 2003 490 2007
rect 490 2003 493 2007
rect 518 1938 522 1942
rect 482 1803 486 1807
rect 489 1803 490 1807
rect 490 1803 493 1807
rect 482 1603 486 1607
rect 489 1603 490 1607
rect 490 1603 493 1607
rect 598 2128 602 2132
rect 582 1858 586 1862
rect 478 1458 482 1462
rect 482 1403 486 1407
rect 489 1403 490 1407
rect 490 1403 493 1407
rect 482 1203 486 1207
rect 489 1203 490 1207
rect 490 1203 493 1207
rect 482 1003 486 1007
rect 489 1003 490 1007
rect 490 1003 493 1007
rect 482 803 486 807
rect 489 803 490 807
rect 490 803 493 807
rect 494 668 498 672
rect 462 658 466 662
rect 482 603 486 607
rect 489 603 490 607
rect 490 603 493 607
rect 454 558 458 562
rect 482 403 486 407
rect 489 403 490 407
rect 490 403 493 407
rect 534 678 538 682
rect 566 638 570 642
rect 638 1948 642 1952
rect 606 1768 610 1772
rect 606 638 610 642
rect 590 578 594 582
rect 702 1948 706 1952
rect 854 2018 858 2022
rect 822 1958 826 1962
rect 742 1868 746 1872
rect 646 868 650 872
rect 646 668 650 672
rect 686 1058 690 1062
rect 678 938 682 942
rect 694 358 698 362
rect 598 238 602 242
rect 790 1148 794 1152
rect 750 728 754 732
rect 766 658 770 662
rect 830 678 834 682
rect 822 658 826 662
rect 1222 2338 1226 2342
rect 986 2303 990 2307
rect 993 2303 994 2307
rect 994 2303 997 2307
rect 950 1958 954 1962
rect 806 258 810 262
rect 482 203 486 207
rect 489 203 490 207
rect 490 203 493 207
rect 986 2103 990 2107
rect 993 2103 994 2107
rect 994 2103 997 2107
rect 942 1078 946 1082
rect 926 1048 930 1052
rect 918 858 922 862
rect 986 1903 990 1907
rect 993 1903 994 1907
rect 994 1903 997 1907
rect 986 1703 990 1707
rect 993 1703 994 1707
rect 994 1703 997 1707
rect 986 1503 990 1507
rect 993 1503 994 1507
rect 994 1503 997 1507
rect 986 1303 990 1307
rect 993 1303 994 1307
rect 994 1303 997 1307
rect 966 1148 970 1152
rect 986 1103 990 1107
rect 993 1103 994 1107
rect 994 1103 997 1107
rect 986 903 990 907
rect 993 903 994 907
rect 994 903 997 907
rect 1006 728 1010 732
rect 986 703 990 707
rect 993 703 994 707
rect 994 703 997 707
rect 1078 1658 1082 1662
rect 1054 738 1058 742
rect 1150 2238 1154 2242
rect 1358 2268 1362 2272
rect 1550 2268 1554 2272
rect 1134 2058 1138 2062
rect 1118 2018 1122 2022
rect 1174 1828 1178 1832
rect 986 503 990 507
rect 993 503 994 507
rect 994 503 997 507
rect 986 303 990 307
rect 993 303 994 307
rect 994 303 997 307
rect 1030 158 1034 162
rect 986 103 990 107
rect 993 103 994 107
rect 994 103 997 107
rect 1102 1048 1106 1052
rect 1142 948 1146 952
rect 1118 848 1122 852
rect 1110 758 1114 762
rect 1102 658 1106 662
rect 1246 2248 1250 2252
rect 1446 2248 1450 2252
rect 1310 2128 1314 2132
rect 1302 1938 1306 1942
rect 1190 1058 1194 1062
rect 1214 1038 1218 1042
rect 1238 1648 1242 1652
rect 1342 1858 1346 1862
rect 1334 1748 1338 1752
rect 1310 1058 1314 1062
rect 1318 1058 1322 1062
rect 1254 858 1258 862
rect 1222 778 1226 782
rect 1158 698 1162 702
rect 1142 648 1146 652
rect 1142 578 1146 582
rect 1238 728 1242 732
rect 1198 558 1202 562
rect 1150 368 1154 372
rect 1142 348 1146 352
rect 1294 868 1298 872
rect 1350 1038 1354 1042
rect 1358 938 1362 942
rect 1318 748 1322 752
rect 1374 658 1378 662
rect 1446 1958 1450 1962
rect 1454 1928 1458 1932
rect 1498 2203 1502 2207
rect 1505 2203 1506 2207
rect 1506 2203 1509 2207
rect 1498 2003 1502 2007
rect 1505 2003 1506 2007
rect 1506 2003 1509 2007
rect 1502 1868 1506 1872
rect 1542 1838 1546 1842
rect 1498 1803 1502 1807
rect 1505 1803 1506 1807
rect 1506 1803 1509 1807
rect 1502 1768 1506 1772
rect 1498 1603 1502 1607
rect 1505 1603 1506 1607
rect 1506 1603 1509 1607
rect 1498 1403 1502 1407
rect 1505 1403 1506 1407
rect 1506 1403 1509 1407
rect 1498 1203 1502 1207
rect 1505 1203 1506 1207
rect 1506 1203 1509 1207
rect 1438 1078 1442 1082
rect 1498 1003 1502 1007
rect 1505 1003 1506 1007
rect 1506 1003 1509 1007
rect 1390 838 1394 842
rect 1494 848 1498 852
rect 1498 803 1502 807
rect 1505 803 1506 807
rect 1506 803 1509 807
rect 2366 2348 2370 2352
rect 1590 1848 1594 1852
rect 1598 1668 1602 1672
rect 1498 603 1502 607
rect 1505 603 1506 607
rect 1506 603 1509 607
rect 1498 403 1502 407
rect 1505 403 1506 407
rect 1506 403 1509 407
rect 1382 238 1386 242
rect 678 58 682 62
rect 1094 58 1098 62
rect 1606 868 1610 872
rect 1606 748 1610 752
rect 1678 1658 1682 1662
rect 1646 728 1650 732
rect 1598 368 1602 372
rect 1498 203 1502 207
rect 1505 203 1506 207
rect 1506 203 1509 207
rect 1694 738 1698 742
rect 2018 2303 2022 2307
rect 2025 2303 2026 2307
rect 2026 2303 2029 2307
rect 1766 1658 1770 1662
rect 1750 1648 1754 1652
rect 1902 2058 1906 2062
rect 1846 1838 1850 1842
rect 1718 868 1722 872
rect 1734 668 1738 672
rect 1854 1738 1858 1742
rect 1878 1868 1882 1872
rect 1910 1928 1914 1932
rect 1878 1388 1882 1392
rect 1918 1388 1922 1392
rect 1934 1668 1938 1672
rect 1910 1038 1914 1042
rect 1902 658 1906 662
rect 2018 2103 2022 2107
rect 2025 2103 2026 2107
rect 2026 2103 2029 2107
rect 2018 1903 2022 1907
rect 2025 1903 2026 1907
rect 2026 1903 2029 1907
rect 2094 1828 2098 1832
rect 2094 1768 2098 1772
rect 2102 1738 2106 1742
rect 2018 1703 2022 1707
rect 2025 1703 2026 1707
rect 2026 1703 2029 1707
rect 2018 1503 2022 1507
rect 2025 1503 2026 1507
rect 2026 1503 2029 1507
rect 2022 1458 2026 1462
rect 2018 1303 2022 1307
rect 2025 1303 2026 1307
rect 2026 1303 2029 1307
rect 2018 1103 2022 1107
rect 2025 1103 2026 1107
rect 2026 1103 2029 1107
rect 1942 748 1946 752
rect 2014 1058 2018 1062
rect 2046 1058 2050 1062
rect 2086 1058 2090 1062
rect 2018 903 2022 907
rect 2025 903 2026 907
rect 2026 903 2029 907
rect 2062 748 2066 752
rect 1998 658 2002 662
rect 2054 728 2058 732
rect 2018 703 2022 707
rect 2025 703 2026 707
rect 2026 703 2029 707
rect 2038 668 2042 672
rect 2018 503 2022 507
rect 2025 503 2026 507
rect 2026 503 2029 507
rect 2158 1748 2162 1752
rect 2134 1458 2138 1462
rect 2018 303 2022 307
rect 2025 303 2026 307
rect 2026 303 2029 307
rect 1614 258 1618 262
rect 1574 158 1578 162
rect 2158 1058 2162 1062
rect 2198 1848 2202 1852
rect 2262 2248 2266 2252
rect 2246 658 2250 662
rect 2294 1048 2298 1052
rect 2374 2128 2378 2132
rect 2374 1608 2378 1612
rect 2390 1608 2394 1612
rect 2390 1598 2394 1602
rect 2414 1598 2418 1602
rect 2414 1268 2418 1272
rect 2438 948 2442 952
rect 2478 2258 2482 2262
rect 2018 103 2022 107
rect 2025 103 2026 107
rect 2026 103 2029 107
rect 2486 1238 2490 1242
rect 482 3 486 7
rect 489 3 490 7
rect 490 3 493 7
rect 1498 3 1502 7
rect 1505 3 1506 7
rect 1506 3 1509 7
<< metal5 >>
rect 486 2403 489 2407
rect 485 2402 490 2403
rect 495 2402 496 2407
rect 1502 2403 1505 2407
rect 1501 2402 1506 2403
rect 1511 2402 1512 2407
rect 2366 2342 2369 2348
rect 58 2338 1222 2341
rect 990 2303 993 2307
rect 989 2302 994 2303
rect 999 2302 1000 2307
rect 2022 2303 2025 2307
rect 2021 2302 2026 2303
rect 2031 2302 2032 2307
rect 1362 2268 1550 2271
rect 402 2258 590 2261
rect 2478 2252 2481 2258
rect 442 2248 1246 2251
rect 1450 2248 2262 2251
rect 762 2238 1150 2241
rect 486 2203 489 2207
rect 485 2202 490 2203
rect 495 2202 496 2207
rect 1502 2203 1505 2207
rect 1501 2202 1506 2203
rect 1511 2202 1512 2207
rect 602 2128 1310 2131
rect 1314 2128 2374 2131
rect 990 2103 993 2107
rect 989 2102 994 2103
rect 999 2102 1000 2107
rect 2022 2103 2025 2107
rect 2021 2102 2026 2103
rect 2031 2102 2032 2107
rect 1138 2058 1902 2061
rect 858 2018 1118 2021
rect 486 2003 489 2007
rect 485 2002 490 2003
rect 495 2002 496 2007
rect 1502 2003 1505 2007
rect 1501 2002 1506 2003
rect 1511 2002 1512 2007
rect 826 1958 950 1961
rect 954 1958 1446 1961
rect 642 1948 702 1951
rect 522 1938 1302 1941
rect 1458 1928 1910 1931
rect 990 1903 993 1907
rect 989 1902 994 1903
rect 999 1902 1000 1907
rect 2022 1903 2025 1907
rect 2021 1902 2026 1903
rect 2031 1902 2032 1907
rect 746 1868 1502 1871
rect 1506 1868 1878 1871
rect 586 1858 1342 1861
rect 1594 1848 2198 1851
rect 1546 1838 1846 1841
rect 1178 1828 2094 1831
rect 486 1803 489 1807
rect 485 1802 490 1803
rect 495 1802 496 1807
rect 1502 1803 1505 1807
rect 1501 1802 1506 1803
rect 1511 1802 1512 1807
rect 610 1768 1502 1771
rect 1506 1768 2094 1771
rect 1338 1748 2158 1751
rect 1858 1738 2102 1741
rect 990 1703 993 1707
rect 989 1702 994 1703
rect 999 1702 1000 1707
rect 2022 1703 2025 1707
rect 2021 1702 2026 1703
rect 2031 1702 2032 1707
rect 1602 1668 1934 1671
rect 190 1661 193 1668
rect 190 1658 1078 1661
rect 1682 1658 1766 1661
rect 1242 1648 1750 1651
rect 2378 1608 2390 1611
rect 486 1603 489 1607
rect 485 1602 490 1603
rect 495 1602 496 1607
rect 1502 1603 1505 1607
rect 1501 1602 1506 1603
rect 1511 1602 1512 1607
rect 2394 1598 2414 1601
rect 990 1503 993 1507
rect 989 1502 994 1503
rect 999 1502 1000 1507
rect 2022 1503 2025 1507
rect 2021 1502 2026 1503
rect 2031 1502 2032 1507
rect 2026 1458 2134 1461
rect 478 1451 481 1458
rect 378 1448 481 1451
rect 486 1403 489 1407
rect 485 1402 490 1403
rect 495 1402 496 1407
rect 1502 1403 1505 1407
rect 1501 1402 1506 1403
rect 1511 1402 1512 1407
rect 1882 1388 1918 1391
rect 990 1303 993 1307
rect 989 1302 994 1303
rect 999 1302 1000 1307
rect 2022 1303 2025 1307
rect 2021 1302 2026 1303
rect 2031 1302 2032 1307
rect 2370 1268 2414 1271
rect 2482 1238 2486 1241
rect 486 1203 489 1207
rect 485 1202 490 1203
rect 495 1202 496 1207
rect 1502 1203 1505 1207
rect 1501 1202 1506 1203
rect 1511 1202 1512 1207
rect 794 1148 966 1151
rect 990 1103 993 1107
rect 989 1102 994 1103
rect 999 1102 1000 1107
rect 2022 1103 2025 1107
rect 2021 1102 2026 1103
rect 2031 1102 2032 1107
rect 946 1078 1438 1081
rect 690 1058 1190 1061
rect 1322 1058 2014 1061
rect 2018 1058 2046 1061
rect 2090 1058 2158 1061
rect 930 1048 1102 1051
rect 1310 1051 1313 1058
rect 1106 1048 1313 1051
rect 1910 1048 2294 1051
rect 1910 1042 1913 1048
rect 1218 1038 1350 1041
rect 486 1003 489 1007
rect 485 1002 490 1003
rect 495 1002 496 1007
rect 1502 1003 1505 1007
rect 1501 1002 1506 1003
rect 1511 1002 1512 1007
rect 1146 948 2438 951
rect 682 938 1358 941
rect 990 903 993 907
rect 989 902 994 903
rect 999 902 1000 907
rect 2022 903 2025 907
rect 2021 902 2026 903
rect 2031 902 2032 907
rect 650 868 1294 871
rect 1610 868 1718 871
rect 922 858 1254 861
rect 1122 848 1494 851
rect 338 838 1390 841
rect 486 803 489 807
rect 485 802 490 803
rect 495 802 496 807
rect 1502 803 1505 807
rect 1501 802 1506 803
rect 1511 802 1512 807
rect 162 778 1222 781
rect 338 758 1110 761
rect 130 748 1318 751
rect 1946 748 2062 751
rect 322 738 1054 741
rect 1606 741 1609 748
rect 1606 738 1694 741
rect 754 728 1006 731
rect 1010 728 1238 731
rect 1242 728 1646 731
rect 1650 728 2054 731
rect 990 703 993 707
rect 989 702 994 703
rect 999 702 1000 707
rect 2022 703 2025 707
rect 2021 702 2026 703
rect 2031 702 2032 707
rect 1158 691 1161 698
rect 354 688 1161 691
rect 538 678 830 681
rect 834 678 841 681
rect 346 668 406 671
rect 498 668 646 671
rect 1738 668 2038 671
rect 290 658 374 661
rect 466 658 766 661
rect 826 658 1102 661
rect 1378 658 1902 661
rect 2002 658 2246 661
rect 50 648 1142 651
rect 570 638 606 641
rect 486 603 489 607
rect 485 602 490 603
rect 495 602 496 607
rect 1502 603 1505 607
rect 1501 602 1506 603
rect 1511 602 1512 607
rect 594 578 1142 581
rect 458 558 1198 561
rect 990 503 993 507
rect 989 502 994 503
rect 999 502 1000 507
rect 2022 503 2025 507
rect 2021 502 2026 503
rect 2031 502 2032 507
rect 486 403 489 407
rect 485 402 490 403
rect 495 402 496 407
rect 1502 403 1505 407
rect 1501 402 1506 403
rect 1511 402 1512 407
rect 1154 368 1598 371
rect 694 351 697 358
rect 694 348 1142 351
rect 990 303 993 307
rect 989 302 994 303
rect 999 302 1000 307
rect 2022 303 2025 307
rect 2021 302 2026 303
rect 2031 302 2032 307
rect 810 258 1614 261
rect 602 238 1382 241
rect 486 203 489 207
rect 485 202 490 203
rect 495 202 496 207
rect 1502 203 1505 207
rect 1501 202 1506 203
rect 1511 202 1512 207
rect 1034 158 1574 161
rect 990 103 993 107
rect 989 102 994 103
rect 999 102 1000 107
rect 2022 103 2025 107
rect 2021 102 2026 103
rect 2031 102 2032 107
rect 682 58 1094 61
rect 486 3 489 7
rect 485 2 490 3
rect 495 2 496 7
rect 1502 3 1505 7
rect 1501 2 1506 3
rect 1511 2 1512 7
<< m6contact >>
rect 480 2403 482 2407
rect 482 2403 485 2407
rect 490 2403 493 2407
rect 493 2403 495 2407
rect 480 2402 485 2403
rect 490 2402 495 2403
rect 1496 2403 1498 2407
rect 1498 2403 1501 2407
rect 1506 2403 1509 2407
rect 1509 2403 1511 2407
rect 1496 2402 1501 2403
rect 1506 2402 1511 2403
rect 2365 2337 2370 2342
rect 984 2303 986 2307
rect 986 2303 989 2307
rect 994 2303 997 2307
rect 997 2303 999 2307
rect 984 2302 989 2303
rect 994 2302 999 2303
rect 2016 2303 2018 2307
rect 2018 2303 2021 2307
rect 2026 2303 2029 2307
rect 2029 2303 2031 2307
rect 2016 2302 2021 2303
rect 2026 2302 2031 2303
rect 2477 2247 2482 2252
rect 480 2203 482 2207
rect 482 2203 485 2207
rect 490 2203 493 2207
rect 493 2203 495 2207
rect 480 2202 485 2203
rect 490 2202 495 2203
rect 1496 2203 1498 2207
rect 1498 2203 1501 2207
rect 1506 2203 1509 2207
rect 1509 2203 1511 2207
rect 1496 2202 1501 2203
rect 1506 2202 1511 2203
rect 984 2103 986 2107
rect 986 2103 989 2107
rect 994 2103 997 2107
rect 997 2103 999 2107
rect 984 2102 989 2103
rect 994 2102 999 2103
rect 2016 2103 2018 2107
rect 2018 2103 2021 2107
rect 2026 2103 2029 2107
rect 2029 2103 2031 2107
rect 2016 2102 2021 2103
rect 2026 2102 2031 2103
rect 480 2003 482 2007
rect 482 2003 485 2007
rect 490 2003 493 2007
rect 493 2003 495 2007
rect 480 2002 485 2003
rect 490 2002 495 2003
rect 1496 2003 1498 2007
rect 1498 2003 1501 2007
rect 1506 2003 1509 2007
rect 1509 2003 1511 2007
rect 1496 2002 1501 2003
rect 1506 2002 1511 2003
rect 984 1903 986 1907
rect 986 1903 989 1907
rect 994 1903 997 1907
rect 997 1903 999 1907
rect 984 1902 989 1903
rect 994 1902 999 1903
rect 2016 1903 2018 1907
rect 2018 1903 2021 1907
rect 2026 1903 2029 1907
rect 2029 1903 2031 1907
rect 2016 1902 2021 1903
rect 2026 1902 2031 1903
rect 480 1803 482 1807
rect 482 1803 485 1807
rect 490 1803 493 1807
rect 493 1803 495 1807
rect 480 1802 485 1803
rect 490 1802 495 1803
rect 1496 1803 1498 1807
rect 1498 1803 1501 1807
rect 1506 1803 1509 1807
rect 1509 1803 1511 1807
rect 1496 1802 1501 1803
rect 1506 1802 1511 1803
rect 984 1703 986 1707
rect 986 1703 989 1707
rect 994 1703 997 1707
rect 997 1703 999 1707
rect 984 1702 989 1703
rect 994 1702 999 1703
rect 2016 1703 2018 1707
rect 2018 1703 2021 1707
rect 2026 1703 2029 1707
rect 2029 1703 2031 1707
rect 2016 1702 2021 1703
rect 2026 1702 2031 1703
rect 480 1603 482 1607
rect 482 1603 485 1607
rect 490 1603 493 1607
rect 493 1603 495 1607
rect 480 1602 485 1603
rect 490 1602 495 1603
rect 1496 1603 1498 1607
rect 1498 1603 1501 1607
rect 1506 1603 1509 1607
rect 1509 1603 1511 1607
rect 1496 1602 1501 1603
rect 1506 1602 1511 1603
rect 984 1503 986 1507
rect 986 1503 989 1507
rect 994 1503 997 1507
rect 997 1503 999 1507
rect 984 1502 989 1503
rect 994 1502 999 1503
rect 2016 1503 2018 1507
rect 2018 1503 2021 1507
rect 2026 1503 2029 1507
rect 2029 1503 2031 1507
rect 2016 1502 2021 1503
rect 2026 1502 2031 1503
rect 480 1403 482 1407
rect 482 1403 485 1407
rect 490 1403 493 1407
rect 493 1403 495 1407
rect 480 1402 485 1403
rect 490 1402 495 1403
rect 1496 1403 1498 1407
rect 1498 1403 1501 1407
rect 1506 1403 1509 1407
rect 1509 1403 1511 1407
rect 1496 1402 1501 1403
rect 1506 1402 1511 1403
rect 984 1303 986 1307
rect 986 1303 989 1307
rect 994 1303 997 1307
rect 997 1303 999 1307
rect 984 1302 989 1303
rect 994 1302 999 1303
rect 2016 1303 2018 1307
rect 2018 1303 2021 1307
rect 2026 1303 2029 1307
rect 2029 1303 2031 1307
rect 2016 1302 2021 1303
rect 2026 1302 2031 1303
rect 2365 1267 2370 1272
rect 2477 1237 2482 1242
rect 480 1203 482 1207
rect 482 1203 485 1207
rect 490 1203 493 1207
rect 493 1203 495 1207
rect 480 1202 485 1203
rect 490 1202 495 1203
rect 1496 1203 1498 1207
rect 1498 1203 1501 1207
rect 1506 1203 1509 1207
rect 1509 1203 1511 1207
rect 1496 1202 1501 1203
rect 1506 1202 1511 1203
rect 984 1103 986 1107
rect 986 1103 989 1107
rect 994 1103 997 1107
rect 997 1103 999 1107
rect 984 1102 989 1103
rect 994 1102 999 1103
rect 2016 1103 2018 1107
rect 2018 1103 2021 1107
rect 2026 1103 2029 1107
rect 2029 1103 2031 1107
rect 2016 1102 2021 1103
rect 2026 1102 2031 1103
rect 480 1003 482 1007
rect 482 1003 485 1007
rect 490 1003 493 1007
rect 493 1003 495 1007
rect 480 1002 485 1003
rect 490 1002 495 1003
rect 1496 1003 1498 1007
rect 1498 1003 1501 1007
rect 1506 1003 1509 1007
rect 1509 1003 1511 1007
rect 1496 1002 1501 1003
rect 1506 1002 1511 1003
rect 984 903 986 907
rect 986 903 989 907
rect 994 903 997 907
rect 997 903 999 907
rect 984 902 989 903
rect 994 902 999 903
rect 2016 903 2018 907
rect 2018 903 2021 907
rect 2026 903 2029 907
rect 2029 903 2031 907
rect 2016 902 2021 903
rect 2026 902 2031 903
rect 480 803 482 807
rect 482 803 485 807
rect 490 803 493 807
rect 493 803 495 807
rect 480 802 485 803
rect 490 802 495 803
rect 1496 803 1498 807
rect 1498 803 1501 807
rect 1506 803 1509 807
rect 1509 803 1511 807
rect 1496 802 1501 803
rect 1506 802 1511 803
rect 984 703 986 707
rect 986 703 989 707
rect 994 703 997 707
rect 997 703 999 707
rect 984 702 989 703
rect 994 702 999 703
rect 2016 703 2018 707
rect 2018 703 2021 707
rect 2026 703 2029 707
rect 2029 703 2031 707
rect 2016 702 2021 703
rect 2026 702 2031 703
rect 480 603 482 607
rect 482 603 485 607
rect 490 603 493 607
rect 493 603 495 607
rect 480 602 485 603
rect 490 602 495 603
rect 1496 603 1498 607
rect 1498 603 1501 607
rect 1506 603 1509 607
rect 1509 603 1511 607
rect 1496 602 1501 603
rect 1506 602 1511 603
rect 984 503 986 507
rect 986 503 989 507
rect 994 503 997 507
rect 997 503 999 507
rect 984 502 989 503
rect 994 502 999 503
rect 2016 503 2018 507
rect 2018 503 2021 507
rect 2026 503 2029 507
rect 2029 503 2031 507
rect 2016 502 2021 503
rect 2026 502 2031 503
rect 480 403 482 407
rect 482 403 485 407
rect 490 403 493 407
rect 493 403 495 407
rect 480 402 485 403
rect 490 402 495 403
rect 1496 403 1498 407
rect 1498 403 1501 407
rect 1506 403 1509 407
rect 1509 403 1511 407
rect 1496 402 1501 403
rect 1506 402 1511 403
rect 984 303 986 307
rect 986 303 989 307
rect 994 303 997 307
rect 997 303 999 307
rect 984 302 989 303
rect 994 302 999 303
rect 2016 303 2018 307
rect 2018 303 2021 307
rect 2026 303 2029 307
rect 2029 303 2031 307
rect 2016 302 2021 303
rect 2026 302 2031 303
rect 480 203 482 207
rect 482 203 485 207
rect 490 203 493 207
rect 493 203 495 207
rect 480 202 485 203
rect 490 202 495 203
rect 1496 203 1498 207
rect 1498 203 1501 207
rect 1506 203 1509 207
rect 1509 203 1511 207
rect 1496 202 1501 203
rect 1506 202 1511 203
rect 984 103 986 107
rect 986 103 989 107
rect 994 103 997 107
rect 997 103 999 107
rect 984 102 989 103
rect 994 102 999 103
rect 2016 103 2018 107
rect 2018 103 2021 107
rect 2026 103 2029 107
rect 2029 103 2031 107
rect 2016 102 2021 103
rect 2026 102 2031 103
rect 480 3 482 7
rect 482 3 485 7
rect 490 3 493 7
rect 493 3 495 7
rect 480 2 485 3
rect 490 2 495 3
rect 1496 3 1498 7
rect 1498 3 1501 7
rect 1506 3 1509 7
rect 1509 3 1511 7
rect 1496 2 1501 3
rect 1506 2 1511 3
<< metal6 >>
rect 480 2407 496 2430
rect 485 2402 490 2407
rect 495 2402 496 2407
rect 480 2207 496 2402
rect 485 2202 490 2207
rect 495 2202 496 2207
rect 480 2007 496 2202
rect 485 2002 490 2007
rect 495 2002 496 2007
rect 480 1807 496 2002
rect 485 1802 490 1807
rect 495 1802 496 1807
rect 480 1607 496 1802
rect 485 1602 490 1607
rect 495 1602 496 1607
rect 480 1407 496 1602
rect 485 1402 490 1407
rect 495 1402 496 1407
rect 480 1207 496 1402
rect 485 1202 490 1207
rect 495 1202 496 1207
rect 480 1007 496 1202
rect 485 1002 490 1007
rect 495 1002 496 1007
rect 480 807 496 1002
rect 485 802 490 807
rect 495 802 496 807
rect 480 607 496 802
rect 485 602 490 607
rect 495 602 496 607
rect 480 407 496 602
rect 485 402 490 407
rect 495 402 496 407
rect 480 207 496 402
rect 485 202 490 207
rect 495 202 496 207
rect 480 7 496 202
rect 485 2 490 7
rect 495 2 496 7
rect 480 -30 496 2
rect 984 2307 1000 2430
rect 989 2302 994 2307
rect 999 2302 1000 2307
rect 984 2107 1000 2302
rect 989 2102 994 2107
rect 999 2102 1000 2107
rect 984 1907 1000 2102
rect 989 1902 994 1907
rect 999 1902 1000 1907
rect 984 1707 1000 1902
rect 989 1702 994 1707
rect 999 1702 1000 1707
rect 984 1507 1000 1702
rect 989 1502 994 1507
rect 999 1502 1000 1507
rect 984 1307 1000 1502
rect 989 1302 994 1307
rect 999 1302 1000 1307
rect 984 1107 1000 1302
rect 989 1102 994 1107
rect 999 1102 1000 1107
rect 984 907 1000 1102
rect 989 902 994 907
rect 999 902 1000 907
rect 984 707 1000 902
rect 989 702 994 707
rect 999 702 1000 707
rect 984 507 1000 702
rect 989 502 994 507
rect 999 502 1000 507
rect 984 307 1000 502
rect 989 302 994 307
rect 999 302 1000 307
rect 984 107 1000 302
rect 989 102 994 107
rect 999 102 1000 107
rect 984 -30 1000 102
rect 1496 2407 1512 2430
rect 1501 2402 1506 2407
rect 1511 2402 1512 2407
rect 1496 2207 1512 2402
rect 1501 2202 1506 2207
rect 1511 2202 1512 2207
rect 1496 2007 1512 2202
rect 1501 2002 1506 2007
rect 1511 2002 1512 2007
rect 1496 1807 1512 2002
rect 1501 1802 1506 1807
rect 1511 1802 1512 1807
rect 1496 1607 1512 1802
rect 1501 1602 1506 1607
rect 1511 1602 1512 1607
rect 1496 1407 1512 1602
rect 1501 1402 1506 1407
rect 1511 1402 1512 1407
rect 1496 1207 1512 1402
rect 1501 1202 1506 1207
rect 1511 1202 1512 1207
rect 1496 1007 1512 1202
rect 1501 1002 1506 1007
rect 1511 1002 1512 1007
rect 1496 807 1512 1002
rect 1501 802 1506 807
rect 1511 802 1512 807
rect 1496 607 1512 802
rect 1501 602 1506 607
rect 1511 602 1512 607
rect 1496 407 1512 602
rect 1501 402 1506 407
rect 1511 402 1512 407
rect 1496 207 1512 402
rect 1501 202 1506 207
rect 1511 202 1512 207
rect 1496 7 1512 202
rect 1501 2 1506 7
rect 1511 2 1512 7
rect 1496 -30 1512 2
rect 2016 2307 2032 2430
rect 2021 2302 2026 2307
rect 2031 2302 2032 2307
rect 2016 2107 2032 2302
rect 2021 2102 2026 2107
rect 2031 2102 2032 2107
rect 2016 1907 2032 2102
rect 2021 1902 2026 1907
rect 2031 1902 2032 1907
rect 2016 1707 2032 1902
rect 2021 1702 2026 1707
rect 2031 1702 2032 1707
rect 2016 1507 2032 1702
rect 2021 1502 2026 1507
rect 2031 1502 2032 1507
rect 2016 1307 2032 1502
rect 2021 1302 2026 1307
rect 2031 1302 2032 1307
rect 2016 1107 2032 1302
rect 2365 1272 2370 2337
rect 2477 1242 2482 2247
rect 2021 1102 2026 1107
rect 2031 1102 2032 1107
rect 2016 907 2032 1102
rect 2021 902 2026 907
rect 2031 902 2032 907
rect 2016 707 2032 902
rect 2021 702 2026 707
rect 2031 702 2032 707
rect 2016 507 2032 702
rect 2021 502 2026 507
rect 2031 502 2032 507
rect 2016 307 2032 502
rect 2021 302 2026 307
rect 2031 302 2032 307
rect 2016 107 2032 302
rect 2021 102 2026 107
rect 2031 102 2032 107
rect 2016 -30 2032 102
use CLKBUF1  CLKBUF1_37
timestamp 1732942936
transform 1 0 4 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_8
timestamp 1732942936
transform 1 0 76 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1732942936
transform -1 0 100 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_31
timestamp 1732942936
transform 1 0 100 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_189
timestamp 1732942936
transform 1 0 148 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1732942936
transform 1 0 180 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_27
timestamp 1732942936
transform -1 0 156 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_231
timestamp 1732942936
transform -1 0 180 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_5
timestamp 1732942936
transform 1 0 180 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1732942936
transform -1 0 300 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_7
timestamp 1732942936
transform -1 0 332 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1732942936
transform -1 0 236 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1732942936
transform 1 0 236 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1732942936
transform 1 0 332 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_14
timestamp 1732942936
transform 1 0 332 0 1 105
box -2 -3 74 103
use INVX8  INVX8_5
timestamp 1732942936
transform -1 0 444 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_29
timestamp 1732942936
transform 1 0 428 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_33
timestamp 1732942936
transform -1 0 484 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1732942936
transform -1 0 492 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1732942936
transform -1 0 500 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1732942936
transform -1 0 596 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_151
timestamp 1732942936
transform -1 0 492 0 1 105
box -2 -3 50 103
use FILL  FILL_1_0_0
timestamp 1732942936
transform 1 0 492 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1732942936
transform 1 0 500 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_7
timestamp 1732942936
transform 1 0 508 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1732942936
transform -1 0 692 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_6
timestamp 1732942936
transform 1 0 532 0 1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_49
timestamp 1732942936
transform 1 0 604 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_5
timestamp 1732942936
transform 1 0 692 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1732942936
transform -1 0 660 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_110
timestamp 1732942936
transform -1 0 708 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1732942936
transform 1 0 708 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1732942936
transform 1 0 724 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_123
timestamp 1732942936
transform 1 0 804 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_166
timestamp 1732942936
transform 1 0 820 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_147
timestamp 1732942936
transform -1 0 876 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1732942936
transform 1 0 876 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1732942936
transform -1 0 1004 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_109
timestamp 1732942936
transform -1 0 860 0 1 105
box -2 -3 34 103
use INVX8  INVX8_7
timestamp 1732942936
transform -1 0 900 0 1 105
box -2 -3 42 103
use CLKBUF1  CLKBUF1_35
timestamp 1732942936
transform 1 0 900 0 1 105
box -2 -3 74 103
use FILL  FILL_0_1_0
timestamp 1732942936
transform 1 0 1004 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1732942936
transform 1 0 1012 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_1_0
timestamp 1732942936
transform -1 0 980 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1732942936
transform -1 0 988 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_166
timestamp 1732942936
transform -1 0 1036 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_148
timestamp 1732942936
transform 1 0 1020 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_131
timestamp 1732942936
transform -1 0 1076 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_13
timestamp 1732942936
transform 1 0 1076 0 -1 105
box -2 -3 74 103
use MUX2X1  MUX2X1_118
timestamp 1732942936
transform -1 0 1084 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_114
timestamp 1732942936
transform 1 0 1084 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_101
timestamp 1732942936
transform -1 0 1140 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1732942936
transform 1 0 1148 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1732942936
transform -1 0 1236 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_121
timestamp 1732942936
transform 1 0 1244 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_107
timestamp 1732942936
transform -1 0 1300 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1732942936
transform 1 0 1300 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_168
timestamp 1732942936
transform 1 0 1236 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1732942936
transform -1 0 1380 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_133
timestamp 1732942936
transform -1 0 1428 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1732942936
transform 1 0 1380 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_99
timestamp 1732942936
transform -1 0 1436 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1732942936
transform 1 0 1428 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1732942936
transform -1 0 1468 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1732942936
transform -1 0 1476 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1732942936
transform -1 0 1572 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_150
timestamp 1732942936
transform -1 0 1460 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_177
timestamp 1732942936
transform -1 0 1484 0 1 105
box -2 -3 26 103
use FILL  FILL_1_2_0
timestamp 1732942936
transform -1 0 1492 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1732942936
transform -1 0 1500 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_167
timestamp 1732942936
transform -1 0 1548 0 1 105
box -2 -3 50 103
use CLKBUF1  CLKBUF1_7
timestamp 1732942936
transform -1 0 1644 0 -1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_141
timestamp 1732942936
transform 1 0 1548 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_125
timestamp 1732942936
transform -1 0 1604 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1732942936
transform 1 0 1604 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_117
timestamp 1732942936
transform 1 0 1644 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_132
timestamp 1732942936
transform 1 0 1676 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1732942936
transform -1 0 1796 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_230
timestamp 1732942936
transform -1 0 1724 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_149
timestamp 1732942936
transform -1 0 1820 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_132
timestamp 1732942936
transform -1 0 1852 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_188
timestamp 1732942936
transform -1 0 1756 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1732942936
transform -1 0 1852 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1732942936
transform 1 0 1852 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_156
timestamp 1732942936
transform 1 0 1852 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_176
timestamp 1732942936
transform -1 0 1908 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1732942936
transform 1 0 1908 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_148
timestamp 1732942936
transform 1 0 1948 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1732942936
transform -1 0 2004 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_3_0
timestamp 1732942936
transform 1 0 2004 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1732942936
transform 1 0 2012 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1732942936
transform 1 0 2020 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_3_0
timestamp 1732942936
transform -1 0 2012 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1732942936
transform -1 0 2020 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_134
timestamp 1732942936
transform -1 0 2068 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1732942936
transform 1 0 2116 0 -1 105
box -2 -3 98 103
use BUFX4  BUFX4_27
timestamp 1732942936
transform -1 0 2100 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_143
timestamp 1732942936
transform 1 0 2100 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_116
timestamp 1732942936
transform 1 0 2212 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1732942936
transform 1 0 2148 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1732942936
transform -1 0 2204 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_124
timestamp 1732942936
transform 1 0 2204 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1732942936
transform -1 0 2268 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1732942936
transform -1 0 2364 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_140
timestamp 1732942936
transform -1 0 2260 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1732942936
transform -1 0 2356 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_36
timestamp 1732942936
transform 1 0 2364 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_11
timestamp 1732942936
transform -1 0 2428 0 1 105
box -2 -3 74 103
use INVX8  INVX8_6
timestamp 1732942936
transform -1 0 2476 0 -1 105
box -2 -3 42 103
use INVX8  INVX8_4
timestamp 1732942936
transform -1 0 2516 0 -1 105
box -2 -3 42 103
use FILL  FILL_1_1
timestamp 1732942936
transform -1 0 2524 0 -1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_45
timestamp 1732942936
transform -1 0 2500 0 1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_25
timestamp 1732942936
transform -1 0 2524 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_229
timestamp 1732942936
transform 1 0 4 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_187
timestamp 1732942936
transform -1 0 60 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1732942936
transform 1 0 60 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_173
timestamp 1732942936
transform -1 0 116 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1732942936
transform 1 0 116 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1732942936
transform 1 0 212 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1732942936
transform -1 0 404 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1732942936
transform -1 0 500 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1732942936
transform 1 0 500 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1732942936
transform 1 0 508 0 -1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_100
timestamp 1732942936
transform 1 0 516 0 -1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_155
timestamp 1732942936
transform 1 0 564 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1732942936
transform -1 0 620 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1732942936
transform 1 0 620 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_109
timestamp 1732942936
transform -1 0 764 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_157
timestamp 1732942936
transform 1 0 764 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_139
timestamp 1732942936
transform -1 0 820 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1732942936
transform 1 0 820 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1732942936
transform -1 0 948 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_1_0
timestamp 1732942936
transform -1 0 956 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1732942936
transform -1 0 964 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1732942936
transform -1 0 1060 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_58
timestamp 1732942936
transform 1 0 1060 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_51
timestamp 1732942936
transform -1 0 1116 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1732942936
transform 1 0 1116 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_168
timestamp 1732942936
transform -1 0 1172 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1732942936
transform 1 0 1172 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_123
timestamp 1732942936
transform 1 0 1268 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1732942936
transform -1 0 1324 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1732942936
transform 1 0 1324 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_115
timestamp 1732942936
transform -1 0 1452 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_158
timestamp 1732942936
transform 1 0 1452 0 -1 305
box -2 -3 50 103
use FILL  FILL_2_2_0
timestamp 1732942936
transform 1 0 1500 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1732942936
transform 1 0 1508 0 -1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_157
timestamp 1732942936
transform 1 0 1516 0 -1 305
box -2 -3 50 103
use BUFX4  BUFX4_44
timestamp 1732942936
transform 1 0 1564 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1732942936
transform 1 0 1596 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_141
timestamp 1732942936
transform -1 0 1652 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1732942936
transform 1 0 1652 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1732942936
transform -1 0 1716 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1732942936
transform -1 0 1812 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_113
timestamp 1732942936
transform 1 0 1812 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_100
timestamp 1732942936
transform -1 0 1868 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1732942936
transform -1 0 1964 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_133
timestamp 1732942936
transform 1 0 1964 0 -1 305
box -2 -3 50 103
use FILL  FILL_2_3_0
timestamp 1732942936
transform 1 0 2012 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1732942936
transform 1 0 2020 0 -1 305
box -2 -3 10 103
use BUFX4  BUFX4_36
timestamp 1732942936
transform 1 0 2028 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_158
timestamp 1732942936
transform 1 0 2060 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_140
timestamp 1732942936
transform -1 0 2116 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1732942936
transform 1 0 2116 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_28
timestamp 1732942936
transform -1 0 2180 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1732942936
transform -1 0 2276 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_151
timestamp 1732942936
transform 1 0 2276 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1732942936
transform -1 0 2396 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1732942936
transform -1 0 2492 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_166
timestamp 1732942936
transform 1 0 2492 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1732942936
transform 1 0 4 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_103
timestamp 1732942936
transform -1 0 148 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_91
timestamp 1732942936
transform 1 0 148 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1732942936
transform -1 0 204 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1732942936
transform 1 0 204 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_146
timestamp 1732942936
transform 1 0 300 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_98
timestamp 1732942936
transform -1 0 396 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_193
timestamp 1732942936
transform 1 0 396 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_171
timestamp 1732942936
transform -1 0 452 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1732942936
transform -1 0 484 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1732942936
transform 1 0 484 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1732942936
transform 1 0 492 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_3
timestamp 1732942936
transform 1 0 500 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_3
timestamp 1732942936
transform -1 0 556 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_102
timestamp 1732942936
transform 1 0 556 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_101
timestamp 1732942936
transform -1 0 652 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_111
timestamp 1732942936
transform -1 0 700 0 1 305
box -2 -3 50 103
use BUFX4  BUFX4_41
timestamp 1732942936
transform -1 0 732 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1732942936
transform 1 0 732 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_40
timestamp 1732942936
transform 1 0 828 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_15
timestamp 1732942936
transform 1 0 852 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_17
timestamp 1732942936
transform 1 0 884 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_160
timestamp 1732942936
transform -1 0 956 0 1 305
box -2 -3 50 103
use BUFX4  BUFX4_43
timestamp 1732942936
transform -1 0 988 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1732942936
transform -1 0 996 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1732942936
transform -1 0 1004 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_120
timestamp 1732942936
transform -1 0 1052 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_5
timestamp 1732942936
transform 1 0 1052 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_5
timestamp 1732942936
transform -1 0 1108 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1732942936
transform 1 0 1108 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_148
timestamp 1732942936
transform 1 0 1204 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_119
timestamp 1732942936
transform -1 0 1300 0 1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1732942936
transform -1 0 1396 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_130
timestamp 1732942936
transform 1 0 1396 0 1 305
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1732942936
transform 1 0 1420 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_159
timestamp 1732942936
transform -1 0 1492 0 1 305
box -2 -3 50 103
use FILL  FILL_3_2_0
timestamp 1732942936
transform -1 0 1500 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1732942936
transform -1 0 1508 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1732942936
transform -1 0 1604 0 1 305
box -2 -3 98 103
use BUFX4  BUFX4_34
timestamp 1732942936
transform -1 0 1636 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1732942936
transform 1 0 1636 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1732942936
transform -1 0 1692 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_127
timestamp 1732942936
transform 1 0 1692 0 1 305
box -2 -3 50 103
use BUFX4  BUFX4_29
timestamp 1732942936
transform 1 0 1740 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_142
timestamp 1732942936
transform 1 0 1772 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_122
timestamp 1732942936
transform 1 0 1820 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_108
timestamp 1732942936
transform -1 0 1876 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1732942936
transform -1 0 1972 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_135
timestamp 1732942936
transform 1 0 1972 0 1 305
box -2 -3 50 103
use FILL  FILL_3_3_0
timestamp 1732942936
transform -1 0 2028 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1732942936
transform -1 0 2036 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1732942936
transform -1 0 2132 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_59
timestamp 1732942936
transform -1 0 2156 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_125
timestamp 1732942936
transform 1 0 2156 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_92
timestamp 1732942936
transform 1 0 2204 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1732942936
transform -1 0 2260 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_121
timestamp 1732942936
transform -1 0 2308 0 1 305
box -2 -3 50 103
use NOR2X1  NOR2X1_8
timestamp 1732942936
transform 1 0 2308 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1732942936
transform -1 0 2364 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1732942936
transform 1 0 2364 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1732942936
transform -1 0 2420 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1732942936
transform 1 0 2420 0 1 305
box -2 -3 98 103
use FILL  FILL_4_1
timestamp 1732942936
transform 1 0 2516 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_5
timestamp 1732942936
transform -1 0 28 0 -1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_16
timestamp 1732942936
transform -1 0 100 0 -1 505
box -2 -3 74 103
use NAND2X1  NAND2X1_24
timestamp 1732942936
transform 1 0 100 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1732942936
transform -1 0 156 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1732942936
transform 1 0 156 0 -1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_97
timestamp 1732942936
transform -1 0 300 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_22
timestamp 1732942936
transform 1 0 300 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_19
timestamp 1732942936
transform -1 0 356 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1732942936
transform -1 0 452 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_209
timestamp 1732942936
transform -1 0 476 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1732942936
transform 1 0 476 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1732942936
transform 1 0 484 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_215
timestamp 1732942936
transform 1 0 492 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1732942936
transform -1 0 612 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1732942936
transform 1 0 612 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_37
timestamp 1732942936
transform 1 0 708 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1732942936
transform -1 0 764 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1732942936
transform 1 0 764 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_15
timestamp 1732942936
transform 1 0 860 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_13
timestamp 1732942936
transform -1 0 916 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1732942936
transform -1 0 1012 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_1_0
timestamp 1732942936
transform 1 0 1012 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1732942936
transform 1 0 1020 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_186
timestamp 1732942936
transform 1 0 1028 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_165
timestamp 1732942936
transform -1 0 1084 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1732942936
transform -1 0 1116 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_5
timestamp 1732942936
transform -1 0 1188 0 -1 505
box -2 -3 74 103
use OAI21X1  OAI21X1_45
timestamp 1732942936
transform 1 0 1188 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1732942936
transform -1 0 1244 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1732942936
transform -1 0 1340 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_42
timestamp 1732942936
transform 1 0 1340 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_222
timestamp 1732942936
transform 1 0 1372 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1732942936
transform 1 0 1396 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_2_0
timestamp 1732942936
transform -1 0 1500 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1732942936
transform -1 0 1508 0 -1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_164
timestamp 1732942936
transform -1 0 1556 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_96
timestamp 1732942936
transform 1 0 1556 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_85
timestamp 1732942936
transform -1 0 1612 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1732942936
transform -1 0 1644 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1732942936
transform -1 0 1676 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1732942936
transform -1 0 1708 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1732942936
transform 1 0 1708 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_37
timestamp 1732942936
transform 1 0 1740 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1732942936
transform -1 0 1804 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_12
timestamp 1732942936
transform 1 0 1804 0 -1 505
box -2 -3 74 103
use MUX2X1  MUX2X1_144
timestamp 1732942936
transform 1 0 1876 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1732942936
transform -1 0 2020 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_3_0
timestamp 1732942936
transform -1 0 2028 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1732942936
transform -1 0 2036 0 -1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_136
timestamp 1732942936
transform -1 0 2084 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1732942936
transform -1 0 2180 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_185
timestamp 1732942936
transform 1 0 2180 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_164
timestamp 1732942936
transform -1 0 2236 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_16
timestamp 1732942936
transform 1 0 2236 0 -1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_123
timestamp 1732942936
transform 1 0 2260 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_122
timestamp 1732942936
transform -1 0 2356 0 -1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_172
timestamp 1732942936
transform 1 0 2356 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_194
timestamp 1732942936
transform -1 0 2412 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1732942936
transform 1 0 2412 0 -1 505
box -2 -3 98 103
use FILL  FILL_5_1
timestamp 1732942936
transform -1 0 2516 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1732942936
transform -1 0 2524 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_67
timestamp 1732942936
transform 1 0 4 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_59
timestamp 1732942936
transform -1 0 60 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1732942936
transform 1 0 60 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1732942936
transform 1 0 156 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_105
timestamp 1732942936
transform 1 0 252 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_93
timestamp 1732942936
transform -1 0 308 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1732942936
transform -1 0 404 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_145
timestamp 1732942936
transform -1 0 452 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_99
timestamp 1732942936
transform 1 0 452 0 1 505
box -2 -3 50 103
use FILL  FILL_5_0_0
timestamp 1732942936
transform 1 0 500 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1732942936
transform 1 0 508 0 1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_105
timestamp 1732942936
transform 1 0 516 0 1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_29
timestamp 1732942936
transform 1 0 564 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1732942936
transform -1 0 628 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1732942936
transform 1 0 628 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1732942936
transform -1 0 684 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1732942936
transform 1 0 684 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_149
timestamp 1732942936
transform -1 0 828 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_150
timestamp 1732942936
transform -1 0 876 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_153
timestamp 1732942936
transform 1 0 876 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_152
timestamp 1732942936
transform 1 0 924 0 1 505
box -2 -3 50 103
use FILL  FILL_5_1_0
timestamp 1732942936
transform -1 0 980 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1732942936
transform -1 0 988 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1732942936
transform -1 0 1084 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_60
timestamp 1732942936
transform 1 0 1084 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_53
timestamp 1732942936
transform -1 0 1140 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1732942936
transform 1 0 1140 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_223
timestamp 1732942936
transform -1 0 1188 0 1 505
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1732942936
transform -1 0 1204 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_162
timestamp 1732942936
transform 1 0 1204 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_69
timestamp 1732942936
transform -1 0 1276 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_61
timestamp 1732942936
transform -1 0 1308 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1732942936
transform 1 0 1308 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_23
timestamp 1732942936
transform 1 0 1404 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1732942936
transform -1 0 1460 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_161
timestamp 1732942936
transform -1 0 1508 0 1 505
box -2 -3 50 103
use FILL  FILL_5_2_0
timestamp 1732942936
transform 1 0 1508 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1732942936
transform 1 0 1516 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_221
timestamp 1732942936
transform 1 0 1524 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_270
timestamp 1732942936
transform -1 0 1580 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1732942936
transform 1 0 1580 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1732942936
transform -1 0 1772 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1732942936
transform 1 0 1772 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_36
timestamp 1732942936
transform -1 0 1900 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1732942936
transform -1 0 1924 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_89
timestamp 1732942936
transform -1 0 1972 0 1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_24
timestamp 1732942936
transform 1 0 1972 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_20
timestamp 1732942936
transform -1 0 2028 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1732942936
transform 1 0 2028 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1732942936
transform 1 0 2036 0 1 505
box -2 -3 10 103
use BUFX4  BUFX4_32
timestamp 1732942936
transform 1 0 2044 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_9
timestamp 1732942936
transform 1 0 2076 0 1 505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1732942936
transform -1 0 2244 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_14
timestamp 1732942936
transform -1 0 2276 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1732942936
transform -1 0 2372 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_220
timestamp 1732942936
transform -1 0 2404 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1732942936
transform -1 0 2500 0 1 505
box -2 -3 98 103
use FILL  FILL_6_1
timestamp 1732942936
transform 1 0 2500 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1732942936
transform 1 0 2508 0 1 505
box -2 -3 10 103
use FILL  FILL_6_3
timestamp 1732942936
transform 1 0 2516 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_248
timestamp 1732942936
transform 1 0 4 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_203
timestamp 1732942936
transform -1 0 60 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_107
timestamp 1732942936
transform -1 0 108 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1732942936
transform 1 0 108 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1732942936
transform 1 0 204 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_113
timestamp 1732942936
transform 1 0 300 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_108
timestamp 1732942936
transform 1 0 348 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_147
timestamp 1732942936
transform -1 0 444 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_114
timestamp 1732942936
transform -1 0 492 0 -1 705
box -2 -3 50 103
use FILL  FILL_6_0_0
timestamp 1732942936
transform -1 0 500 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1732942936
transform -1 0 508 0 -1 705
box -2 -3 10 103
use AOI22X1  AOI22X1_18
timestamp 1732942936
transform -1 0 548 0 -1 705
box -2 -3 42 103
use AOI22X1  AOI22X1_17
timestamp 1732942936
transform 1 0 548 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_210
timestamp 1732942936
transform 1 0 588 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_179
timestamp 1732942936
transform 1 0 612 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1732942936
transform -1 0 684 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_211
timestamp 1732942936
transform 1 0 684 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_104
timestamp 1732942936
transform -1 0 756 0 -1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_25
timestamp 1732942936
transform 1 0 756 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_181
timestamp 1732942936
transform -1 0 828 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_216
timestamp 1732942936
transform 1 0 828 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1732942936
transform 1 0 852 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_26
timestamp 1732942936
transform 1 0 884 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_224
timestamp 1732942936
transform 1 0 924 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_1_0
timestamp 1732942936
transform -1 0 956 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1732942936
transform -1 0 964 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1732942936
transform -1 0 1060 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_3
timestamp 1732942936
transform 1 0 1060 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_7
timestamp 1732942936
transform 1 0 1076 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_252
timestamp 1732942936
transform 1 0 1100 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_217
timestamp 1732942936
transform -1 0 1148 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_27
timestamp 1732942936
transform -1 0 1188 0 -1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1732942936
transform -1 0 1284 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_250
timestamp 1732942936
transform 1 0 1284 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_205
timestamp 1732942936
transform -1 0 1340 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1732942936
transform 1 0 1340 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_41
timestamp 1732942936
transform -1 0 1396 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1732942936
transform 1 0 1396 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_2_0
timestamp 1732942936
transform 1 0 1492 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1732942936
transform 1 0 1500 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1732942936
transform 1 0 1508 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_259
timestamp 1732942936
transform 1 0 1604 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_212
timestamp 1732942936
transform -1 0 1660 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_22
timestamp 1732942936
transform -1 0 1700 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_129
timestamp 1732942936
transform 1 0 1700 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1732942936
transform 1 0 1748 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_213
timestamp 1732942936
transform -1 0 1868 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_138
timestamp 1732942936
transform -1 0 1916 0 -1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_23
timestamp 1732942936
transform -1 0 1956 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_90
timestamp 1732942936
transform -1 0 2004 0 -1 705
box -2 -3 50 103
use FILL  FILL_6_3_0
timestamp 1732942936
transform -1 0 2012 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1732942936
transform -1 0 2020 0 -1 705
box -2 -3 10 103
use AOI22X1  AOI22X1_21
timestamp 1732942936
transform -1 0 2060 0 -1 705
box -2 -3 42 103
use BUFX4  BUFX4_26
timestamp 1732942936
transform -1 0 2092 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_25
timestamp 1732942936
transform 1 0 2092 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_58
timestamp 1732942936
transform 1 0 2124 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1732942936
transform -1 0 2252 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_88
timestamp 1732942936
transform -1 0 2300 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_269
timestamp 1732942936
transform 1 0 2300 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1732942936
transform -1 0 2420 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1732942936
transform 1 0 2420 0 -1 705
box -2 -3 98 103
use FILL  FILL_7_1
timestamp 1732942936
transform -1 0 2524 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1732942936
transform 1 0 4 0 1 705
box -2 -3 98 103
use BUFX2  BUFX2_6
timestamp 1732942936
transform -1 0 124 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1732942936
transform 1 0 124 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1732942936
transform -1 0 180 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_211
timestamp 1732942936
transform 1 0 180 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_258
timestamp 1732942936
transform -1 0 236 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1732942936
transform 1 0 236 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_25
timestamp 1732942936
transform -1 0 292 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_163
timestamp 1732942936
transform 1 0 292 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_184
timestamp 1732942936
transform -1 0 348 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1732942936
transform 1 0 348 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_112
timestamp 1732942936
transform 1 0 444 0 1 705
box -2 -3 50 103
use FILL  FILL_7_0_0
timestamp 1732942936
transform 1 0 492 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1732942936
transform 1 0 500 0 1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_15
timestamp 1732942936
transform 1 0 508 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1732942936
transform -1 0 564 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1732942936
transform -1 0 660 0 1 705
box -2 -3 98 103
use BUFX4  BUFX4_1
timestamp 1732942936
transform -1 0 692 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1732942936
transform 1 0 692 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1732942936
transform 1 0 724 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_278
timestamp 1732942936
transform -1 0 780 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1732942936
transform 1 0 780 0 1 705
box -2 -3 98 103
use AOI22X1  AOI22X1_20
timestamp 1732942936
transform 1 0 876 0 1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_98
timestamp 1732942936
transform 1 0 916 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_116
timestamp 1732942936
transform -1 0 964 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_280
timestamp 1732942936
transform 1 0 964 0 1 705
box -2 -3 26 103
use FILL  FILL_7_1_0
timestamp 1732942936
transform -1 0 996 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1732942936
transform -1 0 1004 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_229
timestamp 1732942936
transform -1 0 1036 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1732942936
transform 1 0 1036 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1732942936
transform 1 0 1068 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1732942936
transform -1 0 1116 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_33
timestamp 1732942936
transform -1 0 1140 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_156
timestamp 1732942936
transform -1 0 1188 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_242
timestamp 1732942936
transform 1 0 1188 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_32
timestamp 1732942936
transform -1 0 1236 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_155
timestamp 1732942936
transform -1 0 1284 0 1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_28
timestamp 1732942936
transform -1 0 1324 0 1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_165
timestamp 1732942936
transform 1 0 1324 0 1 705
box -2 -3 50 103
use AND2X2  AND2X2_1
timestamp 1732942936
transform 1 0 1372 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_243
timestamp 1732942936
transform 1 0 1404 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_11
timestamp 1732942936
transform 1 0 1428 0 1 705
box -2 -3 34 103
use FILL  FILL_7_2_0
timestamp 1732942936
transform -1 0 1468 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1732942936
transform -1 0 1476 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1732942936
transform -1 0 1572 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_212
timestamp 1732942936
transform -1 0 1596 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1732942936
transform 1 0 1596 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1732942936
transform -1 0 1660 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_196
timestamp 1732942936
transform 1 0 1660 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_239
timestamp 1732942936
transform -1 0 1716 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1732942936
transform 1 0 1716 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_180
timestamp 1732942936
transform -1 0 1844 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_130
timestamp 1732942936
transform 1 0 1844 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_132
timestamp 1732942936
transform 1 0 1892 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_12
timestamp 1732942936
transform 1 0 1940 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1732942936
transform -1 0 1996 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_214
timestamp 1732942936
transform 1 0 1996 0 1 705
box -2 -3 26 103
use FILL  FILL_7_3_0
timestamp 1732942936
transform -1 0 2028 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1732942936
transform -1 0 2036 0 1 705
box -2 -3 10 103
use AOI22X1  AOI22X1_24
timestamp 1732942936
transform -1 0 2076 0 1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_128
timestamp 1732942936
transform 1 0 2076 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_66
timestamp 1732942936
transform 1 0 2124 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_279
timestamp 1732942936
transform 1 0 2148 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_228
timestamp 1732942936
transform 1 0 2172 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_126
timestamp 1732942936
transform -1 0 2252 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1732942936
transform -1 0 2348 0 1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_20
timestamp 1732942936
transform 1 0 2348 0 1 705
box -2 -3 74 103
use NOR2X1  NOR2X1_14
timestamp 1732942936
transform 1 0 2420 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1732942936
transform -1 0 2476 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1732942936
transform -1 0 2508 0 1 705
box -2 -3 34 103
use FILL  FILL_8_1
timestamp 1732942936
transform 1 0 2508 0 1 705
box -2 -3 10 103
use FILL  FILL_8_2
timestamp 1732942936
transform 1 0 2516 0 1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_46
timestamp 1732942936
transform 1 0 4 0 -1 905
box -2 -3 74 103
use NAND2X1  NAND2X1_64
timestamp 1732942936
transform -1 0 100 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1732942936
transform 1 0 100 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1732942936
transform -1 0 292 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_106
timestamp 1732942936
transform -1 0 340 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_94
timestamp 1732942936
transform -1 0 364 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_116
timestamp 1732942936
transform 1 0 364 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_268
timestamp 1732942936
transform 1 0 412 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_0_0
timestamp 1732942936
transform -1 0 444 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1732942936
transform -1 0 452 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1732942936
transform -1 0 548 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_75
timestamp 1732942936
transform 1 0 548 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1732942936
transform -1 0 604 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_117
timestamp 1732942936
transform -1 0 652 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1732942936
transform -1 0 748 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_15
timestamp 1732942936
transform -1 0 820 0 -1 905
box -2 -3 74 103
use NAND2X1  NAND2X1_44
timestamp 1732942936
transform -1 0 844 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_152
timestamp 1732942936
transform -1 0 868 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_233
timestamp 1732942936
transform -1 0 892 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_80
timestamp 1732942936
transform 1 0 892 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_188
timestamp 1732942936
transform -1 0 940 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_125
timestamp 1732942936
transform 1 0 940 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_283
timestamp 1732942936
transform -1 0 988 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1732942936
transform 1 0 988 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1732942936
transform 1 0 996 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_17
timestamp 1732942936
transform 1 0 1004 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1732942936
transform 1 0 1028 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1732942936
transform 1 0 1052 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_213
timestamp 1732942936
transform 1 0 1148 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_260
timestamp 1732942936
transform -1 0 1204 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_154
timestamp 1732942936
transform 1 0 1204 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_197
timestamp 1732942936
transform 1 0 1252 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_240
timestamp 1732942936
transform -1 0 1308 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1732942936
transform -1 0 1404 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1732942936
transform -1 0 1500 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_2_0
timestamp 1732942936
transform 1 0 1500 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1732942936
transform 1 0 1508 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_86
timestamp 1732942936
transform 1 0 1516 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_76
timestamp 1732942936
transform -1 0 1572 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1732942936
transform 1 0 1572 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_137
timestamp 1732942936
transform -1 0 1652 0 -1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_26
timestamp 1732942936
transform 1 0 1652 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1732942936
transform -1 0 1708 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1732942936
transform -1 0 1804 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_139
timestamp 1732942936
transform -1 0 1852 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_141
timestamp 1732942936
transform 1 0 1852 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_131
timestamp 1732942936
transform 1 0 1900 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_249
timestamp 1732942936
transform 1 0 1948 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_68
timestamp 1732942936
transform 1 0 1972 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_60
timestamp 1732942936
transform -1 0 2028 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_3_0
timestamp 1732942936
transform -1 0 2036 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1732942936
transform -1 0 2044 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1732942936
transform -1 0 2140 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_140
timestamp 1732942936
transform -1 0 2188 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_95
timestamp 1732942936
transform 1 0 2188 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_124
timestamp 1732942936
transform 1 0 2212 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_50
timestamp 1732942936
transform 1 0 2260 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1732942936
transform -1 0 2316 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1732942936
transform 1 0 2316 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_18
timestamp 1732942936
transform 1 0 2412 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_4
timestamp 1732942936
transform -1 0 2516 0 -1 905
box -2 -3 74 103
use FILL  FILL_9_1
timestamp 1732942936
transform -1 0 2524 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_56
timestamp 1732942936
transform -1 0 36 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1732942936
transform 1 0 36 0 1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_43
timestamp 1732942936
transform -1 0 180 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_73
timestamp 1732942936
transform 1 0 180 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_64
timestamp 1732942936
transform -1 0 236 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_238
timestamp 1732942936
transform 1 0 236 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_195
timestamp 1732942936
transform -1 0 292 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1732942936
transform 1 0 292 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1732942936
transform 1 0 324 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_219
timestamp 1732942936
transform -1 0 452 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_45
timestamp 1732942936
transform 1 0 452 0 1 905
box -2 -3 50 103
use FILL  FILL_9_0_0
timestamp 1732942936
transform 1 0 500 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1732942936
transform 1 0 508 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1732942936
transform 1 0 516 0 1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_115
timestamp 1732942936
transform 1 0 612 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_76
timestamp 1732942936
transform 1 0 660 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1732942936
transform -1 0 716 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_232
timestamp 1732942936
transform 1 0 716 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1732942936
transform 1 0 748 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1732942936
transform 1 0 844 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_8
timestamp 1732942936
transform -1 0 964 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_87
timestamp 1732942936
transform -1 0 988 0 1 905
box -2 -3 26 103
use FILL  FILL_9_1_0
timestamp 1732942936
transform -1 0 996 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1732942936
transform -1 0 1004 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_77
timestamp 1732942936
transform -1 0 1036 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1732942936
transform 1 0 1036 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_253
timestamp 1732942936
transform 1 0 1132 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_179
timestamp 1732942936
transform 1 0 1156 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_163
timestamp 1732942936
transform -1 0 1228 0 1 905
box -2 -3 50 103
use AND2X2  AND2X2_4
timestamp 1732942936
transform -1 0 1260 0 1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_47
timestamp 1732942936
transform 1 0 1260 0 1 905
box -2 -3 74 103
use NAND2X1  NAND2X1_35
timestamp 1732942936
transform 1 0 1332 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_7
timestamp 1732942936
transform -1 0 1388 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1732942936
transform -1 0 1420 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1732942936
transform -1 0 1452 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1732942936
transform 1 0 1452 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1732942936
transform -1 0 1516 0 1 905
box -2 -3 34 103
use FILL  FILL_9_2_0
timestamp 1732942936
transform -1 0 1524 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1732942936
transform -1 0 1532 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_83
timestamp 1732942936
transform -1 0 1580 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_40
timestamp 1732942936
transform -1 0 1604 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1732942936
transform -1 0 1700 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1732942936
transform 1 0 1700 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1732942936
transform -1 0 1892 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_77
timestamp 1732942936
transform 1 0 1892 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_68
timestamp 1732942936
transform -1 0 1948 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1732942936
transform -1 0 2044 0 1 905
box -2 -3 98 103
use FILL  FILL_9_3_0
timestamp 1732942936
transform -1 0 2052 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1732942936
transform -1 0 2060 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_204
timestamp 1732942936
transform -1 0 2092 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_77
timestamp 1732942936
transform 1 0 2092 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_39
timestamp 1732942936
transform -1 0 2164 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1732942936
transform -1 0 2260 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_84
timestamp 1732942936
transform -1 0 2292 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1732942936
transform 1 0 2292 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1732942936
transform -1 0 2348 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1732942936
transform 1 0 2348 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_21
timestamp 1732942936
transform -1 0 2468 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_73
timestamp 1732942936
transform 1 0 2468 0 1 905
box -2 -3 50 103
use FILL  FILL_10_1
timestamp 1732942936
transform 1 0 2516 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1732942936
transform 1 0 4 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_54
timestamp 1732942936
transform -1 0 132 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1732942936
transform -1 0 228 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_82
timestamp 1732942936
transform 1 0 228 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1732942936
transform -1 0 284 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1732942936
transform -1 0 380 0 -1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_40
timestamp 1732942936
transform -1 0 452 0 -1 1105
box -2 -3 74 103
use NAND2X1  NAND2X1_91
timestamp 1732942936
transform -1 0 476 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_0_0
timestamp 1732942936
transform 1 0 476 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1732942936
transform 1 0 484 0 -1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_44
timestamp 1732942936
transform 1 0 492 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1732942936
transform -1 0 636 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_265
timestamp 1732942936
transform -1 0 660 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_216
timestamp 1732942936
transform -1 0 692 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1732942936
transform 1 0 692 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1732942936
transform -1 0 748 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1732942936
transform -1 0 844 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1732942936
transform 1 0 844 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_32
timestamp 1732942936
transform 1 0 940 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1732942936
transform -1 0 996 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1732942936
transform -1 0 1004 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1732942936
transform -1 0 1012 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_89
timestamp 1732942936
transform -1 0 1036 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_143
timestamp 1732942936
transform -1 0 1060 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_26
timestamp 1732942936
transform 1 0 1060 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_107
timestamp 1732942936
transform -1 0 1108 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_71
timestamp 1732942936
transform 1 0 1108 0 -1 1105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_39
timestamp 1732942936
transform 1 0 1132 0 -1 1105
box -2 -3 74 103
use NAND2X1  NAND2X1_170
timestamp 1732942936
transform 1 0 1204 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_78
timestamp 1732942936
transform 1 0 1228 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1732942936
transform -1 0 1284 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_263
timestamp 1732942936
transform 1 0 1284 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_134
timestamp 1732942936
transform -1 0 1332 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_273
timestamp 1732942936
transform 1 0 1332 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1732942936
transform -1 0 1452 0 -1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_10
timestamp 1732942936
transform 1 0 1452 0 -1 1105
box -2 -3 74 103
use FILL  FILL_10_2_0
timestamp 1732942936
transform 1 0 1524 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1732942936
transform 1 0 1532 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_247
timestamp 1732942936
transform 1 0 1540 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_84
timestamp 1732942936
transform 1 0 1564 0 -1 1105
box -2 -3 50 103
use AOI22X1  AOI22X1_14
timestamp 1732942936
transform -1 0 1652 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_207
timestamp 1732942936
transform -1 0 1676 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_178
timestamp 1732942936
transform 1 0 1676 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1732942936
transform -1 0 1740 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_206
timestamp 1732942936
transform 1 0 1740 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1732942936
transform -1 0 1860 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_50
timestamp 1732942936
transform -1 0 1892 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1732942936
transform -1 0 1988 0 -1 1105
box -2 -3 98 103
use AOI22X1  AOI22X1_13
timestamp 1732942936
transform -1 0 2028 0 -1 1105
box -2 -3 42 103
use FILL  FILL_10_3_0
timestamp 1732942936
transform -1 0 2036 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1732942936
transform -1 0 2044 0 -1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_78
timestamp 1732942936
transform -1 0 2092 0 -1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_34
timestamp 1732942936
transform 1 0 2092 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1732942936
transform 1 0 2124 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_2
timestamp 1732942936
transform -1 0 2244 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_76
timestamp 1732942936
transform 1 0 2244 0 -1 1105
box -2 -3 50 103
use BUFX2  BUFX2_4
timestamp 1732942936
transform 1 0 2292 0 -1 1105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_19
timestamp 1732942936
transform 1 0 2316 0 -1 1105
box -2 -3 74 103
use NAND2X1  NAND2X1_48
timestamp 1732942936
transform 1 0 2388 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_42
timestamp 1732942936
transform -1 0 2444 0 -1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_33
timestamp 1732942936
transform 1 0 2444 0 -1 1105
box -2 -3 74 103
use FILL  FILL_11_1
timestamp 1732942936
transform -1 0 2524 0 -1 1105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_26
timestamp 1732942936
transform -1 0 76 0 1 1105
box -2 -3 74 103
use NAND2X1  NAND2X1_255
timestamp 1732942936
transform 1 0 76 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1732942936
transform -1 0 132 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1732942936
transform 1 0 132 0 1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_34
timestamp 1732942936
transform 1 0 228 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_235
timestamp 1732942936
transform 1 0 276 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_192
timestamp 1732942936
transform 1 0 300 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1732942936
transform 1 0 332 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_80
timestamp 1732942936
transform -1 0 460 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1732942936
transform -1 0 468 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1732942936
transform -1 0 476 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1732942936
transform -1 0 572 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_40
timestamp 1732942936
transform 1 0 572 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1732942936
transform -1 0 628 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_28
timestamp 1732942936
transform -1 0 676 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_30
timestamp 1732942936
transform 1 0 676 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_285
timestamp 1732942936
transform 1 0 724 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_46
timestamp 1732942936
transform -1 0 796 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_136
timestamp 1732942936
transform 1 0 796 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1732942936
transform -1 0 852 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1732942936
transform 1 0 852 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_37
timestamp 1732942936
transform 1 0 948 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_163
timestamp 1732942936
transform 1 0 972 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1732942936
transform -1 0 1004 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1732942936
transform -1 0 1012 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_144
timestamp 1732942936
transform -1 0 1044 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_109
timestamp 1732942936
transform 1 0 1044 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_96
timestamp 1732942936
transform -1 0 1100 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1732942936
transform -1 0 1196 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1732942936
transform -1 0 1292 0 1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_18
timestamp 1732942936
transform 1 0 1292 0 1 1105
box -2 -3 74 103
use MUX2X1  MUX2X1_82
timestamp 1732942936
transform 1 0 1364 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_237
timestamp 1732942936
transform 1 0 1412 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_194
timestamp 1732942936
transform -1 0 1468 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_2_0
timestamp 1732942936
transform -1 0 1476 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1732942936
transform -1 0 1484 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1732942936
transform -1 0 1580 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_202
timestamp 1732942936
transform -1 0 1612 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1732942936
transform 1 0 1612 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_10
timestamp 1732942936
transform 1 0 1708 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1732942936
transform -1 0 1764 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_80
timestamp 1732942936
transform 1 0 1764 0 1 1105
box -2 -3 50 103
use BUFX4  BUFX4_48
timestamp 1732942936
transform -1 0 1844 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1732942936
transform 1 0 1844 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_174
timestamp 1732942936
transform -1 0 1892 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_154
timestamp 1732942936
transform -1 0 1924 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_226
timestamp 1732942936
transform 1 0 1924 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1732942936
transform -1 0 1980 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_3_0
timestamp 1732942936
transform -1 0 1988 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1732942936
transform -1 0 1996 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1732942936
transform -1 0 2092 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1732942936
transform 1 0 2092 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_2
timestamp 1732942936
transform 1 0 2188 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1732942936
transform -1 0 2252 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_75
timestamp 1732942936
transform 1 0 2252 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_74
timestamp 1732942936
transform 1 0 2300 0 1 1105
box -2 -3 50 103
use BUFX4  BUFX4_49
timestamp 1732942936
transform 1 0 2348 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_192
timestamp 1732942936
transform 1 0 2380 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1732942936
transform 1 0 2404 0 1 1105
box -2 -3 98 103
use FILL  FILL_12_1
timestamp 1732942936
transform 1 0 2500 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1732942936
transform 1 0 2508 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_3
timestamp 1732942936
transform 1 0 2516 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1732942936
transform 1 0 4 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_245
timestamp 1732942936
transform -1 0 124 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_200
timestamp 1732942936
transform -1 0 156 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1732942936
transform 1 0 156 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1732942936
transform 1 0 188 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_35
timestamp 1732942936
transform -1 0 332 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_36
timestamp 1732942936
transform 1 0 332 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_26
timestamp 1732942936
transform 1 0 380 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_4
timestamp 1732942936
transform -1 0 452 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1732942936
transform -1 0 484 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1732942936
transform -1 0 492 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1732942936
transform -1 0 500 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1732942936
transform -1 0 596 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_10
timestamp 1732942936
transform 1 0 596 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_8
timestamp 1732942936
transform -1 0 652 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_51
timestamp 1732942936
transform 1 0 652 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_25
timestamp 1732942936
transform 1 0 684 0 -1 1305
box -2 -3 74 103
use MUX2X1  MUX2X1_48
timestamp 1732942936
transform -1 0 804 0 -1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_8
timestamp 1732942936
transform 1 0 804 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_202
timestamp 1732942936
transform -1 0 868 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_53
timestamp 1732942936
transform 1 0 868 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_29
timestamp 1732942936
transform -1 0 948 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_38
timestamp 1732942936
transform 1 0 948 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_1_0
timestamp 1732942936
transform -1 0 1004 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1732942936
transform -1 0 1012 0 -1 1305
box -2 -3 10 103
use AOI22X1  AOI22X1_7
timestamp 1732942936
transform -1 0 1052 0 -1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_39
timestamp 1732942936
transform -1 0 1100 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_37
timestamp 1732942936
transform -1 0 1148 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_48
timestamp 1732942936
transform 1 0 1148 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1732942936
transform -1 0 1204 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1732942936
transform 1 0 1204 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1732942936
transform -1 0 1396 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_257
timestamp 1732942936
transform 1 0 1396 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1732942936
transform -1 0 1452 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_186
timestamp 1732942936
transform 1 0 1452 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_2_0
timestamp 1732942936
transform -1 0 1492 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1732942936
transform -1 0 1500 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1732942936
transform -1 0 1596 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_30
timestamp 1732942936
transform 1 0 1596 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_26
timestamp 1732942936
transform -1 0 1652 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_81
timestamp 1732942936
transform 1 0 1652 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_146
timestamp 1732942936
transform 1 0 1700 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_165
timestamp 1732942936
transform -1 0 1756 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1732942936
transform 1 0 1756 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_86
timestamp 1732942936
transform 1 0 1852 0 -1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_15
timestamp 1732942936
transform -1 0 1940 0 -1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_87
timestamp 1732942936
transform -1 0 1988 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_3_0
timestamp 1732942936
transform -1 0 1996 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1732942936
transform -1 0 2004 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1732942936
transform -1 0 2100 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_129
timestamp 1732942936
transform 1 0 2100 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_114
timestamp 1732942936
transform -1 0 2156 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_85
timestamp 1732942936
transform 1 0 2156 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_156
timestamp 1732942936
transform -1 0 2228 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_138
timestamp 1732942936
transform -1 0 2260 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1732942936
transform -1 0 2356 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_147
timestamp 1732942936
transform 1 0 2356 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1732942936
transform 1 0 2380 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1732942936
transform -1 0 2508 0 -1 1305
box -2 -3 98 103
use FILL  FILL_13_1
timestamp 1732942936
transform -1 0 2516 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1732942936
transform -1 0 2524 0 -1 1305
box -2 -3 10 103
use INVX8  INVX8_2
timestamp 1732942936
transform 1 0 4 0 1 1305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1732942936
transform 1 0 44 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_168
timestamp 1732942936
transform 1 0 140 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1732942936
transform -1 0 196 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_100
timestamp 1732942936
transform -1 0 220 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_25
timestamp 1732942936
transform 1 0 220 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_52
timestamp 1732942936
transform 1 0 268 0 1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_42
timestamp 1732942936
transform 1 0 300 0 1 1305
box -2 -3 74 103
use MUX2X1  MUX2X1_32
timestamp 1732942936
transform -1 0 420 0 1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_6
timestamp 1732942936
transform 1 0 420 0 1 1305
box -2 -3 42 103
use FILL  FILL_13_0_0
timestamp 1732942936
transform 1 0 460 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1732942936
transform 1 0 468 0 1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_27
timestamp 1732942936
transform 1 0 476 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1732942936
transform -1 0 620 0 1 1305
box -2 -3 98 103
use AOI22X1  AOI22X1_5
timestamp 1732942936
transform 1 0 620 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_201
timestamp 1732942936
transform 1 0 660 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_176
timestamp 1732942936
transform 1 0 684 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_50
timestamp 1732942936
transform 1 0 716 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1732942936
transform 1 0 748 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_127
timestamp 1732942936
transform 1 0 796 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_112
timestamp 1732942936
transform -1 0 852 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1732942936
transform 1 0 852 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_172
timestamp 1732942936
transform -1 0 908 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1732942936
transform 1 0 908 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_1_0
timestamp 1732942936
transform 1 0 1004 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1732942936
transform 1 0 1012 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1732942936
transform 1 0 1020 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_136
timestamp 1732942936
transform 1 0 1116 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_120
timestamp 1732942936
transform -1 0 1172 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_42
timestamp 1732942936
transform -1 0 1220 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_145
timestamp 1732942936
transform 1 0 1220 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_128
timestamp 1732942936
transform -1 0 1276 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1732942936
transform -1 0 1372 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1732942936
transform 1 0 1372 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_228
timestamp 1732942936
transform 1 0 1468 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_2_0
timestamp 1732942936
transform -1 0 1500 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1732942936
transform -1 0 1508 0 1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_79
timestamp 1732942936
transform -1 0 1556 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1732942936
transform 1 0 1556 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_94
timestamp 1732942936
transform 1 0 1652 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_120
timestamp 1732942936
transform 1 0 1700 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_106
timestamp 1732942936
transform -1 0 1756 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_96
timestamp 1732942936
transform 1 0 1756 0 1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_16
timestamp 1732942936
transform -1 0 1844 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_208
timestamp 1732942936
transform -1 0 1868 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_45
timestamp 1732942936
transform 1 0 1868 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_95
timestamp 1732942936
transform -1 0 1948 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_66
timestamp 1732942936
transform 1 0 1948 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1732942936
transform -1 0 2004 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_3_0
timestamp 1732942936
transform -1 0 2012 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1732942936
transform -1 0 2020 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1732942936
transform -1 0 2116 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_138
timestamp 1732942936
transform 1 0 2116 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_122
timestamp 1732942936
transform -1 0 2172 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1732942936
transform -1 0 2268 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1732942936
transform -1 0 2364 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_130
timestamp 1732942936
transform -1 0 2396 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1732942936
transform -1 0 2428 0 1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_17
timestamp 1732942936
transform -1 0 2500 0 1 1305
box -2 -3 74 103
use FILL  FILL_14_1
timestamp 1732942936
transform 1 0 2500 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1732942936
transform 1 0 2508 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_3
timestamp 1732942936
transform 1 0 2516 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1732942936
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_19
timestamp 1732942936
transform 1 0 100 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_16
timestamp 1732942936
transform -1 0 156 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1732942936
transform 1 0 156 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_224
timestamp 1732942936
transform 1 0 252 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_275
timestamp 1732942936
transform -1 0 308 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1732942936
transform 1 0 308 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_221
timestamp 1732942936
transform 1 0 324 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_282
timestamp 1732942936
transform -1 0 372 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1732942936
transform -1 0 388 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_33
timestamp 1732942936
transform -1 0 436 0 -1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_272
timestamp 1732942936
transform 1 0 436 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_262
timestamp 1732942936
transform 1 0 460 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_0_0
timestamp 1732942936
transform 1 0 484 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1732942936
transform 1 0 492 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_34
timestamp 1732942936
transform 1 0 500 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_19
timestamp 1732942936
transform -1 0 548 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_20
timestamp 1732942936
transform 1 0 548 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_1
timestamp 1732942936
transform 1 0 572 0 -1 1505
box -2 -3 34 103
use INVX8  INVX8_9
timestamp 1732942936
transform 1 0 604 0 -1 1505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1732942936
transform 1 0 644 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_26
timestamp 1732942936
transform -1 0 772 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_200
timestamp 1732942936
transform -1 0 796 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1732942936
transform -1 0 892 0 -1 1505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_27
timestamp 1732942936
transform 1 0 892 0 -1 1505
box -2 -3 74 103
use FILL  FILL_14_1_0
timestamp 1732942936
transform 1 0 964 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1732942936
transform 1 0 972 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1732942936
transform 1 0 980 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1732942936
transform 1 0 1076 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_41
timestamp 1732942936
transform 1 0 1172 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1732942936
transform 1 0 1220 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_40
timestamp 1732942936
transform -1 0 1364 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1732942936
transform -1 0 1460 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_160
timestamp 1732942936
transform 1 0 1460 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1732942936
transform 1 0 1492 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_2_0
timestamp 1732942936
transform -1 0 1524 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1732942936
transform -1 0 1532 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_198
timestamp 1732942936
transform -1 0 1564 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_98
timestamp 1732942936
transform 1 0 1564 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_111
timestamp 1732942936
transform -1 0 1620 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1732942936
transform 1 0 1620 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_214
timestamp 1732942936
transform -1 0 1748 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1732942936
transform -1 0 1844 0 -1 1505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_38
timestamp 1732942936
transform -1 0 1916 0 -1 1505
box -2 -3 74 103
use MUX2X1  MUX2X1_93
timestamp 1732942936
transform 1 0 1916 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_74
timestamp 1732942936
transform 1 0 1964 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1732942936
transform -1 0 2020 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_3_0
timestamp 1732942936
transform 1 0 2020 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1732942936
transform 1 0 2028 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_91
timestamp 1732942936
transform 1 0 2036 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1732942936
transform -1 0 2180 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_92
timestamp 1732942936
transform -1 0 2228 0 -1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_93
timestamp 1732942936
transform 1 0 2228 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_82
timestamp 1732942936
transform -1 0 2284 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1732942936
transform -1 0 2380 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_218
timestamp 1732942936
transform 1 0 2380 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1732942936
transform 1 0 2412 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1732942936
transform -1 0 2516 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1732942936
transform -1 0 2524 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1732942936
transform 1 0 4 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_226
timestamp 1732942936
transform 1 0 100 0 1 1505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_28
timestamp 1732942936
transform -1 0 76 0 -1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1732942936
transform 1 0 76 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_184
timestamp 1732942936
transform -1 0 156 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_31
timestamp 1732942936
transform -1 0 204 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_191
timestamp 1732942936
transform 1 0 204 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1732942936
transform -1 0 204 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1732942936
transform 1 0 204 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_234
timestamp 1732942936
transform -1 0 260 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1732942936
transform -1 0 356 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_244
timestamp 1732942936
transform 1 0 300 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_29
timestamp 1732942936
transform -1 0 380 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_31
timestamp 1732942936
transform -1 0 404 0 1 1505
box -2 -3 26 103
use INVX2  INVX2_1
timestamp 1732942936
transform -1 0 420 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_199
timestamp 1732942936
transform -1 0 356 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_11
timestamp 1732942936
transform -1 0 404 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_63
timestamp 1732942936
transform 1 0 404 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_10
timestamp 1732942936
transform -1 0 468 0 1 1505
box -2 -3 50 103
use NOR2X1  NOR2X1_43
timestamp 1732942936
transform -1 0 492 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_0_0
timestamp 1732942936
transform -1 0 500 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1732942936
transform -1 0 508 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_2
timestamp 1732942936
transform -1 0 532 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_12
timestamp 1732942936
transform -1 0 476 0 -1 1705
box -2 -3 50 103
use FILL  FILL_16_0_0
timestamp 1732942936
transform -1 0 484 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1732942936
transform -1 0 492 0 -1 1705
box -2 -3 10 103
use AOI22X1  AOI22X1_2
timestamp 1732942936
transform -1 0 532 0 -1 1705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1732942936
transform -1 0 628 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1732942936
transform 1 0 532 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_254
timestamp 1732942936
transform 1 0 628 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_207
timestamp 1732942936
transform -1 0 684 0 1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_31
timestamp 1732942936
transform 1 0 684 0 1 1505
box -2 -3 74 103
use OAI21X1  OAI21X1_151
timestamp 1732942936
transform 1 0 628 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_171
timestamp 1732942936
transform -1 0 684 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_9
timestamp 1732942936
transform 1 0 684 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_143
timestamp 1732942936
transform 1 0 756 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_162
timestamp 1732942936
transform 1 0 788 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_14
timestamp 1732942936
transform -1 0 780 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_135
timestamp 1732942936
transform 1 0 780 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1732942936
transform -1 0 908 0 1 1505
box -2 -3 98 103
use BUFX2  BUFX2_2
timestamp 1732942936
transform 1 0 908 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_153
timestamp 1732942936
transform -1 0 836 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_10
timestamp 1732942936
transform -1 0 876 0 -1 1705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1732942936
transform -1 0 972 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_10
timestamp 1732942936
transform 1 0 932 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_12
timestamp 1732942936
transform -1 0 988 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_1_0
timestamp 1732942936
transform 1 0 988 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1732942936
transform 1 0 996 0 1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_18
timestamp 1732942936
transform 1 0 1004 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_276
timestamp 1732942936
transform 1 0 972 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_1_0
timestamp 1732942936
transform -1 0 1004 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1732942936
transform -1 0 1012 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_225
timestamp 1732942936
transform -1 0 1044 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1732942936
transform -1 0 1060 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1732942936
transform 1 0 1060 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1732942936
transform -1 0 1116 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1732942936
transform 1 0 1044 0 -1 1705
box -2 -3 98 103
use INVX4  INVX4_2
timestamp 1732942936
transform -1 0 1140 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1732942936
transform 1 0 1140 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_153
timestamp 1732942936
transform 1 0 1140 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1732942936
transform -1 0 1196 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_62
timestamp 1732942936
transform -1 0 1244 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_20
timestamp 1732942936
transform 1 0 1236 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_17
timestamp 1732942936
transform -1 0 1292 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_49
timestamp 1732942936
transform 1 0 1292 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_164
timestamp 1732942936
transform 1 0 1244 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_145
timestamp 1732942936
transform -1 0 1300 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_204
timestamp 1732942936
transform -1 0 1324 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1732942936
transform 1 0 1340 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1732942936
transform -1 0 1420 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_101
timestamp 1732942936
transform -1 0 1460 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_241
timestamp 1732942936
transform 1 0 1460 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_2_0
timestamp 1732942936
transform -1 0 1492 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1732942936
transform -1 0 1500 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_178
timestamp 1732942936
transform -1 0 1548 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_89
timestamp 1732942936
transform 1 0 1420 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1732942936
transform -1 0 1548 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_30
timestamp 1732942936
transform 1 0 1548 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1732942936
transform -1 0 1604 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1732942936
transform -1 0 1700 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_2_0
timestamp 1732942936
transform 1 0 1548 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1732942936
transform 1 0 1556 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_180
timestamp 1732942936
transform 1 0 1564 0 -1 1705
box -2 -3 50 103
use AOI22X1  AOI22X1_30
timestamp 1732942936
transform -1 0 1652 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_261
timestamp 1732942936
transform 1 0 1700 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_190
timestamp 1732942936
transform 1 0 1652 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_232
timestamp 1732942936
transform -1 0 1708 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_175
timestamp 1732942936
transform 1 0 1708 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_14
timestamp 1732942936
transform 1 0 1724 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1732942936
transform -1 0 1780 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_176
timestamp 1732942936
transform 1 0 1780 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_177
timestamp 1732942936
transform 1 0 1756 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_219
timestamp 1732942936
transform -1 0 1828 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1732942936
transform -1 0 1924 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1732942936
transform -1 0 1924 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_281
timestamp 1732942936
transform 1 0 1924 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_230
timestamp 1732942936
transform -1 0 1980 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_158
timestamp 1732942936
transform 1 0 1980 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_3_0
timestamp 1732942936
transform -1 0 2020 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1732942936
transform -1 0 2028 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_150
timestamp 1732942936
transform 1 0 1924 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1732942936
transform -1 0 1980 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_182
timestamp 1732942936
transform 1 0 1980 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_178
timestamp 1732942936
transform -1 0 2052 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1732942936
transform -1 0 2148 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_3_0
timestamp 1732942936
transform 1 0 2028 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1732942936
transform 1 0 2036 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_179
timestamp 1732942936
transform 1 0 2044 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_70
timestamp 1732942936
transform 1 0 2092 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_251
timestamp 1732942936
transform 1 0 2116 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1732942936
transform -1 0 2244 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_206
timestamp 1732942936
transform -1 0 2172 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1732942936
transform -1 0 2268 0 -1 1705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_43
timestamp 1732942936
transform 1 0 2244 0 1 1505
box -2 -3 74 103
use OAI21X1  OAI21X1_6
timestamp 1732942936
transform 1 0 2316 0 1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_3
timestamp 1732942936
transform -1 0 2340 0 -1 1705
box -2 -3 74 103
use NAND2X1  NAND2X1_6
timestamp 1732942936
transform -1 0 2372 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1732942936
transform -1 0 2468 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1732942936
transform -1 0 2436 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_6
timestamp 1732942936
transform 1 0 2468 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_183
timestamp 1732942936
transform 1 0 2492 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_1
timestamp 1732942936
transform 1 0 2516 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_24
timestamp 1732942936
transform -1 0 2468 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1732942936
transform -1 0 2500 0 -1 1705
box -2 -3 34 103
use FILL  FILL_17_1
timestamp 1732942936
transform -1 0 2508 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_2
timestamp 1732942936
transform -1 0 2516 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_3
timestamp 1732942936
transform -1 0 2524 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1732942936
transform -1 0 100 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_87
timestamp 1732942936
transform -1 0 132 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_99
timestamp 1732942936
transform -1 0 156 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_28
timestamp 1732942936
transform 1 0 156 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_15
timestamp 1732942936
transform 1 0 180 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1732942936
transform -1 0 236 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1732942936
transform 1 0 236 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1732942936
transform -1 0 428 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_55
timestamp 1732942936
transform -1 0 460 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_0_0
timestamp 1732942936
transform 1 0 460 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1732942936
transform 1 0 468 0 1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_3
timestamp 1732942936
transform 1 0 476 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_198
timestamp 1732942936
transform -1 0 548 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_1
timestamp 1732942936
transform 1 0 548 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_189
timestamp 1732942936
transform 1 0 588 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_167
timestamp 1732942936
transform -1 0 644 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1732942936
transform -1 0 740 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_15
timestamp 1732942936
transform -1 0 788 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1732942936
transform 1 0 788 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_13
timestamp 1732942936
transform -1 0 932 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_57
timestamp 1732942936
transform -1 0 980 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_1_0
timestamp 1732942936
transform -1 0 988 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1732942936
transform -1 0 996 0 1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_56
timestamp 1732942936
transform -1 0 1044 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1732942936
transform -1 0 1140 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_11
timestamp 1732942936
transform 1 0 1140 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1732942936
transform -1 0 1196 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_144
timestamp 1732942936
transform -1 0 1220 0 1 1705
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1732942936
transform -1 0 1252 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_51
timestamp 1732942936
transform -1 0 1300 0 1 1705
box -2 -3 50 103
use AOI22X1  AOI22X1_9
timestamp 1732942936
transform 1 0 1300 0 1 1705
box -2 -3 42 103
use MUX2X1  MUX2X1_54
timestamp 1732942936
transform -1 0 1388 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_63
timestamp 1732942936
transform -1 0 1436 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_52
timestamp 1732942936
transform -1 0 1484 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_47
timestamp 1732942936
transform 1 0 1484 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_2_0
timestamp 1732942936
transform -1 0 1516 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1732942936
transform -1 0 1524 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_41
timestamp 1732942936
transform -1 0 1556 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1732942936
transform -1 0 1652 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_61
timestamp 1732942936
transform -1 0 1700 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_146
timestamp 1732942936
transform 1 0 1700 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_129
timestamp 1732942936
transform -1 0 1756 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1732942936
transform -1 0 1852 0 1 1705
box -2 -3 98 103
use BUFX4  BUFX4_57
timestamp 1732942936
transform 1 0 1852 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1732942936
transform 1 0 1884 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_183
timestamp 1732942936
transform 1 0 1980 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_3_0
timestamp 1732942936
transform -1 0 2036 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1732942936
transform -1 0 2044 0 1 1705
box -2 -3 10 103
use AOI22X1  AOI22X1_29
timestamp 1732942936
transform -1 0 2084 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_62
timestamp 1732942936
transform 1 0 2084 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1732942936
transform -1 0 2212 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_171
timestamp 1732942936
transform -1 0 2260 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_169
timestamp 1732942936
transform 1 0 2260 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_172
timestamp 1732942936
transform -1 0 2356 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_52
timestamp 1732942936
transform 1 0 2356 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1732942936
transform -1 0 2476 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_22
timestamp 1732942936
transform 1 0 2476 0 1 1705
box -2 -3 34 103
use FILL  FILL_18_1
timestamp 1732942936
transform 1 0 2508 0 1 1705
box -2 -3 10 103
use FILL  FILL_18_2
timestamp 1732942936
transform 1 0 2516 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_246
timestamp 1732942936
transform 1 0 4 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_201
timestamp 1732942936
transform -1 0 60 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_57
timestamp 1732942936
transform 1 0 60 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1732942936
transform -1 0 116 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_59
timestamp 1732942936
transform -1 0 164 0 -1 1905
box -2 -3 50 103
use CLKBUF1  CLKBUF1_29
timestamp 1732942936
transform -1 0 236 0 -1 1905
box -2 -3 74 103
use MUX2X1  MUX2X1_1
timestamp 1732942936
transform -1 0 284 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_60
timestamp 1732942936
transform -1 0 332 0 -1 1905
box -2 -3 50 103
use CLKBUF1  CLKBUF1_30
timestamp 1732942936
transform -1 0 404 0 -1 1905
box -2 -3 74 103
use NOR2X1  NOR2X1_11
timestamp 1732942936
transform 1 0 404 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1732942936
transform -1 0 460 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_0_0
timestamp 1732942936
transform -1 0 468 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1732942936
transform -1 0 476 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1732942936
transform -1 0 572 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_2
timestamp 1732942936
transform 1 0 572 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_4
timestamp 1732942936
transform -1 0 668 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_6
timestamp 1732942936
transform 1 0 668 0 -1 1905
box -2 -3 50 103
use AOI22X1  AOI22X1_3
timestamp 1732942936
transform -1 0 756 0 -1 1905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1732942936
transform 1 0 756 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_274
timestamp 1732942936
transform 1 0 852 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_223
timestamp 1732942936
transform -1 0 908 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_284
timestamp 1732942936
transform 1 0 908 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_231
timestamp 1732942936
transform -1 0 964 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_8
timestamp 1732942936
transform -1 0 1012 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_1_0
timestamp 1732942936
transform 1 0 1012 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1732942936
transform 1 0 1020 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1732942936
transform 1 0 1028 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_9
timestamp 1732942936
transform 1 0 1124 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1732942936
transform -1 0 1180 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_127
timestamp 1732942936
transform 1 0 1180 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1732942936
transform -1 0 1308 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_177
timestamp 1732942936
transform 1 0 1308 0 -1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_24
timestamp 1732942936
transform -1 0 1412 0 -1 1905
box -2 -3 74 103
use NOR2X1  NOR2X1_23
timestamp 1732942936
transform 1 0 1412 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1732942936
transform -1 0 1468 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_205
timestamp 1732942936
transform -1 0 1492 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_2_0
timestamp 1732942936
transform 1 0 1492 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1732942936
transform 1 0 1500 0 -1 1905
box -2 -3 10 103
use AOI22X1  AOI22X1_11
timestamp 1732942936
transform 1 0 1508 0 -1 1905
box -2 -3 42 103
use BUFX4  BUFX4_15
timestamp 1732942936
transform 1 0 1548 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_155
timestamp 1732942936
transform -1 0 1604 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1732942936
transform 1 0 1604 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_1
timestamp 1732942936
transform 1 0 1628 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1732942936
transform -1 0 1756 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_53
timestamp 1732942936
transform 1 0 1756 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_33
timestamp 1732942936
transform 1 0 1804 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1732942936
transform -1 0 1860 0 -1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_31
timestamp 1732942936
transform -1 0 1900 0 -1 1905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1732942936
transform -1 0 1996 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_115
timestamp 1732942936
transform -1 0 2020 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_3_0
timestamp 1732942936
transform -1 0 2028 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1732942936
transform -1 0 2036 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1732942936
transform -1 0 2132 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_124
timestamp 1732942936
transform 1 0 2132 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_181
timestamp 1732942936
transform 1 0 2156 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_174
timestamp 1732942936
transform -1 0 2252 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_94
timestamp 1732942936
transform 1 0 2252 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1732942936
transform -1 0 2308 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1732942936
transform 1 0 2308 0 -1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_44
timestamp 1732942936
transform -1 0 2476 0 -1 1905
box -2 -3 74 103
use BUFX4  BUFX4_58
timestamp 1732942936
transform -1 0 2508 0 -1 1905
box -2 -3 34 103
use FILL  FILL_19_1
timestamp 1732942936
transform -1 0 2516 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_2
timestamp 1732942936
transform -1 0 2524 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1732942936
transform -1 0 100 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1732942936
transform 1 0 100 0 1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_41
timestamp 1732942936
transform -1 0 268 0 1 1905
box -2 -3 74 103
use NAND2X1  NAND2X1_180
timestamp 1732942936
transform 1 0 268 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_159
timestamp 1732942936
transform -1 0 324 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1732942936
transform 1 0 324 0 1 1905
box -2 -3 98 103
use BUFX4  BUFX4_19
timestamp 1732942936
transform -1 0 452 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_16
timestamp 1732942936
transform 1 0 452 0 1 1905
box -2 -3 50 103
use FILL  FILL_19_0_0
timestamp 1732942936
transform 1 0 500 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1732942936
transform 1 0 508 0 1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_18
timestamp 1732942936
transform 1 0 516 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_45
timestamp 1732942936
transform 1 0 564 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_39
timestamp 1732942936
transform -1 0 620 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_175
timestamp 1732942936
transform 1 0 620 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1732942936
transform 1 0 652 0 1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_199
timestamp 1732942936
transform -1 0 716 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_23
timestamp 1732942936
transform -1 0 748 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1732942936
transform 1 0 748 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1732942936
transform -1 0 812 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1732942936
transform -1 0 908 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_24
timestamp 1732942936
transform -1 0 956 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_31
timestamp 1732942936
transform 1 0 956 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_1_0
timestamp 1732942936
transform -1 0 996 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1732942936
transform -1 0 1004 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_36
timestamp 1732942936
transform -1 0 1028 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1732942936
transform -1 0 1124 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_65
timestamp 1732942936
transform -1 0 1172 0 1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1732942936
transform -1 0 1268 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_66
timestamp 1732942936
transform -1 0 1316 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_64
timestamp 1732942936
transform -1 0 1364 0 1 1905
box -2 -3 50 103
use AOI22X1  AOI22X1_12
timestamp 1732942936
transform 1 0 1364 0 1 1905
box -2 -3 42 103
use MUX2X1  MUX2X1_72
timestamp 1732942936
transform -1 0 1452 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_137
timestamp 1732942936
transform 1 0 1452 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1732942936
transform 1 0 1484 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1732942936
transform 1 0 1492 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1732942936
transform 1 0 1500 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1732942936
transform -1 0 1692 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_182
timestamp 1732942936
transform 1 0 1692 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_161
timestamp 1732942936
transform -1 0 1748 0 1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_48
timestamp 1732942936
transform -1 0 1820 0 1 1905
box -2 -3 74 103
use OAI21X1  OAI21X1_182
timestamp 1732942936
transform -1 0 1852 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1732942936
transform -1 0 1876 0 1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_32
timestamp 1732942936
transform -1 0 1916 0 1 1905
box -2 -3 42 103
use MUX2X1  MUX2X1_192
timestamp 1732942936
transform 1 0 1916 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_190
timestamp 1732942936
transform -1 0 2012 0 1 1905
box -2 -3 50 103
use FILL  FILL_19_3_0
timestamp 1732942936
transform -1 0 2020 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1732942936
transform -1 0 2028 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1732942936
transform -1 0 2124 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_110
timestamp 1732942936
transform 1 0 2124 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1732942936
transform 1 0 2156 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1732942936
transform -1 0 2212 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1732942936
transform -1 0 2308 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_134
timestamp 1732942936
transform 1 0 2308 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1732942936
transform -1 0 2436 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_170
timestamp 1732942936
transform -1 0 2468 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_55
timestamp 1732942936
transform 1 0 2468 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1732942936
transform 1 0 2500 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1732942936
transform 1 0 2508 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_3
timestamp 1732942936
transform 1 0 2516 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1732942936
transform -1 0 100 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_209
timestamp 1732942936
transform 1 0 100 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_256
timestamp 1732942936
transform -1 0 156 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_73
timestamp 1732942936
transform 1 0 156 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_83
timestamp 1732942936
transform -1 0 212 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_58
timestamp 1732942936
transform 1 0 212 0 -1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1732942936
transform -1 0 356 0 -1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_236
timestamp 1732942936
transform 1 0 356 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_193
timestamp 1732942936
transform -1 0 412 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1732942936
transform 1 0 412 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_0_0
timestamp 1732942936
transform -1 0 516 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1732942936
transform -1 0 524 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_197
timestamp 1732942936
transform -1 0 548 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1732942936
transform 1 0 548 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_67
timestamp 1732942936
transform -1 0 628 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_74
timestamp 1732942936
transform 1 0 628 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1732942936
transform -1 0 748 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_3
timestamp 1732942936
transform 1 0 748 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_126
timestamp 1732942936
transform 1 0 772 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1732942936
transform 1 0 796 0 -1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_23
timestamp 1732942936
transform 1 0 892 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_5
timestamp 1732942936
transform -1 0 988 0 -1 2105
box -2 -3 50 103
use FILL  FILL_20_1_0
timestamp 1732942936
transform 1 0 988 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1732942936
transform 1 0 996 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_54
timestamp 1732942936
transform 1 0 1004 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1732942936
transform -1 0 1124 0 -1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_69
timestamp 1732942936
transform 1 0 1124 0 -1 2105
box -2 -3 50 103
use BUFX4  BUFX4_17
timestamp 1732942936
transform 1 0 1172 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1732942936
transform 1 0 1204 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_50
timestamp 1732942936
transform 1 0 1236 0 -1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1732942936
transform -1 0 1380 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_5
timestamp 1732942936
transform 1 0 1380 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1732942936
transform -1 0 1436 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1732942936
transform -1 0 1460 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1732942936
transform -1 0 1492 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_2_0
timestamp 1732942936
transform 1 0 1492 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1732942936
transform 1 0 1500 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1732942936
transform 1 0 1508 0 -1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_71
timestamp 1732942936
transform 1 0 1604 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_49
timestamp 1732942936
transform 1 0 1652 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1732942936
transform -1 0 1708 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1732942936
transform 1 0 1708 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_32
timestamp 1732942936
transform -1 0 1836 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_186
timestamp 1732942936
transform -1 0 1884 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_184
timestamp 1732942936
transform -1 0 1932 0 -1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_18
timestamp 1732942936
transform -1 0 1956 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1732942936
transform -1 0 1988 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1732942936
transform 1 0 1988 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_3_0
timestamp 1732942936
transform -1 0 2028 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1732942936
transform -1 0 2036 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1732942936
transform -1 0 2132 0 -1 2105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_2
timestamp 1732942936
transform -1 0 2204 0 -1 2105
box -2 -3 74 103
use MUX2X1  MUX2X1_191
timestamp 1732942936
transform -1 0 2252 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_170
timestamp 1732942936
transform 1 0 2252 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_133
timestamp 1732942936
transform 1 0 2300 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1732942936
transform -1 0 2420 0 -1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_187
timestamp 1732942936
transform 1 0 2420 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1732942936
transform 1 0 2444 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1732942936
transform 1 0 2468 0 -1 2105
box -2 -3 34 103
use FILL  FILL_21_1
timestamp 1732942936
transform -1 0 2508 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_2
timestamp 1732942936
transform -1 0 2516 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_3
timestamp 1732942936
transform -1 0 2524 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1732942936
transform -1 0 100 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_185
timestamp 1732942936
transform 1 0 100 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_227
timestamp 1732942936
transform -1 0 156 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1732942936
transform 1 0 156 0 1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_17
timestamp 1732942936
transform -1 0 300 0 1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_21
timestamp 1732942936
transform -1 0 324 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1732942936
transform -1 0 356 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1732942936
transform -1 0 452 0 1 2105
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1732942936
transform -1 0 476 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_0_0
timestamp 1732942936
transform -1 0 484 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1732942936
transform -1 0 492 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1732942936
transform -1 0 588 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1732942936
transform -1 0 684 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_65
timestamp 1732942936
transform -1 0 716 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1732942936
transform 1 0 716 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1732942936
transform 1 0 748 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1732942936
transform -1 0 812 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1732942936
transform 1 0 812 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_119
timestamp 1732942936
transform 1 0 908 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1732942936
transform 1 0 940 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_55
timestamp 1732942936
transform -1 0 1012 0 1 2105
box -2 -3 50 103
use FILL  FILL_21_1_0
timestamp 1732942936
transform -1 0 1020 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1732942936
transform -1 0 1028 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_47
timestamp 1732942936
transform -1 0 1060 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1732942936
transform 1 0 1060 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1732942936
transform -1 0 1180 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_203
timestamp 1732942936
transform 1 0 1180 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1732942936
transform -1 0 1300 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_169
timestamp 1732942936
transform 1 0 1300 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_191
timestamp 1732942936
transform -1 0 1356 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1732942936
transform 1 0 1356 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1732942936
transform -1 0 1548 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_2_0
timestamp 1732942936
transform 1 0 1548 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1732942936
transform 1 0 1556 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_113
timestamp 1732942936
transform 1 0 1564 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_128
timestamp 1732942936
transform -1 0 1620 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_121
timestamp 1732942936
transform 1 0 1620 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_137
timestamp 1732942936
transform -1 0 1676 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1732942936
transform 1 0 1676 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_56
timestamp 1732942936
transform -1 0 1804 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_218
timestamp 1732942936
transform 1 0 1804 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1732942936
transform -1 0 1924 0 1 2105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_34
timestamp 1732942936
transform 1 0 1924 0 1 2105
box -2 -3 74 103
use BUFX4  BUFX4_59
timestamp 1732942936
transform 1 0 1996 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_3_0
timestamp 1732942936
transform 1 0 2028 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1732942936
transform 1 0 2036 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_54
timestamp 1732942936
transform 1 0 2044 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1732942936
transform -1 0 2100 0 1 2105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_1
timestamp 1732942936
transform 1 0 2100 0 1 2105
box -2 -3 74 103
use NAND2X1  NAND2X1_142
timestamp 1732942936
transform -1 0 2196 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_126
timestamp 1732942936
transform -1 0 2228 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1732942936
transform 1 0 2228 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_118
timestamp 1732942936
transform -1 0 2356 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_196
timestamp 1732942936
transform 1 0 2356 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_174
timestamp 1732942936
transform -1 0 2412 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1732942936
transform -1 0 2508 0 1 2105
box -2 -3 98 103
use FILL  FILL_22_1
timestamp 1732942936
transform 1 0 2508 0 1 2105
box -2 -3 10 103
use FILL  FILL_22_2
timestamp 1732942936
transform 1 0 2516 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1732942936
transform -1 0 100 0 -1 2305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_22
timestamp 1732942936
transform -1 0 172 0 -1 2305
box -2 -3 74 103
use OAI21X1  OAI21X1_63
timestamp 1732942936
transform 1 0 172 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_72
timestamp 1732942936
transform -1 0 228 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1732942936
transform 1 0 228 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_19
timestamp 1732942936
transform 1 0 324 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_79
timestamp 1732942936
transform 1 0 372 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_90
timestamp 1732942936
transform -1 0 428 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1732942936
transform 1 0 428 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_0_0
timestamp 1732942936
transform 1 0 524 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1732942936
transform 1 0 532 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_20
timestamp 1732942936
transform 1 0 540 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_21
timestamp 1732942936
transform 1 0 588 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_7
timestamp 1732942936
transform 1 0 636 0 -1 2305
box -2 -3 50 103
use CLKBUF1  CLKBUF1_32
timestamp 1732942936
transform 1 0 684 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1732942936
transform -1 0 852 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_225
timestamp 1732942936
transform 1 0 852 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_183
timestamp 1732942936
transform -1 0 908 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_22
timestamp 1732942936
transform -1 0 956 0 -1 2305
box -2 -3 50 103
use FILL  FILL_22_1_0
timestamp 1732942936
transform -1 0 964 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1732942936
transform -1 0 972 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1732942936
transform -1 0 1068 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_95
timestamp 1732942936
transform 1 0 1068 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_108
timestamp 1732942936
transform 1 0 1100 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_25
timestamp 1732942936
transform -1 0 1156 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1732942936
transform 1 0 1156 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_35
timestamp 1732942936
transform -1 0 1212 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_266
timestamp 1732942936
transform -1 0 1236 0 -1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_68
timestamp 1732942936
transform -1 0 1284 0 -1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1732942936
transform -1 0 1380 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_81
timestamp 1732942936
transform 1 0 1380 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1732942936
transform 1 0 1412 0 -1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_70
timestamp 1732942936
transform -1 0 1484 0 -1 2305
box -2 -3 50 103
use FILL  FILL_22_2_0
timestamp 1732942936
transform -1 0 1492 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1732942936
transform -1 0 1500 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1732942936
transform -1 0 1596 0 -1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_24
timestamp 1732942936
transform 1 0 1596 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1732942936
transform -1 0 1652 0 -1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_21
timestamp 1732942936
transform -1 0 1724 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1732942936
transform 1 0 1724 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_185
timestamp 1732942936
transform 1 0 1820 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_187
timestamp 1732942936
transform -1 0 1916 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_189
timestamp 1732942936
transform 1 0 1916 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_70
timestamp 1732942936
transform 1 0 1964 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1732942936
transform -1 0 2020 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_3_0
timestamp 1732942936
transform 1 0 2020 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1732942936
transform 1 0 2028 0 -1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_43
timestamp 1732942936
transform 1 0 2036 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1732942936
transform 1 0 2060 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_173
timestamp 1732942936
transform 1 0 2156 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_188
timestamp 1732942936
transform -1 0 2252 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_86
timestamp 1732942936
transform 1 0 2252 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_97
timestamp 1732942936
transform -1 0 2308 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1732942936
transform -1 0 2404 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1732942936
transform -1 0 2500 0 -1 2305
box -2 -3 98 103
use FILL  FILL_23_1
timestamp 1732942936
transform -1 0 2508 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_2
timestamp 1732942936
transform -1 0 2516 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_3
timestamp 1732942936
transform -1 0 2524 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_35
timestamp 1732942936
transform 1 0 4 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_33
timestamp 1732942936
transform -1 0 60 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_71
timestamp 1732942936
transform 1 0 60 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_81
timestamp 1732942936
transform -1 0 116 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1732942936
transform -1 0 212 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_21
timestamp 1732942936
transform -1 0 244 0 1 2305
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1732942936
transform 1 0 244 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_23
timestamp 1732942936
transform 1 0 284 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1732942936
transform -1 0 340 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1732942936
transform 1 0 340 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_0_0
timestamp 1732942936
transform -1 0 444 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1732942936
transform -1 0 452 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1732942936
transform -1 0 548 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_264
timestamp 1732942936
transform 1 0 548 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_215
timestamp 1732942936
transform -1 0 604 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1732942936
transform 1 0 604 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_117
timestamp 1732942936
transform 1 0 700 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_103
timestamp 1732942936
transform -1 0 756 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1732942936
transform -1 0 852 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_16
timestamp 1732942936
transform 1 0 852 0 1 2305
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1732942936
transform -1 0 908 0 1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_23
timestamp 1732942936
transform 1 0 908 0 1 2305
box -2 -3 74 103
use FILL  FILL_23_1_0
timestamp 1732942936
transform 1 0 980 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1732942936
transform 1 0 988 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1732942936
transform 1 0 996 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_217
timestamp 1732942936
transform 1 0 1092 0 1 2305
box -2 -3 34 103
use INVX8  INVX8_3
timestamp 1732942936
transform -1 0 1164 0 1 2305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1732942936
transform 1 0 1164 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_119
timestamp 1732942936
transform 1 0 1260 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_105
timestamp 1732942936
transform -1 0 1316 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1732942936
transform 1 0 1316 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_110
timestamp 1732942936
transform -1 0 1372 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1732942936
transform 1 0 1372 0 1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_40
timestamp 1732942936
transform 1 0 1468 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_2_0
timestamp 1732942936
transform -1 0 1508 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1732942936
transform -1 0 1516 0 1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_42
timestamp 1732942936
transform -1 0 1540 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1732942936
transform -1 0 1564 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_78
timestamp 1732942936
transform 1 0 1564 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_88
timestamp 1732942936
transform -1 0 1620 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1732942936
transform -1 0 1716 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1732942936
transform -1 0 1812 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1732942936
transform 1 0 1812 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_38
timestamp 1732942936
transform 1 0 1908 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1732942936
transform 1 0 1940 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_3_0
timestamp 1732942936
transform 1 0 2036 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1732942936
transform 1 0 2044 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_271
timestamp 1732942936
transform 1 0 2052 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_222
timestamp 1732942936
transform -1 0 2108 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1732942936
transform 1 0 2108 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_267
timestamp 1732942936
transform -1 0 2228 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1732942936
transform 1 0 2228 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1732942936
transform 1 0 2324 0 1 2305
box -2 -3 98 103
use INVX8  INVX8_8
timestamp 1732942936
transform -1 0 2460 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_90
timestamp 1732942936
transform 1 0 2460 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1732942936
transform -1 0 2516 0 1 2305
box -2 -3 26 103
use FILL  FILL_24_1
timestamp 1732942936
transform 1 0 2516 0 1 2305
box -2 -3 10 103
<< labels >>
flabel metal6 s 480 -30 496 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 984 -30 1000 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1422 -22 1426 -18 7 FreeSans 24 270 0 0 enable
port 2 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 clk
port 3 nsew
flabel metal2 s 1806 2428 1810 2432 3 FreeSans 24 90 0 0 r_w
port 4 nsew
flabel metal2 s 262 2428 266 2432 3 FreeSans 24 90 0 0 datain[0]
port 5 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 0 0 0 datain[1]
port 6 nsew
flabel metal2 s 1142 2428 1146 2432 3 FreeSans 24 90 0 0 datain[2]
port 7 nsew
flabel metal3 s 2550 68 2554 72 3 FreeSans 24 0 0 0 datain[3]
port 8 nsew
flabel metal2 s 422 -22 426 -18 7 FreeSans 24 270 0 0 datain[4]
port 9 nsew
flabel metal3 s 2550 48 2554 52 3 FreeSans 24 270 0 0 datain[5]
port 10 nsew
flabel metal2 s 878 -22 882 -18 7 FreeSans 24 270 0 0 datain[6]
port 11 nsew
flabel metal3 s 2550 2348 2554 2352 3 FreeSans 24 90 0 0 datain[7]
port 12 nsew
flabel metal2 s 2038 -22 2042 -18 7 FreeSans 24 270 0 0 address[0]
port 13 nsew
flabel metal2 s 1654 -22 1658 -18 7 FreeSans 24 270 0 0 address[1]
port 14 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 address[2]
port 15 nsew
flabel metal3 s -26 1448 -22 1452 7 FreeSans 24 0 0 0 address[3]
port 16 nsew
flabel metal3 s -26 1468 -22 1472 7 FreeSans 24 0 0 0 address[4]
port 17 nsew
flabel metal2 s 462 2428 466 2432 3 FreeSans 24 90 0 0 dataout[0]
port 18 nsew
flabel metal2 s 918 2428 922 2432 3 FreeSans 24 90 0 0 dataout[1]
port 19 nsew
flabel metal2 s 894 2428 898 2432 3 FreeSans 24 90 0 0 dataout[2]
port 20 nsew
flabel metal3 s 2550 1048 2554 1052 3 FreeSans 24 0 0 0 dataout[3]
port 21 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 dataout[4]
port 22 nsew
flabel metal3 s -26 748 -22 752 7 FreeSans 24 0 0 0 dataout[5]
port 23 nsew
flabel metal2 s 518 -22 522 -18 7 FreeSans 24 270 0 0 dataout[6]
port 24 nsew
flabel metal2 s 1550 2428 1554 2432 3 FreeSans 24 90 0 0 dataout[7]
port 25 nsew
<< end >>
