magic
tech scmos
timestamp 1732942776
<< metal1 >>
rect 544 2403 546 2407
rect 550 2403 553 2407
rect 557 2403 560 2407
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1573 2403 1576 2407
rect 1374 2368 1382 2371
rect 646 2351 649 2361
rect 1086 2358 1094 2361
rect 626 2348 633 2351
rect 646 2348 665 2351
rect 878 2348 897 2351
rect 966 2348 974 2351
rect 1034 2348 1041 2351
rect 1046 2348 1078 2351
rect 1166 2348 1182 2351
rect 1254 2351 1257 2361
rect 1254 2348 1273 2351
rect 1406 2351 1409 2361
rect 1614 2358 1633 2361
rect 1390 2348 1409 2351
rect 1430 2348 1441 2351
rect 1538 2348 1553 2351
rect 1430 2342 1433 2348
rect 1830 2351 1833 2361
rect 1842 2358 1846 2362
rect 1790 2348 1801 2351
rect 1814 2348 1833 2351
rect 538 2338 553 2341
rect 890 2338 897 2341
rect 1054 2338 1078 2341
rect 1402 2338 1409 2341
rect 1462 2338 1481 2341
rect 1798 2341 1801 2348
rect 2002 2348 2017 2351
rect 2066 2348 2073 2351
rect 2238 2351 2241 2361
rect 2238 2348 2257 2351
rect 2374 2348 2382 2351
rect 2490 2348 2497 2351
rect 1798 2338 1806 2341
rect 606 2332 610 2334
rect 862 2331 866 2333
rect 862 2328 870 2331
rect 1462 2328 1465 2338
rect 1778 2318 1779 2322
rect 1056 2303 1058 2307
rect 1062 2303 1065 2307
rect 1069 2303 1072 2307
rect 2080 2303 2082 2307
rect 2086 2303 2089 2307
rect 2093 2303 2096 2307
rect 1138 2288 1139 2292
rect 198 2278 217 2281
rect 846 2278 865 2281
rect 1734 2278 1753 2281
rect 1958 2278 1977 2281
rect 2106 2278 2121 2281
rect 2126 2278 2145 2281
rect 434 2268 449 2271
rect 690 2268 697 2271
rect 1118 2268 1129 2271
rect 1178 2268 1185 2271
rect 1362 2268 1369 2271
rect 1562 2268 1593 2271
rect 1854 2271 1858 2274
rect 1786 2268 1793 2271
rect 1846 2268 1858 2271
rect 110 2258 126 2261
rect 358 2258 377 2261
rect 386 2258 393 2261
rect 694 2261 697 2268
rect 662 2258 681 2261
rect 694 2258 705 2261
rect 998 2258 1006 2261
rect 1118 2261 1121 2268
rect 1114 2258 1121 2261
rect 1226 2258 1233 2261
rect 1350 2258 1366 2261
rect 1374 2258 1393 2261
rect 1846 2262 1849 2268
rect 1774 2258 1782 2261
rect 1906 2258 1913 2261
rect 2206 2258 2214 2261
rect 2382 2258 2401 2261
rect 2422 2258 2441 2261
rect 662 2248 665 2258
rect 1390 2248 1393 2258
rect 1402 2248 1406 2252
rect 2382 2248 2385 2258
rect 2438 2248 2441 2258
rect 299 2238 302 2242
rect 346 2238 347 2242
rect 1054 2238 1070 2241
rect 410 2218 411 2222
rect 717 2218 718 2222
rect 1538 2218 1539 2222
rect 544 2203 546 2207
rect 550 2203 553 2207
rect 557 2203 560 2207
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1573 2203 1576 2207
rect 1845 2188 1846 2192
rect 555 2168 558 2172
rect 706 2168 713 2171
rect 2378 2168 2381 2172
rect 126 2142 129 2151
rect 374 2151 377 2161
rect 202 2148 217 2151
rect 358 2148 377 2151
rect 518 2148 534 2151
rect 622 2151 625 2161
rect 606 2148 625 2151
rect 678 2151 681 2161
rect 678 2148 697 2151
rect 742 2148 750 2151
rect 1386 2148 1393 2151
rect 1798 2151 1801 2161
rect 1782 2148 1801 2151
rect 1958 2151 1961 2161
rect 1958 2148 1977 2151
rect 2034 2148 2049 2151
rect 2154 2148 2161 2151
rect 398 2138 414 2141
rect 574 2138 601 2141
rect 650 2138 657 2141
rect 678 2138 686 2141
rect 894 2138 906 2141
rect 1002 2138 1009 2141
rect 1186 2138 1193 2141
rect 1717 2138 1718 2142
rect 1794 2138 1801 2141
rect 2090 2138 2106 2141
rect 574 2136 578 2138
rect 110 2128 129 2131
rect 1142 2128 1145 2138
rect 2390 2132 2393 2142
rect 2446 2138 2458 2141
rect 2526 2132 2530 2136
rect 1166 2128 1185 2131
rect 574 2118 590 2121
rect 1056 2103 1058 2107
rect 1062 2103 1065 2107
rect 1069 2103 1072 2107
rect 2080 2103 2082 2107
rect 2086 2103 2089 2107
rect 2093 2103 2096 2107
rect 197 2088 198 2092
rect 2109 2088 2110 2092
rect 434 2078 435 2082
rect 630 2078 641 2081
rect 630 2077 634 2078
rect 638 2072 641 2078
rect 750 2072 753 2081
rect 758 2078 777 2081
rect 2142 2078 2161 2081
rect 2454 2078 2466 2081
rect 2462 2077 2466 2078
rect 138 2068 145 2071
rect 530 2068 546 2071
rect 658 2068 665 2071
rect 1222 2071 1226 2074
rect 1214 2068 1226 2071
rect 1622 2068 1630 2071
rect 2430 2068 2438 2071
rect 38 2058 46 2061
rect 118 2058 137 2061
rect 158 2058 185 2061
rect 226 2058 233 2061
rect 446 2058 465 2061
rect 510 2058 518 2061
rect 646 2058 665 2061
rect 838 2058 846 2061
rect 1102 2058 1110 2061
rect 1190 2058 1209 2061
rect 1438 2058 1457 2061
rect 1502 2058 1510 2061
rect 1514 2058 1521 2061
rect 1534 2058 1542 2061
rect 1566 2058 1598 2061
rect 1622 2058 1641 2061
rect 1686 2058 1694 2061
rect 1794 2058 1809 2061
rect 1966 2058 1985 2061
rect 2038 2058 2046 2061
rect 2062 2058 2097 2061
rect 2182 2058 2185 2068
rect 2222 2058 2230 2061
rect 2254 2058 2273 2061
rect 2354 2058 2361 2061
rect 2430 2058 2449 2061
rect 134 2052 137 2058
rect 1190 2048 1193 2058
rect 1438 2048 1441 2058
rect 1518 2048 1521 2058
rect 1530 2048 1534 2052
rect 1622 2048 1625 2058
rect 1966 2048 1969 2058
rect 2270 2048 2273 2058
rect 1426 2038 1427 2042
rect 1650 2038 1657 2041
rect 293 2018 294 2022
rect 498 2018 499 2022
rect 725 2018 726 2022
rect 954 2018 955 2022
rect 1090 2018 1091 2022
rect 2026 2018 2027 2022
rect 2210 2018 2211 2022
rect 544 2003 546 2007
rect 550 2003 553 2007
rect 557 2003 560 2007
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1573 2003 1576 2007
rect 1781 1988 1782 1992
rect 1845 1988 1846 1992
rect 2482 1988 2483 1992
rect 2626 1988 2627 1992
rect 1106 1968 1109 1972
rect 1610 1968 1617 1971
rect 2322 1968 2329 1971
rect 2538 1968 2541 1972
rect 6 1938 9 1948
rect 198 1942 201 1951
rect 254 1951 257 1961
rect 266 1958 270 1962
rect 958 1953 962 1958
rect 238 1948 257 1951
rect 494 1948 518 1951
rect 578 1948 585 1951
rect 910 1948 929 1951
rect 1062 1948 1078 1951
rect 1206 1951 1209 1961
rect 1278 1958 1297 1961
rect 1306 1958 1310 1962
rect 1566 1958 1574 1961
rect 1190 1948 1209 1951
rect 1470 1948 1481 1951
rect 1558 1948 1582 1951
rect 1750 1948 1769 1951
rect 1830 1951 1833 1961
rect 1814 1948 1833 1951
rect 1894 1948 1913 1951
rect 2158 1951 2161 1961
rect 502 1938 510 1941
rect 646 1938 665 1941
rect 910 1938 918 1941
rect 1234 1938 1249 1941
rect 1470 1941 1473 1948
rect 2142 1948 2161 1951
rect 2294 1951 2297 1961
rect 2638 1958 2646 1961
rect 2274 1948 2281 1951
rect 2294 1948 2313 1951
rect 2498 1948 2505 1951
rect 1454 1938 1473 1941
rect 1578 1938 1601 1941
rect 1894 1938 1902 1941
rect 2122 1938 2137 1941
rect 2154 1938 2161 1941
rect 2294 1938 2302 1941
rect 2454 1938 2462 1941
rect 150 1932 154 1936
rect 166 1931 170 1933
rect 166 1928 177 1931
rect 182 1928 201 1931
rect 646 1928 649 1938
rect 942 1931 946 1933
rect 934 1928 946 1931
rect 1926 1931 1930 1933
rect 1922 1928 1930 1931
rect 2518 1931 2522 1933
rect 2514 1928 2522 1931
rect 2210 1918 2211 1922
rect 1056 1903 1058 1907
rect 1062 1903 1065 1907
rect 1069 1903 1072 1907
rect 2080 1903 2082 1907
rect 2086 1903 2089 1907
rect 2093 1903 2096 1907
rect 482 1888 483 1892
rect 2613 1888 2614 1892
rect 94 1878 105 1881
rect 141 1878 142 1882
rect 282 1878 283 1882
rect 442 1878 443 1882
rect 2005 1878 2006 1882
rect 94 1877 98 1878
rect 1518 1872 1522 1874
rect 526 1868 550 1871
rect 710 1868 718 1871
rect 1178 1868 1185 1871
rect 1666 1868 1673 1871
rect 1918 1868 1937 1871
rect 2126 1868 2134 1871
rect 2338 1868 2345 1871
rect 102 1861 105 1868
rect 94 1858 105 1861
rect 294 1858 313 1861
rect 638 1858 646 1861
rect 710 1858 729 1861
rect 894 1858 913 1861
rect 954 1858 961 1861
rect 1038 1858 1046 1861
rect 1166 1858 1185 1861
rect 1406 1858 1425 1861
rect 1582 1858 1598 1861
rect 1654 1858 1673 1861
rect 1714 1858 1721 1861
rect 1802 1858 1809 1861
rect 1934 1861 1937 1868
rect 2382 1862 2385 1871
rect 2622 1868 2638 1871
rect 1934 1858 1945 1861
rect 2222 1858 2238 1861
rect 2326 1858 2334 1861
rect 2390 1858 2409 1861
rect 2422 1858 2430 1861
rect 94 1857 98 1858
rect 1182 1848 1185 1858
rect 1406 1848 1409 1858
rect 2406 1848 2409 1858
rect 2418 1848 2422 1852
rect 1619 1838 1622 1842
rect 349 1818 350 1822
rect 397 1818 398 1822
rect 973 1818 974 1822
rect 1733 1818 1734 1822
rect 1826 1818 1827 1822
rect 1957 1818 1958 1822
rect 544 1803 546 1807
rect 550 1803 553 1807
rect 557 1803 560 1807
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1573 1803 1576 1807
rect 317 1778 318 1782
rect 525 1768 526 1772
rect 2062 1768 2070 1771
rect 2378 1768 2385 1771
rect 1526 1766 1530 1768
rect 182 1748 190 1751
rect 198 1748 209 1751
rect 286 1748 294 1751
rect 362 1748 369 1751
rect 498 1748 513 1751
rect 562 1748 569 1751
rect 598 1748 609 1751
rect 686 1751 689 1761
rect 1054 1758 1062 1761
rect 1838 1753 1842 1758
rect 670 1748 689 1751
rect 770 1748 777 1751
rect 198 1741 201 1748
rect 182 1738 201 1741
rect 358 1738 366 1741
rect 390 1738 398 1741
rect 606 1741 609 1748
rect 606 1738 625 1741
rect 838 1738 846 1741
rect 982 1741 985 1751
rect 1138 1748 1145 1751
rect 1438 1748 1457 1751
rect 1526 1748 1537 1751
rect 1670 1748 1689 1751
rect 1526 1742 1529 1748
rect 2114 1748 2121 1751
rect 2154 1748 2161 1751
rect 2190 1748 2198 1751
rect 2294 1751 2297 1761
rect 2306 1758 2310 1762
rect 2282 1748 2297 1751
rect 982 1738 1001 1741
rect 1058 1738 1089 1741
rect 1146 1738 1153 1741
rect 1306 1738 1313 1741
rect 1318 1738 1326 1741
rect 1450 1738 1457 1741
rect 1682 1738 1689 1741
rect 2622 1738 2638 1741
rect 221 1728 222 1732
rect 1286 1728 1305 1731
rect 1406 1731 1410 1736
rect 1394 1728 1410 1731
rect 1422 1731 1426 1733
rect 1422 1728 1433 1731
rect 1654 1731 1658 1733
rect 1654 1728 1665 1731
rect 349 1718 350 1722
rect 389 1718 390 1722
rect 429 1718 430 1722
rect 1050 1718 1051 1722
rect 2101 1718 2102 1722
rect 2170 1718 2171 1722
rect 2266 1718 2267 1722
rect 2613 1718 2614 1722
rect 1056 1703 1058 1707
rect 1062 1703 1065 1707
rect 1069 1703 1072 1707
rect 2080 1703 2082 1707
rect 2086 1703 2089 1707
rect 2093 1703 2096 1707
rect 1989 1688 1990 1692
rect 246 1678 257 1681
rect 1142 1678 1153 1681
rect 1365 1678 1366 1682
rect 246 1677 250 1678
rect 1142 1677 1146 1678
rect 94 1671 98 1674
rect 94 1668 105 1671
rect 122 1668 129 1671
rect 1022 1668 1046 1671
rect 1170 1668 1177 1671
rect 1278 1668 1286 1671
rect 1326 1668 1345 1671
rect 1438 1668 1457 1671
rect 1510 1668 1526 1671
rect 1838 1671 1841 1681
rect 2150 1672 2153 1681
rect 1838 1668 1857 1671
rect 110 1658 129 1661
rect 190 1658 206 1661
rect 262 1658 281 1661
rect 310 1658 318 1661
rect 326 1658 345 1661
rect 526 1658 534 1661
rect 602 1658 609 1661
rect 654 1658 673 1661
rect 686 1658 694 1661
rect 870 1661 873 1668
rect 870 1658 881 1661
rect 1150 1661 1153 1668
rect 1142 1658 1153 1661
rect 1158 1658 1177 1661
rect 1342 1661 1345 1668
rect 1342 1658 1353 1661
rect 1566 1658 1582 1661
rect 1670 1658 1678 1661
rect 1934 1661 1937 1671
rect 1970 1668 1977 1671
rect 2170 1668 2177 1671
rect 2414 1671 2417 1681
rect 2398 1668 2417 1671
rect 1918 1658 1937 1661
rect 1962 1658 1969 1661
rect 2158 1658 2177 1661
rect 2314 1658 2321 1661
rect 2502 1658 2510 1661
rect 126 1648 129 1658
rect 342 1648 345 1658
rect 386 1648 390 1652
rect 670 1648 673 1658
rect 1142 1657 1146 1658
rect 2006 1648 2009 1658
rect 2638 1638 2646 1641
rect 1658 1628 1659 1632
rect 2021 1618 2022 1622
rect 544 1603 546 1607
rect 550 1603 553 1607
rect 557 1603 560 1607
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1573 1603 1576 1607
rect 1018 1588 1019 1592
rect 1762 1588 1763 1592
rect 2266 1588 2267 1592
rect 94 1568 102 1571
rect 877 1568 878 1572
rect 1274 1568 1275 1572
rect 2414 1568 2426 1571
rect 2422 1566 2426 1568
rect 438 1541 441 1551
rect 510 1548 529 1551
rect 750 1548 761 1551
rect 822 1551 825 1561
rect 806 1548 825 1551
rect 1030 1548 1046 1551
rect 1086 1551 1089 1561
rect 1054 1548 1089 1551
rect 1198 1548 1206 1551
rect 1286 1551 1289 1561
rect 1286 1548 1305 1551
rect 1470 1551 1473 1561
rect 1646 1558 1665 1561
rect 1982 1558 2001 1561
rect 1454 1548 1473 1551
rect 1486 1548 1494 1551
rect 1498 1548 1513 1551
rect 750 1542 753 1548
rect 438 1538 457 1541
rect 798 1538 801 1548
rect 1666 1548 1673 1551
rect 1678 1548 1686 1551
rect 1042 1538 1049 1541
rect 1074 1538 1089 1541
rect 1466 1538 1473 1541
rect 1686 1538 1694 1541
rect 1710 1541 1713 1551
rect 1942 1548 1950 1551
rect 2018 1548 2025 1551
rect 2050 1548 2057 1551
rect 2182 1548 2190 1551
rect 2470 1551 2473 1561
rect 2422 1548 2433 1551
rect 2454 1548 2473 1551
rect 2526 1551 2529 1561
rect 2510 1548 2529 1551
rect 2602 1548 2617 1551
rect 2422 1542 2425 1548
rect 1710 1538 1726 1541
rect 398 1528 417 1531
rect 2170 1528 2171 1532
rect 114 1518 115 1522
rect 1130 1518 1131 1522
rect 1056 1503 1058 1507
rect 1062 1503 1065 1507
rect 1069 1503 1072 1507
rect 2080 1503 2082 1507
rect 2086 1503 2089 1507
rect 2093 1503 2096 1507
rect 330 1488 331 1492
rect 986 1488 988 1492
rect 1558 1488 1574 1491
rect 126 1468 134 1471
rect 602 1468 609 1471
rect 654 1462 657 1471
rect 874 1468 881 1471
rect 1322 1468 1329 1471
rect 1358 1471 1361 1481
rect 1354 1468 1361 1471
rect 2446 1468 2454 1471
rect 2630 1468 2646 1471
rect 158 1458 177 1461
rect 342 1458 361 1461
rect 630 1458 649 1461
rect 694 1458 702 1461
rect 862 1458 881 1461
rect 910 1458 918 1461
rect 926 1458 945 1461
rect 1274 1458 1281 1461
rect 1342 1458 1350 1461
rect 1806 1458 1825 1461
rect 2278 1458 2297 1461
rect 2446 1458 2465 1461
rect 146 1448 150 1452
rect 158 1448 161 1458
rect 630 1448 633 1458
rect 1006 1448 1014 1451
rect 1438 1448 1446 1451
rect 1558 1448 1582 1451
rect 2038 1448 2041 1458
rect 2294 1448 2297 1458
rect 2446 1448 2449 1458
rect 1494 1446 1498 1448
rect 2494 1442 2498 1444
rect 1422 1438 1430 1441
rect 1434 1438 1465 1441
rect 2522 1438 2525 1442
rect 1022 1428 1025 1438
rect 682 1418 683 1422
rect 957 1418 958 1422
rect 544 1403 546 1407
rect 550 1403 553 1407
rect 557 1403 560 1407
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1573 1403 1576 1407
rect 2630 1388 2638 1391
rect 334 1368 342 1371
rect 570 1358 574 1362
rect 126 1342 129 1351
rect 162 1348 169 1351
rect 210 1348 217 1351
rect 758 1348 766 1351
rect 806 1348 814 1351
rect 874 1348 881 1351
rect 1230 1351 1233 1361
rect 1422 1358 1430 1361
rect 1230 1348 1249 1351
rect 1526 1351 1529 1361
rect 1586 1358 1593 1361
rect 1510 1348 1529 1351
rect 1638 1351 1641 1358
rect 1610 1348 1625 1351
rect 1630 1348 1641 1351
rect 1814 1348 1833 1351
rect 2038 1348 2046 1351
rect 1506 1338 1513 1341
rect 2130 1338 2145 1341
rect 2214 1341 2217 1351
rect 2582 1348 2590 1351
rect 2606 1342 2609 1351
rect 2202 1338 2217 1341
rect 2594 1338 2601 1341
rect 94 1331 98 1333
rect 94 1328 105 1331
rect 110 1328 129 1331
rect 229 1328 230 1332
rect 309 1328 310 1332
rect 350 1331 354 1333
rect 598 1332 602 1334
rect 342 1328 354 1331
rect 1478 1331 1481 1338
rect 1478 1328 1489 1331
rect 1494 1328 1502 1331
rect 1981 1328 1982 1332
rect 2218 1328 2225 1331
rect 2582 1331 2585 1338
rect 2582 1328 2593 1331
rect 181 1318 182 1322
rect 1042 1318 1043 1322
rect 1082 1318 1083 1322
rect 1389 1318 1390 1322
rect 1437 1318 1438 1322
rect 1597 1318 1598 1322
rect 2058 1318 2059 1322
rect 1056 1303 1058 1307
rect 1062 1303 1065 1307
rect 1069 1303 1072 1307
rect 2080 1303 2082 1307
rect 2086 1303 2089 1307
rect 2093 1303 2096 1307
rect 253 1288 254 1292
rect 858 1288 859 1292
rect 2274 1288 2275 1292
rect 2634 1288 2641 1291
rect 541 1278 542 1282
rect 626 1278 627 1282
rect 166 1271 170 1274
rect 74 1268 82 1271
rect 166 1268 177 1271
rect 194 1268 201 1271
rect 1590 1268 1601 1271
rect 1674 1268 1681 1271
rect 1702 1268 1710 1271
rect 1790 1268 1798 1271
rect 2126 1268 2134 1271
rect 2470 1268 2478 1271
rect 2502 1271 2506 1274
rect 2494 1268 2506 1271
rect 182 1258 201 1261
rect 234 1258 241 1261
rect 310 1258 318 1261
rect 398 1258 417 1261
rect 426 1258 433 1261
rect 462 1258 470 1261
rect 510 1258 518 1261
rect 902 1258 922 1261
rect 1198 1258 1201 1268
rect 1646 1262 1650 1264
rect 1438 1258 1457 1261
rect 1658 1258 1665 1261
rect 1674 1258 1681 1261
rect 1738 1258 1745 1261
rect 1794 1258 1801 1261
rect 2126 1258 2145 1261
rect 2298 1258 2313 1261
rect 2470 1258 2489 1261
rect 2534 1258 2542 1261
rect 198 1248 201 1258
rect 398 1248 401 1258
rect 918 1257 922 1258
rect 570 1248 582 1251
rect 814 1248 833 1251
rect 1050 1248 1057 1251
rect 1062 1248 1078 1251
rect 1202 1248 1209 1251
rect 1438 1248 1441 1258
rect 1614 1248 1625 1251
rect 2470 1248 2473 1258
rect 2614 1238 2630 1241
rect 1094 1228 1097 1238
rect 802 1218 803 1222
rect 890 1218 891 1222
rect 2058 1218 2059 1222
rect 544 1203 546 1207
rect 550 1203 553 1207
rect 557 1203 560 1207
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1573 1203 1576 1207
rect 770 1188 771 1192
rect 858 1188 859 1192
rect 1530 1188 1531 1192
rect 186 1168 187 1172
rect 1227 1168 1230 1172
rect 2278 1168 2286 1171
rect 110 1148 118 1151
rect 198 1151 201 1161
rect 718 1158 737 1161
rect 198 1148 217 1151
rect 262 1148 270 1151
rect 326 1148 334 1151
rect 398 1148 417 1151
rect 630 1148 646 1151
rect 870 1151 873 1161
rect 870 1148 889 1151
rect 1094 1148 1110 1151
rect 1270 1148 1286 1151
rect 1310 1151 1313 1161
rect 1310 1148 1329 1151
rect 1478 1148 1486 1151
rect 1598 1151 1601 1161
rect 1542 1148 1553 1151
rect 1566 1148 1601 1151
rect 1682 1148 1689 1151
rect 302 1138 321 1141
rect 398 1138 406 1141
rect 1038 1138 1066 1141
rect 1310 1138 1318 1141
rect 1550 1141 1553 1148
rect 2006 1148 2014 1151
rect 2114 1148 2121 1151
rect 2310 1151 2313 1161
rect 2294 1148 2313 1151
rect 2422 1142 2425 1151
rect 1550 1138 1558 1141
rect 1794 1138 1801 1141
rect 2106 1138 2113 1141
rect 2306 1138 2313 1141
rect 302 1128 305 1138
rect 430 1131 434 1133
rect 422 1128 434 1131
rect 550 1128 585 1131
rect 2142 1128 2161 1131
rect 2414 1128 2422 1131
rect 1056 1103 1058 1107
rect 1062 1103 1065 1107
rect 1069 1103 1072 1107
rect 2080 1103 2082 1107
rect 2086 1103 2089 1107
rect 2093 1103 2096 1107
rect 2058 1088 2059 1092
rect 2314 1088 2315 1092
rect 166 1078 185 1081
rect 854 1078 873 1081
rect 326 1068 334 1071
rect 554 1068 577 1071
rect 718 1068 726 1071
rect 1002 1068 1009 1071
rect 1054 1071 1057 1081
rect 1066 1078 1081 1081
rect 1430 1072 1433 1081
rect 1478 1078 1486 1081
rect 1886 1078 1905 1081
rect 1910 1078 1922 1081
rect 2106 1078 2113 1081
rect 1918 1077 1922 1078
rect 1054 1068 1089 1071
rect 1374 1068 1382 1071
rect 1422 1068 1430 1071
rect 1854 1068 1865 1071
rect 2254 1071 2257 1078
rect 2326 1077 2330 1078
rect 2606 1072 2610 1074
rect 2246 1068 2257 1071
rect 230 1058 246 1061
rect 326 1058 342 1061
rect 350 1058 369 1061
rect 718 1058 737 1061
rect 1134 1058 1153 1061
rect 1506 1058 1513 1061
rect 1546 1058 1553 1061
rect 1582 1058 1590 1061
rect 1862 1062 1865 1068
rect 1814 1058 1833 1061
rect 1886 1058 1889 1068
rect 2126 1058 2129 1068
rect 2178 1058 2193 1061
rect 2622 1061 2625 1068
rect 2622 1058 2633 1061
rect 2638 1058 2646 1061
rect 718 1048 721 1058
rect 1830 1048 1833 1058
rect 2062 1048 2065 1058
rect 2122 1018 2123 1022
rect 544 1003 546 1007
rect 550 1003 553 1007
rect 557 1003 560 1007
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1573 1003 1576 1007
rect 429 988 430 992
rect 1549 988 1550 992
rect 318 968 326 971
rect 674 968 677 972
rect 2646 971 2649 978
rect 2638 968 2649 971
rect 2190 966 2194 968
rect 2614 966 2618 968
rect 38 948 54 951
rect 126 951 129 961
rect 110 948 129 951
rect 190 948 201 951
rect 350 951 353 961
rect 334 948 353 951
rect 398 948 406 951
rect 478 951 481 961
rect 634 958 638 962
rect 478 948 497 951
rect 854 948 865 951
rect 950 948 969 951
rect 1090 948 1097 951
rect 1126 948 1145 951
rect 198 942 201 948
rect 94 938 105 941
rect 202 938 209 941
rect 374 938 382 941
rect 478 938 486 941
rect 502 938 518 941
rect 862 941 865 948
rect 1274 948 1281 951
rect 1526 948 1537 951
rect 1566 948 1582 951
rect 1734 951 1737 961
rect 1718 948 1737 951
rect 2026 948 2033 951
rect 1526 942 1529 948
rect 862 938 881 941
rect 950 938 958 941
rect 1126 938 1134 941
rect 1578 938 1593 941
rect 1702 938 1713 941
rect 1730 938 1737 941
rect 1758 938 1766 941
rect 1866 938 1873 941
rect 1910 938 1913 948
rect 2350 948 2369 951
rect 2590 942 2593 951
rect 2514 938 2529 941
rect 94 936 98 938
rect 974 931 977 938
rect 1702 936 1706 938
rect 982 931 986 933
rect 1686 932 1690 936
rect 974 928 986 931
rect 1262 928 1273 931
rect 2398 931 2402 933
rect 2390 928 2402 931
rect 2582 928 2590 931
rect 218 918 219 922
rect 522 918 529 921
rect 842 918 843 922
rect 1922 918 1923 922
rect 2186 918 2187 922
rect 2610 918 2611 922
rect 1056 903 1058 907
rect 1062 903 1065 907
rect 1069 903 1072 907
rect 2080 903 2082 907
rect 2086 903 2089 907
rect 2093 903 2096 907
rect 821 888 822 892
rect 1677 888 1678 892
rect 94 878 102 881
rect 1050 878 1051 882
rect 1182 878 1190 881
rect 1342 878 1353 881
rect 94 877 98 878
rect 1182 877 1186 878
rect 1342 877 1346 878
rect 1350 872 1353 878
rect 122 868 129 871
rect 510 868 529 871
rect 578 868 585 871
rect 1210 868 1217 871
rect 1370 868 1377 871
rect 1614 871 1617 878
rect 1614 868 1625 871
rect 110 858 129 861
rect 326 858 334 861
rect 426 858 433 861
rect 510 861 513 868
rect 502 858 513 861
rect 558 858 566 861
rect 802 858 809 861
rect 1198 858 1217 861
rect 1358 858 1377 861
rect 1406 858 1414 861
rect 1650 858 1665 861
rect 1734 858 1750 861
rect 1814 858 1822 861
rect 1862 861 1865 871
rect 1850 858 1865 861
rect 2058 858 2074 861
rect 710 848 729 851
rect 922 848 929 851
rect 1790 851 1794 854
rect 1610 848 1625 851
rect 1790 848 1801 851
rect 1813 838 1814 842
rect 2133 838 2134 842
rect 2379 838 2382 842
rect 2229 818 2230 822
rect 544 803 546 807
rect 550 803 553 807
rect 557 803 560 807
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1573 803 1576 807
rect 1653 788 1654 792
rect 1981 788 1982 792
rect 2101 778 2102 782
rect 94 768 102 771
rect 1282 768 1289 771
rect 2317 768 2318 772
rect 126 751 129 761
rect 894 761 897 768
rect 110 748 129 751
rect 342 748 358 751
rect 438 748 457 751
rect 702 751 705 761
rect 894 758 905 761
rect 954 758 961 761
rect 686 748 705 751
rect 766 748 785 751
rect 998 748 1006 751
rect 1062 751 1065 761
rect 1062 748 1097 751
rect 942 746 946 748
rect 1274 748 1281 751
rect 1502 748 1510 751
rect 1674 748 1681 751
rect 1766 751 1770 753
rect 1750 748 1770 751
rect 122 738 129 741
rect 262 738 281 741
rect 438 738 446 741
rect 558 738 574 741
rect 766 738 774 741
rect 1022 738 1038 741
rect 1278 738 1281 748
rect 1922 748 1929 751
rect 2150 748 2158 751
rect 2218 748 2225 751
rect 2254 748 2270 751
rect 2386 748 2393 751
rect 1602 738 1609 741
rect 2454 742 2457 751
rect 2506 748 2521 751
rect 2266 738 2273 741
rect 278 728 281 738
rect 1782 733 1786 738
rect 470 731 474 733
rect 466 728 474 731
rect 798 731 802 733
rect 790 728 802 731
rect 1390 731 1394 733
rect 1390 728 1401 731
rect 1870 728 1889 731
rect 1738 718 1739 722
rect 1056 703 1058 707
rect 1062 703 1065 707
rect 1069 703 1072 707
rect 2080 703 2082 707
rect 2086 703 2089 707
rect 2093 703 2096 707
rect 533 688 534 692
rect 586 688 587 692
rect 970 688 971 692
rect 1306 688 1307 692
rect 1658 688 1659 692
rect 270 678 289 681
rect 914 678 915 682
rect 1578 678 1590 681
rect 2042 678 2046 682
rect 2162 678 2166 682
rect 2258 678 2259 682
rect 2346 678 2362 681
rect 2450 678 2451 682
rect 2358 674 2362 678
rect 534 668 542 671
rect 606 668 625 671
rect 694 668 702 671
rect 742 668 761 671
rect 954 668 969 671
rect 990 668 1009 671
rect 1094 668 1110 671
rect 1166 668 1174 671
rect 1214 668 1222 671
rect 1298 668 1305 671
rect 1326 668 1345 671
rect 1518 668 1529 671
rect 1598 668 1606 671
rect 1854 668 1873 671
rect 1990 668 2006 671
rect 2022 668 2030 671
rect 2074 668 2097 671
rect 2142 668 2150 671
rect 2182 668 2201 671
rect 2386 668 2393 671
rect 182 658 198 661
rect 298 658 313 661
rect 382 658 401 661
rect 606 661 609 668
rect 598 658 609 661
rect 758 658 761 668
rect 926 658 945 661
rect 990 658 993 668
rect 1094 658 1102 661
rect 1326 658 1329 668
rect 1518 662 1521 668
rect 1602 658 1609 661
rect 1814 658 1833 661
rect 2062 658 2078 661
rect 2182 658 2185 668
rect 2194 658 2201 661
rect 2230 658 2238 661
rect 2270 658 2278 661
rect 2338 658 2345 661
rect 2374 658 2393 661
rect 2610 658 2617 661
rect 1830 648 1833 658
rect 2374 657 2378 658
rect 2538 648 2542 652
rect 437 638 438 642
rect 485 638 486 642
rect 325 628 326 632
rect 544 603 546 607
rect 550 603 553 607
rect 557 603 560 607
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1573 603 1576 607
rect 661 588 662 592
rect 1365 588 1366 592
rect 1458 588 1459 592
rect 2274 588 2275 592
rect 2618 588 2619 592
rect 2586 568 2593 571
rect 710 558 729 561
rect 862 558 881 561
rect 326 548 345 551
rect 366 548 385 551
rect 454 548 462 551
rect 502 548 510 551
rect 578 548 585 551
rect 642 548 649 551
rect 606 538 625 541
rect 718 538 721 548
rect 842 548 849 551
rect 974 548 982 551
rect 1098 548 1113 551
rect 1222 548 1230 551
rect 1310 551 1313 561
rect 1294 548 1313 551
rect 1434 548 1441 551
rect 1622 551 1625 561
rect 1622 548 1641 551
rect 1654 548 1665 551
rect 1706 548 1713 551
rect 1858 548 1865 551
rect 1934 548 1953 551
rect 2066 548 2073 551
rect 2078 548 2094 551
rect 1126 538 1134 541
rect 1278 538 1289 541
rect 1654 541 1657 548
rect 2210 548 2217 551
rect 2298 548 2305 551
rect 2334 548 2350 551
rect 2502 551 2505 561
rect 2502 548 2521 551
rect 2598 551 2601 558
rect 2598 548 2617 551
rect 1650 538 1657 541
rect 2058 538 2065 541
rect 2346 538 2353 541
rect 2578 538 2585 541
rect 314 528 315 532
rect 606 528 609 538
rect 1278 536 1282 538
rect 1142 528 1161 531
rect 1758 528 1777 531
rect 2322 528 2323 532
rect 1922 518 1923 522
rect 1056 503 1058 507
rect 1062 503 1065 507
rect 1069 503 1072 507
rect 2080 503 2082 507
rect 2086 503 2089 507
rect 2093 503 2096 507
rect 2274 488 2275 492
rect 94 478 102 481
rect 2026 478 2042 481
rect 94 477 98 478
rect 2038 474 2042 478
rect 2054 478 2065 481
rect 2070 478 2105 481
rect 2054 477 2058 478
rect 950 472 954 474
rect 122 468 129 471
rect 254 468 265 471
rect 282 468 289 471
rect 546 468 561 471
rect 958 471 962 474
rect 958 468 969 471
rect 1742 468 1750 471
rect 1774 471 1778 474
rect 1766 468 1778 471
rect 2326 468 2334 471
rect 2618 468 2625 471
rect 58 458 65 461
rect 110 458 129 461
rect 198 458 206 461
rect 262 462 265 468
rect 270 458 289 461
rect 526 458 561 461
rect 838 458 857 461
rect 974 458 993 461
rect 1006 458 1030 461
rect 1166 458 1174 461
rect 1414 458 1433 461
rect 1486 458 1505 461
rect 1526 458 1545 461
rect 1742 458 1761 461
rect 1902 458 1918 461
rect 2178 458 2185 461
rect 2326 458 2345 461
rect 2614 458 2633 461
rect 558 448 561 458
rect 826 448 830 452
rect 838 448 841 458
rect 990 448 993 458
rect 1414 448 1417 458
rect 1542 448 1545 458
rect 1554 448 1558 452
rect 1742 448 1745 458
rect 2182 448 2185 458
rect 2326 448 2329 458
rect 2614 452 2617 458
rect 75 438 78 442
rect 2602 438 2609 441
rect 1402 428 1403 432
rect 1474 418 1475 422
rect 2634 418 2635 422
rect 544 403 546 407
rect 550 403 553 407
rect 557 403 560 407
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1573 403 1576 407
rect 909 388 910 392
rect 2013 388 2014 392
rect 2133 388 2134 392
rect 2181 388 2182 392
rect 2282 388 2283 392
rect 1851 368 1854 372
rect 2349 368 2350 372
rect 2514 368 2521 371
rect 94 348 110 351
rect 262 348 270 351
rect 294 351 297 361
rect 294 348 313 351
rect 350 351 353 361
rect 350 348 369 351
rect 426 348 433 351
rect 542 351 546 353
rect 506 348 513 351
rect 542 348 577 351
rect 682 348 694 351
rect 710 351 713 361
rect 710 348 729 351
rect 890 348 897 351
rect 966 348 974 351
rect 1038 348 1073 351
rect 1366 348 1382 351
rect 1710 348 1718 351
rect 1910 348 1929 351
rect 1994 348 2001 351
rect 2162 348 2169 351
rect 2334 351 2337 361
rect 2294 348 2305 351
rect 2318 348 2337 351
rect 2418 348 2425 351
rect 2486 351 2489 361
rect 2486 348 2505 351
rect 2618 348 2625 351
rect 22 338 30 341
rect 226 338 233 341
rect 710 338 718 341
rect 1058 338 1073 341
rect 2302 341 2305 348
rect 2230 338 2249 341
rect 2302 338 2310 341
rect 2486 338 2494 341
rect 30 328 49 331
rect 1022 331 1026 333
rect 1030 331 1033 338
rect 1022 328 1033 331
rect 1390 328 1409 331
rect 1734 328 1753 331
rect 1934 328 1937 338
rect 2062 328 2081 331
rect 2086 328 2094 331
rect 2230 328 2233 338
rect 589 318 590 322
rect 1056 303 1058 307
rect 1062 303 1065 307
rect 1069 303 1072 307
rect 2080 303 2082 307
rect 2086 303 2089 307
rect 2093 303 2096 307
rect 245 288 246 292
rect 582 288 598 291
rect 954 288 955 292
rect 1082 288 1089 291
rect 2194 288 2195 292
rect 2506 288 2507 292
rect 870 272 873 281
rect 1290 278 1298 281
rect 1294 277 1298 278
rect 206 268 225 271
rect 478 268 486 271
rect 658 268 673 271
rect 222 261 225 268
rect 222 258 233 261
rect 718 262 721 271
rect 890 268 897 271
rect 1038 268 1046 271
rect 1062 268 1078 271
rect 1262 268 1270 271
rect 1534 268 1550 271
rect 1710 271 1714 274
rect 1702 268 1714 271
rect 2450 268 2457 271
rect 694 258 713 261
rect 878 258 897 261
rect 966 258 982 261
rect 1038 258 1057 261
rect 1262 258 1281 261
rect 1510 258 1529 261
rect 1678 258 1697 261
rect 1762 258 1769 261
rect 1870 258 1889 261
rect 2022 258 2041 261
rect 2266 258 2281 261
rect 2438 258 2457 261
rect 2518 258 2526 261
rect 618 248 622 252
rect 694 248 697 258
rect 1038 248 1041 258
rect 1510 248 1513 258
rect 1678 248 1681 258
rect 2022 248 2025 258
rect 2454 248 2457 258
rect 1410 238 1413 242
rect 1666 238 1667 242
rect 682 218 683 222
rect 544 203 546 207
rect 550 203 553 207
rect 557 203 560 207
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1573 203 1576 207
rect 754 188 755 192
rect 1165 188 1166 192
rect 1213 188 1214 192
rect 2570 168 2573 172
rect 158 151 161 161
rect 158 148 177 151
rect 238 151 242 153
rect 222 148 242 151
rect 126 138 134 141
rect 182 138 185 148
rect 606 151 609 161
rect 606 148 625 151
rect 886 148 905 151
rect 1110 142 1113 151
rect 1138 148 1153 151
rect 1622 148 1641 151
rect 1766 151 1769 161
rect 1766 148 1785 151
rect 1798 148 1809 151
rect 1798 142 1801 148
rect 2094 151 2097 161
rect 2106 158 2110 162
rect 2050 148 2057 151
rect 2062 148 2097 151
rect 2310 148 2318 151
rect 2510 148 2518 151
rect 606 138 614 141
rect 1766 138 1774 141
rect 1790 138 1798 141
rect 1958 138 1966 141
rect 2246 141 2249 148
rect 2238 138 2249 141
rect 342 128 361 131
rect 1110 128 1129 131
rect 1610 128 1611 132
rect 2266 118 2267 122
rect 1056 103 1058 107
rect 1062 103 1065 107
rect 1069 103 1072 107
rect 2080 103 2082 107
rect 2086 103 2089 107
rect 2093 103 2096 107
rect 90 88 91 92
rect 1054 88 1065 91
rect 1062 81 1065 88
rect 1062 78 1078 81
rect 1654 78 1665 81
rect 1822 78 1834 81
rect 1654 77 1658 78
rect 1830 77 1834 78
rect 314 68 321 71
rect 558 68 585 71
rect 686 68 694 71
rect 930 68 937 71
rect 1166 68 1174 71
rect 1198 71 1202 74
rect 1190 68 1202 71
rect 1798 68 1806 71
rect 558 62 561 68
rect 134 58 150 61
rect 302 58 321 61
rect 686 58 705 61
rect 918 58 937 61
rect 998 58 1014 61
rect 1086 58 1105 61
rect 1166 58 1185 61
rect 1302 58 1321 61
rect 1394 58 1409 61
rect 1598 58 1614 61
rect 1670 58 1689 61
rect 1730 58 1737 61
rect 1798 58 1817 61
rect 2158 58 2177 61
rect 318 48 321 58
rect 934 48 937 58
rect 1166 48 1169 58
rect 1318 48 1321 58
rect 2158 48 2161 58
rect 544 3 546 7
rect 550 3 553 7
rect 557 3 560 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1573 3 1576 7
<< m2contact >>
rect 546 2403 550 2407
rect 553 2403 557 2407
rect 1562 2403 1566 2407
rect 1569 2403 1573 2407
rect 278 2368 282 2372
rect 1382 2368 1386 2372
rect 1750 2368 1754 2372
rect 1950 2368 1954 2372
rect 2438 2368 2442 2372
rect 470 2348 474 2352
rect 622 2348 626 2352
rect 654 2358 658 2362
rect 1030 2358 1034 2362
rect 1078 2358 1082 2362
rect 1094 2358 1098 2362
rect 1126 2358 1130 2362
rect 710 2348 714 2352
rect 806 2348 810 2352
rect 830 2348 834 2352
rect 918 2348 922 2352
rect 926 2348 930 2352
rect 974 2348 978 2352
rect 1030 2348 1034 2352
rect 1078 2348 1082 2352
rect 1110 2348 1114 2352
rect 1182 2348 1186 2352
rect 1238 2348 1242 2352
rect 1246 2348 1250 2352
rect 1262 2358 1266 2362
rect 1398 2358 1402 2362
rect 1318 2348 1322 2352
rect 1462 2358 1466 2362
rect 1606 2358 1610 2362
rect 1822 2358 1826 2362
rect 1422 2348 1426 2352
rect 1486 2348 1490 2352
rect 1526 2348 1530 2352
rect 1534 2348 1538 2352
rect 1638 2348 1642 2352
rect 1646 2348 1650 2352
rect 1686 2347 1690 2351
rect 1758 2348 1762 2352
rect 1766 2348 1770 2352
rect 1846 2358 1850 2362
rect 1846 2348 1850 2352
rect 6 2338 10 2342
rect 78 2338 82 2342
rect 214 2338 218 2342
rect 222 2338 226 2342
rect 294 2338 298 2342
rect 358 2338 362 2342
rect 366 2338 370 2342
rect 446 2338 450 2342
rect 494 2338 498 2342
rect 534 2338 538 2342
rect 622 2338 626 2342
rect 646 2338 650 2342
rect 670 2338 674 2342
rect 686 2338 690 2342
rect 886 2338 890 2342
rect 974 2338 978 2342
rect 1078 2338 1082 2342
rect 1094 2338 1098 2342
rect 1102 2338 1106 2342
rect 1118 2338 1122 2342
rect 1230 2338 1234 2342
rect 1278 2338 1282 2342
rect 1294 2338 1298 2342
rect 1382 2338 1386 2342
rect 1398 2338 1402 2342
rect 1430 2338 1434 2342
rect 1446 2338 1450 2342
rect 1622 2338 1626 2342
rect 1654 2338 1658 2342
rect 1886 2347 1890 2351
rect 1998 2348 2002 2352
rect 2062 2348 2066 2352
rect 2222 2348 2226 2352
rect 2246 2358 2250 2362
rect 2534 2358 2538 2362
rect 2382 2348 2386 2352
rect 2486 2348 2490 2352
rect 1806 2338 1810 2342
rect 1854 2338 1858 2342
rect 1870 2338 1874 2342
rect 2038 2338 2042 2342
rect 2134 2338 2138 2342
rect 2142 2338 2146 2342
rect 2206 2338 2210 2342
rect 2214 2338 2218 2342
rect 2262 2338 2266 2342
rect 2270 2338 2274 2342
rect 2334 2338 2338 2342
rect 2374 2338 2378 2342
rect 2518 2338 2522 2342
rect 2550 2338 2554 2342
rect 2558 2338 2562 2342
rect 606 2328 610 2332
rect 870 2328 874 2332
rect 1158 2328 1162 2332
rect 1470 2328 1474 2332
rect 1686 2328 1690 2332
rect 2502 2328 2506 2332
rect 62 2318 66 2322
rect 134 2318 138 2322
rect 158 2318 162 2322
rect 422 2318 426 2322
rect 526 2318 530 2322
rect 766 2318 770 2322
rect 1022 2318 1026 2322
rect 1222 2318 1226 2322
rect 1494 2318 1498 2322
rect 1774 2318 1778 2322
rect 1958 2318 1962 2322
rect 2238 2318 2242 2322
rect 2430 2318 2434 2322
rect 2534 2318 2538 2322
rect 2614 2318 2618 2322
rect 1058 2303 1062 2307
rect 1065 2303 1069 2307
rect 2082 2303 2086 2307
rect 2089 2303 2093 2307
rect 318 2288 322 2292
rect 630 2288 634 2292
rect 950 2288 954 2292
rect 1102 2288 1106 2292
rect 1134 2288 1138 2292
rect 1166 2288 1170 2292
rect 1422 2288 1426 2292
rect 1630 2288 1634 2292
rect 1982 2288 1986 2292
rect 2006 2288 2010 2292
rect 2262 2288 2266 2292
rect 2382 2288 2386 2292
rect 2438 2288 2442 2292
rect 2622 2288 2626 2292
rect 222 2278 226 2282
rect 254 2278 258 2282
rect 382 2278 386 2282
rect 478 2278 482 2282
rect 838 2278 842 2282
rect 1726 2278 1730 2282
rect 1950 2278 1954 2282
rect 2102 2278 2106 2282
rect 2150 2278 2154 2282
rect 6 2268 10 2272
rect 70 2268 74 2272
rect 86 2268 90 2272
rect 182 2268 186 2272
rect 190 2268 194 2272
rect 430 2268 434 2272
rect 486 2268 490 2272
rect 566 2268 570 2272
rect 638 2268 642 2272
rect 654 2268 658 2272
rect 686 2268 690 2272
rect 798 2268 802 2272
rect 870 2268 874 2272
rect 878 2268 882 2272
rect 894 2268 898 2272
rect 974 2268 978 2272
rect 1174 2268 1178 2272
rect 1358 2268 1362 2272
rect 1414 2268 1418 2272
rect 1486 2268 1490 2272
rect 1558 2268 1562 2272
rect 1686 2268 1690 2272
rect 1766 2268 1770 2272
rect 1782 2268 1786 2272
rect 1910 2268 1914 2272
rect 1934 2268 1938 2272
rect 1990 2268 1994 2272
rect 2086 2268 2090 2272
rect 2158 2268 2162 2272
rect 2206 2268 2210 2272
rect 2302 2268 2306 2272
rect 2358 2268 2362 2272
rect 2406 2268 2410 2272
rect 2414 2268 2418 2272
rect 2462 2268 2466 2272
rect 2534 2268 2538 2272
rect 2558 2268 2562 2272
rect 2566 2268 2570 2272
rect 126 2258 130 2262
rect 174 2258 178 2262
rect 206 2258 210 2262
rect 262 2258 266 2262
rect 326 2258 330 2262
rect 334 2258 338 2262
rect 382 2258 386 2262
rect 398 2258 402 2262
rect 422 2258 426 2262
rect 462 2258 466 2262
rect 510 2258 514 2262
rect 574 2258 578 2262
rect 646 2258 650 2262
rect 726 2258 730 2262
rect 734 2258 738 2262
rect 806 2259 810 2263
rect 854 2258 858 2262
rect 886 2258 890 2262
rect 1006 2258 1010 2262
rect 1078 2258 1082 2262
rect 1086 2258 1090 2262
rect 1110 2258 1114 2262
rect 1150 2258 1154 2262
rect 1222 2258 1226 2262
rect 1254 2258 1258 2262
rect 1262 2258 1266 2262
rect 1270 2258 1274 2262
rect 1278 2258 1282 2262
rect 1302 2258 1306 2262
rect 1318 2258 1322 2262
rect 1326 2258 1330 2262
rect 1366 2258 1370 2262
rect 1406 2258 1410 2262
rect 1478 2258 1482 2262
rect 1518 2258 1522 2262
rect 1526 2258 1530 2262
rect 1550 2258 1554 2262
rect 1590 2258 1594 2262
rect 1614 2258 1618 2262
rect 1622 2258 1626 2262
rect 1662 2258 1666 2262
rect 1694 2259 1698 2263
rect 1742 2258 1746 2262
rect 1750 2258 1754 2262
rect 1782 2258 1786 2262
rect 1790 2258 1794 2262
rect 1814 2258 1818 2262
rect 1822 2258 1826 2262
rect 1846 2258 1850 2262
rect 1902 2258 1906 2262
rect 1966 2258 1970 2262
rect 1998 2258 2002 2262
rect 2070 2259 2074 2263
rect 2134 2258 2138 2262
rect 2166 2258 2170 2262
rect 2214 2258 2218 2262
rect 2318 2258 2322 2262
rect 2342 2258 2346 2262
rect 2350 2258 2354 2262
rect 2366 2258 2370 2262
rect 2454 2258 2458 2262
rect 670 2248 674 2252
rect 1142 2248 1146 2252
rect 1382 2248 1386 2252
rect 1406 2248 1410 2252
rect 1830 2248 1834 2252
rect 2390 2248 2394 2252
rect 2430 2248 2434 2252
rect 2542 2248 2546 2252
rect 166 2238 170 2242
rect 302 2238 306 2242
rect 342 2238 346 2242
rect 1070 2238 1074 2242
rect 406 2218 410 2222
rect 470 2218 474 2222
rect 718 2218 722 2222
rect 742 2218 746 2222
rect 950 2218 954 2222
rect 1190 2218 1194 2222
rect 1238 2218 1242 2222
rect 1294 2218 1298 2222
rect 1342 2218 1346 2222
rect 1534 2218 1538 2222
rect 1838 2218 1842 2222
rect 2262 2218 2266 2222
rect 2278 2218 2282 2222
rect 2326 2218 2330 2222
rect 2478 2218 2482 2222
rect 2550 2218 2554 2222
rect 546 2203 550 2207
rect 553 2203 557 2207
rect 1562 2203 1566 2207
rect 1569 2203 1573 2207
rect 462 2188 466 2192
rect 1406 2188 1410 2192
rect 1846 2188 1850 2192
rect 1870 2188 1874 2192
rect 2238 2188 2242 2192
rect 2542 2188 2546 2192
rect 558 2168 562 2172
rect 702 2168 706 2172
rect 1678 2168 1682 2172
rect 2190 2168 2194 2172
rect 2374 2168 2378 2172
rect 366 2158 370 2162
rect 70 2147 74 2151
rect 118 2148 122 2152
rect 150 2148 154 2152
rect 198 2148 202 2152
rect 614 2158 618 2162
rect 318 2147 322 2151
rect 390 2148 394 2152
rect 430 2148 434 2152
rect 438 2148 442 2152
rect 446 2148 450 2152
rect 470 2148 474 2152
rect 534 2148 538 2152
rect 638 2148 642 2152
rect 662 2148 666 2152
rect 686 2158 690 2162
rect 1790 2158 1794 2162
rect 750 2148 754 2152
rect 766 2148 770 2152
rect 838 2148 842 2152
rect 862 2148 866 2152
rect 934 2148 938 2152
rect 1022 2148 1026 2152
rect 1078 2148 1082 2152
rect 1110 2147 1114 2151
rect 1174 2148 1178 2152
rect 1206 2148 1210 2152
rect 1270 2148 1274 2152
rect 1318 2148 1322 2152
rect 1342 2148 1346 2152
rect 1350 2148 1354 2152
rect 1382 2148 1386 2152
rect 1526 2148 1530 2152
rect 1550 2148 1554 2152
rect 1606 2148 1610 2152
rect 1830 2158 1834 2162
rect 1742 2147 1746 2151
rect 1814 2148 1818 2152
rect 1846 2148 1850 2152
rect 1942 2148 1946 2152
rect 1966 2158 1970 2162
rect 2030 2148 2034 2152
rect 2126 2147 2130 2151
rect 2150 2148 2154 2152
rect 2198 2148 2202 2152
rect 2254 2148 2258 2152
rect 2318 2148 2322 2152
rect 2414 2148 2418 2152
rect 2478 2147 2482 2151
rect 2582 2148 2586 2152
rect 62 2138 66 2142
rect 126 2138 130 2142
rect 142 2138 146 2142
rect 238 2138 242 2142
rect 302 2138 306 2142
rect 350 2138 354 2142
rect 374 2138 378 2142
rect 414 2138 418 2142
rect 494 2138 498 2142
rect 622 2138 626 2142
rect 646 2138 650 2142
rect 686 2138 690 2142
rect 702 2138 706 2142
rect 998 2138 1002 2142
rect 1014 2138 1018 2142
rect 1142 2138 1146 2142
rect 1182 2138 1186 2142
rect 1198 2138 1202 2142
rect 1294 2138 1298 2142
rect 1422 2138 1426 2142
rect 1486 2138 1490 2142
rect 1670 2138 1674 2142
rect 1718 2138 1722 2142
rect 1758 2138 1762 2142
rect 1774 2138 1778 2142
rect 1790 2138 1794 2142
rect 1822 2138 1826 2142
rect 1854 2138 1858 2142
rect 1926 2138 1930 2142
rect 1934 2138 1938 2142
rect 1958 2138 1962 2142
rect 1982 2138 1986 2142
rect 2038 2138 2042 2142
rect 2086 2138 2090 2142
rect 2342 2138 2346 2142
rect 102 2128 106 2132
rect 998 2128 1002 2132
rect 2438 2138 2442 2142
rect 2590 2138 2594 2142
rect 1158 2128 1162 2132
rect 2390 2128 2394 2132
rect 2526 2128 2530 2132
rect 6 2118 10 2122
rect 158 2118 162 2122
rect 254 2118 258 2122
rect 590 2118 594 2122
rect 806 2118 810 2122
rect 990 2118 994 2122
rect 1046 2118 1050 2122
rect 1150 2118 1154 2122
rect 1214 2118 1218 2122
rect 1326 2118 1330 2122
rect 1366 2118 1370 2122
rect 1494 2118 1498 2122
rect 1990 2118 1994 2122
rect 2214 2118 2218 2122
rect 2262 2118 2266 2122
rect 2358 2118 2362 2122
rect 2638 2118 2642 2122
rect 1058 2103 1062 2107
rect 1065 2103 1069 2107
rect 2082 2103 2086 2107
rect 2089 2103 2093 2107
rect 94 2088 98 2092
rect 198 2088 202 2092
rect 406 2088 410 2092
rect 782 2088 786 2092
rect 990 2088 994 2092
rect 1142 2088 1146 2092
rect 1222 2088 1226 2092
rect 1406 2088 1410 2092
rect 1550 2088 1554 2092
rect 1846 2088 1850 2092
rect 1966 2088 1970 2092
rect 2110 2088 2114 2092
rect 2166 2088 2170 2092
rect 2302 2088 2306 2092
rect 2614 2088 2618 2092
rect 166 2078 170 2082
rect 430 2078 434 2082
rect 470 2078 474 2082
rect 982 2078 986 2082
rect 1190 2078 1194 2082
rect 1718 2078 1722 2082
rect 1910 2078 1914 2082
rect 2054 2078 2058 2082
rect 2134 2078 2138 2082
rect 126 2068 130 2072
rect 134 2068 138 2072
rect 150 2068 154 2072
rect 326 2068 330 2072
rect 374 2068 378 2072
rect 526 2068 530 2072
rect 638 2068 642 2072
rect 654 2068 658 2072
rect 750 2068 754 2072
rect 790 2068 794 2072
rect 814 2068 818 2072
rect 902 2068 906 2072
rect 926 2068 930 2072
rect 1166 2068 1170 2072
rect 1302 2068 1306 2072
rect 1358 2068 1362 2072
rect 1414 2068 1418 2072
rect 1462 2068 1466 2072
rect 1502 2068 1506 2072
rect 1542 2068 1546 2072
rect 1574 2068 1578 2072
rect 1598 2068 1602 2072
rect 1630 2068 1634 2072
rect 1646 2068 1650 2072
rect 1830 2068 1834 2072
rect 1942 2068 1946 2072
rect 1998 2068 2002 2072
rect 2174 2068 2178 2072
rect 2182 2068 2186 2072
rect 2238 2068 2242 2072
rect 2294 2068 2298 2072
rect 2382 2068 2386 2072
rect 2438 2068 2442 2072
rect 2542 2068 2546 2072
rect 2558 2068 2562 2072
rect 46 2058 50 2062
rect 62 2058 66 2062
rect 110 2058 114 2062
rect 206 2058 210 2062
rect 214 2058 218 2062
rect 222 2058 226 2062
rect 254 2058 258 2062
rect 262 2058 266 2062
rect 278 2058 282 2062
rect 302 2058 306 2062
rect 310 2058 314 2062
rect 350 2058 354 2062
rect 414 2058 418 2062
rect 422 2058 426 2062
rect 478 2058 482 2062
rect 486 2058 490 2062
rect 518 2058 522 2062
rect 574 2058 578 2062
rect 598 2058 602 2062
rect 686 2058 690 2062
rect 694 2058 698 2062
rect 710 2058 714 2062
rect 734 2058 738 2062
rect 742 2058 746 2062
rect 766 2058 770 2062
rect 798 2058 802 2062
rect 846 2058 850 2062
rect 918 2058 922 2062
rect 934 2058 938 2062
rect 942 2058 946 2062
rect 966 2058 970 2062
rect 998 2058 1002 2062
rect 1014 2058 1018 2062
rect 1038 2058 1042 2062
rect 1046 2058 1050 2062
rect 1070 2058 1074 2062
rect 1078 2058 1082 2062
rect 1110 2058 1114 2062
rect 1118 2058 1122 2062
rect 1126 2058 1130 2062
rect 1150 2058 1154 2062
rect 1174 2058 1178 2062
rect 1278 2058 1282 2062
rect 1350 2058 1354 2062
rect 1422 2058 1426 2062
rect 1470 2058 1474 2062
rect 1478 2058 1482 2062
rect 1510 2058 1514 2062
rect 1542 2058 1546 2062
rect 1598 2058 1602 2062
rect 1606 2058 1610 2062
rect 1694 2058 1698 2062
rect 1710 2058 1714 2062
rect 1790 2058 1794 2062
rect 1902 2058 1906 2062
rect 1950 2058 1954 2062
rect 1990 2058 1994 2062
rect 2006 2058 2010 2062
rect 2014 2058 2018 2062
rect 2046 2058 2050 2062
rect 2118 2058 2122 2062
rect 2126 2058 2130 2062
rect 2150 2058 2154 2062
rect 2190 2058 2194 2062
rect 2198 2058 2202 2062
rect 2230 2058 2234 2062
rect 2246 2058 2250 2062
rect 2278 2058 2282 2062
rect 2286 2058 2290 2062
rect 2350 2058 2354 2062
rect 2398 2058 2402 2062
rect 2406 2058 2410 2062
rect 2518 2058 2522 2062
rect 102 2048 106 2052
rect 134 2048 138 2052
rect 902 2048 906 2052
rect 1198 2048 1202 2052
rect 1446 2048 1450 2052
rect 1534 2048 1538 2052
rect 1550 2048 1554 2052
rect 1630 2048 1634 2052
rect 1974 2048 1978 2052
rect 2262 2048 2266 2052
rect 1422 2038 1426 2042
rect 1646 2038 1650 2042
rect 238 2018 242 2022
rect 294 2018 298 2022
rect 494 2018 498 2022
rect 726 2018 730 2022
rect 894 2018 898 2022
rect 950 2018 954 2022
rect 1022 2018 1026 2022
rect 1086 2018 1090 2022
rect 1750 2018 1754 2022
rect 2022 2018 2026 2022
rect 2206 2018 2210 2022
rect 2462 2018 2466 2022
rect 546 2003 550 2007
rect 553 2003 557 2007
rect 1562 2003 1566 2007
rect 1569 2003 1573 2007
rect 862 1988 866 1992
rect 1534 1988 1538 1992
rect 1782 1988 1786 1992
rect 1846 1988 1850 1992
rect 2478 1988 2482 1992
rect 2622 1988 2626 1992
rect 1102 1968 1106 1972
rect 1414 1968 1418 1972
rect 1606 1968 1610 1972
rect 2318 1968 2322 1972
rect 2534 1968 2538 1972
rect 246 1958 250 1962
rect 6 1948 10 1952
rect 110 1948 114 1952
rect 190 1948 194 1952
rect 222 1948 226 1952
rect 270 1958 274 1962
rect 478 1958 482 1962
rect 678 1958 682 1962
rect 854 1958 858 1962
rect 958 1958 962 1962
rect 1198 1958 1202 1962
rect 270 1948 274 1952
rect 342 1948 346 1952
rect 414 1948 418 1952
rect 518 1948 522 1952
rect 574 1948 578 1952
rect 622 1948 626 1952
rect 638 1948 642 1952
rect 670 1948 674 1952
rect 686 1948 690 1952
rect 694 1948 698 1952
rect 766 1948 770 1952
rect 806 1948 810 1952
rect 814 1948 818 1952
rect 838 1948 842 1952
rect 878 1948 882 1952
rect 886 1948 890 1952
rect 998 1948 1002 1952
rect 1078 1948 1082 1952
rect 1270 1958 1274 1962
rect 1310 1958 1314 1962
rect 1574 1958 1578 1962
rect 1590 1958 1594 1962
rect 1822 1958 1826 1962
rect 1150 1947 1154 1951
rect 1214 1948 1218 1952
rect 1222 1948 1226 1952
rect 1262 1948 1266 1952
rect 1310 1948 1314 1952
rect 1350 1947 1354 1951
rect 1422 1948 1426 1952
rect 1430 1948 1434 1952
rect 1454 1948 1458 1952
rect 1502 1948 1506 1952
rect 1510 1948 1514 1952
rect 1518 1948 1522 1952
rect 1550 1948 1554 1952
rect 1582 1948 1586 1952
rect 1670 1948 1674 1952
rect 1734 1948 1738 1952
rect 1790 1948 1794 1952
rect 1798 1948 1802 1952
rect 2150 1958 2154 1962
rect 1846 1948 1850 1952
rect 1862 1948 1866 1952
rect 1870 1948 1874 1952
rect 1982 1948 1986 1952
rect 86 1938 90 1942
rect 198 1938 202 1942
rect 214 1938 218 1942
rect 230 1938 234 1942
rect 278 1938 282 1942
rect 366 1938 370 1942
rect 390 1938 394 1942
rect 486 1938 490 1942
rect 510 1938 514 1942
rect 582 1938 586 1942
rect 630 1938 634 1942
rect 702 1938 706 1942
rect 774 1938 778 1942
rect 870 1938 874 1942
rect 918 1938 922 1942
rect 1006 1938 1010 1942
rect 1142 1938 1146 1942
rect 1182 1938 1186 1942
rect 1230 1938 1234 1942
rect 1286 1938 1290 1942
rect 1318 1938 1322 1942
rect 1334 1938 1338 1942
rect 1358 1938 1362 1942
rect 2086 1947 2090 1951
rect 2174 1948 2178 1952
rect 2190 1948 2194 1952
rect 2198 1948 2202 1952
rect 2222 1948 2226 1952
rect 2238 1948 2242 1952
rect 2270 1948 2274 1952
rect 2302 1958 2306 1962
rect 2494 1958 2498 1962
rect 2646 1958 2650 1962
rect 2382 1948 2386 1952
rect 2422 1948 2426 1952
rect 2430 1948 2434 1952
rect 2454 1948 2458 1952
rect 2478 1948 2482 1952
rect 2494 1948 2498 1952
rect 2574 1948 2578 1952
rect 2622 1948 2626 1952
rect 1542 1938 1546 1942
rect 1574 1938 1578 1942
rect 1606 1938 1610 1942
rect 1694 1938 1698 1942
rect 1806 1938 1810 1942
rect 1854 1938 1858 1942
rect 1902 1938 1906 1942
rect 2006 1938 2010 1942
rect 2070 1938 2074 1942
rect 2118 1938 2122 1942
rect 2150 1938 2154 1942
rect 2182 1938 2186 1942
rect 2270 1938 2274 1942
rect 2302 1938 2306 1942
rect 2318 1938 2322 1942
rect 2406 1938 2410 1942
rect 2462 1938 2466 1942
rect 2470 1938 2474 1942
rect 2598 1938 2602 1942
rect 2614 1938 2618 1942
rect 150 1928 154 1932
rect 654 1928 658 1932
rect 1742 1928 1746 1932
rect 1918 1928 1922 1932
rect 2510 1928 2514 1932
rect 62 1918 66 1922
rect 286 1918 290 1922
rect 470 1918 474 1922
rect 526 1918 530 1922
rect 710 1918 714 1922
rect 830 1918 834 1922
rect 1046 1918 1050 1922
rect 1086 1918 1090 1922
rect 1486 1918 1490 1922
rect 1718 1918 1722 1922
rect 2022 1918 2026 1922
rect 2206 1918 2210 1922
rect 2254 1918 2258 1922
rect 1058 1903 1062 1907
rect 1065 1903 1069 1907
rect 2082 1903 2086 1907
rect 2089 1903 2093 1907
rect 254 1888 258 1892
rect 478 1888 482 1892
rect 670 1888 674 1892
rect 830 1888 834 1892
rect 1062 1888 1066 1892
rect 1374 1888 1378 1892
rect 1638 1888 1642 1892
rect 1870 1888 1874 1892
rect 2438 1888 2442 1892
rect 2614 1888 2618 1892
rect 142 1878 146 1882
rect 278 1878 282 1882
rect 318 1878 322 1882
rect 438 1878 442 1882
rect 734 1878 738 1882
rect 886 1878 890 1882
rect 1310 1878 1314 1882
rect 1462 1878 1466 1882
rect 1646 1878 1650 1882
rect 2006 1878 2010 1882
rect 102 1868 106 1872
rect 174 1868 178 1872
rect 470 1868 474 1872
rect 550 1868 554 1872
rect 654 1868 658 1872
rect 718 1868 722 1872
rect 1142 1868 1146 1872
rect 1158 1868 1162 1872
rect 1174 1868 1178 1872
rect 1206 1868 1210 1872
rect 1214 1868 1218 1872
rect 1382 1868 1386 1872
rect 1430 1868 1434 1872
rect 1518 1868 1522 1872
rect 1558 1868 1562 1872
rect 1662 1868 1666 1872
rect 2134 1868 2138 1872
rect 2222 1868 2226 1872
rect 2334 1868 2338 1872
rect 38 1858 42 1862
rect 62 1858 66 1862
rect 126 1858 130 1862
rect 150 1858 154 1862
rect 158 1858 162 1862
rect 198 1858 202 1862
rect 262 1858 266 1862
rect 270 1858 274 1862
rect 334 1858 338 1862
rect 358 1858 362 1862
rect 366 1858 370 1862
rect 382 1858 386 1862
rect 406 1858 410 1862
rect 414 1858 418 1862
rect 422 1858 426 1862
rect 430 1858 434 1862
rect 454 1858 458 1862
rect 494 1858 498 1862
rect 502 1858 506 1862
rect 526 1858 530 1862
rect 558 1858 562 1862
rect 566 1858 570 1862
rect 590 1858 594 1862
rect 606 1858 610 1862
rect 614 1858 618 1862
rect 630 1858 634 1862
rect 646 1858 650 1862
rect 678 1858 682 1862
rect 686 1858 690 1862
rect 766 1859 770 1863
rect 798 1858 802 1862
rect 838 1858 842 1862
rect 846 1858 850 1862
rect 870 1858 874 1862
rect 934 1858 938 1862
rect 942 1858 946 1862
rect 950 1858 954 1862
rect 982 1858 986 1862
rect 990 1858 994 1862
rect 1006 1858 1010 1862
rect 1030 1858 1034 1862
rect 1046 1858 1050 1862
rect 1094 1858 1098 1862
rect 1126 1859 1130 1863
rect 1198 1858 1202 1862
rect 1318 1858 1322 1862
rect 1390 1858 1394 1862
rect 1398 1858 1402 1862
rect 1470 1858 1474 1862
rect 1598 1858 1602 1862
rect 1694 1858 1698 1862
rect 1702 1858 1706 1862
rect 1710 1858 1714 1862
rect 1742 1858 1746 1862
rect 1750 1858 1754 1862
rect 1758 1858 1762 1862
rect 1766 1858 1770 1862
rect 1790 1858 1794 1862
rect 1798 1858 1802 1862
rect 1814 1858 1818 1862
rect 1838 1858 1842 1862
rect 1854 1858 1858 1862
rect 1886 1858 1890 1862
rect 1894 1858 1898 1862
rect 1918 1858 1922 1862
rect 2430 1868 2434 1872
rect 2518 1868 2522 1872
rect 2534 1868 2538 1872
rect 2598 1868 2602 1872
rect 2638 1868 2642 1872
rect 1966 1858 1970 1862
rect 1974 1858 1978 1862
rect 1990 1858 1994 1862
rect 2014 1858 2018 1862
rect 2022 1858 2026 1862
rect 2030 1858 2034 1862
rect 2038 1858 2042 1862
rect 2062 1858 2066 1862
rect 2094 1858 2098 1862
rect 2102 1858 2106 1862
rect 2126 1858 2130 1862
rect 2142 1858 2146 1862
rect 2150 1858 2154 1862
rect 2174 1858 2178 1862
rect 2238 1858 2242 1862
rect 2246 1858 2250 1862
rect 2294 1858 2298 1862
rect 2318 1858 2322 1862
rect 2334 1858 2338 1862
rect 2342 1858 2346 1862
rect 2366 1858 2370 1862
rect 2374 1858 2378 1862
rect 2382 1858 2386 1862
rect 2430 1858 2434 1862
rect 2494 1858 2498 1862
rect 486 1848 490 1852
rect 670 1848 674 1852
rect 1174 1848 1178 1852
rect 1414 1848 1418 1852
rect 2398 1848 2402 1852
rect 2422 1848 2426 1852
rect 2606 1848 2610 1852
rect 1622 1838 1626 1842
rect 110 1818 114 1822
rect 350 1818 354 1822
rect 398 1818 402 1822
rect 582 1818 586 1822
rect 862 1818 866 1822
rect 918 1818 922 1822
rect 974 1818 978 1822
rect 1014 1818 1018 1822
rect 1270 1818 1274 1822
rect 1526 1818 1530 1822
rect 1734 1818 1738 1822
rect 1782 1818 1786 1822
rect 1822 1818 1826 1822
rect 1958 1818 1962 1822
rect 2054 1818 2058 1822
rect 2166 1818 2170 1822
rect 2278 1818 2282 1822
rect 2302 1818 2306 1822
rect 2590 1818 2594 1822
rect 546 1803 550 1807
rect 553 1803 557 1807
rect 1562 1803 1566 1807
rect 1569 1803 1573 1807
rect 118 1788 122 1792
rect 854 1788 858 1792
rect 1518 1788 1522 1792
rect 1654 1788 1658 1792
rect 1814 1788 1818 1792
rect 2214 1788 2218 1792
rect 318 1778 322 1782
rect 526 1768 530 1772
rect 718 1768 722 1772
rect 1526 1768 1530 1772
rect 2070 1768 2074 1772
rect 2374 1768 2378 1772
rect 262 1758 266 1762
rect 342 1758 346 1762
rect 678 1758 682 1762
rect 70 1747 74 1751
rect 110 1748 114 1752
rect 134 1748 138 1752
rect 142 1748 146 1752
rect 150 1748 154 1752
rect 158 1748 162 1752
rect 190 1748 194 1752
rect 230 1748 234 1752
rect 238 1748 242 1752
rect 254 1748 258 1752
rect 278 1748 282 1752
rect 294 1748 298 1752
rect 302 1748 306 1752
rect 326 1748 330 1752
rect 334 1748 338 1752
rect 358 1748 362 1752
rect 398 1748 402 1752
rect 406 1748 410 1752
rect 438 1748 442 1752
rect 470 1748 474 1752
rect 478 1748 482 1752
rect 494 1748 498 1752
rect 534 1748 538 1752
rect 542 1748 546 1752
rect 558 1748 562 1752
rect 574 1748 578 1752
rect 622 1748 626 1752
rect 646 1748 650 1752
rect 654 1748 658 1752
rect 1062 1758 1066 1762
rect 1086 1758 1090 1762
rect 1134 1758 1138 1762
rect 1150 1758 1154 1762
rect 1838 1758 1842 1762
rect 1942 1758 1946 1762
rect 2094 1758 2098 1762
rect 702 1748 706 1752
rect 766 1748 770 1752
rect 814 1748 818 1752
rect 846 1748 850 1752
rect 886 1748 890 1752
rect 86 1738 90 1742
rect 366 1738 370 1742
rect 374 1738 378 1742
rect 398 1738 402 1742
rect 414 1738 418 1742
rect 430 1738 434 1742
rect 918 1747 922 1751
rect 950 1748 954 1752
rect 662 1738 666 1742
rect 694 1738 698 1742
rect 710 1738 714 1742
rect 798 1738 802 1742
rect 822 1738 826 1742
rect 846 1738 850 1742
rect 934 1738 938 1742
rect 958 1738 962 1742
rect 974 1738 978 1742
rect 998 1748 1002 1752
rect 1022 1748 1026 1752
rect 1030 1748 1034 1752
rect 1078 1748 1082 1752
rect 1110 1748 1114 1752
rect 1134 1748 1138 1752
rect 1174 1748 1178 1752
rect 1246 1747 1250 1751
rect 1294 1748 1298 1752
rect 1326 1748 1330 1752
rect 1366 1748 1370 1752
rect 1478 1748 1482 1752
rect 1486 1748 1490 1752
rect 1494 1748 1498 1752
rect 1598 1748 1602 1752
rect 1710 1748 1714 1752
rect 1718 1748 1722 1752
rect 1758 1748 1762 1752
rect 1854 1748 1858 1752
rect 1878 1748 1882 1752
rect 1918 1748 1922 1752
rect 1926 1748 1930 1752
rect 1950 1748 1954 1752
rect 1990 1747 1994 1751
rect 2110 1748 2114 1752
rect 2150 1748 2154 1752
rect 2198 1748 2202 1752
rect 2206 1748 2210 1752
rect 2230 1748 2234 1752
rect 2238 1748 2242 1752
rect 2246 1748 2250 1752
rect 2254 1748 2258 1752
rect 2278 1748 2282 1752
rect 2310 1758 2314 1762
rect 2326 1758 2330 1762
rect 2358 1758 2362 1762
rect 2478 1758 2482 1762
rect 2606 1758 2610 1762
rect 2310 1748 2314 1752
rect 2334 1748 2338 1752
rect 2342 1748 2346 1752
rect 2438 1748 2442 1752
rect 2486 1748 2490 1752
rect 2494 1748 2498 1752
rect 2566 1748 2570 1752
rect 1038 1738 1042 1742
rect 1054 1738 1058 1742
rect 1102 1738 1106 1742
rect 1118 1738 1122 1742
rect 1142 1738 1146 1742
rect 1166 1738 1170 1742
rect 1262 1738 1266 1742
rect 1302 1738 1306 1742
rect 1326 1738 1330 1742
rect 1342 1738 1346 1742
rect 1446 1738 1450 1742
rect 1502 1738 1506 1742
rect 1526 1738 1530 1742
rect 1542 1738 1546 1742
rect 1678 1738 1682 1742
rect 1902 1738 1906 1742
rect 1974 1738 1978 1742
rect 2110 1738 2114 1742
rect 2126 1738 2130 1742
rect 2142 1738 2146 1742
rect 2166 1738 2170 1742
rect 2182 1738 2186 1742
rect 2318 1738 2322 1742
rect 2350 1738 2354 1742
rect 2374 1738 2378 1742
rect 2502 1738 2506 1742
rect 2590 1738 2594 1742
rect 2638 1738 2642 1742
rect 222 1728 226 1732
rect 494 1728 498 1732
rect 1278 1728 1282 1732
rect 1390 1728 1394 1732
rect 1518 1728 1522 1732
rect 1590 1728 1594 1732
rect 1750 1728 1754 1732
rect 2070 1728 2074 1732
rect 2134 1728 2138 1732
rect 2446 1728 2450 1732
rect 6 1718 10 1722
rect 350 1718 354 1722
rect 390 1718 394 1722
rect 430 1718 434 1722
rect 454 1718 458 1722
rect 486 1718 490 1722
rect 590 1718 594 1722
rect 830 1718 834 1722
rect 966 1718 970 1722
rect 1046 1718 1050 1722
rect 1134 1718 1138 1722
rect 1182 1718 1186 1722
rect 1814 1718 1818 1722
rect 1822 1718 1826 1722
rect 2054 1718 2058 1722
rect 2102 1718 2106 1722
rect 2166 1718 2170 1722
rect 2262 1718 2266 1722
rect 2358 1718 2362 1722
rect 2510 1718 2514 1722
rect 2614 1718 2618 1722
rect 1058 1703 1062 1707
rect 1065 1703 1069 1707
rect 2082 1703 2086 1707
rect 2089 1703 2093 1707
rect 94 1688 98 1692
rect 246 1688 250 1692
rect 406 1688 410 1692
rect 550 1688 554 1692
rect 702 1688 706 1692
rect 854 1688 858 1692
rect 1478 1688 1482 1692
rect 1606 1688 1610 1692
rect 1710 1688 1714 1692
rect 1790 1688 1794 1692
rect 1830 1688 1834 1692
rect 1958 1688 1962 1692
rect 1990 1688 1994 1692
rect 2054 1688 2058 1692
rect 2462 1688 2466 1692
rect 2470 1688 2474 1692
rect 342 1678 346 1682
rect 502 1678 506 1682
rect 766 1678 770 1682
rect 1366 1678 1370 1682
rect 14 1668 18 1672
rect 118 1668 122 1672
rect 150 1668 154 1672
rect 166 1668 170 1672
rect 318 1668 322 1672
rect 366 1668 370 1672
rect 398 1668 402 1672
rect 486 1668 490 1672
rect 518 1668 522 1672
rect 646 1668 650 1672
rect 694 1668 698 1672
rect 798 1668 802 1672
rect 870 1668 874 1672
rect 966 1668 970 1672
rect 1046 1668 1050 1672
rect 1062 1668 1066 1672
rect 1150 1668 1154 1672
rect 1166 1668 1170 1672
rect 1230 1668 1234 1672
rect 1286 1668 1290 1672
rect 1398 1668 1402 1672
rect 1406 1668 1410 1672
rect 1414 1668 1418 1672
rect 1430 1668 1434 1672
rect 1494 1668 1498 1672
rect 1502 1668 1506 1672
rect 1526 1668 1530 1672
rect 1686 1668 1690 1672
rect 1822 1668 1826 1672
rect 1846 1678 1850 1682
rect 2406 1678 2410 1682
rect 1878 1668 1882 1672
rect 1894 1668 1898 1672
rect 1926 1668 1930 1672
rect 38 1658 42 1662
rect 142 1658 146 1662
rect 206 1658 210 1662
rect 302 1658 306 1662
rect 318 1658 322 1662
rect 358 1658 362 1662
rect 390 1658 394 1662
rect 462 1658 466 1662
rect 510 1658 514 1662
rect 534 1658 538 1662
rect 582 1658 586 1662
rect 598 1658 602 1662
rect 678 1658 682 1662
rect 694 1658 698 1662
rect 758 1658 762 1662
rect 902 1658 906 1662
rect 910 1658 914 1662
rect 926 1658 930 1662
rect 934 1658 938 1662
rect 950 1658 954 1662
rect 958 1658 962 1662
rect 990 1658 994 1662
rect 998 1658 1002 1662
rect 1022 1658 1026 1662
rect 1086 1658 1090 1662
rect 1198 1658 1202 1662
rect 1206 1658 1210 1662
rect 1214 1658 1218 1662
rect 1246 1658 1250 1662
rect 1254 1658 1258 1662
rect 1278 1658 1282 1662
rect 1294 1658 1298 1662
rect 1302 1658 1306 1662
rect 1326 1658 1330 1662
rect 1374 1658 1378 1662
rect 1382 1658 1386 1662
rect 1390 1658 1394 1662
rect 1422 1658 1426 1662
rect 1462 1658 1466 1662
rect 1486 1658 1490 1662
rect 1518 1658 1522 1662
rect 1534 1658 1538 1662
rect 1558 1658 1562 1662
rect 1582 1658 1586 1662
rect 1598 1658 1602 1662
rect 1622 1658 1626 1662
rect 1630 1658 1634 1662
rect 1638 1658 1642 1662
rect 1646 1658 1650 1662
rect 1678 1658 1682 1662
rect 1694 1658 1698 1662
rect 1718 1658 1722 1662
rect 1726 1658 1730 1662
rect 1750 1658 1754 1662
rect 1766 1658 1770 1662
rect 1774 1658 1778 1662
rect 1798 1658 1802 1662
rect 1814 1658 1818 1662
rect 1862 1658 1866 1662
rect 1870 1658 1874 1662
rect 1902 1658 1906 1662
rect 1966 1668 1970 1672
rect 1990 1668 1994 1672
rect 2030 1668 2034 1672
rect 2134 1668 2138 1672
rect 2150 1668 2154 1672
rect 2166 1668 2170 1672
rect 2318 1668 2322 1672
rect 2366 1668 2370 1672
rect 2382 1668 2386 1672
rect 2566 1678 2570 1682
rect 2430 1668 2434 1672
rect 2446 1668 2450 1672
rect 2526 1668 2530 1672
rect 2582 1668 2586 1672
rect 2614 1668 2618 1672
rect 1942 1658 1946 1662
rect 1958 1658 1962 1662
rect 1998 1658 2002 1662
rect 2006 1658 2010 1662
rect 2022 1658 2026 1662
rect 2118 1659 2122 1663
rect 2198 1658 2202 1662
rect 2206 1658 2210 1662
rect 2222 1658 2226 1662
rect 2246 1658 2250 1662
rect 2254 1658 2258 1662
rect 2270 1658 2274 1662
rect 2294 1658 2298 1662
rect 2302 1658 2306 1662
rect 2310 1658 2314 1662
rect 2342 1658 2346 1662
rect 2350 1658 2354 1662
rect 2374 1658 2378 1662
rect 2390 1658 2394 1662
rect 2422 1658 2426 1662
rect 2438 1658 2442 1662
rect 2510 1658 2514 1662
rect 2526 1658 2530 1662
rect 2590 1658 2594 1662
rect 2598 1658 2602 1662
rect 2622 1658 2626 1662
rect 118 1648 122 1652
rect 286 1648 290 1652
rect 334 1648 338 1652
rect 374 1648 378 1652
rect 390 1648 394 1652
rect 662 1648 666 1652
rect 886 1648 890 1652
rect 982 1648 986 1652
rect 1446 1648 1450 1652
rect 1478 1648 1482 1652
rect 1542 1648 1546 1652
rect 1710 1648 1714 1652
rect 1742 1648 1746 1652
rect 1894 1648 1898 1652
rect 1910 1648 1914 1652
rect 1958 1648 1962 1652
rect 2358 1648 2362 1652
rect 2462 1648 2466 1652
rect 2230 1638 2234 1642
rect 2646 1638 2650 1642
rect 974 1628 978 1632
rect 1654 1628 1658 1632
rect 2022 1618 2026 1622
rect 2054 1618 2058 1622
rect 2278 1618 2282 1622
rect 2566 1618 2570 1622
rect 546 1603 550 1607
rect 553 1603 557 1607
rect 1562 1603 1566 1607
rect 1569 1603 1573 1607
rect 766 1588 770 1592
rect 1014 1588 1018 1592
rect 1126 1588 1130 1592
rect 1430 1588 1434 1592
rect 1758 1588 1762 1592
rect 1798 1588 1802 1592
rect 1918 1588 1922 1592
rect 2214 1588 2218 1592
rect 2262 1588 2266 1592
rect 2414 1588 2418 1592
rect 1254 1578 1258 1582
rect 1542 1578 1546 1582
rect 102 1568 106 1572
rect 646 1568 650 1572
rect 742 1568 746 1572
rect 878 1568 882 1572
rect 990 1568 994 1572
rect 1270 1568 1274 1572
rect 1294 1568 1298 1572
rect 1414 1568 1418 1572
rect 1774 1568 1778 1572
rect 2014 1568 2018 1572
rect 2558 1568 2562 1572
rect 118 1558 122 1562
rect 454 1558 458 1562
rect 814 1558 818 1562
rect 38 1548 42 1552
rect 62 1548 66 1552
rect 230 1548 234 1552
rect 254 1548 258 1552
rect 326 1548 330 1552
rect 406 1548 410 1552
rect 102 1538 106 1542
rect 126 1538 130 1542
rect 190 1538 194 1542
rect 206 1538 210 1542
rect 302 1538 306 1542
rect 430 1538 434 1542
rect 470 1548 474 1552
rect 478 1548 482 1552
rect 486 1548 490 1552
rect 582 1547 586 1551
rect 686 1548 690 1552
rect 782 1548 786 1552
rect 790 1548 794 1552
rect 798 1548 802 1552
rect 1062 1558 1066 1562
rect 838 1548 842 1552
rect 862 1548 866 1552
rect 886 1548 890 1552
rect 894 1548 898 1552
rect 934 1548 938 1552
rect 998 1548 1002 1552
rect 1006 1548 1010 1552
rect 1046 1548 1050 1552
rect 1134 1558 1138 1562
rect 1102 1548 1106 1552
rect 1158 1548 1162 1552
rect 1206 1548 1210 1552
rect 1270 1548 1274 1552
rect 1422 1558 1426 1562
rect 1462 1558 1466 1562
rect 1310 1548 1314 1552
rect 1358 1548 1362 1552
rect 1502 1558 1506 1562
rect 1638 1558 1642 1562
rect 1950 1558 1954 1562
rect 2006 1558 2010 1562
rect 2462 1558 2466 1562
rect 1494 1548 1498 1552
rect 510 1538 514 1542
rect 566 1538 570 1542
rect 662 1538 666 1542
rect 750 1538 754 1542
rect 1606 1547 1610 1551
rect 1662 1548 1666 1552
rect 1686 1548 1690 1552
rect 822 1538 826 1542
rect 846 1538 850 1542
rect 910 1538 914 1542
rect 1038 1538 1042 1542
rect 1070 1538 1074 1542
rect 1110 1538 1114 1542
rect 1118 1538 1122 1542
rect 1174 1538 1178 1542
rect 1222 1538 1226 1542
rect 1262 1538 1266 1542
rect 1318 1538 1322 1542
rect 1334 1538 1338 1542
rect 1438 1538 1442 1542
rect 1446 1538 1450 1542
rect 1462 1538 1466 1542
rect 1494 1538 1498 1542
rect 1518 1538 1522 1542
rect 1622 1538 1626 1542
rect 1654 1538 1658 1542
rect 1694 1538 1698 1542
rect 1718 1548 1722 1552
rect 1758 1548 1762 1552
rect 1790 1548 1794 1552
rect 1814 1548 1818 1552
rect 1822 1548 1826 1552
rect 1862 1548 1866 1552
rect 1934 1548 1938 1552
rect 1950 1548 1954 1552
rect 1966 1548 1970 1552
rect 2014 1548 2018 1552
rect 2030 1548 2034 1552
rect 2046 1548 2050 1552
rect 2062 1548 2066 1552
rect 2078 1548 2082 1552
rect 2086 1548 2090 1552
rect 2110 1548 2114 1552
rect 2142 1548 2146 1552
rect 2150 1548 2154 1552
rect 2158 1548 2162 1552
rect 2190 1548 2194 1552
rect 2206 1548 2210 1552
rect 2230 1548 2234 1552
rect 2238 1548 2242 1552
rect 2246 1548 2250 1552
rect 2254 1548 2258 1552
rect 2278 1548 2282 1552
rect 2302 1548 2306 1552
rect 2318 1548 2322 1552
rect 2518 1558 2522 1562
rect 2350 1547 2354 1551
rect 2486 1548 2490 1552
rect 2542 1548 2546 1552
rect 2590 1548 2594 1552
rect 2598 1548 2602 1552
rect 1726 1538 1730 1542
rect 1750 1538 1754 1542
rect 1870 1538 1874 1542
rect 1926 1538 1930 1542
rect 1958 1538 1962 1542
rect 1990 1538 1994 1542
rect 2038 1538 2042 1542
rect 2118 1538 2122 1542
rect 2134 1538 2138 1542
rect 2310 1538 2314 1542
rect 2334 1538 2338 1542
rect 2422 1538 2426 1542
rect 2438 1538 2442 1542
rect 2446 1538 2450 1542
rect 2494 1538 2498 1542
rect 2502 1538 2506 1542
rect 2534 1538 2538 1542
rect 2550 1538 2554 1542
rect 390 1528 394 1532
rect 422 1528 426 1532
rect 534 1528 538 1532
rect 1142 1528 1146 1532
rect 1694 1528 1698 1532
rect 1702 1528 1706 1532
rect 1742 1528 1746 1532
rect 2166 1528 2170 1532
rect 2294 1528 2298 1532
rect 110 1518 114 1522
rect 286 1518 290 1522
rect 382 1518 386 1522
rect 1126 1518 1130 1522
rect 1150 1518 1154 1522
rect 1734 1518 1738 1522
rect 1982 1518 1986 1522
rect 2126 1518 2130 1522
rect 2470 1518 2474 1522
rect 1058 1503 1062 1507
rect 1065 1503 1069 1507
rect 2082 1503 2086 1507
rect 2089 1503 2093 1507
rect 94 1488 98 1492
rect 326 1488 330 1492
rect 398 1488 402 1492
rect 582 1488 586 1492
rect 758 1488 762 1492
rect 982 1488 986 1492
rect 1222 1488 1226 1492
rect 1366 1488 1370 1492
rect 1398 1488 1402 1492
rect 1526 1488 1530 1492
rect 1574 1488 1578 1492
rect 1598 1488 1602 1492
rect 1646 1488 1650 1492
rect 1678 1488 1682 1492
rect 1870 1488 1874 1492
rect 2206 1488 2210 1492
rect 2414 1488 2418 1492
rect 2502 1488 2506 1492
rect 102 1478 106 1482
rect 366 1478 370 1482
rect 854 1478 858 1482
rect 918 1478 922 1482
rect 1190 1478 1194 1482
rect 14 1468 18 1472
rect 134 1468 138 1472
rect 182 1468 186 1472
rect 238 1468 242 1472
rect 302 1468 306 1472
rect 422 1468 426 1472
rect 486 1468 490 1472
rect 502 1468 506 1472
rect 598 1468 602 1472
rect 806 1468 810 1472
rect 870 1468 874 1472
rect 1102 1468 1106 1472
rect 1206 1468 1210 1472
rect 1270 1468 1274 1472
rect 1318 1468 1322 1472
rect 1334 1468 1338 1472
rect 1350 1468 1354 1472
rect 1830 1478 1834 1482
rect 1542 1468 1546 1472
rect 1582 1468 1586 1472
rect 1670 1468 1674 1472
rect 1742 1468 1746 1472
rect 1854 1468 1858 1472
rect 1918 1468 1922 1472
rect 2014 1468 2018 1472
rect 2054 1468 2058 1472
rect 2070 1468 2074 1472
rect 2174 1468 2178 1472
rect 2230 1468 2234 1472
rect 2270 1468 2274 1472
rect 2318 1468 2322 1472
rect 2334 1468 2338 1472
rect 2422 1468 2426 1472
rect 2454 1468 2458 1472
rect 2470 1468 2474 1472
rect 2478 1468 2482 1472
rect 2582 1468 2586 1472
rect 2646 1468 2650 1472
rect 38 1458 42 1462
rect 118 1458 122 1462
rect 142 1458 146 1462
rect 190 1458 194 1462
rect 198 1458 202 1462
rect 222 1458 226 1462
rect 310 1458 314 1462
rect 318 1458 322 1462
rect 374 1458 378 1462
rect 382 1458 386 1462
rect 406 1458 410 1462
rect 526 1458 530 1462
rect 614 1458 618 1462
rect 622 1458 626 1462
rect 654 1458 658 1462
rect 662 1458 666 1462
rect 670 1458 674 1462
rect 702 1458 706 1462
rect 710 1458 714 1462
rect 718 1458 722 1462
rect 742 1458 746 1462
rect 822 1459 826 1463
rect 902 1458 906 1462
rect 918 1458 922 1462
rect 966 1458 970 1462
rect 974 1458 978 1462
rect 998 1458 1002 1462
rect 1022 1458 1026 1462
rect 1070 1458 1074 1462
rect 1126 1458 1130 1462
rect 1198 1458 1202 1462
rect 1214 1458 1218 1462
rect 1270 1458 1274 1462
rect 1350 1458 1354 1462
rect 1374 1458 1378 1462
rect 1382 1458 1386 1462
rect 1430 1458 1434 1462
rect 1454 1458 1458 1462
rect 1486 1458 1490 1462
rect 1510 1458 1514 1462
rect 1614 1458 1618 1462
rect 1734 1458 1738 1462
rect 1774 1458 1778 1462
rect 1782 1458 1786 1462
rect 1838 1458 1842 1462
rect 1934 1459 1938 1463
rect 1974 1458 1978 1462
rect 1998 1458 2002 1462
rect 2006 1458 2010 1462
rect 2022 1458 2026 1462
rect 2030 1458 2034 1462
rect 2038 1458 2042 1462
rect 2062 1458 2066 1462
rect 2150 1458 2154 1462
rect 2190 1458 2194 1462
rect 2230 1458 2234 1462
rect 2254 1458 2258 1462
rect 2262 1458 2266 1462
rect 2302 1458 2306 1462
rect 2310 1458 2314 1462
rect 2358 1458 2362 1462
rect 2430 1458 2434 1462
rect 2558 1458 2562 1462
rect 102 1448 106 1452
rect 142 1448 146 1452
rect 166 1448 170 1452
rect 638 1448 642 1452
rect 1014 1448 1018 1452
rect 1062 1448 1066 1452
rect 1318 1448 1322 1452
rect 1446 1448 1450 1452
rect 1478 1448 1482 1452
rect 1494 1448 1498 1452
rect 1582 1448 1586 1452
rect 1598 1448 1602 1452
rect 1630 1448 1634 1452
rect 2046 1448 2050 1452
rect 2286 1448 2290 1452
rect 2454 1448 2458 1452
rect 990 1438 994 1442
rect 1022 1438 1026 1442
rect 1030 1438 1034 1442
rect 1078 1438 1082 1442
rect 1430 1438 1434 1442
rect 1614 1438 1618 1442
rect 2094 1438 2098 1442
rect 2494 1438 2498 1442
rect 2518 1438 2522 1442
rect 1622 1428 1626 1432
rect 214 1418 218 1422
rect 678 1418 682 1422
rect 734 1418 738 1422
rect 958 1418 962 1422
rect 1070 1418 1074 1422
rect 1182 1418 1186 1422
rect 1398 1418 1402 1422
rect 1430 1418 1434 1422
rect 1454 1418 1458 1422
rect 1486 1418 1490 1422
rect 1526 1418 1530 1422
rect 1550 1418 1554 1422
rect 1662 1418 1666 1422
rect 1798 1418 1802 1422
rect 1982 1418 1986 1422
rect 2486 1418 2490 1422
rect 2606 1418 2610 1422
rect 546 1403 550 1407
rect 553 1403 557 1407
rect 1562 1403 1566 1407
rect 1569 1403 1573 1407
rect 94 1388 98 1392
rect 350 1388 354 1392
rect 702 1388 706 1392
rect 750 1388 754 1392
rect 902 1388 906 1392
rect 1318 1388 1322 1392
rect 1342 1388 1346 1392
rect 1374 1388 1378 1392
rect 1390 1388 1394 1392
rect 1414 1388 1418 1392
rect 1438 1388 1442 1392
rect 1462 1388 1466 1392
rect 1534 1388 1538 1392
rect 1558 1388 1562 1392
rect 1598 1388 1602 1392
rect 1686 1388 1690 1392
rect 1950 1388 1954 1392
rect 2070 1388 2074 1392
rect 2118 1388 2122 1392
rect 2238 1388 2242 1392
rect 2638 1388 2642 1392
rect 1038 1378 1042 1382
rect 342 1368 346 1372
rect 1006 1368 1010 1372
rect 1934 1368 1938 1372
rect 566 1358 570 1362
rect 582 1358 586 1362
rect 870 1358 874 1362
rect 998 1358 1002 1362
rect 1022 1358 1026 1362
rect 1046 1358 1050 1362
rect 38 1348 42 1352
rect 118 1348 122 1352
rect 150 1348 154 1352
rect 158 1348 162 1352
rect 190 1348 194 1352
rect 198 1348 202 1352
rect 206 1348 210 1352
rect 238 1348 242 1352
rect 246 1348 250 1352
rect 278 1348 282 1352
rect 294 1348 298 1352
rect 318 1348 322 1352
rect 326 1348 330 1352
rect 406 1348 410 1352
rect 478 1348 482 1352
rect 566 1348 570 1352
rect 686 1348 690 1352
rect 718 1348 722 1352
rect 726 1348 730 1352
rect 734 1348 738 1352
rect 766 1348 770 1352
rect 814 1348 818 1352
rect 870 1348 874 1352
rect 886 1348 890 1352
rect 958 1348 962 1352
rect 1014 1348 1018 1352
rect 1070 1348 1074 1352
rect 1102 1348 1106 1352
rect 1142 1348 1146 1352
rect 1214 1348 1218 1352
rect 1222 1348 1226 1352
rect 1238 1358 1242 1362
rect 1382 1358 1386 1362
rect 1430 1358 1434 1362
rect 1470 1358 1474 1362
rect 1358 1348 1362 1352
rect 1478 1348 1482 1352
rect 1502 1348 1506 1352
rect 1550 1358 1554 1362
rect 1582 1358 1586 1362
rect 1638 1358 1642 1362
rect 2062 1358 2066 1362
rect 2574 1358 2578 1362
rect 1606 1348 1610 1352
rect 1678 1348 1682 1352
rect 1750 1347 1754 1351
rect 1782 1348 1786 1352
rect 1790 1348 1794 1352
rect 1870 1347 1874 1351
rect 1902 1348 1906 1352
rect 1966 1348 1970 1352
rect 1990 1348 1994 1352
rect 1998 1348 2002 1352
rect 2006 1348 2010 1352
rect 2046 1348 2050 1352
rect 2102 1348 2106 1352
rect 2142 1348 2146 1352
rect 2166 1348 2170 1352
rect 2174 1348 2178 1352
rect 2206 1348 2210 1352
rect 14 1338 18 1342
rect 126 1338 130 1342
rect 142 1338 146 1342
rect 454 1338 458 1342
rect 558 1338 562 1342
rect 654 1338 658 1342
rect 782 1338 786 1342
rect 894 1338 898 1342
rect 982 1338 986 1342
rect 1030 1338 1034 1342
rect 1078 1338 1082 1342
rect 1094 1338 1098 1342
rect 1150 1338 1154 1342
rect 1206 1338 1210 1342
rect 1254 1338 1258 1342
rect 1262 1338 1266 1342
rect 1366 1338 1370 1342
rect 1398 1338 1402 1342
rect 1406 1338 1410 1342
rect 1446 1338 1450 1342
rect 1454 1338 1458 1342
rect 1478 1338 1482 1342
rect 1502 1338 1506 1342
rect 1542 1338 1546 1342
rect 1566 1338 1570 1342
rect 1606 1338 1610 1342
rect 1654 1338 1658 1342
rect 1742 1338 1746 1342
rect 1766 1338 1770 1342
rect 1942 1338 1946 1342
rect 2014 1338 2018 1342
rect 2030 1338 2034 1342
rect 2046 1338 2050 1342
rect 2078 1338 2082 1342
rect 2126 1338 2130 1342
rect 2198 1338 2202 1342
rect 2302 1347 2306 1351
rect 2334 1348 2338 1352
rect 2406 1348 2410 1352
rect 2422 1348 2426 1352
rect 2502 1347 2506 1351
rect 2534 1348 2538 1352
rect 2550 1348 2554 1352
rect 2590 1348 2594 1352
rect 2614 1348 2618 1352
rect 2318 1338 2322 1342
rect 2398 1338 2402 1342
rect 2414 1338 2418 1342
rect 2518 1338 2522 1342
rect 2542 1338 2546 1342
rect 2582 1338 2586 1342
rect 2590 1338 2594 1342
rect 2606 1338 2610 1342
rect 30 1328 34 1332
rect 230 1328 234 1332
rect 310 1328 314 1332
rect 414 1328 418 1332
rect 598 1328 602 1332
rect 1502 1328 1506 1332
rect 1518 1328 1522 1332
rect 1614 1328 1618 1332
rect 1646 1328 1650 1332
rect 1662 1328 1666 1332
rect 1838 1328 1842 1332
rect 1982 1328 1986 1332
rect 2022 1328 2026 1332
rect 2182 1328 2186 1332
rect 2214 1328 2218 1332
rect 2230 1328 2234 1332
rect 2430 1328 2434 1332
rect 2558 1328 2562 1332
rect 2566 1328 2570 1332
rect 182 1318 186 1322
rect 262 1318 266 1322
rect 534 1318 538 1322
rect 670 1318 674 1322
rect 702 1318 706 1322
rect 862 1318 866 1322
rect 1038 1318 1042 1322
rect 1078 1318 1082 1322
rect 1198 1318 1202 1322
rect 1342 1318 1346 1322
rect 1390 1318 1394 1322
rect 1422 1318 1426 1322
rect 1438 1318 1442 1322
rect 1550 1318 1554 1322
rect 1598 1318 1602 1322
rect 1670 1318 1674 1322
rect 1806 1318 1810 1322
rect 2054 1318 2058 1322
rect 2118 1318 2122 1322
rect 2190 1318 2194 1322
rect 2438 1318 2442 1322
rect 1058 1303 1062 1307
rect 1065 1303 1069 1307
rect 2082 1303 2086 1307
rect 2089 1303 2093 1307
rect 14 1288 18 1292
rect 166 1288 170 1292
rect 254 1288 258 1292
rect 366 1288 370 1292
rect 582 1288 586 1292
rect 782 1288 786 1292
rect 854 1288 858 1292
rect 1030 1288 1034 1292
rect 1302 1288 1306 1292
rect 1406 1288 1410 1292
rect 1590 1288 1594 1292
rect 1622 1288 1626 1292
rect 1718 1288 1722 1292
rect 1758 1288 1762 1292
rect 1942 1288 1946 1292
rect 2038 1288 2042 1292
rect 2246 1288 2250 1292
rect 2270 1288 2274 1292
rect 2422 1288 2426 1292
rect 2502 1288 2506 1292
rect 2630 1288 2634 1292
rect 302 1278 306 1282
rect 542 1278 546 1282
rect 622 1278 626 1282
rect 718 1278 722 1282
rect 982 1278 986 1282
rect 1654 1278 1658 1282
rect 1822 1278 1826 1282
rect 2150 1278 2154 1282
rect 2302 1278 2306 1282
rect 70 1268 74 1272
rect 190 1268 194 1272
rect 222 1268 226 1272
rect 374 1268 378 1272
rect 422 1268 426 1272
rect 438 1268 442 1272
rect 454 1268 458 1272
rect 598 1268 602 1272
rect 662 1268 666 1272
rect 670 1268 674 1272
rect 678 1268 682 1272
rect 790 1268 794 1272
rect 822 1268 826 1272
rect 846 1268 850 1272
rect 1046 1268 1050 1272
rect 1118 1268 1122 1272
rect 1150 1268 1154 1272
rect 1166 1268 1170 1272
rect 1198 1268 1202 1272
rect 1214 1268 1218 1272
rect 1278 1268 1282 1272
rect 1326 1268 1330 1272
rect 1414 1268 1418 1272
rect 1462 1268 1466 1272
rect 1582 1268 1586 1272
rect 1670 1268 1674 1272
rect 1710 1268 1714 1272
rect 1798 1268 1802 1272
rect 1806 1268 1810 1272
rect 1830 1268 1834 1272
rect 2014 1268 2018 1272
rect 2046 1268 2050 1272
rect 2134 1268 2138 1272
rect 2446 1268 2450 1272
rect 2478 1268 2482 1272
rect 110 1258 114 1262
rect 214 1258 218 1262
rect 230 1258 234 1262
rect 262 1258 266 1262
rect 270 1258 274 1262
rect 318 1258 322 1262
rect 382 1258 386 1262
rect 390 1258 394 1262
rect 422 1258 426 1262
rect 470 1258 474 1262
rect 478 1258 482 1262
rect 502 1258 506 1262
rect 518 1258 522 1262
rect 526 1258 530 1262
rect 550 1258 554 1262
rect 558 1258 562 1262
rect 606 1258 610 1262
rect 614 1258 618 1262
rect 638 1258 642 1262
rect 654 1258 658 1262
rect 686 1258 690 1262
rect 726 1258 730 1262
rect 798 1258 802 1262
rect 870 1258 874 1262
rect 878 1258 882 1262
rect 974 1258 978 1262
rect 1014 1258 1018 1262
rect 1094 1258 1098 1262
rect 1142 1258 1146 1262
rect 1174 1258 1178 1262
rect 1294 1258 1298 1262
rect 1350 1258 1354 1262
rect 1422 1258 1426 1262
rect 1430 1258 1434 1262
rect 1470 1258 1474 1262
rect 1478 1258 1482 1262
rect 1502 1258 1506 1262
rect 1526 1258 1530 1262
rect 1550 1258 1554 1262
rect 1558 1258 1562 1262
rect 1638 1258 1642 1262
rect 1646 1258 1650 1262
rect 1654 1258 1658 1262
rect 1670 1258 1674 1262
rect 1686 1258 1690 1262
rect 1734 1258 1738 1262
rect 1790 1258 1794 1262
rect 1838 1258 1842 1262
rect 1878 1259 1882 1263
rect 1910 1258 1914 1262
rect 1950 1258 1954 1262
rect 2022 1258 2026 1262
rect 2054 1258 2058 1262
rect 2094 1258 2098 1262
rect 2102 1258 2106 1262
rect 2190 1258 2194 1262
rect 2214 1258 2218 1262
rect 2254 1258 2258 1262
rect 2262 1258 2266 1262
rect 2286 1258 2290 1262
rect 2294 1258 2298 1262
rect 2350 1258 2354 1262
rect 2374 1258 2378 1262
rect 2438 1258 2442 1262
rect 2454 1258 2458 1262
rect 2542 1258 2546 1262
rect 2558 1258 2562 1262
rect 2598 1258 2602 1262
rect 2638 1258 2642 1262
rect 190 1248 194 1252
rect 406 1248 410 1252
rect 486 1248 490 1252
rect 566 1248 570 1252
rect 582 1248 586 1252
rect 838 1248 842 1252
rect 862 1248 866 1252
rect 1046 1248 1050 1252
rect 1078 1248 1082 1252
rect 1086 1248 1090 1252
rect 1134 1248 1138 1252
rect 1150 1248 1154 1252
rect 1198 1248 1202 1252
rect 1286 1248 1290 1252
rect 1446 1248 1450 1252
rect 1534 1248 1538 1252
rect 1702 1248 1706 1252
rect 1782 1248 1786 1252
rect 1846 1248 1850 1252
rect 2070 1248 2074 1252
rect 2478 1248 2482 1252
rect 2622 1248 2626 1252
rect 454 1238 458 1242
rect 1094 1238 1098 1242
rect 1102 1238 1106 1242
rect 1182 1238 1186 1242
rect 1190 1238 1194 1242
rect 1302 1238 1306 1242
rect 2630 1238 2634 1242
rect 2638 1238 2642 1242
rect 798 1218 802 1222
rect 886 1218 890 1222
rect 918 1218 922 1222
rect 1030 1218 1034 1222
rect 1126 1218 1130 1222
rect 1310 1218 1314 1222
rect 1494 1218 1498 1222
rect 1606 1218 1610 1222
rect 1758 1218 1762 1222
rect 1822 1218 1826 1222
rect 2054 1218 2058 1222
rect 2318 1218 2322 1222
rect 2422 1218 2426 1222
rect 546 1203 550 1207
rect 553 1203 557 1207
rect 1562 1203 1566 1207
rect 1569 1203 1573 1207
rect 254 1188 258 1192
rect 766 1188 770 1192
rect 854 1188 858 1192
rect 926 1188 930 1192
rect 1486 1188 1490 1192
rect 1526 1188 1530 1192
rect 1854 1188 1858 1192
rect 1990 1188 1994 1192
rect 2062 1188 2066 1192
rect 2118 1188 2122 1192
rect 2462 1188 2466 1192
rect 2646 1188 2650 1192
rect 2390 1178 2394 1182
rect 166 1168 170 1172
rect 182 1168 186 1172
rect 1230 1168 1234 1172
rect 1246 1168 1250 1172
rect 1430 1168 1434 1172
rect 1630 1168 1634 1172
rect 2286 1168 2290 1172
rect 70 1148 74 1152
rect 118 1148 122 1152
rect 182 1148 186 1152
rect 206 1158 210 1162
rect 742 1158 746 1162
rect 230 1148 234 1152
rect 238 1148 242 1152
rect 270 1148 274 1152
rect 278 1148 282 1152
rect 334 1148 338 1152
rect 358 1148 362 1152
rect 366 1148 370 1152
rect 374 1148 378 1152
rect 486 1148 490 1152
rect 526 1148 530 1152
rect 574 1148 578 1152
rect 646 1148 650 1152
rect 702 1148 706 1152
rect 710 1148 714 1152
rect 750 1148 754 1152
rect 758 1148 762 1152
rect 782 1148 786 1152
rect 798 1148 802 1152
rect 806 1148 810 1152
rect 830 1148 834 1152
rect 854 1148 858 1152
rect 878 1158 882 1162
rect 1278 1158 1282 1162
rect 902 1148 906 1152
rect 910 1148 914 1152
rect 934 1148 938 1152
rect 1014 1147 1018 1151
rect 1110 1148 1114 1152
rect 1190 1148 1194 1152
rect 1214 1148 1218 1152
rect 1262 1148 1266 1152
rect 1286 1148 1290 1152
rect 1294 1148 1298 1152
rect 1318 1158 1322 1162
rect 1470 1158 1474 1162
rect 1574 1158 1578 1162
rect 1366 1147 1370 1151
rect 1454 1148 1458 1152
rect 1486 1148 1490 1152
rect 1510 1148 1514 1152
rect 1518 1148 1522 1152
rect 2126 1158 2130 1162
rect 2302 1158 2306 1162
rect 1614 1148 1618 1152
rect 1678 1148 1682 1152
rect 1918 1148 1922 1152
rect 6 1138 10 1142
rect 86 1138 90 1142
rect 174 1138 178 1142
rect 222 1138 226 1142
rect 286 1138 290 1142
rect 342 1138 346 1142
rect 406 1138 410 1142
rect 494 1138 498 1142
rect 510 1138 514 1142
rect 534 1138 538 1142
rect 606 1138 610 1142
rect 694 1138 698 1142
rect 726 1138 730 1142
rect 846 1138 850 1142
rect 894 1138 898 1142
rect 1094 1138 1098 1142
rect 1166 1138 1170 1142
rect 1254 1138 1258 1142
rect 1286 1138 1290 1142
rect 1318 1138 1322 1142
rect 1334 1138 1338 1142
rect 1382 1138 1386 1142
rect 1950 1147 1954 1151
rect 2014 1148 2018 1152
rect 2038 1148 2042 1152
rect 2054 1148 2058 1152
rect 2078 1148 2082 1152
rect 2086 1148 2090 1152
rect 2110 1148 2114 1152
rect 2150 1148 2154 1152
rect 2182 1148 2186 1152
rect 2222 1148 2226 1152
rect 2454 1158 2458 1162
rect 2326 1148 2330 1152
rect 2342 1148 2346 1152
rect 2374 1148 2378 1152
rect 2430 1148 2434 1152
rect 2518 1148 2522 1152
rect 2582 1147 2586 1151
rect 1558 1138 1562 1142
rect 1606 1138 1610 1142
rect 1622 1138 1626 1142
rect 1710 1138 1714 1142
rect 1790 1138 1794 1142
rect 1870 1138 1874 1142
rect 2022 1138 2026 1142
rect 2102 1138 2106 1142
rect 2174 1138 2178 1142
rect 2286 1138 2290 1142
rect 2302 1138 2306 1142
rect 2334 1138 2338 1142
rect 2350 1138 2354 1142
rect 2422 1138 2426 1142
rect 2438 1138 2442 1142
rect 2542 1138 2546 1142
rect 2566 1138 2570 1142
rect 310 1128 314 1132
rect 590 1128 594 1132
rect 822 1128 826 1132
rect 1438 1128 1442 1132
rect 1462 1128 1466 1132
rect 1502 1128 1506 1132
rect 2134 1128 2138 1132
rect 2214 1128 2218 1132
rect 2358 1128 2362 1132
rect 2366 1128 2370 1132
rect 2406 1128 2410 1132
rect 2422 1128 2426 1132
rect 2454 1128 2458 1132
rect 294 1118 298 1122
rect 430 1118 434 1122
rect 542 1118 546 1122
rect 686 1118 690 1122
rect 950 1118 954 1122
rect 1150 1118 1154 1122
rect 1446 1118 1450 1122
rect 1734 1118 1738 1122
rect 1878 1118 1882 1122
rect 1886 1118 1890 1122
rect 1990 1118 1994 1122
rect 2166 1118 2170 1122
rect 1058 1103 1062 1107
rect 1065 1103 1069 1107
rect 2082 1103 2086 1107
rect 2089 1103 2093 1107
rect 134 1088 138 1092
rect 286 1088 290 1092
rect 422 1088 426 1092
rect 454 1088 458 1092
rect 686 1088 690 1092
rect 990 1088 994 1092
rect 1046 1088 1050 1092
rect 1126 1088 1130 1092
rect 1174 1088 1178 1092
rect 1246 1088 1250 1092
rect 1270 1088 1274 1092
rect 1398 1088 1402 1092
rect 1438 1088 1442 1092
rect 1526 1088 1530 1092
rect 1662 1088 1666 1092
rect 1830 1088 1834 1092
rect 2030 1088 2034 1092
rect 2054 1088 2058 1092
rect 2134 1088 2138 1092
rect 2230 1088 2234 1092
rect 2310 1088 2314 1092
rect 2462 1088 2466 1092
rect 70 1078 74 1082
rect 190 1078 194 1082
rect 342 1078 346 1082
rect 846 1078 850 1082
rect 6 1068 10 1072
rect 86 1068 90 1072
rect 150 1068 154 1072
rect 206 1068 210 1072
rect 334 1068 338 1072
rect 510 1068 514 1072
rect 550 1068 554 1072
rect 606 1068 610 1072
rect 694 1068 698 1072
rect 726 1068 730 1072
rect 742 1068 746 1072
rect 886 1068 890 1072
rect 926 1068 930 1072
rect 998 1068 1002 1072
rect 1038 1068 1042 1072
rect 1062 1078 1066 1082
rect 1158 1078 1162 1082
rect 1486 1078 1490 1082
rect 1502 1078 1506 1082
rect 2070 1078 2074 1082
rect 2102 1078 2106 1082
rect 2254 1078 2258 1082
rect 2326 1078 2330 1082
rect 2446 1078 2450 1082
rect 2622 1078 2626 1082
rect 1230 1068 1234 1072
rect 1286 1068 1290 1072
rect 1382 1068 1386 1072
rect 1430 1068 1434 1072
rect 1470 1068 1474 1072
rect 1614 1068 1618 1072
rect 1630 1068 1634 1072
rect 1646 1068 1650 1072
rect 1678 1068 1682 1072
rect 1694 1068 1698 1072
rect 1790 1068 1794 1072
rect 1806 1068 1810 1072
rect 1870 1068 1874 1072
rect 1886 1068 1890 1072
rect 1998 1068 2002 1072
rect 2046 1068 2050 1072
rect 2126 1068 2130 1072
rect 2182 1068 2186 1072
rect 2214 1068 2218 1072
rect 2278 1068 2282 1072
rect 2302 1068 2306 1072
rect 2382 1068 2386 1072
rect 2430 1068 2434 1072
rect 2518 1068 2522 1072
rect 2534 1068 2538 1072
rect 2606 1068 2610 1072
rect 2622 1068 2626 1072
rect 78 1058 82 1062
rect 142 1058 146 1062
rect 158 1058 162 1062
rect 174 1058 178 1062
rect 246 1058 250 1062
rect 294 1058 298 1062
rect 302 1058 306 1062
rect 342 1058 346 1062
rect 390 1058 394 1062
rect 398 1058 402 1062
rect 414 1058 418 1062
rect 438 1058 442 1062
rect 446 1058 450 1062
rect 510 1058 514 1062
rect 590 1058 594 1062
rect 622 1059 626 1063
rect 654 1058 658 1062
rect 702 1058 706 1062
rect 774 1059 778 1063
rect 806 1058 810 1062
rect 862 1058 866 1062
rect 878 1058 882 1062
rect 894 1058 898 1062
rect 934 1058 938 1062
rect 1022 1058 1026 1062
rect 1030 1058 1034 1062
rect 1094 1058 1098 1062
rect 1102 1058 1106 1062
rect 1110 1058 1114 1062
rect 1262 1058 1266 1062
rect 1294 1058 1298 1062
rect 1302 1058 1306 1062
rect 1326 1058 1330 1062
rect 1342 1058 1346 1062
rect 1350 1058 1354 1062
rect 1374 1058 1378 1062
rect 1446 1058 1450 1062
rect 1486 1058 1490 1062
rect 1502 1058 1506 1062
rect 1542 1058 1546 1062
rect 1558 1058 1562 1062
rect 1574 1058 1578 1062
rect 1590 1058 1594 1062
rect 1606 1058 1610 1062
rect 1638 1058 1642 1062
rect 1670 1058 1674 1062
rect 1686 1058 1690 1062
rect 1702 1058 1706 1062
rect 1774 1059 1778 1063
rect 1846 1058 1850 1062
rect 1862 1058 1866 1062
rect 1894 1058 1898 1062
rect 1974 1058 1978 1062
rect 2014 1058 2018 1062
rect 2062 1058 2066 1062
rect 2086 1058 2090 1062
rect 2174 1058 2178 1062
rect 2270 1058 2274 1062
rect 2390 1059 2394 1063
rect 2422 1058 2426 1062
rect 2438 1058 2442 1062
rect 2558 1058 2562 1062
rect 2646 1058 2650 1062
rect 374 1048 378 1052
rect 726 1048 730 1052
rect 1270 1048 1274 1052
rect 1318 1048 1322 1052
rect 1454 1048 1458 1052
rect 1630 1048 1634 1052
rect 1662 1048 1666 1052
rect 1822 1048 1826 1052
rect 2230 1048 2234 1052
rect 2262 1048 2266 1052
rect 2294 1048 2298 1052
rect 2318 1048 2322 1052
rect 838 1038 842 1042
rect 1710 1038 1714 1042
rect 2286 1038 2290 1042
rect 14 1028 18 1032
rect 1174 1018 1178 1022
rect 1486 1018 1490 1022
rect 1918 1018 1922 1022
rect 2030 1018 2034 1022
rect 2086 1018 2090 1022
rect 2118 1018 2122 1022
rect 2614 1018 2618 1022
rect 546 1003 550 1007
rect 553 1003 557 1007
rect 1562 1003 1566 1007
rect 1569 1003 1573 1007
rect 182 988 186 992
rect 430 988 434 992
rect 758 988 762 992
rect 1318 988 1322 992
rect 1550 988 1554 992
rect 1782 988 1786 992
rect 1830 988 1834 992
rect 1942 988 1946 992
rect 1974 988 1978 992
rect 2302 988 2306 992
rect 2398 988 2402 992
rect 2566 988 2570 992
rect 2646 978 2650 982
rect 94 968 98 972
rect 326 968 330 972
rect 670 968 674 972
rect 1246 968 1250 972
rect 1494 968 1498 972
rect 2190 968 2194 972
rect 2286 968 2290 972
rect 2614 968 2618 972
rect 118 958 122 962
rect 54 948 58 952
rect 222 958 226 962
rect 342 958 346 962
rect 142 948 146 952
rect 158 948 162 952
rect 166 948 170 952
rect 262 948 266 952
rect 366 948 370 952
rect 406 948 410 952
rect 414 948 418 952
rect 438 948 442 952
rect 446 948 450 952
rect 462 948 466 952
rect 486 958 490 962
rect 622 958 626 962
rect 638 958 642 962
rect 1510 958 1514 962
rect 1606 958 1610 962
rect 1726 958 1730 962
rect 582 948 586 952
rect 638 948 642 952
rect 710 948 714 952
rect 822 948 826 952
rect 830 948 834 952
rect 878 948 882 952
rect 902 948 906 952
rect 910 948 914 952
rect 918 948 922 952
rect 926 948 930 952
rect 1038 948 1042 952
rect 1086 948 1090 952
rect 1102 948 1106 952
rect 30 938 34 942
rect 126 938 130 942
rect 150 938 154 942
rect 198 938 202 942
rect 238 938 242 942
rect 326 938 330 942
rect 350 938 354 942
rect 382 938 386 942
rect 454 938 458 942
rect 486 938 490 942
rect 518 938 522 942
rect 606 938 610 942
rect 646 938 650 942
rect 734 938 738 942
rect 750 938 754 942
rect 814 938 818 942
rect 1182 947 1186 951
rect 1270 948 1274 952
rect 1286 948 1290 952
rect 1294 948 1298 952
rect 1302 948 1306 952
rect 1326 948 1330 952
rect 1342 948 1346 952
rect 1374 948 1378 952
rect 1398 948 1402 952
rect 1430 947 1434 951
rect 1518 948 1522 952
rect 1558 948 1562 952
rect 1582 948 1586 952
rect 1646 948 1650 952
rect 1926 958 1930 962
rect 2374 958 2378 962
rect 2510 958 2514 962
rect 1750 948 1754 952
rect 1774 948 1778 952
rect 1798 948 1802 952
rect 1806 948 1810 952
rect 1822 948 1826 952
rect 1846 948 1850 952
rect 1854 948 1858 952
rect 1870 948 1874 952
rect 1894 948 1898 952
rect 1902 948 1906 952
rect 1910 948 1914 952
rect 1958 948 1962 952
rect 1990 948 1994 952
rect 2022 948 2026 952
rect 958 938 962 942
rect 974 938 978 942
rect 1014 938 1018 942
rect 1062 938 1066 942
rect 1134 938 1138 942
rect 1198 938 1202 942
rect 1382 938 1386 942
rect 1526 938 1530 942
rect 1574 938 1578 942
rect 1726 938 1730 942
rect 1766 938 1770 942
rect 1862 938 1866 942
rect 2142 947 2146 951
rect 2230 948 2234 952
rect 2318 948 2322 952
rect 2382 948 2386 952
rect 2430 948 2434 952
rect 2462 947 2466 951
rect 2518 948 2522 952
rect 2550 948 2554 952
rect 2622 948 2626 952
rect 2158 938 2162 942
rect 2174 938 2178 942
rect 2342 938 2346 942
rect 2358 938 2362 942
rect 2494 938 2498 942
rect 2510 938 2514 942
rect 2590 938 2594 942
rect 2598 938 2602 942
rect 382 928 386 932
rect 1150 928 1154 932
rect 1254 928 1258 932
rect 1398 928 1402 932
rect 1430 928 1434 932
rect 1502 928 1506 932
rect 1638 928 1642 932
rect 1686 928 1690 932
rect 2222 928 2226 932
rect 2326 928 2330 932
rect 2534 928 2538 932
rect 2542 928 2546 932
rect 2574 928 2578 932
rect 2590 928 2594 932
rect 214 918 218 922
rect 390 918 394 922
rect 518 918 522 922
rect 654 918 658 922
rect 838 918 842 922
rect 1358 918 1362 922
rect 1606 918 1610 922
rect 1918 918 1922 922
rect 1942 918 1946 922
rect 1974 918 1978 922
rect 2006 918 2010 922
rect 2046 918 2050 922
rect 2078 918 2082 922
rect 2182 918 2186 922
rect 2334 918 2338 922
rect 2510 918 2514 922
rect 2606 918 2610 922
rect 1058 903 1062 907
rect 1065 903 1069 907
rect 2082 903 2086 907
rect 2089 903 2093 907
rect 166 888 170 892
rect 494 888 498 892
rect 598 888 602 892
rect 606 888 610 892
rect 822 888 826 892
rect 902 888 906 892
rect 934 888 938 892
rect 1486 888 1490 892
rect 1510 888 1514 892
rect 1678 888 1682 892
rect 1790 888 1794 892
rect 1894 888 1898 892
rect 2070 888 2074 892
rect 2150 888 2154 892
rect 2198 888 2202 892
rect 2398 888 2402 892
rect 2414 888 2418 892
rect 2558 888 2562 892
rect 2638 888 2642 892
rect 102 878 106 882
rect 390 878 394 882
rect 918 878 922 882
rect 1046 878 1050 882
rect 1190 878 1194 882
rect 1278 878 1282 882
rect 1614 878 1618 882
rect 1886 878 1890 882
rect 2206 878 2210 882
rect 2550 878 2554 882
rect 14 868 18 872
rect 118 868 122 872
rect 246 868 250 872
rect 262 868 266 872
rect 286 868 290 872
rect 318 868 322 872
rect 406 868 410 872
rect 574 868 578 872
rect 718 868 722 872
rect 726 868 730 872
rect 750 868 754 872
rect 766 868 770 872
rect 782 868 786 872
rect 846 868 850 872
rect 990 868 994 872
rect 1102 868 1106 872
rect 1206 868 1210 872
rect 1350 868 1354 872
rect 1366 868 1370 872
rect 1462 868 1466 872
rect 1494 868 1498 872
rect 1590 868 1594 872
rect 1646 868 1650 872
rect 1734 868 1738 872
rect 1822 868 1826 872
rect 1830 868 1834 872
rect 1854 868 1858 872
rect 38 858 42 862
rect 150 858 154 862
rect 158 858 162 862
rect 222 858 226 862
rect 278 858 282 862
rect 334 858 338 862
rect 390 858 394 862
rect 414 858 418 862
rect 422 858 426 862
rect 454 858 458 862
rect 462 858 466 862
rect 470 858 474 862
rect 478 858 482 862
rect 526 858 530 862
rect 550 858 554 862
rect 566 858 570 862
rect 638 858 642 862
rect 670 859 674 863
rect 742 858 746 862
rect 758 858 762 862
rect 790 858 794 862
rect 798 858 802 862
rect 830 858 834 862
rect 838 858 842 862
rect 998 859 1002 863
rect 1030 858 1034 862
rect 1038 858 1042 862
rect 1062 858 1066 862
rect 1126 858 1130 862
rect 1238 858 1242 862
rect 1246 858 1250 862
rect 1286 858 1290 862
rect 1398 858 1402 862
rect 1414 858 1418 862
rect 1422 858 1426 862
rect 1446 858 1450 862
rect 1454 858 1458 862
rect 1470 858 1474 862
rect 1542 858 1546 862
rect 1574 859 1578 863
rect 1638 858 1642 862
rect 1646 858 1650 862
rect 1686 858 1690 862
rect 1694 858 1698 862
rect 1750 858 1754 862
rect 1822 858 1826 862
rect 1846 858 1850 862
rect 1974 868 1978 872
rect 1990 868 1994 872
rect 2054 868 2058 872
rect 2062 868 2066 872
rect 2142 868 2146 872
rect 2174 868 2178 872
rect 2190 868 2194 872
rect 2238 868 2242 872
rect 2278 868 2282 872
rect 2318 868 2322 872
rect 2470 868 2474 872
rect 2478 868 2482 872
rect 2566 868 2570 872
rect 2582 868 2586 872
rect 1870 858 1874 862
rect 1950 858 1954 862
rect 2054 858 2058 862
rect 2134 858 2138 862
rect 2166 858 2170 862
rect 2182 858 2186 862
rect 2230 858 2234 862
rect 2270 858 2274 862
rect 2286 858 2290 862
rect 2294 858 2298 862
rect 2334 859 2338 863
rect 2574 858 2578 862
rect 262 848 266 852
rect 438 848 442 852
rect 598 848 602 852
rect 702 848 706 852
rect 918 848 922 852
rect 1606 848 1610 852
rect 1830 848 1834 852
rect 1886 848 1890 852
rect 2118 848 2122 852
rect 2150 848 2154 852
rect 2214 848 2218 852
rect 2302 848 2306 852
rect 382 838 386 842
rect 1814 838 1818 842
rect 2134 838 2138 842
rect 2382 838 2386 842
rect 766 818 770 822
rect 1430 818 1434 822
rect 1502 818 1506 822
rect 2230 818 2234 822
rect 2254 818 2258 822
rect 2534 818 2538 822
rect 2638 818 2642 822
rect 546 803 550 807
rect 553 803 557 807
rect 1562 803 1566 807
rect 1569 803 1573 807
rect 798 788 802 792
rect 918 788 922 792
rect 982 788 986 792
rect 1214 788 1218 792
rect 1390 788 1394 792
rect 1446 788 1450 792
rect 1590 788 1594 792
rect 1630 788 1634 792
rect 1654 788 1658 792
rect 1982 788 1986 792
rect 2006 788 2010 792
rect 2206 788 2210 792
rect 2102 778 2106 782
rect 2334 778 2338 782
rect 102 768 106 772
rect 894 768 898 772
rect 1278 768 1282 772
rect 2318 768 2322 772
rect 118 758 122 762
rect 38 748 42 752
rect 694 758 698 762
rect 142 748 146 752
rect 190 748 194 752
rect 254 748 258 752
rect 302 748 306 752
rect 358 748 362 752
rect 406 748 410 752
rect 414 748 418 752
rect 526 748 530 752
rect 638 748 642 752
rect 910 758 914 762
rect 950 758 954 762
rect 966 758 970 762
rect 718 748 722 752
rect 734 748 738 752
rect 742 748 746 752
rect 854 748 858 752
rect 934 748 938 752
rect 942 748 946 752
rect 1006 748 1010 752
rect 1046 748 1050 752
rect 1086 758 1090 762
rect 1294 758 1298 762
rect 1598 758 1602 762
rect 1638 758 1642 762
rect 1966 758 1970 762
rect 2086 758 2090 762
rect 2214 758 2218 762
rect 2262 758 2266 762
rect 2294 758 2298 762
rect 2302 758 2306 762
rect 1134 747 1138 751
rect 1166 748 1170 752
rect 1270 748 1274 752
rect 1334 748 1338 752
rect 1414 748 1418 752
rect 1422 748 1426 752
rect 1430 748 1434 752
rect 1454 748 1458 752
rect 1510 748 1514 752
rect 1654 748 1658 752
rect 1670 748 1674 752
rect 1702 748 1706 752
rect 1710 748 1714 752
rect 1718 748 1722 752
rect 1726 748 1730 752
rect 14 738 18 742
rect 102 738 106 742
rect 118 738 122 742
rect 150 738 154 742
rect 294 738 298 742
rect 446 738 450 742
rect 526 738 530 742
rect 574 738 578 742
rect 662 738 666 742
rect 678 738 682 742
rect 726 738 730 742
rect 774 738 778 742
rect 878 738 882 742
rect 894 738 898 742
rect 950 738 954 742
rect 1038 738 1042 742
rect 1062 738 1066 742
rect 1102 738 1106 742
rect 1118 738 1122 742
rect 1270 738 1274 742
rect 1830 747 1834 751
rect 1878 748 1882 752
rect 1910 748 1914 752
rect 1918 748 1922 752
rect 1950 748 1954 752
rect 1958 748 1962 752
rect 1982 748 1986 752
rect 2102 748 2106 752
rect 2158 748 2162 752
rect 2214 748 2218 752
rect 2230 748 2234 752
rect 2270 748 2274 752
rect 2278 748 2282 752
rect 2318 748 2322 752
rect 2382 748 2386 752
rect 2430 748 2434 752
rect 1478 738 1482 742
rect 1582 738 1586 742
rect 1598 738 1602 742
rect 1614 740 1618 744
rect 2502 748 2506 752
rect 2614 748 2618 752
rect 1662 738 1666 742
rect 1678 738 1682 742
rect 1782 738 1786 742
rect 1846 738 1850 742
rect 1894 738 1898 742
rect 1902 738 1906 742
rect 1926 738 1930 742
rect 1990 738 1994 742
rect 1998 738 2002 742
rect 2062 738 2066 742
rect 2110 738 2114 742
rect 2126 738 2130 742
rect 2238 738 2242 742
rect 2246 738 2250 742
rect 2262 738 2266 742
rect 2326 738 2330 742
rect 2414 738 2418 742
rect 2438 738 2442 742
rect 2454 738 2458 742
rect 2526 738 2530 742
rect 2638 738 2642 742
rect 182 728 186 732
rect 270 728 274 732
rect 286 728 290 732
rect 334 728 338 732
rect 462 728 466 732
rect 702 728 706 732
rect 1326 728 1330 732
rect 1862 728 1866 732
rect 2454 728 2458 732
rect 246 718 250 722
rect 398 718 402 722
rect 582 718 586 722
rect 918 718 922 722
rect 1022 718 1026 722
rect 1198 718 1202 722
rect 1406 718 1410 722
rect 1558 718 1562 722
rect 1734 718 1738 722
rect 2206 718 2210 722
rect 2294 718 2298 722
rect 2462 718 2466 722
rect 2558 718 2562 722
rect 1058 703 1062 707
rect 1065 703 1069 707
rect 2082 703 2086 707
rect 2089 703 2093 707
rect 14 688 18 692
rect 238 688 242 692
rect 262 688 266 692
rect 374 688 378 692
rect 534 688 538 692
rect 582 688 586 692
rect 886 688 890 692
rect 966 688 970 692
rect 1246 688 1250 692
rect 1302 688 1306 692
rect 1398 688 1402 692
rect 1422 688 1426 692
rect 1510 688 1514 692
rect 1654 688 1658 692
rect 1686 688 1690 692
rect 1710 688 1714 692
rect 1870 688 1874 692
rect 2006 688 2010 692
rect 2126 688 2130 692
rect 2558 688 2562 692
rect 294 678 298 682
rect 406 678 410 682
rect 910 678 914 682
rect 950 678 954 682
rect 1406 678 1410 682
rect 1574 678 1578 682
rect 2038 678 2042 682
rect 2158 678 2162 682
rect 2254 678 2258 682
rect 2310 678 2314 682
rect 2342 678 2346 682
rect 2446 678 2450 682
rect 70 668 74 672
rect 78 668 82 672
rect 182 668 186 672
rect 254 668 258 672
rect 518 668 522 672
rect 542 668 546 672
rect 702 668 706 672
rect 766 668 770 672
rect 782 668 786 672
rect 806 668 810 672
rect 950 668 954 672
rect 982 668 986 672
rect 1110 668 1114 672
rect 1126 668 1130 672
rect 1174 668 1178 672
rect 1222 668 1226 672
rect 1230 668 1234 672
rect 1262 668 1266 672
rect 1278 668 1282 672
rect 1294 668 1298 672
rect 1318 668 1322 672
rect 1390 668 1394 672
rect 1478 668 1482 672
rect 1486 668 1490 672
rect 1606 668 1610 672
rect 1614 668 1618 672
rect 1622 668 1626 672
rect 1630 668 1634 672
rect 1646 668 1650 672
rect 1678 668 1682 672
rect 1694 668 1698 672
rect 1806 668 1810 672
rect 1830 668 1834 672
rect 1894 668 1898 672
rect 1974 668 1978 672
rect 2006 668 2010 672
rect 2030 668 2034 672
rect 2038 668 2042 672
rect 2054 668 2058 672
rect 2070 668 2074 672
rect 2110 668 2114 672
rect 2150 668 2154 672
rect 2158 668 2162 672
rect 2174 668 2178 672
rect 2382 668 2386 672
rect 2550 668 2554 672
rect 2622 668 2626 672
rect 2638 668 2642 672
rect 6 658 10 662
rect 142 658 146 662
rect 198 658 202 662
rect 206 658 210 662
rect 246 658 250 662
rect 278 658 282 662
rect 294 658 298 662
rect 334 658 338 662
rect 342 658 346 662
rect 350 658 354 662
rect 358 658 362 662
rect 422 658 426 662
rect 446 658 450 662
rect 454 658 458 662
rect 470 658 474 662
rect 494 658 498 662
rect 502 658 506 662
rect 510 658 514 662
rect 542 658 546 662
rect 566 658 570 662
rect 574 658 578 662
rect 622 658 626 662
rect 646 658 650 662
rect 654 658 658 662
rect 662 658 666 662
rect 670 658 674 662
rect 694 658 698 662
rect 710 658 714 662
rect 718 658 722 662
rect 742 658 746 662
rect 790 658 794 662
rect 830 658 834 662
rect 894 658 898 662
rect 902 658 906 662
rect 958 658 962 662
rect 1006 658 1010 662
rect 1030 658 1034 662
rect 1038 658 1042 662
rect 1062 658 1066 662
rect 1070 658 1074 662
rect 1102 658 1106 662
rect 1134 658 1138 662
rect 1142 658 1146 662
rect 1166 658 1170 662
rect 1182 658 1186 662
rect 1190 658 1194 662
rect 1214 658 1218 662
rect 1254 658 1258 662
rect 1286 658 1290 662
rect 1294 658 1298 662
rect 1342 658 1346 662
rect 1366 658 1370 662
rect 1374 658 1378 662
rect 1382 658 1386 662
rect 1494 658 1498 662
rect 1518 658 1522 662
rect 1526 658 1530 662
rect 1550 658 1554 662
rect 1558 658 1562 662
rect 1598 658 1602 662
rect 1638 658 1642 662
rect 1670 658 1674 662
rect 1702 658 1706 662
rect 1742 658 1746 662
rect 1774 659 1778 663
rect 1846 658 1850 662
rect 1886 658 1890 662
rect 1966 658 1970 662
rect 1998 658 2002 662
rect 2030 658 2034 662
rect 2078 658 2082 662
rect 2086 658 2090 662
rect 2118 658 2122 662
rect 2150 658 2154 662
rect 2190 658 2194 662
rect 2222 658 2226 662
rect 2238 658 2242 662
rect 2246 658 2250 662
rect 2278 658 2282 662
rect 2318 658 2322 662
rect 2334 658 2338 662
rect 2414 658 2418 662
rect 2422 658 2426 662
rect 2430 658 2434 662
rect 2438 658 2442 662
rect 2462 658 2466 662
rect 2478 658 2482 662
rect 2486 658 2490 662
rect 2510 658 2514 662
rect 2542 658 2546 662
rect 2606 658 2610 662
rect 1110 648 1114 652
rect 1246 648 1250 652
rect 1510 648 1514 652
rect 1582 648 1586 652
rect 1662 648 1666 652
rect 1822 648 1826 652
rect 1990 648 1994 652
rect 2006 648 2010 652
rect 2126 648 2130 652
rect 2502 648 2506 652
rect 2526 648 2530 652
rect 2542 648 2546 652
rect 438 638 442 642
rect 486 638 490 642
rect 1262 638 1266 642
rect 2110 638 2114 642
rect 326 628 330 632
rect 782 628 786 632
rect 1118 618 1122 622
rect 1950 618 1954 622
rect 546 603 550 607
rect 553 603 557 607
rect 1562 603 1566 607
rect 1569 603 1573 607
rect 134 588 138 592
rect 174 588 178 592
rect 446 588 450 592
rect 662 588 666 592
rect 918 588 922 592
rect 966 588 970 592
rect 1078 588 1082 592
rect 1366 588 1370 592
rect 1414 588 1418 592
rect 1454 588 1458 592
rect 1670 588 1674 592
rect 1718 588 1722 592
rect 2038 588 2042 592
rect 2222 588 2226 592
rect 2270 588 2274 592
rect 2558 588 2562 592
rect 2614 588 2618 592
rect 1278 578 1282 582
rect 742 568 746 572
rect 1574 568 1578 572
rect 2582 568 2586 572
rect 606 558 610 562
rect 734 558 738 562
rect 886 558 890 562
rect 1102 558 1106 562
rect 1302 558 1306 562
rect 150 548 154 552
rect 158 548 162 552
rect 182 548 186 552
rect 230 548 234 552
rect 294 548 298 552
rect 302 548 306 552
rect 406 548 410 552
rect 414 548 418 552
rect 422 548 426 552
rect 430 548 434 552
rect 462 548 466 552
rect 510 548 514 552
rect 574 548 578 552
rect 630 548 634 552
rect 638 548 642 552
rect 670 548 674 552
rect 678 548 682 552
rect 694 548 698 552
rect 718 548 722 552
rect 6 538 10 542
rect 70 538 74 542
rect 78 538 82 542
rect 206 538 210 542
rect 382 538 386 542
rect 502 538 506 542
rect 590 538 594 542
rect 686 538 690 542
rect 806 547 810 551
rect 838 548 842 552
rect 854 548 858 552
rect 894 548 898 552
rect 902 548 906 552
rect 926 548 930 552
rect 942 548 946 552
rect 950 548 954 552
rect 982 548 986 552
rect 1022 548 1026 552
rect 1094 548 1098 552
rect 1118 548 1122 552
rect 1150 548 1154 552
rect 1182 548 1186 552
rect 1230 548 1234 552
rect 1318 548 1322 552
rect 1326 548 1330 552
rect 1350 548 1354 552
rect 1374 548 1378 552
rect 1382 548 1386 552
rect 1390 548 1394 552
rect 1398 548 1402 552
rect 1422 548 1426 552
rect 1430 548 1434 552
rect 1446 548 1450 552
rect 1470 548 1474 552
rect 1518 548 1522 552
rect 1606 548 1610 552
rect 1614 548 1618 552
rect 1630 558 1634 562
rect 1990 558 1994 562
rect 2086 558 2090 562
rect 2374 558 2378 562
rect 1686 548 1690 552
rect 1694 548 1698 552
rect 1702 548 1706 552
rect 1734 548 1738 552
rect 1742 548 1746 552
rect 1766 548 1770 552
rect 1782 548 1786 552
rect 1798 548 1802 552
rect 1854 548 1858 552
rect 1902 548 1906 552
rect 1910 548 1914 552
rect 1966 548 1970 552
rect 1974 548 1978 552
rect 1998 548 2002 552
rect 2014 548 2018 552
rect 2022 548 2026 552
rect 2046 548 2050 552
rect 2062 548 2066 552
rect 2094 548 2098 552
rect 798 538 802 542
rect 838 538 842 542
rect 870 538 874 542
rect 1014 538 1018 542
rect 1046 538 1050 542
rect 1134 538 1138 542
rect 1174 538 1178 542
rect 1198 538 1202 542
rect 1334 538 1338 542
rect 1494 538 1498 542
rect 1598 538 1602 542
rect 1646 538 1650 542
rect 2134 547 2138 551
rect 2206 548 2210 552
rect 2238 548 2242 552
rect 2246 548 2250 552
rect 2254 548 2258 552
rect 2262 548 2266 552
rect 2286 548 2290 552
rect 2294 548 2298 552
rect 2310 548 2314 552
rect 2350 548 2354 552
rect 2358 548 2362 552
rect 2366 548 2370 552
rect 2406 547 2410 551
rect 2486 548 2490 552
rect 2510 558 2514 562
rect 2598 558 2602 562
rect 2630 558 2634 562
rect 2534 548 2538 552
rect 2542 548 2546 552
rect 2566 548 2570 552
rect 1790 538 1794 542
rect 1854 538 1858 542
rect 2054 538 2058 542
rect 2118 538 2122 542
rect 2342 538 2346 542
rect 2390 538 2394 542
rect 2478 538 2482 542
rect 2526 538 2530 542
rect 2574 538 2578 542
rect 2606 538 2610 542
rect 310 528 314 532
rect 350 528 354 532
rect 358 528 362 532
rect 614 528 618 532
rect 1134 528 1138 532
rect 1750 528 1754 532
rect 1958 528 1962 532
rect 2318 528 2322 532
rect 286 518 290 522
rect 558 518 562 522
rect 710 518 714 522
rect 1166 518 1170 522
rect 1806 518 1810 522
rect 1918 518 1922 522
rect 2198 518 2202 522
rect 2470 518 2474 522
rect 2502 518 2506 522
rect 1058 503 1062 507
rect 1065 503 1069 507
rect 2082 503 2086 507
rect 2089 503 2093 507
rect 166 488 170 492
rect 326 488 330 492
rect 422 488 426 492
rect 598 488 602 492
rect 622 488 626 492
rect 718 488 722 492
rect 1038 488 1042 492
rect 1590 488 1594 492
rect 1702 488 1706 492
rect 1774 488 1778 492
rect 1958 488 1962 492
rect 2158 488 2162 492
rect 2182 488 2186 492
rect 2230 488 2234 492
rect 2270 488 2274 492
rect 2374 488 2378 492
rect 2382 488 2386 492
rect 2486 488 2490 492
rect 2590 488 2594 492
rect 102 478 106 482
rect 262 478 266 482
rect 390 478 394 482
rect 990 478 994 482
rect 1318 478 1322 482
rect 1510 478 1514 482
rect 2022 478 2026 482
rect 2110 478 2114 482
rect 2494 478 2498 482
rect 2526 478 2530 482
rect 118 468 122 472
rect 278 468 282 472
rect 502 468 506 472
rect 518 468 522 472
rect 542 468 546 472
rect 582 468 586 472
rect 702 468 706 472
rect 798 468 802 472
rect 814 468 818 472
rect 862 468 866 472
rect 878 468 882 472
rect 950 468 954 472
rect 1014 468 1018 472
rect 1102 468 1106 472
rect 1142 468 1146 472
rect 1230 468 1234 472
rect 1254 468 1258 472
rect 1262 468 1266 472
rect 1286 468 1290 472
rect 1390 468 1394 472
rect 1446 468 1450 472
rect 1518 468 1522 472
rect 1566 468 1570 472
rect 1670 468 1674 472
rect 1718 468 1722 472
rect 1750 468 1754 472
rect 1854 468 1858 472
rect 1878 468 1882 472
rect 1990 468 1994 472
rect 2118 468 2122 472
rect 2198 468 2202 472
rect 2302 468 2306 472
rect 2334 468 2338 472
rect 2350 468 2354 472
rect 2358 468 2362 472
rect 2598 468 2602 472
rect 2614 468 2618 472
rect 38 458 42 462
rect 54 458 58 462
rect 150 458 154 462
rect 158 458 162 462
rect 206 458 210 462
rect 230 459 234 463
rect 262 458 266 462
rect 310 458 314 462
rect 318 458 322 462
rect 382 458 386 462
rect 486 459 490 463
rect 574 458 578 462
rect 614 458 618 462
rect 686 459 690 463
rect 782 459 786 463
rect 822 458 826 462
rect 902 458 906 462
rect 926 458 930 462
rect 1030 458 1034 462
rect 1094 458 1098 462
rect 1174 458 1178 462
rect 1246 458 1250 462
rect 1278 458 1282 462
rect 1326 458 1330 462
rect 1398 458 1402 462
rect 1438 458 1442 462
rect 1454 458 1458 462
rect 1462 458 1466 462
rect 1558 458 1562 462
rect 1646 458 1650 462
rect 1686 458 1690 462
rect 1726 458 1730 462
rect 1830 458 1834 462
rect 1918 458 1922 462
rect 1998 458 2002 462
rect 2078 458 2082 462
rect 2126 458 2130 462
rect 2134 458 2138 462
rect 2142 458 2146 462
rect 2166 458 2170 462
rect 2174 458 2178 462
rect 2206 458 2210 462
rect 2214 458 2218 462
rect 2238 458 2242 462
rect 2254 458 2258 462
rect 2262 458 2266 462
rect 2286 458 2290 462
rect 2310 458 2314 462
rect 2414 458 2418 462
rect 2438 458 2442 462
rect 2478 458 2482 462
rect 2526 459 2530 463
rect 534 448 538 452
rect 822 448 826 452
rect 846 448 850 452
rect 982 448 986 452
rect 1230 448 1234 452
rect 1422 448 1426 452
rect 1534 448 1538 452
rect 1558 448 1562 452
rect 1750 448 1754 452
rect 2334 448 2338 452
rect 2374 448 2378 452
rect 2614 448 2618 452
rect 2646 448 2650 452
rect 78 438 82 442
rect 1262 438 1266 442
rect 1382 438 1386 442
rect 2598 438 2602 442
rect 1398 428 1402 432
rect 1222 418 1226 422
rect 1470 418 1474 422
rect 2630 418 2634 422
rect 546 403 550 407
rect 553 403 557 407
rect 1562 403 1566 407
rect 1569 403 1573 407
rect 86 388 90 392
rect 406 388 410 392
rect 662 388 666 392
rect 862 388 866 392
rect 910 388 914 392
rect 1118 388 1122 392
rect 1190 388 1194 392
rect 1278 388 1282 392
rect 1318 388 1322 392
rect 1358 388 1362 392
rect 1526 388 1530 392
rect 1558 388 1562 392
rect 1670 388 1674 392
rect 1702 388 1706 392
rect 1966 388 1970 392
rect 2014 388 2018 392
rect 2134 388 2138 392
rect 2182 388 2186 392
rect 2278 388 2282 392
rect 830 368 834 372
rect 1854 368 1858 372
rect 2350 368 2354 372
rect 2366 368 2370 372
rect 2510 368 2514 372
rect 6 348 10 352
rect 38 348 42 352
rect 62 348 66 352
rect 70 348 74 352
rect 110 348 114 352
rect 118 348 122 352
rect 190 347 194 351
rect 230 348 234 352
rect 254 348 258 352
rect 270 348 274 352
rect 278 348 282 352
rect 302 358 306 362
rect 334 348 338 352
rect 358 358 362 362
rect 630 358 634 362
rect 382 348 386 352
rect 390 348 394 352
rect 414 348 418 352
rect 422 348 426 352
rect 478 347 482 351
rect 502 348 506 352
rect 598 348 602 352
rect 606 348 610 352
rect 638 348 642 352
rect 646 348 650 352
rect 670 348 674 352
rect 678 348 682 352
rect 694 348 698 352
rect 718 358 722 362
rect 2326 358 2330 362
rect 766 347 770 351
rect 798 348 802 352
rect 838 348 842 352
rect 846 348 850 352
rect 870 348 874 352
rect 886 348 890 352
rect 918 348 922 352
rect 926 348 930 352
rect 974 348 978 352
rect 1094 348 1098 352
rect 1102 348 1106 352
rect 1254 348 1258 352
rect 1262 348 1266 352
rect 1286 348 1290 352
rect 1302 348 1306 352
rect 1334 348 1338 352
rect 1342 348 1346 352
rect 1382 348 1386 352
rect 1398 348 1402 352
rect 1430 348 1434 352
rect 1470 348 1474 352
rect 1494 348 1498 352
rect 1614 348 1618 352
rect 1678 348 1682 352
rect 1686 348 1690 352
rect 1718 348 1722 352
rect 1742 348 1746 352
rect 1774 348 1778 352
rect 1814 348 1818 352
rect 1878 348 1882 352
rect 1886 348 1890 352
rect 1942 348 1946 352
rect 1950 348 1954 352
rect 1974 348 1978 352
rect 1990 348 1994 352
rect 2022 348 2026 352
rect 2030 348 2034 352
rect 2038 348 2042 352
rect 2070 348 2074 352
rect 2118 348 2122 352
rect 2142 348 2146 352
rect 2150 348 2154 352
rect 2158 348 2162 352
rect 2190 348 2194 352
rect 2198 348 2202 352
rect 2206 348 2210 352
rect 2254 348 2258 352
rect 2262 348 2266 352
rect 2270 348 2274 352
rect 2350 348 2354 352
rect 2414 348 2418 352
rect 2470 348 2474 352
rect 2494 358 2498 362
rect 2638 358 2642 362
rect 2574 348 2578 352
rect 2614 348 2618 352
rect 14 338 18 342
rect 30 338 34 342
rect 206 338 210 342
rect 222 338 226 342
rect 270 338 274 342
rect 318 338 322 342
rect 326 338 330 342
rect 374 338 378 342
rect 614 338 618 342
rect 686 338 690 342
rect 718 338 722 342
rect 734 338 738 342
rect 782 338 786 342
rect 966 338 970 342
rect 1030 338 1034 342
rect 1054 338 1058 342
rect 1174 338 1178 342
rect 1246 338 1250 342
rect 1422 338 1426 342
rect 1446 338 1450 342
rect 1542 338 1546 342
rect 1590 338 1594 342
rect 1766 338 1770 342
rect 1790 338 1794 342
rect 1934 338 1938 342
rect 2046 338 2050 342
rect 2214 338 2218 342
rect 2310 338 2314 342
rect 2358 338 2362 342
rect 2398 338 2402 342
rect 2446 338 2450 342
rect 2462 338 2466 342
rect 2494 338 2498 342
rect 2510 338 2514 342
rect 2566 338 2570 342
rect 2614 338 2618 342
rect 2630 338 2634 342
rect 54 328 58 332
rect 110 328 114 332
rect 446 328 450 332
rect 1382 328 1386 332
rect 1534 328 1538 332
rect 1726 328 1730 332
rect 1758 328 1762 332
rect 1902 328 1906 332
rect 2094 328 2098 332
rect 2238 328 2242 332
rect 126 318 130 322
rect 294 318 298 322
rect 350 318 354 322
rect 438 318 442 322
rect 542 318 546 322
rect 590 318 594 322
rect 630 318 634 322
rect 1414 318 1418 322
rect 1870 318 1874 322
rect 2054 318 2058 322
rect 2222 318 2226 322
rect 1058 303 1062 307
rect 1065 303 1069 307
rect 2082 303 2086 307
rect 2089 303 2093 307
rect 94 288 98 292
rect 246 288 250 292
rect 358 288 362 292
rect 454 288 458 292
rect 470 288 474 292
rect 598 288 602 292
rect 726 288 730 292
rect 838 288 842 292
rect 950 288 954 292
rect 990 288 994 292
rect 1078 288 1082 292
rect 1206 288 1210 292
rect 1390 288 1394 292
rect 1646 288 1650 292
rect 1710 288 1714 292
rect 1814 288 1818 292
rect 1902 288 1906 292
rect 2022 288 2026 292
rect 2166 288 2170 292
rect 2190 288 2194 292
rect 2222 288 2226 292
rect 2334 288 2338 292
rect 2502 288 2506 292
rect 2534 288 2538 292
rect 462 278 466 282
rect 1286 278 1290 282
rect 1894 278 1898 282
rect 2326 278 2330 282
rect 102 268 106 272
rect 166 268 170 272
rect 294 268 298 272
rect 486 268 490 272
rect 502 268 506 272
rect 606 268 610 272
rect 654 268 658 272
rect 30 259 34 263
rect 62 258 66 262
rect 174 258 178 262
rect 182 258 186 262
rect 206 258 210 262
rect 254 258 258 262
rect 262 258 266 262
rect 302 258 306 262
rect 390 259 394 263
rect 782 268 786 272
rect 870 268 874 272
rect 886 268 890 272
rect 1014 268 1018 272
rect 1046 268 1050 272
rect 1078 268 1082 272
rect 1166 268 1170 272
rect 1270 268 1274 272
rect 1374 268 1378 272
rect 1486 268 1490 272
rect 1510 268 1514 272
rect 1550 268 1554 272
rect 1566 268 1570 272
rect 1654 268 1658 272
rect 1790 268 1794 272
rect 1966 268 1970 272
rect 1998 268 2002 272
rect 2054 268 2058 272
rect 2302 268 2306 272
rect 2382 268 2386 272
rect 2430 268 2434 272
rect 2446 268 2450 272
rect 2478 268 2482 272
rect 2614 268 2618 272
rect 422 258 426 262
rect 486 258 490 262
rect 526 258 530 262
rect 614 258 618 262
rect 638 258 642 262
rect 678 258 682 262
rect 718 258 722 262
rect 790 259 794 263
rect 830 258 834 262
rect 854 258 858 262
rect 862 258 866 262
rect 918 258 922 262
rect 926 258 930 262
rect 934 258 938 262
rect 942 258 946 262
rect 982 258 986 262
rect 1006 258 1010 262
rect 1022 258 1026 262
rect 1142 258 1146 262
rect 1182 258 1186 262
rect 1190 258 1194 262
rect 1214 258 1218 262
rect 1230 258 1234 262
rect 1238 258 1242 262
rect 1350 258 1354 262
rect 1422 258 1426 262
rect 1446 258 1450 262
rect 1494 258 1498 262
rect 1582 259 1586 263
rect 1662 258 1666 262
rect 1758 258 1762 262
rect 1830 258 1834 262
rect 1838 258 1842 262
rect 1846 258 1850 262
rect 1958 258 1962 262
rect 2006 258 2010 262
rect 2046 258 2050 262
rect 2102 259 2106 263
rect 2134 258 2138 262
rect 2174 258 2178 262
rect 2182 258 2186 262
rect 2206 258 2210 262
rect 2262 258 2266 262
rect 2398 259 2402 263
rect 2470 258 2474 262
rect 2486 258 2490 262
rect 2494 258 2498 262
rect 2526 258 2530 262
rect 2598 259 2602 263
rect 614 248 618 252
rect 630 248 634 252
rect 702 248 706 252
rect 1046 248 1050 252
rect 1518 248 1522 252
rect 1686 248 1690 252
rect 2030 248 2034 252
rect 2446 248 2450 252
rect 1406 238 1410 242
rect 1662 238 1666 242
rect 678 218 682 222
rect 1086 218 1090 222
rect 1862 218 1866 222
rect 2318 218 2322 222
rect 546 203 550 207
rect 553 203 557 207
rect 1562 203 1566 207
rect 1569 203 1573 207
rect 6 188 10 192
rect 214 188 218 192
rect 478 188 482 192
rect 750 188 754 192
rect 870 188 874 192
rect 1046 188 1050 192
rect 1166 188 1170 192
rect 1214 188 1218 192
rect 1390 188 1394 192
rect 1678 188 1682 192
rect 1710 188 1714 192
rect 1814 188 1818 192
rect 1982 188 1986 192
rect 2326 188 2330 192
rect 2534 188 2538 192
rect 2550 188 2554 192
rect 518 178 522 182
rect 726 168 730 172
rect 942 168 946 172
rect 2070 168 2074 172
rect 2126 168 2130 172
rect 2566 168 2570 172
rect 102 158 106 162
rect 70 147 74 151
rect 110 148 114 152
rect 118 148 122 152
rect 142 148 146 152
rect 166 158 170 162
rect 182 148 186 152
rect 190 148 194 152
rect 198 148 202 152
rect 134 138 138 142
rect 150 138 154 142
rect 302 147 306 151
rect 350 148 354 152
rect 382 148 386 152
rect 414 148 418 152
rect 574 148 578 152
rect 590 148 594 152
rect 614 158 618 162
rect 910 158 914 162
rect 662 147 666 151
rect 734 148 738 152
rect 742 148 746 152
rect 766 148 770 152
rect 806 147 810 151
rect 838 148 842 152
rect 926 148 930 152
rect 934 148 938 152
rect 974 148 978 152
rect 998 148 1002 152
rect 1062 148 1066 152
rect 1086 148 1090 152
rect 1118 148 1122 152
rect 1134 148 1138 152
rect 1174 148 1178 152
rect 1182 148 1186 152
rect 1198 148 1202 152
rect 1222 148 1226 152
rect 1230 148 1234 152
rect 1294 148 1298 152
rect 1406 148 1410 152
rect 1510 148 1514 152
rect 1590 148 1594 152
rect 1598 148 1602 152
rect 1654 148 1658 152
rect 1662 148 1666 152
rect 1686 148 1690 152
rect 1750 148 1754 152
rect 1774 158 1778 162
rect 1830 148 1834 152
rect 1838 148 1842 152
rect 1870 147 1874 151
rect 1942 148 1946 152
rect 2046 148 2050 152
rect 2110 158 2114 162
rect 2270 158 2274 162
rect 2518 158 2522 162
rect 2542 158 2546 162
rect 2110 148 2114 152
rect 2182 148 2186 152
rect 2222 148 2226 152
rect 2246 148 2250 152
rect 2278 148 2282 152
rect 2286 148 2290 152
rect 2318 148 2322 152
rect 2382 148 2386 152
rect 2502 148 2506 152
rect 2518 148 2522 152
rect 2606 148 2610 152
rect 294 138 298 142
rect 374 138 378 142
rect 422 138 426 142
rect 526 138 530 142
rect 582 138 586 142
rect 614 138 618 142
rect 630 138 634 142
rect 646 138 650 142
rect 1094 138 1098 142
rect 1110 138 1114 142
rect 1318 138 1322 142
rect 1334 138 1338 142
rect 1470 138 1474 142
rect 1486 138 1490 142
rect 1702 138 1706 142
rect 1742 138 1746 142
rect 1774 138 1778 142
rect 1798 138 1802 142
rect 1854 138 1858 142
rect 1966 138 1970 142
rect 2038 138 2042 142
rect 2046 138 2050 142
rect 2118 138 2122 142
rect 2254 138 2258 142
rect 2310 138 2314 142
rect 2390 138 2394 142
rect 2422 138 2426 142
rect 2494 138 2498 142
rect 2526 138 2530 142
rect 70 128 74 132
rect 334 128 338 132
rect 398 128 402 132
rect 878 128 882 132
rect 1134 128 1138 132
rect 1606 128 1610 132
rect 1646 128 1650 132
rect 2190 128 2194 132
rect 2614 128 2618 132
rect 238 118 242 122
rect 366 118 370 122
rect 558 118 562 122
rect 1046 118 1050 122
rect 1238 118 1242 122
rect 1566 118 1570 122
rect 1934 118 1938 122
rect 1982 118 1986 122
rect 2262 118 2266 122
rect 2478 118 2482 122
rect 1058 103 1062 107
rect 1065 103 1069 107
rect 2082 103 2086 107
rect 2089 103 2093 107
rect 62 88 66 92
rect 86 88 90 92
rect 190 88 194 92
rect 198 88 202 92
rect 502 88 506 92
rect 806 88 810 92
rect 814 88 818 92
rect 1198 88 1202 92
rect 1350 88 1354 92
rect 1526 88 1530 92
rect 1654 88 1658 92
rect 1750 88 1754 92
rect 1830 88 1834 92
rect 2014 88 2018 92
rect 2110 88 2114 92
rect 2294 88 2298 92
rect 2446 88 2450 92
rect 2534 88 2538 92
rect 126 78 130 82
rect 710 78 714 82
rect 1078 78 1082 82
rect 6 68 10 72
rect 78 68 82 72
rect 278 68 282 72
rect 294 68 298 72
rect 310 68 314 72
rect 342 68 346 72
rect 414 68 418 72
rect 422 68 426 72
rect 486 68 490 72
rect 646 68 650 72
rect 694 68 698 72
rect 726 68 730 72
rect 870 68 874 72
rect 910 68 914 72
rect 926 68 930 72
rect 958 68 962 72
rect 974 68 978 72
rect 1102 68 1106 72
rect 1142 68 1146 72
rect 1174 68 1178 72
rect 1278 68 1282 72
rect 1294 68 1298 72
rect 1342 68 1346 72
rect 1430 68 1434 72
rect 1446 68 1450 72
rect 1510 68 1514 72
rect 1574 68 1578 72
rect 1686 68 1690 72
rect 1758 68 1762 72
rect 1806 68 1810 72
rect 1910 68 1914 72
rect 1982 68 1986 72
rect 2062 68 2066 72
rect 2134 68 2138 72
rect 2182 68 2186 72
rect 2190 68 2194 72
rect 2254 68 2258 72
rect 2286 68 2290 72
rect 2374 68 2378 72
rect 2390 68 2394 72
rect 2462 68 2466 72
rect 2614 68 2618 72
rect 150 58 154 62
rect 254 58 258 62
rect 334 58 338 62
rect 350 58 354 62
rect 558 58 562 62
rect 654 58 658 62
rect 662 58 666 62
rect 742 59 746 63
rect 878 59 882 63
rect 950 58 954 62
rect 1014 58 1018 62
rect 1126 58 1130 62
rect 1134 58 1138 62
rect 1150 58 1154 62
rect 1254 58 1258 62
rect 1326 58 1330 62
rect 1334 58 1338 62
rect 1390 58 1394 62
rect 1542 58 1546 62
rect 1614 58 1618 62
rect 1710 58 1714 62
rect 1718 58 1722 62
rect 1726 58 1730 62
rect 1766 58 1770 62
rect 1774 58 1778 62
rect 1886 58 1890 62
rect 1958 58 1962 62
rect 2054 58 2058 62
rect 2142 58 2146 62
rect 2150 58 2154 62
rect 2270 58 2274 62
rect 2278 58 2282 62
rect 2350 58 2354 62
rect 2526 58 2530 62
rect 2566 58 2570 62
rect 2598 59 2602 63
rect 94 48 98 52
rect 310 48 314 52
rect 926 48 930 52
rect 1174 48 1178 52
rect 1310 48 1314 52
rect 2166 48 2170 52
rect 2262 48 2266 52
rect 546 3 550 7
rect 553 3 557 7
rect 1562 3 1566 7
rect 1569 3 1573 7
<< metal2 >>
rect 502 2428 506 2432
rect 1198 2428 1202 2432
rect 1526 2428 1530 2432
rect 2286 2428 2290 2432
rect 502 2402 505 2428
rect 544 2403 546 2407
rect 550 2403 553 2407
rect 557 2403 560 2407
rect 1198 2402 1201 2428
rect 1526 2402 1529 2428
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1573 2403 1576 2407
rect 2286 2402 2289 2428
rect 282 2368 286 2371
rect 214 2342 217 2368
rect 294 2342 297 2368
rect 358 2342 361 2348
rect 366 2342 369 2368
rect 446 2342 449 2348
rect 10 2338 14 2341
rect 74 2338 78 2341
rect 226 2338 230 2341
rect 58 2318 62 2321
rect 6 2272 9 2318
rect 6 2132 9 2268
rect 62 2142 65 2288
rect 70 2262 73 2268
rect 86 2262 89 2268
rect 126 2262 129 2268
rect 70 2151 73 2158
rect 10 2118 14 2121
rect 62 2062 65 2128
rect 50 2058 54 2061
rect 6 1942 9 1948
rect 62 1942 65 2058
rect 86 2052 89 2258
rect 118 2142 121 2148
rect 126 2142 129 2148
rect 102 2122 105 2128
rect 98 2088 102 2091
rect 134 2082 137 2318
rect 158 2292 161 2318
rect 190 2272 193 2278
rect 182 2262 185 2268
rect 174 2252 177 2258
rect 150 2152 153 2248
rect 170 2238 174 2241
rect 146 2138 150 2141
rect 162 2118 169 2121
rect 150 2072 153 2088
rect 166 2082 169 2118
rect 190 2082 193 2138
rect 198 2092 201 2148
rect 206 2112 209 2258
rect 138 2068 142 2071
rect 102 2052 105 2068
rect 114 2058 118 2061
rect 114 1948 118 1951
rect 86 1942 89 1948
rect 62 1912 65 1918
rect 62 1862 65 1908
rect 126 1901 129 2068
rect 166 2062 169 2078
rect 134 2042 137 2048
rect 126 1898 134 1901
rect 102 1862 105 1868
rect 122 1858 126 1861
rect 38 1852 41 1858
rect 10 1718 14 1721
rect 14 1472 17 1668
rect 38 1662 41 1668
rect 62 1652 65 1858
rect 110 1752 113 1818
rect 118 1792 121 1848
rect 134 1752 137 1898
rect 142 1872 145 1878
rect 150 1862 153 1928
rect 174 1872 177 2078
rect 190 1952 193 2078
rect 214 2071 217 2248
rect 206 2068 217 2071
rect 222 2242 225 2278
rect 206 2062 209 2068
rect 222 2062 225 2238
rect 238 2142 241 2338
rect 254 2282 257 2288
rect 318 2272 321 2288
rect 422 2282 425 2318
rect 382 2272 385 2278
rect 398 2262 401 2268
rect 422 2262 425 2268
rect 430 2262 433 2268
rect 322 2258 326 2261
rect 338 2258 342 2261
rect 458 2258 462 2261
rect 262 2242 265 2258
rect 334 2252 337 2258
rect 346 2238 350 2241
rect 302 2192 305 2238
rect 254 2122 257 2128
rect 254 2062 257 2118
rect 262 2062 265 2168
rect 302 2142 305 2188
rect 318 2151 321 2158
rect 366 2152 369 2158
rect 374 2142 377 2158
rect 350 2132 353 2138
rect 302 2062 305 2118
rect 274 2058 278 2061
rect 190 1932 193 1948
rect 198 1942 201 1948
rect 206 1942 209 2058
rect 214 2032 217 2058
rect 158 1852 161 1858
rect 142 1752 145 1768
rect 70 1711 73 1747
rect 86 1742 89 1748
rect 70 1708 81 1711
rect 78 1682 81 1708
rect 94 1692 97 1708
rect 122 1668 126 1671
rect 118 1652 121 1658
rect 62 1552 65 1648
rect 38 1482 41 1548
rect 102 1542 105 1568
rect 122 1558 126 1561
rect 102 1502 105 1538
rect 98 1488 102 1491
rect 102 1472 105 1478
rect 14 1342 17 1468
rect 38 1452 41 1458
rect 110 1451 113 1518
rect 118 1462 121 1558
rect 134 1541 137 1738
rect 150 1702 153 1748
rect 158 1712 161 1748
rect 174 1742 177 1868
rect 190 1752 193 1918
rect 198 1862 201 1878
rect 206 1672 209 1938
rect 214 1932 217 1938
rect 214 1782 217 1928
rect 222 1902 225 1948
rect 230 1932 233 1938
rect 238 1761 241 2018
rect 262 1962 265 2058
rect 310 2022 313 2058
rect 326 2052 329 2068
rect 350 2062 353 2078
rect 374 2072 377 2128
rect 382 2122 385 2258
rect 390 2042 393 2148
rect 406 2102 409 2218
rect 454 2182 457 2258
rect 470 2251 473 2348
rect 478 2272 481 2278
rect 486 2272 489 2398
rect 534 2342 537 2368
rect 1034 2358 1038 2361
rect 1090 2358 1094 2361
rect 654 2352 657 2358
rect 926 2352 929 2358
rect 1078 2352 1081 2358
rect 614 2348 622 2351
rect 810 2348 814 2351
rect 978 2348 982 2351
rect 1026 2348 1030 2351
rect 494 2302 497 2338
rect 606 2322 609 2328
rect 526 2272 529 2318
rect 506 2258 510 2261
rect 462 2248 473 2251
rect 462 2192 465 2248
rect 454 2162 457 2178
rect 430 2152 433 2158
rect 470 2152 473 2218
rect 414 2142 417 2148
rect 410 2088 414 2091
rect 426 2078 430 2081
rect 438 2062 441 2148
rect 446 2142 449 2148
rect 494 2132 497 2138
rect 510 2132 513 2138
rect 410 2058 414 2061
rect 270 1962 273 1968
rect 246 1922 249 1958
rect 270 1922 273 1948
rect 278 1942 281 1948
rect 286 1922 289 1928
rect 258 1888 262 1891
rect 270 1862 273 1898
rect 282 1878 286 1881
rect 294 1862 297 2018
rect 318 1882 321 1888
rect 262 1851 265 1858
rect 262 1848 270 1851
rect 230 1758 241 1761
rect 262 1762 265 1768
rect 230 1752 233 1758
rect 238 1742 241 1748
rect 218 1728 222 1731
rect 254 1712 257 1748
rect 250 1688 254 1691
rect 146 1668 150 1671
rect 146 1658 150 1661
rect 166 1652 169 1668
rect 206 1652 209 1658
rect 254 1552 257 1578
rect 130 1538 137 1541
rect 190 1542 193 1548
rect 206 1542 209 1548
rect 134 1482 137 1538
rect 230 1532 233 1548
rect 138 1468 142 1471
rect 138 1458 142 1461
rect 106 1448 113 1451
rect 142 1442 145 1448
rect 94 1392 97 1408
rect 118 1352 121 1358
rect 42 1348 46 1351
rect 126 1342 129 1348
rect 142 1342 145 1358
rect 150 1352 153 1468
rect 158 1352 161 1498
rect 182 1472 185 1488
rect 238 1472 241 1478
rect 186 1468 190 1471
rect 198 1462 201 1468
rect 186 1458 190 1461
rect 166 1452 169 1458
rect 166 1442 169 1448
rect 198 1352 201 1378
rect 214 1352 217 1418
rect 222 1412 225 1458
rect 270 1422 273 1848
rect 314 1778 318 1781
rect 294 1752 297 1768
rect 302 1752 305 1758
rect 326 1752 329 1978
rect 390 1972 393 2038
rect 342 1952 345 1958
rect 366 1942 369 1948
rect 414 1942 417 1948
rect 334 1852 337 1858
rect 342 1762 345 1918
rect 390 1912 393 1938
rect 422 1902 425 2058
rect 438 1992 441 2058
rect 382 1862 385 1868
rect 406 1862 409 1868
rect 430 1862 433 1888
rect 438 1872 441 1878
rect 454 1862 457 2088
rect 470 2082 473 2088
rect 490 2058 494 2061
rect 478 2052 481 2058
rect 494 1982 497 2018
rect 470 1872 473 1918
rect 478 1892 481 1958
rect 510 1942 513 2128
rect 518 2062 521 2218
rect 544 2203 546 2207
rect 550 2203 553 2207
rect 557 2203 560 2207
rect 566 2191 569 2268
rect 574 2262 577 2268
rect 558 2188 569 2191
rect 598 2232 601 2278
rect 558 2172 561 2188
rect 534 2142 537 2148
rect 558 2102 561 2168
rect 526 1952 529 2068
rect 570 2058 574 2061
rect 544 2003 546 2007
rect 550 2003 553 2007
rect 557 2003 560 2007
rect 574 1952 577 1958
rect 490 1938 494 1941
rect 470 1862 473 1868
rect 502 1862 505 1868
rect 354 1858 358 1861
rect 366 1842 369 1858
rect 414 1842 417 1858
rect 422 1852 425 1858
rect 486 1842 489 1848
rect 494 1822 497 1858
rect 518 1842 521 1948
rect 582 1942 585 2098
rect 530 1918 534 1921
rect 526 1862 529 1918
rect 338 1758 342 1761
rect 282 1748 286 1751
rect 350 1751 353 1818
rect 398 1761 401 1818
rect 398 1758 409 1761
rect 350 1748 358 1751
rect 278 1722 281 1748
rect 318 1672 321 1748
rect 334 1742 337 1748
rect 342 1672 345 1678
rect 302 1662 305 1668
rect 350 1662 353 1718
rect 366 1712 369 1738
rect 374 1732 377 1738
rect 366 1672 369 1678
rect 382 1661 385 1758
rect 406 1752 409 1758
rect 394 1748 398 1751
rect 430 1742 433 1778
rect 526 1752 529 1768
rect 534 1752 537 1908
rect 590 1892 593 2118
rect 598 2062 601 2228
rect 614 2162 617 2348
rect 710 2342 713 2348
rect 650 2338 654 2341
rect 622 2242 625 2338
rect 670 2322 673 2338
rect 686 2332 689 2338
rect 762 2318 766 2321
rect 634 2288 638 2291
rect 686 2272 689 2288
rect 658 2268 662 2271
rect 638 2242 641 2268
rect 726 2262 729 2318
rect 750 2282 753 2298
rect 646 2252 649 2258
rect 734 2252 737 2258
rect 670 2162 673 2248
rect 738 2218 742 2221
rect 682 2158 686 2161
rect 614 2152 617 2158
rect 662 2152 665 2158
rect 638 2142 641 2148
rect 618 2138 622 2141
rect 646 2132 649 2138
rect 638 2072 641 2078
rect 654 2062 657 2068
rect 642 1948 646 1951
rect 622 1942 625 1948
rect 654 1941 657 1978
rect 646 1938 657 1941
rect 630 1932 633 1938
rect 550 1852 553 1868
rect 558 1862 561 1868
rect 606 1862 609 1868
rect 614 1862 617 1888
rect 646 1862 649 1938
rect 654 1922 657 1928
rect 662 1922 665 2148
rect 686 2142 689 2148
rect 702 2142 705 2168
rect 682 2058 686 2061
rect 694 2032 697 2058
rect 670 1952 673 1998
rect 702 1982 705 2138
rect 710 2062 713 2078
rect 718 1982 721 2218
rect 742 2172 745 2208
rect 734 2062 737 2078
rect 742 2062 745 2168
rect 750 2152 753 2278
rect 798 2272 801 2328
rect 830 2312 833 2348
rect 886 2342 889 2348
rect 918 2341 921 2348
rect 1110 2342 1113 2348
rect 918 2338 929 2341
rect 870 2302 873 2328
rect 798 2172 801 2268
rect 806 2263 809 2268
rect 806 2258 809 2259
rect 838 2222 841 2278
rect 866 2268 870 2271
rect 878 2262 881 2268
rect 886 2262 889 2288
rect 898 2268 902 2271
rect 850 2258 854 2261
rect 886 2242 889 2258
rect 762 2148 766 2151
rect 750 2082 753 2098
rect 750 2072 753 2078
rect 766 2062 769 2068
rect 746 2058 753 2061
rect 670 1932 673 1948
rect 678 1921 681 1958
rect 686 1952 689 1958
rect 694 1952 697 1968
rect 670 1918 681 1921
rect 654 1872 657 1908
rect 670 1892 673 1918
rect 694 1882 697 1948
rect 594 1858 598 1861
rect 634 1858 638 1861
rect 566 1852 569 1858
rect 670 1852 673 1878
rect 702 1862 705 1938
rect 710 1912 713 1918
rect 718 1862 721 1868
rect 666 1848 670 1851
rect 544 1803 546 1807
rect 550 1803 553 1807
rect 557 1803 560 1807
rect 582 1782 585 1818
rect 558 1752 561 1768
rect 442 1748 446 1751
rect 482 1748 486 1751
rect 570 1748 574 1751
rect 470 1742 473 1748
rect 402 1738 406 1741
rect 414 1732 417 1738
rect 426 1718 430 1721
rect 390 1682 393 1718
rect 454 1712 457 1718
rect 406 1692 409 1708
rect 394 1668 398 1671
rect 382 1658 390 1661
rect 458 1658 462 1661
rect 282 1648 286 1651
rect 318 1542 321 1658
rect 334 1652 337 1658
rect 358 1652 361 1658
rect 374 1652 377 1658
rect 338 1648 342 1651
rect 382 1562 385 1658
rect 398 1651 401 1658
rect 394 1648 401 1651
rect 454 1562 457 1568
rect 470 1552 473 1738
rect 494 1732 497 1748
rect 542 1742 545 1748
rect 494 1722 497 1728
rect 586 1718 590 1721
rect 486 1692 489 1718
rect 502 1682 505 1688
rect 522 1668 526 1671
rect 486 1592 489 1668
rect 534 1662 537 1708
rect 550 1692 553 1718
rect 514 1658 518 1661
rect 594 1658 598 1661
rect 582 1622 585 1658
rect 544 1603 546 1607
rect 550 1603 553 1607
rect 557 1603 560 1607
rect 582 1582 585 1618
rect 486 1552 489 1558
rect 410 1548 414 1551
rect 290 1518 294 1521
rect 302 1472 305 1538
rect 326 1492 329 1548
rect 430 1542 433 1548
rect 478 1542 481 1548
rect 514 1538 518 1541
rect 390 1522 393 1528
rect 422 1522 425 1528
rect 278 1352 281 1368
rect 294 1352 297 1368
rect 234 1348 238 1351
rect 250 1348 254 1351
rect 14 1292 17 1338
rect 10 1138 14 1141
rect 30 1072 33 1328
rect 150 1282 153 1348
rect 170 1288 174 1291
rect 70 1152 73 1268
rect 114 1258 118 1261
rect 118 1152 121 1168
rect 166 1152 169 1168
rect 70 1082 73 1148
rect 174 1142 177 1278
rect 182 1272 185 1318
rect 190 1292 193 1348
rect 190 1262 193 1268
rect 194 1248 198 1251
rect 206 1241 209 1348
rect 302 1341 305 1468
rect 366 1462 369 1478
rect 382 1462 385 1518
rect 390 1502 393 1518
rect 394 1488 398 1491
rect 418 1468 422 1471
rect 386 1458 390 1461
rect 310 1422 313 1458
rect 318 1352 321 1458
rect 350 1392 353 1448
rect 374 1432 377 1458
rect 406 1452 409 1458
rect 338 1368 342 1371
rect 430 1362 433 1538
rect 534 1532 537 1548
rect 566 1542 569 1578
rect 582 1542 585 1547
rect 318 1342 321 1348
rect 302 1338 310 1341
rect 226 1328 230 1331
rect 306 1328 310 1331
rect 214 1262 217 1298
rect 250 1288 254 1291
rect 262 1282 265 1318
rect 326 1312 329 1348
rect 302 1282 305 1288
rect 366 1282 369 1288
rect 382 1281 385 1338
rect 406 1332 409 1348
rect 414 1312 417 1328
rect 374 1278 385 1281
rect 222 1272 225 1278
rect 374 1272 377 1278
rect 422 1272 425 1278
rect 230 1262 233 1268
rect 270 1262 273 1268
rect 254 1258 262 1261
rect 322 1258 326 1261
rect 214 1252 217 1258
rect 198 1238 209 1241
rect 186 1168 190 1171
rect 182 1152 185 1158
rect 86 1072 89 1138
rect 198 1132 201 1238
rect 254 1192 257 1258
rect 210 1158 214 1161
rect 242 1148 246 1151
rect 222 1142 225 1148
rect 230 1132 233 1148
rect 270 1132 273 1148
rect 278 1142 281 1148
rect 290 1138 294 1141
rect 306 1128 310 1131
rect 138 1088 142 1091
rect 150 1072 153 1078
rect 6 1052 9 1068
rect 18 1028 22 1031
rect 30 942 33 1068
rect 174 1062 177 1078
rect 82 1058 86 1061
rect 146 1058 153 1061
rect 162 1058 166 1061
rect 98 968 102 971
rect 118 962 121 998
rect 142 952 145 998
rect 54 942 57 948
rect 14 742 17 868
rect 42 858 46 861
rect 42 748 46 751
rect 14 692 17 738
rect 6 662 9 668
rect 6 542 9 658
rect 42 458 46 461
rect 6 352 9 388
rect 14 342 17 368
rect 38 352 41 368
rect 54 341 57 458
rect 62 352 65 948
rect 150 942 153 1058
rect 182 992 185 1128
rect 190 1082 193 1088
rect 206 1062 209 1068
rect 246 1062 249 1118
rect 286 1092 289 1128
rect 294 1112 297 1118
rect 302 1062 305 1088
rect 294 992 297 1058
rect 326 972 329 1248
rect 358 1152 361 1168
rect 374 1161 377 1268
rect 382 1262 385 1268
rect 394 1258 398 1261
rect 406 1252 409 1268
rect 374 1158 385 1161
rect 334 1142 337 1148
rect 342 1142 345 1148
rect 334 1112 337 1138
rect 366 1132 369 1148
rect 374 1142 377 1148
rect 342 1082 345 1088
rect 334 1062 337 1068
rect 342 1062 345 1078
rect 374 1052 377 1058
rect 158 952 161 958
rect 166 952 169 968
rect 222 952 225 958
rect 262 952 265 958
rect 122 938 126 941
rect 154 938 158 941
rect 102 882 105 918
rect 118 862 121 868
rect 150 862 153 938
rect 198 892 201 938
rect 238 932 241 938
rect 170 888 174 891
rect 162 858 166 861
rect 214 852 217 918
rect 266 868 270 871
rect 222 862 225 868
rect 78 681 81 818
rect 246 812 249 868
rect 278 862 281 948
rect 326 942 329 968
rect 342 962 345 978
rect 350 942 353 958
rect 366 952 369 978
rect 382 942 385 1158
rect 406 1142 409 1148
rect 390 1062 393 1138
rect 398 1062 401 1118
rect 422 1092 425 1258
rect 430 1172 433 1358
rect 454 1342 457 1508
rect 486 1462 489 1468
rect 502 1462 505 1468
rect 478 1352 481 1358
rect 454 1322 457 1338
rect 438 1262 441 1268
rect 414 1062 417 1068
rect 390 942 393 1058
rect 430 1042 433 1118
rect 446 1062 449 1298
rect 454 1272 457 1278
rect 486 1261 489 1458
rect 502 1262 505 1268
rect 518 1262 521 1478
rect 582 1472 585 1488
rect 530 1458 534 1461
rect 544 1403 546 1407
rect 550 1403 553 1407
rect 557 1403 560 1407
rect 566 1362 569 1368
rect 554 1338 558 1341
rect 486 1258 497 1261
rect 454 1232 457 1238
rect 462 1162 465 1228
rect 470 1222 473 1258
rect 478 1252 481 1258
rect 486 1242 489 1248
rect 454 1092 457 1098
rect 406 952 409 958
rect 414 952 417 1038
rect 438 1031 441 1058
rect 430 1028 441 1031
rect 430 992 433 1028
rect 462 962 465 1158
rect 462 952 465 958
rect 286 872 289 938
rect 262 852 265 858
rect 102 742 105 768
rect 122 758 126 761
rect 142 752 145 758
rect 254 752 257 828
rect 118 742 121 748
rect 150 721 153 738
rect 190 732 193 748
rect 150 718 161 721
rect 70 678 81 681
rect 70 672 73 678
rect 78 662 81 668
rect 70 542 73 548
rect 78 442 81 538
rect 86 392 89 658
rect 134 592 137 668
rect 102 482 105 528
rect 142 482 145 658
rect 158 652 161 718
rect 182 712 185 728
rect 270 722 273 728
rect 250 718 254 721
rect 182 672 185 708
rect 270 702 273 718
rect 258 688 262 691
rect 198 662 201 688
rect 238 682 241 688
rect 278 672 281 768
rect 294 742 297 748
rect 286 722 289 728
rect 294 682 297 688
rect 258 668 262 671
rect 278 662 281 668
rect 290 658 294 661
rect 174 592 177 638
rect 150 552 153 558
rect 206 552 209 658
rect 246 652 249 658
rect 234 548 238 551
rect 158 532 161 548
rect 118 462 121 468
rect 150 462 153 518
rect 182 492 185 548
rect 206 542 209 548
rect 246 522 249 648
rect 254 511 257 588
rect 302 582 305 748
rect 246 508 257 511
rect 170 488 174 491
rect 162 458 166 461
rect 226 459 230 462
rect 150 392 153 458
rect 118 352 121 358
rect 54 338 65 341
rect 30 263 33 338
rect 50 328 54 331
rect 62 272 65 338
rect 70 332 73 348
rect 110 332 113 348
rect 94 292 97 328
rect 126 322 129 328
rect 62 262 65 268
rect 102 262 105 268
rect 10 188 14 191
rect 62 92 65 258
rect 106 158 110 161
rect 70 142 73 147
rect 70 122 73 128
rect 86 92 89 158
rect 118 152 121 158
rect 106 148 110 151
rect 126 132 129 258
rect 134 142 137 388
rect 166 262 169 268
rect 174 262 177 338
rect 190 332 193 347
rect 206 342 209 458
rect 226 348 230 351
rect 206 292 209 338
rect 222 332 225 338
rect 246 292 249 508
rect 262 482 265 488
rect 262 462 265 468
rect 270 352 273 568
rect 294 552 297 558
rect 302 552 305 578
rect 310 532 313 548
rect 290 518 294 521
rect 318 472 321 868
rect 338 858 342 861
rect 382 842 385 928
rect 390 882 393 918
rect 406 872 409 948
rect 438 922 441 948
rect 394 858 398 861
rect 386 838 390 841
rect 406 772 409 868
rect 414 862 417 908
rect 422 842 425 858
rect 438 852 441 858
rect 446 851 449 948
rect 454 912 457 938
rect 454 862 457 868
rect 470 862 473 1178
rect 482 1148 486 1151
rect 494 1142 497 1258
rect 518 1182 521 1258
rect 526 1252 529 1258
rect 534 1252 537 1318
rect 542 1272 545 1278
rect 550 1262 553 1278
rect 558 1262 561 1288
rect 566 1252 569 1348
rect 582 1292 585 1358
rect 590 1332 593 1588
rect 598 1522 601 1558
rect 598 1472 601 1518
rect 606 1372 609 1698
rect 614 1462 617 1838
rect 678 1832 681 1858
rect 686 1852 689 1858
rect 714 1768 718 1771
rect 658 1748 662 1751
rect 622 1742 625 1748
rect 646 1692 649 1748
rect 670 1742 673 1768
rect 682 1758 686 1761
rect 702 1752 705 1758
rect 666 1738 670 1741
rect 690 1738 694 1741
rect 710 1712 713 1738
rect 646 1672 649 1688
rect 694 1672 697 1708
rect 726 1702 729 2018
rect 734 1882 737 1888
rect 750 1752 753 2058
rect 762 1948 766 1951
rect 774 1942 777 2158
rect 782 2092 785 2108
rect 790 2072 793 2148
rect 806 2102 809 2118
rect 814 2072 817 2188
rect 838 2152 841 2168
rect 862 2112 865 2148
rect 926 2072 929 2338
rect 1086 2338 1094 2341
rect 934 2142 937 2148
rect 786 2068 790 2071
rect 902 2062 905 2068
rect 926 2062 929 2068
rect 942 2062 945 2298
rect 950 2292 953 2308
rect 974 2272 977 2338
rect 974 2232 977 2268
rect 1006 2262 1009 2328
rect 1026 2318 1030 2321
rect 1056 2303 1058 2307
rect 1062 2303 1065 2307
rect 1069 2303 1072 2307
rect 1078 2302 1081 2338
rect 1086 2322 1089 2338
rect 950 2162 953 2218
rect 1022 2152 1025 2288
rect 1086 2262 1089 2318
rect 1102 2302 1105 2338
rect 1118 2332 1121 2338
rect 1126 2321 1129 2358
rect 1142 2342 1145 2358
rect 1126 2318 1137 2321
rect 1134 2292 1137 2318
rect 1098 2288 1102 2291
rect 1070 2242 1073 2258
rect 1078 2252 1081 2258
rect 1078 2212 1081 2248
rect 1078 2152 1081 2158
rect 1002 2138 1006 2141
rect 982 2118 990 2121
rect 982 2082 985 2118
rect 998 2111 1001 2128
rect 990 2108 1001 2111
rect 990 2092 993 2108
rect 1014 2102 1017 2138
rect 998 2062 1001 2098
rect 1022 2082 1025 2148
rect 1050 2118 1054 2121
rect 1056 2103 1058 2107
rect 1062 2103 1065 2107
rect 1069 2103 1072 2107
rect 1014 2062 1017 2078
rect 1038 2062 1041 2088
rect 1070 2062 1073 2068
rect 1078 2062 1081 2118
rect 794 2058 798 2061
rect 850 2058 854 2061
rect 902 2042 905 2048
rect 862 1992 865 2038
rect 894 2012 897 2018
rect 838 1952 841 1968
rect 850 1958 854 1961
rect 818 1948 822 1951
rect 766 1852 769 1859
rect 766 1742 769 1748
rect 774 1701 777 1938
rect 806 1932 809 1948
rect 870 1942 873 2008
rect 878 1952 881 1988
rect 918 1962 921 2058
rect 934 2052 937 2058
rect 966 2051 969 2058
rect 958 2048 969 2051
rect 934 1962 937 2048
rect 950 1992 953 2018
rect 886 1942 889 1948
rect 918 1942 921 1948
rect 830 1912 833 1918
rect 826 1888 830 1891
rect 846 1862 849 1888
rect 870 1862 873 1938
rect 798 1752 801 1858
rect 838 1852 841 1858
rect 854 1792 857 1798
rect 818 1748 822 1751
rect 842 1748 846 1751
rect 798 1742 801 1748
rect 822 1722 825 1738
rect 846 1732 849 1738
rect 834 1718 838 1721
rect 766 1698 777 1701
rect 702 1692 705 1698
rect 682 1658 686 1661
rect 694 1652 697 1658
rect 666 1648 670 1651
rect 694 1602 697 1648
rect 646 1552 649 1568
rect 686 1552 689 1558
rect 662 1512 665 1538
rect 654 1462 657 1468
rect 670 1462 673 1488
rect 710 1471 713 1698
rect 766 1682 769 1698
rect 754 1658 758 1661
rect 766 1652 769 1678
rect 806 1671 809 1708
rect 802 1668 809 1671
rect 766 1592 769 1628
rect 746 1568 750 1571
rect 798 1552 801 1568
rect 750 1542 753 1548
rect 782 1502 785 1548
rect 790 1542 793 1548
rect 798 1542 801 1548
rect 806 1532 809 1668
rect 846 1612 849 1728
rect 854 1692 857 1738
rect 862 1682 865 1818
rect 886 1802 889 1878
rect 934 1862 937 1878
rect 950 1862 953 1978
rect 958 1962 961 2048
rect 998 2002 1001 2058
rect 1046 2022 1049 2058
rect 1086 2031 1089 2188
rect 1078 2028 1089 2031
rect 994 1948 998 1951
rect 1006 1942 1009 1948
rect 982 1862 985 1868
rect 1006 1862 1009 1888
rect 1022 1862 1025 2018
rect 1078 1982 1081 2028
rect 1078 1952 1081 1978
rect 1086 1972 1089 2018
rect 1102 1972 1105 2268
rect 1114 2258 1118 2261
rect 1142 2252 1145 2338
rect 1158 2332 1161 2338
rect 1158 2272 1161 2328
rect 1166 2292 1169 2298
rect 1174 2272 1177 2398
rect 1754 2368 1758 2371
rect 1946 2368 1950 2371
rect 1182 2352 1185 2368
rect 1246 2352 1249 2368
rect 1262 2362 1265 2368
rect 1262 2352 1265 2358
rect 1322 2348 1326 2351
rect 1230 2322 1233 2338
rect 1110 2142 1113 2147
rect 1110 2062 1113 2128
rect 1126 2062 1129 2168
rect 1142 2162 1145 2248
rect 1150 2192 1153 2258
rect 1194 2218 1198 2221
rect 1206 2172 1209 2318
rect 1222 2312 1225 2318
rect 1238 2311 1241 2348
rect 1382 2342 1385 2368
rect 1606 2362 1609 2368
rect 1394 2358 1398 2361
rect 1466 2358 1470 2361
rect 1422 2352 1425 2358
rect 1534 2352 1537 2358
rect 1398 2342 1401 2348
rect 1230 2308 1241 2311
rect 1278 2312 1281 2338
rect 1294 2332 1297 2338
rect 1222 2262 1225 2288
rect 1206 2152 1209 2168
rect 1170 2148 1174 2151
rect 1198 2142 1201 2148
rect 1178 2138 1182 2141
rect 1142 2132 1145 2138
rect 1158 2122 1161 2128
rect 1214 2122 1217 2128
rect 1142 2092 1145 2108
rect 1150 2062 1153 2118
rect 1222 2092 1225 2098
rect 1190 2082 1193 2088
rect 1166 2072 1169 2078
rect 1170 2058 1174 2061
rect 1118 2032 1121 2058
rect 1194 2048 1198 2051
rect 1082 1918 1086 1921
rect 1030 1862 1033 1918
rect 1046 1902 1049 1918
rect 1056 1903 1058 1907
rect 1062 1903 1065 1907
rect 1069 1903 1072 1907
rect 1066 1888 1070 1891
rect 886 1712 889 1748
rect 870 1662 873 1668
rect 902 1662 905 1798
rect 910 1662 913 1858
rect 942 1852 945 1858
rect 918 1751 921 1818
rect 934 1742 937 1838
rect 950 1742 953 1748
rect 958 1742 961 1778
rect 974 1772 977 1818
rect 990 1792 993 1858
rect 1014 1762 1017 1818
rect 1046 1812 1049 1858
rect 1094 1842 1097 1858
rect 1118 1851 1121 2028
rect 1150 1951 1153 1958
rect 1198 1952 1201 1958
rect 1214 1952 1217 1958
rect 1230 1951 1233 2308
rect 1254 2262 1257 2268
rect 1278 2262 1281 2308
rect 1358 2272 1361 2288
rect 1302 2262 1305 2268
rect 1358 2262 1361 2268
rect 1366 2262 1369 2328
rect 1382 2272 1385 2338
rect 1430 2322 1433 2338
rect 1418 2288 1422 2291
rect 1414 2262 1417 2268
rect 1314 2258 1318 2261
rect 1330 2258 1334 2261
rect 1402 2258 1406 2261
rect 1262 2252 1265 2258
rect 1270 2242 1273 2258
rect 1382 2252 1385 2258
rect 1422 2251 1425 2258
rect 1410 2248 1425 2251
rect 1382 2242 1385 2248
rect 1238 2212 1241 2218
rect 1270 2212 1273 2238
rect 1430 2232 1433 2318
rect 1446 2302 1449 2338
rect 1466 2328 1470 2331
rect 1486 2302 1489 2348
rect 1494 2322 1497 2328
rect 1526 2292 1529 2348
rect 1606 2342 1609 2358
rect 1622 2342 1625 2368
rect 1638 2352 1641 2358
rect 1686 2351 1689 2358
rect 1766 2352 1769 2368
rect 1646 2342 1649 2348
rect 1758 2342 1761 2348
rect 1806 2342 1809 2368
rect 1850 2358 1854 2361
rect 1822 2352 1825 2358
rect 1842 2348 1846 2351
rect 1886 2351 1889 2358
rect 2066 2348 2070 2351
rect 1654 2332 1657 2338
rect 1486 2272 1489 2288
rect 1474 2258 1478 2261
rect 1226 1948 1233 1951
rect 1262 1952 1265 2178
rect 1294 2152 1297 2218
rect 1342 2152 1345 2218
rect 1382 2152 1385 2218
rect 1406 2192 1409 2228
rect 1486 2152 1489 2268
rect 1550 2262 1553 2288
rect 1630 2272 1633 2288
rect 1558 2262 1561 2268
rect 1590 2262 1593 2268
rect 1662 2262 1665 2278
rect 1686 2272 1689 2328
rect 1726 2272 1729 2278
rect 1530 2258 1534 2261
rect 1690 2259 1694 2261
rect 1742 2262 1745 2298
rect 1766 2272 1769 2298
rect 1774 2292 1777 2318
rect 1778 2268 1782 2271
rect 1790 2262 1793 2278
rect 1814 2262 1817 2268
rect 1822 2262 1825 2338
rect 1854 2332 1857 2338
rect 1846 2262 1849 2268
rect 1854 2262 1857 2328
rect 1690 2258 1697 2259
rect 1754 2258 1758 2261
rect 1518 2252 1521 2258
rect 1534 2202 1537 2218
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1573 2203 1576 2207
rect 1614 2172 1617 2258
rect 1526 2152 1529 2158
rect 1314 2148 1318 2151
rect 1602 2148 1606 2151
rect 1270 2112 1273 2148
rect 1350 2142 1353 2148
rect 1486 2142 1489 2148
rect 1294 2132 1297 2138
rect 1422 2132 1425 2138
rect 1330 2118 1334 2121
rect 1498 2118 1502 2121
rect 1366 2082 1369 2118
rect 1410 2088 1414 2091
rect 1278 2062 1281 2078
rect 1270 1952 1273 1958
rect 1142 1872 1145 1938
rect 1182 1922 1185 1938
rect 1158 1872 1161 1888
rect 1206 1872 1209 1878
rect 1178 1868 1182 1871
rect 1126 1863 1129 1868
rect 1142 1862 1145 1868
rect 1214 1862 1217 1868
rect 1198 1852 1201 1858
rect 1222 1852 1225 1948
rect 1230 1872 1233 1938
rect 1262 1902 1265 1948
rect 1286 1942 1289 1968
rect 1302 1932 1305 2068
rect 1350 2042 1353 2058
rect 1314 1958 1318 1961
rect 1350 1951 1353 1958
rect 1310 1942 1313 1948
rect 1318 1942 1321 1948
rect 1358 1942 1361 2068
rect 1366 1942 1369 2078
rect 1414 2072 1417 2078
rect 1462 2072 1465 2078
rect 1478 2062 1481 2078
rect 1466 2058 1470 2061
rect 1422 2052 1425 2058
rect 1446 2042 1449 2048
rect 1422 2032 1425 2038
rect 1410 1968 1414 1971
rect 1422 1952 1425 2018
rect 1454 1952 1457 1968
rect 1502 1952 1505 2068
rect 1510 2062 1513 2118
rect 1550 2092 1553 2148
rect 1542 2072 1545 2078
rect 1622 2072 1625 2258
rect 1682 2168 1686 2171
rect 1742 2151 1745 2158
rect 1758 2142 1761 2158
rect 1774 2142 1777 2168
rect 1674 2138 1678 2141
rect 1718 2082 1721 2138
rect 1782 2132 1785 2258
rect 1790 2162 1793 2238
rect 1814 2152 1817 2238
rect 1822 2232 1825 2258
rect 1830 2242 1833 2248
rect 1838 2161 1841 2218
rect 1846 2192 1849 2248
rect 1870 2192 1873 2338
rect 1958 2282 1961 2318
rect 1966 2282 1969 2298
rect 1998 2292 2001 2348
rect 2038 2342 2041 2348
rect 2214 2342 2217 2348
rect 2222 2342 2225 2348
rect 2246 2342 2249 2358
rect 1986 2288 1990 2291
rect 2010 2288 2014 2291
rect 1954 2278 1958 2281
rect 1902 2252 1905 2258
rect 1834 2158 1841 2161
rect 1870 2162 1873 2188
rect 1842 2148 1846 2151
rect 1790 2142 1793 2148
rect 1822 2132 1825 2138
rect 1830 2072 1833 2078
rect 1634 2068 1638 2071
rect 1534 2042 1537 2048
rect 1542 2032 1545 2058
rect 1550 2042 1553 2048
rect 1534 1992 1537 2028
rect 1574 2022 1577 2068
rect 1598 2062 1601 2068
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1573 2003 1576 2007
rect 1554 1948 1558 1951
rect 1310 1882 1313 1888
rect 1322 1858 1326 1861
rect 1118 1848 1129 1851
rect 1178 1848 1182 1851
rect 998 1752 1001 1758
rect 1014 1748 1022 1751
rect 974 1742 977 1748
rect 966 1682 969 1718
rect 926 1662 929 1678
rect 962 1668 966 1671
rect 938 1658 942 1661
rect 962 1658 966 1661
rect 886 1652 889 1658
rect 910 1582 913 1658
rect 950 1632 953 1658
rect 982 1652 985 1678
rect 990 1652 993 1658
rect 998 1642 1001 1658
rect 974 1632 977 1638
rect 874 1568 878 1571
rect 814 1552 817 1558
rect 822 1542 825 1558
rect 702 1468 713 1471
rect 702 1462 705 1468
rect 718 1462 721 1468
rect 742 1462 745 1498
rect 758 1492 761 1498
rect 806 1472 809 1528
rect 802 1468 806 1471
rect 822 1463 825 1468
rect 626 1458 630 1461
rect 614 1452 617 1458
rect 662 1452 665 1458
rect 710 1452 713 1458
rect 594 1328 598 1331
rect 598 1252 601 1268
rect 606 1262 609 1368
rect 638 1321 641 1448
rect 658 1338 662 1341
rect 638 1318 649 1321
rect 626 1278 630 1281
rect 614 1252 617 1258
rect 582 1232 585 1248
rect 544 1203 546 1207
rect 550 1203 553 1207
rect 557 1203 560 1207
rect 638 1182 641 1258
rect 646 1242 649 1318
rect 670 1292 673 1318
rect 678 1281 681 1418
rect 702 1392 705 1448
rect 734 1352 737 1418
rect 750 1392 753 1448
rect 838 1422 841 1548
rect 862 1542 865 1548
rect 846 1512 849 1538
rect 886 1502 889 1548
rect 894 1542 897 1548
rect 934 1542 937 1548
rect 910 1532 913 1538
rect 854 1482 857 1498
rect 870 1462 873 1468
rect 886 1392 889 1498
rect 902 1462 905 1518
rect 918 1482 921 1498
rect 966 1472 969 1508
rect 982 1492 985 1598
rect 1014 1592 1017 1748
rect 990 1552 993 1568
rect 998 1552 1001 1578
rect 1022 1572 1025 1658
rect 1030 1602 1033 1748
rect 1054 1742 1057 1768
rect 1066 1758 1070 1761
rect 1090 1758 1094 1761
rect 1114 1748 1118 1751
rect 1078 1742 1081 1748
rect 1102 1742 1105 1748
rect 1038 1732 1041 1738
rect 1046 1712 1049 1718
rect 1056 1703 1058 1707
rect 1062 1703 1065 1707
rect 1069 1703 1072 1707
rect 1046 1672 1049 1678
rect 1062 1622 1065 1668
rect 1062 1552 1065 1558
rect 1010 1548 1014 1551
rect 998 1482 1001 1548
rect 1038 1542 1041 1548
rect 1046 1532 1049 1548
rect 1066 1538 1070 1541
rect 1056 1503 1058 1507
rect 1062 1503 1065 1507
rect 1069 1503 1072 1507
rect 966 1462 969 1468
rect 922 1458 926 1461
rect 978 1458 982 1461
rect 1002 1458 1006 1461
rect 1022 1452 1025 1458
rect 1070 1452 1073 1458
rect 994 1438 998 1441
rect 906 1388 910 1391
rect 866 1358 870 1361
rect 818 1348 822 1351
rect 686 1292 689 1348
rect 702 1302 705 1318
rect 718 1292 721 1348
rect 726 1302 729 1348
rect 678 1278 689 1281
rect 722 1278 726 1281
rect 670 1272 673 1278
rect 658 1268 662 1271
rect 678 1262 681 1268
rect 686 1262 689 1278
rect 654 1252 657 1258
rect 654 1222 657 1248
rect 530 1148 534 1151
rect 510 1072 513 1138
rect 534 1112 537 1138
rect 542 1112 545 1118
rect 534 1102 537 1108
rect 550 1072 553 1148
rect 574 1102 577 1148
rect 590 1132 593 1178
rect 606 1132 609 1138
rect 510 1052 513 1058
rect 590 1042 593 1058
rect 544 1003 546 1007
rect 550 1003 553 1007
rect 557 1003 560 1007
rect 482 958 486 961
rect 482 938 486 941
rect 518 922 521 938
rect 490 888 494 891
rect 518 862 521 918
rect 526 862 529 878
rect 550 862 553 868
rect 566 862 569 988
rect 582 942 585 948
rect 606 942 609 1068
rect 622 1063 625 1108
rect 638 1092 641 1178
rect 650 1148 654 1151
rect 678 1112 681 1258
rect 726 1222 729 1258
rect 742 1162 745 1248
rect 766 1192 769 1348
rect 782 1332 785 1338
rect 854 1292 857 1358
rect 886 1352 889 1358
rect 958 1352 961 1418
rect 998 1362 1001 1368
rect 1006 1362 1009 1368
rect 1014 1361 1017 1448
rect 1034 1438 1038 1441
rect 1022 1432 1025 1438
rect 1038 1382 1041 1388
rect 1046 1362 1049 1368
rect 1014 1358 1022 1361
rect 1022 1352 1025 1358
rect 1062 1352 1065 1448
rect 1078 1442 1081 1738
rect 1102 1732 1105 1738
rect 1118 1722 1121 1738
rect 1086 1662 1089 1668
rect 1126 1592 1129 1848
rect 1150 1762 1153 1768
rect 1138 1758 1142 1761
rect 1178 1748 1182 1751
rect 1134 1742 1137 1748
rect 1134 1702 1137 1718
rect 1142 1662 1145 1738
rect 1166 1732 1169 1738
rect 1182 1722 1185 1728
rect 1198 1692 1201 1848
rect 1270 1782 1273 1818
rect 1334 1782 1337 1938
rect 1374 1882 1377 1888
rect 1270 1771 1273 1778
rect 1262 1768 1273 1771
rect 1162 1668 1166 1671
rect 1150 1662 1153 1668
rect 1106 1548 1110 1551
rect 1106 1538 1110 1541
rect 1110 1512 1113 1538
rect 1102 1472 1105 1488
rect 1118 1482 1121 1538
rect 1134 1532 1137 1558
rect 1158 1542 1161 1548
rect 1174 1542 1177 1688
rect 1230 1682 1233 1748
rect 1246 1742 1249 1747
rect 1262 1742 1265 1768
rect 1322 1748 1326 1751
rect 1294 1732 1297 1748
rect 1342 1742 1345 1778
rect 1382 1752 1385 1868
rect 1398 1862 1401 1868
rect 1390 1832 1393 1858
rect 1422 1852 1425 1948
rect 1430 1882 1433 1948
rect 1462 1882 1465 1888
rect 1430 1872 1433 1878
rect 1474 1858 1478 1861
rect 1414 1832 1417 1848
rect 1486 1772 1489 1918
rect 1510 1832 1513 1948
rect 1518 1872 1521 1948
rect 1574 1942 1577 1958
rect 1582 1952 1585 1958
rect 1590 1952 1593 1958
rect 1598 1942 1601 2058
rect 1606 2052 1609 2058
rect 1606 1942 1609 1968
rect 1538 1938 1542 1941
rect 1558 1872 1561 1928
rect 1598 1862 1601 1868
rect 1518 1792 1521 1858
rect 1526 1772 1529 1818
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1573 1803 1576 1807
rect 1606 1772 1609 1938
rect 1622 1862 1625 2068
rect 1630 2042 1633 2048
rect 1646 2042 1649 2068
rect 1710 2062 1713 2068
rect 1846 2062 1849 2088
rect 1782 2058 1790 2061
rect 1646 1912 1649 2038
rect 1670 1952 1673 1958
rect 1694 1942 1697 2058
rect 1742 2018 1750 2021
rect 1734 1952 1737 1978
rect 1742 1932 1745 2018
rect 1782 1992 1785 2058
rect 1790 1952 1793 2008
rect 1790 1932 1793 1948
rect 1798 1942 1801 1948
rect 1806 1942 1809 2058
rect 1846 1992 1849 2038
rect 1854 2012 1857 2138
rect 1910 2082 1913 2268
rect 1934 2262 1937 2268
rect 1966 2262 1969 2278
rect 1990 2272 1993 2278
rect 2038 2272 2041 2338
rect 2134 2332 2137 2338
rect 2080 2303 2082 2307
rect 2086 2303 2089 2307
rect 2093 2303 2096 2307
rect 1998 2222 2001 2258
rect 1926 2142 1929 2178
rect 1934 2132 1937 2138
rect 1942 2122 1945 2148
rect 1902 2042 1905 2058
rect 1942 2022 1945 2068
rect 1950 2062 1953 2218
rect 1958 2142 1961 2148
rect 1966 2122 1969 2158
rect 1982 2142 1985 2168
rect 1990 2112 1993 2118
rect 1966 2092 1969 2098
rect 1822 1952 1825 1958
rect 1870 1952 1873 1988
rect 1842 1948 1846 1951
rect 1718 1922 1721 1928
rect 1638 1882 1641 1888
rect 1650 1878 1654 1881
rect 1658 1868 1662 1871
rect 1694 1862 1697 1918
rect 1710 1862 1713 1878
rect 1742 1862 1745 1928
rect 1750 1862 1753 1888
rect 1790 1862 1793 1878
rect 1806 1861 1809 1938
rect 1806 1858 1814 1861
rect 1622 1792 1625 1838
rect 1654 1792 1657 1808
rect 1694 1772 1697 1858
rect 1366 1742 1369 1748
rect 1306 1738 1310 1741
rect 1326 1732 1329 1738
rect 1198 1662 1201 1668
rect 1214 1662 1217 1678
rect 1230 1672 1233 1678
rect 1246 1662 1249 1708
rect 1278 1662 1281 1728
rect 1362 1678 1366 1681
rect 1390 1672 1393 1728
rect 1398 1672 1401 1678
rect 1406 1672 1409 1678
rect 1286 1662 1289 1668
rect 1326 1662 1329 1668
rect 1370 1658 1374 1661
rect 1394 1658 1398 1661
rect 1206 1652 1209 1658
rect 1246 1582 1249 1658
rect 1254 1652 1257 1658
rect 1294 1642 1297 1658
rect 1258 1578 1262 1581
rect 1302 1581 1305 1658
rect 1298 1578 1305 1581
rect 1294 1572 1297 1578
rect 1274 1568 1278 1571
rect 1206 1552 1209 1568
rect 1270 1552 1273 1558
rect 1358 1552 1361 1558
rect 1142 1532 1145 1538
rect 1130 1518 1134 1521
rect 1142 1502 1145 1528
rect 1150 1482 1153 1518
rect 1186 1478 1190 1481
rect 1206 1472 1209 1538
rect 1222 1532 1225 1538
rect 1262 1512 1265 1538
rect 1130 1458 1134 1461
rect 1194 1458 1198 1461
rect 1206 1442 1209 1468
rect 1214 1462 1217 1508
rect 1222 1492 1225 1498
rect 1270 1472 1273 1478
rect 1266 1458 1270 1461
rect 1070 1402 1073 1418
rect 1078 1362 1081 1438
rect 1182 1412 1185 1418
rect 1242 1358 1246 1361
rect 1070 1352 1073 1358
rect 1214 1352 1217 1358
rect 866 1348 870 1351
rect 1010 1348 1014 1351
rect 1098 1348 1102 1351
rect 1146 1348 1150 1351
rect 1226 1348 1230 1351
rect 782 1282 785 1288
rect 862 1282 865 1318
rect 790 1262 793 1268
rect 798 1242 801 1258
rect 794 1218 798 1221
rect 702 1152 705 1158
rect 798 1152 801 1208
rect 806 1152 809 1278
rect 822 1272 825 1278
rect 846 1272 849 1278
rect 838 1242 841 1248
rect 846 1222 849 1258
rect 862 1252 865 1268
rect 878 1262 881 1278
rect 886 1272 889 1348
rect 1254 1342 1257 1348
rect 1154 1338 1158 1341
rect 870 1252 873 1258
rect 894 1222 897 1338
rect 982 1322 985 1338
rect 1030 1332 1033 1338
rect 1078 1332 1081 1338
rect 1094 1332 1097 1338
rect 982 1312 985 1318
rect 778 1148 782 1151
rect 710 1142 713 1148
rect 690 1138 694 1141
rect 730 1138 734 1141
rect 686 1122 689 1128
rect 682 1088 686 1091
rect 694 1072 697 1138
rect 726 1132 729 1138
rect 742 1072 745 1148
rect 750 1132 753 1148
rect 758 1142 761 1148
rect 722 1068 726 1071
rect 622 1058 625 1059
rect 706 1058 710 1061
rect 654 1052 657 1058
rect 670 972 673 1058
rect 642 958 646 961
rect 574 862 577 868
rect 462 851 465 858
rect 446 848 465 851
rect 406 752 409 758
rect 334 712 337 728
rect 342 662 345 708
rect 358 682 361 748
rect 374 682 377 688
rect 350 662 353 668
rect 390 662 393 738
rect 398 682 401 718
rect 402 678 406 681
rect 334 642 337 658
rect 358 652 361 658
rect 330 628 334 631
rect 350 532 353 538
rect 358 532 361 638
rect 414 582 417 748
rect 446 742 449 748
rect 446 662 449 698
rect 454 662 457 848
rect 422 642 425 658
rect 434 638 438 641
rect 454 622 457 658
rect 446 592 449 608
rect 406 552 409 578
rect 414 552 417 568
rect 422 552 425 558
rect 462 552 465 728
rect 470 722 473 858
rect 478 852 481 858
rect 590 851 593 928
rect 622 902 625 958
rect 702 952 705 1058
rect 726 1052 729 1058
rect 742 1052 745 1068
rect 774 1063 777 1068
rect 758 992 761 1018
rect 710 952 713 958
rect 638 932 641 948
rect 734 942 737 948
rect 750 942 753 948
rect 646 932 649 938
rect 646 912 649 928
rect 598 892 601 898
rect 606 882 609 888
rect 654 862 657 918
rect 590 848 598 851
rect 544 803 546 807
rect 550 803 553 807
rect 557 803 560 807
rect 522 748 526 751
rect 574 742 577 798
rect 598 772 601 848
rect 638 802 641 858
rect 670 852 673 859
rect 702 852 705 938
rect 750 912 753 928
rect 782 922 785 1108
rect 798 1002 801 1148
rect 822 1132 825 1138
rect 830 1112 833 1148
rect 846 1142 849 1218
rect 854 1192 857 1198
rect 854 1152 857 1158
rect 838 1138 846 1141
rect 838 1072 841 1138
rect 846 1082 849 1108
rect 854 1062 857 1148
rect 862 1062 865 1168
rect 878 1162 881 1168
rect 886 1152 889 1218
rect 894 1142 897 1208
rect 902 1162 905 1298
rect 982 1282 985 1308
rect 1038 1302 1041 1318
rect 1056 1303 1058 1307
rect 1062 1303 1065 1307
rect 1069 1303 1072 1307
rect 1034 1288 1038 1291
rect 918 1212 921 1218
rect 926 1192 929 1278
rect 1014 1262 1017 1288
rect 1042 1268 1046 1271
rect 974 1202 977 1258
rect 1078 1252 1081 1318
rect 1094 1262 1097 1298
rect 1050 1248 1054 1251
rect 1090 1248 1094 1251
rect 1102 1242 1105 1308
rect 1150 1272 1153 1278
rect 1166 1272 1169 1328
rect 1198 1322 1201 1328
rect 1206 1312 1209 1338
rect 1198 1272 1201 1298
rect 1214 1272 1217 1338
rect 1254 1332 1257 1338
rect 1262 1332 1265 1338
rect 1114 1268 1118 1271
rect 1170 1268 1174 1271
rect 1198 1262 1201 1268
rect 1178 1258 1182 1261
rect 1134 1252 1137 1258
rect 1094 1232 1097 1238
rect 1030 1162 1033 1218
rect 902 1152 905 1158
rect 930 1148 934 1151
rect 910 1142 913 1148
rect 1014 1142 1017 1147
rect 874 1058 878 1061
rect 718 872 721 878
rect 750 872 753 908
rect 766 872 769 888
rect 782 872 785 918
rect 726 862 729 868
rect 742 852 745 858
rect 638 782 641 798
rect 694 762 697 768
rect 718 752 721 768
rect 734 752 737 758
rect 750 751 753 868
rect 790 862 793 898
rect 806 892 809 1058
rect 862 1052 865 1058
rect 886 1052 889 1068
rect 894 1062 897 1068
rect 838 1042 841 1048
rect 822 952 825 968
rect 818 938 822 941
rect 762 858 766 861
rect 766 832 769 858
rect 766 802 769 818
rect 746 748 753 751
rect 470 662 473 688
rect 518 672 521 678
rect 502 662 505 668
rect 490 658 494 661
rect 482 638 486 641
rect 510 632 513 658
rect 510 552 513 558
rect 430 542 433 548
rect 350 522 353 528
rect 358 492 361 528
rect 330 488 334 491
rect 278 462 281 468
rect 382 462 385 538
rect 390 482 393 488
rect 322 458 326 461
rect 310 452 313 458
rect 298 358 302 361
rect 278 352 281 358
rect 254 322 257 348
rect 270 332 273 338
rect 310 322 313 448
rect 358 362 361 458
rect 358 352 361 358
rect 382 352 385 418
rect 406 392 409 518
rect 426 488 430 491
rect 502 472 505 538
rect 518 492 521 628
rect 518 472 521 488
rect 526 482 529 738
rect 638 732 641 748
rect 662 742 665 748
rect 774 742 777 748
rect 678 722 681 738
rect 706 728 710 731
rect 586 718 590 721
rect 534 692 537 698
rect 542 672 545 688
rect 566 662 569 718
rect 586 688 590 691
rect 698 668 702 671
rect 646 662 649 668
rect 654 662 657 668
rect 662 662 665 668
rect 578 658 582 661
rect 706 658 710 661
rect 542 652 545 658
rect 622 632 625 658
rect 670 651 673 658
rect 662 648 673 651
rect 544 603 546 607
rect 550 603 553 607
rect 557 603 560 607
rect 662 592 665 648
rect 694 582 697 658
rect 718 642 721 658
rect 574 552 577 578
rect 602 558 606 561
rect 678 552 681 558
rect 694 552 697 568
rect 558 522 561 528
rect 574 512 577 548
rect 630 542 633 548
rect 586 538 590 541
rect 638 532 641 548
rect 670 542 673 548
rect 718 542 721 548
rect 618 528 622 531
rect 598 492 601 508
rect 670 492 673 538
rect 686 512 689 538
rect 710 492 713 518
rect 718 492 721 498
rect 626 488 630 491
rect 538 468 542 471
rect 486 463 489 468
rect 502 352 505 468
rect 574 462 577 468
rect 534 452 537 458
rect 582 452 585 468
rect 686 463 689 488
rect 726 472 729 738
rect 766 682 769 728
rect 766 672 769 678
rect 778 668 782 671
rect 790 662 793 828
rect 798 792 801 858
rect 806 672 809 778
rect 814 742 817 938
rect 830 931 833 948
rect 822 928 833 931
rect 878 932 881 948
rect 822 892 825 928
rect 838 902 841 918
rect 830 862 833 888
rect 838 862 841 868
rect 846 832 849 868
rect 886 842 889 1048
rect 910 1032 913 1128
rect 950 1092 953 1118
rect 990 1092 993 1108
rect 1046 1092 1049 1148
rect 1056 1103 1058 1107
rect 1062 1103 1065 1107
rect 1069 1103 1072 1107
rect 902 952 905 978
rect 910 952 913 1028
rect 926 1022 929 1068
rect 934 1052 937 1058
rect 950 982 953 1088
rect 1062 1082 1065 1088
rect 1038 1072 1041 1078
rect 998 1062 1001 1068
rect 1022 1052 1025 1058
rect 918 952 921 958
rect 902 892 905 938
rect 926 912 929 948
rect 958 942 961 948
rect 974 932 977 938
rect 930 888 934 891
rect 918 882 921 888
rect 922 848 926 851
rect 918 792 921 838
rect 982 792 985 908
rect 990 872 993 998
rect 998 863 1001 878
rect 894 762 897 768
rect 914 758 918 761
rect 934 752 937 768
rect 942 762 945 778
rect 954 758 958 761
rect 942 752 945 758
rect 850 748 854 751
rect 878 742 881 748
rect 894 732 897 738
rect 918 702 921 718
rect 890 688 894 691
rect 914 678 918 681
rect 830 662 833 678
rect 894 662 897 668
rect 934 662 937 748
rect 950 712 953 738
rect 966 692 969 758
rect 1014 752 1017 938
rect 1030 912 1033 1058
rect 1038 1042 1041 1068
rect 1086 952 1089 1208
rect 1094 1112 1097 1138
rect 1102 1132 1105 1238
rect 1142 1232 1145 1258
rect 1154 1248 1158 1251
rect 1202 1248 1206 1251
rect 1182 1242 1185 1248
rect 1190 1232 1193 1238
rect 1130 1218 1134 1221
rect 1214 1152 1217 1268
rect 1194 1148 1198 1151
rect 1110 1092 1113 1148
rect 1122 1088 1126 1091
rect 1102 1062 1105 1078
rect 1150 1071 1153 1118
rect 1158 1072 1161 1078
rect 1150 1068 1158 1071
rect 1114 1058 1118 1061
rect 1094 1042 1097 1058
rect 1110 951 1113 1058
rect 1106 948 1113 951
rect 1038 942 1041 948
rect 1062 932 1065 938
rect 1056 903 1058 907
rect 1062 903 1065 907
rect 1069 903 1072 907
rect 1050 878 1054 881
rect 1030 862 1033 868
rect 1006 732 1009 748
rect 1038 742 1041 858
rect 1062 852 1065 858
rect 1086 812 1089 948
rect 1134 942 1137 948
rect 1150 932 1153 968
rect 1102 792 1105 868
rect 1126 862 1129 868
rect 950 682 953 688
rect 982 672 985 678
rect 942 668 950 671
rect 738 658 742 661
rect 790 652 793 658
rect 902 652 905 658
rect 782 632 785 638
rect 918 592 921 638
rect 942 592 945 668
rect 954 658 958 661
rect 966 592 969 648
rect 1006 642 1009 658
rect 746 568 750 571
rect 734 562 737 568
rect 838 552 841 578
rect 802 548 806 551
rect 850 548 854 551
rect 870 542 873 568
rect 886 562 889 578
rect 902 552 905 568
rect 942 552 945 558
rect 890 548 894 551
rect 926 542 929 548
rect 798 482 801 538
rect 798 472 801 478
rect 838 472 841 538
rect 862 492 865 538
rect 862 472 865 488
rect 878 472 881 478
rect 818 468 822 471
rect 614 452 617 458
rect 544 403 546 407
rect 550 403 553 407
rect 557 403 560 407
rect 662 382 665 388
rect 634 358 638 361
rect 338 348 342 351
rect 410 348 414 351
rect 374 342 377 348
rect 382 342 385 348
rect 262 262 265 308
rect 294 291 297 318
rect 318 292 321 338
rect 326 332 329 338
rect 294 288 305 291
rect 250 258 254 261
rect 182 192 185 258
rect 170 158 174 161
rect 142 152 145 158
rect 190 152 193 168
rect 182 142 185 148
rect 198 142 201 148
rect 134 132 137 138
rect 126 82 129 128
rect 6 72 9 78
rect 82 68 86 71
rect 150 62 153 138
rect 190 92 193 138
rect 206 92 209 258
rect 214 192 217 258
rect 238 122 241 138
rect 202 88 206 91
rect 278 72 281 288
rect 294 272 297 278
rect 294 142 297 268
rect 302 262 305 288
rect 326 282 329 328
rect 302 122 305 147
rect 334 132 337 138
rect 294 72 297 88
rect 342 72 345 318
rect 350 262 353 318
rect 390 302 393 348
rect 414 302 417 348
rect 358 292 361 298
rect 422 292 425 348
rect 610 348 614 351
rect 446 322 449 328
rect 438 292 441 318
rect 478 311 481 347
rect 470 308 481 311
rect 454 292 457 298
rect 470 292 473 308
rect 350 142 353 148
rect 374 142 377 288
rect 422 272 425 288
rect 462 282 465 288
rect 390 263 393 268
rect 478 262 481 278
rect 486 272 489 278
rect 502 272 505 348
rect 598 332 601 348
rect 614 332 617 338
rect 538 318 542 321
rect 586 318 590 321
rect 598 292 601 328
rect 610 268 614 271
rect 482 258 486 261
rect 422 232 425 258
rect 502 252 505 268
rect 606 262 609 268
rect 622 261 625 358
rect 694 352 697 378
rect 634 348 638 351
rect 618 258 625 261
rect 526 252 529 258
rect 478 192 481 248
rect 414 152 417 178
rect 370 118 374 121
rect 382 92 385 148
rect 414 138 422 141
rect 398 132 401 138
rect 382 72 385 88
rect 414 72 417 138
rect 502 122 505 228
rect 544 203 546 207
rect 550 203 553 207
rect 557 203 560 207
rect 522 178 526 181
rect 574 152 577 178
rect 586 148 590 151
rect 606 142 609 258
rect 614 242 617 248
rect 622 162 625 258
rect 630 252 633 318
rect 638 262 641 338
rect 646 322 649 348
rect 658 268 662 271
rect 638 212 641 258
rect 670 222 673 348
rect 678 262 681 348
rect 690 338 694 341
rect 702 322 705 468
rect 782 452 785 459
rect 718 362 721 378
rect 718 342 721 348
rect 734 342 737 368
rect 766 351 769 358
rect 798 352 801 358
rect 814 342 817 468
rect 826 458 830 461
rect 846 452 849 458
rect 850 448 854 451
rect 822 442 825 448
rect 826 368 830 371
rect 838 352 841 408
rect 862 392 865 398
rect 870 352 873 368
rect 730 288 734 291
rect 782 272 785 338
rect 838 292 841 338
rect 718 262 721 268
rect 790 263 793 278
rect 830 262 833 268
rect 678 252 681 258
rect 698 248 702 251
rect 678 192 681 218
rect 750 192 753 218
rect 830 192 833 258
rect 846 252 849 348
rect 862 262 865 278
rect 870 272 873 278
rect 730 168 734 171
rect 614 152 617 158
rect 586 138 590 141
rect 502 92 505 118
rect 422 72 425 78
rect 314 68 318 71
rect 346 68 350 71
rect 410 68 414 71
rect 490 68 494 71
rect 254 62 257 68
rect 94 52 97 58
rect 278 52 281 68
rect 330 58 334 61
rect 310 52 313 58
rect 350 52 353 58
rect 526 12 529 138
rect 614 132 617 138
rect 558 92 561 118
rect 558 62 561 68
rect 622 42 625 158
rect 630 142 633 168
rect 734 152 737 158
rect 742 152 745 168
rect 806 151 809 188
rect 854 172 857 258
rect 866 188 870 191
rect 878 181 881 468
rect 902 462 905 478
rect 910 392 913 518
rect 950 472 953 548
rect 982 502 985 548
rect 1014 542 1017 738
rect 1046 722 1049 748
rect 1062 742 1065 748
rect 1086 722 1089 758
rect 1118 742 1121 748
rect 1138 748 1142 751
rect 1102 732 1105 738
rect 1022 572 1025 718
rect 1030 652 1033 658
rect 1038 622 1041 658
rect 1022 542 1025 548
rect 990 482 993 488
rect 1010 468 1014 471
rect 926 442 929 458
rect 982 452 985 458
rect 926 352 929 428
rect 886 342 889 348
rect 918 312 921 348
rect 890 268 894 271
rect 926 262 929 338
rect 950 292 953 308
rect 942 262 945 278
rect 918 251 921 258
rect 934 252 937 258
rect 918 248 929 251
rect 870 178 881 181
rect 838 152 841 158
rect 662 142 665 147
rect 646 82 649 138
rect 646 72 649 78
rect 654 62 657 108
rect 766 102 769 148
rect 814 92 817 98
rect 802 88 806 91
rect 662 62 665 88
rect 710 82 713 88
rect 726 72 729 78
rect 870 72 873 178
rect 878 132 881 168
rect 914 158 918 161
rect 926 152 929 248
rect 938 168 942 171
rect 934 152 937 158
rect 958 152 961 358
rect 974 342 977 348
rect 966 192 969 338
rect 990 292 993 468
rect 1030 462 1033 608
rect 1046 582 1049 718
rect 1056 703 1058 707
rect 1062 703 1065 707
rect 1069 703 1072 707
rect 1062 662 1065 668
rect 1070 662 1073 688
rect 1110 662 1113 668
rect 1098 658 1102 661
rect 1078 592 1081 638
rect 1102 552 1105 558
rect 1110 552 1113 648
rect 1126 642 1129 668
rect 1134 662 1137 698
rect 1142 662 1145 668
rect 1118 562 1121 618
rect 1090 548 1094 551
rect 1122 548 1126 551
rect 1038 502 1041 528
rect 1038 492 1041 498
rect 1046 362 1049 538
rect 1056 503 1058 507
rect 1062 503 1065 507
rect 1069 503 1072 507
rect 1094 462 1097 508
rect 1102 442 1105 468
rect 1118 452 1121 548
rect 1134 542 1137 568
rect 1150 552 1153 898
rect 1166 752 1169 1138
rect 1174 1092 1177 1108
rect 1230 1072 1233 1168
rect 1246 1162 1249 1168
rect 1254 1142 1257 1308
rect 1278 1282 1281 1318
rect 1278 1272 1281 1278
rect 1286 1252 1289 1338
rect 1294 1262 1297 1308
rect 1302 1292 1305 1548
rect 1310 1542 1313 1548
rect 1318 1482 1321 1538
rect 1334 1532 1337 1538
rect 1366 1522 1369 1548
rect 1366 1492 1369 1518
rect 1382 1502 1385 1658
rect 1414 1622 1417 1668
rect 1422 1662 1425 1768
rect 1486 1752 1489 1758
rect 1474 1748 1478 1751
rect 1498 1748 1502 1751
rect 1602 1748 1606 1751
rect 1450 1738 1454 1741
rect 1430 1672 1433 1678
rect 1398 1492 1401 1598
rect 1430 1592 1433 1648
rect 1418 1568 1422 1571
rect 1422 1552 1425 1558
rect 1438 1542 1441 1658
rect 1446 1652 1449 1668
rect 1462 1662 1465 1698
rect 1446 1572 1449 1628
rect 1470 1572 1473 1748
rect 1486 1742 1489 1748
rect 1526 1742 1529 1748
rect 1502 1732 1505 1738
rect 1522 1728 1526 1731
rect 1478 1692 1481 1728
rect 1494 1672 1497 1678
rect 1526 1672 1529 1688
rect 1542 1672 1545 1738
rect 1590 1722 1593 1728
rect 1502 1662 1505 1668
rect 1582 1662 1585 1698
rect 1482 1658 1486 1661
rect 1562 1658 1566 1661
rect 1478 1642 1481 1648
rect 1518 1622 1521 1658
rect 1446 1542 1449 1568
rect 1466 1558 1470 1561
rect 1454 1551 1457 1558
rect 1454 1548 1465 1551
rect 1462 1542 1465 1548
rect 1486 1541 1489 1568
rect 1494 1552 1497 1558
rect 1502 1552 1505 1558
rect 1518 1542 1521 1618
rect 1486 1538 1494 1541
rect 1438 1532 1441 1538
rect 1334 1472 1337 1488
rect 1322 1468 1326 1471
rect 1346 1468 1350 1471
rect 1354 1458 1358 1461
rect 1350 1452 1353 1458
rect 1318 1441 1321 1448
rect 1310 1438 1321 1441
rect 1310 1292 1313 1438
rect 1318 1392 1321 1398
rect 1342 1392 1345 1418
rect 1358 1352 1361 1408
rect 1374 1392 1377 1458
rect 1382 1412 1385 1458
rect 1390 1392 1393 1438
rect 1398 1382 1401 1418
rect 1406 1372 1409 1468
rect 1414 1392 1417 1518
rect 1426 1458 1430 1461
rect 1430 1452 1433 1458
rect 1426 1438 1430 1441
rect 1430 1422 1433 1428
rect 1438 1392 1441 1508
rect 1454 1462 1457 1468
rect 1446 1452 1449 1458
rect 1366 1342 1369 1348
rect 1382 1342 1385 1358
rect 1406 1342 1409 1368
rect 1362 1338 1366 1341
rect 1398 1332 1401 1338
rect 1430 1332 1433 1358
rect 1446 1352 1449 1448
rect 1454 1402 1457 1418
rect 1462 1392 1465 1478
rect 1478 1452 1481 1478
rect 1486 1452 1489 1458
rect 1494 1452 1497 1508
rect 1474 1448 1478 1451
rect 1454 1342 1457 1368
rect 1470 1352 1473 1358
rect 1478 1352 1481 1388
rect 1486 1362 1489 1418
rect 1494 1412 1497 1448
rect 1510 1442 1513 1458
rect 1502 1352 1505 1388
rect 1510 1372 1513 1438
rect 1518 1422 1521 1538
rect 1526 1492 1529 1648
rect 1534 1632 1537 1658
rect 1542 1652 1545 1658
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1573 1603 1576 1607
rect 1546 1578 1550 1581
rect 1526 1342 1529 1418
rect 1534 1392 1537 1508
rect 1574 1492 1577 1568
rect 1582 1512 1585 1658
rect 1590 1592 1593 1718
rect 1610 1688 1614 1691
rect 1646 1662 1649 1768
rect 1678 1742 1681 1748
rect 1686 1662 1689 1668
rect 1598 1652 1601 1658
rect 1622 1632 1625 1658
rect 1630 1602 1633 1658
rect 1638 1652 1641 1658
rect 1658 1628 1662 1631
rect 1642 1558 1646 1561
rect 1602 1547 1606 1550
rect 1654 1542 1657 1578
rect 1666 1548 1670 1551
rect 1598 1492 1601 1518
rect 1622 1482 1625 1538
rect 1646 1492 1649 1528
rect 1542 1472 1545 1478
rect 1670 1472 1673 1538
rect 1678 1492 1681 1658
rect 1694 1652 1697 1658
rect 1686 1552 1689 1558
rect 1694 1542 1697 1608
rect 1702 1541 1705 1858
rect 1710 1752 1713 1768
rect 1718 1752 1721 1828
rect 1758 1822 1761 1858
rect 1710 1692 1713 1738
rect 1718 1692 1721 1748
rect 1734 1661 1737 1818
rect 1766 1812 1769 1858
rect 1758 1742 1761 1748
rect 1750 1722 1753 1728
rect 1750 1662 1753 1688
rect 1774 1662 1777 1728
rect 1782 1692 1785 1818
rect 1798 1702 1801 1858
rect 1814 1792 1817 1808
rect 1822 1732 1825 1818
rect 1838 1762 1841 1858
rect 1846 1802 1849 1948
rect 1854 1902 1857 1938
rect 1854 1862 1857 1868
rect 1854 1752 1857 1788
rect 1862 1762 1865 1948
rect 1870 1892 1873 1898
rect 1886 1862 1889 2008
rect 1950 1992 1953 2058
rect 1974 2052 1977 2108
rect 2030 2092 2033 2148
rect 2038 2142 2041 2268
rect 1994 2068 1998 2071
rect 2046 2062 2049 2288
rect 2102 2282 2105 2288
rect 2070 2263 2073 2278
rect 2142 2272 2145 2338
rect 2206 2332 2209 2338
rect 2150 2282 2153 2288
rect 2206 2272 2209 2328
rect 2238 2302 2241 2318
rect 2146 2268 2153 2271
rect 2086 2262 2089 2268
rect 2138 2258 2142 2261
rect 2126 2151 2129 2158
rect 2150 2152 2153 2268
rect 2158 2262 2161 2268
rect 2054 2082 2057 2128
rect 2086 2122 2089 2138
rect 2054 2062 2057 2078
rect 2018 2058 2022 2061
rect 1974 2002 1977 2048
rect 1990 2032 1993 2058
rect 2006 2052 2009 2058
rect 1978 1948 1982 1951
rect 1902 1942 1905 1948
rect 1918 1862 1921 1928
rect 1886 1852 1889 1858
rect 1874 1748 1878 1751
rect 1794 1688 1798 1691
rect 1814 1681 1817 1718
rect 1822 1712 1825 1718
rect 1830 1692 1833 1748
rect 1806 1678 1817 1681
rect 1846 1682 1849 1708
rect 1730 1658 1737 1661
rect 1718 1652 1721 1658
rect 1742 1652 1745 1658
rect 1766 1652 1769 1658
rect 1710 1592 1713 1648
rect 1762 1588 1766 1591
rect 1774 1572 1777 1648
rect 1798 1592 1801 1658
rect 1806 1652 1809 1678
rect 1878 1672 1881 1678
rect 1826 1668 1830 1671
rect 1862 1662 1865 1668
rect 1870 1662 1873 1668
rect 1814 1632 1817 1658
rect 1814 1612 1817 1628
rect 1714 1548 1718 1551
rect 1726 1542 1729 1558
rect 1790 1552 1793 1578
rect 1822 1552 1825 1608
rect 1862 1572 1865 1658
rect 1886 1602 1889 1848
rect 1894 1812 1897 1858
rect 1918 1752 1921 1758
rect 1926 1752 1929 1898
rect 1966 1862 1969 1928
rect 1990 1862 1993 1998
rect 2006 1942 2009 1948
rect 2022 1932 2025 2018
rect 2070 1952 2073 2118
rect 2080 2103 2082 2107
rect 2086 2103 2089 2107
rect 2093 2103 2096 2107
rect 2110 2092 2113 2098
rect 2134 2082 2137 2118
rect 2118 2062 2121 2078
rect 2086 1951 2089 1958
rect 2070 1942 2073 1948
rect 2026 1918 2030 1921
rect 2006 1872 2009 1878
rect 2014 1862 2017 1918
rect 2080 1903 2082 1907
rect 2086 1903 2089 1907
rect 2093 1903 2096 1907
rect 2038 1862 2041 1868
rect 2062 1862 2065 1878
rect 2102 1862 2105 1988
rect 2118 1972 2121 2058
rect 2126 2052 2129 2058
rect 2118 1922 2121 1938
rect 2134 1881 2137 2078
rect 2158 2062 2161 2258
rect 2166 2222 2169 2258
rect 2206 2182 2209 2268
rect 2214 2262 2217 2298
rect 2262 2292 2265 2338
rect 2270 2332 2273 2338
rect 2302 2272 2305 2398
rect 2434 2368 2438 2371
rect 2334 2322 2337 2338
rect 2318 2262 2321 2278
rect 2362 2268 2366 2271
rect 2342 2262 2345 2268
rect 2350 2252 2353 2258
rect 2366 2252 2369 2258
rect 2238 2192 2241 2218
rect 2186 2168 2190 2171
rect 2254 2152 2257 2188
rect 2262 2172 2265 2218
rect 2278 2192 2281 2218
rect 2314 2148 2318 2151
rect 2174 2111 2177 2148
rect 2198 2142 2201 2148
rect 2166 2108 2177 2111
rect 2166 2092 2169 2108
rect 2174 2062 2177 2068
rect 2182 2062 2185 2068
rect 2198 2062 2201 2108
rect 2214 2082 2217 2118
rect 2214 2062 2217 2078
rect 2146 2058 2150 2061
rect 2190 2012 2193 2058
rect 2146 1958 2150 1961
rect 2174 1952 2177 1958
rect 2150 1942 2153 1948
rect 2182 1942 2185 1968
rect 2206 1951 2209 2018
rect 2202 1948 2209 1951
rect 2222 1952 2225 2138
rect 2234 2068 2238 2071
rect 2234 2058 2238 2061
rect 2246 2032 2249 2058
rect 2254 1982 2257 2148
rect 2326 2142 2329 2218
rect 2342 2142 2345 2148
rect 2358 2122 2361 2128
rect 2266 2118 2270 2121
rect 2366 2111 2369 2248
rect 2374 2172 2377 2338
rect 2382 2292 2385 2348
rect 2406 2272 2409 2278
rect 2414 2272 2417 2368
rect 2482 2348 2486 2351
rect 2430 2282 2433 2318
rect 2438 2292 2441 2348
rect 2534 2342 2537 2358
rect 2518 2332 2521 2338
rect 2414 2262 2417 2268
rect 2454 2252 2457 2258
rect 2386 2248 2390 2251
rect 2434 2248 2438 2251
rect 2390 2132 2393 2138
rect 2414 2122 2417 2148
rect 2438 2142 2441 2158
rect 2358 2108 2369 2111
rect 2262 2062 2265 2088
rect 2286 2082 2289 2098
rect 2298 2088 2302 2091
rect 2286 2062 2289 2078
rect 2298 2068 2302 2071
rect 2274 2058 2278 2061
rect 2346 2058 2350 2061
rect 2262 2052 2265 2058
rect 2238 1952 2241 1978
rect 2190 1942 2193 1948
rect 2206 1901 2209 1918
rect 2126 1878 2137 1881
rect 2198 1898 2209 1901
rect 2126 1862 2129 1878
rect 2134 1862 2137 1868
rect 2150 1862 2153 1868
rect 2178 1858 2182 1861
rect 1958 1812 1961 1818
rect 1974 1792 1977 1858
rect 1942 1762 1945 1768
rect 1950 1752 1953 1768
rect 1990 1751 1993 1758
rect 1902 1742 1905 1748
rect 1926 1701 1929 1748
rect 1974 1742 1977 1748
rect 1926 1698 1937 1701
rect 1894 1672 1897 1688
rect 1926 1672 1929 1688
rect 1898 1658 1902 1661
rect 1898 1648 1910 1651
rect 1934 1632 1937 1698
rect 1990 1692 1993 1728
rect 2022 1712 2025 1858
rect 2030 1852 2033 1858
rect 2094 1822 2097 1858
rect 2054 1782 2057 1818
rect 2066 1768 2070 1771
rect 2070 1732 2073 1758
rect 2094 1732 2097 1758
rect 2110 1752 2113 1778
rect 2122 1738 2126 1741
rect 2134 1741 2137 1808
rect 2142 1792 2145 1858
rect 2146 1748 2150 1751
rect 2166 1742 2169 1818
rect 2134 1738 2142 1741
rect 2110 1732 2113 1738
rect 2182 1732 2185 1738
rect 2138 1728 2142 1731
rect 2070 1722 2073 1728
rect 2058 1718 2062 1721
rect 2080 1703 2082 1707
rect 2086 1703 2089 1707
rect 2093 1703 2096 1707
rect 1962 1688 1966 1691
rect 2054 1682 2057 1688
rect 1966 1672 1969 1678
rect 2102 1672 2105 1718
rect 2166 1702 2169 1718
rect 2134 1672 2137 1688
rect 2150 1672 2153 1678
rect 2034 1668 2038 1671
rect 1954 1658 1958 1661
rect 1942 1652 1945 1658
rect 1954 1648 1958 1651
rect 1966 1632 1969 1668
rect 1922 1588 1926 1591
rect 1934 1582 1937 1628
rect 1990 1622 1993 1668
rect 1998 1662 2001 1668
rect 2118 1663 2121 1668
rect 2018 1658 2022 1661
rect 2166 1662 2169 1668
rect 1998 1642 2001 1658
rect 2006 1652 2009 1658
rect 1934 1552 1937 1578
rect 1950 1562 1953 1568
rect 1762 1548 1766 1551
rect 1866 1548 1870 1551
rect 1946 1548 1950 1551
rect 1702 1538 1713 1541
rect 1746 1538 1750 1541
rect 1694 1492 1697 1528
rect 1702 1522 1705 1528
rect 1682 1488 1686 1491
rect 1586 1468 1590 1471
rect 1674 1468 1678 1471
rect 1594 1448 1598 1451
rect 1542 1342 1545 1418
rect 1550 1402 1553 1418
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1573 1403 1576 1407
rect 1558 1382 1561 1388
rect 1550 1371 1553 1378
rect 1550 1368 1561 1371
rect 1550 1352 1553 1358
rect 1498 1338 1502 1341
rect 1434 1318 1438 1321
rect 1326 1272 1329 1278
rect 1294 1252 1297 1258
rect 1282 1248 1286 1251
rect 1302 1242 1305 1268
rect 1306 1238 1310 1241
rect 1262 1152 1265 1178
rect 1270 1158 1278 1161
rect 1246 1138 1254 1141
rect 1246 1092 1249 1138
rect 1246 1062 1249 1088
rect 1262 1071 1265 1148
rect 1270 1092 1273 1158
rect 1294 1152 1297 1158
rect 1282 1148 1286 1151
rect 1282 1138 1286 1141
rect 1286 1072 1289 1108
rect 1262 1068 1273 1071
rect 1262 1052 1265 1058
rect 1270 1052 1273 1068
rect 1174 1002 1177 1018
rect 1246 972 1249 1008
rect 1242 968 1246 971
rect 1182 942 1185 947
rect 1198 932 1201 938
rect 1254 932 1257 1018
rect 1262 972 1265 1048
rect 1270 952 1273 1038
rect 1190 882 1193 918
rect 1198 912 1201 928
rect 1198 862 1201 908
rect 1210 868 1214 871
rect 1238 862 1241 888
rect 1278 882 1281 998
rect 1286 982 1289 1068
rect 1294 992 1297 1058
rect 1302 1012 1305 1058
rect 1310 1012 1313 1218
rect 1322 1158 1326 1161
rect 1318 1152 1321 1158
rect 1326 1141 1329 1148
rect 1322 1138 1329 1141
rect 1334 1142 1337 1188
rect 1342 1171 1345 1318
rect 1354 1258 1358 1261
rect 1366 1172 1369 1188
rect 1342 1168 1350 1171
rect 1370 1148 1374 1151
rect 1382 1102 1385 1138
rect 1326 1062 1329 1068
rect 1342 1062 1345 1068
rect 1382 1062 1385 1068
rect 1318 1052 1321 1058
rect 1350 1052 1353 1058
rect 1374 1042 1377 1058
rect 1286 952 1289 958
rect 1246 862 1249 868
rect 1286 862 1289 868
rect 1214 792 1217 858
rect 1294 852 1297 948
rect 1302 922 1305 948
rect 1270 752 1273 798
rect 1282 768 1286 771
rect 1190 721 1193 728
rect 1190 718 1198 721
rect 1174 662 1177 668
rect 1190 662 1193 718
rect 1246 692 1249 738
rect 1270 732 1273 738
rect 1294 721 1297 758
rect 1294 718 1305 721
rect 1302 692 1305 718
rect 1218 668 1222 671
rect 1258 668 1262 671
rect 1274 668 1278 671
rect 1158 658 1166 661
rect 1150 542 1153 548
rect 1130 528 1134 531
rect 1118 392 1121 438
rect 1102 352 1105 368
rect 974 152 977 288
rect 1014 272 1017 348
rect 1050 338 1054 341
rect 1030 332 1033 338
rect 1056 303 1058 307
rect 1062 303 1065 307
rect 1069 303 1072 307
rect 1078 272 1081 288
rect 910 72 913 98
rect 926 92 929 148
rect 934 112 937 148
rect 974 122 977 148
rect 982 122 985 258
rect 1006 182 1009 258
rect 1014 202 1017 268
rect 1046 262 1049 268
rect 1022 252 1025 258
rect 1042 248 1046 251
rect 1006 172 1009 178
rect 994 148 998 151
rect 958 72 961 88
rect 974 72 977 78
rect 690 68 694 71
rect 930 68 934 71
rect 742 63 745 68
rect 878 63 881 68
rect 1014 62 1017 68
rect 1022 62 1025 248
rect 1094 242 1097 348
rect 1142 292 1145 468
rect 1158 402 1161 658
rect 1182 652 1185 658
rect 1214 642 1217 658
rect 1230 632 1233 668
rect 1286 662 1289 678
rect 1294 672 1297 688
rect 1258 658 1262 661
rect 1298 658 1302 661
rect 1246 642 1249 648
rect 1262 632 1265 638
rect 1310 612 1313 1008
rect 1318 992 1321 1038
rect 1326 952 1329 978
rect 1342 952 1345 968
rect 1374 952 1377 978
rect 1390 962 1393 1318
rect 1410 1288 1414 1291
rect 1422 1282 1425 1318
rect 1446 1312 1449 1338
rect 1478 1332 1481 1338
rect 1498 1328 1502 1331
rect 1414 1142 1417 1268
rect 1422 1262 1425 1278
rect 1434 1258 1438 1261
rect 1446 1252 1449 1278
rect 1434 1168 1438 1171
rect 1446 1142 1449 1248
rect 1454 1152 1457 1278
rect 1462 1272 1465 1288
rect 1478 1262 1481 1288
rect 1518 1272 1521 1328
rect 1542 1282 1545 1338
rect 1550 1292 1553 1318
rect 1502 1262 1505 1268
rect 1558 1262 1561 1368
rect 1582 1362 1585 1448
rect 1598 1392 1601 1428
rect 1566 1332 1569 1338
rect 1574 1272 1577 1298
rect 1582 1292 1585 1358
rect 1606 1352 1609 1468
rect 1614 1462 1617 1468
rect 1630 1452 1633 1458
rect 1614 1422 1617 1438
rect 1622 1432 1625 1438
rect 1710 1432 1713 1538
rect 1750 1532 1753 1538
rect 1738 1528 1742 1531
rect 1734 1462 1737 1518
rect 1814 1502 1817 1548
rect 1642 1358 1646 1361
rect 1606 1332 1609 1338
rect 1618 1328 1622 1331
rect 1590 1292 1593 1308
rect 1578 1268 1582 1271
rect 1466 1258 1470 1261
rect 1470 1162 1473 1228
rect 1482 1188 1486 1191
rect 1494 1182 1497 1218
rect 1526 1192 1529 1258
rect 1538 1248 1542 1251
rect 1518 1152 1521 1168
rect 1490 1148 1494 1151
rect 1506 1148 1510 1151
rect 1398 1092 1401 1128
rect 1414 982 1417 1138
rect 1438 1132 1441 1138
rect 1438 1092 1441 1118
rect 1446 1072 1449 1118
rect 1430 1052 1433 1068
rect 1454 1061 1457 1148
rect 1466 1128 1470 1131
rect 1470 1072 1473 1128
rect 1502 1122 1505 1128
rect 1502 1082 1505 1118
rect 1486 1062 1489 1078
rect 1450 1058 1465 1061
rect 1450 1048 1454 1051
rect 1454 1002 1457 1028
rect 1394 948 1398 951
rect 1382 932 1385 938
rect 1398 932 1401 938
rect 1358 892 1361 918
rect 1382 902 1385 928
rect 1350 872 1353 878
rect 1358 862 1361 888
rect 1370 868 1374 871
rect 1414 862 1417 958
rect 1434 948 1438 951
rect 1430 912 1433 928
rect 1446 862 1449 878
rect 1454 862 1457 998
rect 1462 882 1465 1058
rect 1490 1018 1494 1021
rect 1502 972 1505 1058
rect 1510 1002 1513 1148
rect 1526 1092 1529 1108
rect 1542 1062 1545 1178
rect 1494 951 1497 968
rect 1510 962 1513 968
rect 1542 962 1545 1008
rect 1550 992 1553 1258
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1573 1203 1576 1207
rect 1558 1142 1561 1168
rect 1570 1158 1574 1161
rect 1558 1052 1561 1058
rect 1574 1022 1577 1058
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1573 1003 1576 1007
rect 1582 952 1585 1258
rect 1598 1242 1601 1318
rect 1606 1312 1609 1328
rect 1626 1288 1630 1291
rect 1638 1262 1641 1348
rect 1654 1342 1657 1388
rect 1662 1352 1665 1418
rect 1686 1392 1689 1408
rect 1678 1352 1681 1388
rect 1662 1342 1665 1348
rect 1666 1328 1670 1331
rect 1646 1302 1649 1328
rect 1670 1312 1673 1318
rect 1718 1292 1721 1338
rect 1654 1282 1657 1288
rect 1662 1268 1670 1271
rect 1646 1262 1649 1268
rect 1654 1262 1657 1268
rect 1606 1222 1609 1228
rect 1626 1168 1630 1171
rect 1614 1152 1617 1158
rect 1602 1138 1606 1141
rect 1622 1112 1625 1138
rect 1610 1068 1614 1071
rect 1602 1058 1606 1061
rect 1590 1042 1593 1058
rect 1602 958 1606 961
rect 1494 948 1502 951
rect 1562 948 1566 951
rect 1502 932 1505 948
rect 1394 858 1398 861
rect 1338 748 1342 751
rect 1330 728 1334 731
rect 1318 672 1321 688
rect 1366 662 1369 668
rect 1374 662 1377 668
rect 1382 662 1385 858
rect 1390 792 1393 838
rect 1414 822 1417 858
rect 1422 842 1425 858
rect 1414 812 1417 818
rect 1390 672 1393 758
rect 1414 752 1417 758
rect 1422 752 1425 758
rect 1430 752 1433 818
rect 1398 692 1401 748
rect 1406 682 1409 718
rect 1422 702 1425 728
rect 1422 692 1425 698
rect 1338 658 1342 661
rect 1366 592 1369 608
rect 1390 602 1393 668
rect 1414 592 1417 648
rect 1282 578 1286 581
rect 1302 562 1305 568
rect 1326 552 1329 558
rect 1234 548 1238 551
rect 1314 548 1318 551
rect 1174 542 1177 548
rect 1166 512 1169 518
rect 1174 462 1177 468
rect 1182 372 1185 548
rect 1198 521 1201 538
rect 1190 518 1201 521
rect 1190 392 1193 518
rect 1190 382 1193 388
rect 1174 342 1177 358
rect 1206 292 1209 508
rect 1254 472 1257 498
rect 1318 482 1321 488
rect 1286 472 1289 478
rect 1230 462 1233 468
rect 1234 448 1238 451
rect 1246 442 1249 458
rect 1262 452 1265 468
rect 1282 458 1286 461
rect 1262 422 1265 438
rect 1226 418 1230 421
rect 1166 272 1169 278
rect 1182 262 1185 268
rect 1230 262 1233 388
rect 1262 352 1265 418
rect 1278 392 1281 448
rect 1318 392 1321 438
rect 1326 432 1329 458
rect 1334 442 1337 538
rect 1342 361 1345 568
rect 1382 552 1385 558
rect 1390 552 1393 568
rect 1398 552 1401 578
rect 1430 552 1433 588
rect 1438 572 1441 858
rect 1446 792 1449 838
rect 1462 782 1465 868
rect 1470 862 1473 868
rect 1478 792 1481 918
rect 1486 892 1489 928
rect 1510 892 1513 938
rect 1518 932 1521 948
rect 1526 942 1529 948
rect 1558 942 1561 948
rect 1574 942 1577 948
rect 1494 872 1497 878
rect 1454 592 1457 748
rect 1478 742 1481 788
rect 1502 782 1505 818
rect 1518 752 1521 928
rect 1598 902 1601 958
rect 1622 942 1625 1108
rect 1646 1082 1649 1258
rect 1662 1092 1665 1268
rect 1674 1258 1678 1261
rect 1686 1252 1689 1258
rect 1678 1142 1681 1148
rect 1694 1111 1697 1278
rect 1702 1252 1705 1288
rect 1710 1272 1713 1278
rect 1706 1248 1710 1251
rect 1710 1142 1713 1228
rect 1694 1108 1705 1111
rect 1630 1072 1633 1078
rect 1678 1072 1681 1078
rect 1638 1062 1641 1068
rect 1646 1062 1649 1068
rect 1666 1058 1670 1061
rect 1630 1052 1633 1058
rect 1686 1052 1689 1058
rect 1694 1052 1697 1068
rect 1702 1062 1705 1108
rect 1666 1048 1670 1051
rect 1702 1012 1705 1058
rect 1714 1038 1718 1041
rect 1726 962 1729 1438
rect 1734 1262 1737 1368
rect 1742 1342 1745 1468
rect 1786 1458 1790 1461
rect 1774 1432 1777 1458
rect 1822 1452 1825 1548
rect 1958 1542 1961 1578
rect 2014 1572 2017 1588
rect 2022 1582 2025 1618
rect 2054 1562 2057 1618
rect 2006 1552 2009 1558
rect 2014 1552 2017 1558
rect 2078 1552 2081 1558
rect 2110 1552 2113 1638
rect 2022 1548 2030 1551
rect 2066 1548 2070 1551
rect 1870 1522 1873 1538
rect 1870 1492 1873 1498
rect 1830 1482 1833 1488
rect 1918 1482 1921 1518
rect 1926 1512 1929 1538
rect 1926 1482 1929 1508
rect 1794 1418 1798 1421
rect 1750 1351 1753 1418
rect 1830 1412 1833 1478
rect 1918 1472 1921 1478
rect 1854 1462 1857 1468
rect 1782 1352 1785 1358
rect 1790 1352 1793 1398
rect 1758 1292 1761 1308
rect 1766 1242 1769 1338
rect 1806 1312 1809 1318
rect 1806 1272 1809 1278
rect 1798 1262 1801 1268
rect 1782 1252 1785 1258
rect 1790 1251 1793 1258
rect 1806 1251 1809 1258
rect 1790 1248 1809 1251
rect 1734 1101 1737 1118
rect 1734 1098 1742 1101
rect 1758 972 1761 1218
rect 1774 1063 1777 1088
rect 1790 1082 1793 1138
rect 1790 1072 1793 1078
rect 1806 1042 1809 1068
rect 1814 1051 1817 1318
rect 1822 1292 1825 1378
rect 1838 1372 1841 1458
rect 1838 1332 1841 1358
rect 1870 1312 1873 1347
rect 1902 1312 1905 1348
rect 1918 1311 1921 1468
rect 1930 1459 1934 1462
rect 1934 1372 1937 1448
rect 1966 1442 1969 1548
rect 1982 1462 1985 1518
rect 1990 1502 1993 1538
rect 2014 1472 2017 1528
rect 1998 1462 2001 1468
rect 2022 1462 2025 1548
rect 2038 1532 2041 1538
rect 2046 1492 2049 1548
rect 2086 1532 2089 1548
rect 2118 1542 2121 1638
rect 2134 1542 2137 1628
rect 2150 1552 2153 1568
rect 2158 1552 2161 1558
rect 2190 1552 2193 1788
rect 2198 1752 2201 1898
rect 2214 1792 2217 1858
rect 2206 1752 2209 1758
rect 2198 1662 2201 1718
rect 2222 1692 2225 1868
rect 2246 1862 2249 1968
rect 2270 1952 2273 1998
rect 2302 1962 2305 1998
rect 2302 1942 2305 1948
rect 2318 1942 2321 1968
rect 2254 1912 2257 1918
rect 2238 1772 2241 1858
rect 2258 1748 2262 1751
rect 2230 1742 2233 1748
rect 2206 1662 2209 1668
rect 2142 1532 2145 1548
rect 2198 1541 2201 1658
rect 2222 1622 2225 1658
rect 2238 1651 2241 1748
rect 2246 1742 2249 1748
rect 2270 1722 2273 1938
rect 2318 1872 2321 1938
rect 2294 1862 2297 1868
rect 2326 1861 2329 1898
rect 2334 1872 2337 1878
rect 2322 1858 2329 1861
rect 2334 1852 2337 1858
rect 2278 1752 2281 1818
rect 2246 1662 2249 1668
rect 2238 1648 2249 1651
rect 2230 1642 2233 1648
rect 2214 1592 2217 1618
rect 2206 1552 2209 1568
rect 2238 1552 2241 1558
rect 2246 1552 2249 1648
rect 2254 1562 2257 1658
rect 2262 1632 2265 1718
rect 2270 1632 2273 1658
rect 2262 1592 2265 1618
rect 2278 1572 2281 1618
rect 2198 1538 2209 1541
rect 2170 1528 2174 1531
rect 2080 1503 2082 1507
rect 2086 1503 2089 1507
rect 2093 1503 2096 1507
rect 2070 1472 2073 1478
rect 2050 1468 2054 1471
rect 2038 1462 2041 1468
rect 1974 1452 1977 1458
rect 2006 1452 2009 1458
rect 1982 1412 1985 1418
rect 1950 1392 1953 1398
rect 1934 1362 1937 1368
rect 1942 1342 1945 1358
rect 1966 1352 1969 1408
rect 1998 1352 2001 1358
rect 2022 1352 2025 1458
rect 2030 1452 2033 1458
rect 2038 1452 2041 1458
rect 2046 1452 2049 1458
rect 2062 1422 2065 1458
rect 2094 1442 2097 1448
rect 2062 1412 2065 1418
rect 2074 1388 2078 1391
rect 2102 1372 2105 1458
rect 2110 1372 2113 1398
rect 2118 1392 2121 1408
rect 2066 1358 2070 1361
rect 2102 1352 2105 1368
rect 2126 1362 2129 1518
rect 2206 1492 2209 1538
rect 2174 1472 2177 1478
rect 2230 1472 2233 1548
rect 2246 1522 2249 1548
rect 2254 1512 2257 1548
rect 2150 1462 2153 1468
rect 2190 1452 2193 1458
rect 2190 1412 2193 1448
rect 2162 1358 2169 1361
rect 2166 1352 2169 1358
rect 2174 1352 2177 1358
rect 2206 1352 2209 1358
rect 2010 1348 2014 1351
rect 2050 1348 2054 1351
rect 1942 1332 1945 1338
rect 1978 1328 1982 1331
rect 1910 1308 1921 1311
rect 1822 1282 1825 1288
rect 1910 1272 1913 1308
rect 1942 1282 1945 1288
rect 1822 1212 1825 1218
rect 1830 1142 1833 1268
rect 1838 1262 1841 1268
rect 1846 1252 1849 1268
rect 1910 1262 1913 1268
rect 1854 1222 1857 1238
rect 1854 1192 1857 1218
rect 1878 1212 1881 1259
rect 1954 1258 1958 1261
rect 1990 1242 1993 1348
rect 2126 1342 2129 1348
rect 2142 1342 2145 1348
rect 2198 1342 2201 1348
rect 2026 1338 2030 1341
rect 2082 1338 2086 1341
rect 2014 1332 2017 1338
rect 2046 1332 2049 1338
rect 2230 1332 2233 1458
rect 2238 1392 2241 1508
rect 2254 1462 2257 1468
rect 2262 1462 2265 1518
rect 2270 1472 2273 1508
rect 2278 1502 2281 1548
rect 2262 1432 2265 1458
rect 2286 1452 2289 1838
rect 2302 1792 2305 1818
rect 2342 1812 2345 1858
rect 2294 1662 2297 1778
rect 2314 1758 2318 1761
rect 2322 1758 2326 1761
rect 2334 1752 2337 1768
rect 2358 1762 2361 2108
rect 2462 2102 2465 2268
rect 2478 2162 2481 2218
rect 2466 2098 2473 2101
rect 2382 2072 2385 2078
rect 2406 2062 2409 2098
rect 2438 2062 2441 2068
rect 2398 2052 2401 2058
rect 2462 1992 2465 2018
rect 2378 1948 2382 1951
rect 2458 1948 2462 1951
rect 2406 1922 2409 1938
rect 2422 1921 2425 1948
rect 2430 1942 2433 1948
rect 2470 1942 2473 2098
rect 2478 1992 2481 2147
rect 2494 1962 2497 2278
rect 2502 1972 2505 2328
rect 2534 2282 2537 2318
rect 2538 2268 2542 2271
rect 2538 2248 2542 2251
rect 2550 2231 2553 2338
rect 2558 2322 2561 2338
rect 2614 2272 2617 2318
rect 2622 2292 2625 2328
rect 2542 2228 2553 2231
rect 2542 2192 2545 2228
rect 2558 2222 2561 2268
rect 2550 2172 2553 2218
rect 2566 2211 2569 2268
rect 2558 2208 2569 2211
rect 2526 2112 2529 2128
rect 2558 2072 2561 2208
rect 2586 2148 2590 2151
rect 2590 2112 2593 2138
rect 2614 2092 2617 2108
rect 2514 2058 2518 2061
rect 2542 2021 2545 2068
rect 2534 2018 2545 2021
rect 2534 1972 2537 2018
rect 2622 1992 2625 2148
rect 2478 1952 2481 1958
rect 2498 1948 2502 1951
rect 2574 1942 2577 1948
rect 2458 1938 2462 1941
rect 2414 1918 2425 1921
rect 2366 1862 2369 1868
rect 2382 1862 2385 1868
rect 2374 1852 2377 1858
rect 2398 1852 2401 1858
rect 2414 1832 2417 1918
rect 2430 1912 2433 1928
rect 2430 1872 2433 1908
rect 2510 1902 2513 1928
rect 2438 1872 2441 1888
rect 2518 1872 2521 1878
rect 2534 1872 2537 1918
rect 2598 1872 2601 1938
rect 2614 1932 2617 1938
rect 2614 1892 2617 1918
rect 2434 1858 2438 1861
rect 2494 1852 2497 1858
rect 2426 1848 2430 1851
rect 2534 1841 2537 1868
rect 2526 1838 2537 1841
rect 2606 1842 2609 1848
rect 2622 1842 2625 1948
rect 2638 1872 2641 2118
rect 2646 1922 2649 1958
rect 2374 1772 2377 1808
rect 2306 1748 2310 1751
rect 2314 1738 2318 1741
rect 2342 1722 2345 1748
rect 2350 1732 2353 1738
rect 2358 1732 2361 1758
rect 2310 1662 2313 1688
rect 2318 1662 2321 1668
rect 2342 1662 2345 1698
rect 2294 1532 2297 1638
rect 2302 1602 2305 1658
rect 2350 1652 2353 1658
rect 2358 1652 2361 1718
rect 2366 1672 2369 1748
rect 2374 1742 2377 1768
rect 2434 1748 2438 1751
rect 2374 1662 2377 1718
rect 2438 1712 2441 1738
rect 2446 1722 2449 1728
rect 2406 1682 2409 1688
rect 2382 1672 2385 1678
rect 2426 1668 2430 1671
rect 2390 1662 2393 1668
rect 2438 1662 2441 1708
rect 2446 1702 2449 1708
rect 2446 1672 2449 1698
rect 2462 1692 2465 1758
rect 2478 1752 2481 1758
rect 2486 1752 2489 1758
rect 2494 1752 2497 1798
rect 2498 1738 2502 1741
rect 2510 1712 2513 1718
rect 2470 1682 2473 1688
rect 2526 1672 2529 1838
rect 2562 1748 2566 1751
rect 2590 1742 2593 1818
rect 2638 1782 2641 1868
rect 2382 1658 2390 1661
rect 2426 1658 2430 1661
rect 2522 1658 2526 1661
rect 2302 1552 2305 1558
rect 2310 1542 2313 1578
rect 2350 1551 2353 1558
rect 2318 1542 2321 1548
rect 2286 1442 2289 1448
rect 2294 1382 2297 1528
rect 2334 1482 2337 1538
rect 2334 1472 2337 1478
rect 2314 1468 2318 1471
rect 2302 1351 2305 1458
rect 2310 1442 2313 1458
rect 2334 1352 2337 1468
rect 2358 1462 2361 1508
rect 2318 1342 2321 1348
rect 2334 1342 2337 1348
rect 2026 1328 2030 1331
rect 2186 1328 2190 1331
rect 2218 1328 2222 1331
rect 1998 1272 2001 1308
rect 2010 1268 2014 1271
rect 1990 1192 1993 1208
rect 1918 1152 1921 1158
rect 1870 1122 1873 1138
rect 1950 1132 1953 1147
rect 1878 1122 1881 1128
rect 1830 1082 1833 1088
rect 1870 1082 1873 1118
rect 1886 1082 1889 1118
rect 1990 1112 1993 1118
rect 1998 1072 2001 1268
rect 2022 1262 2025 1278
rect 2014 1142 2017 1148
rect 2022 1142 2025 1148
rect 1842 1058 1846 1061
rect 1822 1052 1825 1058
rect 1814 1048 1822 1051
rect 1782 992 1785 1018
rect 1806 981 1809 1038
rect 1830 992 1833 1048
rect 1798 978 1809 981
rect 1750 952 1753 958
rect 1798 952 1801 978
rect 1806 952 1809 958
rect 1650 948 1654 951
rect 1754 948 1761 951
rect 1726 942 1729 948
rect 1638 922 1641 928
rect 1590 872 1593 888
rect 1574 863 1577 868
rect 1510 692 1513 748
rect 1478 672 1481 678
rect 1486 662 1489 668
rect 1494 662 1497 668
rect 1350 452 1353 548
rect 1374 422 1377 548
rect 1422 532 1425 548
rect 1446 512 1449 548
rect 1390 472 1393 478
rect 1398 462 1401 488
rect 1430 452 1433 508
rect 1462 492 1465 658
rect 1510 652 1513 678
rect 1518 662 1521 668
rect 1526 652 1529 658
rect 1522 548 1526 551
rect 1470 522 1473 548
rect 1442 468 1446 471
rect 1438 452 1441 458
rect 1426 448 1430 451
rect 1382 442 1385 448
rect 1430 432 1433 438
rect 1398 422 1401 428
rect 1358 392 1361 418
rect 1334 358 1345 361
rect 1334 352 1337 358
rect 1430 352 1433 428
rect 1438 382 1441 448
rect 1446 402 1449 468
rect 1462 462 1465 488
rect 1454 422 1457 458
rect 1454 392 1457 418
rect 1470 352 1473 418
rect 1494 352 1497 538
rect 1510 482 1513 518
rect 1518 492 1521 528
rect 1510 392 1513 478
rect 1518 472 1521 488
rect 1534 452 1537 458
rect 1522 388 1526 391
rect 1326 348 1334 351
rect 1402 348 1406 351
rect 1242 338 1246 341
rect 1138 258 1142 261
rect 1046 192 1049 238
rect 1086 212 1089 218
rect 1062 192 1065 208
rect 1062 152 1065 188
rect 1086 152 1089 198
rect 1110 142 1113 148
rect 1118 142 1121 148
rect 1090 138 1094 141
rect 1134 132 1137 148
rect 1134 122 1137 128
rect 1046 92 1049 118
rect 1056 103 1058 107
rect 1062 103 1065 107
rect 1069 103 1072 107
rect 1046 62 1049 88
rect 1078 82 1081 118
rect 1142 72 1145 198
rect 1166 192 1169 258
rect 1190 252 1193 258
rect 1182 152 1185 178
rect 1198 152 1201 208
rect 1214 192 1217 258
rect 1238 242 1241 258
rect 1254 162 1257 348
rect 1286 282 1289 348
rect 1302 312 1305 348
rect 1270 262 1273 268
rect 1302 192 1305 308
rect 1326 182 1329 348
rect 1230 152 1233 158
rect 1290 148 1294 151
rect 1174 92 1177 148
rect 1222 102 1225 148
rect 1334 142 1337 338
rect 1342 332 1345 348
rect 1382 332 1385 348
rect 1422 342 1425 348
rect 1446 342 1449 348
rect 1534 332 1537 398
rect 1542 392 1545 858
rect 1606 852 1609 918
rect 1614 872 1617 878
rect 1638 862 1641 898
rect 1646 872 1649 938
rect 1678 892 1681 908
rect 1686 862 1689 928
rect 1734 872 1737 888
rect 1694 862 1697 868
rect 1750 862 1753 868
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1573 803 1576 807
rect 1590 792 1593 828
rect 1630 792 1633 808
rect 1638 792 1641 858
rect 1598 762 1601 778
rect 1582 742 1585 758
rect 1598 742 1601 758
rect 1614 722 1617 740
rect 1558 692 1561 718
rect 1578 678 1582 681
rect 1598 662 1601 708
rect 1606 672 1609 688
rect 1622 672 1625 678
rect 1630 672 1633 768
rect 1638 762 1641 768
rect 1550 632 1553 658
rect 1558 642 1561 658
rect 1582 652 1585 658
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1573 603 1576 607
rect 1582 602 1585 648
rect 1614 622 1617 668
rect 1638 662 1641 738
rect 1646 692 1649 858
rect 1654 792 1657 818
rect 1654 752 1657 758
rect 1702 752 1705 758
rect 1710 752 1713 798
rect 1718 752 1721 778
rect 1654 738 1662 741
rect 1654 692 1657 738
rect 1670 732 1673 748
rect 1682 738 1686 741
rect 1726 692 1729 748
rect 1734 712 1737 718
rect 1690 688 1694 691
rect 1714 688 1718 691
rect 1646 672 1649 678
rect 1662 652 1665 688
rect 1678 672 1681 678
rect 1694 662 1697 668
rect 1702 662 1705 668
rect 1742 662 1745 698
rect 1674 658 1678 661
rect 1590 592 1593 608
rect 1670 592 1673 638
rect 1718 592 1721 628
rect 1758 582 1761 948
rect 1766 942 1769 948
rect 1766 922 1769 938
rect 1774 892 1777 948
rect 1822 912 1825 948
rect 1786 888 1790 891
rect 1822 872 1825 878
rect 1830 862 1833 868
rect 1822 852 1825 858
rect 1814 842 1817 848
rect 1830 842 1833 848
rect 1838 802 1841 1058
rect 1862 1032 1865 1058
rect 1870 1042 1873 1068
rect 1886 1062 1889 1068
rect 1970 1058 1974 1061
rect 1894 1042 1897 1058
rect 1854 952 1857 968
rect 1918 952 1921 1018
rect 1942 992 1945 1018
rect 1974 982 1977 988
rect 1930 958 1934 961
rect 1874 948 1878 951
rect 1846 942 1849 948
rect 1862 942 1865 948
rect 1894 942 1897 948
rect 1846 862 1849 918
rect 1894 892 1897 938
rect 1902 922 1905 948
rect 1910 942 1913 948
rect 1918 902 1921 918
rect 1890 878 1897 881
rect 1894 871 1897 878
rect 1894 868 1902 871
rect 1854 832 1857 868
rect 1874 858 1878 861
rect 1886 852 1889 868
rect 1926 862 1929 958
rect 1962 948 1966 951
rect 1986 948 1990 951
rect 1942 912 1945 918
rect 1854 812 1857 828
rect 1926 821 1929 838
rect 1918 818 1929 821
rect 1778 738 1782 741
rect 1806 672 1809 688
rect 1774 663 1777 668
rect 1822 662 1825 788
rect 1918 752 1921 818
rect 1874 748 1878 751
rect 1830 722 1833 747
rect 1902 742 1905 748
rect 1890 738 1894 741
rect 1846 732 1849 738
rect 1862 732 1865 738
rect 1910 722 1913 748
rect 1926 742 1929 758
rect 1870 692 1873 718
rect 1834 668 1838 671
rect 1886 662 1889 708
rect 1894 672 1897 698
rect 1842 658 1846 661
rect 1822 652 1825 658
rect 1574 562 1577 568
rect 1606 552 1609 568
rect 1630 562 1633 568
rect 1618 548 1622 551
rect 1646 542 1649 558
rect 1694 552 1697 568
rect 1742 552 1745 568
rect 1766 552 1769 558
rect 1706 548 1710 551
rect 1778 548 1782 551
rect 1586 488 1590 491
rect 1550 391 1553 478
rect 1558 462 1561 468
rect 1558 442 1561 448
rect 1566 432 1569 468
rect 1598 432 1601 538
rect 1686 512 1689 548
rect 1694 542 1697 548
rect 1702 492 1705 538
rect 1734 532 1737 548
rect 1750 532 1753 548
rect 1790 542 1793 558
rect 1798 552 1801 618
rect 1798 542 1801 548
rect 1750 522 1753 528
rect 1670 472 1673 478
rect 1646 452 1649 458
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1573 403 1576 407
rect 1550 388 1558 391
rect 1558 382 1561 388
rect 1542 342 1545 378
rect 1382 291 1385 328
rect 1414 302 1417 318
rect 1382 288 1390 291
rect 1374 262 1377 268
rect 1422 262 1425 268
rect 1446 262 1449 298
rect 1550 272 1553 288
rect 1566 282 1569 388
rect 1590 322 1593 338
rect 1614 332 1617 348
rect 1566 272 1569 278
rect 1346 258 1350 261
rect 1390 192 1393 238
rect 1406 152 1409 238
rect 1234 118 1238 121
rect 1198 82 1201 88
rect 1278 72 1281 78
rect 1294 72 1297 98
rect 1318 82 1321 138
rect 1342 72 1345 148
rect 1406 142 1409 148
rect 1470 142 1473 178
rect 1486 152 1489 268
rect 1494 262 1497 268
rect 1510 252 1513 268
rect 1518 252 1521 258
rect 1582 252 1585 259
rect 1590 242 1593 318
rect 1642 288 1646 291
rect 1654 272 1657 428
rect 1674 388 1678 391
rect 1686 382 1689 458
rect 1702 392 1705 398
rect 1674 348 1678 351
rect 1686 341 1689 348
rect 1678 338 1689 341
rect 1658 258 1662 261
rect 1662 242 1665 248
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1573 203 1576 207
rect 1590 152 1593 178
rect 1654 162 1657 198
rect 1678 192 1681 338
rect 1702 312 1705 378
rect 1686 252 1689 258
rect 1702 191 1705 308
rect 1710 292 1713 508
rect 1774 492 1777 528
rect 1802 518 1806 521
rect 1746 468 1750 471
rect 1718 432 1721 468
rect 1726 452 1729 458
rect 1754 448 1758 451
rect 1718 222 1721 348
rect 1726 332 1729 388
rect 1766 362 1769 458
rect 1822 452 1825 648
rect 1910 632 1913 718
rect 1902 552 1905 588
rect 1850 548 1854 551
rect 1854 482 1857 538
rect 1854 472 1857 478
rect 1830 462 1833 468
rect 1878 452 1881 468
rect 1854 372 1857 448
rect 1910 372 1913 548
rect 1942 542 1945 888
rect 1950 862 1953 868
rect 1950 752 1953 788
rect 1958 782 1961 898
rect 1974 892 1977 918
rect 1990 872 1993 888
rect 1998 871 2001 1068
rect 2014 1062 2017 1138
rect 2030 1092 2033 1308
rect 2042 1288 2046 1291
rect 2054 1271 2057 1318
rect 2080 1303 2082 1307
rect 2086 1303 2089 1307
rect 2093 1303 2096 1307
rect 2050 1268 2057 1271
rect 2094 1262 2097 1288
rect 2118 1262 2121 1318
rect 2134 1262 2137 1268
rect 2050 1258 2054 1261
rect 2106 1258 2110 1261
rect 2066 1248 2070 1251
rect 2054 1172 2057 1218
rect 2062 1192 2065 1238
rect 2094 1202 2097 1258
rect 2118 1192 2121 1198
rect 2150 1192 2153 1278
rect 2190 1262 2193 1318
rect 2230 1292 2233 1328
rect 2270 1292 2273 1338
rect 2242 1288 2246 1291
rect 2262 1262 2265 1288
rect 2374 1282 2377 1658
rect 2382 1532 2385 1658
rect 2458 1648 2462 1651
rect 2398 1342 2401 1608
rect 2414 1592 2417 1618
rect 2422 1542 2425 1548
rect 2414 1492 2417 1498
rect 2422 1472 2425 1528
rect 2418 1468 2422 1471
rect 2430 1462 2433 1648
rect 2502 1572 2505 1628
rect 2510 1612 2513 1658
rect 2566 1642 2569 1678
rect 2578 1668 2582 1671
rect 2590 1662 2593 1688
rect 2606 1661 2609 1758
rect 2614 1692 2617 1718
rect 2614 1672 2617 1678
rect 2602 1658 2609 1661
rect 2554 1568 2558 1571
rect 2462 1552 2465 1558
rect 2490 1548 2494 1551
rect 2502 1542 2505 1568
rect 2518 1552 2521 1558
rect 2546 1548 2550 1551
rect 2490 1538 2494 1541
rect 2530 1538 2534 1541
rect 2438 1482 2441 1538
rect 2446 1492 2449 1538
rect 2550 1532 2553 1538
rect 2470 1512 2473 1518
rect 2498 1488 2502 1491
rect 2470 1472 2473 1488
rect 2478 1472 2481 1478
rect 2450 1468 2454 1471
rect 2470 1462 2473 1468
rect 2558 1462 2561 1468
rect 2430 1452 2433 1458
rect 2450 1448 2454 1451
rect 2398 1282 2401 1338
rect 2406 1332 2409 1348
rect 2414 1342 2417 1368
rect 2422 1352 2425 1418
rect 2422 1292 2425 1338
rect 2430 1332 2433 1358
rect 2302 1272 2305 1278
rect 2078 1152 2081 1158
rect 2086 1152 2089 1178
rect 2150 1162 2153 1188
rect 2038 1142 2041 1148
rect 2054 1142 2057 1148
rect 2102 1122 2105 1138
rect 2054 1092 2057 1108
rect 2080 1103 2082 1107
rect 2086 1103 2089 1107
rect 2093 1103 2096 1107
rect 2102 1082 2105 1118
rect 2066 1078 2070 1081
rect 2046 1072 2049 1078
rect 2090 1058 2094 1061
rect 2014 982 2017 1058
rect 2062 1052 2065 1058
rect 2014 952 2017 978
rect 2018 948 2022 951
rect 2006 922 2009 928
rect 1998 868 2006 871
rect 1974 862 1977 868
rect 1990 862 1993 868
rect 1982 792 1985 818
rect 2006 792 2009 868
rect 1958 752 1961 778
rect 1966 762 1969 768
rect 1978 748 1982 751
rect 1986 738 1990 741
rect 1998 732 2001 738
rect 1974 682 1977 698
rect 2006 692 2009 738
rect 2030 692 2033 1018
rect 2046 902 2049 918
rect 2070 892 2073 1028
rect 2110 1022 2113 1148
rect 2126 1102 2129 1158
rect 2182 1152 2185 1248
rect 2214 1232 2217 1258
rect 2254 1212 2257 1258
rect 2286 1172 2289 1258
rect 2146 1148 2150 1151
rect 2226 1148 2230 1151
rect 2174 1142 2177 1148
rect 2182 1142 2185 1148
rect 2286 1142 2289 1168
rect 2134 1132 2137 1138
rect 2134 1092 2137 1128
rect 2126 1062 2129 1068
rect 2166 1061 2169 1118
rect 2214 1072 2217 1128
rect 2230 1082 2233 1088
rect 2258 1078 2262 1081
rect 2278 1072 2281 1078
rect 2186 1068 2190 1071
rect 2166 1058 2174 1061
rect 2266 1058 2270 1061
rect 2126 1042 2129 1058
rect 2230 1052 2233 1058
rect 2258 1048 2262 1051
rect 2082 1018 2086 1021
rect 2118 1012 2121 1018
rect 2082 918 2086 921
rect 2080 903 2082 907
rect 2086 903 2089 907
rect 2093 903 2096 907
rect 2050 868 2054 871
rect 2062 862 2065 868
rect 2054 682 2057 858
rect 2118 852 2121 918
rect 2118 842 2121 848
rect 2102 772 2105 778
rect 2082 758 2086 761
rect 2098 748 2102 751
rect 2126 742 2129 868
rect 2134 862 2137 1018
rect 2278 1012 2281 1068
rect 2294 1052 2297 1258
rect 2318 1192 2321 1218
rect 2326 1162 2329 1278
rect 2438 1262 2441 1318
rect 2370 1258 2374 1261
rect 2306 1158 2310 1161
rect 2326 1152 2329 1158
rect 2302 1142 2305 1148
rect 2334 1142 2337 1238
rect 2350 1222 2353 1258
rect 2438 1252 2441 1258
rect 2374 1152 2377 1248
rect 2446 1242 2449 1268
rect 2478 1262 2481 1268
rect 2454 1252 2457 1258
rect 2474 1248 2478 1251
rect 2346 1148 2350 1151
rect 2330 1138 2334 1141
rect 2350 1122 2353 1138
rect 2358 1132 2361 1138
rect 2366 1132 2369 1138
rect 2310 1092 2313 1108
rect 2326 1082 2329 1088
rect 2302 1072 2305 1078
rect 2302 1062 2305 1068
rect 2298 1048 2302 1051
rect 2290 1038 2294 1041
rect 2302 992 2305 1028
rect 2194 968 2198 971
rect 2270 952 2273 978
rect 2282 968 2286 971
rect 2310 952 2313 1018
rect 2318 1002 2321 1048
rect 2374 1022 2377 1148
rect 2382 1072 2385 1218
rect 2390 1182 2393 1188
rect 2422 1182 2425 1218
rect 2430 1152 2433 1208
rect 2462 1192 2465 1198
rect 2406 1132 2409 1148
rect 2422 1142 2425 1148
rect 2438 1142 2441 1168
rect 2454 1162 2457 1168
rect 2418 1128 2422 1131
rect 2406 1082 2409 1128
rect 2454 1122 2457 1128
rect 2386 1059 2390 1062
rect 2422 1062 2425 1078
rect 2430 1052 2433 1068
rect 2446 1062 2449 1078
rect 2438 1052 2441 1058
rect 2314 948 2318 951
rect 2142 891 2145 947
rect 2178 938 2182 941
rect 2158 912 2161 938
rect 2142 888 2150 891
rect 2142 872 2145 878
rect 2162 858 2166 861
rect 2150 842 2153 848
rect 2134 832 2137 838
rect 2174 812 2177 868
rect 2182 862 2185 918
rect 2198 892 2201 898
rect 2206 882 2209 928
rect 2190 862 2193 868
rect 2206 848 2214 851
rect 2206 792 2209 848
rect 2222 822 2225 928
rect 2230 902 2233 948
rect 2238 872 2241 878
rect 2270 862 2273 948
rect 2362 938 2366 941
rect 2330 928 2334 931
rect 2342 922 2345 938
rect 2278 872 2281 878
rect 2318 872 2321 888
rect 2334 863 2337 918
rect 2374 902 2377 958
rect 2382 952 2385 998
rect 2398 992 2401 1008
rect 2386 948 2390 951
rect 2398 892 2401 898
rect 2414 892 2417 908
rect 2230 852 2233 858
rect 2286 852 2289 858
rect 2230 762 2233 818
rect 2254 812 2257 818
rect 2218 758 2222 761
rect 2238 752 2241 808
rect 2162 748 2166 751
rect 2210 748 2214 751
rect 2066 738 2070 741
rect 2110 732 2113 738
rect 2080 703 2082 707
rect 2086 703 2089 707
rect 2093 703 2096 707
rect 2030 678 2038 681
rect 1974 672 1977 678
rect 2030 672 2033 678
rect 2054 672 2057 678
rect 2070 672 2073 698
rect 2126 692 2129 728
rect 2230 722 2233 748
rect 2238 742 2241 748
rect 2246 742 2249 778
rect 2262 762 2265 798
rect 2270 752 2273 768
rect 2294 762 2297 858
rect 2302 832 2305 848
rect 2302 762 2305 768
rect 2262 742 2265 748
rect 2102 678 2129 681
rect 2010 668 2017 671
rect 2102 671 2105 678
rect 2126 672 2129 678
rect 2150 678 2158 681
rect 2150 672 2153 678
rect 2174 672 2177 678
rect 2078 668 2105 671
rect 1998 662 2001 668
rect 1962 658 1966 661
rect 1994 648 2006 651
rect 1918 462 1921 518
rect 1742 352 1745 358
rect 1766 342 1769 358
rect 1818 348 1822 351
rect 1774 342 1777 348
rect 1758 332 1761 338
rect 1790 322 1793 338
rect 1818 288 1822 291
rect 1758 242 1761 258
rect 1702 188 1710 191
rect 1750 162 1753 228
rect 1770 158 1774 161
rect 1654 152 1657 158
rect 1750 152 1753 158
rect 1602 148 1606 151
rect 1350 92 1353 98
rect 1430 72 1433 78
rect 1446 72 1449 138
rect 1486 132 1489 138
rect 1510 132 1513 148
rect 1526 92 1529 148
rect 1662 142 1665 148
rect 1566 122 1569 138
rect 1646 132 1649 138
rect 1610 128 1614 131
rect 1686 92 1689 148
rect 1658 88 1662 91
rect 1510 72 1513 78
rect 1574 72 1577 78
rect 1098 68 1102 71
rect 1134 62 1137 68
rect 1174 62 1177 68
rect 1614 62 1617 78
rect 1686 72 1689 78
rect 946 58 950 61
rect 1122 58 1126 61
rect 1250 58 1254 61
rect 1338 58 1342 61
rect 1546 58 1550 61
rect 926 52 929 58
rect 1150 42 1153 58
rect 1310 52 1313 58
rect 1326 52 1329 58
rect 1390 52 1393 58
rect 1306 48 1310 51
rect 1174 42 1177 48
rect 510 -18 513 8
rect 544 3 546 7
rect 550 3 553 7
rect 557 3 560 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1573 3 1576 7
rect 510 -22 514 -18
rect 1702 -19 1705 138
rect 1710 82 1713 148
rect 1742 142 1745 148
rect 1770 138 1774 141
rect 1754 88 1758 91
rect 1790 82 1793 268
rect 1838 262 1841 358
rect 1846 292 1849 308
rect 1846 262 1849 288
rect 1830 222 1833 258
rect 1814 192 1817 218
rect 1830 172 1833 218
rect 1838 152 1841 158
rect 1798 122 1801 138
rect 1830 92 1833 148
rect 1854 142 1857 368
rect 1878 352 1881 358
rect 1886 342 1889 348
rect 1870 322 1873 328
rect 1862 192 1865 218
rect 1870 151 1873 158
rect 1886 152 1889 338
rect 1894 282 1897 348
rect 1902 332 1905 338
rect 1910 312 1913 368
rect 1942 352 1945 538
rect 1950 532 1953 618
rect 1966 552 1969 608
rect 2014 572 2017 668
rect 2026 658 2030 661
rect 2038 592 2041 668
rect 2078 662 2081 668
rect 2086 652 2089 658
rect 2110 651 2113 668
rect 2118 662 2121 668
rect 2146 658 2150 661
rect 2110 648 2121 651
rect 2110 632 2113 638
rect 2118 632 2121 648
rect 2126 642 2129 648
rect 1990 562 1993 568
rect 2022 552 2025 558
rect 2010 548 2014 551
rect 1958 522 1961 528
rect 1974 522 1977 548
rect 1998 522 2001 548
rect 1958 492 1961 518
rect 1966 392 1969 438
rect 1990 421 1993 468
rect 1998 462 2001 478
rect 2014 472 2017 548
rect 2022 482 2025 518
rect 1982 418 1993 421
rect 1970 348 1974 351
rect 1950 342 1953 348
rect 1934 332 1937 338
rect 1950 292 1953 338
rect 1906 288 1910 291
rect 1894 92 1897 278
rect 1958 262 1961 288
rect 1966 242 1969 268
rect 1982 192 1985 418
rect 2014 392 2017 448
rect 2046 442 2049 548
rect 2054 542 2057 628
rect 2062 552 2065 578
rect 2090 558 2094 561
rect 2098 548 2102 551
rect 2062 492 2065 548
rect 2138 547 2142 550
rect 2118 532 2121 538
rect 2080 503 2082 507
rect 2086 503 2089 507
rect 2093 503 2096 507
rect 2158 492 2161 668
rect 2190 652 2193 658
rect 2182 492 2185 558
rect 2198 531 2201 688
rect 2206 552 2209 718
rect 2238 662 2241 708
rect 2278 692 2281 748
rect 2294 712 2297 718
rect 2310 682 2313 818
rect 2330 778 2334 781
rect 2322 768 2326 771
rect 2318 752 2321 758
rect 2326 742 2329 748
rect 2246 662 2249 678
rect 2254 672 2257 678
rect 2222 592 2225 658
rect 2270 592 2273 628
rect 2254 552 2257 588
rect 2198 528 2209 531
rect 2114 478 2118 481
rect 2118 462 2121 468
rect 2134 462 2137 468
rect 2174 462 2177 488
rect 2198 472 2201 518
rect 2206 462 2209 528
rect 2230 492 2233 548
rect 2238 492 2241 548
rect 2246 542 2249 548
rect 2254 462 2257 548
rect 2262 542 2265 548
rect 2270 492 2273 568
rect 2074 458 2078 461
rect 2030 352 2033 358
rect 2038 352 2041 408
rect 2046 362 2049 418
rect 2126 412 2129 458
rect 2142 451 2145 458
rect 2134 448 2145 451
rect 2166 452 2169 458
rect 2134 392 2137 448
rect 2174 402 2177 458
rect 2214 452 2217 458
rect 2182 392 2185 438
rect 1990 332 1993 348
rect 2022 332 2025 348
rect 2038 312 2041 348
rect 2046 342 2049 358
rect 2070 352 2073 358
rect 2118 352 2121 388
rect 2150 352 2153 378
rect 2198 352 2201 358
rect 2070 342 2073 348
rect 2098 328 2102 331
rect 2002 268 2006 271
rect 1942 132 1945 148
rect 1930 118 1934 121
rect 1710 62 1713 78
rect 1762 68 1766 71
rect 1718 62 1721 68
rect 1730 58 1734 61
rect 1742 -18 1745 68
rect 1774 62 1777 78
rect 1910 72 1913 78
rect 1806 62 1809 68
rect 1958 62 1961 188
rect 1966 142 1969 148
rect 1998 142 2001 268
rect 2014 261 2017 308
rect 2054 292 2057 318
rect 2026 288 2030 291
rect 2054 272 2057 278
rect 2010 258 2017 261
rect 2030 252 2033 268
rect 2042 258 2046 261
rect 2046 152 2049 258
rect 2054 141 2057 268
rect 2070 172 2073 328
rect 2142 322 2145 348
rect 2158 332 2161 348
rect 2190 332 2193 348
rect 2162 328 2169 331
rect 2080 303 2082 307
rect 2086 303 2089 307
rect 2093 303 2096 307
rect 2166 292 2169 328
rect 2190 292 2193 298
rect 2206 292 2209 348
rect 2218 338 2222 341
rect 2238 332 2241 458
rect 2262 442 2265 458
rect 2254 352 2257 418
rect 2278 392 2281 658
rect 2294 552 2297 668
rect 2318 662 2321 708
rect 2326 622 2329 738
rect 2342 682 2345 828
rect 2382 792 2385 838
rect 2382 752 2385 768
rect 2414 742 2417 848
rect 2430 802 2433 948
rect 2454 932 2457 1118
rect 2470 1092 2473 1228
rect 2486 1212 2489 1418
rect 2494 1272 2497 1438
rect 2502 1342 2505 1347
rect 2518 1342 2521 1438
rect 2534 1332 2537 1348
rect 2542 1342 2545 1388
rect 2566 1372 2569 1618
rect 2590 1552 2593 1558
rect 2590 1491 2593 1548
rect 2598 1542 2601 1548
rect 2582 1488 2593 1491
rect 2582 1472 2585 1488
rect 2606 1432 2609 1658
rect 2622 1622 2625 1658
rect 2638 1482 2641 1738
rect 2646 1642 2649 1648
rect 2646 1452 2649 1468
rect 2606 1412 2609 1418
rect 2642 1388 2646 1391
rect 2574 1352 2577 1358
rect 2590 1352 2593 1368
rect 2550 1342 2553 1348
rect 2606 1342 2609 1348
rect 2594 1338 2598 1341
rect 2558 1332 2561 1338
rect 2582 1332 2585 1338
rect 2570 1328 2574 1331
rect 2502 1282 2505 1288
rect 2582 1282 2585 1328
rect 2614 1301 2617 1348
rect 2606 1298 2617 1301
rect 2494 1192 2497 1268
rect 2598 1262 2601 1268
rect 2554 1258 2558 1261
rect 2518 1152 2521 1158
rect 2542 1142 2545 1258
rect 2566 1142 2569 1168
rect 2586 1147 2590 1150
rect 2542 1132 2545 1138
rect 2466 1088 2470 1091
rect 2534 1072 2537 1088
rect 2514 1068 2518 1071
rect 2506 958 2510 961
rect 2462 932 2465 947
rect 2470 852 2473 868
rect 2434 748 2438 751
rect 2430 692 2433 748
rect 2454 742 2457 748
rect 2478 742 2481 868
rect 2494 762 2497 938
rect 2502 762 2505 958
rect 2550 952 2553 968
rect 2522 948 2526 951
rect 2510 942 2513 948
rect 2546 928 2550 931
rect 2534 922 2537 928
rect 2498 748 2502 751
rect 2438 732 2441 738
rect 2458 728 2462 731
rect 2466 718 2470 721
rect 2450 678 2454 681
rect 2382 672 2385 678
rect 2478 662 2481 668
rect 2486 662 2489 668
rect 2286 542 2289 548
rect 2302 472 2305 558
rect 2310 522 2313 548
rect 2318 532 2321 538
rect 2334 532 2337 658
rect 2342 542 2345 558
rect 2358 552 2361 598
rect 2366 552 2369 558
rect 2350 522 2353 548
rect 2358 521 2361 548
rect 2358 518 2369 521
rect 2350 511 2353 518
rect 2350 508 2361 511
rect 2350 472 2353 488
rect 2358 472 2361 508
rect 2330 468 2334 471
rect 2310 462 2313 468
rect 2286 432 2289 458
rect 2334 452 2337 458
rect 2366 451 2369 518
rect 2374 492 2377 558
rect 2406 551 2409 558
rect 2390 532 2393 538
rect 2414 512 2417 658
rect 2422 652 2425 658
rect 2422 572 2425 648
rect 2430 592 2433 658
rect 2438 652 2441 658
rect 2462 632 2465 658
rect 2494 622 2497 718
rect 2510 682 2513 918
rect 2502 652 2505 658
rect 2510 622 2513 658
rect 2482 548 2486 551
rect 2466 518 2470 521
rect 2478 492 2481 538
rect 2486 492 2489 538
rect 2382 482 2385 488
rect 2438 462 2441 468
rect 2366 448 2374 451
rect 2414 442 2417 458
rect 2262 352 2265 358
rect 2254 342 2257 348
rect 2222 302 2225 318
rect 2238 292 2241 328
rect 2226 288 2230 291
rect 2102 263 2105 288
rect 2134 262 2137 278
rect 2182 262 2185 268
rect 2262 262 2265 298
rect 2270 292 2273 348
rect 2302 272 2305 438
rect 2354 368 2358 371
rect 2326 362 2329 368
rect 2350 352 2353 358
rect 2366 352 2369 368
rect 2414 352 2417 368
rect 2310 342 2313 348
rect 2446 342 2449 478
rect 2462 342 2465 488
rect 2494 482 2497 618
rect 2510 552 2513 558
rect 2502 491 2505 518
rect 2518 501 2521 908
rect 2558 892 2561 1058
rect 2566 982 2569 988
rect 2574 952 2577 1078
rect 2606 1072 2609 1298
rect 2626 1288 2630 1291
rect 2638 1262 2641 1318
rect 2614 1248 2622 1251
rect 2614 1172 2617 1248
rect 2630 1242 2633 1248
rect 2646 1241 2649 1278
rect 2642 1238 2649 1241
rect 2642 1188 2646 1191
rect 2614 1082 2617 1168
rect 2618 1078 2622 1081
rect 2622 1062 2625 1068
rect 2574 932 2577 948
rect 2590 942 2593 948
rect 2598 942 2601 1048
rect 2614 972 2617 1018
rect 2586 928 2590 931
rect 2554 878 2558 881
rect 2562 868 2566 871
rect 2574 862 2577 868
rect 2582 852 2585 868
rect 2606 862 2609 918
rect 2622 902 2625 948
rect 2638 892 2641 1138
rect 2646 1052 2649 1058
rect 2646 972 2649 978
rect 2534 822 2537 848
rect 2526 818 2534 821
rect 2526 742 2529 818
rect 2526 652 2529 678
rect 2542 662 2545 758
rect 2562 718 2566 721
rect 2550 672 2553 688
rect 2558 672 2561 688
rect 2542 642 2545 648
rect 2550 582 2553 668
rect 2558 592 2561 628
rect 2534 552 2537 568
rect 2574 552 2577 718
rect 2606 652 2609 658
rect 2614 592 2617 748
rect 2638 742 2641 818
rect 2638 672 2641 738
rect 2586 568 2590 571
rect 2594 558 2598 561
rect 2546 548 2550 551
rect 2566 542 2569 548
rect 2574 542 2577 548
rect 2606 542 2609 578
rect 2610 538 2617 541
rect 2526 512 2529 538
rect 2518 498 2529 501
rect 2502 488 2513 491
rect 2510 462 2513 488
rect 2526 482 2529 498
rect 2590 492 2593 508
rect 2598 472 2601 538
rect 2614 472 2617 538
rect 2526 463 2529 468
rect 2598 462 2601 468
rect 2478 422 2481 458
rect 2470 352 2473 398
rect 2494 362 2497 398
rect 2494 342 2497 348
rect 2326 282 2329 318
rect 2358 312 2361 338
rect 2338 288 2342 291
rect 2398 282 2401 338
rect 2462 312 2465 338
rect 2170 258 2174 261
rect 2074 168 2086 171
rect 2122 168 2126 171
rect 2114 158 2118 161
rect 2182 152 2185 158
rect 2106 148 2110 151
rect 2050 138 2057 141
rect 2114 138 2118 141
rect 2038 131 2041 138
rect 2038 128 2049 131
rect 1982 72 1985 118
rect 2046 92 2049 128
rect 2010 88 2014 91
rect 2062 72 2065 118
rect 2080 103 2082 107
rect 2086 103 2089 107
rect 2093 103 2096 107
rect 2110 82 2113 88
rect 2134 72 2137 148
rect 2190 122 2193 128
rect 2182 72 2185 78
rect 2190 72 2193 118
rect 2206 102 2209 258
rect 2222 152 2225 218
rect 2270 162 2273 168
rect 2246 142 2249 148
rect 2254 102 2257 138
rect 2254 72 2257 88
rect 2150 62 2153 68
rect 1762 58 1766 61
rect 1882 58 1886 61
rect 2058 58 2062 61
rect 2142 52 2145 58
rect 2262 52 2265 118
rect 2270 81 2273 158
rect 2278 152 2281 208
rect 2286 152 2289 158
rect 2270 78 2281 81
rect 2270 62 2273 68
rect 2278 62 2281 78
rect 2286 72 2289 148
rect 2302 102 2305 268
rect 2318 152 2321 218
rect 2326 192 2329 278
rect 2430 272 2433 288
rect 2478 272 2481 308
rect 2386 268 2390 271
rect 2378 148 2382 151
rect 2310 142 2313 148
rect 2390 142 2393 268
rect 2398 263 2401 268
rect 2446 262 2449 268
rect 2470 252 2473 258
rect 2442 248 2446 251
rect 2478 142 2481 268
rect 2486 262 2489 298
rect 2502 292 2505 428
rect 2510 342 2513 368
rect 2510 262 2513 338
rect 2534 292 2537 458
rect 2610 448 2614 451
rect 2602 438 2606 441
rect 2614 352 2617 448
rect 2570 348 2574 351
rect 2498 258 2502 261
rect 2502 152 2505 178
rect 2518 162 2521 168
rect 2514 148 2518 151
rect 2490 138 2494 141
rect 2294 92 2297 98
rect 2374 72 2377 98
rect 2422 92 2425 138
rect 2478 102 2481 118
rect 2442 88 2446 91
rect 2390 72 2393 78
rect 2462 72 2465 88
rect 2346 58 2350 61
rect 2502 52 2505 148
rect 2526 142 2529 258
rect 2534 192 2537 278
rect 2566 242 2569 338
rect 2598 263 2601 348
rect 2614 312 2617 338
rect 2622 291 2625 668
rect 2630 562 2633 568
rect 2646 442 2649 448
rect 2630 352 2633 418
rect 2614 288 2625 291
rect 2614 272 2617 288
rect 2550 192 2553 198
rect 2542 162 2545 178
rect 2566 172 2569 238
rect 2602 148 2606 151
rect 2526 91 2529 138
rect 2526 88 2534 91
rect 2614 72 2617 128
rect 2566 62 2569 68
rect 2598 63 2601 68
rect 2522 58 2526 61
rect 2630 62 2633 338
rect 2638 282 2641 358
rect 2170 48 2174 51
rect 1718 -19 1722 -18
rect 1702 -22 1722 -19
rect 1742 -22 1746 -18
<< m3contact >>
rect 546 2403 550 2407
rect 553 2403 557 2407
rect 1562 2403 1566 2407
rect 1569 2403 1573 2407
rect 486 2398 490 2402
rect 502 2398 506 2402
rect 1174 2398 1178 2402
rect 1198 2398 1202 2402
rect 1526 2398 1530 2402
rect 2286 2398 2290 2402
rect 2302 2398 2306 2402
rect 214 2368 218 2372
rect 286 2368 290 2372
rect 294 2368 298 2372
rect 366 2368 370 2372
rect 358 2348 362 2352
rect 446 2348 450 2352
rect 14 2338 18 2342
rect 70 2338 74 2342
rect 230 2338 234 2342
rect 238 2338 242 2342
rect 6 2318 10 2322
rect 54 2318 58 2322
rect 62 2288 66 2292
rect 126 2268 130 2272
rect 70 2258 74 2262
rect 86 2258 90 2262
rect 70 2158 74 2162
rect 6 2128 10 2132
rect 62 2128 66 2132
rect 14 2118 18 2122
rect 54 2058 58 2062
rect 126 2148 130 2152
rect 118 2138 122 2142
rect 102 2118 106 2122
rect 102 2088 106 2092
rect 158 2288 162 2292
rect 190 2278 194 2282
rect 182 2258 186 2262
rect 206 2258 210 2262
rect 150 2248 154 2252
rect 174 2248 178 2252
rect 174 2238 178 2242
rect 150 2138 154 2142
rect 190 2138 194 2142
rect 150 2088 154 2092
rect 134 2078 138 2082
rect 214 2248 218 2252
rect 206 2108 210 2112
rect 174 2078 178 2082
rect 190 2078 194 2082
rect 102 2068 106 2072
rect 142 2068 146 2072
rect 118 2058 122 2062
rect 86 2048 90 2052
rect 86 1948 90 1952
rect 118 1948 122 1952
rect 6 1938 10 1942
rect 62 1938 66 1942
rect 62 1908 66 1912
rect 166 2058 170 2062
rect 134 2038 138 2042
rect 134 1898 138 1902
rect 102 1858 106 1862
rect 118 1858 122 1862
rect 38 1848 42 1852
rect 14 1718 18 1722
rect 38 1668 42 1672
rect 118 1848 122 1852
rect 142 1868 146 1872
rect 222 2238 226 2242
rect 254 2288 258 2292
rect 422 2278 426 2282
rect 318 2268 322 2272
rect 382 2268 386 2272
rect 398 2268 402 2272
rect 422 2268 426 2272
rect 318 2258 322 2262
rect 342 2258 346 2262
rect 430 2258 434 2262
rect 454 2258 458 2262
rect 334 2248 338 2252
rect 262 2238 266 2242
rect 350 2238 354 2242
rect 302 2188 306 2192
rect 262 2168 266 2172
rect 254 2128 258 2132
rect 318 2158 322 2162
rect 374 2158 378 2162
rect 366 2148 370 2152
rect 350 2128 354 2132
rect 374 2128 378 2132
rect 302 2118 306 2122
rect 350 2078 354 2082
rect 270 2058 274 2062
rect 198 1948 202 1952
rect 214 2028 218 2032
rect 206 1938 210 1942
rect 190 1928 194 1932
rect 190 1918 194 1922
rect 158 1848 162 1852
rect 142 1768 146 1772
rect 86 1748 90 1752
rect 134 1738 138 1742
rect 94 1708 98 1712
rect 78 1678 82 1682
rect 126 1668 130 1672
rect 118 1658 122 1662
rect 62 1648 66 1652
rect 126 1558 130 1562
rect 102 1498 106 1502
rect 102 1488 106 1492
rect 38 1478 42 1482
rect 102 1468 106 1472
rect 38 1448 42 1452
rect 198 1878 202 1882
rect 174 1738 178 1742
rect 158 1708 162 1712
rect 150 1698 154 1702
rect 214 1928 218 1932
rect 230 1928 234 1932
rect 222 1898 226 1902
rect 214 1778 218 1782
rect 390 2148 394 2152
rect 382 2118 386 2122
rect 326 2048 330 2052
rect 534 2368 538 2372
rect 926 2358 930 2362
rect 1038 2358 1042 2362
rect 1086 2358 1090 2362
rect 1142 2358 1146 2362
rect 622 2348 626 2352
rect 654 2348 658 2352
rect 814 2348 818 2352
rect 886 2348 890 2352
rect 982 2348 986 2352
rect 1022 2348 1026 2352
rect 1078 2348 1082 2352
rect 606 2318 610 2322
rect 494 2298 498 2302
rect 598 2278 602 2282
rect 478 2268 482 2272
rect 526 2268 530 2272
rect 574 2268 578 2272
rect 502 2258 506 2262
rect 518 2218 522 2222
rect 454 2178 458 2182
rect 430 2158 434 2162
rect 454 2158 458 2162
rect 414 2148 418 2152
rect 406 2098 410 2102
rect 414 2088 418 2092
rect 422 2078 426 2082
rect 446 2138 450 2142
rect 510 2138 514 2142
rect 494 2128 498 2132
rect 510 2128 514 2132
rect 454 2088 458 2092
rect 470 2088 474 2092
rect 406 2058 410 2062
rect 438 2058 442 2062
rect 390 2038 394 2042
rect 310 2018 314 2022
rect 270 1968 274 1972
rect 262 1958 266 1962
rect 278 1948 282 1952
rect 286 1928 290 1932
rect 246 1918 250 1922
rect 270 1918 274 1922
rect 270 1898 274 1902
rect 262 1888 266 1892
rect 286 1878 290 1882
rect 326 1978 330 1982
rect 318 1888 322 1892
rect 294 1858 298 1862
rect 270 1848 274 1852
rect 262 1768 266 1772
rect 238 1738 242 1742
rect 214 1728 218 1732
rect 254 1708 258 1712
rect 254 1688 258 1692
rect 142 1668 146 1672
rect 206 1668 210 1672
rect 150 1658 154 1662
rect 166 1648 170 1652
rect 206 1648 210 1652
rect 254 1578 258 1582
rect 190 1548 194 1552
rect 206 1548 210 1552
rect 230 1528 234 1532
rect 158 1498 162 1502
rect 134 1478 138 1482
rect 142 1468 146 1472
rect 150 1468 154 1472
rect 134 1458 138 1462
rect 142 1438 146 1442
rect 94 1408 98 1412
rect 118 1358 122 1362
rect 142 1358 146 1362
rect 46 1348 50 1352
rect 126 1348 130 1352
rect 182 1488 186 1492
rect 238 1478 242 1482
rect 190 1468 194 1472
rect 198 1468 202 1472
rect 238 1468 242 1472
rect 166 1458 170 1462
rect 182 1458 186 1462
rect 166 1438 170 1442
rect 198 1378 202 1382
rect 310 1778 314 1782
rect 294 1768 298 1772
rect 302 1758 306 1762
rect 390 1968 394 1972
rect 342 1958 346 1962
rect 366 1948 370 1952
rect 414 1938 418 1942
rect 342 1918 346 1922
rect 334 1848 338 1852
rect 390 1908 394 1912
rect 438 1988 442 1992
rect 422 1898 426 1902
rect 430 1888 434 1892
rect 382 1868 386 1872
rect 406 1868 410 1872
rect 438 1868 442 1872
rect 494 2058 498 2062
rect 478 2048 482 2052
rect 494 1978 498 1982
rect 546 2203 550 2207
rect 553 2203 557 2207
rect 598 2228 602 2232
rect 534 2138 538 2142
rect 558 2098 562 2102
rect 582 2098 586 2102
rect 566 2058 570 2062
rect 546 2003 550 2007
rect 553 2003 557 2007
rect 574 1958 578 1962
rect 526 1948 530 1952
rect 494 1938 498 1942
rect 510 1938 514 1942
rect 502 1868 506 1872
rect 350 1858 354 1862
rect 470 1858 474 1862
rect 422 1848 426 1852
rect 366 1838 370 1842
rect 414 1838 418 1842
rect 486 1838 490 1842
rect 534 1918 538 1922
rect 534 1908 538 1912
rect 518 1838 522 1842
rect 494 1818 498 1822
rect 334 1758 338 1762
rect 286 1748 290 1752
rect 318 1748 322 1752
rect 382 1758 386 1762
rect 430 1778 434 1782
rect 278 1718 282 1722
rect 334 1738 338 1742
rect 302 1668 306 1672
rect 342 1668 346 1672
rect 374 1728 378 1732
rect 366 1708 370 1712
rect 366 1678 370 1682
rect 334 1658 338 1662
rect 350 1658 354 1662
rect 374 1658 378 1662
rect 390 1748 394 1752
rect 654 2338 658 2342
rect 710 2338 714 2342
rect 686 2328 690 2332
rect 798 2328 802 2332
rect 670 2318 674 2322
rect 726 2318 730 2322
rect 758 2318 762 2322
rect 638 2288 642 2292
rect 686 2288 690 2292
rect 662 2268 666 2272
rect 750 2298 754 2302
rect 750 2278 754 2282
rect 646 2248 650 2252
rect 670 2248 674 2252
rect 734 2248 738 2252
rect 622 2238 626 2242
rect 638 2238 642 2242
rect 734 2218 738 2222
rect 662 2158 666 2162
rect 670 2158 674 2162
rect 678 2158 682 2162
rect 614 2148 618 2152
rect 686 2148 690 2152
rect 614 2138 618 2142
rect 638 2138 642 2142
rect 646 2128 650 2132
rect 638 2078 642 2082
rect 654 2058 658 2062
rect 654 1978 658 1982
rect 646 1948 650 1952
rect 622 1938 626 1942
rect 630 1928 634 1932
rect 590 1888 594 1892
rect 614 1888 618 1892
rect 558 1868 562 1872
rect 606 1868 610 1872
rect 678 2058 682 2062
rect 694 2028 698 2032
rect 670 1998 674 2002
rect 710 2078 714 2082
rect 742 2208 746 2212
rect 742 2168 746 2172
rect 734 2078 738 2082
rect 830 2308 834 2312
rect 870 2298 874 2302
rect 886 2288 890 2292
rect 806 2268 810 2272
rect 862 2268 866 2272
rect 902 2268 906 2272
rect 846 2258 850 2262
rect 878 2258 882 2262
rect 886 2238 890 2242
rect 838 2218 842 2222
rect 814 2188 818 2192
rect 798 2168 802 2172
rect 774 2158 778 2162
rect 758 2148 762 2152
rect 750 2098 754 2102
rect 750 2078 754 2082
rect 766 2068 770 2072
rect 702 1978 706 1982
rect 718 1978 722 1982
rect 694 1968 698 1972
rect 686 1958 690 1962
rect 670 1928 674 1932
rect 654 1918 658 1922
rect 662 1918 666 1922
rect 654 1908 658 1912
rect 702 1938 706 1942
rect 670 1878 674 1882
rect 694 1878 698 1882
rect 598 1858 602 1862
rect 638 1858 642 1862
rect 710 1908 714 1912
rect 702 1858 706 1862
rect 718 1858 722 1862
rect 550 1848 554 1852
rect 566 1848 570 1852
rect 662 1848 666 1852
rect 614 1838 618 1842
rect 546 1803 550 1807
rect 553 1803 557 1807
rect 582 1778 586 1782
rect 558 1768 562 1772
rect 446 1748 450 1752
rect 486 1748 490 1752
rect 526 1748 530 1752
rect 566 1748 570 1752
rect 406 1738 410 1742
rect 470 1738 474 1742
rect 414 1728 418 1732
rect 422 1718 426 1722
rect 406 1708 410 1712
rect 454 1708 458 1712
rect 390 1678 394 1682
rect 390 1668 394 1672
rect 398 1658 402 1662
rect 454 1658 458 1662
rect 278 1648 282 1652
rect 342 1648 346 1652
rect 358 1648 362 1652
rect 454 1568 458 1572
rect 382 1558 386 1562
rect 542 1738 546 1742
rect 494 1718 498 1722
rect 550 1718 554 1722
rect 582 1718 586 1722
rect 534 1708 538 1712
rect 486 1688 490 1692
rect 502 1688 506 1692
rect 526 1668 530 1672
rect 606 1698 610 1702
rect 518 1658 522 1662
rect 590 1658 594 1662
rect 582 1618 586 1622
rect 546 1603 550 1607
rect 553 1603 557 1607
rect 486 1588 490 1592
rect 590 1588 594 1592
rect 566 1578 570 1582
rect 582 1578 586 1582
rect 486 1558 490 1562
rect 414 1548 418 1552
rect 430 1548 434 1552
rect 534 1548 538 1552
rect 318 1538 322 1542
rect 294 1518 298 1522
rect 478 1538 482 1542
rect 518 1538 522 1542
rect 390 1518 394 1522
rect 422 1518 426 1522
rect 270 1418 274 1422
rect 222 1408 226 1412
rect 278 1368 282 1372
rect 294 1368 298 1372
rect 214 1348 218 1352
rect 230 1348 234 1352
rect 254 1348 258 1352
rect 14 1138 18 1142
rect 174 1288 178 1292
rect 150 1278 154 1282
rect 174 1278 178 1282
rect 118 1258 122 1262
rect 118 1168 122 1172
rect 166 1148 170 1152
rect 190 1288 194 1292
rect 182 1268 186 1272
rect 190 1258 194 1262
rect 198 1248 202 1252
rect 390 1498 394 1502
rect 390 1488 394 1492
rect 414 1468 418 1472
rect 366 1458 370 1462
rect 390 1458 394 1462
rect 310 1418 314 1422
rect 350 1448 354 1452
rect 406 1448 410 1452
rect 374 1428 378 1432
rect 334 1368 338 1372
rect 582 1538 586 1542
rect 454 1508 458 1512
rect 430 1358 434 1362
rect 310 1338 314 1342
rect 318 1338 322 1342
rect 222 1328 226 1332
rect 302 1328 306 1332
rect 214 1298 218 1302
rect 246 1288 250 1292
rect 382 1338 386 1342
rect 326 1308 330 1312
rect 302 1288 306 1292
rect 222 1278 226 1282
rect 262 1278 266 1282
rect 366 1278 370 1282
rect 406 1328 410 1332
rect 414 1308 418 1312
rect 422 1278 426 1282
rect 230 1268 234 1272
rect 270 1268 274 1272
rect 382 1268 386 1272
rect 406 1268 410 1272
rect 422 1268 426 1272
rect 326 1258 330 1262
rect 214 1248 218 1252
rect 190 1168 194 1172
rect 182 1158 186 1162
rect 174 1138 178 1142
rect 326 1248 330 1252
rect 214 1158 218 1162
rect 222 1148 226 1152
rect 246 1148 250 1152
rect 278 1138 282 1142
rect 294 1138 298 1142
rect 182 1128 186 1132
rect 198 1128 202 1132
rect 230 1128 234 1132
rect 270 1128 274 1132
rect 286 1128 290 1132
rect 302 1128 306 1132
rect 142 1088 146 1092
rect 150 1078 154 1082
rect 174 1078 178 1082
rect 30 1068 34 1072
rect 6 1048 10 1052
rect 22 1028 26 1032
rect 86 1058 90 1062
rect 166 1058 170 1062
rect 118 998 122 1002
rect 142 998 146 1002
rect 102 968 106 972
rect 62 948 66 952
rect 54 938 58 942
rect 46 858 50 862
rect 46 748 50 752
rect 6 668 10 672
rect 46 458 50 462
rect 6 388 10 392
rect 14 368 18 372
rect 38 368 42 372
rect 246 1118 250 1122
rect 190 1088 194 1092
rect 294 1108 298 1112
rect 302 1088 306 1092
rect 206 1058 210 1062
rect 294 988 298 992
rect 358 1168 362 1172
rect 398 1258 402 1262
rect 342 1148 346 1152
rect 334 1138 338 1142
rect 374 1138 378 1142
rect 366 1128 370 1132
rect 334 1108 338 1112
rect 342 1088 346 1092
rect 334 1058 338 1062
rect 374 1058 378 1062
rect 342 978 346 982
rect 366 978 370 982
rect 166 968 170 972
rect 158 958 162 962
rect 262 958 266 962
rect 222 948 226 952
rect 278 948 282 952
rect 118 938 122 942
rect 158 938 162 942
rect 102 918 106 922
rect 238 928 242 932
rect 174 888 178 892
rect 198 888 202 892
rect 118 858 122 862
rect 166 858 170 862
rect 222 868 226 872
rect 270 868 274 872
rect 214 848 218 852
rect 78 818 82 822
rect 350 958 354 962
rect 406 1148 410 1152
rect 390 1138 394 1142
rect 398 1118 402 1122
rect 518 1478 522 1482
rect 486 1458 490 1462
rect 502 1458 506 1462
rect 478 1358 482 1362
rect 454 1318 458 1322
rect 446 1298 450 1302
rect 438 1258 442 1262
rect 430 1168 434 1172
rect 414 1068 418 1072
rect 454 1278 458 1282
rect 502 1268 506 1272
rect 582 1468 586 1472
rect 534 1458 538 1462
rect 546 1403 550 1407
rect 553 1403 557 1407
rect 566 1368 570 1372
rect 550 1338 554 1342
rect 454 1228 458 1232
rect 462 1228 466 1232
rect 478 1248 482 1252
rect 486 1238 490 1242
rect 470 1218 474 1222
rect 470 1178 474 1182
rect 462 1158 466 1162
rect 454 1098 458 1102
rect 414 1038 418 1042
rect 430 1038 434 1042
rect 406 958 410 962
rect 462 958 466 962
rect 286 938 290 942
rect 390 938 394 942
rect 262 858 266 862
rect 254 828 258 832
rect 246 808 250 812
rect 126 758 130 762
rect 142 758 146 762
rect 278 768 282 772
rect 118 748 122 752
rect 254 748 258 752
rect 102 738 106 742
rect 190 728 194 732
rect 134 668 138 672
rect 78 658 82 662
rect 86 658 90 662
rect 70 548 74 552
rect 102 528 106 532
rect 254 718 258 722
rect 270 718 274 722
rect 182 708 186 712
rect 270 698 274 702
rect 198 688 202 692
rect 254 688 258 692
rect 238 678 242 682
rect 294 748 298 752
rect 286 718 290 722
rect 294 688 298 692
rect 294 678 298 682
rect 262 668 266 672
rect 278 668 282 672
rect 286 658 290 662
rect 158 648 162 652
rect 174 638 178 642
rect 150 558 154 562
rect 246 648 250 652
rect 206 548 210 552
rect 238 548 242 552
rect 158 528 162 532
rect 150 518 154 522
rect 142 478 146 482
rect 254 588 258 592
rect 246 518 250 522
rect 302 578 306 582
rect 270 568 274 572
rect 174 488 178 492
rect 182 488 186 492
rect 118 458 122 462
rect 166 458 170 462
rect 222 459 226 463
rect 134 388 138 392
rect 150 388 154 392
rect 118 358 122 362
rect 46 328 50 332
rect 70 328 74 332
rect 94 328 98 332
rect 110 328 114 332
rect 126 328 130 332
rect 62 268 66 272
rect 102 258 106 262
rect 126 258 130 262
rect 14 188 18 192
rect 86 158 90 162
rect 110 158 114 162
rect 118 158 122 162
rect 70 138 74 142
rect 70 118 74 122
rect 102 148 106 152
rect 174 338 178 342
rect 222 348 226 352
rect 190 328 194 332
rect 222 328 226 332
rect 262 488 266 492
rect 262 468 266 472
rect 294 558 298 562
rect 310 548 314 552
rect 294 518 298 522
rect 342 858 346 862
rect 438 918 442 922
rect 414 908 418 912
rect 398 858 402 862
rect 390 838 394 842
rect 438 858 442 862
rect 454 908 458 912
rect 454 868 458 872
rect 478 1148 482 1152
rect 558 1288 562 1292
rect 550 1278 554 1282
rect 542 1268 546 1272
rect 598 1558 602 1562
rect 598 1518 602 1522
rect 686 1848 690 1852
rect 678 1828 682 1832
rect 670 1768 674 1772
rect 710 1768 714 1772
rect 662 1748 666 1752
rect 622 1738 626 1742
rect 686 1758 690 1762
rect 702 1758 706 1762
rect 670 1738 674 1742
rect 686 1738 690 1742
rect 694 1708 698 1712
rect 710 1708 714 1712
rect 646 1688 650 1692
rect 734 1888 738 1892
rect 758 1948 762 1952
rect 790 2148 794 2152
rect 782 2108 786 2112
rect 806 2098 810 2102
rect 838 2168 842 2172
rect 862 2108 866 2112
rect 1110 2338 1114 2342
rect 950 2308 954 2312
rect 942 2298 946 2302
rect 934 2138 938 2142
rect 782 2068 786 2072
rect 1006 2328 1010 2332
rect 1030 2318 1034 2322
rect 1058 2303 1062 2307
rect 1065 2303 1069 2307
rect 1086 2318 1090 2322
rect 1078 2298 1082 2302
rect 1022 2288 1026 2292
rect 974 2228 978 2232
rect 950 2158 954 2162
rect 1118 2328 1122 2332
rect 1142 2338 1146 2342
rect 1158 2338 1162 2342
rect 1102 2298 1106 2302
rect 1094 2288 1098 2292
rect 1102 2268 1106 2272
rect 1070 2258 1074 2262
rect 1078 2248 1082 2252
rect 1078 2208 1082 2212
rect 1086 2188 1090 2192
rect 1078 2158 1082 2162
rect 1006 2138 1010 2142
rect 998 2098 1002 2102
rect 1014 2098 1018 2102
rect 982 2078 986 2082
rect 1054 2118 1058 2122
rect 1078 2118 1082 2122
rect 1058 2103 1062 2107
rect 1065 2103 1069 2107
rect 1038 2088 1042 2092
rect 1014 2078 1018 2082
rect 1022 2078 1026 2082
rect 1070 2068 1074 2072
rect 790 2058 794 2062
rect 854 2058 858 2062
rect 902 2058 906 2062
rect 926 2058 930 2062
rect 862 2038 866 2042
rect 902 2038 906 2042
rect 870 2008 874 2012
rect 894 2008 898 2012
rect 838 1968 842 1972
rect 846 1958 850 1962
rect 822 1948 826 1952
rect 766 1848 770 1852
rect 750 1748 754 1752
rect 766 1738 770 1742
rect 702 1698 706 1702
rect 710 1698 714 1702
rect 726 1698 730 1702
rect 878 1988 882 1992
rect 934 2048 938 2052
rect 950 1988 954 1992
rect 950 1978 954 1982
rect 918 1958 922 1962
rect 934 1958 938 1962
rect 918 1948 922 1952
rect 886 1938 890 1942
rect 806 1928 810 1932
rect 830 1908 834 1912
rect 822 1888 826 1892
rect 846 1888 850 1892
rect 934 1878 938 1882
rect 838 1848 842 1852
rect 854 1798 858 1802
rect 798 1748 802 1752
rect 822 1748 826 1752
rect 838 1748 842 1752
rect 854 1738 858 1742
rect 846 1728 850 1732
rect 822 1718 826 1722
rect 838 1718 842 1722
rect 806 1708 810 1712
rect 686 1658 690 1662
rect 670 1648 674 1652
rect 694 1648 698 1652
rect 694 1598 698 1602
rect 686 1558 690 1562
rect 646 1548 650 1552
rect 662 1508 666 1512
rect 670 1488 674 1492
rect 654 1468 658 1472
rect 750 1658 754 1662
rect 766 1648 770 1652
rect 766 1628 770 1632
rect 750 1568 754 1572
rect 798 1568 802 1572
rect 750 1548 754 1552
rect 790 1538 794 1542
rect 798 1538 802 1542
rect 854 1688 858 1692
rect 1046 2018 1050 2022
rect 998 1998 1002 2002
rect 990 1948 994 1952
rect 1006 1948 1010 1952
rect 1006 1888 1010 1892
rect 982 1868 986 1872
rect 1078 1978 1082 1982
rect 1118 2258 1122 2262
rect 1166 2298 1170 2302
rect 1182 2368 1186 2372
rect 1246 2368 1250 2372
rect 1262 2368 1266 2372
rect 1606 2368 1610 2372
rect 1622 2368 1626 2372
rect 1758 2368 1762 2372
rect 1766 2368 1770 2372
rect 1806 2368 1810 2372
rect 1942 2368 1946 2372
rect 1238 2348 1242 2352
rect 1262 2348 1266 2352
rect 1326 2348 1330 2352
rect 1206 2318 1210 2322
rect 1230 2318 1234 2322
rect 1158 2268 1162 2272
rect 1126 2168 1130 2172
rect 1110 2138 1114 2142
rect 1110 2128 1114 2132
rect 1198 2218 1202 2222
rect 1150 2188 1154 2192
rect 1222 2308 1226 2312
rect 1390 2358 1394 2362
rect 1422 2358 1426 2362
rect 1470 2358 1474 2362
rect 1534 2358 1538 2362
rect 1398 2348 1402 2352
rect 1422 2348 1426 2352
rect 1294 2328 1298 2332
rect 1366 2328 1370 2332
rect 1278 2308 1282 2312
rect 1222 2288 1226 2292
rect 1206 2168 1210 2172
rect 1142 2158 1146 2162
rect 1166 2148 1170 2152
rect 1198 2148 1202 2152
rect 1174 2138 1178 2142
rect 1142 2128 1146 2132
rect 1214 2128 1218 2132
rect 1158 2118 1162 2122
rect 1142 2108 1146 2112
rect 1222 2098 1226 2102
rect 1190 2088 1194 2092
rect 1166 2078 1170 2082
rect 1126 2058 1130 2062
rect 1166 2058 1170 2062
rect 1190 2048 1194 2052
rect 1118 2028 1122 2032
rect 1086 1968 1090 1972
rect 1030 1918 1034 1922
rect 1078 1918 1082 1922
rect 1058 1903 1062 1907
rect 1065 1903 1069 1907
rect 1046 1898 1050 1902
rect 1070 1888 1074 1892
rect 910 1858 914 1862
rect 1022 1858 1026 1862
rect 886 1798 890 1802
rect 902 1798 906 1802
rect 886 1708 890 1712
rect 862 1678 866 1682
rect 942 1848 946 1852
rect 934 1838 938 1842
rect 958 1778 962 1782
rect 990 1788 994 1792
rect 974 1768 978 1772
rect 1150 1958 1154 1962
rect 1214 1958 1218 1962
rect 1198 1948 1202 1952
rect 1222 1948 1226 1952
rect 1254 2268 1258 2272
rect 1358 2288 1362 2292
rect 1302 2268 1306 2272
rect 1430 2318 1434 2322
rect 1414 2288 1418 2292
rect 1382 2268 1386 2272
rect 1310 2258 1314 2262
rect 1334 2258 1338 2262
rect 1358 2258 1362 2262
rect 1382 2258 1386 2262
rect 1398 2258 1402 2262
rect 1414 2258 1418 2262
rect 1422 2258 1426 2262
rect 1262 2248 1266 2252
rect 1270 2238 1274 2242
rect 1382 2238 1386 2242
rect 1462 2328 1466 2332
rect 1494 2328 1498 2332
rect 1446 2298 1450 2302
rect 1486 2298 1490 2302
rect 1638 2358 1642 2362
rect 1686 2358 1690 2362
rect 1854 2358 1858 2362
rect 1886 2358 1890 2362
rect 1822 2348 1826 2352
rect 1838 2348 1842 2352
rect 2038 2348 2042 2352
rect 2070 2348 2074 2352
rect 2214 2348 2218 2352
rect 1606 2338 1610 2342
rect 1646 2338 1650 2342
rect 1758 2338 1762 2342
rect 1822 2338 1826 2342
rect 1854 2338 1858 2342
rect 1654 2328 1658 2332
rect 1486 2288 1490 2292
rect 1526 2288 1530 2292
rect 1550 2288 1554 2292
rect 1470 2258 1474 2262
rect 1406 2228 1410 2232
rect 1430 2228 1434 2232
rect 1382 2218 1386 2222
rect 1238 2208 1242 2212
rect 1270 2208 1274 2212
rect 1262 2178 1266 2182
rect 1662 2278 1666 2282
rect 1590 2268 1594 2272
rect 1630 2268 1634 2272
rect 1742 2298 1746 2302
rect 1766 2298 1770 2302
rect 1726 2268 1730 2272
rect 1534 2258 1538 2262
rect 1558 2258 1562 2262
rect 1686 2258 1690 2262
rect 1774 2288 1778 2292
rect 1790 2278 1794 2282
rect 1774 2268 1778 2272
rect 1814 2268 1818 2272
rect 1854 2328 1858 2332
rect 1846 2268 1850 2272
rect 1758 2258 1762 2262
rect 1782 2258 1786 2262
rect 1854 2258 1858 2262
rect 1518 2248 1522 2252
rect 1562 2203 1566 2207
rect 1569 2203 1573 2207
rect 1534 2198 1538 2202
rect 1614 2168 1618 2172
rect 1526 2158 1530 2162
rect 1294 2148 1298 2152
rect 1310 2148 1314 2152
rect 1486 2148 1490 2152
rect 1598 2148 1602 2152
rect 1350 2138 1354 2142
rect 1294 2128 1298 2132
rect 1422 2128 1426 2132
rect 1334 2118 1338 2122
rect 1502 2118 1506 2122
rect 1510 2118 1514 2122
rect 1270 2108 1274 2112
rect 1414 2088 1418 2092
rect 1278 2078 1282 2082
rect 1366 2078 1370 2082
rect 1414 2078 1418 2082
rect 1462 2078 1466 2082
rect 1478 2078 1482 2082
rect 1286 1968 1290 1972
rect 1270 1948 1274 1952
rect 1182 1918 1186 1922
rect 1158 1888 1162 1892
rect 1206 1878 1210 1882
rect 1126 1868 1130 1872
rect 1182 1868 1186 1872
rect 1142 1858 1146 1862
rect 1214 1858 1218 1862
rect 1350 2038 1354 2042
rect 1318 1958 1322 1962
rect 1350 1958 1354 1962
rect 1318 1948 1322 1952
rect 1462 2058 1466 2062
rect 1422 2048 1426 2052
rect 1446 2038 1450 2042
rect 1422 2028 1426 2032
rect 1422 2018 1426 2022
rect 1406 1968 1410 1972
rect 1454 1968 1458 1972
rect 1542 2078 1546 2082
rect 1686 2168 1690 2172
rect 1774 2168 1778 2172
rect 1742 2158 1746 2162
rect 1758 2158 1762 2162
rect 1678 2138 1682 2142
rect 1790 2238 1794 2242
rect 1814 2238 1818 2242
rect 1846 2248 1850 2252
rect 1830 2238 1834 2242
rect 1822 2228 1826 2232
rect 1966 2298 1970 2302
rect 2222 2338 2226 2342
rect 2246 2338 2250 2342
rect 1990 2288 1994 2292
rect 1998 2288 2002 2292
rect 2014 2288 2018 2292
rect 1958 2278 1962 2282
rect 1966 2278 1970 2282
rect 1990 2278 1994 2282
rect 1902 2248 1906 2252
rect 1870 2158 1874 2162
rect 1790 2148 1794 2152
rect 1814 2148 1818 2152
rect 1838 2148 1842 2152
rect 1854 2138 1858 2142
rect 1782 2128 1786 2132
rect 1822 2128 1826 2132
rect 1830 2078 1834 2082
rect 1622 2068 1626 2072
rect 1638 2068 1642 2072
rect 1710 2068 1714 2072
rect 1534 2038 1538 2042
rect 1550 2038 1554 2042
rect 1534 2028 1538 2032
rect 1542 2028 1546 2032
rect 1574 2018 1578 2022
rect 1562 2003 1566 2007
rect 1569 2003 1573 2007
rect 1582 1958 1586 1962
rect 1558 1948 1562 1952
rect 1310 1938 1314 1942
rect 1366 1938 1370 1942
rect 1302 1928 1306 1932
rect 1262 1898 1266 1902
rect 1310 1888 1314 1892
rect 1230 1868 1234 1872
rect 1326 1858 1330 1862
rect 1182 1848 1186 1852
rect 1198 1848 1202 1852
rect 1222 1848 1226 1852
rect 1094 1838 1098 1842
rect 1046 1808 1050 1812
rect 1054 1768 1058 1772
rect 998 1758 1002 1762
rect 1014 1758 1018 1762
rect 974 1748 978 1752
rect 950 1738 954 1742
rect 926 1678 930 1682
rect 966 1678 970 1682
rect 982 1678 986 1682
rect 958 1668 962 1672
rect 870 1658 874 1662
rect 886 1658 890 1662
rect 942 1658 946 1662
rect 966 1658 970 1662
rect 846 1608 850 1612
rect 990 1648 994 1652
rect 974 1638 978 1642
rect 998 1638 1002 1642
rect 950 1628 954 1632
rect 982 1598 986 1602
rect 910 1578 914 1582
rect 870 1568 874 1572
rect 822 1558 826 1562
rect 814 1548 818 1552
rect 838 1548 842 1552
rect 806 1528 810 1532
rect 742 1498 746 1502
rect 758 1498 762 1502
rect 782 1498 786 1502
rect 718 1468 722 1472
rect 798 1468 802 1472
rect 822 1468 826 1472
rect 630 1458 634 1462
rect 614 1448 618 1452
rect 638 1448 642 1452
rect 662 1448 666 1452
rect 702 1448 706 1452
rect 710 1448 714 1452
rect 750 1448 754 1452
rect 606 1368 610 1372
rect 590 1328 594 1332
rect 662 1338 666 1342
rect 630 1278 634 1282
rect 526 1248 530 1252
rect 534 1248 538 1252
rect 598 1248 602 1252
rect 614 1248 618 1252
rect 582 1228 586 1232
rect 546 1203 550 1207
rect 553 1203 557 1207
rect 670 1288 674 1292
rect 670 1278 674 1282
rect 862 1538 866 1542
rect 846 1508 850 1512
rect 894 1538 898 1542
rect 934 1538 938 1542
rect 910 1528 914 1532
rect 902 1518 906 1522
rect 854 1498 858 1502
rect 886 1498 890 1502
rect 870 1458 874 1462
rect 838 1418 842 1422
rect 966 1508 970 1512
rect 918 1498 922 1502
rect 998 1578 1002 1582
rect 1070 1758 1074 1762
rect 1094 1758 1098 1762
rect 1102 1748 1106 1752
rect 1118 1748 1122 1752
rect 1078 1738 1082 1742
rect 1038 1728 1042 1732
rect 1046 1708 1050 1712
rect 1058 1703 1062 1707
rect 1065 1703 1069 1707
rect 1046 1678 1050 1682
rect 1062 1618 1066 1622
rect 1030 1598 1034 1602
rect 1022 1568 1026 1572
rect 990 1548 994 1552
rect 1014 1548 1018 1552
rect 1038 1548 1042 1552
rect 1062 1548 1066 1552
rect 1062 1538 1066 1542
rect 1046 1528 1050 1532
rect 1058 1503 1062 1507
rect 1065 1503 1069 1507
rect 998 1478 1002 1482
rect 966 1468 970 1472
rect 926 1458 930 1462
rect 982 1458 986 1462
rect 1006 1458 1010 1462
rect 1022 1448 1026 1452
rect 1070 1448 1074 1452
rect 998 1438 1002 1442
rect 886 1388 890 1392
rect 910 1388 914 1392
rect 854 1358 858 1362
rect 862 1358 866 1362
rect 886 1358 890 1362
rect 726 1348 730 1352
rect 822 1348 826 1352
rect 702 1298 706 1302
rect 726 1298 730 1302
rect 686 1288 690 1292
rect 718 1288 722 1292
rect 726 1278 730 1282
rect 654 1268 658 1272
rect 678 1258 682 1262
rect 654 1248 658 1252
rect 646 1238 650 1242
rect 654 1218 658 1222
rect 518 1178 522 1182
rect 590 1178 594 1182
rect 638 1178 642 1182
rect 534 1148 538 1152
rect 550 1148 554 1152
rect 510 1138 514 1142
rect 534 1108 538 1112
rect 542 1108 546 1112
rect 534 1098 538 1102
rect 606 1128 610 1132
rect 622 1108 626 1112
rect 574 1098 578 1102
rect 510 1048 514 1052
rect 590 1038 594 1042
rect 546 1003 550 1007
rect 553 1003 557 1007
rect 566 988 570 992
rect 478 958 482 962
rect 478 938 482 942
rect 486 888 490 892
rect 526 878 530 882
rect 550 868 554 872
rect 654 1148 658 1152
rect 742 1248 746 1252
rect 726 1218 730 1222
rect 782 1328 786 1332
rect 998 1368 1002 1372
rect 1006 1358 1010 1362
rect 1038 1438 1042 1442
rect 1022 1428 1026 1432
rect 1038 1388 1042 1392
rect 1046 1368 1050 1372
rect 1102 1728 1106 1732
rect 1118 1718 1122 1722
rect 1086 1668 1090 1672
rect 1150 1768 1154 1772
rect 1142 1758 1146 1762
rect 1182 1748 1186 1752
rect 1134 1738 1138 1742
rect 1134 1698 1138 1702
rect 1166 1728 1170 1732
rect 1182 1728 1186 1732
rect 1374 1878 1378 1882
rect 1398 1868 1402 1872
rect 1270 1778 1274 1782
rect 1334 1778 1338 1782
rect 1342 1778 1346 1782
rect 1230 1748 1234 1752
rect 1174 1688 1178 1692
rect 1198 1688 1202 1692
rect 1158 1668 1162 1672
rect 1142 1658 1146 1662
rect 1150 1658 1154 1662
rect 1110 1548 1114 1552
rect 1102 1538 1106 1542
rect 1110 1508 1114 1512
rect 1102 1488 1106 1492
rect 1318 1748 1322 1752
rect 1246 1738 1250 1742
rect 1462 1888 1466 1892
rect 1430 1878 1434 1882
rect 1478 1858 1482 1862
rect 1422 1848 1426 1852
rect 1390 1828 1394 1832
rect 1414 1828 1418 1832
rect 1590 1948 1594 1952
rect 1606 2048 1610 2052
rect 1534 1938 1538 1942
rect 1598 1938 1602 1942
rect 1558 1928 1562 1932
rect 1598 1868 1602 1872
rect 1518 1858 1522 1862
rect 1510 1828 1514 1832
rect 1562 1803 1566 1807
rect 1569 1803 1573 1807
rect 1806 2058 1810 2062
rect 1846 2058 1850 2062
rect 1630 2038 1634 2042
rect 1670 1958 1674 1962
rect 1734 1978 1738 1982
rect 1790 2008 1794 2012
rect 1846 2038 1850 2042
rect 2134 2328 2138 2332
rect 2082 2303 2086 2307
rect 2089 2303 2093 2307
rect 2046 2288 2050 2292
rect 2102 2288 2106 2292
rect 2038 2268 2042 2272
rect 1934 2258 1938 2262
rect 1950 2218 1954 2222
rect 1998 2218 2002 2222
rect 1926 2178 1930 2182
rect 1934 2128 1938 2132
rect 1942 2118 1946 2122
rect 1910 2078 1914 2082
rect 1902 2038 1906 2042
rect 1982 2168 1986 2172
rect 1958 2148 1962 2152
rect 1966 2118 1970 2122
rect 1974 2108 1978 2112
rect 1990 2108 1994 2112
rect 1966 2098 1970 2102
rect 1942 2018 1946 2022
rect 1854 2008 1858 2012
rect 1886 2008 1890 2012
rect 1870 1988 1874 1992
rect 1822 1948 1826 1952
rect 1838 1948 1842 1952
rect 1798 1938 1802 1942
rect 1718 1928 1722 1932
rect 1790 1928 1794 1932
rect 1694 1918 1698 1922
rect 1646 1908 1650 1912
rect 1638 1878 1642 1882
rect 1654 1878 1658 1882
rect 1654 1868 1658 1872
rect 1710 1878 1714 1882
rect 1750 1888 1754 1892
rect 1790 1878 1794 1882
rect 1622 1858 1626 1862
rect 1654 1808 1658 1812
rect 1622 1788 1626 1792
rect 1422 1768 1426 1772
rect 1486 1768 1490 1772
rect 1606 1768 1610 1772
rect 1646 1768 1650 1772
rect 1694 1768 1698 1772
rect 1382 1748 1386 1752
rect 1310 1738 1314 1742
rect 1366 1738 1370 1742
rect 1278 1728 1282 1732
rect 1294 1728 1298 1732
rect 1326 1728 1330 1732
rect 1246 1708 1250 1712
rect 1214 1678 1218 1682
rect 1230 1678 1234 1682
rect 1198 1668 1202 1672
rect 1358 1678 1362 1682
rect 1398 1678 1402 1682
rect 1406 1678 1410 1682
rect 1326 1668 1330 1672
rect 1390 1668 1394 1672
rect 1286 1658 1290 1662
rect 1366 1658 1370 1662
rect 1398 1658 1402 1662
rect 1206 1648 1210 1652
rect 1254 1648 1258 1652
rect 1294 1638 1298 1642
rect 1246 1578 1250 1582
rect 1262 1578 1266 1582
rect 1294 1578 1298 1582
rect 1206 1568 1210 1572
rect 1278 1568 1282 1572
rect 1270 1558 1274 1562
rect 1358 1558 1362 1562
rect 1302 1548 1306 1552
rect 1366 1548 1370 1552
rect 1142 1538 1146 1542
rect 1158 1538 1162 1542
rect 1206 1538 1210 1542
rect 1134 1528 1138 1532
rect 1134 1518 1138 1522
rect 1142 1498 1146 1502
rect 1118 1478 1122 1482
rect 1150 1478 1154 1482
rect 1182 1478 1186 1482
rect 1222 1528 1226 1532
rect 1214 1508 1218 1512
rect 1262 1508 1266 1512
rect 1134 1458 1138 1462
rect 1190 1458 1194 1462
rect 1222 1498 1226 1502
rect 1270 1478 1274 1482
rect 1262 1458 1266 1462
rect 1206 1438 1210 1442
rect 1070 1398 1074 1402
rect 1182 1408 1186 1412
rect 1070 1358 1074 1362
rect 1078 1358 1082 1362
rect 1214 1358 1218 1362
rect 1246 1358 1250 1362
rect 862 1348 866 1352
rect 1006 1348 1010 1352
rect 1022 1348 1026 1352
rect 1062 1348 1066 1352
rect 1094 1348 1098 1352
rect 1150 1348 1154 1352
rect 1230 1348 1234 1352
rect 1254 1348 1258 1352
rect 782 1278 786 1282
rect 806 1278 810 1282
rect 822 1278 826 1282
rect 846 1278 850 1282
rect 862 1278 866 1282
rect 878 1278 882 1282
rect 790 1258 794 1262
rect 798 1238 802 1242
rect 790 1218 794 1222
rect 798 1208 802 1212
rect 702 1158 706 1162
rect 742 1158 746 1162
rect 862 1268 866 1272
rect 846 1258 850 1262
rect 838 1238 842 1242
rect 1158 1338 1162 1342
rect 1214 1338 1218 1342
rect 1286 1338 1290 1342
rect 886 1268 890 1272
rect 862 1248 866 1252
rect 870 1248 874 1252
rect 1030 1328 1034 1332
rect 1078 1328 1082 1332
rect 1094 1328 1098 1332
rect 1166 1328 1170 1332
rect 1198 1328 1202 1332
rect 982 1318 986 1322
rect 982 1308 986 1312
rect 902 1298 906 1302
rect 846 1218 850 1222
rect 894 1218 898 1222
rect 742 1148 746 1152
rect 774 1148 778 1152
rect 686 1138 690 1142
rect 710 1138 714 1142
rect 734 1138 738 1142
rect 686 1128 690 1132
rect 678 1108 682 1112
rect 638 1088 642 1092
rect 678 1088 682 1092
rect 726 1128 730 1132
rect 758 1138 762 1142
rect 750 1128 754 1132
rect 782 1108 786 1112
rect 718 1068 722 1072
rect 774 1068 778 1072
rect 670 1058 674 1062
rect 710 1058 714 1062
rect 726 1058 730 1062
rect 654 1048 658 1052
rect 646 958 650 962
rect 582 938 586 942
rect 590 928 594 932
rect 518 858 522 862
rect 574 858 578 862
rect 422 838 426 842
rect 406 768 410 772
rect 406 758 410 762
rect 446 748 450 752
rect 334 708 338 712
rect 342 708 346 712
rect 390 738 394 742
rect 358 678 362 682
rect 374 678 378 682
rect 350 668 354 672
rect 398 678 402 682
rect 390 658 394 662
rect 358 648 362 652
rect 334 638 338 642
rect 358 638 362 642
rect 334 628 338 632
rect 350 538 354 542
rect 446 698 450 702
rect 422 638 426 642
rect 430 638 434 642
rect 454 618 458 622
rect 446 608 450 612
rect 406 578 410 582
rect 414 578 418 582
rect 414 568 418 572
rect 422 558 426 562
rect 478 848 482 852
rect 742 1048 746 1052
rect 758 1018 762 1022
rect 710 958 714 962
rect 702 948 706 952
rect 734 948 738 952
rect 750 948 754 952
rect 702 938 706 942
rect 638 928 642 932
rect 646 928 650 932
rect 646 908 650 912
rect 598 898 602 902
rect 622 898 626 902
rect 606 878 610 882
rect 654 858 658 862
rect 546 803 550 807
rect 553 803 557 807
rect 574 798 578 802
rect 518 748 522 752
rect 750 928 754 932
rect 822 1138 826 1142
rect 854 1198 858 1202
rect 862 1168 866 1172
rect 878 1168 882 1172
rect 854 1158 858 1162
rect 830 1108 834 1112
rect 846 1108 850 1112
rect 838 1068 842 1072
rect 894 1208 898 1212
rect 886 1148 890 1152
rect 1058 1303 1062 1307
rect 1065 1303 1069 1307
rect 1038 1298 1042 1302
rect 1014 1288 1018 1292
rect 1038 1288 1042 1292
rect 926 1278 930 1282
rect 918 1208 922 1212
rect 1038 1268 1042 1272
rect 1102 1308 1106 1312
rect 1094 1298 1098 1302
rect 1054 1248 1058 1252
rect 1094 1248 1098 1252
rect 1150 1278 1154 1282
rect 1206 1308 1210 1312
rect 1198 1298 1202 1302
rect 1254 1328 1258 1332
rect 1262 1328 1266 1332
rect 1278 1318 1282 1322
rect 1254 1308 1258 1312
rect 1110 1268 1114 1272
rect 1174 1268 1178 1272
rect 1134 1258 1138 1262
rect 1182 1258 1186 1262
rect 1198 1258 1202 1262
rect 1094 1228 1098 1232
rect 974 1198 978 1202
rect 1086 1208 1090 1212
rect 902 1158 906 1162
rect 1030 1158 1034 1162
rect 926 1148 930 1152
rect 1046 1148 1050 1152
rect 910 1138 914 1142
rect 1014 1138 1018 1142
rect 910 1128 914 1132
rect 894 1068 898 1072
rect 854 1058 858 1062
rect 870 1058 874 1062
rect 798 998 802 1002
rect 782 918 786 922
rect 750 908 754 912
rect 718 878 722 882
rect 766 888 770 892
rect 790 898 794 902
rect 726 858 730 862
rect 670 848 674 852
rect 702 848 706 852
rect 742 848 746 852
rect 638 798 642 802
rect 638 778 642 782
rect 598 768 602 772
rect 694 768 698 772
rect 718 768 722 772
rect 734 758 738 762
rect 662 748 666 752
rect 838 1048 842 1052
rect 862 1048 866 1052
rect 886 1048 890 1052
rect 822 968 826 972
rect 822 938 826 942
rect 806 888 810 892
rect 766 858 770 862
rect 766 828 770 832
rect 790 828 794 832
rect 766 798 770 802
rect 774 748 778 752
rect 470 718 474 722
rect 470 688 474 692
rect 518 678 522 682
rect 502 668 506 672
rect 486 658 490 662
rect 478 638 482 642
rect 510 628 514 632
rect 518 628 522 632
rect 510 558 514 562
rect 430 538 434 542
rect 350 518 354 522
rect 334 488 338 492
rect 358 488 362 492
rect 318 468 322 472
rect 406 518 410 522
rect 390 488 394 492
rect 278 458 282 462
rect 326 458 330 462
rect 358 458 362 462
rect 310 448 314 452
rect 278 358 282 362
rect 294 358 298 362
rect 270 328 274 332
rect 382 418 386 422
rect 430 488 434 492
rect 518 488 522 492
rect 638 728 642 732
rect 710 728 714 732
rect 566 718 570 722
rect 590 718 594 722
rect 678 718 682 722
rect 534 698 538 702
rect 542 688 546 692
rect 590 688 594 692
rect 646 668 650 672
rect 654 668 658 672
rect 662 668 666 672
rect 694 668 698 672
rect 566 658 570 662
rect 582 658 586 662
rect 702 658 706 662
rect 542 648 546 652
rect 622 628 626 632
rect 546 603 550 607
rect 553 603 557 607
rect 718 638 722 642
rect 574 578 578 582
rect 694 578 698 582
rect 694 568 698 572
rect 598 558 602 562
rect 678 558 682 562
rect 558 528 562 532
rect 582 538 586 542
rect 630 538 634 542
rect 670 538 674 542
rect 718 538 722 542
rect 622 528 626 532
rect 638 528 642 532
rect 574 508 578 512
rect 598 508 602 512
rect 686 508 690 512
rect 718 498 722 502
rect 630 488 634 492
rect 670 488 674 492
rect 686 488 690 492
rect 710 488 714 492
rect 526 478 530 482
rect 486 468 490 472
rect 534 468 538 472
rect 574 468 578 472
rect 534 458 538 462
rect 766 728 770 732
rect 766 678 770 682
rect 774 668 778 672
rect 806 778 810 782
rect 878 928 882 932
rect 838 898 842 902
rect 830 888 834 892
rect 838 868 842 872
rect 990 1108 994 1112
rect 1058 1103 1062 1107
rect 1065 1103 1069 1107
rect 950 1088 954 1092
rect 1062 1088 1066 1092
rect 910 1028 914 1032
rect 902 978 906 982
rect 934 1048 938 1052
rect 926 1018 930 1022
rect 1038 1078 1042 1082
rect 998 1058 1002 1062
rect 1022 1048 1026 1052
rect 990 998 994 1002
rect 950 978 954 982
rect 918 958 922 962
rect 958 948 962 952
rect 902 938 906 942
rect 974 928 978 932
rect 926 908 930 912
rect 982 908 986 912
rect 918 888 922 892
rect 926 888 930 892
rect 926 848 930 852
rect 886 838 890 842
rect 918 838 922 842
rect 846 828 850 832
rect 998 878 1002 882
rect 942 778 946 782
rect 934 768 938 772
rect 894 758 898 762
rect 918 758 922 762
rect 942 758 946 762
rect 958 758 962 762
rect 846 748 850 752
rect 878 748 882 752
rect 814 738 818 742
rect 894 728 898 732
rect 918 698 922 702
rect 894 688 898 692
rect 830 678 834 682
rect 918 678 922 682
rect 894 668 898 672
rect 950 708 954 712
rect 1038 1038 1042 1042
rect 1158 1248 1162 1252
rect 1182 1248 1186 1252
rect 1206 1248 1210 1252
rect 1142 1228 1146 1232
rect 1190 1228 1194 1232
rect 1134 1218 1138 1222
rect 1198 1148 1202 1152
rect 1102 1128 1106 1132
rect 1094 1108 1098 1112
rect 1110 1088 1114 1092
rect 1118 1088 1122 1092
rect 1102 1078 1106 1082
rect 1158 1068 1162 1072
rect 1118 1058 1122 1062
rect 1094 1038 1098 1042
rect 1150 968 1154 972
rect 1134 948 1138 952
rect 1038 938 1042 942
rect 1062 928 1066 932
rect 1030 908 1034 912
rect 1058 903 1062 907
rect 1065 903 1069 907
rect 1054 878 1058 882
rect 1030 868 1034 872
rect 1014 748 1018 752
rect 1062 848 1066 852
rect 1150 898 1154 902
rect 1126 868 1130 872
rect 1086 808 1090 812
rect 1102 788 1106 792
rect 1062 748 1066 752
rect 1014 738 1018 742
rect 1006 728 1010 732
rect 950 688 954 692
rect 982 678 986 682
rect 734 658 738 662
rect 934 658 938 662
rect 790 648 794 652
rect 902 648 906 652
rect 782 638 786 642
rect 918 638 922 642
rect 950 658 954 662
rect 966 648 970 652
rect 1006 638 1010 642
rect 942 588 946 592
rect 838 578 842 582
rect 886 578 890 582
rect 734 568 738 572
rect 750 568 754 572
rect 870 568 874 572
rect 798 548 802 552
rect 846 548 850 552
rect 902 568 906 572
rect 942 558 946 562
rect 886 548 890 552
rect 862 538 866 542
rect 926 538 930 542
rect 798 478 802 482
rect 910 518 914 522
rect 862 488 866 492
rect 878 478 882 482
rect 902 478 906 482
rect 726 468 730 472
rect 822 468 826 472
rect 838 468 842 472
rect 582 448 586 452
rect 614 448 618 452
rect 546 403 550 407
rect 553 403 557 407
rect 662 378 666 382
rect 694 378 698 382
rect 622 358 626 362
rect 638 358 642 362
rect 342 348 346 352
rect 358 348 362 352
rect 374 348 378 352
rect 406 348 410 352
rect 382 338 386 342
rect 254 318 258 322
rect 310 318 314 322
rect 262 308 266 312
rect 206 288 210 292
rect 278 288 282 292
rect 326 328 330 332
rect 318 288 322 292
rect 166 258 170 262
rect 214 258 218 262
rect 246 258 250 262
rect 182 188 186 192
rect 190 168 194 172
rect 142 158 146 162
rect 174 158 178 162
rect 182 138 186 142
rect 190 138 194 142
rect 198 138 202 142
rect 126 128 130 132
rect 134 128 138 132
rect 6 78 10 82
rect 86 68 90 72
rect 238 138 242 142
rect 206 88 210 92
rect 294 278 298 282
rect 342 318 346 322
rect 326 278 330 282
rect 334 138 338 142
rect 302 118 306 122
rect 294 88 298 92
rect 358 298 362 302
rect 390 298 394 302
rect 414 298 418 302
rect 614 348 618 352
rect 446 318 450 322
rect 454 298 458 302
rect 374 288 378 292
rect 422 288 426 292
rect 438 288 442 292
rect 462 288 466 292
rect 350 258 354 262
rect 478 278 482 282
rect 486 278 490 282
rect 390 268 394 272
rect 422 268 426 272
rect 598 328 602 332
rect 614 328 618 332
rect 534 318 538 322
rect 582 318 586 322
rect 614 268 618 272
rect 478 258 482 262
rect 606 258 610 262
rect 630 348 634 352
rect 638 338 642 342
rect 478 248 482 252
rect 502 248 506 252
rect 526 248 530 252
rect 422 228 426 232
rect 502 228 506 232
rect 414 178 418 182
rect 350 138 354 142
rect 374 138 378 142
rect 374 118 378 122
rect 398 138 402 142
rect 382 88 386 92
rect 546 203 550 207
rect 553 203 557 207
rect 526 178 530 182
rect 574 178 578 182
rect 582 148 586 152
rect 614 238 618 242
rect 646 318 650 322
rect 662 268 666 272
rect 694 338 698 342
rect 782 448 786 452
rect 718 378 722 382
rect 734 368 738 372
rect 718 348 722 352
rect 766 358 770 362
rect 798 358 802 362
rect 830 458 834 462
rect 846 458 850 462
rect 854 448 858 452
rect 822 438 826 442
rect 838 408 842 412
rect 822 368 826 372
rect 862 398 866 402
rect 870 368 874 372
rect 814 338 818 342
rect 838 338 842 342
rect 702 318 706 322
rect 734 288 738 292
rect 790 278 794 282
rect 718 268 722 272
rect 830 268 834 272
rect 678 248 682 252
rect 694 248 698 252
rect 670 218 674 222
rect 750 218 754 222
rect 638 208 642 212
rect 862 278 866 282
rect 870 278 874 282
rect 846 248 850 252
rect 678 188 682 192
rect 806 188 810 192
rect 830 188 834 192
rect 630 168 634 172
rect 734 168 738 172
rect 742 168 746 172
rect 622 158 626 162
rect 614 148 618 152
rect 590 138 594 142
rect 606 138 610 142
rect 502 118 506 122
rect 422 78 426 82
rect 254 68 258 72
rect 318 68 322 72
rect 350 68 354 72
rect 382 68 386 72
rect 406 68 410 72
rect 494 68 498 72
rect 94 58 98 62
rect 310 58 314 62
rect 326 58 330 62
rect 278 48 282 52
rect 350 48 354 52
rect 614 128 618 132
rect 558 88 562 92
rect 558 68 562 72
rect 734 158 738 162
rect 862 188 866 192
rect 1118 748 1122 752
rect 1142 748 1146 752
rect 1102 728 1106 732
rect 1046 718 1050 722
rect 1086 718 1090 722
rect 1030 648 1034 652
rect 1038 618 1042 622
rect 1030 608 1034 612
rect 1022 568 1026 572
rect 1022 538 1026 542
rect 982 498 986 502
rect 990 488 994 492
rect 990 468 994 472
rect 1006 468 1010 472
rect 982 458 986 462
rect 926 438 930 442
rect 926 428 930 432
rect 958 358 962 362
rect 886 338 890 342
rect 926 338 930 342
rect 918 308 922 312
rect 894 268 898 272
rect 950 308 954 312
rect 942 278 946 282
rect 934 248 938 252
rect 854 168 858 172
rect 838 158 842 162
rect 662 138 666 142
rect 654 108 658 112
rect 646 78 650 82
rect 766 98 770 102
rect 814 98 818 102
rect 662 88 666 92
rect 710 88 714 92
rect 798 88 802 92
rect 726 78 730 82
rect 878 168 882 172
rect 918 158 922 162
rect 934 168 938 172
rect 934 158 938 162
rect 974 338 978 342
rect 1058 703 1062 707
rect 1065 703 1069 707
rect 1134 698 1138 702
rect 1070 688 1074 692
rect 1062 668 1066 672
rect 1094 658 1098 662
rect 1110 658 1114 662
rect 1078 638 1082 642
rect 1046 578 1050 582
rect 1142 668 1146 672
rect 1126 638 1130 642
rect 1134 568 1138 572
rect 1118 558 1122 562
rect 1086 548 1090 552
rect 1102 548 1106 552
rect 1110 548 1114 552
rect 1126 548 1130 552
rect 1038 528 1042 532
rect 1038 498 1042 502
rect 1030 458 1034 462
rect 1094 508 1098 512
rect 1058 503 1062 507
rect 1065 503 1069 507
rect 1174 1108 1178 1112
rect 1246 1158 1250 1162
rect 1278 1278 1282 1282
rect 1294 1308 1298 1312
rect 1310 1538 1314 1542
rect 1334 1528 1338 1532
rect 1366 1518 1370 1522
rect 1486 1758 1490 1762
rect 1470 1748 1474 1752
rect 1502 1748 1506 1752
rect 1526 1748 1530 1752
rect 1606 1748 1610 1752
rect 1454 1738 1458 1742
rect 1462 1698 1466 1702
rect 1430 1678 1434 1682
rect 1446 1668 1450 1672
rect 1438 1658 1442 1662
rect 1430 1648 1434 1652
rect 1414 1618 1418 1622
rect 1398 1598 1402 1602
rect 1382 1498 1386 1502
rect 1422 1568 1426 1572
rect 1422 1548 1426 1552
rect 1446 1628 1450 1632
rect 1486 1738 1490 1742
rect 1478 1728 1482 1732
rect 1502 1728 1506 1732
rect 1526 1728 1530 1732
rect 1526 1688 1530 1692
rect 1494 1678 1498 1682
rect 1590 1718 1594 1722
rect 1582 1698 1586 1702
rect 1542 1668 1546 1672
rect 1478 1658 1482 1662
rect 1502 1658 1506 1662
rect 1542 1658 1546 1662
rect 1566 1658 1570 1662
rect 1478 1638 1482 1642
rect 1526 1648 1530 1652
rect 1518 1618 1522 1622
rect 1446 1568 1450 1572
rect 1470 1568 1474 1572
rect 1486 1568 1490 1572
rect 1454 1558 1458 1562
rect 1470 1558 1474 1562
rect 1494 1558 1498 1562
rect 1502 1548 1506 1552
rect 1438 1528 1442 1532
rect 1414 1518 1418 1522
rect 1334 1488 1338 1492
rect 1318 1478 1322 1482
rect 1326 1468 1330 1472
rect 1342 1468 1346 1472
rect 1406 1468 1410 1472
rect 1358 1458 1362 1462
rect 1350 1448 1354 1452
rect 1342 1418 1346 1422
rect 1318 1398 1322 1402
rect 1358 1408 1362 1412
rect 1390 1438 1394 1442
rect 1382 1408 1386 1412
rect 1374 1388 1378 1392
rect 1398 1378 1402 1382
rect 1438 1508 1442 1512
rect 1494 1508 1498 1512
rect 1422 1458 1426 1462
rect 1430 1448 1434 1452
rect 1422 1438 1426 1442
rect 1430 1428 1434 1432
rect 1462 1478 1466 1482
rect 1478 1478 1482 1482
rect 1454 1468 1458 1472
rect 1446 1458 1450 1462
rect 1406 1368 1410 1372
rect 1366 1348 1370 1352
rect 1358 1338 1362 1342
rect 1382 1338 1386 1342
rect 1454 1398 1458 1402
rect 1470 1448 1474 1452
rect 1486 1448 1490 1452
rect 1478 1388 1482 1392
rect 1454 1368 1458 1372
rect 1446 1348 1450 1352
rect 1510 1438 1514 1442
rect 1494 1408 1498 1412
rect 1502 1388 1506 1392
rect 1486 1358 1490 1362
rect 1534 1628 1538 1632
rect 1562 1603 1566 1607
rect 1569 1603 1573 1607
rect 1550 1578 1554 1582
rect 1574 1568 1578 1572
rect 1534 1508 1538 1512
rect 1518 1418 1522 1422
rect 1510 1368 1514 1372
rect 1470 1348 1474 1352
rect 1614 1688 1618 1692
rect 1678 1748 1682 1752
rect 1686 1658 1690 1662
rect 1598 1648 1602 1652
rect 1622 1628 1626 1632
rect 1638 1648 1642 1652
rect 1662 1628 1666 1632
rect 1630 1598 1634 1602
rect 1590 1588 1594 1592
rect 1654 1578 1658 1582
rect 1646 1558 1650 1562
rect 1598 1547 1602 1551
rect 1670 1548 1674 1552
rect 1670 1538 1674 1542
rect 1598 1518 1602 1522
rect 1582 1508 1586 1512
rect 1646 1528 1650 1532
rect 1542 1478 1546 1482
rect 1622 1478 1626 1482
rect 1694 1648 1698 1652
rect 1694 1608 1698 1612
rect 1686 1558 1690 1562
rect 1718 1828 1722 1832
rect 1710 1768 1714 1772
rect 1758 1818 1762 1822
rect 1710 1738 1714 1742
rect 1718 1688 1722 1692
rect 1766 1808 1770 1812
rect 1758 1738 1762 1742
rect 1774 1728 1778 1732
rect 1750 1718 1754 1722
rect 1750 1688 1754 1692
rect 1814 1808 1818 1812
rect 1854 1898 1858 1902
rect 1854 1868 1858 1872
rect 1846 1798 1850 1802
rect 1854 1788 1858 1792
rect 1870 1898 1874 1902
rect 2030 2088 2034 2092
rect 1990 2068 1994 2072
rect 2070 2278 2074 2282
rect 2206 2328 2210 2332
rect 2150 2288 2154 2292
rect 2214 2298 2218 2302
rect 2238 2298 2242 2302
rect 2142 2268 2146 2272
rect 2086 2258 2090 2262
rect 2142 2258 2146 2262
rect 2126 2158 2130 2162
rect 2158 2258 2162 2262
rect 2054 2128 2058 2132
rect 2070 2118 2074 2122
rect 2086 2118 2090 2122
rect 2134 2118 2138 2122
rect 2022 2058 2026 2062
rect 2054 2058 2058 2062
rect 2006 2048 2010 2052
rect 1990 2028 1994 2032
rect 1974 1998 1978 2002
rect 1990 1998 1994 2002
rect 1950 1988 1954 1992
rect 1902 1948 1906 1952
rect 1974 1948 1978 1952
rect 1966 1928 1970 1932
rect 1926 1898 1930 1902
rect 1886 1848 1890 1852
rect 1862 1758 1866 1762
rect 1830 1748 1834 1752
rect 1870 1748 1874 1752
rect 1822 1728 1826 1732
rect 1798 1698 1802 1702
rect 1782 1688 1786 1692
rect 1798 1688 1802 1692
rect 1822 1708 1826 1712
rect 1846 1708 1850 1712
rect 1878 1678 1882 1682
rect 1742 1658 1746 1662
rect 1718 1648 1722 1652
rect 1766 1648 1770 1652
rect 1774 1648 1778 1652
rect 1710 1588 1714 1592
rect 1766 1588 1770 1592
rect 1830 1668 1834 1672
rect 1862 1668 1866 1672
rect 1870 1668 1874 1672
rect 1806 1648 1810 1652
rect 1814 1628 1818 1632
rect 1814 1608 1818 1612
rect 1822 1608 1826 1612
rect 1790 1578 1794 1582
rect 1726 1558 1730 1562
rect 1710 1548 1714 1552
rect 1894 1808 1898 1812
rect 1918 1758 1922 1762
rect 2006 1948 2010 1952
rect 2082 2103 2086 2107
rect 2089 2103 2093 2107
rect 2110 2098 2114 2102
rect 2118 2078 2122 2082
rect 2102 1988 2106 1992
rect 2086 1958 2090 1962
rect 2070 1948 2074 1952
rect 2022 1928 2026 1932
rect 2014 1918 2018 1922
rect 2030 1918 2034 1922
rect 2006 1868 2010 1872
rect 2082 1903 2086 1907
rect 2089 1903 2093 1907
rect 2062 1878 2066 1882
rect 2038 1868 2042 1872
rect 2126 2048 2130 2052
rect 2118 1968 2122 1972
rect 2118 1918 2122 1922
rect 2166 2218 2170 2222
rect 2270 2328 2274 2332
rect 2414 2368 2418 2372
rect 2430 2368 2434 2372
rect 2334 2318 2338 2322
rect 2318 2278 2322 2282
rect 2342 2268 2346 2272
rect 2366 2268 2370 2272
rect 2350 2248 2354 2252
rect 2366 2248 2370 2252
rect 2238 2218 2242 2222
rect 2254 2188 2258 2192
rect 2206 2178 2210 2182
rect 2182 2168 2186 2172
rect 2278 2188 2282 2192
rect 2262 2168 2266 2172
rect 2174 2148 2178 2152
rect 2310 2148 2314 2152
rect 2198 2138 2202 2142
rect 2222 2138 2226 2142
rect 2198 2108 2202 2112
rect 2214 2078 2218 2082
rect 2142 2058 2146 2062
rect 2158 2058 2162 2062
rect 2174 2058 2178 2062
rect 2182 2058 2186 2062
rect 2214 2058 2218 2062
rect 2190 2008 2194 2012
rect 2182 1968 2186 1972
rect 2142 1958 2146 1962
rect 2174 1958 2178 1962
rect 2150 1948 2154 1952
rect 2230 2068 2234 2072
rect 2238 2058 2242 2062
rect 2246 2028 2250 2032
rect 2342 2148 2346 2152
rect 2326 2138 2330 2142
rect 2358 2128 2362 2132
rect 2270 2118 2274 2122
rect 2406 2278 2410 2282
rect 2438 2348 2442 2352
rect 2478 2348 2482 2352
rect 2534 2338 2538 2342
rect 2518 2328 2522 2332
rect 2430 2278 2434 2282
rect 2494 2278 2498 2282
rect 2462 2268 2466 2272
rect 2414 2258 2418 2262
rect 2382 2248 2386 2252
rect 2438 2248 2442 2252
rect 2454 2248 2458 2252
rect 2438 2158 2442 2162
rect 2390 2138 2394 2142
rect 2414 2118 2418 2122
rect 2286 2098 2290 2102
rect 2262 2088 2266 2092
rect 2294 2088 2298 2092
rect 2286 2078 2290 2082
rect 2302 2068 2306 2072
rect 2262 2058 2266 2062
rect 2270 2058 2274 2062
rect 2342 2058 2346 2062
rect 2270 1998 2274 2002
rect 2302 1998 2306 2002
rect 2238 1978 2242 1982
rect 2254 1978 2258 1982
rect 2246 1968 2250 1972
rect 2190 1938 2194 1942
rect 2150 1868 2154 1872
rect 2022 1858 2026 1862
rect 2134 1858 2138 1862
rect 2182 1858 2186 1862
rect 1958 1808 1962 1812
rect 1974 1788 1978 1792
rect 1942 1768 1946 1772
rect 1950 1768 1954 1772
rect 1990 1758 1994 1762
rect 1902 1748 1906 1752
rect 1974 1748 1978 1752
rect 1990 1728 1994 1732
rect 1894 1688 1898 1692
rect 1926 1688 1930 1692
rect 1894 1658 1898 1662
rect 2030 1848 2034 1852
rect 2094 1818 2098 1822
rect 2134 1808 2138 1812
rect 2054 1778 2058 1782
rect 2110 1778 2114 1782
rect 2062 1768 2066 1772
rect 2070 1758 2074 1762
rect 2118 1738 2122 1742
rect 2142 1788 2146 1792
rect 2142 1748 2146 1752
rect 2190 1788 2194 1792
rect 2094 1728 2098 1732
rect 2110 1728 2114 1732
rect 2142 1728 2146 1732
rect 2182 1728 2186 1732
rect 2062 1718 2066 1722
rect 2070 1718 2074 1722
rect 2022 1708 2026 1712
rect 2082 1703 2086 1707
rect 2089 1703 2093 1707
rect 1966 1688 1970 1692
rect 1966 1678 1970 1682
rect 2054 1678 2058 1682
rect 2166 1698 2170 1702
rect 2134 1688 2138 1692
rect 2150 1678 2154 1682
rect 1998 1668 2002 1672
rect 2038 1668 2042 1672
rect 2102 1668 2106 1672
rect 2118 1668 2122 1672
rect 1950 1658 1954 1662
rect 1942 1648 1946 1652
rect 1950 1648 1954 1652
rect 1934 1628 1938 1632
rect 1966 1628 1970 1632
rect 1886 1598 1890 1602
rect 1926 1588 1930 1592
rect 2014 1658 2018 1662
rect 2166 1658 2170 1662
rect 2006 1648 2010 1652
rect 1998 1638 2002 1642
rect 2110 1638 2114 1642
rect 2118 1638 2122 1642
rect 1990 1618 1994 1622
rect 2014 1588 2018 1592
rect 1934 1578 1938 1582
rect 1958 1578 1962 1582
rect 1862 1568 1866 1572
rect 1950 1568 1954 1572
rect 1766 1548 1770 1552
rect 1870 1548 1874 1552
rect 1942 1548 1946 1552
rect 1742 1538 1746 1542
rect 1702 1518 1706 1522
rect 1686 1488 1690 1492
rect 1694 1488 1698 1492
rect 1590 1468 1594 1472
rect 1606 1468 1610 1472
rect 1614 1468 1618 1472
rect 1678 1468 1682 1472
rect 1582 1448 1586 1452
rect 1590 1448 1594 1452
rect 1542 1418 1546 1422
rect 1562 1403 1566 1407
rect 1569 1403 1573 1407
rect 1550 1398 1554 1402
rect 1550 1378 1554 1382
rect 1558 1378 1562 1382
rect 1550 1348 1554 1352
rect 1494 1338 1498 1342
rect 1526 1338 1530 1342
rect 1398 1328 1402 1332
rect 1430 1328 1434 1332
rect 1430 1318 1434 1322
rect 1310 1288 1314 1292
rect 1326 1278 1330 1282
rect 1302 1268 1306 1272
rect 1278 1248 1282 1252
rect 1294 1248 1298 1252
rect 1310 1238 1314 1242
rect 1262 1178 1266 1182
rect 1294 1158 1298 1162
rect 1254 1138 1258 1142
rect 1278 1148 1282 1152
rect 1278 1138 1282 1142
rect 1286 1108 1290 1112
rect 1246 1058 1250 1062
rect 1262 1048 1266 1052
rect 1254 1018 1258 1022
rect 1246 1008 1250 1012
rect 1174 998 1178 1002
rect 1238 968 1242 972
rect 1182 938 1186 942
rect 1270 1038 1274 1042
rect 1262 968 1266 972
rect 1278 998 1282 1002
rect 1198 928 1202 932
rect 1190 918 1194 922
rect 1198 908 1202 912
rect 1238 888 1242 892
rect 1214 868 1218 872
rect 1334 1188 1338 1192
rect 1326 1158 1330 1162
rect 1318 1148 1322 1152
rect 1326 1148 1330 1152
rect 1358 1258 1362 1262
rect 1366 1188 1370 1192
rect 1350 1168 1354 1172
rect 1366 1168 1370 1172
rect 1374 1148 1378 1152
rect 1382 1098 1386 1102
rect 1326 1068 1330 1072
rect 1342 1068 1346 1072
rect 1318 1058 1322 1062
rect 1382 1058 1386 1062
rect 1350 1048 1354 1052
rect 1318 1038 1322 1042
rect 1374 1038 1378 1042
rect 1302 1008 1306 1012
rect 1310 1008 1314 1012
rect 1294 988 1298 992
rect 1286 978 1290 982
rect 1286 958 1290 962
rect 1246 868 1250 872
rect 1286 868 1290 872
rect 1198 858 1202 862
rect 1214 858 1218 862
rect 1302 918 1306 922
rect 1294 848 1298 852
rect 1270 798 1274 802
rect 1286 768 1290 772
rect 1246 738 1250 742
rect 1190 728 1194 732
rect 1270 728 1274 732
rect 1294 688 1298 692
rect 1286 678 1290 682
rect 1214 668 1218 672
rect 1254 668 1258 672
rect 1270 668 1274 672
rect 1174 658 1178 662
rect 1150 538 1154 542
rect 1126 528 1130 532
rect 1118 448 1122 452
rect 1102 438 1106 442
rect 1118 438 1122 442
rect 1102 368 1106 372
rect 1046 358 1050 362
rect 1014 348 1018 352
rect 974 288 978 292
rect 966 188 970 192
rect 1046 338 1050 342
rect 1030 328 1034 332
rect 1058 303 1062 307
rect 1065 303 1069 307
rect 958 148 962 152
rect 910 98 914 102
rect 1046 258 1050 262
rect 1022 248 1026 252
rect 1038 248 1042 252
rect 1014 198 1018 202
rect 1006 178 1010 182
rect 1006 168 1010 172
rect 990 148 994 152
rect 974 118 978 122
rect 982 118 986 122
rect 934 108 938 112
rect 926 88 930 92
rect 958 88 962 92
rect 974 78 978 82
rect 686 68 690 72
rect 742 68 746 72
rect 878 68 882 72
rect 934 68 938 72
rect 1014 68 1018 72
rect 1182 648 1186 652
rect 1214 638 1218 642
rect 1262 658 1266 662
rect 1302 658 1306 662
rect 1246 638 1250 642
rect 1230 628 1234 632
rect 1262 628 1266 632
rect 1326 978 1330 982
rect 1374 978 1378 982
rect 1342 968 1346 972
rect 1414 1288 1418 1292
rect 1478 1328 1482 1332
rect 1494 1328 1498 1332
rect 1446 1308 1450 1312
rect 1462 1288 1466 1292
rect 1478 1288 1482 1292
rect 1422 1278 1426 1282
rect 1446 1278 1450 1282
rect 1454 1278 1458 1282
rect 1438 1258 1442 1262
rect 1438 1168 1442 1172
rect 1550 1288 1554 1292
rect 1542 1278 1546 1282
rect 1502 1268 1506 1272
rect 1518 1268 1522 1272
rect 1598 1428 1602 1432
rect 1566 1328 1570 1332
rect 1574 1298 1578 1302
rect 1630 1458 1634 1462
rect 1622 1438 1626 1442
rect 1734 1528 1738 1532
rect 1750 1528 1754 1532
rect 1814 1498 1818 1502
rect 1726 1438 1730 1442
rect 1710 1428 1714 1432
rect 1614 1418 1618 1422
rect 1654 1388 1658 1392
rect 1646 1358 1650 1362
rect 1638 1348 1642 1352
rect 1606 1328 1610 1332
rect 1622 1328 1626 1332
rect 1590 1308 1594 1312
rect 1582 1288 1586 1292
rect 1574 1268 1578 1272
rect 1462 1258 1466 1262
rect 1582 1258 1586 1262
rect 1470 1228 1474 1232
rect 1478 1188 1482 1192
rect 1542 1248 1546 1252
rect 1494 1178 1498 1182
rect 1542 1178 1546 1182
rect 1518 1168 1522 1172
rect 1494 1148 1498 1152
rect 1502 1148 1506 1152
rect 1414 1138 1418 1142
rect 1438 1138 1442 1142
rect 1446 1138 1450 1142
rect 1398 1128 1402 1132
rect 1438 1118 1442 1122
rect 1446 1068 1450 1072
rect 1470 1128 1474 1132
rect 1502 1118 1506 1122
rect 1486 1078 1490 1082
rect 1430 1048 1434 1052
rect 1446 1048 1450 1052
rect 1454 1028 1458 1032
rect 1454 998 1458 1002
rect 1414 978 1418 982
rect 1390 958 1394 962
rect 1414 958 1418 962
rect 1390 948 1394 952
rect 1398 938 1402 942
rect 1382 928 1386 932
rect 1382 898 1386 902
rect 1358 888 1362 892
rect 1350 878 1354 882
rect 1374 868 1378 872
rect 1438 948 1442 952
rect 1430 908 1434 912
rect 1446 878 1450 882
rect 1494 1018 1498 1022
rect 1526 1108 1530 1112
rect 1542 1008 1546 1012
rect 1510 998 1514 1002
rect 1502 968 1506 972
rect 1510 968 1514 972
rect 1562 1203 1566 1207
rect 1569 1203 1573 1207
rect 1558 1168 1562 1172
rect 1566 1158 1570 1162
rect 1558 1048 1562 1052
rect 1574 1018 1578 1022
rect 1562 1003 1566 1007
rect 1569 1003 1573 1007
rect 1542 958 1546 962
rect 1606 1308 1610 1312
rect 1630 1288 1634 1292
rect 1686 1408 1690 1412
rect 1678 1388 1682 1392
rect 1662 1348 1666 1352
rect 1662 1338 1666 1342
rect 1718 1338 1722 1342
rect 1670 1328 1674 1332
rect 1670 1308 1674 1312
rect 1646 1298 1650 1302
rect 1654 1288 1658 1292
rect 1702 1288 1706 1292
rect 1694 1278 1698 1282
rect 1646 1268 1650 1272
rect 1654 1268 1658 1272
rect 1638 1258 1642 1262
rect 1598 1238 1602 1242
rect 1606 1228 1610 1232
rect 1622 1168 1626 1172
rect 1614 1158 1618 1162
rect 1598 1138 1602 1142
rect 1622 1108 1626 1112
rect 1606 1068 1610 1072
rect 1598 1058 1602 1062
rect 1590 1038 1594 1042
rect 1598 958 1602 962
rect 1502 948 1506 952
rect 1526 948 1530 952
rect 1566 948 1570 952
rect 1574 948 1578 952
rect 1510 938 1514 942
rect 1486 928 1490 932
rect 1478 918 1482 922
rect 1462 878 1466 882
rect 1470 868 1474 872
rect 1358 858 1362 862
rect 1382 858 1386 862
rect 1390 858 1394 862
rect 1438 858 1442 862
rect 1342 748 1346 752
rect 1334 728 1338 732
rect 1318 688 1322 692
rect 1318 668 1322 672
rect 1366 668 1370 672
rect 1374 668 1378 672
rect 1390 838 1394 842
rect 1422 838 1426 842
rect 1414 818 1418 822
rect 1414 808 1418 812
rect 1390 758 1394 762
rect 1414 758 1418 762
rect 1422 758 1426 762
rect 1398 748 1402 752
rect 1422 728 1426 732
rect 1422 698 1426 702
rect 1334 658 1338 662
rect 1382 658 1386 662
rect 1310 608 1314 612
rect 1366 608 1370 612
rect 1414 648 1418 652
rect 1390 598 1394 602
rect 1430 588 1434 592
rect 1286 578 1290 582
rect 1398 578 1402 582
rect 1302 568 1306 572
rect 1342 568 1346 572
rect 1390 568 1394 572
rect 1326 558 1330 562
rect 1174 548 1178 552
rect 1238 548 1242 552
rect 1310 548 1314 552
rect 1166 508 1170 512
rect 1174 468 1178 472
rect 1158 398 1162 402
rect 1206 508 1210 512
rect 1190 378 1194 382
rect 1182 368 1186 372
rect 1174 358 1178 362
rect 1174 338 1178 342
rect 1254 498 1258 502
rect 1318 488 1322 492
rect 1286 478 1290 482
rect 1230 458 1234 462
rect 1238 448 1242 452
rect 1286 458 1290 462
rect 1262 448 1266 452
rect 1278 448 1282 452
rect 1246 438 1250 442
rect 1230 418 1234 422
rect 1262 418 1266 422
rect 1230 388 1234 392
rect 1142 288 1146 292
rect 1166 278 1170 282
rect 1182 268 1186 272
rect 1318 438 1322 442
rect 1334 438 1338 442
rect 1326 428 1330 432
rect 1382 558 1386 562
rect 1446 838 1450 842
rect 1558 938 1562 942
rect 1518 928 1522 932
rect 1494 878 1498 882
rect 1478 788 1482 792
rect 1462 778 1466 782
rect 1502 778 1506 782
rect 1678 1258 1682 1262
rect 1686 1248 1690 1252
rect 1678 1138 1682 1142
rect 1710 1278 1714 1282
rect 1710 1248 1714 1252
rect 1710 1228 1714 1232
rect 1630 1078 1634 1082
rect 1646 1078 1650 1082
rect 1678 1078 1682 1082
rect 1638 1068 1642 1072
rect 1630 1058 1634 1062
rect 1646 1058 1650 1062
rect 1662 1058 1666 1062
rect 1670 1048 1674 1052
rect 1686 1048 1690 1052
rect 1694 1048 1698 1052
rect 1718 1038 1722 1042
rect 1702 1008 1706 1012
rect 1734 1368 1738 1372
rect 1790 1458 1794 1462
rect 2022 1578 2026 1582
rect 2014 1558 2018 1562
rect 2054 1558 2058 1562
rect 2078 1558 2082 1562
rect 1966 1548 1970 1552
rect 2006 1548 2010 1552
rect 2030 1548 2034 1552
rect 2070 1548 2074 1552
rect 1870 1518 1874 1522
rect 1918 1518 1922 1522
rect 1870 1498 1874 1502
rect 1830 1488 1834 1492
rect 1926 1508 1930 1512
rect 1918 1478 1922 1482
rect 1926 1478 1930 1482
rect 1822 1448 1826 1452
rect 1774 1428 1778 1432
rect 1750 1418 1754 1422
rect 1790 1418 1794 1422
rect 1854 1458 1858 1462
rect 1830 1408 1834 1412
rect 1790 1398 1794 1402
rect 1782 1358 1786 1362
rect 1822 1378 1826 1382
rect 1758 1308 1762 1312
rect 1814 1318 1818 1322
rect 1806 1308 1810 1312
rect 1806 1278 1810 1282
rect 1782 1258 1786 1262
rect 1798 1258 1802 1262
rect 1806 1258 1810 1262
rect 1766 1238 1770 1242
rect 1742 1098 1746 1102
rect 1774 1088 1778 1092
rect 1790 1078 1794 1082
rect 1838 1368 1842 1372
rect 1838 1358 1842 1362
rect 1870 1308 1874 1312
rect 1902 1308 1906 1312
rect 1926 1459 1930 1463
rect 1934 1448 1938 1452
rect 2014 1528 2018 1532
rect 1990 1498 1994 1502
rect 1998 1468 2002 1472
rect 2038 1528 2042 1532
rect 2134 1628 2138 1632
rect 2150 1568 2154 1572
rect 2158 1558 2162 1562
rect 2214 1858 2218 1862
rect 2206 1758 2210 1762
rect 2198 1718 2202 1722
rect 2302 1948 2306 1952
rect 2270 1938 2274 1942
rect 2254 1908 2258 1912
rect 2238 1768 2242 1772
rect 2262 1748 2266 1752
rect 2230 1738 2234 1742
rect 2222 1688 2226 1692
rect 2206 1668 2210 1672
rect 2230 1648 2234 1652
rect 2246 1738 2250 1742
rect 2326 1898 2330 1902
rect 2294 1868 2298 1872
rect 2318 1868 2322 1872
rect 2334 1878 2338 1882
rect 2334 1848 2338 1852
rect 2286 1838 2290 1842
rect 2270 1718 2274 1722
rect 2246 1668 2250 1672
rect 2214 1618 2218 1622
rect 2222 1618 2226 1622
rect 2206 1568 2210 1572
rect 2238 1558 2242 1562
rect 2262 1628 2266 1632
rect 2270 1628 2274 1632
rect 2262 1618 2266 1622
rect 2278 1568 2282 1572
rect 2254 1558 2258 1562
rect 2086 1528 2090 1532
rect 2142 1528 2146 1532
rect 2174 1528 2178 1532
rect 2082 1503 2086 1507
rect 2089 1503 2093 1507
rect 2046 1488 2050 1492
rect 2070 1478 2074 1482
rect 2038 1468 2042 1472
rect 2046 1468 2050 1472
rect 1982 1458 1986 1462
rect 2046 1458 2050 1462
rect 2102 1458 2106 1462
rect 1974 1448 1978 1452
rect 2006 1448 2010 1452
rect 1966 1438 1970 1442
rect 1966 1408 1970 1412
rect 1982 1408 1986 1412
rect 1950 1398 1954 1402
rect 1934 1358 1938 1362
rect 1942 1358 1946 1362
rect 1998 1358 2002 1362
rect 2030 1448 2034 1452
rect 2038 1448 2042 1452
rect 2094 1448 2098 1452
rect 2062 1418 2066 1422
rect 2062 1408 2066 1412
rect 2078 1388 2082 1392
rect 2118 1408 2122 1412
rect 2110 1398 2114 1402
rect 2102 1368 2106 1372
rect 2110 1368 2114 1372
rect 2070 1358 2074 1362
rect 2174 1478 2178 1482
rect 2246 1518 2250 1522
rect 2262 1518 2266 1522
rect 2238 1508 2242 1512
rect 2254 1508 2258 1512
rect 2150 1468 2154 1472
rect 2190 1448 2194 1452
rect 2190 1408 2194 1412
rect 2126 1358 2130 1362
rect 2158 1358 2162 1362
rect 2174 1358 2178 1362
rect 2206 1358 2210 1362
rect 2014 1348 2018 1352
rect 2022 1348 2026 1352
rect 2054 1348 2058 1352
rect 2126 1348 2130 1352
rect 2198 1348 2202 1352
rect 1942 1328 1946 1332
rect 1974 1328 1978 1332
rect 1822 1288 1826 1292
rect 1942 1278 1946 1282
rect 1830 1268 1834 1272
rect 1838 1268 1842 1272
rect 1846 1268 1850 1272
rect 1910 1268 1914 1272
rect 1822 1208 1826 1212
rect 1854 1238 1858 1242
rect 1854 1218 1858 1222
rect 1958 1258 1962 1262
rect 2022 1338 2026 1342
rect 2086 1338 2090 1342
rect 2142 1338 2146 1342
rect 2254 1468 2258 1472
rect 2270 1508 2274 1512
rect 2278 1498 2282 1502
rect 2342 1808 2346 1812
rect 2302 1788 2306 1792
rect 2294 1778 2298 1782
rect 2334 1768 2338 1772
rect 2318 1758 2322 1762
rect 2478 2158 2482 2162
rect 2406 2098 2410 2102
rect 2462 2098 2466 2102
rect 2382 2078 2386 2082
rect 2438 2058 2442 2062
rect 2398 2048 2402 2052
rect 2462 1988 2466 1992
rect 2374 1948 2378 1952
rect 2462 1948 2466 1952
rect 2406 1918 2410 1922
rect 2534 2278 2538 2282
rect 2542 2268 2546 2272
rect 2534 2248 2538 2252
rect 2622 2328 2626 2332
rect 2558 2318 2562 2322
rect 2566 2268 2570 2272
rect 2614 2268 2618 2272
rect 2558 2218 2562 2222
rect 2550 2168 2554 2172
rect 2526 2108 2530 2112
rect 2590 2148 2594 2152
rect 2622 2148 2626 2152
rect 2590 2108 2594 2112
rect 2614 2108 2618 2112
rect 2558 2068 2562 2072
rect 2510 2058 2514 2062
rect 2502 1968 2506 1972
rect 2478 1958 2482 1962
rect 2502 1948 2506 1952
rect 2430 1938 2434 1942
rect 2454 1938 2458 1942
rect 2574 1938 2578 1942
rect 2430 1928 2434 1932
rect 2366 1868 2370 1872
rect 2382 1868 2386 1872
rect 2398 1858 2402 1862
rect 2374 1848 2378 1852
rect 2430 1908 2434 1912
rect 2534 1918 2538 1922
rect 2510 1898 2514 1902
rect 2518 1878 2522 1882
rect 2614 1928 2618 1932
rect 2614 1918 2618 1922
rect 2438 1868 2442 1872
rect 2598 1868 2602 1872
rect 2438 1858 2442 1862
rect 2430 1848 2434 1852
rect 2494 1848 2498 1852
rect 2646 1918 2650 1922
rect 2606 1838 2610 1842
rect 2622 1838 2626 1842
rect 2414 1828 2418 1832
rect 2374 1808 2378 1812
rect 2494 1798 2498 1802
rect 2302 1748 2306 1752
rect 2310 1738 2314 1742
rect 2366 1748 2370 1752
rect 2350 1728 2354 1732
rect 2358 1728 2362 1732
rect 2342 1718 2346 1722
rect 2342 1698 2346 1702
rect 2310 1688 2314 1692
rect 2318 1658 2322 1662
rect 2294 1638 2298 1642
rect 2462 1758 2466 1762
rect 2486 1758 2490 1762
rect 2430 1748 2434 1752
rect 2438 1738 2442 1742
rect 2374 1718 2378 1722
rect 2446 1718 2450 1722
rect 2438 1708 2442 1712
rect 2446 1708 2450 1712
rect 2406 1688 2410 1692
rect 2382 1678 2386 1682
rect 2390 1668 2394 1672
rect 2422 1668 2426 1672
rect 2446 1698 2450 1702
rect 2478 1748 2482 1752
rect 2494 1738 2498 1742
rect 2510 1708 2514 1712
rect 2470 1678 2474 1682
rect 2558 1748 2562 1752
rect 2638 1778 2642 1782
rect 2590 1688 2594 1692
rect 2430 1658 2434 1662
rect 2518 1658 2522 1662
rect 2350 1648 2354 1652
rect 2302 1598 2306 1602
rect 2310 1578 2314 1582
rect 2302 1558 2306 1562
rect 2350 1558 2354 1562
rect 2318 1538 2322 1542
rect 2286 1438 2290 1442
rect 2262 1428 2266 1432
rect 2358 1508 2362 1512
rect 2334 1478 2338 1482
rect 2310 1468 2314 1472
rect 2294 1378 2298 1382
rect 2310 1438 2314 1442
rect 2318 1348 2322 1352
rect 2270 1338 2274 1342
rect 2334 1338 2338 1342
rect 2014 1328 2018 1332
rect 2030 1328 2034 1332
rect 2046 1328 2050 1332
rect 2190 1328 2194 1332
rect 2222 1328 2226 1332
rect 1998 1308 2002 1312
rect 2030 1308 2034 1312
rect 2022 1278 2026 1282
rect 1998 1268 2002 1272
rect 2006 1268 2010 1272
rect 1990 1238 1994 1242
rect 1878 1208 1882 1212
rect 1990 1208 1994 1212
rect 1918 1158 1922 1162
rect 1830 1138 1834 1142
rect 1878 1128 1882 1132
rect 1950 1128 1954 1132
rect 1870 1118 1874 1122
rect 1990 1108 1994 1112
rect 1830 1078 1834 1082
rect 1870 1078 1874 1082
rect 1886 1078 1890 1082
rect 2022 1148 2026 1152
rect 2014 1138 2018 1142
rect 1998 1068 2002 1072
rect 1822 1058 1826 1062
rect 1838 1058 1842 1062
rect 1830 1048 1834 1052
rect 1806 1038 1810 1042
rect 1782 1018 1786 1022
rect 1758 968 1762 972
rect 1726 958 1730 962
rect 1750 958 1754 962
rect 1806 958 1810 962
rect 1654 948 1658 952
rect 1726 948 1730 952
rect 1622 938 1626 942
rect 1646 938 1650 942
rect 1638 918 1642 922
rect 1598 898 1602 902
rect 1590 888 1594 892
rect 1574 868 1578 872
rect 1518 748 1522 752
rect 1478 678 1482 682
rect 1510 678 1514 682
rect 1494 668 1498 672
rect 1462 658 1466 662
rect 1486 658 1490 662
rect 1438 568 1442 572
rect 1350 448 1354 452
rect 1422 528 1426 532
rect 1430 508 1434 512
rect 1446 508 1450 512
rect 1398 488 1402 492
rect 1390 478 1394 482
rect 1518 668 1522 672
rect 1526 648 1530 652
rect 1526 548 1530 552
rect 1470 518 1474 522
rect 1462 488 1466 492
rect 1438 468 1442 472
rect 1382 448 1386 452
rect 1430 448 1434 452
rect 1438 448 1442 452
rect 1430 438 1434 442
rect 1430 428 1434 432
rect 1358 418 1362 422
rect 1374 418 1378 422
rect 1398 418 1402 422
rect 1454 418 1458 422
rect 1446 398 1450 402
rect 1454 388 1458 392
rect 1438 378 1442 382
rect 1518 528 1522 532
rect 1510 518 1514 522
rect 1518 488 1522 492
rect 1534 458 1538 462
rect 1534 398 1538 402
rect 1510 388 1514 392
rect 1518 388 1522 392
rect 1254 348 1258 352
rect 1406 348 1410 352
rect 1422 348 1426 352
rect 1446 348 1450 352
rect 1238 338 1242 342
rect 1134 258 1138 262
rect 1166 258 1170 262
rect 1046 238 1050 242
rect 1094 238 1098 242
rect 1062 208 1066 212
rect 1086 208 1090 212
rect 1086 198 1090 202
rect 1142 198 1146 202
rect 1062 188 1066 192
rect 1110 148 1114 152
rect 1086 138 1090 142
rect 1118 138 1122 142
rect 1078 118 1082 122
rect 1134 118 1138 122
rect 1058 103 1062 107
rect 1065 103 1069 107
rect 1046 88 1050 92
rect 1190 248 1194 252
rect 1198 208 1202 212
rect 1182 178 1186 182
rect 1238 238 1242 242
rect 1302 308 1306 312
rect 1270 258 1274 262
rect 1302 188 1306 192
rect 1334 338 1338 342
rect 1326 178 1330 182
rect 1230 158 1234 162
rect 1254 158 1258 162
rect 1286 148 1290 152
rect 1638 898 1642 902
rect 1614 868 1618 872
rect 1678 908 1682 912
rect 1734 888 1738 892
rect 1694 868 1698 872
rect 1750 868 1754 872
rect 1590 828 1594 832
rect 1562 803 1566 807
rect 1569 803 1573 807
rect 1630 808 1634 812
rect 1638 788 1642 792
rect 1598 778 1602 782
rect 1630 768 1634 772
rect 1638 768 1642 772
rect 1582 758 1586 762
rect 1614 718 1618 722
rect 1598 708 1602 712
rect 1558 688 1562 692
rect 1582 678 1586 682
rect 1606 688 1610 692
rect 1622 678 1626 682
rect 1638 738 1642 742
rect 1582 658 1586 662
rect 1558 638 1562 642
rect 1550 628 1554 632
rect 1562 603 1566 607
rect 1569 603 1573 607
rect 1654 818 1658 822
rect 1710 798 1714 802
rect 1654 758 1658 762
rect 1702 758 1706 762
rect 1718 778 1722 782
rect 1686 738 1690 742
rect 1670 728 1674 732
rect 1734 708 1738 712
rect 1742 698 1746 702
rect 1646 688 1650 692
rect 1662 688 1666 692
rect 1694 688 1698 692
rect 1718 688 1722 692
rect 1726 688 1730 692
rect 1646 678 1650 682
rect 1678 678 1682 682
rect 1702 668 1706 672
rect 1678 658 1682 662
rect 1694 658 1698 662
rect 1670 638 1674 642
rect 1614 618 1618 622
rect 1590 608 1594 612
rect 1582 598 1586 602
rect 1718 628 1722 632
rect 1590 588 1594 592
rect 1766 948 1770 952
rect 1766 918 1770 922
rect 1822 908 1826 912
rect 1774 888 1778 892
rect 1782 888 1786 892
rect 1822 878 1826 882
rect 1830 858 1834 862
rect 1814 848 1818 852
rect 1822 848 1826 852
rect 1830 838 1834 842
rect 1886 1058 1890 1062
rect 1966 1058 1970 1062
rect 1870 1038 1874 1042
rect 1894 1038 1898 1042
rect 1862 1028 1866 1032
rect 1942 1018 1946 1022
rect 1854 968 1858 972
rect 1974 978 1978 982
rect 1934 958 1938 962
rect 1862 948 1866 952
rect 1878 948 1882 952
rect 1918 948 1922 952
rect 1846 938 1850 942
rect 1894 938 1898 942
rect 1846 918 1850 922
rect 1910 938 1914 942
rect 1902 918 1906 922
rect 1918 898 1922 902
rect 1886 868 1890 872
rect 1902 868 1906 872
rect 1878 858 1882 862
rect 1966 948 1970 952
rect 1982 948 1986 952
rect 1942 908 1946 912
rect 1958 898 1962 902
rect 1942 888 1946 892
rect 1926 858 1930 862
rect 1926 838 1930 842
rect 1854 828 1858 832
rect 1854 808 1858 812
rect 1838 798 1842 802
rect 1822 788 1826 792
rect 1774 738 1778 742
rect 1806 688 1810 692
rect 1774 668 1778 672
rect 1926 758 1930 762
rect 1870 748 1874 752
rect 1902 748 1906 752
rect 1862 738 1866 742
rect 1886 738 1890 742
rect 1846 728 1850 732
rect 1830 718 1834 722
rect 1870 718 1874 722
rect 1910 718 1914 722
rect 1886 708 1890 712
rect 1838 668 1842 672
rect 1894 698 1898 702
rect 1822 658 1826 662
rect 1838 658 1842 662
rect 1798 618 1802 622
rect 1758 578 1762 582
rect 1606 568 1610 572
rect 1630 568 1634 572
rect 1694 568 1698 572
rect 1742 568 1746 572
rect 1574 558 1578 562
rect 1646 558 1650 562
rect 1622 548 1626 552
rect 1766 558 1770 562
rect 1790 558 1794 562
rect 1710 548 1714 552
rect 1750 548 1754 552
rect 1774 548 1778 552
rect 1582 488 1586 492
rect 1550 478 1554 482
rect 1542 388 1546 392
rect 1558 468 1562 472
rect 1558 438 1562 442
rect 1694 538 1698 542
rect 1702 538 1706 542
rect 1686 508 1690 512
rect 1798 538 1802 542
rect 1734 528 1738 532
rect 1774 528 1778 532
rect 1750 518 1754 522
rect 1710 508 1714 512
rect 1670 478 1674 482
rect 1646 448 1650 452
rect 1566 428 1570 432
rect 1598 428 1602 432
rect 1654 428 1658 432
rect 1562 403 1566 407
rect 1569 403 1573 407
rect 1566 388 1570 392
rect 1542 378 1546 382
rect 1558 378 1562 382
rect 1542 338 1546 342
rect 1342 328 1346 332
rect 1534 328 1538 332
rect 1414 298 1418 302
rect 1446 298 1450 302
rect 1422 268 1426 272
rect 1550 288 1554 292
rect 1614 328 1618 332
rect 1590 318 1594 322
rect 1566 278 1570 282
rect 1494 268 1498 272
rect 1342 258 1346 262
rect 1374 258 1378 262
rect 1390 238 1394 242
rect 1470 178 1474 182
rect 1342 148 1346 152
rect 1230 118 1234 122
rect 1222 98 1226 102
rect 1294 98 1298 102
rect 1174 88 1178 92
rect 1198 78 1202 82
rect 1278 78 1282 82
rect 1318 78 1322 82
rect 1518 258 1522 262
rect 1510 248 1514 252
rect 1582 248 1586 252
rect 1638 288 1642 292
rect 1678 388 1682 392
rect 1702 398 1706 402
rect 1686 378 1690 382
rect 1702 378 1706 382
rect 1670 348 1674 352
rect 1654 258 1658 262
rect 1662 248 1666 252
rect 1590 238 1594 242
rect 1562 203 1566 207
rect 1569 203 1573 207
rect 1654 198 1658 202
rect 1590 178 1594 182
rect 1702 308 1706 312
rect 1686 258 1690 262
rect 1686 248 1690 252
rect 1798 518 1802 522
rect 1742 468 1746 472
rect 1766 458 1770 462
rect 1726 448 1730 452
rect 1758 448 1762 452
rect 1718 428 1722 432
rect 1726 388 1730 392
rect 1910 628 1914 632
rect 1902 588 1906 592
rect 1846 548 1850 552
rect 1854 478 1858 482
rect 1830 468 1834 472
rect 1822 448 1826 452
rect 1854 448 1858 452
rect 1878 448 1882 452
rect 1950 868 1954 872
rect 1950 788 1954 792
rect 1974 888 1978 892
rect 1990 888 1994 892
rect 2046 1288 2050 1292
rect 2082 1303 2086 1307
rect 2089 1303 2093 1307
rect 2094 1288 2098 1292
rect 2046 1258 2050 1262
rect 2110 1258 2114 1262
rect 2118 1258 2122 1262
rect 2134 1258 2138 1262
rect 2062 1248 2066 1252
rect 2062 1238 2066 1242
rect 2094 1198 2098 1202
rect 2118 1198 2122 1202
rect 2230 1288 2234 1292
rect 2238 1288 2242 1292
rect 2262 1288 2266 1292
rect 2430 1648 2434 1652
rect 2454 1648 2458 1652
rect 2414 1618 2418 1622
rect 2398 1608 2402 1612
rect 2382 1528 2386 1532
rect 2422 1548 2426 1552
rect 2422 1528 2426 1532
rect 2414 1498 2418 1502
rect 2414 1468 2418 1472
rect 2502 1628 2506 1632
rect 2574 1668 2578 1672
rect 2638 1738 2642 1742
rect 2614 1688 2618 1692
rect 2614 1678 2618 1682
rect 2566 1638 2570 1642
rect 2510 1608 2514 1612
rect 2502 1568 2506 1572
rect 2550 1568 2554 1572
rect 2462 1548 2466 1552
rect 2494 1548 2498 1552
rect 2518 1548 2522 1552
rect 2550 1548 2554 1552
rect 2486 1538 2490 1542
rect 2526 1538 2530 1542
rect 2550 1528 2554 1532
rect 2470 1508 2474 1512
rect 2446 1488 2450 1492
rect 2470 1488 2474 1492
rect 2494 1488 2498 1492
rect 2438 1478 2442 1482
rect 2478 1478 2482 1482
rect 2446 1468 2450 1472
rect 2558 1468 2562 1472
rect 2470 1458 2474 1462
rect 2430 1448 2434 1452
rect 2446 1448 2450 1452
rect 2422 1418 2426 1422
rect 2414 1368 2418 1372
rect 2430 1358 2434 1362
rect 2422 1338 2426 1342
rect 2406 1328 2410 1332
rect 2326 1278 2330 1282
rect 2374 1278 2378 1282
rect 2398 1278 2402 1282
rect 2302 1268 2306 1272
rect 2182 1248 2186 1252
rect 2150 1188 2154 1192
rect 2086 1178 2090 1182
rect 2054 1168 2058 1172
rect 2078 1158 2082 1162
rect 2150 1158 2154 1162
rect 2038 1138 2042 1142
rect 2054 1138 2058 1142
rect 2102 1118 2106 1122
rect 2054 1108 2058 1112
rect 2082 1103 2086 1107
rect 2089 1103 2093 1107
rect 2046 1078 2050 1082
rect 2062 1078 2066 1082
rect 2094 1058 2098 1062
rect 2062 1048 2066 1052
rect 2070 1028 2074 1032
rect 2014 978 2018 982
rect 2014 948 2018 952
rect 2006 928 2010 932
rect 2006 868 2010 872
rect 1974 858 1978 862
rect 1990 858 1994 862
rect 1982 818 1986 822
rect 1958 778 1962 782
rect 1966 768 1970 772
rect 1974 748 1978 752
rect 1982 738 1986 742
rect 2006 738 2010 742
rect 1998 728 2002 732
rect 1974 698 1978 702
rect 2046 898 2050 902
rect 2214 1228 2218 1232
rect 2254 1208 2258 1212
rect 2142 1148 2146 1152
rect 2174 1148 2178 1152
rect 2230 1148 2234 1152
rect 2134 1138 2138 1142
rect 2182 1138 2186 1142
rect 2126 1098 2130 1102
rect 2126 1058 2130 1062
rect 2230 1078 2234 1082
rect 2262 1078 2266 1082
rect 2278 1078 2282 1082
rect 2190 1068 2194 1072
rect 2230 1058 2234 1062
rect 2262 1058 2266 1062
rect 2254 1048 2258 1052
rect 2126 1038 2130 1042
rect 2078 1018 2082 1022
rect 2110 1018 2114 1022
rect 2134 1018 2138 1022
rect 2118 1008 2122 1012
rect 2086 918 2090 922
rect 2118 918 2122 922
rect 2082 903 2086 907
rect 2089 903 2093 907
rect 2046 868 2050 872
rect 2062 858 2066 862
rect 2030 688 2034 692
rect 2126 868 2130 872
rect 2118 838 2122 842
rect 2102 768 2106 772
rect 2078 758 2082 762
rect 2094 748 2098 752
rect 2318 1188 2322 1192
rect 2366 1258 2370 1262
rect 2334 1238 2338 1242
rect 2310 1158 2314 1162
rect 2326 1158 2330 1162
rect 2302 1148 2306 1152
rect 2374 1248 2378 1252
rect 2438 1248 2442 1252
rect 2350 1218 2354 1222
rect 2478 1258 2482 1262
rect 2454 1248 2458 1252
rect 2470 1248 2474 1252
rect 2446 1238 2450 1242
rect 2470 1228 2474 1232
rect 2382 1218 2386 1222
rect 2350 1148 2354 1152
rect 2326 1138 2330 1142
rect 2358 1138 2362 1142
rect 2366 1138 2370 1142
rect 2350 1118 2354 1122
rect 2310 1108 2314 1112
rect 2326 1088 2330 1092
rect 2302 1078 2306 1082
rect 2302 1058 2306 1062
rect 2302 1048 2306 1052
rect 2294 1038 2298 1042
rect 2302 1028 2306 1032
rect 2278 1008 2282 1012
rect 2310 1018 2314 1022
rect 2270 978 2274 982
rect 2198 968 2202 972
rect 2278 968 2282 972
rect 2390 1188 2394 1192
rect 2430 1208 2434 1212
rect 2422 1178 2426 1182
rect 2462 1198 2466 1202
rect 2438 1168 2442 1172
rect 2454 1168 2458 1172
rect 2406 1148 2410 1152
rect 2422 1148 2426 1152
rect 2414 1128 2418 1132
rect 2454 1118 2458 1122
rect 2406 1078 2410 1082
rect 2422 1078 2426 1082
rect 2382 1059 2386 1063
rect 2446 1058 2450 1062
rect 2430 1048 2434 1052
rect 2438 1048 2442 1052
rect 2374 1018 2378 1022
rect 2398 1008 2402 1012
rect 2318 998 2322 1002
rect 2382 998 2386 1002
rect 2270 948 2274 952
rect 2310 948 2314 952
rect 2182 938 2186 942
rect 2206 928 2210 932
rect 2158 908 2162 912
rect 2142 878 2146 882
rect 2134 858 2138 862
rect 2158 858 2162 862
rect 2150 838 2154 842
rect 2134 828 2138 832
rect 2198 898 2202 902
rect 2190 858 2194 862
rect 2174 808 2178 812
rect 2230 898 2234 902
rect 2238 878 2242 882
rect 2366 938 2370 942
rect 2334 928 2338 932
rect 2342 918 2346 922
rect 2318 888 2322 892
rect 2278 878 2282 882
rect 2390 948 2394 952
rect 2414 908 2418 912
rect 2374 898 2378 902
rect 2398 898 2402 902
rect 2230 848 2234 852
rect 2286 848 2290 852
rect 2222 818 2226 822
rect 2238 808 2242 812
rect 2254 808 2258 812
rect 2222 758 2226 762
rect 2230 758 2234 762
rect 2262 798 2266 802
rect 2246 778 2250 782
rect 2166 748 2170 752
rect 2206 748 2210 752
rect 2238 748 2242 752
rect 2070 738 2074 742
rect 2110 728 2114 732
rect 2126 728 2130 732
rect 2082 703 2086 707
rect 2089 703 2093 707
rect 2070 698 2074 702
rect 1974 678 1978 682
rect 2054 678 2058 682
rect 2270 768 2274 772
rect 2262 758 2266 762
rect 2414 848 2418 852
rect 2302 828 2306 832
rect 2342 828 2346 832
rect 2310 818 2314 822
rect 2302 768 2306 772
rect 2262 748 2266 752
rect 2230 718 2234 722
rect 2198 688 2202 692
rect 1998 668 2002 672
rect 2174 678 2178 682
rect 2118 668 2122 672
rect 2126 668 2130 672
rect 1958 658 1962 662
rect 1942 538 1946 542
rect 1910 368 1914 372
rect 1742 358 1746 362
rect 1766 358 1770 362
rect 1838 358 1842 362
rect 1822 348 1826 352
rect 1758 338 1762 342
rect 1774 338 1778 342
rect 1790 318 1794 322
rect 1822 288 1826 292
rect 1758 238 1762 242
rect 1750 228 1754 232
rect 1718 218 1722 222
rect 1654 158 1658 162
rect 1750 158 1754 162
rect 1766 158 1770 162
rect 1486 148 1490 152
rect 1526 148 1530 152
rect 1606 148 1610 152
rect 1710 148 1714 152
rect 1742 148 1746 152
rect 1406 138 1410 142
rect 1446 138 1450 142
rect 1350 98 1354 102
rect 1430 78 1434 82
rect 1486 128 1490 132
rect 1510 128 1514 132
rect 1566 138 1570 142
rect 1646 138 1650 142
rect 1662 138 1666 142
rect 1614 128 1618 132
rect 1662 88 1666 92
rect 1686 88 1690 92
rect 1510 78 1514 82
rect 1574 78 1578 82
rect 1614 78 1618 82
rect 1686 78 1690 82
rect 1094 68 1098 72
rect 1134 68 1138 72
rect 926 58 930 62
rect 942 58 946 62
rect 1022 58 1026 62
rect 1046 58 1050 62
rect 1118 58 1122 62
rect 1174 58 1178 62
rect 1246 58 1250 62
rect 1310 58 1314 62
rect 1342 58 1346 62
rect 1550 58 1554 62
rect 1302 48 1306 52
rect 1326 48 1330 52
rect 1390 48 1394 52
rect 622 38 626 42
rect 1150 38 1154 42
rect 1174 38 1178 42
rect 510 8 514 12
rect 526 8 530 12
rect 546 3 550 7
rect 553 3 557 7
rect 1562 3 1566 7
rect 1569 3 1573 7
rect 1766 138 1770 142
rect 1758 88 1762 92
rect 1846 308 1850 312
rect 1846 288 1850 292
rect 1814 218 1818 222
rect 1830 218 1834 222
rect 1830 168 1834 172
rect 1838 158 1842 162
rect 1798 118 1802 122
rect 1878 358 1882 362
rect 1894 348 1898 352
rect 1886 338 1890 342
rect 1870 328 1874 332
rect 1862 188 1866 192
rect 1870 158 1874 162
rect 1902 338 1906 342
rect 1966 608 1970 612
rect 2022 658 2026 662
rect 2086 648 2090 652
rect 2142 658 2146 662
rect 2126 638 2130 642
rect 2054 628 2058 632
rect 2110 628 2114 632
rect 2118 628 2122 632
rect 1990 568 1994 572
rect 2014 568 2018 572
rect 2022 558 2026 562
rect 2006 548 2010 552
rect 1950 528 1954 532
rect 1958 518 1962 522
rect 1974 518 1978 522
rect 1998 518 2002 522
rect 1998 478 2002 482
rect 1990 468 1994 472
rect 1966 438 1970 442
rect 2022 518 2026 522
rect 2014 468 2018 472
rect 2014 448 2018 452
rect 1966 348 1970 352
rect 1950 338 1954 342
rect 1934 328 1938 332
rect 1910 308 1914 312
rect 1910 288 1914 292
rect 1950 288 1954 292
rect 1958 288 1962 292
rect 1886 148 1890 152
rect 1966 238 1970 242
rect 2062 578 2066 582
rect 2094 558 2098 562
rect 2102 548 2106 552
rect 2142 547 2146 551
rect 2118 528 2122 532
rect 2082 503 2086 507
rect 2089 503 2093 507
rect 2190 648 2194 652
rect 2182 558 2186 562
rect 2238 708 2242 712
rect 2294 708 2298 712
rect 2278 688 2282 692
rect 2326 778 2330 782
rect 2326 768 2330 772
rect 2318 758 2322 762
rect 2326 748 2330 752
rect 2318 708 2322 712
rect 2246 678 2250 682
rect 2254 668 2258 672
rect 2294 668 2298 672
rect 2270 628 2274 632
rect 2254 588 2258 592
rect 2270 568 2274 572
rect 2230 548 2234 552
rect 2198 518 2202 522
rect 2062 488 2066 492
rect 2174 488 2178 492
rect 2118 478 2122 482
rect 2134 468 2138 472
rect 2246 538 2250 542
rect 2238 488 2242 492
rect 2262 538 2266 542
rect 2070 458 2074 462
rect 2118 458 2122 462
rect 2046 438 2050 442
rect 2046 418 2050 422
rect 2038 408 2042 412
rect 2030 358 2034 362
rect 2166 448 2170 452
rect 2126 408 2130 412
rect 2214 448 2218 452
rect 2182 438 2186 442
rect 2174 398 2178 402
rect 2118 388 2122 392
rect 2046 358 2050 362
rect 2070 358 2074 362
rect 1990 328 1994 332
rect 2022 328 2026 332
rect 2150 378 2154 382
rect 2198 358 2202 362
rect 2070 338 2074 342
rect 2070 328 2074 332
rect 2102 328 2106 332
rect 2014 308 2018 312
rect 2038 308 2042 312
rect 2006 268 2010 272
rect 1958 188 1962 192
rect 1942 128 1946 132
rect 1926 118 1930 122
rect 1894 88 1898 92
rect 1710 78 1714 82
rect 1774 78 1778 82
rect 1790 78 1794 82
rect 1910 78 1914 82
rect 1718 68 1722 72
rect 1742 68 1746 72
rect 1766 68 1770 72
rect 1734 58 1738 62
rect 1966 148 1970 152
rect 2030 288 2034 292
rect 2054 288 2058 292
rect 2054 278 2058 282
rect 2030 268 2034 272
rect 2038 258 2042 262
rect 1998 138 2002 142
rect 2158 328 2162 332
rect 2190 328 2194 332
rect 2142 318 2146 322
rect 2082 303 2086 307
rect 2089 303 2093 307
rect 2190 298 2194 302
rect 2222 338 2226 342
rect 2262 438 2266 442
rect 2254 418 2258 422
rect 2382 788 2386 792
rect 2382 768 2386 772
rect 2542 1388 2546 1392
rect 2502 1338 2506 1342
rect 2590 1558 2594 1562
rect 2598 1538 2602 1542
rect 2622 1618 2626 1622
rect 2646 1648 2650 1652
rect 2638 1478 2642 1482
rect 2646 1448 2650 1452
rect 2606 1428 2610 1432
rect 2606 1408 2610 1412
rect 2646 1388 2650 1392
rect 2566 1368 2570 1372
rect 2590 1368 2594 1372
rect 2574 1348 2578 1352
rect 2606 1348 2610 1352
rect 2550 1338 2554 1342
rect 2558 1338 2562 1342
rect 2598 1338 2602 1342
rect 2534 1328 2538 1332
rect 2574 1328 2578 1332
rect 2582 1328 2586 1332
rect 2638 1318 2642 1322
rect 2502 1278 2506 1282
rect 2582 1278 2586 1282
rect 2494 1268 2498 1272
rect 2598 1268 2602 1272
rect 2486 1208 2490 1212
rect 2550 1258 2554 1262
rect 2494 1188 2498 1192
rect 2518 1158 2522 1162
rect 2566 1168 2570 1172
rect 2590 1147 2594 1151
rect 2542 1128 2546 1132
rect 2470 1088 2474 1092
rect 2534 1088 2538 1092
rect 2574 1078 2578 1082
rect 2510 1068 2514 1072
rect 2550 968 2554 972
rect 2502 958 2506 962
rect 2454 928 2458 932
rect 2462 928 2466 932
rect 2470 848 2474 852
rect 2430 798 2434 802
rect 2438 748 2442 752
rect 2454 748 2458 752
rect 2510 948 2514 952
rect 2526 948 2530 952
rect 2550 928 2554 932
rect 2534 918 2538 922
rect 2494 758 2498 762
rect 2502 758 2506 762
rect 2494 748 2498 752
rect 2478 738 2482 742
rect 2438 728 2442 732
rect 2462 728 2466 732
rect 2470 718 2474 722
rect 2494 718 2498 722
rect 2430 688 2434 692
rect 2382 678 2386 682
rect 2454 678 2458 682
rect 2478 668 2482 672
rect 2486 668 2490 672
rect 2326 618 2330 622
rect 2302 558 2306 562
rect 2286 538 2290 542
rect 2318 538 2322 542
rect 2358 598 2362 602
rect 2342 558 2346 562
rect 2366 558 2370 562
rect 2406 558 2410 562
rect 2334 528 2338 532
rect 2310 518 2314 522
rect 2350 518 2354 522
rect 2350 488 2354 492
rect 2310 468 2314 472
rect 2326 468 2330 472
rect 2334 458 2338 462
rect 2390 528 2394 532
rect 2422 648 2426 652
rect 2438 648 2442 652
rect 2462 628 2466 632
rect 2518 908 2522 912
rect 2510 678 2514 682
rect 2502 658 2506 662
rect 2494 618 2498 622
rect 2510 618 2514 622
rect 2430 588 2434 592
rect 2422 568 2426 572
rect 2478 548 2482 552
rect 2486 538 2490 542
rect 2462 518 2466 522
rect 2414 508 2418 512
rect 2462 488 2466 492
rect 2478 488 2482 492
rect 2382 478 2386 482
rect 2446 478 2450 482
rect 2438 468 2442 472
rect 2374 448 2378 452
rect 2302 438 2306 442
rect 2414 438 2418 442
rect 2286 428 2290 432
rect 2262 358 2266 362
rect 2254 338 2258 342
rect 2222 298 2226 302
rect 2262 298 2266 302
rect 2102 288 2106 292
rect 2206 288 2210 292
rect 2230 288 2234 292
rect 2238 288 2242 292
rect 2134 278 2138 282
rect 2182 268 2186 272
rect 2270 288 2274 292
rect 2326 368 2330 372
rect 2358 368 2362 372
rect 2414 368 2418 372
rect 2350 358 2354 362
rect 2310 348 2314 352
rect 2366 348 2370 352
rect 2510 548 2514 552
rect 2566 978 2570 982
rect 2622 1288 2626 1292
rect 2646 1278 2650 1282
rect 2630 1248 2634 1252
rect 2638 1188 2642 1192
rect 2614 1168 2618 1172
rect 2638 1138 2642 1142
rect 2614 1078 2618 1082
rect 2622 1058 2626 1062
rect 2598 1048 2602 1052
rect 2574 948 2578 952
rect 2590 948 2594 952
rect 2598 938 2602 942
rect 2582 928 2586 932
rect 2558 878 2562 882
rect 2558 868 2562 872
rect 2574 868 2578 872
rect 2622 898 2626 902
rect 2646 1048 2650 1052
rect 2646 968 2650 972
rect 2606 858 2610 862
rect 2534 848 2538 852
rect 2582 848 2586 852
rect 2542 758 2546 762
rect 2526 678 2530 682
rect 2566 718 2570 722
rect 2574 718 2578 722
rect 2550 688 2554 692
rect 2558 668 2562 672
rect 2542 658 2546 662
rect 2542 638 2546 642
rect 2558 628 2562 632
rect 2550 578 2554 582
rect 2534 568 2538 572
rect 2606 648 2610 652
rect 2606 578 2610 582
rect 2590 568 2594 572
rect 2590 558 2594 562
rect 2550 548 2554 552
rect 2574 548 2578 552
rect 2566 538 2570 542
rect 2598 538 2602 542
rect 2526 508 2530 512
rect 2590 508 2594 512
rect 2526 478 2530 482
rect 2526 468 2530 472
rect 2510 458 2514 462
rect 2534 458 2538 462
rect 2598 458 2602 462
rect 2502 428 2506 432
rect 2478 418 2482 422
rect 2470 398 2474 402
rect 2494 398 2498 402
rect 2494 348 2498 352
rect 2326 318 2330 322
rect 2358 308 2362 312
rect 2342 288 2346 292
rect 2462 308 2466 312
rect 2478 308 2482 312
rect 2430 288 2434 292
rect 2398 278 2402 282
rect 2166 258 2170 262
rect 2086 168 2090 172
rect 2118 168 2122 172
rect 2118 158 2122 162
rect 2182 158 2186 162
rect 2102 148 2106 152
rect 2134 148 2138 152
rect 2110 138 2114 142
rect 2062 118 2066 122
rect 2006 88 2010 92
rect 2046 88 2050 92
rect 2082 103 2086 107
rect 2089 103 2093 107
rect 2110 78 2114 82
rect 2190 118 2194 122
rect 2182 78 2186 82
rect 2222 218 2226 222
rect 2278 208 2282 212
rect 2270 168 2274 172
rect 2246 138 2250 142
rect 2206 98 2210 102
rect 2254 98 2258 102
rect 2254 88 2258 92
rect 2062 68 2066 72
rect 2150 68 2154 72
rect 1758 58 1762 62
rect 1806 58 1810 62
rect 1878 58 1882 62
rect 2062 58 2066 62
rect 2286 158 2290 162
rect 2270 68 2274 72
rect 2486 298 2490 302
rect 2390 268 2394 272
rect 2398 268 2402 272
rect 2310 148 2314 152
rect 2374 148 2378 152
rect 2446 258 2450 262
rect 2438 248 2442 252
rect 2470 248 2474 252
rect 2606 448 2610 452
rect 2606 438 2610 442
rect 2566 348 2570 352
rect 2598 348 2602 352
rect 2534 278 2538 282
rect 2502 258 2506 262
rect 2510 258 2514 262
rect 2502 178 2506 182
rect 2518 168 2522 172
rect 2510 148 2514 152
rect 2478 138 2482 142
rect 2486 138 2490 142
rect 2294 98 2298 102
rect 2302 98 2306 102
rect 2374 98 2378 102
rect 2478 98 2482 102
rect 2422 88 2426 92
rect 2438 88 2442 92
rect 2462 88 2466 92
rect 2390 78 2394 82
rect 2342 58 2346 62
rect 2614 308 2618 312
rect 2630 568 2634 572
rect 2646 438 2650 442
rect 2630 348 2634 352
rect 2566 238 2570 242
rect 2550 198 2554 202
rect 2542 178 2546 182
rect 2598 148 2602 152
rect 2566 68 2570 72
rect 2598 68 2602 72
rect 2518 58 2522 62
rect 2638 278 2642 282
rect 2630 58 2634 62
rect 2142 48 2146 52
rect 2174 48 2178 52
rect 2502 48 2506 52
<< metal3 >>
rect 544 2403 546 2407
rect 550 2403 553 2407
rect 558 2403 560 2407
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1574 2403 1576 2407
rect 490 2398 502 2401
rect 1178 2398 1198 2401
rect 1530 2398 1534 2401
rect 2290 2398 2302 2401
rect 218 2368 286 2371
rect 290 2368 294 2371
rect 298 2368 366 2371
rect 370 2368 534 2371
rect 1186 2368 1246 2371
rect 1266 2368 1606 2371
rect 1626 2368 1758 2371
rect 1762 2368 1766 2371
rect 1810 2368 1942 2371
rect 2418 2368 2430 2371
rect 330 2358 926 2361
rect 1042 2358 1086 2361
rect 1146 2358 1390 2361
rect 1394 2358 1422 2361
rect 1474 2358 1534 2361
rect 1642 2358 1686 2361
rect 1846 2358 1854 2361
rect 1858 2358 1886 2361
rect 626 2348 654 2351
rect 818 2348 886 2351
rect 986 2348 1022 2351
rect 1082 2348 1238 2351
rect 1242 2348 1262 2351
rect 1330 2348 1398 2351
rect 1426 2348 1822 2351
rect 1826 2348 1838 2351
rect 2042 2348 2070 2351
rect 2442 2348 2478 2351
rect -26 2341 -22 2342
rect -26 2338 6 2341
rect 10 2338 14 2341
rect 18 2338 70 2341
rect 74 2338 230 2341
rect 358 2341 361 2348
rect 446 2341 449 2348
rect 242 2338 449 2341
rect 658 2338 710 2341
rect 1114 2338 1142 2341
rect 1162 2338 1297 2341
rect 1610 2338 1646 2341
rect 1762 2338 1822 2341
rect 2214 2341 2217 2348
rect 1858 2338 2217 2341
rect 2226 2338 2230 2341
rect 2234 2338 2246 2341
rect 2250 2338 2534 2341
rect 1294 2332 1297 2338
rect 606 2328 686 2331
rect 690 2328 798 2331
rect 1010 2328 1118 2331
rect 1370 2328 1462 2331
rect 1466 2328 1494 2331
rect 1658 2328 1854 2331
rect 2138 2328 2206 2331
rect 2210 2328 2270 2331
rect 2522 2328 2622 2331
rect 606 2322 609 2328
rect 10 2318 54 2321
rect 674 2318 726 2321
rect 730 2318 758 2321
rect 1034 2318 1086 2321
rect 1210 2318 1230 2321
rect 1234 2318 1430 2321
rect 1714 2318 2334 2321
rect 2338 2318 2558 2321
rect 834 2308 950 2311
rect 1226 2308 1278 2311
rect 1056 2303 1058 2307
rect 1062 2303 1065 2307
rect 1070 2303 1072 2307
rect 2080 2303 2082 2307
rect 2086 2303 2089 2307
rect 2094 2303 2096 2307
rect 498 2298 750 2301
rect 874 2298 942 2301
rect 1082 2298 1102 2301
rect 1106 2298 1166 2301
rect 1298 2298 1446 2301
rect 1450 2298 1486 2301
rect 1490 2298 1742 2301
rect 1746 2298 1766 2301
rect 1770 2298 1966 2301
rect 2218 2298 2238 2301
rect 66 2288 158 2291
rect 162 2288 254 2291
rect 642 2288 686 2291
rect 890 2288 1022 2291
rect 1078 2291 1081 2298
rect 1026 2288 1081 2291
rect 1098 2288 1222 2291
rect 1362 2288 1414 2291
rect 1490 2288 1526 2291
rect 1554 2288 1774 2291
rect 1994 2288 1998 2291
rect 2018 2288 2046 2291
rect 2050 2288 2102 2291
rect 426 2278 598 2281
rect 754 2278 1662 2281
rect 1794 2278 1958 2281
rect 1970 2278 1990 2281
rect 2150 2281 2153 2288
rect 2074 2278 2153 2281
rect 2322 2278 2406 2281
rect 2410 2278 2430 2281
rect 2498 2278 2534 2281
rect 70 2268 89 2271
rect 190 2271 193 2278
rect 130 2268 193 2271
rect 322 2268 382 2271
rect 386 2268 398 2271
rect 426 2268 478 2271
rect 482 2268 526 2271
rect 578 2268 662 2271
rect 810 2268 862 2271
rect 906 2268 1102 2271
rect 1106 2268 1158 2271
rect 1306 2268 1382 2271
rect 1594 2268 1630 2271
rect 1634 2268 1726 2271
rect 1738 2268 1774 2271
rect 1818 2268 1846 2271
rect 1934 2268 2038 2271
rect 2086 2268 2142 2271
rect 2370 2268 2462 2271
rect 2546 2268 2566 2271
rect 2570 2268 2614 2271
rect 70 2262 73 2268
rect 86 2262 89 2268
rect 1254 2262 1257 2268
rect 1414 2262 1417 2268
rect 1934 2262 1937 2268
rect 2086 2262 2089 2268
rect 186 2258 206 2261
rect 322 2258 326 2261
rect 346 2258 430 2261
rect 458 2258 502 2261
rect 522 2258 846 2261
rect 850 2258 878 2261
rect 1074 2258 1118 2261
rect 1314 2258 1318 2261
rect 1338 2258 1358 2261
rect 1386 2258 1398 2261
rect 1426 2258 1470 2261
rect 1538 2258 1558 2261
rect 1690 2258 1758 2261
rect 1786 2258 1854 2261
rect 2146 2258 2158 2261
rect 2342 2261 2345 2268
rect 2342 2258 2414 2261
rect 2454 2258 2470 2261
rect 2454 2252 2457 2258
rect 154 2248 174 2251
rect 178 2248 214 2251
rect 218 2248 334 2251
rect 650 2248 670 2251
rect 738 2248 897 2251
rect 1082 2248 1174 2251
rect 1266 2248 1350 2251
rect 1354 2248 1518 2251
rect 1850 2248 1902 2251
rect 2346 2248 2350 2251
rect 2370 2248 2382 2251
rect 2442 2248 2454 2251
rect 2466 2248 2534 2251
rect 178 2238 222 2241
rect 266 2238 350 2241
rect 626 2238 638 2241
rect 642 2238 886 2241
rect 894 2241 897 2248
rect 894 2238 1270 2241
rect 1362 2238 1382 2241
rect 1386 2238 1790 2241
rect 1794 2238 1814 2241
rect 1818 2238 1830 2241
rect 602 2228 974 2231
rect 1410 2228 1430 2231
rect 1826 2228 2374 2231
rect 522 2218 734 2221
rect 738 2218 838 2221
rect 1202 2218 1214 2221
rect 1218 2218 1382 2221
rect 1954 2218 1998 2221
rect 2002 2218 2118 2221
rect 2122 2218 2166 2221
rect 2170 2218 2238 2221
rect 2554 2218 2558 2221
rect 746 2208 1078 2211
rect 1114 2208 1238 2211
rect 1274 2208 1278 2211
rect 544 2203 546 2207
rect 550 2203 553 2207
rect 558 2203 560 2207
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1574 2203 1576 2207
rect 1122 2198 1534 2201
rect 306 2188 814 2191
rect 1090 2188 1150 2191
rect 2258 2188 2278 2191
rect 458 2178 1262 2181
rect 1930 2178 2206 2181
rect 266 2168 742 2171
rect 802 2168 838 2171
rect 1130 2168 1206 2171
rect 1618 2168 1686 2171
rect 1690 2168 1774 2171
rect 1794 2168 1982 2171
rect 1986 2168 2182 2171
rect 2530 2168 2550 2171
rect 2262 2162 2265 2168
rect 322 2158 374 2161
rect 434 2158 454 2161
rect 666 2158 670 2161
rect 674 2158 678 2161
rect 778 2158 950 2161
rect 954 2158 1078 2161
rect 1146 2158 1150 2161
rect 1762 2158 1870 2161
rect 2442 2158 2478 2161
rect 70 2151 73 2158
rect 70 2148 126 2151
rect 370 2148 390 2151
rect 418 2148 449 2151
rect 618 2148 638 2151
rect 690 2148 758 2151
rect 794 2148 1166 2151
rect 1170 2148 1198 2151
rect 1298 2148 1310 2151
rect 1526 2151 1529 2158
rect 1490 2148 1598 2151
rect 1742 2151 1745 2158
rect 1742 2148 1790 2151
rect 1818 2148 1838 2151
rect 2126 2151 2129 2158
rect 1962 2148 2129 2151
rect 2178 2148 2310 2151
rect 2594 2148 2622 2151
rect 446 2142 449 2148
rect 638 2142 641 2148
rect 1350 2142 1353 2148
rect 122 2138 150 2141
rect 154 2138 190 2141
rect 450 2138 510 2141
rect 538 2138 614 2141
rect 938 2138 1006 2141
rect 1114 2138 1174 2141
rect 1682 2138 1710 2141
rect 1858 2138 1937 2141
rect 2002 2138 2198 2141
rect 2226 2138 2326 2141
rect 2342 2141 2345 2148
rect 2342 2138 2390 2141
rect 1822 2132 1825 2138
rect 1934 2132 1937 2138
rect 10 2128 62 2131
rect 258 2128 350 2131
rect 378 2128 494 2131
rect 514 2128 646 2131
rect 1114 2128 1142 2131
rect 1146 2128 1214 2131
rect 1298 2128 1302 2131
rect 1306 2128 1422 2131
rect 1786 2128 1822 2131
rect 2058 2128 2358 2131
rect 18 2118 102 2121
rect 106 2118 302 2121
rect 314 2118 382 2121
rect 386 2118 798 2121
rect 1058 2118 1078 2121
rect 1082 2118 1158 2121
rect 1186 2118 1334 2121
rect 1506 2118 1510 2121
rect 1706 2118 1942 2121
rect 1946 2118 1966 2121
rect 1970 2118 2062 2121
rect 2074 2118 2086 2121
rect 2138 2118 2270 2121
rect 2282 2118 2414 2121
rect 210 2108 518 2111
rect 786 2108 862 2111
rect 1146 2108 1270 2111
rect 1978 2108 1990 2111
rect 2202 2108 2526 2111
rect 2594 2108 2614 2111
rect 1056 2103 1058 2107
rect 1062 2103 1065 2107
rect 1070 2103 1072 2107
rect 2080 2103 2082 2107
rect 2086 2103 2089 2107
rect 2094 2103 2096 2107
rect 362 2098 406 2101
rect 562 2098 582 2101
rect 754 2098 806 2101
rect 1002 2098 1014 2101
rect 1078 2098 1222 2101
rect 2114 2098 2278 2101
rect 2290 2098 2406 2101
rect 2410 2098 2462 2101
rect 106 2088 150 2091
rect 154 2088 302 2091
rect 418 2088 454 2091
rect 458 2088 470 2091
rect 1078 2091 1081 2098
rect 1042 2088 1081 2091
rect 1966 2091 1969 2098
rect 1418 2088 1465 2091
rect 1966 2088 2030 2091
rect 2266 2088 2294 2091
rect 138 2078 174 2081
rect 194 2078 345 2081
rect 354 2078 422 2081
rect 426 2078 433 2081
rect 642 2078 710 2081
rect 738 2078 750 2081
rect 986 2078 1014 2081
rect 1026 2078 1166 2081
rect 1190 2081 1193 2088
rect 1462 2082 1465 2088
rect 2118 2082 2121 2088
rect 1190 2078 1278 2081
rect 1370 2078 1414 2081
rect 1466 2078 1478 2081
rect 1546 2078 1582 2081
rect 1586 2078 1825 2081
rect 1834 2078 1910 2081
rect 2218 2078 2286 2081
rect 106 2068 142 2071
rect 342 2071 345 2078
rect 342 2068 766 2071
rect 770 2068 782 2071
rect 802 2068 1070 2071
rect 1074 2068 1622 2071
rect 1630 2068 1638 2071
rect 1642 2068 1710 2071
rect 1822 2071 1825 2078
rect 1822 2068 1990 2071
rect 1994 2068 2230 2071
rect 2234 2068 2278 2071
rect 2298 2068 2302 2071
rect 2382 2071 2385 2078
rect 2382 2068 2558 2071
rect 58 2058 118 2061
rect 170 2058 270 2061
rect 322 2058 406 2061
rect 410 2058 438 2061
rect 458 2058 494 2061
rect 570 2058 654 2061
rect 682 2058 782 2061
rect 786 2058 790 2061
rect 858 2058 902 2061
rect 930 2058 1126 2061
rect 1178 2058 1462 2061
rect 1466 2058 1641 2061
rect 1810 2058 1846 2061
rect 2026 2058 2054 2061
rect 2122 2058 2142 2061
rect 2146 2058 2158 2061
rect 2162 2058 2174 2061
rect 2186 2058 2214 2061
rect 2242 2058 2262 2061
rect 2274 2058 2342 2061
rect 2442 2058 2510 2061
rect 1166 2052 1169 2058
rect 90 2048 326 2051
rect 338 2048 478 2051
rect 482 2048 934 2051
rect 1170 2048 1190 2051
rect 1426 2048 1446 2051
rect 1534 2048 1553 2051
rect 1610 2048 1630 2051
rect 1638 2051 1641 2058
rect 2006 2052 2009 2058
rect 1638 2048 2006 2051
rect 2106 2048 2126 2051
rect 2130 2048 2398 2051
rect 1446 2042 1449 2048
rect 1534 2042 1537 2048
rect 1550 2042 1553 2048
rect 1630 2042 1633 2048
rect 138 2038 390 2041
rect 866 2038 902 2041
rect 1354 2038 1425 2041
rect 1850 2038 1902 2041
rect 1422 2032 1425 2038
rect 178 2028 214 2031
rect 218 2028 694 2031
rect 698 2028 1118 2031
rect 1530 2028 1534 2031
rect 1546 2028 1990 2031
rect 1994 2028 2246 2031
rect 2250 2028 2310 2031
rect 1542 2022 1545 2028
rect 314 2018 526 2021
rect 906 2018 1046 2021
rect 1050 2018 1318 2021
rect 1322 2018 1422 2021
rect 1578 2018 1942 2021
rect 1946 2018 2294 2021
rect 874 2008 894 2011
rect 1794 2008 1854 2011
rect 1890 2008 2190 2011
rect 544 2003 546 2007
rect 550 2003 553 2007
rect 558 2003 560 2007
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1574 2003 1576 2007
rect 674 1998 998 2001
rect 1978 1998 1990 2001
rect 2066 1998 2270 2001
rect 2274 1998 2302 2001
rect 442 1988 878 1991
rect 890 1988 950 1991
rect 1874 1988 1950 1991
rect 2106 1988 2462 1991
rect 330 1978 494 1981
rect 658 1978 702 1981
rect 722 1978 950 1981
rect 1082 1978 1734 1981
rect 1738 1978 2238 1981
rect 2242 1978 2254 1981
rect 394 1968 694 1971
rect 842 1968 1086 1971
rect 1290 1968 1406 1971
rect 1410 1968 1454 1971
rect 2122 1968 2182 1971
rect 2250 1968 2502 1971
rect 2506 1968 2558 1971
rect 194 1958 262 1961
rect 270 1961 273 1968
rect 270 1958 342 1961
rect 850 1958 854 1961
rect 858 1958 918 1961
rect 938 1958 1126 1961
rect 1154 1958 1214 1961
rect 1310 1958 1318 1961
rect 1322 1958 1350 1961
rect 1586 1958 1670 1961
rect 2138 1958 2142 1961
rect 2146 1958 2174 1961
rect 2178 1958 2222 1961
rect 2226 1958 2478 1961
rect 122 1948 198 1951
rect 370 1948 526 1951
rect 574 1951 577 1958
rect 574 1948 646 1951
rect 686 1951 689 1958
rect 686 1948 758 1951
rect 826 1948 886 1951
rect 922 1948 990 1951
rect 1202 1948 1222 1951
rect 1274 1948 1310 1951
rect 1554 1948 1558 1951
rect 1562 1948 1590 1951
rect 1594 1948 1822 1951
rect 1826 1948 1838 1951
rect 1906 1948 1974 1951
rect 2010 1948 2070 1951
rect 2086 1951 2089 1958
rect 2086 1948 2150 1951
rect 2306 1948 2374 1951
rect 2466 1948 2502 1951
rect 10 1938 62 1941
rect 86 1941 89 1948
rect 66 1938 89 1941
rect 278 1941 281 1948
rect 210 1938 281 1941
rect 418 1938 494 1941
rect 514 1938 622 1941
rect 706 1938 886 1941
rect 1006 1941 1009 1948
rect 1310 1942 1313 1948
rect 1006 1938 1302 1941
rect 1318 1941 1321 1948
rect 1318 1938 1366 1941
rect 1370 1938 1534 1941
rect 1538 1938 1598 1941
rect 1666 1938 1798 1941
rect 2042 1938 2158 1941
rect 2162 1938 2190 1941
rect 2274 1938 2430 1941
rect 2458 1938 2574 1941
rect 194 1928 214 1931
rect 234 1928 286 1931
rect 442 1928 630 1931
rect 634 1928 670 1931
rect 802 1928 806 1931
rect 1306 1928 1326 1931
rect 1330 1928 1558 1931
rect 1722 1928 1790 1931
rect 1970 1928 2022 1931
rect 2434 1928 2614 1931
rect 230 1921 233 1928
rect 194 1918 233 1921
rect 250 1918 270 1921
rect 274 1918 342 1921
rect 538 1918 654 1921
rect 666 1918 878 1921
rect 1034 1918 1078 1921
rect 1082 1918 1182 1921
rect 1718 1921 1721 1928
rect 1698 1918 1721 1921
rect 2018 1918 2030 1921
rect 2034 1918 2118 1921
rect 2410 1918 2534 1921
rect 2618 1918 2646 1921
rect 66 1908 390 1911
rect 538 1908 654 1911
rect 658 1908 710 1911
rect 834 1908 846 1911
rect 1594 1908 1646 1911
rect 2258 1908 2382 1911
rect 2386 1908 2430 1911
rect 1056 1903 1058 1907
rect 1062 1903 1065 1907
rect 1070 1903 1072 1907
rect 2080 1903 2082 1907
rect 2086 1903 2089 1907
rect 2094 1903 2096 1907
rect 138 1898 222 1901
rect 226 1898 270 1901
rect 274 1898 366 1901
rect 370 1898 422 1901
rect 426 1898 1046 1901
rect 1266 1898 1670 1901
rect 1858 1898 1870 1901
rect 1874 1898 1926 1901
rect 2330 1898 2510 1901
rect 266 1888 318 1891
rect 322 1888 430 1891
rect 594 1888 614 1891
rect 738 1888 822 1891
rect 826 1888 846 1891
rect 1010 1888 1070 1891
rect 1074 1888 1158 1891
rect 1314 1888 1462 1891
rect 1738 1888 1750 1891
rect 1754 1888 2342 1891
rect 202 1878 286 1881
rect 674 1878 694 1881
rect 938 1878 1102 1881
rect 1106 1878 1206 1881
rect 1310 1881 1313 1888
rect 1306 1878 1313 1881
rect 1378 1878 1430 1881
rect 1642 1878 1654 1881
rect 1658 1878 1710 1881
rect 1794 1878 1798 1881
rect 2066 1878 2334 1881
rect 146 1868 382 1871
rect 410 1868 438 1871
rect 610 1868 841 1871
rect 106 1858 118 1861
rect 158 1858 230 1861
rect 298 1858 337 1861
rect 354 1858 358 1861
rect 418 1858 425 1861
rect 502 1861 505 1868
rect 474 1858 505 1861
rect 558 1861 561 1868
rect 558 1858 566 1861
rect 602 1858 638 1861
rect 690 1858 702 1861
rect 838 1861 841 1868
rect 1130 1868 1182 1871
rect 1206 1871 1209 1878
rect 1206 1868 1230 1871
rect 1602 1868 1654 1871
rect 1674 1868 1854 1871
rect 1858 1868 1998 1871
rect 2010 1868 2038 1871
rect 2298 1868 2318 1871
rect 2370 1868 2382 1871
rect 2386 1868 2438 1871
rect 2518 1871 2521 1878
rect 2518 1868 2598 1871
rect 722 1858 769 1861
rect 158 1852 161 1858
rect 334 1852 337 1858
rect 422 1852 425 1858
rect 686 1852 689 1858
rect 766 1852 769 1858
rect 838 1858 910 1861
rect 982 1861 985 1868
rect 938 1858 945 1861
rect 982 1858 1022 1861
rect 1146 1858 1214 1861
rect 1218 1858 1262 1861
rect 1398 1861 1401 1868
rect 1330 1858 1401 1861
rect 1482 1858 1518 1861
rect 1626 1858 2022 1861
rect 2150 1861 2153 1868
rect 2138 1858 2153 1861
rect 2186 1858 2214 1861
rect 2334 1858 2342 1861
rect 2402 1858 2438 1861
rect 2442 1858 2470 1861
rect 838 1852 841 1858
rect 942 1852 945 1858
rect 2334 1852 2337 1858
rect 2374 1852 2377 1858
rect 42 1848 118 1851
rect 274 1848 326 1851
rect 554 1848 566 1851
rect 650 1848 662 1851
rect 1146 1848 1182 1851
rect 1186 1848 1198 1851
rect 1226 1848 1398 1851
rect 1426 1848 1886 1851
rect 1986 1848 2030 1851
rect 2034 1848 2038 1851
rect 2422 1848 2430 1851
rect 2434 1848 2494 1851
rect 370 1838 414 1841
rect 418 1838 422 1841
rect 490 1838 518 1841
rect 522 1838 614 1841
rect 938 1838 1094 1841
rect 2290 1838 2606 1841
rect 2610 1838 2622 1841
rect 682 1828 974 1831
rect 1394 1828 1414 1831
rect 1514 1828 1518 1831
rect 1722 1828 2414 1831
rect 1414 1822 1417 1828
rect 498 1818 790 1821
rect 1426 1818 1758 1821
rect 1762 1818 2094 1821
rect 2098 1818 2350 1821
rect 722 1808 1046 1811
rect 1050 1808 1422 1811
rect 1658 1808 1766 1811
rect 1818 1808 1894 1811
rect 1962 1808 2134 1811
rect 2346 1808 2374 1811
rect 544 1803 546 1807
rect 550 1803 553 1807
rect 558 1803 560 1807
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1574 1803 1576 1807
rect 858 1798 886 1801
rect 890 1798 902 1801
rect 1850 1798 2462 1801
rect 2466 1798 2494 1801
rect 570 1788 990 1791
rect 1626 1788 1854 1791
rect 1978 1788 2142 1791
rect 2194 1788 2302 1791
rect 1974 1782 1977 1788
rect 218 1778 254 1781
rect 314 1778 430 1781
rect 586 1778 958 1781
rect 1274 1778 1334 1781
rect 1338 1778 1342 1781
rect 2058 1778 2110 1781
rect 2298 1778 2638 1781
rect 146 1768 174 1771
rect 298 1768 310 1771
rect 394 1768 558 1771
rect 674 1768 710 1771
rect 978 1768 1054 1771
rect 1426 1768 1486 1771
rect 1610 1768 1646 1771
rect 1698 1768 1710 1771
rect 1954 1768 2062 1771
rect 2242 1768 2334 1771
rect 262 1761 265 1768
rect 262 1758 302 1761
rect 338 1758 382 1761
rect 386 1758 686 1761
rect 690 1758 702 1761
rect 706 1758 710 1761
rect 1002 1758 1014 1761
rect 1074 1758 1094 1761
rect 1150 1761 1153 1768
rect 1146 1758 1153 1761
rect 1490 1758 1782 1761
rect 1786 1758 1862 1761
rect 1866 1758 1918 1761
rect 1942 1761 1945 1768
rect 1942 1758 1990 1761
rect 2074 1758 2206 1761
rect 2310 1758 2318 1761
rect 2466 1758 2481 1761
rect 2262 1752 2265 1758
rect 2478 1752 2481 1758
rect 290 1748 318 1751
rect 394 1748 446 1751
rect 450 1748 454 1751
rect 490 1748 518 1751
rect 530 1748 566 1751
rect 666 1748 750 1751
rect 818 1748 822 1751
rect 842 1748 846 1751
rect 978 1748 1102 1751
rect 1114 1748 1118 1751
rect 1186 1748 1190 1751
rect 1234 1748 1318 1751
rect 1322 1748 1382 1751
rect 1386 1748 1470 1751
rect 1506 1748 1526 1751
rect 1610 1748 1678 1751
rect 1834 1748 1870 1751
rect 2002 1748 2142 1751
rect 2306 1748 2310 1751
rect 2370 1748 2430 1751
rect 2486 1751 2489 1758
rect 2486 1748 2558 1751
rect 86 1741 89 1748
rect 470 1742 473 1748
rect 86 1738 134 1741
rect 138 1738 174 1741
rect 242 1738 310 1741
rect 314 1738 334 1741
rect 338 1738 390 1741
rect 402 1738 406 1741
rect 530 1738 542 1741
rect 626 1738 670 1741
rect 690 1738 766 1741
rect 798 1741 801 1748
rect 798 1738 854 1741
rect 954 1738 1078 1741
rect 1082 1738 1134 1741
rect 1250 1738 1310 1741
rect 1370 1738 1454 1741
rect 1482 1738 1486 1741
rect 1714 1738 1758 1741
rect 1902 1741 1905 1748
rect 1902 1738 1918 1741
rect 1974 1741 1977 1748
rect 2230 1742 2233 1748
rect 2246 1742 2249 1748
rect 1922 1738 1977 1741
rect 1994 1738 2118 1741
rect 2122 1738 2185 1741
rect 2282 1738 2310 1741
rect 2442 1738 2486 1741
rect 2490 1738 2494 1741
rect 2678 1741 2682 1742
rect 2642 1738 2682 1741
rect 2182 1732 2185 1738
rect 218 1728 358 1731
rect 378 1728 414 1731
rect 418 1728 846 1731
rect 1034 1728 1038 1731
rect 1106 1728 1158 1731
rect 1162 1728 1166 1731
rect 1186 1728 1278 1731
rect 1298 1728 1326 1731
rect 1330 1728 1366 1731
rect 1482 1728 1502 1731
rect 1530 1728 1678 1731
rect 1778 1728 1822 1731
rect 1994 1728 2094 1731
rect 2114 1728 2142 1731
rect 2242 1728 2294 1731
rect 2298 1728 2350 1731
rect 18 1718 278 1721
rect 426 1718 486 1721
rect 498 1718 550 1721
rect 586 1718 822 1721
rect 830 1718 838 1721
rect 842 1718 1118 1721
rect 1594 1718 1750 1721
rect 2066 1718 2070 1721
rect 2202 1718 2270 1721
rect 2274 1718 2342 1721
rect 2358 1721 2361 1728
rect 2446 1722 2449 1728
rect 2358 1718 2374 1721
rect 98 1708 158 1711
rect 258 1708 366 1711
rect 370 1708 406 1711
rect 458 1708 534 1711
rect 538 1708 686 1711
rect 690 1708 694 1711
rect 698 1708 710 1711
rect 810 1708 886 1711
rect 1250 1708 1270 1711
rect 1274 1708 1734 1711
rect 1738 1708 1814 1711
rect 1826 1708 1846 1711
rect 2342 1711 2345 1718
rect 2342 1708 2438 1711
rect 2450 1708 2510 1711
rect 1046 1702 1049 1708
rect 1056 1703 1058 1707
rect 1062 1703 1065 1707
rect 1070 1703 1072 1707
rect 2022 1702 2025 1708
rect 2080 1703 2082 1707
rect 2086 1703 2089 1707
rect 2094 1703 2096 1707
rect 154 1698 158 1701
rect 162 1698 606 1701
rect 714 1698 726 1701
rect 1138 1698 1462 1701
rect 1586 1698 1798 1701
rect 2130 1698 2166 1701
rect 2346 1698 2446 1701
rect 258 1688 390 1691
rect 490 1688 502 1691
rect 702 1691 705 1698
rect 650 1688 705 1691
rect 858 1688 1174 1691
rect 1202 1688 1206 1691
rect 1530 1688 1614 1691
rect 1674 1688 1718 1691
rect 1754 1688 1782 1691
rect 1790 1688 1798 1691
rect 1802 1688 1894 1691
rect 1930 1688 1934 1691
rect 1958 1688 1966 1691
rect 1970 1688 2110 1691
rect 2138 1688 2222 1691
rect 2314 1688 2406 1691
rect 2410 1688 2473 1691
rect 2594 1688 2614 1691
rect 1214 1682 1217 1688
rect 2470 1682 2473 1688
rect 82 1678 345 1681
rect 370 1678 374 1681
rect 394 1678 857 1681
rect 866 1678 926 1681
rect 970 1678 982 1681
rect 1050 1678 1190 1681
rect 1362 1678 1398 1681
rect 1498 1678 1598 1681
rect 1602 1678 1878 1681
rect 1882 1678 1966 1681
rect 2058 1678 2150 1681
rect 342 1672 345 1678
rect 42 1668 126 1671
rect 146 1668 206 1671
rect 210 1668 302 1671
rect 374 1671 377 1678
rect 374 1668 390 1671
rect 522 1668 526 1671
rect 854 1671 857 1678
rect 854 1668 958 1671
rect 1090 1668 1158 1671
rect 1162 1668 1169 1671
rect 1230 1671 1233 1678
rect 1202 1668 1270 1671
rect 1330 1668 1390 1671
rect 1406 1671 1409 1678
rect 1430 1671 1433 1678
rect 2382 1672 2385 1678
rect 1406 1668 1433 1671
rect 1450 1668 1505 1671
rect 1546 1668 1798 1671
rect 1834 1668 1862 1671
rect 1902 1668 1998 1671
rect 2042 1668 2102 1671
rect 2394 1668 2422 1671
rect 2578 1668 2582 1671
rect 2614 1671 2617 1678
rect 2678 1671 2682 1672
rect 2614 1668 2682 1671
rect 1502 1662 1505 1668
rect 1870 1662 1873 1668
rect 1902 1662 1905 1668
rect 2014 1662 2017 1668
rect 122 1658 150 1661
rect 154 1658 334 1661
rect 354 1658 374 1661
rect 402 1658 454 1661
rect 522 1658 590 1661
rect 678 1658 686 1661
rect 690 1658 750 1661
rect 770 1658 870 1661
rect 934 1658 942 1661
rect 946 1658 950 1661
rect 970 1658 998 1661
rect 1010 1658 1142 1661
rect 1154 1658 1257 1661
rect 1290 1658 1366 1661
rect 1402 1658 1438 1661
rect 1474 1658 1478 1661
rect 1570 1658 1590 1661
rect 1898 1658 1902 1661
rect 1954 1658 1958 1661
rect 2118 1661 2121 1668
rect 2118 1658 2166 1661
rect 2206 1661 2209 1668
rect 2178 1658 2209 1661
rect 2246 1661 2249 1668
rect 2246 1658 2318 1661
rect 2422 1658 2430 1661
rect 2434 1658 2518 1661
rect 66 1648 166 1651
rect 210 1648 278 1651
rect 346 1648 358 1651
rect 362 1648 382 1651
rect 386 1648 670 1651
rect 674 1648 694 1651
rect 770 1648 846 1651
rect 886 1651 889 1658
rect 990 1652 993 1658
rect 1254 1652 1257 1658
rect 886 1648 985 1651
rect 1210 1648 1222 1651
rect 1434 1648 1486 1651
rect 1514 1648 1526 1651
rect 1542 1651 1545 1658
rect 1638 1652 1641 1658
rect 1686 1652 1689 1658
rect 1694 1652 1697 1658
rect 1718 1652 1721 1658
rect 1542 1648 1598 1651
rect 1742 1651 1745 1658
rect 1766 1652 1769 1658
rect 1942 1652 1945 1658
rect 2350 1652 2353 1658
rect 1742 1648 1750 1651
rect 1778 1648 1806 1651
rect 1954 1648 2006 1651
rect 2010 1648 2062 1651
rect 2434 1648 2454 1651
rect 2458 1648 2462 1651
rect 2678 1651 2682 1652
rect 2650 1648 2682 1651
rect 982 1641 985 1648
rect 982 1638 998 1641
rect 1298 1638 1422 1641
rect 1950 1641 1953 1648
rect 1482 1638 1953 1641
rect 2002 1638 2110 1641
rect 2230 1641 2233 1648
rect 2122 1638 2233 1641
rect 2298 1638 2566 1641
rect 2570 1638 2574 1641
rect 770 1628 950 1631
rect 974 1631 977 1638
rect 974 1628 1430 1631
rect 1450 1628 1534 1631
rect 1626 1628 1662 1631
rect 1818 1628 1934 1631
rect 1970 1628 2134 1631
rect 2170 1628 2262 1631
rect 2274 1628 2502 1631
rect 586 1618 1062 1621
rect 1418 1618 1454 1621
rect 1522 1618 1902 1621
rect 1994 1618 2214 1621
rect 2226 1618 2262 1621
rect 2418 1618 2622 1621
rect 850 1608 1038 1611
rect 1698 1608 1814 1611
rect 1826 1608 2246 1611
rect 2402 1608 2510 1611
rect 544 1603 546 1607
rect 550 1603 553 1607
rect 558 1603 560 1607
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1574 1603 1576 1607
rect 698 1598 982 1601
rect 1034 1598 1350 1601
rect 1354 1598 1398 1601
rect 1634 1598 1766 1601
rect 1890 1598 2070 1601
rect 2114 1598 2302 1601
rect 490 1588 590 1591
rect 594 1588 1590 1591
rect 1714 1588 1766 1591
rect 1930 1588 2014 1591
rect 2018 1588 2230 1591
rect 258 1578 566 1581
rect 570 1578 582 1581
rect 890 1578 910 1581
rect 1002 1578 1246 1581
rect 1266 1578 1294 1581
rect 1554 1578 1654 1581
rect 1658 1578 1790 1581
rect 1938 1578 1958 1581
rect 2026 1578 2310 1581
rect 754 1568 798 1571
rect 874 1568 1022 1571
rect 1210 1568 1278 1571
rect 1426 1568 1446 1571
rect 1474 1568 1486 1571
rect 1490 1568 1566 1571
rect 1578 1568 1702 1571
rect 1866 1568 1870 1571
rect 1970 1568 2150 1571
rect 2210 1568 2278 1571
rect 2506 1568 2550 1571
rect 130 1558 382 1561
rect 454 1561 457 1568
rect 454 1558 486 1561
rect 490 1558 598 1561
rect 690 1558 822 1561
rect 1274 1558 1278 1561
rect 1362 1558 1454 1561
rect 1474 1558 1494 1561
rect 1498 1558 1646 1561
rect 1650 1558 1686 1561
rect 1862 1561 1865 1568
rect 1730 1558 1865 1561
rect 1950 1561 1953 1568
rect 1950 1558 2014 1561
rect 2058 1558 2078 1561
rect 2242 1558 2254 1561
rect 2306 1558 2350 1561
rect 418 1548 430 1551
rect 434 1548 438 1551
rect 478 1548 494 1551
rect 538 1548 646 1551
rect 650 1548 750 1551
rect 818 1548 838 1551
rect 842 1548 854 1551
rect 994 1548 1014 1551
rect 1018 1548 1038 1551
rect 1066 1548 1110 1551
rect 1114 1548 1302 1551
rect 1306 1548 1358 1551
rect 1370 1548 1422 1551
rect 1426 1548 1502 1551
rect 190 1541 193 1548
rect 206 1541 209 1548
rect 478 1542 481 1548
rect 790 1542 793 1548
rect 894 1542 897 1548
rect 1602 1548 1670 1551
rect 1706 1548 1710 1551
rect 1762 1548 1766 1551
rect 1874 1548 1942 1551
rect 1970 1548 2006 1551
rect 2034 1548 2038 1551
rect 2062 1548 2070 1551
rect 2158 1551 2161 1558
rect 2238 1551 2241 1558
rect 2590 1552 2593 1558
rect 2074 1548 2161 1551
rect 2166 1548 2241 1551
rect 2318 1548 2422 1551
rect 2466 1548 2494 1551
rect 2498 1548 2518 1551
rect 2522 1548 2542 1551
rect 2546 1548 2550 1551
rect 190 1538 209 1541
rect 322 1538 478 1541
rect 522 1538 582 1541
rect 802 1538 862 1541
rect 938 1538 1062 1541
rect 1098 1538 1102 1541
rect 1126 1538 1142 1541
rect 1162 1538 1206 1541
rect 1210 1538 1294 1541
rect 1314 1538 1422 1541
rect 1426 1538 1670 1541
rect 1706 1538 1742 1541
rect 2166 1541 2169 1548
rect 1770 1538 2169 1541
rect 2318 1542 2321 1548
rect 2482 1538 2486 1541
rect 2530 1538 2598 1541
rect 234 1528 425 1531
rect 810 1528 910 1531
rect 1126 1531 1129 1538
rect 1050 1528 1129 1531
rect 1138 1528 1145 1531
rect 1226 1528 1334 1531
rect 1442 1528 1646 1531
rect 1702 1528 1734 1531
rect 1754 1528 2014 1531
rect 2018 1528 2038 1531
rect 2074 1528 2086 1531
rect 2146 1528 2174 1531
rect 2202 1528 2382 1531
rect 2426 1528 2550 1531
rect 422 1522 425 1528
rect 298 1518 390 1521
rect 602 1518 694 1521
rect 698 1518 902 1521
rect 922 1518 1134 1521
rect 1142 1521 1145 1528
rect 1414 1522 1417 1528
rect 1702 1522 1705 1528
rect 1142 1518 1366 1521
rect 1434 1518 1598 1521
rect 1602 1518 1670 1521
rect 1874 1518 1918 1521
rect 2250 1518 2262 1521
rect 458 1508 662 1511
rect 850 1508 966 1511
rect 1114 1508 1214 1511
rect 1266 1508 1318 1511
rect 1442 1508 1446 1511
rect 1458 1508 1494 1511
rect 1538 1508 1550 1511
rect 1586 1508 1622 1511
rect 1690 1508 1926 1511
rect 2242 1508 2254 1511
rect 2258 1508 2270 1511
rect 2362 1508 2470 1511
rect 1056 1503 1058 1507
rect 1062 1503 1065 1507
rect 1070 1503 1072 1507
rect 2080 1503 2082 1507
rect 2086 1503 2089 1507
rect 2094 1503 2096 1507
rect 106 1498 158 1501
rect 394 1498 742 1501
rect 762 1498 782 1501
rect 786 1498 854 1501
rect 890 1498 918 1501
rect 1146 1498 1222 1501
rect 1386 1498 1670 1501
rect 1818 1498 1870 1501
rect 1874 1498 1990 1501
rect 2282 1498 2414 1501
rect 106 1488 182 1491
rect 394 1488 670 1491
rect 850 1488 1102 1491
rect 1130 1488 1334 1491
rect 1338 1488 1606 1491
rect 1690 1488 1694 1491
rect 1834 1488 2046 1491
rect 2414 1491 2417 1498
rect 2414 1488 2446 1491
rect 2474 1488 2494 1491
rect 42 1478 105 1481
rect 138 1478 238 1481
rect 522 1478 998 1481
rect 1042 1478 1118 1481
rect 1154 1478 1182 1481
rect 1266 1478 1270 1481
rect 1290 1478 1318 1481
rect 1322 1478 1462 1481
rect 1466 1478 1470 1481
rect 1482 1478 1542 1481
rect 1626 1478 1918 1481
rect 1930 1478 2070 1481
rect 2178 1478 2334 1481
rect 2442 1478 2478 1481
rect 2482 1478 2598 1481
rect 2602 1478 2638 1481
rect 102 1472 105 1478
rect 146 1468 150 1471
rect 182 1468 190 1471
rect 194 1468 198 1471
rect 242 1468 414 1471
rect 418 1468 470 1471
rect 486 1468 505 1471
rect 586 1468 654 1471
rect 658 1468 718 1471
rect 802 1468 806 1471
rect 970 1468 1094 1471
rect 1330 1468 1342 1471
rect 1410 1468 1454 1471
rect 1458 1468 1590 1471
rect 1594 1468 1606 1471
rect 1610 1468 1614 1471
rect 1682 1468 1750 1471
rect 2002 1468 2038 1471
rect 2050 1468 2150 1471
rect 2314 1468 2318 1471
rect 2386 1468 2414 1471
rect 2450 1468 2558 1471
rect 486 1462 489 1468
rect 502 1462 505 1468
rect 138 1458 166 1461
rect 186 1458 190 1461
rect 370 1458 390 1461
rect 538 1458 630 1461
rect 710 1458 718 1461
rect 722 1458 750 1461
rect 822 1461 825 1468
rect 822 1458 870 1461
rect 930 1458 934 1461
rect 978 1458 982 1461
rect 1010 1458 1014 1461
rect 1130 1458 1134 1461
rect 1194 1458 1262 1461
rect 1362 1458 1422 1461
rect 1450 1458 1630 1461
rect 1794 1458 1822 1461
rect 1826 1458 1854 1461
rect 1930 1459 1982 1461
rect 1926 1458 1982 1459
rect 2030 1458 2046 1461
rect 2254 1461 2257 1468
rect 2106 1458 2193 1461
rect 2254 1458 2470 1461
rect 710 1452 713 1458
rect 1486 1452 1489 1458
rect 2006 1452 2009 1458
rect 2030 1452 2033 1458
rect 2190 1452 2193 1458
rect 42 1448 145 1451
rect 354 1448 406 1451
rect 618 1448 638 1451
rect 666 1448 702 1451
rect 754 1448 1006 1451
rect 1026 1448 1070 1451
rect 1074 1448 1350 1451
rect 1434 1448 1470 1451
rect 1586 1448 1590 1451
rect 1610 1448 1822 1451
rect 1826 1448 1878 1451
rect 1938 1448 1974 1451
rect 2042 1448 2094 1451
rect 2434 1448 2446 1451
rect 2450 1448 2486 1451
rect 2678 1451 2682 1452
rect 2650 1448 2682 1451
rect 142 1442 145 1448
rect 614 1441 617 1448
rect 170 1438 617 1441
rect 818 1438 998 1441
rect 1002 1438 1038 1441
rect 1042 1438 1078 1441
rect 1210 1438 1214 1441
rect 1226 1438 1390 1441
rect 1426 1438 1430 1441
rect 1466 1438 1510 1441
rect 1626 1438 1630 1441
rect 1634 1438 1726 1441
rect 1730 1438 1966 1441
rect 1970 1438 2286 1441
rect 2290 1438 2310 1441
rect 378 1428 526 1431
rect 530 1428 606 1431
rect 714 1428 1022 1431
rect 1210 1428 1430 1431
rect 1602 1428 1710 1431
rect 1714 1428 1774 1431
rect 2034 1428 2262 1431
rect 2610 1428 2630 1431
rect 170 1418 270 1421
rect 274 1418 310 1421
rect 314 1418 726 1421
rect 842 1418 846 1421
rect 1002 1418 1342 1421
rect 1346 1418 1406 1421
rect 1430 1421 1433 1428
rect 1430 1418 1486 1421
rect 1522 1418 1542 1421
rect 1546 1418 1614 1421
rect 1754 1418 1790 1421
rect 1810 1418 2062 1421
rect 2082 1418 2422 1421
rect 98 1408 222 1411
rect 1026 1408 1182 1411
rect 1186 1408 1358 1411
rect 1362 1408 1382 1411
rect 1386 1408 1462 1411
rect 1498 1408 1550 1411
rect 1690 1408 1830 1411
rect 1970 1408 1982 1411
rect 2066 1408 2118 1411
rect 2194 1408 2606 1411
rect 544 1403 546 1407
rect 550 1403 553 1407
rect 558 1403 560 1407
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1574 1403 1576 1407
rect 882 1398 1070 1401
rect 1322 1398 1326 1401
rect 1402 1398 1454 1401
rect 1466 1398 1550 1401
rect 1794 1398 1806 1401
rect 1826 1398 1950 1401
rect 1954 1398 2110 1401
rect 890 1388 910 1391
rect 1378 1388 1478 1391
rect 1482 1388 1502 1391
rect 1558 1388 1582 1391
rect 1658 1388 1678 1391
rect 1682 1388 2078 1391
rect 2082 1388 2542 1391
rect 2678 1391 2682 1392
rect 2650 1388 2682 1391
rect 202 1378 334 1381
rect 1038 1381 1041 1388
rect 1558 1382 1561 1388
rect 730 1378 1041 1381
rect 1378 1378 1398 1381
rect 1402 1378 1550 1381
rect 1826 1378 2294 1381
rect 282 1368 286 1371
rect 298 1368 334 1371
rect 610 1368 862 1371
rect 866 1368 902 1371
rect 1050 1368 1054 1371
rect 1202 1368 1406 1371
rect 1410 1368 1454 1371
rect 1514 1368 1734 1371
rect 1790 1371 1793 1378
rect 1790 1368 1838 1371
rect 1842 1368 2102 1371
rect 2114 1368 2414 1371
rect 2570 1368 2582 1371
rect 2678 1371 2682 1372
rect 2594 1368 2682 1371
rect 122 1358 142 1361
rect 146 1358 430 1361
rect 566 1361 569 1368
rect 482 1358 569 1361
rect 858 1358 862 1361
rect 998 1361 1001 1368
rect 1782 1362 1785 1368
rect 890 1358 1001 1361
rect 1010 1358 1070 1361
rect 1074 1358 1078 1361
rect 1082 1358 1102 1361
rect 1218 1358 1246 1361
rect 1250 1358 1310 1361
rect 1314 1358 1486 1361
rect 1490 1358 1526 1361
rect 1650 1358 1686 1361
rect 1786 1358 1806 1361
rect 1842 1358 1934 1361
rect 1946 1358 1974 1361
rect 1978 1358 1998 1361
rect 2074 1358 2126 1361
rect 2162 1358 2166 1361
rect 2210 1358 2382 1361
rect 2434 1358 2577 1361
rect 50 1348 126 1351
rect 218 1348 230 1351
rect 258 1348 566 1351
rect 570 1348 630 1351
rect 634 1348 726 1351
rect 826 1348 862 1351
rect 1010 1348 1014 1351
rect 1026 1348 1062 1351
rect 1066 1348 1086 1351
rect 1098 1348 1118 1351
rect 1154 1348 1230 1351
rect 1258 1348 1326 1351
rect 1370 1348 1446 1351
rect 1450 1348 1470 1351
rect 1474 1348 1550 1351
rect 1554 1348 1638 1351
rect 1666 1348 1998 1351
rect 2002 1348 2014 1351
rect 2026 1348 2038 1351
rect 2058 1348 2126 1351
rect 2174 1351 2177 1358
rect 2574 1352 2577 1358
rect 2162 1348 2177 1351
rect 2194 1348 2198 1351
rect 2502 1348 2553 1351
rect 2678 1351 2682 1352
rect 2610 1348 2682 1351
rect 306 1338 310 1341
rect 322 1338 382 1341
rect 386 1338 534 1341
rect 538 1338 550 1341
rect 666 1338 1158 1341
rect 1162 1338 1214 1341
rect 1218 1338 1265 1341
rect 1290 1338 1358 1341
rect 1386 1338 1390 1341
rect 1398 1338 1438 1341
rect 1458 1338 1494 1341
rect 1530 1338 1649 1341
rect 1658 1338 1662 1341
rect 1674 1338 1718 1341
rect 1722 1338 1833 1341
rect 2002 1338 2022 1341
rect 2090 1338 2110 1341
rect 2146 1338 2270 1341
rect 2318 1341 2321 1348
rect 2502 1342 2505 1348
rect 2550 1342 2553 1348
rect 2318 1338 2334 1341
rect 2346 1338 2422 1341
rect 2562 1338 2598 1341
rect 1262 1332 1265 1338
rect 1398 1332 1401 1338
rect 1646 1332 1649 1338
rect 226 1328 286 1331
rect 306 1328 406 1331
rect 594 1328 718 1331
rect 722 1328 782 1331
rect 1034 1328 1038 1331
rect 1074 1328 1078 1331
rect 1098 1328 1158 1331
rect 1162 1328 1166 1331
rect 1202 1328 1254 1331
rect 1434 1328 1478 1331
rect 1498 1328 1542 1331
rect 1570 1328 1606 1331
rect 1618 1328 1622 1331
rect 1626 1328 1638 1331
rect 1650 1328 1670 1331
rect 1830 1331 1833 1338
rect 1830 1328 1942 1331
rect 1978 1328 2014 1331
rect 2022 1328 2030 1331
rect 2034 1328 2046 1331
rect 2194 1328 2222 1331
rect 2410 1328 2534 1331
rect 2538 1328 2574 1331
rect 2578 1328 2582 1331
rect 306 1318 454 1321
rect 986 1318 1278 1321
rect 1434 1318 1814 1321
rect 2678 1321 2682 1322
rect 2642 1318 2682 1321
rect 322 1308 326 1311
rect 418 1308 982 1311
rect 1082 1308 1102 1311
rect 1210 1308 1254 1311
rect 1298 1308 1446 1311
rect 1450 1308 1590 1311
rect 1610 1308 1670 1311
rect 1762 1308 1766 1311
rect 1810 1308 1870 1311
rect 1906 1308 1998 1311
rect 2034 1308 2070 1311
rect 1056 1303 1058 1307
rect 1062 1303 1065 1307
rect 1070 1303 1072 1307
rect 2080 1303 2082 1307
rect 2086 1303 2089 1307
rect 2094 1303 2096 1307
rect 218 1298 382 1301
rect 426 1298 446 1301
rect 450 1298 702 1301
rect 730 1298 902 1301
rect 1034 1298 1038 1301
rect 1098 1298 1198 1301
rect 1578 1298 1646 1301
rect 2678 1301 2682 1302
rect 2650 1298 2682 1301
rect 166 1288 174 1291
rect 178 1288 190 1291
rect 250 1288 294 1291
rect 314 1288 470 1291
rect 474 1288 558 1291
rect 562 1288 670 1291
rect 690 1288 718 1291
rect 722 1288 1014 1291
rect 1018 1288 1022 1291
rect 1030 1288 1038 1291
rect 1042 1288 1310 1291
rect 1418 1288 1462 1291
rect 1466 1288 1478 1291
rect 1534 1288 1550 1291
rect 1586 1288 1630 1291
rect 1658 1288 1702 1291
rect 1722 1288 1822 1291
rect 2038 1288 2046 1291
rect 2050 1288 2078 1291
rect 2098 1288 2102 1291
rect 2234 1288 2238 1291
rect 2266 1288 2505 1291
rect 2578 1288 2622 1291
rect 302 1282 305 1288
rect 154 1278 174 1281
rect 178 1278 222 1281
rect 226 1278 262 1281
rect 370 1278 422 1281
rect 450 1278 454 1281
rect 554 1278 630 1281
rect 722 1278 726 1281
rect 786 1278 806 1281
rect 810 1278 822 1281
rect 850 1278 862 1281
rect 866 1278 878 1281
rect 930 1278 1150 1281
rect 1282 1278 1326 1281
rect 1426 1278 1446 1281
rect 1534 1281 1537 1288
rect 2502 1282 2505 1288
rect 1458 1278 1537 1281
rect 1546 1278 1694 1281
rect 1714 1278 1806 1281
rect 1902 1278 1942 1281
rect 1946 1278 2022 1281
rect 2330 1278 2374 1281
rect 2586 1278 2646 1281
rect 2678 1281 2682 1282
rect 2650 1278 2682 1281
rect 186 1268 230 1271
rect 386 1268 390 1271
rect 394 1268 406 1271
rect 426 1268 502 1271
rect 546 1268 654 1271
rect 670 1271 673 1278
rect 670 1268 857 1271
rect 866 1268 886 1271
rect 1042 1268 1046 1271
rect 1114 1268 1118 1271
rect 1178 1268 1302 1271
rect 1330 1268 1502 1271
rect 1522 1268 1574 1271
rect 1602 1268 1646 1271
rect 1802 1268 1830 1271
rect 1902 1271 1905 1278
rect 2302 1272 2305 1278
rect 2398 1272 2401 1278
rect 1850 1268 1905 1271
rect 2002 1268 2006 1271
rect 2498 1268 2598 1271
rect 122 1258 190 1261
rect 270 1261 273 1268
rect 854 1262 857 1268
rect 270 1258 310 1261
rect 330 1258 398 1261
rect 442 1258 678 1261
rect 786 1258 790 1261
rect 794 1258 846 1261
rect 874 1258 894 1261
rect 1178 1258 1182 1261
rect 1202 1258 1297 1261
rect 1362 1258 1438 1261
rect 1466 1258 1478 1261
rect 1482 1258 1582 1261
rect 1654 1261 1657 1268
rect 1798 1262 1801 1268
rect 1642 1258 1657 1261
rect 1682 1258 1718 1261
rect 1838 1261 1841 1268
rect 1810 1258 1841 1261
rect 1910 1261 1913 1268
rect 1910 1258 1958 1261
rect 2050 1258 2054 1261
rect 2114 1258 2118 1261
rect 2138 1258 2366 1261
rect 2482 1258 2550 1261
rect 870 1252 873 1258
rect 202 1248 214 1251
rect 330 1248 478 1251
rect 486 1248 526 1251
rect 538 1248 598 1251
rect 602 1248 614 1251
rect 658 1248 662 1251
rect 746 1248 862 1251
rect 1058 1248 1078 1251
rect 1090 1248 1094 1251
rect 1134 1251 1137 1258
rect 1294 1252 1297 1258
rect 1134 1248 1158 1251
rect 1202 1248 1206 1251
rect 1210 1248 1278 1251
rect 1450 1248 1542 1251
rect 1682 1248 1686 1251
rect 1782 1251 1785 1258
rect 2062 1252 2065 1258
rect 1714 1248 1966 1251
rect 1970 1248 2062 1251
rect 2118 1251 2121 1258
rect 2118 1248 2182 1251
rect 2378 1248 2438 1251
rect 2458 1248 2470 1251
rect 2678 1251 2682 1252
rect 2634 1248 2682 1251
rect 486 1242 489 1248
rect 454 1238 478 1241
rect 650 1238 670 1241
rect 674 1238 798 1241
rect 802 1238 838 1241
rect 842 1238 1166 1241
rect 1182 1241 1185 1248
rect 2470 1242 2473 1248
rect 1170 1238 1185 1241
rect 1314 1238 1430 1241
rect 1450 1238 1598 1241
rect 1770 1238 1854 1241
rect 1994 1238 2062 1241
rect 2322 1238 2334 1241
rect 2338 1238 2446 1241
rect 454 1232 457 1238
rect 466 1228 582 1231
rect 586 1228 646 1231
rect 650 1228 734 1231
rect 738 1228 1094 1231
rect 1106 1228 1142 1231
rect 1146 1228 1190 1231
rect 1194 1228 1254 1231
rect 1258 1228 1470 1231
rect 1610 1228 1662 1231
rect 1714 1228 2214 1231
rect 2218 1228 2446 1231
rect 2450 1228 2470 1231
rect 474 1218 654 1221
rect 730 1218 790 1221
rect 794 1218 801 1221
rect 850 1218 894 1221
rect 1126 1218 1134 1221
rect 1138 1218 1350 1221
rect 1606 1221 1609 1228
rect 1358 1218 1609 1221
rect 1858 1218 2350 1221
rect 2354 1218 2382 1221
rect 802 1208 886 1211
rect 898 1208 918 1211
rect 930 1208 1086 1211
rect 1358 1211 1361 1218
rect 1090 1208 1361 1211
rect 1826 1208 1878 1211
rect 1994 1208 2022 1211
rect 2026 1208 2254 1211
rect 2434 1208 2486 1211
rect 544 1203 546 1207
rect 550 1203 553 1207
rect 558 1203 560 1207
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1574 1203 1576 1207
rect 858 1198 974 1201
rect 1938 1198 2094 1201
rect 2122 1198 2310 1201
rect 1338 1188 1366 1191
rect 1434 1188 1478 1191
rect 2154 1188 2318 1191
rect 2462 1191 2465 1198
rect 2462 1188 2494 1191
rect 2634 1188 2638 1191
rect 470 1182 473 1188
rect 506 1178 518 1181
rect 594 1178 638 1181
rect 850 1178 1262 1181
rect 1266 1178 1462 1181
rect 1498 1178 1542 1181
rect 2090 1178 2374 1181
rect 2390 1181 2393 1188
rect 2378 1178 2393 1181
rect 2426 1178 2478 1181
rect 358 1172 361 1178
rect 122 1168 190 1171
rect 434 1168 862 1171
rect 1346 1168 1350 1171
rect 1370 1168 1438 1171
rect 1442 1168 1518 1171
rect 1562 1168 1622 1171
rect 2058 1168 2438 1171
rect 2562 1168 2566 1171
rect 2678 1171 2682 1172
rect 2618 1168 2682 1171
rect 878 1162 881 1168
rect 1246 1162 1249 1168
rect 1918 1162 1921 1168
rect 186 1158 214 1161
rect 218 1158 462 1161
rect 474 1158 638 1161
rect 642 1158 702 1161
rect 706 1158 742 1161
rect 858 1158 878 1161
rect 906 1158 1030 1161
rect 1330 1158 1398 1161
rect 1490 1158 1566 1161
rect 1570 1158 1590 1161
rect 1594 1158 1614 1161
rect 2082 1158 2150 1161
rect 2274 1158 2310 1161
rect 2314 1158 2326 1161
rect 2454 1161 2457 1168
rect 2454 1158 2518 1161
rect 2574 1158 2681 1161
rect 170 1148 222 1151
rect 226 1148 246 1151
rect 346 1148 377 1151
rect 410 1148 478 1151
rect 538 1148 550 1151
rect 646 1148 654 1151
rect 658 1148 713 1151
rect 746 1148 774 1151
rect 890 1148 926 1151
rect 1014 1148 1046 1151
rect 1202 1148 1278 1151
rect 1294 1151 1297 1158
rect 1294 1148 1302 1151
rect 1306 1148 1318 1151
rect 1330 1148 1374 1151
rect 1490 1148 1494 1151
rect 1506 1148 2022 1151
rect 2026 1148 2030 1151
rect 2122 1148 2142 1151
rect 2146 1148 2174 1151
rect 2234 1148 2302 1151
rect 2354 1148 2406 1151
rect 2574 1151 2577 1158
rect 2678 1152 2681 1158
rect 2426 1148 2577 1151
rect 2586 1148 2590 1151
rect 374 1142 377 1148
rect 710 1142 713 1148
rect 1014 1142 1017 1148
rect 2678 1148 2682 1152
rect 10 1138 14 1141
rect 178 1138 278 1141
rect 298 1138 334 1141
rect 378 1138 390 1141
rect 514 1138 609 1141
rect 690 1138 694 1141
rect 738 1138 758 1141
rect 826 1138 910 1141
rect 1258 1138 1278 1141
rect 1282 1138 1414 1141
rect 1450 1138 1470 1141
rect 1602 1138 1678 1141
rect 1834 1138 1926 1141
rect 2018 1138 2038 1141
rect 2058 1138 2134 1141
rect 2186 1138 2326 1141
rect 2542 1138 2638 1141
rect 606 1132 609 1138
rect 1438 1132 1441 1138
rect 186 1128 198 1131
rect 274 1128 286 1131
rect 290 1128 302 1131
rect 322 1128 366 1131
rect 690 1128 726 1131
rect 754 1128 790 1131
rect 794 1128 910 1131
rect 1106 1128 1398 1131
rect 1426 1128 1438 1131
rect 1474 1128 1878 1131
rect 2358 1131 2361 1138
rect 1954 1128 2361 1131
rect 2366 1131 2369 1138
rect 2542 1132 2545 1138
rect 2366 1128 2414 1131
rect 230 1122 233 1128
rect 250 1118 297 1121
rect 402 1118 430 1121
rect 434 1118 918 1121
rect 930 1118 1438 1121
rect 1506 1118 1870 1121
rect 1878 1121 1881 1128
rect 1878 1118 2102 1121
rect 2106 1118 2350 1121
rect 2458 1118 2574 1121
rect 294 1112 297 1118
rect 338 1108 422 1111
rect 426 1108 518 1111
rect 522 1108 534 1111
rect 546 1108 622 1111
rect 682 1108 782 1111
rect 834 1108 846 1111
rect 850 1108 990 1111
rect 1098 1108 1174 1111
rect 1250 1108 1286 1111
rect 1530 1108 1622 1111
rect 1730 1108 1990 1111
rect 2042 1108 2054 1111
rect 2106 1108 2310 1111
rect 1056 1103 1058 1107
rect 1062 1103 1065 1107
rect 1070 1103 1072 1107
rect 2080 1103 2082 1107
rect 2086 1103 2089 1107
rect 2094 1103 2096 1107
rect 538 1098 574 1101
rect 578 1098 926 1101
rect 1386 1098 1734 1101
rect 1738 1098 1742 1101
rect 146 1088 190 1091
rect 194 1088 302 1091
rect 454 1091 457 1098
rect 2126 1092 2129 1098
rect 346 1088 457 1091
rect 642 1088 678 1091
rect 954 1088 1062 1091
rect 1114 1088 1118 1091
rect 1778 1088 1833 1091
rect 2462 1088 2470 1091
rect 2474 1088 2534 1091
rect 1830 1082 1833 1088
rect 154 1078 174 1081
rect 178 1078 254 1081
rect 258 1078 1038 1081
rect 1106 1078 1134 1081
rect 1138 1078 1446 1081
rect 1490 1078 1606 1081
rect 1650 1078 1678 1081
rect 1874 1078 1886 1081
rect 1890 1078 2046 1081
rect 2050 1078 2062 1081
rect 2098 1078 2230 1081
rect 2266 1078 2278 1081
rect 2326 1081 2329 1088
rect 2306 1078 2329 1081
rect 2410 1078 2422 1081
rect 2426 1078 2574 1081
rect 2578 1078 2614 1081
rect 1630 1072 1633 1078
rect 34 1068 209 1071
rect 206 1062 209 1068
rect 334 1068 414 1071
rect 722 1068 774 1071
rect 842 1068 894 1071
rect 1162 1068 1326 1071
rect 1370 1068 1414 1071
rect 1418 1068 1446 1071
rect 1554 1068 1606 1071
rect 1642 1068 1654 1071
rect 1790 1071 1793 1078
rect 1790 1068 1998 1071
rect 2002 1068 2190 1071
rect 2194 1068 2398 1071
rect 2402 1068 2510 1071
rect 334 1062 337 1068
rect 90 1058 166 1061
rect 654 1058 670 1061
rect 714 1058 726 1061
rect 730 1058 854 1061
rect 874 1058 886 1061
rect 894 1061 897 1068
rect 1342 1062 1345 1068
rect 894 1058 998 1061
rect 1122 1058 1246 1061
rect 1386 1058 1534 1061
rect 1558 1058 1598 1061
rect 1634 1058 1646 1061
rect 1666 1058 1670 1061
rect 1826 1058 1838 1061
rect 1890 1058 1966 1061
rect 2098 1058 2126 1061
rect 2234 1058 2262 1061
rect 2266 1058 2302 1061
rect 2386 1059 2441 1061
rect 2382 1058 2441 1059
rect 2450 1058 2622 1061
rect -26 1051 -22 1052
rect -26 1048 6 1051
rect 374 1051 377 1058
rect 654 1052 657 1058
rect 374 1048 510 1051
rect 746 1048 838 1051
rect 866 1048 886 1051
rect 898 1048 934 1051
rect 1026 1048 1262 1051
rect 1318 1051 1321 1058
rect 1558 1052 1561 1058
rect 2438 1052 2441 1058
rect 1318 1048 1350 1051
rect 1434 1048 1446 1051
rect 1674 1048 1686 1051
rect 1698 1048 1830 1051
rect 2066 1048 2126 1051
rect 2130 1048 2254 1051
rect 2306 1048 2430 1051
rect 2602 1048 2606 1051
rect 2678 1051 2682 1052
rect 2650 1048 2682 1051
rect 418 1038 430 1041
rect 1022 1041 1025 1048
rect 594 1038 1025 1041
rect 1042 1038 1094 1041
rect 1098 1038 1270 1041
rect 1322 1038 1374 1041
rect 1594 1038 1646 1041
rect 1722 1038 1806 1041
rect 1826 1038 1870 1041
rect 1874 1038 1894 1041
rect 2130 1038 2294 1041
rect 590 1031 593 1038
rect 26 1028 593 1031
rect 914 1028 942 1031
rect 946 1028 1454 1031
rect 1850 1028 1862 1031
rect 2002 1028 2070 1031
rect 2114 1028 2302 1031
rect 762 1018 926 1021
rect 1042 1018 1254 1021
rect 1258 1018 1494 1021
rect 1578 1018 1782 1021
rect 1946 1018 2006 1021
rect 2066 1018 2078 1021
rect 2114 1018 2134 1021
rect 2314 1018 2374 1021
rect 1250 1008 1302 1011
rect 1314 1008 1542 1011
rect 1706 1008 1998 1011
rect 2002 1008 2118 1011
rect 2282 1008 2398 1011
rect 544 1003 546 1007
rect 550 1003 553 1007
rect 558 1003 560 1007
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1574 1003 1576 1007
rect 122 998 142 1001
rect 146 998 470 1001
rect 802 998 806 1001
rect 994 998 1174 1001
rect 1178 998 1278 1001
rect 1458 998 1510 1001
rect 2322 998 2382 1001
rect 194 988 294 991
rect 298 988 414 991
rect 418 988 566 991
rect 570 988 678 991
rect 682 988 870 991
rect 874 988 1294 991
rect 1298 988 1614 991
rect 2678 991 2682 992
rect 1618 988 1977 991
rect 1974 982 1977 988
rect 2566 988 2682 991
rect 2566 982 2569 988
rect 346 978 366 981
rect 370 978 582 981
rect 586 978 710 981
rect 906 978 950 981
rect 1290 978 1326 981
rect 1378 978 1414 981
rect 2018 978 2270 981
rect 106 968 166 971
rect 706 968 822 971
rect 1154 968 1238 971
rect 1266 968 1342 971
rect 1346 968 1502 971
rect 1762 968 1854 971
rect 1858 968 1958 971
rect 2190 968 2198 971
rect 2202 968 2278 971
rect 2282 968 2550 971
rect 2678 971 2682 972
rect 2650 968 2682 971
rect 266 958 350 961
rect 410 958 422 961
rect 466 958 478 961
rect 638 958 646 961
rect 650 958 710 961
rect 1394 958 1414 961
rect 1510 961 1513 968
rect 1426 958 1513 961
rect 1546 958 1598 961
rect 1730 958 1750 961
rect 1938 958 2486 961
rect 2490 958 2502 961
rect 158 952 161 958
rect 918 952 921 958
rect 1286 952 1289 958
rect 66 948 158 951
rect 226 948 278 951
rect 282 948 326 951
rect 330 948 702 951
rect 962 948 1041 951
rect 1138 948 1185 951
rect 1290 948 1310 951
rect 1394 948 1438 951
rect 1506 948 1526 951
rect 1570 948 1574 951
rect 1658 948 1726 951
rect 1806 951 1809 958
rect 1806 948 1814 951
rect 1846 948 1862 951
rect 1882 948 1918 951
rect 1970 948 1982 951
rect 1986 948 2014 951
rect 2018 948 2025 951
rect 2274 948 2310 951
rect 2394 948 2510 951
rect 2530 948 2574 951
rect 2678 951 2682 952
rect 2594 948 2682 951
rect 58 938 118 941
rect 162 938 286 941
rect 290 938 390 941
rect 482 938 582 941
rect 706 938 710 941
rect 734 941 737 948
rect 750 941 753 948
rect 1038 942 1041 948
rect 1182 942 1185 948
rect 734 938 753 941
rect 826 938 902 941
rect 1402 938 1422 941
rect 1514 938 1558 941
rect 1626 938 1646 941
rect 1766 941 1769 948
rect 1650 938 1769 941
rect 1846 942 1849 948
rect 1898 938 1910 941
rect 1930 938 2182 941
rect 2186 938 2366 941
rect 2370 938 2598 941
rect 242 928 246 931
rect 394 928 590 931
rect 594 928 638 931
rect 650 928 750 931
rect 882 928 974 931
rect 1066 928 1198 931
rect 1386 928 1486 931
rect 1490 928 1518 931
rect 2210 928 2334 931
rect 2338 928 2454 931
rect 2466 928 2537 931
rect 2554 928 2582 931
rect 106 918 438 921
rect 786 918 894 921
rect 898 918 1038 921
rect 1194 918 1302 921
rect 1482 918 1638 921
rect 1770 918 1846 921
rect 1874 918 1878 921
rect 1882 918 1902 921
rect 2006 921 2009 928
rect 2534 922 2537 928
rect 1906 918 2009 921
rect 2090 918 2118 921
rect 2218 918 2342 921
rect 418 908 454 911
rect 458 908 646 911
rect 754 908 926 911
rect 930 908 982 911
rect 986 908 1030 911
rect 1202 908 1430 911
rect 1682 908 1822 911
rect 1842 908 1942 911
rect 2162 908 2414 911
rect 2418 908 2518 911
rect 1056 903 1058 907
rect 1062 903 1065 907
rect 1070 903 1072 907
rect 2080 903 2082 907
rect 2086 903 2089 907
rect 2094 903 2096 907
rect 602 898 622 901
rect 794 898 838 901
rect 1154 898 1214 901
rect 1218 898 1382 901
rect 1602 898 1638 901
rect 1890 898 1918 901
rect 1962 898 2046 901
rect 2202 898 2230 901
rect 2378 898 2398 901
rect 2402 898 2622 901
rect 178 888 198 891
rect 490 888 766 891
rect 834 888 918 891
rect 922 888 926 891
rect 1242 888 1358 891
rect 1594 888 1734 891
rect 1738 888 1742 891
rect 1778 888 1782 891
rect 1946 888 1974 891
rect 1994 888 2318 891
rect 806 882 809 888
rect 530 878 606 881
rect 610 878 718 881
rect 1002 878 1054 881
rect 1354 878 1446 881
rect 1466 878 1494 881
rect 1498 878 1822 881
rect 1826 878 2142 881
rect 2146 878 2238 881
rect 2242 878 2278 881
rect 2562 878 2574 881
rect 226 868 270 871
rect 658 868 750 871
rect 754 868 838 871
rect 1130 868 1214 871
rect 1290 868 1374 871
rect 1410 868 1470 871
rect 1474 868 1478 871
rect 1578 868 1614 871
rect 1754 868 1833 871
rect 1890 868 1894 871
rect 1906 868 1950 871
rect 1974 868 1993 871
rect 2010 868 2046 871
rect 2050 868 2126 871
rect 2234 868 2558 871
rect 50 858 118 861
rect 170 858 174 861
rect 346 858 398 861
rect 454 861 457 868
rect 454 858 518 861
rect 550 861 553 868
rect 1030 862 1033 868
rect 550 858 574 861
rect 578 858 654 861
rect 670 858 726 861
rect 762 858 766 861
rect 1202 858 1214 861
rect 1246 861 1249 868
rect 1242 858 1249 861
rect 1362 858 1382 861
rect 1386 858 1390 861
rect 1694 861 1697 868
rect 1830 862 1833 868
rect 1974 862 1977 868
rect 1990 862 1993 868
rect 2190 862 2193 868
rect 1442 858 1726 861
rect 1882 858 1926 861
rect 2066 858 2134 861
rect 2162 858 2166 861
rect 2574 861 2577 868
rect 2574 858 2606 861
rect 262 851 265 858
rect 218 848 265 851
rect 438 851 441 858
rect 670 852 673 858
rect 438 848 478 851
rect 706 848 742 851
rect 930 848 1062 851
rect 1122 848 1294 851
rect 1298 848 1606 851
rect 1610 848 1622 851
rect 2062 851 2065 858
rect 1826 848 2065 851
rect 2134 851 2137 858
rect 2134 848 2230 851
rect 2234 848 2286 851
rect 2418 848 2470 851
rect 2474 848 2534 851
rect 2538 848 2582 851
rect 394 838 422 841
rect 890 838 918 841
rect 1394 838 1422 841
rect 1450 838 1630 841
rect 1814 841 1817 848
rect 1814 838 1830 841
rect 1930 838 2118 841
rect 2134 838 2150 841
rect 254 832 257 838
rect 2134 832 2137 838
rect 770 828 790 831
rect 850 828 1478 831
rect 1594 828 1854 831
rect 2306 828 2342 831
rect 10 818 78 821
rect 846 821 849 828
rect 82 818 849 821
rect 1418 818 1638 821
rect 1658 818 1974 821
rect 1986 818 2214 821
rect 2226 818 2310 821
rect 250 808 254 811
rect 906 808 1086 811
rect 1106 808 1414 811
rect 1634 808 1822 811
rect 1858 808 2174 811
rect 2178 808 2238 811
rect 2258 808 2318 811
rect 2322 808 2350 811
rect 544 803 546 807
rect 550 803 553 807
rect 558 803 560 807
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1574 803 1576 807
rect 578 798 638 801
rect 770 798 1270 801
rect 1650 798 1710 801
rect 1842 798 2262 801
rect 2426 798 2430 801
rect 242 788 1102 791
rect 1106 788 1326 791
rect 1330 788 1478 791
rect 1642 788 1822 791
rect 1954 788 2249 791
rect 2246 782 2249 788
rect 2382 782 2385 788
rect 642 778 806 781
rect 946 778 1462 781
rect 1466 778 1502 781
rect 1506 778 1598 781
rect 1610 778 1718 781
rect 1722 778 1958 781
rect 1962 778 2070 781
rect 2102 778 2230 781
rect 2250 778 2326 781
rect 2102 772 2105 778
rect 282 768 406 771
rect 410 768 470 771
rect 602 768 694 771
rect 698 768 718 771
rect 938 768 1254 771
rect 1290 768 1566 771
rect 1582 768 1630 771
rect 1642 768 1966 771
rect 2274 768 2302 771
rect 2318 768 2326 771
rect 2330 768 2382 771
rect 1582 762 1585 768
rect 1966 762 1969 768
rect 130 758 142 761
rect 146 758 182 761
rect 322 758 406 761
rect 410 758 734 761
rect 738 758 894 761
rect 922 758 942 761
rect 962 758 1278 761
rect 1394 758 1414 761
rect 1554 758 1582 761
rect 1634 758 1654 761
rect 1706 758 1926 761
rect 1970 758 2078 761
rect 2226 758 2230 761
rect 2266 758 2310 761
rect 2314 758 2318 761
rect 2490 758 2494 761
rect 2506 758 2542 761
rect 1414 752 1417 758
rect 1422 752 1425 758
rect 50 748 118 751
rect 130 748 254 751
rect 258 748 294 751
rect 450 748 518 751
rect 778 748 846 751
rect 882 748 1014 751
rect 1066 748 1070 751
rect 1126 748 1142 751
rect 1346 748 1398 751
rect 1522 748 1766 751
rect 1770 748 1870 751
rect 1874 748 1902 751
rect 1978 748 1982 751
rect 2098 748 2102 751
rect 2170 748 2206 751
rect 2242 748 2262 751
rect 2330 748 2438 751
rect 2458 748 2494 751
rect 106 738 390 741
rect 662 741 665 748
rect 662 738 814 741
rect 818 738 1014 741
rect 1118 741 1121 748
rect 1018 738 1121 741
rect 1126 742 1129 748
rect 1250 738 1630 741
rect 1642 738 1686 741
rect 1778 738 1862 741
rect 1890 738 1894 741
rect 1986 738 2006 741
rect 2018 738 2070 741
rect 2074 738 2390 741
rect 2394 738 2478 741
rect 194 728 289 731
rect 642 728 710 731
rect 770 728 886 731
rect 890 728 894 731
rect 1010 728 1094 731
rect 1106 728 1190 731
rect 1274 728 1334 731
rect 1338 728 1422 731
rect 1666 728 1670 731
rect 1850 728 1998 731
rect 2114 728 2126 731
rect 2458 728 2462 731
rect 286 722 289 728
rect 1830 722 1833 728
rect 2438 722 2441 728
rect 258 718 270 721
rect 474 718 566 721
rect 594 718 646 721
rect 650 718 678 721
rect 1050 718 1086 721
rect 1090 718 1302 721
rect 1618 718 1702 721
rect 1874 718 1910 721
rect 1914 718 2230 721
rect 2234 718 2294 721
rect 2474 718 2494 721
rect 2570 718 2574 721
rect 186 708 334 711
rect 346 708 702 711
rect 910 708 950 711
rect 1602 708 1654 711
rect 1666 708 1734 711
rect 1802 708 1886 711
rect 2162 708 2238 711
rect 2298 708 2318 711
rect 274 698 446 701
rect 910 701 913 708
rect 1056 703 1058 707
rect 1062 703 1065 707
rect 1070 703 1072 707
rect 2080 703 2082 707
rect 2086 703 2089 707
rect 2094 703 2096 707
rect 538 698 913 701
rect 922 698 950 701
rect 1090 698 1134 701
rect 1138 698 1342 701
rect 1426 698 1742 701
rect 1746 698 1894 701
rect 1978 698 2062 701
rect 2066 698 2070 701
rect 202 688 254 691
rect 298 688 470 691
rect 546 688 590 691
rect 898 688 950 691
rect 954 688 1070 691
rect 1282 688 1294 691
rect 1322 688 1406 691
rect 1562 688 1606 691
rect 1610 688 1646 691
rect 1666 688 1694 691
rect 1722 688 1726 691
rect 1730 688 1806 691
rect 2034 688 2198 691
rect 2282 688 2422 691
rect 2434 688 2550 691
rect 242 678 294 681
rect 362 678 374 681
rect 402 678 406 681
rect 522 678 766 681
rect 834 678 918 681
rect 986 678 1273 681
rect 1290 678 1294 681
rect 1514 678 1582 681
rect 1682 678 1974 681
rect 2058 678 2174 681
rect 2250 678 2382 681
rect 2410 678 2454 681
rect 2514 678 2526 681
rect 1270 672 1273 678
rect 1478 672 1481 678
rect 10 668 81 671
rect 138 668 238 671
rect 266 668 278 671
rect 698 668 774 671
rect 962 668 1062 671
rect 1066 668 1118 671
rect 1210 668 1214 671
rect 1226 668 1254 671
rect 1274 668 1318 671
rect 1506 668 1518 671
rect 1622 671 1625 678
rect 1646 671 1649 678
rect 1622 668 1649 671
rect 1678 672 1681 678
rect 2478 672 2481 678
rect 1778 668 1838 671
rect 2002 668 2118 671
rect 2130 668 2254 671
rect 2298 668 2478 671
rect 2490 668 2558 671
rect 78 662 81 668
rect 350 662 353 668
rect 502 662 505 668
rect 646 662 649 668
rect 654 662 657 668
rect 662 662 665 668
rect 90 658 286 661
rect 394 658 486 661
rect 562 658 566 661
rect 578 658 582 661
rect 706 658 710 661
rect 738 658 742 661
rect 894 661 897 668
rect 894 658 902 661
rect 906 658 918 661
rect 938 658 950 661
rect 970 658 1094 661
rect 1142 661 1145 668
rect 1334 662 1337 668
rect 1366 662 1369 668
rect 1374 662 1377 668
rect 1494 662 1497 668
rect 1694 662 1697 668
rect 1702 662 1705 668
rect 1998 662 2001 668
rect 2486 662 2489 668
rect 1114 658 1145 661
rect 1178 658 1246 661
rect 1258 658 1262 661
rect 1266 658 1302 661
rect 1386 658 1462 661
rect 1466 658 1486 661
rect 1498 658 1582 661
rect 1666 658 1678 661
rect 1826 658 1838 661
rect 1962 658 1966 661
rect 2026 658 2030 661
rect 2034 658 2142 661
rect 2322 658 2425 661
rect 2522 658 2542 661
rect 2190 652 2193 658
rect 2422 652 2425 658
rect 162 648 246 651
rect 250 648 358 651
rect 546 648 790 651
rect 906 648 910 651
rect 970 648 1030 651
rect 1042 648 1182 651
rect 1186 648 1358 651
rect 1418 648 1526 651
rect 2066 648 2086 651
rect 2502 651 2505 658
rect 2442 648 2505 651
rect 2542 648 2606 651
rect 1670 642 1673 648
rect 2542 642 2545 648
rect 178 638 334 641
rect 362 638 422 641
rect 434 638 454 641
rect 482 638 486 641
rect 538 638 718 641
rect 922 638 1006 641
rect 1082 638 1126 641
rect 1130 638 1214 641
rect 1250 638 1265 641
rect 1378 638 1558 641
rect 2110 638 2126 641
rect 326 628 334 631
rect 338 628 510 631
rect 522 628 622 631
rect 782 631 785 638
rect 1262 632 1265 638
rect 2110 632 2113 638
rect 782 628 1230 631
rect 1554 628 1718 631
rect 1914 628 2054 631
rect 2122 628 2270 631
rect 2466 628 2558 631
rect 458 618 798 621
rect 802 618 894 621
rect 1042 618 1374 621
rect 1550 618 1614 621
rect 1802 618 2166 621
rect 2170 618 2326 621
rect 2498 618 2510 621
rect 450 608 534 611
rect 1034 608 1310 611
rect 1550 611 1553 618
rect 1370 608 1553 611
rect 1594 608 1966 611
rect 1970 608 2110 611
rect 544 603 546 607
rect 550 603 553 607
rect 558 603 560 607
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1574 603 1576 607
rect 1394 598 1398 601
rect 1586 598 2358 601
rect 258 588 942 591
rect 1434 588 1590 591
rect 1642 588 1902 591
rect 1906 588 1934 591
rect 1962 588 2254 591
rect 2258 588 2430 591
rect 306 578 406 581
rect 410 578 414 581
rect 418 578 574 581
rect 690 578 694 581
rect 842 578 886 581
rect 890 578 1046 581
rect 1290 578 1398 581
rect 1762 578 2062 581
rect 2554 578 2606 581
rect 734 572 737 578
rect 274 568 414 571
rect 418 568 430 571
rect 698 568 734 571
rect 754 568 870 571
rect 874 568 902 571
rect 1026 568 1134 571
rect 1346 568 1390 571
rect 1394 568 1438 571
rect 1530 568 1606 571
rect 1610 568 1630 571
rect 1698 568 1742 571
rect 1746 568 1870 571
rect 2018 568 2270 571
rect 2426 568 2534 571
rect 2594 568 2630 571
rect 678 562 681 568
rect 1302 562 1305 568
rect 170 558 294 561
rect 514 558 598 561
rect 686 558 942 561
rect 1102 558 1118 561
rect 1306 558 1326 561
rect 1578 558 1646 561
rect 1770 558 1790 561
rect 1990 561 1993 568
rect 1990 558 2022 561
rect 2098 558 2182 561
rect 2298 558 2302 561
rect 2306 558 2342 561
rect 2370 558 2406 561
rect 2594 558 2598 561
rect 150 551 153 558
rect 150 548 198 551
rect 242 548 310 551
rect 422 551 425 558
rect 686 551 689 558
rect 942 552 945 558
rect 1102 552 1105 558
rect 422 548 689 551
rect 802 548 846 551
rect 890 548 894 551
rect 1022 548 1086 551
rect 1114 548 1126 551
rect 1130 548 1150 551
rect 1242 548 1310 551
rect 1382 551 1385 558
rect 1766 552 1769 558
rect 1382 548 1422 551
rect 1530 548 1622 551
rect 1714 548 1750 551
rect 1778 548 1846 551
rect 1946 548 2006 551
rect 2106 548 2142 551
rect 70 541 73 548
rect 206 541 209 548
rect 1022 542 1025 548
rect 70 538 209 541
rect 354 538 430 541
rect 474 538 582 541
rect 586 538 630 541
rect 674 538 718 541
rect 866 538 926 541
rect 1174 541 1177 548
rect 2234 548 2265 551
rect 2314 548 2478 551
rect 2482 548 2510 551
rect 2554 548 2574 551
rect 2262 542 2265 548
rect 1154 538 1177 541
rect 1362 538 1694 541
rect 1706 538 1798 541
rect 1946 538 2246 541
rect 2290 538 2318 541
rect 2458 538 2486 541
rect 2570 538 2598 541
rect 106 528 158 531
rect 562 528 622 531
rect 626 528 638 531
rect 1042 528 1126 531
rect 1426 528 1518 531
rect 1738 528 1774 531
rect 1954 528 2118 531
rect 2122 528 2334 531
rect 2338 528 2390 531
rect 154 518 246 521
rect 298 518 350 521
rect 410 518 694 521
rect 914 518 1462 521
rect 1474 518 1510 521
rect 1754 518 1798 521
rect 1962 518 1974 521
rect 2002 518 2022 521
rect 2202 518 2310 521
rect 2354 518 2462 521
rect 578 508 598 511
rect 602 508 686 511
rect 1098 508 1166 511
rect 1210 508 1278 511
rect 1434 508 1446 511
rect 1690 508 1710 511
rect 2418 508 2526 511
rect 2530 508 2590 511
rect 1056 503 1058 507
rect 1062 503 1065 507
rect 1070 503 1072 507
rect 2080 503 2082 507
rect 2086 503 2089 507
rect 2094 503 2096 507
rect 986 498 1038 501
rect 1258 498 1294 501
rect 178 488 182 491
rect 186 488 262 491
rect 338 488 358 491
rect 434 488 518 491
rect 634 488 670 491
rect 690 488 710 491
rect 718 491 721 498
rect 718 488 862 491
rect 1322 488 1326 491
rect 1402 488 1462 491
rect 1522 488 1582 491
rect 2066 488 2174 491
rect 2242 488 2350 491
rect 2354 488 2385 491
rect 2426 488 2462 491
rect 2466 488 2478 491
rect 390 481 393 488
rect 146 478 526 481
rect 802 478 878 481
rect 990 481 993 488
rect 2382 482 2385 488
rect 906 478 993 481
rect 1298 478 1318 481
rect 1322 478 1390 481
rect 1394 478 1550 481
rect 1674 478 1854 481
rect 2002 478 2118 481
rect 2450 478 2526 481
rect 266 468 318 471
rect 490 468 534 471
rect 730 468 822 471
rect 826 468 838 471
rect 842 468 910 471
rect 914 468 990 471
rect 994 468 1006 471
rect 1286 471 1289 478
rect 1286 468 1310 471
rect 1314 468 1438 471
rect 1746 468 1830 471
rect 1854 471 1857 478
rect 1854 468 1990 471
rect 2018 468 2134 471
rect 2330 468 2438 471
rect 166 462 169 468
rect 50 458 118 461
rect 226 459 278 461
rect 222 458 278 459
rect 322 458 326 461
rect 362 458 534 461
rect 574 461 577 468
rect 538 458 582 461
rect 834 458 846 461
rect 986 458 1030 461
rect 1174 461 1177 468
rect 1174 458 1230 461
rect 1290 458 1438 461
rect 1558 461 1561 468
rect 2310 462 2313 468
rect 1538 458 1590 461
rect 1770 458 2070 461
rect 2074 458 2118 461
rect 2202 458 2217 461
rect 2314 458 2334 461
rect 2526 461 2529 468
rect 2514 458 2529 461
rect 2538 458 2598 461
rect 1438 452 1441 458
rect 2214 452 2217 458
rect 314 448 582 451
rect 618 448 622 451
rect 786 448 825 451
rect 858 448 1118 451
rect 1242 448 1262 451
rect 1282 448 1350 451
rect 1386 448 1430 451
rect 1558 448 1646 451
rect 1730 448 1758 451
rect 1762 448 1822 451
rect 1858 448 1878 451
rect 2018 448 2166 451
rect 2378 448 2542 451
rect 2546 448 2606 451
rect 822 442 825 448
rect 1558 442 1561 448
rect 930 438 1102 441
rect 1106 438 1118 441
rect 1250 438 1318 441
rect 1322 438 1334 441
rect 1338 438 1430 441
rect 1970 438 2046 441
rect 2186 438 2262 441
rect 2306 438 2414 441
rect 2418 438 2430 441
rect 2610 438 2646 441
rect 930 428 1086 431
rect 1330 428 1401 431
rect 1434 428 1566 431
rect 1570 428 1598 431
rect 1602 428 1654 431
rect 1658 428 1718 431
rect 2290 428 2502 431
rect 1398 422 1401 428
rect 386 418 958 421
rect 1234 418 1262 421
rect 1362 418 1374 421
rect 1458 418 1806 421
rect 1826 418 2046 421
rect 2258 418 2438 421
rect 2442 418 2478 421
rect 842 408 1038 411
rect 2042 408 2126 411
rect 544 403 546 407
rect 550 403 553 407
rect 558 403 560 407
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1574 403 1576 407
rect 866 398 1158 401
rect 1450 398 1534 401
rect 1706 398 2062 401
rect 2178 398 2470 401
rect 2474 398 2494 401
rect 2498 398 2598 401
rect 10 388 134 391
rect 138 388 150 391
rect 662 388 1222 391
rect 1234 388 1454 391
rect 1514 388 1518 391
rect 1546 388 1566 391
rect 1682 388 1726 391
rect 1730 388 2118 391
rect 662 382 665 388
rect 698 378 718 381
rect 722 378 846 381
rect 850 378 886 381
rect 898 378 1190 381
rect 1442 378 1542 381
rect 1562 378 1678 381
rect 1690 378 1702 381
rect 1874 378 2150 381
rect 18 368 38 371
rect 42 368 126 371
rect 738 368 822 371
rect 826 368 870 371
rect 1106 368 1110 371
rect 1186 368 1910 371
rect 2350 368 2358 371
rect 2362 368 2414 371
rect 2262 362 2265 368
rect 2326 362 2329 368
rect 282 358 294 361
rect 298 358 390 361
rect 626 358 638 361
rect 642 358 670 361
rect 802 358 806 361
rect 962 358 1046 361
rect 1050 358 1174 361
rect 1422 358 1742 361
rect 1746 358 1766 361
rect 1810 358 1838 361
rect 1842 358 1878 361
rect 2050 358 2070 361
rect 2330 358 2350 361
rect 118 351 121 358
rect 118 348 222 351
rect 346 348 358 351
rect 378 348 406 351
rect 610 348 614 351
rect 634 348 638 351
rect 766 351 769 358
rect 722 348 769 351
rect 798 351 801 358
rect 1422 352 1425 358
rect 798 348 894 351
rect 1018 348 1022 351
rect 1066 348 1254 351
rect 1402 348 1406 351
rect 1410 348 1422 351
rect 1666 348 1670 351
rect 1826 348 1886 351
rect 1898 348 1966 351
rect 2030 351 2033 358
rect 2198 351 2201 358
rect 2026 348 2201 351
rect 2314 348 2366 351
rect 2498 348 2566 351
rect 2602 348 2630 351
rect 178 338 230 341
rect 234 338 382 341
rect 618 338 638 341
rect 698 338 814 341
rect 842 338 886 341
rect 922 338 926 341
rect 978 338 1046 341
rect 1178 338 1238 341
rect 1242 338 1334 341
rect 1446 341 1449 348
rect 1338 338 1449 341
rect 1546 338 1750 341
rect 1778 338 1886 341
rect 1898 338 1902 341
rect 1954 338 2014 341
rect 2074 338 2222 341
rect 2226 338 2254 341
rect 50 328 70 331
rect 74 328 94 331
rect 114 328 126 331
rect 194 328 222 331
rect 274 328 326 331
rect 602 328 614 331
rect 1034 328 1342 331
rect 1538 328 1606 331
rect 1758 331 1761 338
rect 1618 328 1761 331
rect 1874 328 1934 331
rect 1938 328 1990 331
rect 2026 328 2070 331
rect 2106 328 2158 331
rect 2194 328 2550 331
rect 258 318 310 321
rect 314 318 342 321
rect 450 318 534 321
rect 586 318 646 321
rect 706 318 1246 321
rect 1594 318 1790 321
rect 2146 318 2326 321
rect 266 308 630 311
rect 922 308 950 311
rect 1306 308 1702 311
rect 1850 308 1910 311
rect 1914 308 2014 311
rect 2018 308 2038 311
rect 2362 308 2462 311
rect 2466 308 2478 311
rect 2482 308 2614 311
rect 1056 303 1058 307
rect 1062 303 1065 307
rect 1070 303 1072 307
rect 2080 303 2082 307
rect 2086 303 2089 307
rect 2094 303 2096 307
rect 2190 302 2193 308
rect 362 298 390 301
rect 418 298 454 301
rect 1418 298 1446 301
rect 2226 298 2262 301
rect 2378 298 2486 301
rect 210 288 278 291
rect 358 291 361 298
rect 322 288 361 291
rect 378 288 422 291
rect 442 288 462 291
rect 738 288 873 291
rect 978 288 1142 291
rect 1554 288 1638 291
rect 1642 288 1726 291
rect 1814 288 1822 291
rect 1826 288 1846 291
rect 1914 288 1950 291
rect 1962 288 2030 291
rect 2058 288 2102 291
rect 2210 288 2214 291
rect 2234 288 2238 291
rect 2274 288 2342 291
rect 2346 288 2430 291
rect 870 282 873 288
rect 330 278 478 281
rect 794 278 841 281
rect 858 278 862 281
rect 874 278 942 281
rect 1170 278 1566 281
rect 1610 278 2054 281
rect 2138 278 2398 281
rect 2538 278 2638 281
rect 294 271 297 278
rect 166 268 297 271
rect 486 271 489 278
rect 426 268 542 271
rect 618 268 662 271
rect 722 268 830 271
rect 838 271 841 278
rect 838 268 894 271
rect 1178 268 1182 271
rect 1682 268 2006 271
rect 2018 268 2030 271
rect 2082 268 2182 271
rect 2386 268 2390 271
rect 62 261 65 268
rect 166 262 169 268
rect 62 258 102 261
rect 130 258 166 261
rect 218 258 246 261
rect 390 261 393 268
rect 354 258 393 261
rect 482 258 606 261
rect 738 258 937 261
rect 1050 258 1134 261
rect 1170 258 1193 261
rect 1274 258 1342 261
rect 1422 261 1425 268
rect 1378 258 1425 261
rect 1494 261 1497 268
rect 1474 258 1518 261
rect 1522 258 1654 261
rect 1658 258 1686 261
rect 1754 258 2038 261
rect 2074 258 2166 261
rect 2398 261 2401 268
rect 2398 258 2446 261
rect 2506 258 2510 261
rect 934 252 937 258
rect 1190 252 1193 258
rect 482 248 502 251
rect 530 248 617 251
rect 682 248 694 251
rect 842 248 846 251
rect 1026 248 1038 251
rect 1514 248 1582 251
rect 1690 248 2438 251
rect 2442 248 2470 251
rect 614 242 617 248
rect 1050 238 1094 241
rect 1098 238 1238 241
rect 1250 238 1390 241
rect 1394 238 1590 241
rect 1662 241 1665 248
rect 1662 238 1758 241
rect 1970 238 2566 241
rect 258 228 422 231
rect 426 228 502 231
rect 890 228 1750 231
rect 674 218 750 221
rect 1722 218 1814 221
rect 1834 218 2222 221
rect 642 208 1062 211
rect 1090 208 1198 211
rect 1938 208 2278 211
rect 544 203 546 207
rect 550 203 553 207
rect 558 203 560 207
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1574 203 1576 207
rect 1018 198 1086 201
rect 1090 198 1142 201
rect 1658 198 2374 201
rect 2550 192 2553 198
rect 18 188 78 191
rect 82 188 182 191
rect 682 188 806 191
rect 834 188 862 191
rect 970 188 974 191
rect 1066 188 1302 191
rect 1866 188 1958 191
rect 2542 182 2545 188
rect 418 178 526 181
rect 530 178 574 181
rect 578 178 1006 181
rect 1186 178 1326 181
rect 1474 178 1478 181
rect 1594 178 1598 181
rect 2506 178 2518 181
rect 194 168 198 171
rect 634 168 734 171
rect 738 168 742 171
rect 858 168 878 171
rect 882 168 934 171
rect 1010 168 1830 171
rect 2090 168 2118 171
rect 2274 168 2326 171
rect 90 158 110 161
rect 146 158 174 161
rect 178 158 622 161
rect 910 158 918 161
rect 922 158 926 161
rect 938 158 942 161
rect 1234 158 1254 161
rect 1258 158 1654 161
rect 1754 158 1766 161
rect 2110 158 2118 161
rect 2122 158 2182 161
rect 2518 161 2521 168
rect 2518 158 2526 161
rect 118 152 121 158
rect 734 152 737 158
rect 70 148 102 151
rect 122 148 582 151
rect 586 148 614 151
rect 618 148 622 151
rect 838 151 841 158
rect 1838 152 1841 158
rect 838 148 958 151
rect 994 148 998 151
rect 1114 148 1286 151
rect 1346 148 1486 151
rect 1490 148 1526 151
rect 1530 148 1606 151
rect 1610 148 1710 151
rect 1714 148 1742 151
rect 70 142 73 148
rect 186 138 190 141
rect 194 138 198 141
rect 242 138 334 141
rect 354 138 374 141
rect 594 138 606 141
rect 614 138 662 141
rect 954 138 1086 141
rect 1090 138 1118 141
rect 1410 138 1446 141
rect 1450 138 1489 141
rect 1570 138 1646 141
rect 1650 138 1662 141
rect 1870 141 1873 158
rect 1890 148 1966 151
rect 1970 148 2102 151
rect 2106 148 2134 151
rect 2138 148 2206 151
rect 2286 151 2289 158
rect 2210 148 2289 151
rect 2314 148 2374 151
rect 2514 148 2598 151
rect 1770 138 1873 141
rect 2002 138 2110 141
rect 2250 138 2478 141
rect 2482 138 2486 141
rect 70 128 126 131
rect 398 131 401 138
rect 138 128 401 131
rect 614 132 617 138
rect 1486 132 1489 138
rect 1514 128 1614 131
rect 1794 128 1942 131
rect 70 122 73 128
rect 306 118 374 121
rect 506 118 974 121
rect 986 118 1078 121
rect 1138 118 1230 121
rect 1802 118 1926 121
rect 2066 118 2190 121
rect 658 108 934 111
rect 1056 103 1058 107
rect 1062 103 1065 107
rect 1070 103 1072 107
rect 2080 103 2082 107
rect 2086 103 2089 107
rect 2094 103 2096 107
rect 770 98 814 101
rect 818 98 910 101
rect 1226 98 1294 101
rect 1298 98 1350 101
rect 2210 98 2254 101
rect 2258 98 2294 101
rect 2306 98 2374 101
rect 2378 98 2478 101
rect 210 88 294 91
rect 386 88 558 91
rect 562 88 662 91
rect 714 88 798 91
rect 802 88 846 91
rect 930 88 958 91
rect 962 88 1046 91
rect 1178 88 1201 91
rect 1666 88 1686 91
rect 1762 88 1790 91
rect 1898 88 2006 91
rect 2050 88 2254 91
rect 2258 88 2422 91
rect 2426 88 2438 91
rect 2442 88 2462 91
rect 1198 82 1201 88
rect 10 78 422 81
rect 650 78 726 81
rect 730 78 966 81
rect 970 78 974 81
rect 1282 78 1318 81
rect 1322 78 1430 81
rect 1434 78 1510 81
rect 1514 78 1574 81
rect 1618 78 1686 81
rect 1714 78 1774 81
rect 1794 78 1910 81
rect 2114 78 2182 81
rect 2186 78 2198 81
rect 6 72 9 78
rect 82 68 86 71
rect 258 68 318 71
rect 354 68 382 71
rect 410 68 494 71
rect 498 68 558 71
rect 690 68 742 71
rect 882 68 934 71
rect 1018 68 1094 71
rect 1138 68 1718 71
rect 1746 68 1766 71
rect 1910 71 1913 78
rect 2390 72 2393 78
rect 1910 68 2062 71
rect 326 62 329 68
rect 1134 62 1137 68
rect 314 58 326 61
rect 330 58 926 61
rect 930 58 942 61
rect 946 58 1022 61
rect 1050 58 1118 61
rect 1178 58 1246 61
rect 1314 58 1342 61
rect 1554 58 1734 61
rect 1762 58 1766 61
rect 1810 58 1878 61
rect 2150 61 2153 68
rect 2066 58 2153 61
rect 2270 61 2273 68
rect 2270 58 2342 61
rect 2566 61 2569 68
rect 2522 58 2569 61
rect 2598 61 2601 68
rect 2598 58 2630 61
rect 94 51 97 58
rect 94 48 118 51
rect 282 48 350 51
rect 626 48 1302 51
rect 1330 48 1390 51
rect 2146 48 2174 51
rect 2178 48 2502 51
rect 626 38 1150 41
rect 1154 38 1174 41
rect 514 8 526 11
rect 544 3 546 7
rect 550 3 553 7
rect 558 3 560 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1574 3 1576 7
<< m4contact >>
rect 546 2403 550 2407
rect 554 2403 557 2407
rect 557 2403 558 2407
rect 1562 2403 1566 2407
rect 1570 2403 1573 2407
rect 1573 2403 1574 2407
rect 1534 2398 1538 2402
rect 326 2358 330 2362
rect 6 2338 10 2342
rect 2230 2338 2234 2342
rect 1710 2318 1714 2322
rect 1058 2303 1062 2307
rect 1066 2303 1069 2307
rect 1069 2303 1070 2307
rect 2082 2303 2086 2307
rect 2090 2303 2093 2307
rect 2093 2303 2094 2307
rect 1294 2298 1298 2302
rect 1414 2268 1418 2272
rect 1734 2268 1738 2272
rect 326 2258 330 2262
rect 518 2258 522 2262
rect 1254 2258 1258 2262
rect 1318 2258 1322 2262
rect 2470 2258 2474 2262
rect 1174 2248 1178 2252
rect 1350 2248 1354 2252
rect 2342 2248 2346 2252
rect 2462 2248 2466 2252
rect 1358 2238 1362 2242
rect 2374 2228 2378 2232
rect 1214 2218 1218 2222
rect 2118 2218 2122 2222
rect 2550 2218 2554 2222
rect 1110 2208 1114 2212
rect 1278 2208 1282 2212
rect 546 2203 550 2207
rect 554 2203 557 2207
rect 557 2203 558 2207
rect 1562 2203 1566 2207
rect 1570 2203 1573 2207
rect 1573 2203 1574 2207
rect 1118 2198 1122 2202
rect 1790 2168 1794 2172
rect 2526 2168 2530 2172
rect 1150 2158 1154 2162
rect 2262 2158 2266 2162
rect 638 2148 642 2152
rect 1350 2148 1354 2152
rect 1710 2138 1714 2142
rect 1822 2138 1826 2142
rect 1998 2138 2002 2142
rect 1302 2128 1306 2132
rect 310 2118 314 2122
rect 798 2118 802 2122
rect 1182 2118 1186 2122
rect 1702 2118 1706 2122
rect 2062 2118 2066 2122
rect 2278 2118 2282 2122
rect 518 2108 522 2112
rect 2590 2108 2594 2112
rect 1058 2103 1062 2107
rect 1066 2103 1069 2107
rect 1069 2103 1070 2107
rect 2082 2103 2086 2107
rect 2090 2103 2093 2107
rect 2093 2103 2094 2107
rect 358 2098 362 2102
rect 2278 2098 2282 2102
rect 302 2088 306 2092
rect 2118 2088 2122 2092
rect 1414 2078 1418 2082
rect 1582 2078 1586 2082
rect 798 2068 802 2072
rect 2278 2068 2282 2072
rect 2294 2068 2298 2072
rect 318 2058 322 2062
rect 454 2058 458 2062
rect 782 2058 786 2062
rect 1174 2058 1178 2062
rect 2006 2058 2010 2062
rect 2118 2058 2122 2062
rect 334 2048 338 2052
rect 1166 2048 1170 2052
rect 1446 2048 1450 2052
rect 1630 2048 1634 2052
rect 2102 2048 2106 2052
rect 174 2028 178 2032
rect 1526 2028 1530 2032
rect 2310 2028 2314 2032
rect 526 2018 530 2022
rect 902 2018 906 2022
rect 1318 2018 1322 2022
rect 1542 2018 1546 2022
rect 2294 2018 2298 2022
rect 546 2003 550 2007
rect 554 2003 557 2007
rect 557 2003 558 2007
rect 1562 2003 1566 2007
rect 1570 2003 1573 2007
rect 1573 2003 1574 2007
rect 2062 1998 2066 2002
rect 886 1988 890 1992
rect 2558 1968 2562 1972
rect 190 1958 194 1962
rect 854 1958 858 1962
rect 1126 1958 1130 1962
rect 2134 1958 2138 1962
rect 2222 1958 2226 1962
rect 886 1948 890 1952
rect 1310 1948 1314 1952
rect 1550 1948 1554 1952
rect 1302 1938 1306 1942
rect 1662 1938 1666 1942
rect 2038 1938 2042 1942
rect 2158 1938 2162 1942
rect 438 1928 442 1932
rect 798 1928 802 1932
rect 1326 1928 1330 1932
rect 878 1918 882 1922
rect 846 1908 850 1912
rect 1590 1908 1594 1912
rect 2382 1908 2386 1912
rect 1058 1903 1062 1907
rect 1066 1903 1069 1907
rect 1069 1903 1070 1907
rect 2082 1903 2086 1907
rect 2090 1903 2093 1907
rect 2093 1903 2094 1907
rect 366 1898 370 1902
rect 1670 1898 1674 1902
rect 1734 1888 1738 1892
rect 2342 1888 2346 1892
rect 1102 1878 1106 1882
rect 1302 1878 1306 1882
rect 1798 1878 1802 1882
rect 230 1858 234 1862
rect 358 1858 362 1862
rect 414 1858 418 1862
rect 566 1858 570 1862
rect 686 1858 690 1862
rect 1670 1868 1674 1872
rect 1998 1868 2002 1872
rect 934 1858 938 1862
rect 1262 1858 1266 1862
rect 2342 1858 2346 1862
rect 2374 1858 2378 1862
rect 2470 1858 2474 1862
rect 326 1848 330 1852
rect 646 1848 650 1852
rect 1142 1848 1146 1852
rect 1398 1848 1402 1852
rect 1982 1848 1986 1852
rect 2038 1848 2042 1852
rect 422 1838 426 1842
rect 974 1828 978 1832
rect 1518 1828 1522 1832
rect 790 1818 794 1822
rect 1414 1818 1418 1822
rect 1422 1818 1426 1822
rect 2350 1818 2354 1822
rect 718 1808 722 1812
rect 1422 1808 1426 1812
rect 546 1803 550 1807
rect 554 1803 557 1807
rect 557 1803 558 1807
rect 1562 1803 1566 1807
rect 1570 1803 1573 1807
rect 1573 1803 1574 1807
rect 2462 1798 2466 1802
rect 566 1788 570 1792
rect 254 1778 258 1782
rect 1974 1778 1978 1782
rect 174 1768 178 1772
rect 310 1768 314 1772
rect 390 1768 394 1772
rect 1694 1768 1698 1772
rect 710 1758 714 1762
rect 1782 1758 1786 1762
rect 2262 1758 2266 1762
rect 454 1748 458 1752
rect 470 1748 474 1752
rect 518 1748 522 1752
rect 814 1748 818 1752
rect 846 1748 850 1752
rect 1110 1748 1114 1752
rect 1190 1748 1194 1752
rect 1998 1748 2002 1752
rect 2230 1748 2234 1752
rect 2246 1748 2250 1752
rect 2310 1748 2314 1752
rect 310 1738 314 1742
rect 390 1738 394 1742
rect 398 1738 402 1742
rect 526 1738 530 1742
rect 1478 1738 1482 1742
rect 1918 1738 1922 1742
rect 1990 1738 1994 1742
rect 2278 1738 2282 1742
rect 2486 1738 2490 1742
rect 358 1728 362 1732
rect 1030 1728 1034 1732
rect 1158 1728 1162 1732
rect 1366 1728 1370 1732
rect 1678 1728 1682 1732
rect 2238 1728 2242 1732
rect 2294 1728 2298 1732
rect 2446 1728 2450 1732
rect 486 1718 490 1722
rect 686 1708 690 1712
rect 1270 1708 1274 1712
rect 1734 1708 1738 1712
rect 1814 1708 1818 1712
rect 1058 1703 1062 1707
rect 1066 1703 1069 1707
rect 1069 1703 1070 1707
rect 2082 1703 2086 1707
rect 2090 1703 2093 1707
rect 2093 1703 2094 1707
rect 158 1698 162 1702
rect 1046 1698 1050 1702
rect 2022 1698 2026 1702
rect 2126 1698 2130 1702
rect 390 1688 394 1692
rect 1206 1688 1210 1692
rect 1214 1688 1218 1692
rect 1670 1688 1674 1692
rect 1934 1688 1938 1692
rect 2110 1688 2114 1692
rect 374 1678 378 1682
rect 1190 1678 1194 1682
rect 1598 1678 1602 1682
rect 518 1668 522 1672
rect 1270 1668 1274 1672
rect 1798 1668 1802 1672
rect 2014 1668 2018 1672
rect 2382 1668 2386 1672
rect 2582 1668 2586 1672
rect 766 1658 770 1662
rect 950 1658 954 1662
rect 998 1658 1002 1662
rect 1006 1658 1010 1662
rect 1470 1658 1474 1662
rect 1590 1658 1594 1662
rect 1638 1658 1642 1662
rect 1694 1658 1698 1662
rect 1718 1658 1722 1662
rect 1766 1658 1770 1662
rect 1870 1658 1874 1662
rect 1902 1658 1906 1662
rect 1942 1658 1946 1662
rect 1958 1658 1962 1662
rect 2174 1658 2178 1662
rect 2350 1658 2354 1662
rect 382 1648 386 1652
rect 846 1648 850 1652
rect 1222 1648 1226 1652
rect 1486 1648 1490 1652
rect 1510 1648 1514 1652
rect 1686 1648 1690 1652
rect 1750 1648 1754 1652
rect 2062 1648 2066 1652
rect 2462 1648 2466 1652
rect 1422 1638 1426 1642
rect 2574 1638 2578 1642
rect 1430 1628 1434 1632
rect 2166 1628 2170 1632
rect 1454 1618 1458 1622
rect 1902 1618 1906 1622
rect 1038 1608 1042 1612
rect 2246 1608 2250 1612
rect 546 1603 550 1607
rect 554 1603 557 1607
rect 557 1603 558 1607
rect 1562 1603 1566 1607
rect 1570 1603 1573 1607
rect 1573 1603 1574 1607
rect 1350 1598 1354 1602
rect 1766 1598 1770 1602
rect 2070 1598 2074 1602
rect 2110 1598 2114 1602
rect 2230 1588 2234 1592
rect 886 1578 890 1582
rect 1566 1568 1570 1572
rect 1702 1568 1706 1572
rect 1870 1568 1874 1572
rect 1966 1568 1970 1572
rect 1278 1558 1282 1562
rect 1494 1558 1498 1562
rect 438 1548 442 1552
rect 494 1548 498 1552
rect 790 1548 794 1552
rect 854 1548 858 1552
rect 894 1548 898 1552
rect 1358 1548 1362 1552
rect 1702 1548 1706 1552
rect 1758 1548 1762 1552
rect 2038 1548 2042 1552
rect 2542 1548 2546 1552
rect 2590 1548 2594 1552
rect 1094 1538 1098 1542
rect 1294 1538 1298 1542
rect 1422 1538 1426 1542
rect 1702 1538 1706 1542
rect 1766 1538 1770 1542
rect 2478 1538 2482 1542
rect 1414 1528 1418 1532
rect 1438 1528 1442 1532
rect 2070 1528 2074 1532
rect 2198 1528 2202 1532
rect 694 1518 698 1522
rect 918 1518 922 1522
rect 1430 1518 1434 1522
rect 1670 1518 1674 1522
rect 1318 1508 1322 1512
rect 1446 1508 1450 1512
rect 1454 1508 1458 1512
rect 1550 1508 1554 1512
rect 1622 1508 1626 1512
rect 1686 1508 1690 1512
rect 1058 1503 1062 1507
rect 1066 1503 1069 1507
rect 1069 1503 1070 1507
rect 2082 1503 2086 1507
rect 2090 1503 2093 1507
rect 2093 1503 2094 1507
rect 1670 1498 1674 1502
rect 846 1488 850 1492
rect 1126 1488 1130 1492
rect 1606 1488 1610 1492
rect 1038 1478 1042 1482
rect 1262 1478 1266 1482
rect 1286 1478 1290 1482
rect 1470 1478 1474 1482
rect 2598 1478 2602 1482
rect 470 1468 474 1472
rect 806 1468 810 1472
rect 1094 1468 1098 1472
rect 1750 1468 1754 1472
rect 2318 1468 2322 1472
rect 2382 1468 2386 1472
rect 190 1458 194 1462
rect 718 1458 722 1462
rect 750 1458 754 1462
rect 934 1458 938 1462
rect 974 1458 978 1462
rect 1014 1458 1018 1462
rect 1126 1458 1130 1462
rect 1822 1458 1826 1462
rect 2006 1458 2010 1462
rect 1006 1448 1010 1452
rect 1606 1448 1610 1452
rect 1878 1448 1882 1452
rect 2486 1448 2490 1452
rect 814 1438 818 1442
rect 1078 1438 1082 1442
rect 1214 1438 1218 1442
rect 1222 1438 1226 1442
rect 1430 1438 1434 1442
rect 1462 1438 1466 1442
rect 1630 1438 1634 1442
rect 526 1428 530 1432
rect 606 1428 610 1432
rect 710 1428 714 1432
rect 1206 1428 1210 1432
rect 2030 1428 2034 1432
rect 2262 1428 2266 1432
rect 2630 1428 2634 1432
rect 166 1418 170 1422
rect 726 1418 730 1422
rect 846 1418 850 1422
rect 998 1418 1002 1422
rect 1406 1418 1410 1422
rect 1486 1418 1490 1422
rect 1806 1418 1810 1422
rect 2078 1418 2082 1422
rect 1022 1408 1026 1412
rect 1462 1408 1466 1412
rect 1550 1408 1554 1412
rect 546 1403 550 1407
rect 554 1403 557 1407
rect 557 1403 558 1407
rect 1562 1403 1566 1407
rect 1570 1403 1573 1407
rect 1573 1403 1574 1407
rect 878 1398 882 1402
rect 1326 1398 1330 1402
rect 1398 1398 1402 1402
rect 1462 1398 1466 1402
rect 1806 1398 1810 1402
rect 1822 1398 1826 1402
rect 1582 1388 1586 1392
rect 334 1378 338 1382
rect 726 1378 730 1382
rect 1374 1378 1378 1382
rect 1790 1378 1794 1382
rect 286 1368 290 1372
rect 862 1368 866 1372
rect 902 1368 906 1372
rect 1054 1368 1058 1372
rect 1198 1368 1202 1372
rect 1782 1368 1786 1372
rect 2582 1368 2586 1372
rect 1102 1358 1106 1362
rect 1310 1358 1314 1362
rect 1526 1358 1530 1362
rect 1686 1358 1690 1362
rect 1806 1358 1810 1362
rect 1974 1358 1978 1362
rect 2166 1358 2170 1362
rect 2382 1358 2386 1362
rect 566 1348 570 1352
rect 630 1348 634 1352
rect 1014 1348 1018 1352
rect 1086 1348 1090 1352
rect 1118 1348 1122 1352
rect 1326 1348 1330 1352
rect 1998 1348 2002 1352
rect 2038 1348 2042 1352
rect 2158 1348 2162 1352
rect 2190 1348 2194 1352
rect 302 1338 306 1342
rect 534 1338 538 1342
rect 1390 1338 1394 1342
rect 1438 1338 1442 1342
rect 1454 1338 1458 1342
rect 1654 1338 1658 1342
rect 1670 1338 1674 1342
rect 1998 1338 2002 1342
rect 2110 1338 2114 1342
rect 2342 1338 2346 1342
rect 286 1328 290 1332
rect 718 1328 722 1332
rect 1038 1328 1042 1332
rect 1070 1328 1074 1332
rect 1158 1328 1162 1332
rect 1542 1328 1546 1332
rect 1614 1328 1618 1332
rect 1638 1328 1642 1332
rect 1646 1328 1650 1332
rect 1942 1328 1946 1332
rect 302 1318 306 1322
rect 318 1308 322 1312
rect 1078 1308 1082 1312
rect 1766 1308 1770 1312
rect 2070 1308 2074 1312
rect 1058 1303 1062 1307
rect 1066 1303 1069 1307
rect 1069 1303 1070 1307
rect 2082 1303 2086 1307
rect 2090 1303 2093 1307
rect 2093 1303 2094 1307
rect 382 1298 386 1302
rect 422 1298 426 1302
rect 702 1298 706 1302
rect 1030 1298 1034 1302
rect 2646 1298 2650 1302
rect 294 1288 298 1292
rect 310 1288 314 1292
rect 470 1288 474 1292
rect 1022 1288 1026 1292
rect 1718 1288 1722 1292
rect 2078 1288 2082 1292
rect 2102 1288 2106 1292
rect 2574 1288 2578 1292
rect 302 1278 306 1282
rect 446 1278 450 1282
rect 718 1278 722 1282
rect 2302 1278 2306 1282
rect 390 1268 394 1272
rect 1046 1268 1050 1272
rect 1118 1268 1122 1272
rect 1326 1268 1330 1272
rect 1598 1268 1602 1272
rect 1798 1268 1802 1272
rect 2398 1268 2402 1272
rect 310 1258 314 1262
rect 782 1258 786 1262
rect 854 1258 858 1262
rect 870 1258 874 1262
rect 894 1258 898 1262
rect 1174 1258 1178 1262
rect 1478 1258 1482 1262
rect 1678 1258 1682 1262
rect 1718 1258 1722 1262
rect 2054 1258 2058 1262
rect 2062 1258 2066 1262
rect 662 1248 666 1252
rect 1078 1248 1082 1252
rect 1086 1248 1090 1252
rect 1198 1248 1202 1252
rect 1446 1248 1450 1252
rect 1678 1248 1682 1252
rect 1966 1248 1970 1252
rect 478 1238 482 1242
rect 670 1238 674 1242
rect 1166 1238 1170 1242
rect 1430 1238 1434 1242
rect 1446 1238 1450 1242
rect 2318 1238 2322 1242
rect 2470 1238 2474 1242
rect 646 1228 650 1232
rect 734 1228 738 1232
rect 1102 1228 1106 1232
rect 1254 1228 1258 1232
rect 1662 1228 1666 1232
rect 2446 1228 2450 1232
rect 1350 1218 1354 1222
rect 886 1208 890 1212
rect 926 1208 930 1212
rect 2022 1208 2026 1212
rect 546 1203 550 1207
rect 554 1203 557 1207
rect 557 1203 558 1207
rect 1562 1203 1566 1207
rect 1570 1203 1573 1207
rect 1573 1203 1574 1207
rect 1934 1198 1938 1202
rect 2310 1198 2314 1202
rect 470 1188 474 1192
rect 1430 1188 1434 1192
rect 1478 1188 1482 1192
rect 2630 1188 2634 1192
rect 358 1178 362 1182
rect 502 1178 506 1182
rect 846 1178 850 1182
rect 1462 1178 1466 1182
rect 2374 1178 2378 1182
rect 2478 1178 2482 1182
rect 1246 1168 1250 1172
rect 1342 1168 1346 1172
rect 1918 1168 1922 1172
rect 2558 1168 2562 1172
rect 182 1158 186 1162
rect 470 1158 474 1162
rect 638 1158 642 1162
rect 878 1158 882 1162
rect 1398 1158 1402 1162
rect 1486 1158 1490 1162
rect 1590 1158 1594 1162
rect 2270 1158 2274 1162
rect 2326 1158 2330 1162
rect 534 1148 538 1152
rect 1302 1148 1306 1152
rect 1486 1148 1490 1152
rect 2030 1148 2034 1152
rect 2118 1148 2122 1152
rect 2582 1148 2586 1152
rect 6 1138 10 1142
rect 694 1138 698 1142
rect 1470 1138 1474 1142
rect 1926 1138 1930 1142
rect 318 1128 322 1132
rect 790 1128 794 1132
rect 1422 1128 1426 1132
rect 1438 1128 1442 1132
rect 230 1118 234 1122
rect 430 1118 434 1122
rect 918 1118 922 1122
rect 926 1118 930 1122
rect 2574 1118 2578 1122
rect 422 1108 426 1112
rect 518 1108 522 1112
rect 1246 1108 1250 1112
rect 1726 1108 1730 1112
rect 2038 1108 2042 1112
rect 2102 1108 2106 1112
rect 1058 1103 1062 1107
rect 1066 1103 1069 1107
rect 1069 1103 1070 1107
rect 2082 1103 2086 1107
rect 2090 1103 2093 1107
rect 2093 1103 2094 1107
rect 926 1098 930 1102
rect 1734 1098 1738 1102
rect 2126 1088 2130 1092
rect 254 1078 258 1082
rect 1134 1078 1138 1082
rect 1446 1078 1450 1082
rect 1606 1078 1610 1082
rect 1678 1078 1682 1082
rect 2094 1078 2098 1082
rect 2302 1078 2306 1082
rect 1366 1068 1370 1072
rect 1414 1068 1418 1072
rect 1550 1068 1554 1072
rect 1630 1068 1634 1072
rect 1654 1068 1658 1072
rect 2398 1068 2402 1072
rect 886 1058 890 1062
rect 1342 1058 1346 1062
rect 1534 1058 1538 1062
rect 1670 1058 1674 1062
rect 894 1048 898 1052
rect 2126 1048 2130 1052
rect 2606 1048 2610 1052
rect 1646 1038 1650 1042
rect 1822 1038 1826 1042
rect 1870 1038 1874 1042
rect 942 1028 946 1032
rect 1846 1028 1850 1032
rect 1998 1028 2002 1032
rect 2110 1028 2114 1032
rect 1038 1018 1042 1022
rect 2006 1018 2010 1022
rect 2062 1018 2066 1022
rect 1702 1008 1706 1012
rect 1998 1008 2002 1012
rect 546 1003 550 1007
rect 554 1003 557 1007
rect 557 1003 558 1007
rect 1562 1003 1566 1007
rect 1570 1003 1573 1007
rect 1573 1003 1574 1007
rect 118 998 122 1002
rect 470 998 474 1002
rect 806 998 810 1002
rect 190 988 194 992
rect 414 988 418 992
rect 678 988 682 992
rect 870 988 874 992
rect 1614 988 1618 992
rect 582 978 586 982
rect 710 978 714 982
rect 702 968 706 972
rect 1958 968 1962 972
rect 422 958 426 962
rect 1422 958 1426 962
rect 2486 958 2490 962
rect 158 948 162 952
rect 326 948 330 952
rect 918 948 922 952
rect 1286 948 1290 952
rect 1310 948 1314 952
rect 1814 948 1818 952
rect 710 938 714 942
rect 1422 938 1426 942
rect 1926 938 1930 942
rect 246 928 250 932
rect 390 928 394 932
rect 894 918 898 922
rect 1038 918 1042 922
rect 1846 918 1850 922
rect 1870 918 1874 922
rect 1878 918 1882 922
rect 2214 918 2218 922
rect 1838 908 1842 912
rect 1058 903 1062 907
rect 1066 903 1069 907
rect 1069 903 1070 907
rect 2082 903 2086 907
rect 2090 903 2093 907
rect 2093 903 2094 907
rect 1214 898 1218 902
rect 1886 898 1890 902
rect 1742 888 1746 892
rect 806 878 810 882
rect 2574 878 2578 882
rect 654 868 658 872
rect 750 868 754 872
rect 1406 868 1410 872
rect 1478 868 1482 872
rect 1894 868 1898 872
rect 2190 868 2194 872
rect 2230 868 2234 872
rect 174 858 178 862
rect 758 858 762 862
rect 1030 858 1034 862
rect 1238 858 1242 862
rect 1726 858 1730 862
rect 2166 858 2170 862
rect 1118 848 1122 852
rect 1606 848 1610 852
rect 1622 848 1626 852
rect 254 838 258 842
rect 1630 838 1634 842
rect 1478 828 1482 832
rect 6 818 10 822
rect 1638 818 1642 822
rect 1974 818 1978 822
rect 2214 818 2218 822
rect 254 808 258 812
rect 902 808 906 812
rect 1102 808 1106 812
rect 1822 808 1826 812
rect 2238 808 2242 812
rect 2318 808 2322 812
rect 2350 808 2354 812
rect 546 803 550 807
rect 554 803 557 807
rect 557 803 558 807
rect 1562 803 1566 807
rect 1570 803 1573 807
rect 1573 803 1574 807
rect 1646 798 1650 802
rect 2422 798 2426 802
rect 238 788 242 792
rect 1326 788 1330 792
rect 1606 778 1610 782
rect 2070 778 2074 782
rect 2230 778 2234 782
rect 2382 778 2386 782
rect 470 768 474 772
rect 1254 768 1258 772
rect 1566 768 1570 772
rect 182 758 186 762
rect 318 758 322 762
rect 1278 758 1282 762
rect 1550 758 1554 762
rect 1630 758 1634 762
rect 1966 758 1970 762
rect 2310 758 2314 762
rect 2486 758 2490 762
rect 126 748 130 752
rect 1070 748 1074 752
rect 1414 748 1418 752
rect 1422 748 1426 752
rect 1766 748 1770 752
rect 1982 748 1986 752
rect 2102 748 2106 752
rect 1126 738 1130 742
rect 1630 738 1634 742
rect 1894 738 1898 742
rect 2014 738 2018 742
rect 2390 738 2394 742
rect 886 728 890 732
rect 1094 728 1098 732
rect 1662 728 1666 732
rect 1830 728 1834 732
rect 2454 728 2458 732
rect 646 718 650 722
rect 1302 718 1306 722
rect 1702 718 1706 722
rect 2294 718 2298 722
rect 2438 718 2442 722
rect 702 708 706 712
rect 1654 708 1658 712
rect 1662 708 1666 712
rect 1798 708 1802 712
rect 2158 708 2162 712
rect 1058 703 1062 707
rect 1066 703 1069 707
rect 1069 703 1070 707
rect 2082 703 2086 707
rect 2090 703 2093 707
rect 2093 703 2094 707
rect 950 698 954 702
rect 1086 698 1090 702
rect 1342 698 1346 702
rect 2062 698 2066 702
rect 1278 688 1282 692
rect 1406 688 1410 692
rect 2422 688 2426 692
rect 406 678 410 682
rect 1294 678 1298 682
rect 2406 678 2410 682
rect 2478 678 2482 682
rect 238 668 242 672
rect 958 668 962 672
rect 1118 668 1122 672
rect 1206 668 1210 672
rect 1222 668 1226 672
rect 1334 668 1338 672
rect 1478 668 1482 672
rect 1502 668 1506 672
rect 1678 668 1682 672
rect 1694 668 1698 672
rect 350 658 354 662
rect 502 658 506 662
rect 558 658 562 662
rect 574 658 578 662
rect 646 658 650 662
rect 654 658 658 662
rect 662 658 666 662
rect 710 658 714 662
rect 742 658 746 662
rect 902 658 906 662
rect 918 658 922 662
rect 966 658 970 662
rect 1246 658 1250 662
rect 1254 658 1258 662
rect 1366 658 1370 662
rect 1374 658 1378 662
rect 1494 658 1498 662
rect 1662 658 1666 662
rect 1702 658 1706 662
rect 1966 658 1970 662
rect 1998 658 2002 662
rect 2030 658 2034 662
rect 2190 658 2194 662
rect 2318 658 2322 662
rect 2486 658 2490 662
rect 2518 658 2522 662
rect 910 648 914 652
rect 1038 648 1042 652
rect 1358 648 1362 652
rect 1670 648 1674 652
rect 2062 648 2066 652
rect 454 638 458 642
rect 486 638 490 642
rect 534 638 538 642
rect 1374 638 1378 642
rect 798 618 802 622
rect 894 618 898 622
rect 1374 618 1378 622
rect 2166 618 2170 622
rect 534 608 538 612
rect 2110 608 2114 612
rect 546 603 550 607
rect 554 603 557 607
rect 557 603 558 607
rect 1562 603 1566 607
rect 1570 603 1573 607
rect 1573 603 1574 607
rect 1398 598 1402 602
rect 1430 588 1434 592
rect 1638 588 1642 592
rect 1934 588 1938 592
rect 1958 588 1962 592
rect 686 578 690 582
rect 734 578 738 582
rect 430 568 434 572
rect 678 568 682 572
rect 1022 568 1026 572
rect 1526 568 1530 572
rect 1870 568 1874 572
rect 166 558 170 562
rect 1302 558 1306 562
rect 2294 558 2298 562
rect 2598 558 2602 562
rect 198 548 202 552
rect 894 548 898 552
rect 942 548 946 552
rect 1150 548 1154 552
rect 1422 548 1426 552
rect 1766 548 1770 552
rect 1942 548 1946 552
rect 470 538 474 542
rect 2310 548 2314 552
rect 1358 538 1362 542
rect 2454 538 2458 542
rect 694 518 698 522
rect 1462 518 1466 522
rect 1278 508 1282 512
rect 1058 503 1062 507
rect 1066 503 1069 507
rect 1069 503 1070 507
rect 2082 503 2086 507
rect 2090 503 2093 507
rect 2093 503 2094 507
rect 1294 498 1298 502
rect 1326 488 1330 492
rect 2422 488 2426 492
rect 1294 478 1298 482
rect 1318 478 1322 482
rect 166 468 170 472
rect 910 468 914 472
rect 1310 468 1314 472
rect 318 458 322 462
rect 582 458 586 462
rect 1438 458 1442 462
rect 1590 458 1594 462
rect 2118 458 2122 462
rect 2198 458 2202 462
rect 2310 458 2314 462
rect 622 448 626 452
rect 2542 448 2546 452
rect 2430 438 2434 442
rect 1086 428 1090 432
rect 958 418 962 422
rect 1806 418 1810 422
rect 1822 418 1826 422
rect 2438 418 2442 422
rect 1038 408 1042 412
rect 546 403 550 407
rect 554 403 557 407
rect 557 403 558 407
rect 1562 403 1566 407
rect 1570 403 1573 407
rect 1573 403 1574 407
rect 2062 398 2066 402
rect 2598 398 2602 402
rect 1222 388 1226 392
rect 846 378 850 382
rect 886 378 890 382
rect 894 378 898 382
rect 1678 378 1682 382
rect 1870 378 1874 382
rect 126 368 130 372
rect 1110 368 1114 372
rect 2262 368 2266 372
rect 390 358 394 362
rect 670 358 674 362
rect 806 358 810 362
rect 1806 358 1810 362
rect 2326 358 2330 362
rect 606 348 610 352
rect 638 348 642 352
rect 894 348 898 352
rect 1022 348 1026 352
rect 1062 348 1066 352
rect 1398 348 1402 352
rect 1662 348 1666 352
rect 1886 348 1890 352
rect 2022 348 2026 352
rect 230 338 234 342
rect 614 338 618 342
rect 918 338 922 342
rect 1750 338 1754 342
rect 1894 338 1898 342
rect 2014 338 2018 342
rect 1606 328 1610 332
rect 2550 328 2554 332
rect 1246 318 1250 322
rect 630 308 634 312
rect 2190 308 2194 312
rect 1058 303 1062 307
rect 1066 303 1069 307
rect 1069 303 1070 307
rect 2082 303 2086 307
rect 2090 303 2093 307
rect 2093 303 2094 307
rect 2374 298 2378 302
rect 1726 288 1730 292
rect 2214 288 2218 292
rect 854 278 858 282
rect 1606 278 1610 282
rect 542 268 546 272
rect 1174 268 1178 272
rect 1678 268 1682 272
rect 2014 268 2018 272
rect 2078 268 2082 272
rect 2382 268 2386 272
rect 734 258 738 262
rect 1470 258 1474 262
rect 1750 258 1754 262
rect 2070 258 2074 262
rect 838 248 842 252
rect 2470 248 2474 252
rect 1246 238 1250 242
rect 254 228 258 232
rect 886 228 890 232
rect 1934 208 1938 212
rect 546 203 550 207
rect 554 203 557 207
rect 557 203 558 207
rect 1562 203 1566 207
rect 1570 203 1573 207
rect 1573 203 1574 207
rect 2374 198 2378 202
rect 78 188 82 192
rect 974 188 978 192
rect 2542 188 2546 192
rect 2550 188 2554 192
rect 1478 178 1482 182
rect 1598 178 1602 182
rect 2518 178 2522 182
rect 198 168 202 172
rect 2326 168 2330 172
rect 926 158 930 162
rect 942 158 946 162
rect 2526 158 2530 162
rect 118 148 122 152
rect 622 148 626 152
rect 734 148 738 152
rect 998 148 1002 152
rect 1838 148 1842 152
rect 950 138 954 142
rect 2206 148 2210 152
rect 1790 128 1794 132
rect 1058 103 1062 107
rect 1066 103 1069 107
rect 1069 103 1070 107
rect 2082 103 2086 107
rect 2090 103 2093 107
rect 2093 103 2094 107
rect 846 88 850 92
rect 1790 88 1794 92
rect 966 78 970 82
rect 2198 78 2202 82
rect 6 68 10 72
rect 78 68 82 72
rect 326 68 330 72
rect 2390 68 2394 72
rect 1134 58 1138 62
rect 1766 58 1770 62
rect 118 48 122 52
rect 622 48 626 52
rect 546 3 550 7
rect 554 3 557 7
rect 557 3 558 7
rect 1562 3 1566 7
rect 1570 3 1573 7
rect 1573 3 1574 7
<< metal4 >>
rect 544 2403 546 2407
rect 550 2403 553 2407
rect 558 2403 560 2407
rect 1560 2403 1562 2407
rect 1566 2403 1569 2407
rect 1574 2403 1576 2407
rect 1526 2398 1534 2401
rect 6 1142 9 2338
rect 326 2262 329 2358
rect 1056 2303 1058 2307
rect 1062 2303 1065 2307
rect 1070 2303 1072 2307
rect 1258 2258 1262 2261
rect 302 2062 305 2088
rect 174 1772 177 2028
rect 6 822 9 1138
rect 6 72 9 818
rect 78 72 81 188
rect 118 152 121 998
rect 158 952 161 1698
rect 190 1462 193 1958
rect 194 1458 201 1461
rect 166 861 169 1418
rect 166 858 174 861
rect 126 372 129 748
rect 166 562 169 858
rect 182 762 185 1158
rect 166 472 169 558
rect 190 171 193 988
rect 198 552 201 1458
rect 230 1122 233 1858
rect 198 182 201 548
rect 230 342 233 1118
rect 254 1082 257 1778
rect 310 1772 313 2118
rect 282 1368 286 1371
rect 290 1328 294 1331
rect 302 1322 305 1338
rect 294 1282 297 1288
rect 302 1282 305 1318
rect 310 1292 313 1738
rect 318 1312 321 2058
rect 326 1852 329 2258
rect 518 2112 521 2258
rect 544 2203 546 2207
rect 550 2203 553 2207
rect 558 2203 560 2207
rect 334 1382 337 2048
rect 358 1862 361 2098
rect 450 2058 454 2061
rect 358 1732 361 1738
rect 366 1681 369 1898
rect 390 1742 393 1768
rect 398 1732 401 1738
rect 366 1678 374 1681
rect 390 1662 393 1688
rect 310 1262 313 1288
rect 318 1132 321 1308
rect 358 1182 361 1368
rect 382 1302 385 1648
rect 382 1271 385 1298
rect 382 1268 390 1271
rect 238 928 246 931
rect 238 792 241 928
rect 254 842 257 1078
rect 238 672 241 788
rect 254 232 257 808
rect 318 762 321 1128
rect 318 462 321 758
rect 190 168 198 171
rect 118 52 121 148
rect 326 72 329 948
rect 390 932 393 1268
rect 414 992 417 1858
rect 422 1842 425 1928
rect 422 1302 425 1838
rect 438 1552 441 1928
rect 518 1752 521 2108
rect 450 1748 454 1751
rect 470 1742 473 1748
rect 486 1722 489 1728
rect 518 1672 521 1748
rect 526 1742 529 2018
rect 544 2003 546 2007
rect 550 2003 553 2007
rect 558 2003 560 2007
rect 544 1803 546 1807
rect 550 1803 553 1807
rect 558 1803 560 1807
rect 566 1792 569 1858
rect 474 1468 478 1471
rect 450 1278 454 1281
rect 470 1192 473 1288
rect 478 1242 481 1248
rect 422 962 425 1108
rect 350 632 353 658
rect 390 362 393 928
rect 410 678 414 681
rect 430 572 433 1118
rect 470 1002 473 1158
rect 458 638 462 641
rect 470 542 473 768
rect 486 642 489 648
rect 494 632 497 1548
rect 502 662 505 1178
rect 518 1112 521 1668
rect 526 1432 529 1738
rect 544 1603 546 1607
rect 550 1603 553 1607
rect 558 1603 560 1607
rect 544 1403 546 1407
rect 550 1403 553 1407
rect 558 1403 560 1407
rect 566 1352 569 1788
rect 534 1152 537 1338
rect 544 1203 546 1207
rect 550 1203 553 1207
rect 558 1203 560 1207
rect 544 1003 546 1007
rect 550 1003 553 1007
rect 558 1003 560 1007
rect 544 803 546 807
rect 550 803 553 807
rect 558 803 560 807
rect 562 658 566 661
rect 574 652 577 658
rect 534 612 537 638
rect 544 603 546 607
rect 550 603 553 607
rect 558 603 560 607
rect 582 462 585 978
rect 544 403 546 407
rect 550 403 553 407
rect 558 403 560 407
rect 606 352 609 1428
rect 614 448 622 451
rect 602 348 606 351
rect 614 342 617 448
rect 630 351 633 1348
rect 638 1162 641 2148
rect 798 2072 801 2118
rect 1056 2103 1058 2107
rect 1062 2103 1065 2107
rect 1070 2103 1072 2107
rect 646 1232 649 1848
rect 686 1712 689 1858
rect 654 1251 657 1258
rect 654 1248 662 1251
rect 646 662 649 718
rect 654 662 657 868
rect 662 662 665 668
rect 670 362 673 1238
rect 694 1142 697 1518
rect 710 1432 713 1758
rect 718 1462 721 1808
rect 762 1658 766 1661
rect 678 572 681 988
rect 702 972 705 1298
rect 710 982 713 1428
rect 726 1382 729 1418
rect 718 1282 721 1328
rect 702 712 705 968
rect 710 942 713 978
rect 702 661 705 708
rect 702 658 710 661
rect 734 582 737 1228
rect 750 872 753 1458
rect 782 1262 785 2058
rect 802 1928 806 1931
rect 790 1552 793 1818
rect 846 1752 849 1908
rect 758 862 761 1258
rect 790 1132 793 1548
rect 802 1468 806 1471
rect 814 1442 817 1748
rect 846 1492 849 1648
rect 854 1552 857 1958
rect 886 1952 889 1988
rect 814 1262 817 1438
rect 846 1182 849 1418
rect 878 1402 881 1918
rect 854 1262 857 1268
rect 798 998 806 1001
rect 742 642 745 658
rect 798 622 801 998
rect 690 578 697 581
rect 694 522 697 578
rect 806 362 809 878
rect 846 382 849 1178
rect 630 348 638 351
rect 630 312 633 348
rect 630 282 633 308
rect 862 281 865 1368
rect 870 992 873 1258
rect 878 1162 881 1398
rect 886 1212 889 1578
rect 894 1262 897 1548
rect 902 1372 905 2018
rect 1056 1903 1058 1907
rect 1062 1903 1065 1907
rect 1070 1903 1072 1907
rect 918 1122 921 1518
rect 934 1462 937 1858
rect 954 1658 958 1661
rect 974 1462 977 1828
rect 1034 1728 1038 1731
rect 1056 1703 1058 1707
rect 1062 1703 1065 1707
rect 1070 1703 1072 1707
rect 1046 1672 1049 1698
rect 926 1458 934 1461
rect 978 1458 982 1461
rect 926 1212 929 1458
rect 998 1422 1001 1658
rect 1006 1452 1009 1658
rect 1038 1482 1041 1608
rect 1102 1541 1105 1878
rect 1110 1752 1113 2208
rect 1098 1538 1105 1541
rect 1056 1503 1058 1507
rect 1062 1503 1065 1507
rect 1070 1503 1072 1507
rect 1014 1362 1017 1458
rect 1014 1352 1017 1358
rect 1022 1292 1025 1408
rect 1038 1332 1041 1478
rect 1094 1472 1097 1538
rect 1046 1368 1054 1371
rect 1046 1342 1049 1368
rect 1066 1328 1070 1331
rect 886 1051 889 1058
rect 886 1048 894 1051
rect 918 952 921 1118
rect 926 1102 929 1118
rect 894 731 897 918
rect 890 728 897 731
rect 902 662 905 808
rect 894 552 897 618
rect 898 548 902 551
rect 910 472 913 648
rect 858 278 865 281
rect 546 268 550 271
rect 544 203 546 207
rect 550 203 553 207
rect 558 203 560 207
rect 734 182 737 258
rect 842 248 849 251
rect 734 152 737 178
rect 622 52 625 148
rect 846 92 849 248
rect 886 232 889 378
rect 894 352 897 378
rect 918 342 921 658
rect 918 182 921 338
rect 934 161 937 658
rect 942 552 945 1028
rect 1030 862 1033 1298
rect 1038 1022 1041 1328
rect 1078 1312 1081 1438
rect 1056 1303 1058 1307
rect 1062 1303 1065 1307
rect 1070 1303 1072 1307
rect 1046 1252 1049 1268
rect 1086 1252 1089 1348
rect 1090 1248 1094 1251
rect 1078 1242 1081 1248
rect 1102 1232 1105 1358
rect 1118 1352 1121 2198
rect 1142 2158 1150 2161
rect 1126 1492 1129 1958
rect 1142 1852 1145 2158
rect 1174 2062 1177 2248
rect 1126 1452 1129 1458
rect 1158 1332 1161 1728
rect 1114 1268 1118 1271
rect 1166 1242 1169 2048
rect 1182 1751 1185 2118
rect 1182 1748 1190 1751
rect 1214 1742 1217 2218
rect 1270 2208 1278 2211
rect 1214 1692 1217 1738
rect 1194 1678 1198 1681
rect 1206 1432 1209 1688
rect 1222 1442 1225 1648
rect 1262 1482 1265 1858
rect 1270 1712 1273 2208
rect 1270 1561 1273 1668
rect 1270 1558 1278 1561
rect 1294 1542 1297 2298
rect 1302 1942 1305 2128
rect 1318 2022 1321 2258
rect 1350 2152 1353 2248
rect 1302 1882 1305 1938
rect 1198 1352 1201 1368
rect 1174 1262 1177 1268
rect 1194 1248 1198 1251
rect 1056 1103 1058 1107
rect 1062 1103 1065 1107
rect 1070 1103 1072 1107
rect 1038 922 1041 1018
rect 1056 903 1058 907
rect 1062 903 1065 907
rect 1070 903 1072 907
rect 1066 748 1070 751
rect 1094 712 1097 728
rect 1056 703 1058 707
rect 1062 703 1065 707
rect 1070 703 1072 707
rect 950 272 953 698
rect 958 422 961 668
rect 966 662 969 678
rect 1022 352 1025 568
rect 1038 412 1041 648
rect 1056 503 1058 507
rect 1062 503 1065 507
rect 1070 503 1072 507
rect 1086 432 1089 698
rect 1102 371 1105 808
rect 1118 672 1121 848
rect 1126 742 1129 748
rect 1134 632 1137 1078
rect 1214 902 1217 1438
rect 1238 862 1241 1458
rect 1246 1112 1249 1168
rect 1210 668 1214 671
rect 1102 368 1110 371
rect 1058 348 1062 351
rect 1056 303 1058 307
rect 1062 303 1065 307
rect 1070 303 1072 307
rect 934 158 942 161
rect 926 152 929 158
rect 942 62 945 158
rect 950 142 953 268
rect 966 188 974 191
rect 966 82 969 188
rect 994 148 998 151
rect 1056 103 1058 107
rect 1062 103 1065 107
rect 1070 103 1072 107
rect 1134 62 1137 628
rect 1150 542 1153 548
rect 1222 392 1225 668
rect 1238 662 1241 858
rect 1254 772 1257 1228
rect 1286 952 1289 1478
rect 1310 1362 1313 1948
rect 1318 1512 1321 1588
rect 1254 662 1257 768
rect 1278 752 1281 758
rect 1302 722 1305 1148
rect 1246 652 1249 658
rect 1278 512 1281 688
rect 1290 678 1294 681
rect 1302 562 1305 718
rect 1294 482 1297 498
rect 1310 472 1313 948
rect 1318 482 1321 1508
rect 1326 1402 1329 1928
rect 1350 1602 1353 2148
rect 1358 1552 1361 2238
rect 1414 2082 1417 2268
rect 1446 1962 1449 2048
rect 1526 2032 1529 2398
rect 2222 2338 2230 2341
rect 1560 2203 1562 2207
rect 1566 2203 1569 2207
rect 1574 2203 1576 2207
rect 1710 2142 1713 2318
rect 2080 2303 2082 2307
rect 2086 2303 2089 2307
rect 2094 2303 2096 2307
rect 1734 2262 1737 2268
rect 1326 1272 1329 1348
rect 1350 1222 1353 1248
rect 1342 1062 1345 1168
rect 1366 1072 1369 1728
rect 1398 1402 1401 1848
rect 1406 1422 1409 1648
rect 1414 1532 1417 1818
rect 1422 1812 1425 1818
rect 1422 1642 1425 1808
rect 1422 1552 1425 1638
rect 1434 1628 1438 1631
rect 1326 492 1329 788
rect 1342 702 1345 1058
rect 1334 662 1337 668
rect 1342 362 1345 698
rect 1366 662 1369 668
rect 1374 662 1377 1378
rect 1386 1338 1390 1341
rect 1398 1162 1401 1398
rect 1422 1132 1425 1538
rect 1430 1462 1433 1518
rect 1430 1242 1433 1438
rect 1438 1342 1441 1528
rect 1446 1512 1449 1958
rect 1518 1832 1521 1838
rect 1510 1828 1518 1831
rect 1482 1738 1489 1741
rect 1474 1658 1478 1661
rect 1486 1652 1489 1738
rect 1510 1652 1513 1828
rect 1454 1512 1457 1618
rect 1470 1482 1473 1538
rect 1462 1412 1465 1438
rect 1450 1338 1454 1341
rect 1446 1252 1449 1258
rect 1430 1192 1433 1238
rect 1406 692 1409 868
rect 1414 752 1417 1068
rect 1422 942 1425 958
rect 1422 752 1425 758
rect 1358 542 1361 648
rect 1374 642 1377 658
rect 1374 622 1377 638
rect 1398 352 1401 598
rect 1422 552 1425 748
rect 1430 552 1433 588
rect 1438 462 1441 1128
rect 1446 1082 1449 1238
rect 1462 1182 1465 1398
rect 1478 1262 1481 1548
rect 1462 522 1465 638
rect 1182 271 1185 278
rect 1178 268 1185 271
rect 1246 242 1249 318
rect 1470 262 1473 1138
rect 1478 872 1481 1188
rect 1486 1162 1489 1418
rect 1486 1142 1489 1148
rect 1478 692 1481 828
rect 1478 672 1481 688
rect 1478 182 1481 668
rect 1494 662 1497 1558
rect 1526 1162 1529 1358
rect 1542 1332 1545 2018
rect 1560 2003 1562 2007
rect 1566 2003 1569 2007
rect 1574 2003 1576 2007
rect 1550 1512 1553 1948
rect 1560 1803 1562 1807
rect 1566 1803 1569 1807
rect 1574 1803 1576 1807
rect 1560 1603 1562 1607
rect 1566 1603 1569 1607
rect 1574 1603 1576 1607
rect 1566 1552 1569 1568
rect 1550 1342 1553 1408
rect 1560 1403 1562 1407
rect 1566 1403 1569 1407
rect 1574 1403 1576 1407
rect 1582 1392 1585 2078
rect 1590 1662 1593 1908
rect 1502 672 1505 678
rect 1526 572 1529 1158
rect 1550 1072 1553 1338
rect 1598 1272 1601 1678
rect 1606 1452 1609 1488
rect 1560 1203 1562 1207
rect 1566 1203 1569 1207
rect 1574 1203 1576 1207
rect 1538 1058 1542 1061
rect 1550 762 1553 1068
rect 1560 1003 1562 1007
rect 1566 1003 1569 1007
rect 1574 1003 1576 1007
rect 1560 803 1562 807
rect 1566 803 1569 807
rect 1574 803 1576 807
rect 1570 768 1574 771
rect 1560 603 1562 607
rect 1566 603 1569 607
rect 1574 603 1576 607
rect 1590 542 1593 1158
rect 1602 1078 1606 1081
rect 1614 992 1617 1328
rect 1622 852 1625 1508
rect 1630 1442 1633 2048
rect 1662 1662 1665 1938
rect 1670 1872 1673 1898
rect 1638 1332 1641 1658
rect 1606 782 1609 848
rect 1630 842 1633 1068
rect 1646 1042 1649 1328
rect 1654 1072 1657 1338
rect 1662 1232 1665 1658
rect 1670 1522 1673 1688
rect 1670 1342 1673 1498
rect 1678 1262 1681 1728
rect 1694 1662 1697 1768
rect 1686 1592 1689 1648
rect 1686 1512 1689 1588
rect 1702 1572 1705 2118
rect 1698 1548 1702 1551
rect 1698 1538 1702 1541
rect 1690 1358 1694 1361
rect 1682 1248 1686 1251
rect 1630 742 1633 758
rect 1638 592 1641 818
rect 1646 802 1649 1038
rect 1654 712 1657 1068
rect 1666 1058 1670 1061
rect 1666 728 1673 731
rect 1654 662 1657 708
rect 1662 672 1665 708
rect 1662 642 1665 658
rect 1670 652 1673 728
rect 1678 672 1681 1078
rect 1702 722 1705 1008
rect 1694 672 1697 678
rect 1702 662 1705 718
rect 1710 692 1713 2138
rect 1734 1712 1737 1888
rect 1790 1881 1793 2168
rect 1790 1878 1798 1881
rect 1718 1652 1721 1658
rect 1754 1648 1758 1651
rect 1718 1572 1721 1648
rect 1766 1602 1769 1658
rect 1754 1548 1758 1551
rect 1750 1472 1753 1548
rect 1766 1542 1769 1598
rect 1766 1312 1769 1538
rect 1782 1372 1785 1758
rect 1790 1372 1793 1378
rect 1718 1262 1721 1288
rect 1798 1272 1801 1668
rect 1806 1402 1809 1418
rect 1726 862 1729 1108
rect 1734 891 1737 1098
rect 1734 888 1742 891
rect 1766 552 1769 748
rect 1794 708 1798 711
rect 1590 462 1593 538
rect 1560 403 1562 407
rect 1566 403 1569 407
rect 1574 403 1576 407
rect 1670 351 1673 358
rect 1666 348 1673 351
rect 1606 282 1609 328
rect 1678 272 1681 378
rect 1726 272 1729 288
rect 1750 262 1753 338
rect 1560 203 1562 207
rect 1566 203 1569 207
rect 1574 203 1576 207
rect 1594 178 1598 181
rect 1790 132 1793 708
rect 1806 422 1809 1358
rect 1814 952 1817 1708
rect 1822 1462 1825 2138
rect 1998 1872 2001 2138
rect 1982 1842 1985 1848
rect 1870 1662 1873 1678
rect 1902 1622 1905 1658
rect 1822 1362 1825 1398
rect 1870 1352 1873 1568
rect 1870 1042 1873 1348
rect 1822 812 1825 1038
rect 1846 922 1849 1028
rect 1878 922 1881 1448
rect 1918 1172 1921 1738
rect 1930 1688 1934 1691
rect 1942 1632 1945 1658
rect 1958 1652 1961 1658
rect 1962 1568 1966 1571
rect 1974 1362 1977 1778
rect 1990 1342 1993 1738
rect 1998 1352 2001 1748
rect 2006 1462 2009 2058
rect 2062 2002 2065 2118
rect 2080 2103 2082 2107
rect 2086 2103 2089 2107
rect 2094 2103 2096 2107
rect 2118 2092 2121 2218
rect 2038 1852 2041 1938
rect 2080 1903 2082 1907
rect 2086 1903 2089 1907
rect 2094 1903 2096 1907
rect 2080 1703 2082 1707
rect 2086 1703 2089 1707
rect 2094 1703 2096 1707
rect 2014 1672 2017 1678
rect 1994 1338 1998 1341
rect 1926 942 1929 1138
rect 1822 422 1825 808
rect 1830 732 1833 738
rect 1806 362 1809 418
rect 1838 152 1841 908
rect 1870 572 1873 918
rect 1886 871 1889 898
rect 1886 868 1894 871
rect 1890 738 1894 741
rect 1934 592 1937 1198
rect 1942 762 1945 1328
rect 1870 382 1873 568
rect 1890 348 1897 351
rect 1894 342 1897 348
rect 1934 212 1937 588
rect 1942 552 1945 758
rect 1958 592 1961 968
rect 1966 762 1969 1248
rect 1998 1032 2001 1338
rect 2006 1022 2009 1458
rect 2022 1212 2025 1698
rect 2034 1548 2038 1551
rect 1974 822 1977 868
rect 1978 748 1982 751
rect 1998 662 2001 1008
rect 2014 692 2017 738
rect 1966 652 1969 658
rect 2022 352 2025 1208
rect 2030 1152 2033 1428
rect 2038 1112 2041 1348
rect 2062 1262 2065 1648
rect 2070 1532 2073 1598
rect 2070 1312 2073 1528
rect 2080 1503 2082 1507
rect 2086 1503 2089 1507
rect 2094 1503 2096 1507
rect 2078 1422 2081 1448
rect 2080 1303 2082 1307
rect 2086 1303 2089 1307
rect 2094 1303 2096 1307
rect 2102 1292 2105 2048
rect 2110 1672 2113 1688
rect 2110 1342 2113 1598
rect 2082 1288 2086 1291
rect 2054 1242 2057 1258
rect 2102 1112 2105 1148
rect 2080 1103 2082 1107
rect 2086 1103 2089 1107
rect 2094 1103 2096 1107
rect 2090 1078 2094 1081
rect 2110 1032 2113 1338
rect 2118 1152 2121 2058
rect 2222 1962 2225 2338
rect 2130 1958 2134 1961
rect 2126 1692 2129 1698
rect 2158 1352 2161 1938
rect 2262 1762 2265 2158
rect 2278 2102 2281 2118
rect 2170 1658 2174 1661
rect 2166 1362 2169 1628
rect 2230 1592 2233 1748
rect 2198 1352 2201 1528
rect 2194 1348 2198 1351
rect 2062 702 2065 1018
rect 2080 903 2082 907
rect 2086 903 2089 907
rect 2094 903 2096 907
rect 2030 662 2033 668
rect 2062 402 2065 648
rect 2014 272 2017 338
rect 2070 262 2073 778
rect 2102 752 2105 768
rect 2080 703 2082 707
rect 2086 703 2089 707
rect 2094 703 2096 707
rect 2110 612 2113 1028
rect 2080 503 2082 507
rect 2086 503 2089 507
rect 2094 503 2096 507
rect 2118 462 2121 1148
rect 2126 1052 2129 1088
rect 2158 712 2161 1348
rect 2186 868 2190 871
rect 2166 622 2169 858
rect 2214 822 2217 918
rect 2230 782 2233 868
rect 2238 812 2241 1728
rect 2246 1612 2249 1748
rect 2278 1742 2281 2068
rect 2294 2022 2297 2068
rect 2294 1732 2297 2018
rect 2310 1752 2313 2028
rect 2342 1892 2345 2248
rect 2342 1862 2345 1888
rect 2374 1862 2377 2228
rect 2190 312 2193 658
rect 2080 303 2082 307
rect 2086 303 2089 307
rect 2094 303 2096 307
rect 2078 272 2081 278
rect 1790 92 1793 128
rect 2080 103 2082 107
rect 2086 103 2089 107
rect 2094 103 2096 107
rect 2198 82 2201 458
rect 2262 372 2265 1428
rect 2270 1162 2273 1168
rect 2302 1082 2305 1278
rect 2310 1202 2313 1748
rect 2318 1242 2321 1468
rect 2342 1342 2345 1858
rect 2350 1662 2353 1818
rect 2294 562 2297 718
rect 2310 552 2313 758
rect 2318 662 2321 808
rect 2310 462 2313 548
rect 2326 362 2329 1158
rect 2350 812 2353 1658
rect 2374 1182 2377 1858
rect 2382 1672 2385 1908
rect 2462 1802 2465 2248
rect 2470 1862 2473 2258
rect 2382 1472 2385 1668
rect 2382 1362 2385 1468
rect 2206 288 2214 291
rect 2206 152 2209 288
rect 2326 172 2329 358
rect 2374 302 2377 1178
rect 2398 1072 2401 1268
rect 2446 1232 2449 1728
rect 2462 1652 2465 1798
rect 2470 1242 2473 1858
rect 2486 1541 2489 1738
rect 2482 1538 2489 1541
rect 2426 798 2433 801
rect 2374 202 2377 298
rect 2382 272 2385 778
rect 2390 72 2393 738
rect 2402 678 2406 681
rect 2422 492 2425 688
rect 2430 442 2433 798
rect 2438 422 2441 718
rect 2454 542 2457 728
rect 2470 252 2473 1238
rect 2478 682 2481 1178
rect 2486 962 2489 1448
rect 2486 662 2489 758
rect 2518 182 2521 658
rect 2526 162 2529 2168
rect 2542 452 2545 1548
rect 2542 192 2545 448
rect 2550 332 2553 2218
rect 2558 1172 2561 1968
rect 2578 1668 2582 1671
rect 2574 1292 2577 1638
rect 2590 1552 2593 2108
rect 2574 1122 2577 1288
rect 2582 1152 2585 1368
rect 2574 882 2577 1118
rect 2598 1051 2601 1478
rect 2630 1192 2633 1428
rect 2646 1292 2649 1298
rect 2598 1048 2606 1051
rect 2598 402 2601 558
rect 2550 192 2553 328
rect 1762 58 1766 61
rect 544 3 546 7
rect 550 3 553 7
rect 558 3 560 7
rect 1560 3 1562 7
rect 1566 3 1569 7
rect 1574 3 1576 7
<< m5contact >>
rect 546 2403 550 2407
rect 553 2403 554 2407
rect 554 2403 557 2407
rect 1562 2403 1566 2407
rect 1569 2403 1570 2407
rect 1570 2403 1573 2407
rect 1058 2303 1062 2307
rect 1065 2303 1066 2307
rect 1066 2303 1069 2307
rect 1262 2258 1266 2262
rect 302 2058 306 2062
rect 278 1368 282 1372
rect 294 1328 298 1332
rect 546 2203 550 2207
rect 553 2203 554 2207
rect 554 2203 557 2207
rect 446 2058 450 2062
rect 422 1928 426 1932
rect 358 1738 362 1742
rect 398 1728 402 1732
rect 390 1658 394 1662
rect 358 1368 362 1372
rect 294 1278 298 1282
rect 198 178 202 182
rect 446 1748 450 1752
rect 470 1738 474 1742
rect 486 1728 490 1732
rect 546 2003 550 2007
rect 553 2003 554 2007
rect 554 2003 557 2007
rect 546 1803 550 1807
rect 553 1803 554 1807
rect 554 1803 557 1807
rect 478 1468 482 1472
rect 454 1278 458 1282
rect 478 1248 482 1252
rect 350 628 354 632
rect 414 678 418 682
rect 462 638 466 642
rect 486 648 490 652
rect 546 1603 550 1607
rect 553 1603 554 1607
rect 554 1603 557 1607
rect 546 1403 550 1407
rect 553 1403 554 1407
rect 554 1403 557 1407
rect 546 1203 550 1207
rect 553 1203 554 1207
rect 554 1203 557 1207
rect 546 1003 550 1007
rect 553 1003 554 1007
rect 554 1003 557 1007
rect 546 803 550 807
rect 553 803 554 807
rect 554 803 557 807
rect 566 658 570 662
rect 574 648 578 652
rect 494 628 498 632
rect 546 603 550 607
rect 553 603 554 607
rect 554 603 557 607
rect 546 403 550 407
rect 553 403 554 407
rect 554 403 557 407
rect 598 348 602 352
rect 1058 2103 1062 2107
rect 1065 2103 1066 2107
rect 1066 2103 1069 2107
rect 654 1258 658 1262
rect 662 668 666 672
rect 758 1658 762 1662
rect 806 1928 810 1932
rect 814 1748 818 1752
rect 758 1258 762 1262
rect 798 1468 802 1472
rect 814 1258 818 1262
rect 854 1268 858 1272
rect 742 638 746 642
rect 630 278 634 282
rect 1058 1903 1062 1907
rect 1065 1903 1066 1907
rect 1066 1903 1069 1907
rect 958 1658 962 1662
rect 1038 1728 1042 1732
rect 1058 1703 1062 1707
rect 1065 1703 1066 1707
rect 1066 1703 1069 1707
rect 1046 1668 1050 1672
rect 982 1458 986 1462
rect 1058 1503 1062 1507
rect 1065 1503 1066 1507
rect 1066 1503 1069 1507
rect 1014 1358 1018 1362
rect 1046 1338 1050 1342
rect 1062 1328 1066 1332
rect 934 658 938 662
rect 902 548 906 552
rect 550 268 554 272
rect 546 203 550 207
rect 553 203 554 207
rect 554 203 557 207
rect 734 178 738 182
rect 918 178 922 182
rect 1058 1303 1062 1307
rect 1065 1303 1066 1307
rect 1066 1303 1069 1307
rect 1046 1248 1050 1252
rect 1094 1248 1098 1252
rect 1078 1238 1082 1242
rect 1126 1448 1130 1452
rect 1110 1268 1114 1272
rect 1214 1738 1218 1742
rect 1198 1678 1202 1682
rect 1238 1458 1242 1462
rect 1198 1348 1202 1352
rect 1174 1268 1178 1272
rect 1190 1248 1194 1252
rect 1058 1103 1062 1107
rect 1065 1103 1066 1107
rect 1066 1103 1069 1107
rect 1058 903 1062 907
rect 1065 903 1066 907
rect 1066 903 1069 907
rect 1062 748 1066 752
rect 1094 708 1098 712
rect 1058 703 1062 707
rect 1065 703 1066 707
rect 1066 703 1069 707
rect 966 678 970 682
rect 1058 503 1062 507
rect 1065 503 1066 507
rect 1066 503 1069 507
rect 1126 748 1130 752
rect 1214 668 1218 672
rect 1134 628 1138 632
rect 1054 348 1058 352
rect 1058 303 1062 307
rect 1065 303 1066 307
rect 1066 303 1069 307
rect 950 268 954 272
rect 926 148 930 152
rect 990 148 994 152
rect 1058 103 1062 107
rect 1065 103 1066 107
rect 1066 103 1069 107
rect 1150 538 1154 542
rect 1318 1588 1322 1592
rect 1278 748 1282 752
rect 1238 658 1242 662
rect 1246 648 1250 652
rect 1286 678 1290 682
rect 1562 2203 1566 2207
rect 1569 2203 1570 2207
rect 1570 2203 1573 2207
rect 2082 2303 2086 2307
rect 2089 2303 2090 2307
rect 2090 2303 2093 2307
rect 1734 2258 1738 2262
rect 1446 1958 1450 1962
rect 1350 1248 1354 1252
rect 1406 1648 1410 1652
rect 1438 1628 1442 1632
rect 1422 1548 1426 1552
rect 1334 658 1338 662
rect 1366 668 1370 672
rect 1382 1338 1386 1342
rect 1430 1458 1434 1462
rect 1518 1838 1522 1842
rect 1478 1658 1482 1662
rect 1478 1548 1482 1552
rect 1470 1538 1474 1542
rect 1446 1338 1450 1342
rect 1446 1258 1450 1262
rect 1422 758 1426 762
rect 1342 358 1346 362
rect 1430 548 1434 552
rect 1462 638 1466 642
rect 1182 278 1186 282
rect 1486 1138 1490 1142
rect 1478 688 1482 692
rect 1562 2003 1566 2007
rect 1569 2003 1570 2007
rect 1570 2003 1573 2007
rect 1562 1803 1566 1807
rect 1569 1803 1570 1807
rect 1570 1803 1573 1807
rect 1562 1603 1566 1607
rect 1569 1603 1570 1607
rect 1570 1603 1573 1607
rect 1566 1548 1570 1552
rect 1562 1403 1566 1407
rect 1569 1403 1570 1407
rect 1570 1403 1573 1407
rect 1550 1338 1554 1342
rect 1526 1158 1530 1162
rect 1502 678 1506 682
rect 1562 1203 1566 1207
rect 1569 1203 1570 1207
rect 1570 1203 1573 1207
rect 1542 1058 1546 1062
rect 1562 1003 1566 1007
rect 1569 1003 1570 1007
rect 1570 1003 1573 1007
rect 1562 803 1566 807
rect 1569 803 1570 807
rect 1570 803 1573 807
rect 1574 768 1578 772
rect 1562 603 1566 607
rect 1569 603 1570 607
rect 1570 603 1573 607
rect 1598 1078 1602 1082
rect 1662 1658 1666 1662
rect 1686 1588 1690 1592
rect 1694 1548 1698 1552
rect 1694 1538 1698 1542
rect 1694 1358 1698 1362
rect 1686 1248 1690 1252
rect 1662 1058 1666 1062
rect 1662 668 1666 672
rect 1654 658 1658 662
rect 1694 678 1698 682
rect 1718 1648 1722 1652
rect 1758 1648 1762 1652
rect 1718 1568 1722 1572
rect 1750 1548 1754 1552
rect 1790 1368 1794 1372
rect 1710 688 1714 692
rect 1662 638 1666 642
rect 1790 708 1794 712
rect 1590 538 1594 542
rect 1562 403 1566 407
rect 1569 403 1570 407
rect 1570 403 1573 407
rect 1670 358 1674 362
rect 1726 268 1730 272
rect 1562 203 1566 207
rect 1569 203 1570 207
rect 1570 203 1573 207
rect 1590 178 1594 182
rect 1982 1838 1986 1842
rect 1870 1678 1874 1682
rect 1822 1358 1826 1362
rect 1870 1348 1874 1352
rect 1926 1688 1930 1692
rect 1958 1648 1962 1652
rect 1942 1628 1946 1632
rect 1958 1568 1962 1572
rect 2082 2103 2086 2107
rect 2089 2103 2090 2107
rect 2090 2103 2093 2107
rect 2082 1903 2086 1907
rect 2089 1903 2090 1907
rect 2090 1903 2093 1907
rect 2082 1703 2086 1707
rect 2089 1703 2090 1707
rect 2090 1703 2093 1707
rect 2014 1678 2018 1682
rect 1990 1338 1994 1342
rect 1830 738 1834 742
rect 1886 738 1890 742
rect 1942 758 1946 762
rect 2030 1548 2034 1552
rect 1974 868 1978 872
rect 1974 748 1978 752
rect 2014 688 2018 692
rect 1966 648 1970 652
rect 2082 1503 2086 1507
rect 2089 1503 2090 1507
rect 2090 1503 2093 1507
rect 2078 1448 2082 1452
rect 2082 1303 2086 1307
rect 2089 1303 2090 1307
rect 2090 1303 2093 1307
rect 2110 1668 2114 1672
rect 2086 1288 2090 1292
rect 2054 1238 2058 1242
rect 2102 1148 2106 1152
rect 2082 1103 2086 1107
rect 2089 1103 2090 1107
rect 2090 1103 2093 1107
rect 2086 1078 2090 1082
rect 2126 1958 2130 1962
rect 2126 1688 2130 1692
rect 2166 1658 2170 1662
rect 2198 1348 2202 1352
rect 2082 903 2086 907
rect 2089 903 2090 907
rect 2090 903 2093 907
rect 2030 668 2034 672
rect 2102 768 2106 772
rect 2082 703 2086 707
rect 2089 703 2090 707
rect 2090 703 2093 707
rect 2082 503 2086 507
rect 2089 503 2090 507
rect 2090 503 2093 507
rect 2182 868 2186 872
rect 2082 303 2086 307
rect 2089 303 2090 307
rect 2090 303 2093 307
rect 2078 278 2082 282
rect 2082 103 2086 107
rect 2089 103 2090 107
rect 2090 103 2093 107
rect 2270 1168 2274 1172
rect 2398 678 2402 682
rect 2574 1668 2578 1672
rect 2646 1288 2650 1292
rect 942 58 946 62
rect 1758 58 1762 62
rect 546 3 550 7
rect 553 3 554 7
rect 554 3 557 7
rect 1562 3 1566 7
rect 1569 3 1570 7
rect 1570 3 1573 7
<< metal5 >>
rect 550 2403 553 2407
rect 549 2402 554 2403
rect 559 2402 560 2407
rect 1566 2403 1569 2407
rect 1565 2402 1570 2403
rect 1575 2402 1576 2407
rect 1062 2303 1065 2307
rect 1061 2302 1066 2303
rect 1071 2302 1072 2307
rect 2086 2303 2089 2307
rect 2085 2302 2090 2303
rect 2095 2302 2096 2307
rect 1266 2258 1734 2261
rect 550 2203 553 2207
rect 549 2202 554 2203
rect 559 2202 560 2207
rect 1566 2203 1569 2207
rect 1565 2202 1570 2203
rect 1575 2202 1576 2207
rect 1062 2103 1065 2107
rect 1061 2102 1066 2103
rect 1071 2102 1072 2107
rect 2086 2103 2089 2107
rect 2085 2102 2090 2103
rect 2095 2102 2096 2107
rect 306 2058 446 2061
rect 550 2003 553 2007
rect 549 2002 554 2003
rect 559 2002 560 2007
rect 1566 2003 1569 2007
rect 1565 2002 1570 2003
rect 1575 2002 1576 2007
rect 1450 1958 2126 1961
rect 426 1928 806 1931
rect 1062 1903 1065 1907
rect 1061 1902 1066 1903
rect 1071 1902 1072 1907
rect 2086 1903 2089 1907
rect 2085 1902 2090 1903
rect 2095 1902 2096 1907
rect 1522 1838 1982 1841
rect 550 1803 553 1807
rect 549 1802 554 1803
rect 559 1802 560 1807
rect 1566 1803 1569 1807
rect 1565 1802 1570 1803
rect 1575 1802 1576 1807
rect 450 1748 814 1751
rect 362 1738 401 1741
rect 474 1738 1214 1741
rect 398 1732 401 1738
rect 490 1728 1038 1731
rect 1062 1703 1065 1707
rect 1061 1702 1066 1703
rect 1071 1702 1072 1707
rect 2086 1703 2089 1707
rect 2085 1702 2090 1703
rect 2095 1702 2096 1707
rect 1930 1688 2126 1691
rect 1202 1678 1870 1681
rect 2014 1671 2017 1678
rect 1050 1668 2017 1671
rect 2114 1668 2574 1671
rect 394 1658 758 1661
rect 962 1658 1478 1661
rect 1666 1658 2166 1661
rect 1410 1648 1718 1651
rect 1762 1648 1958 1651
rect 1442 1628 1942 1631
rect 550 1603 553 1607
rect 549 1602 554 1603
rect 559 1602 560 1607
rect 1566 1603 1569 1607
rect 1565 1602 1570 1603
rect 1575 1602 1576 1607
rect 1322 1588 1686 1591
rect 1722 1568 1958 1571
rect 1426 1548 1478 1551
rect 1570 1548 1694 1551
rect 1754 1548 2030 1551
rect 1474 1538 1694 1541
rect 1062 1503 1065 1507
rect 1061 1502 1066 1503
rect 1071 1502 1072 1507
rect 2086 1503 2089 1507
rect 2085 1502 2090 1503
rect 2095 1502 2096 1507
rect 482 1468 798 1471
rect 986 1458 1238 1461
rect 1242 1458 1430 1461
rect 1130 1448 2078 1451
rect 550 1403 553 1407
rect 549 1402 554 1403
rect 559 1402 560 1407
rect 1566 1403 1569 1407
rect 1565 1402 1570 1403
rect 1575 1402 1576 1407
rect 282 1368 358 1371
rect 362 1368 1790 1371
rect 1698 1358 1822 1361
rect 1014 1351 1017 1358
rect 1014 1348 1198 1351
rect 1874 1348 2198 1351
rect 1050 1338 1382 1341
rect 1386 1338 1446 1341
rect 1554 1338 1990 1341
rect 298 1328 1062 1331
rect 1062 1303 1065 1307
rect 1061 1302 1066 1303
rect 1071 1302 1072 1307
rect 2086 1303 2089 1307
rect 2085 1302 2090 1303
rect 2095 1302 2096 1307
rect 2090 1288 2646 1291
rect 298 1278 454 1281
rect 858 1268 1110 1271
rect 658 1258 758 1261
rect 762 1258 814 1261
rect 1174 1261 1177 1268
rect 1174 1258 1446 1261
rect 482 1248 1046 1251
rect 1098 1248 1190 1251
rect 1354 1248 1686 1251
rect 1082 1238 2054 1241
rect 550 1203 553 1207
rect 549 1202 554 1203
rect 559 1202 560 1207
rect 1566 1203 1569 1207
rect 1565 1202 1570 1203
rect 1575 1202 1576 1207
rect 2270 1161 2273 1168
rect 1530 1158 2273 1161
rect 1486 1148 2102 1151
rect 1486 1142 1489 1148
rect 1062 1103 1065 1107
rect 1061 1102 1066 1103
rect 1071 1102 1072 1107
rect 2086 1103 2089 1107
rect 2085 1102 2090 1103
rect 2095 1102 2096 1107
rect 1602 1078 2086 1081
rect 1546 1058 1662 1061
rect 550 1003 553 1007
rect 549 1002 554 1003
rect 559 1002 560 1007
rect 1566 1003 1569 1007
rect 1565 1002 1570 1003
rect 1575 1002 1576 1007
rect 1062 903 1065 907
rect 1061 902 1066 903
rect 1071 902 1072 907
rect 2086 903 2089 907
rect 2085 902 2090 903
rect 2095 902 2096 907
rect 1978 868 2182 871
rect 550 803 553 807
rect 549 802 554 803
rect 559 802 560 807
rect 1566 803 1569 807
rect 1565 802 1570 803
rect 1575 802 1576 807
rect 1578 768 2102 771
rect 1426 758 1942 761
rect 1066 748 1126 751
rect 1282 748 1974 751
rect 1834 738 1886 741
rect 1098 708 1790 711
rect 1062 703 1065 707
rect 1061 702 1066 703
rect 1071 702 1072 707
rect 2086 703 2089 707
rect 2085 702 2090 703
rect 2095 702 2096 707
rect 1482 688 1710 691
rect 1714 688 2014 691
rect 418 678 966 681
rect 1290 678 1502 681
rect 1698 678 2398 681
rect 1218 668 1337 671
rect 1370 668 1662 671
rect 662 661 665 668
rect 1334 662 1337 668
rect 570 658 665 661
rect 938 658 1238 661
rect 2030 661 2033 668
rect 1658 658 2033 661
rect 490 648 574 651
rect 1250 648 1966 651
rect 466 638 742 641
rect 1466 638 1662 641
rect 354 628 494 631
rect 498 628 1134 631
rect 550 603 553 607
rect 549 602 554 603
rect 559 602 560 607
rect 1566 603 1569 607
rect 1565 602 1570 603
rect 1575 602 1576 607
rect 906 548 1430 551
rect 1154 538 1590 541
rect 1062 503 1065 507
rect 1061 502 1066 503
rect 1071 502 1072 507
rect 2086 503 2089 507
rect 2085 502 2090 503
rect 2095 502 2096 507
rect 550 403 553 407
rect 549 402 554 403
rect 559 402 560 407
rect 1566 403 1569 407
rect 1565 402 1570 403
rect 1575 402 1576 407
rect 1346 358 1670 361
rect 602 348 1054 351
rect 1062 303 1065 307
rect 1061 302 1066 303
rect 1071 302 1072 307
rect 2086 303 2089 307
rect 2085 302 2090 303
rect 2095 302 2096 307
rect 634 278 1182 281
rect 554 268 950 271
rect 2078 271 2081 278
rect 1730 268 2081 271
rect 550 203 553 207
rect 549 202 554 203
rect 559 202 560 207
rect 1566 203 1569 207
rect 1565 202 1570 203
rect 1575 202 1576 207
rect 202 178 734 181
rect 922 178 1590 181
rect 930 148 990 151
rect 1062 103 1065 107
rect 1061 102 1066 103
rect 1071 102 1072 107
rect 2086 103 2089 107
rect 2085 102 2090 103
rect 2095 102 2096 107
rect 946 58 1758 61
rect 550 3 553 7
rect 549 2 554 3
rect 559 2 560 7
rect 1566 3 1569 7
rect 1565 2 1570 3
rect 1575 2 1576 7
<< m6contact >>
rect 544 2403 546 2407
rect 546 2403 549 2407
rect 554 2403 557 2407
rect 557 2403 559 2407
rect 544 2402 549 2403
rect 554 2402 559 2403
rect 1560 2403 1562 2407
rect 1562 2403 1565 2407
rect 1570 2403 1573 2407
rect 1573 2403 1575 2407
rect 1560 2402 1565 2403
rect 1570 2402 1575 2403
rect 1056 2303 1058 2307
rect 1058 2303 1061 2307
rect 1066 2303 1069 2307
rect 1069 2303 1071 2307
rect 1056 2302 1061 2303
rect 1066 2302 1071 2303
rect 2080 2303 2082 2307
rect 2082 2303 2085 2307
rect 2090 2303 2093 2307
rect 2093 2303 2095 2307
rect 2080 2302 2085 2303
rect 2090 2302 2095 2303
rect 544 2203 546 2207
rect 546 2203 549 2207
rect 554 2203 557 2207
rect 557 2203 559 2207
rect 544 2202 549 2203
rect 554 2202 559 2203
rect 1560 2203 1562 2207
rect 1562 2203 1565 2207
rect 1570 2203 1573 2207
rect 1573 2203 1575 2207
rect 1560 2202 1565 2203
rect 1570 2202 1575 2203
rect 1056 2103 1058 2107
rect 1058 2103 1061 2107
rect 1066 2103 1069 2107
rect 1069 2103 1071 2107
rect 1056 2102 1061 2103
rect 1066 2102 1071 2103
rect 2080 2103 2082 2107
rect 2082 2103 2085 2107
rect 2090 2103 2093 2107
rect 2093 2103 2095 2107
rect 2080 2102 2085 2103
rect 2090 2102 2095 2103
rect 544 2003 546 2007
rect 546 2003 549 2007
rect 554 2003 557 2007
rect 557 2003 559 2007
rect 544 2002 549 2003
rect 554 2002 559 2003
rect 1560 2003 1562 2007
rect 1562 2003 1565 2007
rect 1570 2003 1573 2007
rect 1573 2003 1575 2007
rect 1560 2002 1565 2003
rect 1570 2002 1575 2003
rect 1056 1903 1058 1907
rect 1058 1903 1061 1907
rect 1066 1903 1069 1907
rect 1069 1903 1071 1907
rect 1056 1902 1061 1903
rect 1066 1902 1071 1903
rect 2080 1903 2082 1907
rect 2082 1903 2085 1907
rect 2090 1903 2093 1907
rect 2093 1903 2095 1907
rect 2080 1902 2085 1903
rect 2090 1902 2095 1903
rect 544 1803 546 1807
rect 546 1803 549 1807
rect 554 1803 557 1807
rect 557 1803 559 1807
rect 544 1802 549 1803
rect 554 1802 559 1803
rect 1560 1803 1562 1807
rect 1562 1803 1565 1807
rect 1570 1803 1573 1807
rect 1573 1803 1575 1807
rect 1560 1802 1565 1803
rect 1570 1802 1575 1803
rect 1056 1703 1058 1707
rect 1058 1703 1061 1707
rect 1066 1703 1069 1707
rect 1069 1703 1071 1707
rect 1056 1702 1061 1703
rect 1066 1702 1071 1703
rect 2080 1703 2082 1707
rect 2082 1703 2085 1707
rect 2090 1703 2093 1707
rect 2093 1703 2095 1707
rect 2080 1702 2085 1703
rect 2090 1702 2095 1703
rect 544 1603 546 1607
rect 546 1603 549 1607
rect 554 1603 557 1607
rect 557 1603 559 1607
rect 544 1602 549 1603
rect 554 1602 559 1603
rect 1560 1603 1562 1607
rect 1562 1603 1565 1607
rect 1570 1603 1573 1607
rect 1573 1603 1575 1607
rect 1560 1602 1565 1603
rect 1570 1602 1575 1603
rect 1056 1503 1058 1507
rect 1058 1503 1061 1507
rect 1066 1503 1069 1507
rect 1069 1503 1071 1507
rect 1056 1502 1061 1503
rect 1066 1502 1071 1503
rect 2080 1503 2082 1507
rect 2082 1503 2085 1507
rect 2090 1503 2093 1507
rect 2093 1503 2095 1507
rect 2080 1502 2085 1503
rect 2090 1502 2095 1503
rect 544 1403 546 1407
rect 546 1403 549 1407
rect 554 1403 557 1407
rect 557 1403 559 1407
rect 544 1402 549 1403
rect 554 1402 559 1403
rect 1560 1403 1562 1407
rect 1562 1403 1565 1407
rect 1570 1403 1573 1407
rect 1573 1403 1575 1407
rect 1560 1402 1565 1403
rect 1570 1402 1575 1403
rect 1056 1303 1058 1307
rect 1058 1303 1061 1307
rect 1066 1303 1069 1307
rect 1069 1303 1071 1307
rect 1056 1302 1061 1303
rect 1066 1302 1071 1303
rect 2080 1303 2082 1307
rect 2082 1303 2085 1307
rect 2090 1303 2093 1307
rect 2093 1303 2095 1307
rect 2080 1302 2085 1303
rect 2090 1302 2095 1303
rect 544 1203 546 1207
rect 546 1203 549 1207
rect 554 1203 557 1207
rect 557 1203 559 1207
rect 544 1202 549 1203
rect 554 1202 559 1203
rect 1560 1203 1562 1207
rect 1562 1203 1565 1207
rect 1570 1203 1573 1207
rect 1573 1203 1575 1207
rect 1560 1202 1565 1203
rect 1570 1202 1575 1203
rect 1056 1103 1058 1107
rect 1058 1103 1061 1107
rect 1066 1103 1069 1107
rect 1069 1103 1071 1107
rect 1056 1102 1061 1103
rect 1066 1102 1071 1103
rect 2080 1103 2082 1107
rect 2082 1103 2085 1107
rect 2090 1103 2093 1107
rect 2093 1103 2095 1107
rect 2080 1102 2085 1103
rect 2090 1102 2095 1103
rect 544 1003 546 1007
rect 546 1003 549 1007
rect 554 1003 557 1007
rect 557 1003 559 1007
rect 544 1002 549 1003
rect 554 1002 559 1003
rect 1560 1003 1562 1007
rect 1562 1003 1565 1007
rect 1570 1003 1573 1007
rect 1573 1003 1575 1007
rect 1560 1002 1565 1003
rect 1570 1002 1575 1003
rect 1056 903 1058 907
rect 1058 903 1061 907
rect 1066 903 1069 907
rect 1069 903 1071 907
rect 1056 902 1061 903
rect 1066 902 1071 903
rect 2080 903 2082 907
rect 2082 903 2085 907
rect 2090 903 2093 907
rect 2093 903 2095 907
rect 2080 902 2085 903
rect 2090 902 2095 903
rect 544 803 546 807
rect 546 803 549 807
rect 554 803 557 807
rect 557 803 559 807
rect 544 802 549 803
rect 554 802 559 803
rect 1560 803 1562 807
rect 1562 803 1565 807
rect 1570 803 1573 807
rect 1573 803 1575 807
rect 1560 802 1565 803
rect 1570 802 1575 803
rect 1056 703 1058 707
rect 1058 703 1061 707
rect 1066 703 1069 707
rect 1069 703 1071 707
rect 1056 702 1061 703
rect 1066 702 1071 703
rect 2080 703 2082 707
rect 2082 703 2085 707
rect 2090 703 2093 707
rect 2093 703 2095 707
rect 2080 702 2085 703
rect 2090 702 2095 703
rect 544 603 546 607
rect 546 603 549 607
rect 554 603 557 607
rect 557 603 559 607
rect 544 602 549 603
rect 554 602 559 603
rect 1560 603 1562 607
rect 1562 603 1565 607
rect 1570 603 1573 607
rect 1573 603 1575 607
rect 1560 602 1565 603
rect 1570 602 1575 603
rect 1056 503 1058 507
rect 1058 503 1061 507
rect 1066 503 1069 507
rect 1069 503 1071 507
rect 1056 502 1061 503
rect 1066 502 1071 503
rect 2080 503 2082 507
rect 2082 503 2085 507
rect 2090 503 2093 507
rect 2093 503 2095 507
rect 2080 502 2085 503
rect 2090 502 2095 503
rect 544 403 546 407
rect 546 403 549 407
rect 554 403 557 407
rect 557 403 559 407
rect 544 402 549 403
rect 554 402 559 403
rect 1560 403 1562 407
rect 1562 403 1565 407
rect 1570 403 1573 407
rect 1573 403 1575 407
rect 1560 402 1565 403
rect 1570 402 1575 403
rect 1056 303 1058 307
rect 1058 303 1061 307
rect 1066 303 1069 307
rect 1069 303 1071 307
rect 1056 302 1061 303
rect 1066 302 1071 303
rect 2080 303 2082 307
rect 2082 303 2085 307
rect 2090 303 2093 307
rect 2093 303 2095 307
rect 2080 302 2085 303
rect 2090 302 2095 303
rect 544 203 546 207
rect 546 203 549 207
rect 554 203 557 207
rect 557 203 559 207
rect 544 202 549 203
rect 554 202 559 203
rect 1560 203 1562 207
rect 1562 203 1565 207
rect 1570 203 1573 207
rect 1573 203 1575 207
rect 1560 202 1565 203
rect 1570 202 1575 203
rect 1056 103 1058 107
rect 1058 103 1061 107
rect 1066 103 1069 107
rect 1069 103 1071 107
rect 1056 102 1061 103
rect 1066 102 1071 103
rect 2080 103 2082 107
rect 2082 103 2085 107
rect 2090 103 2093 107
rect 2093 103 2095 107
rect 2080 102 2085 103
rect 2090 102 2095 103
rect 544 3 546 7
rect 546 3 549 7
rect 554 3 557 7
rect 557 3 559 7
rect 544 2 549 3
rect 554 2 559 3
rect 1560 3 1562 7
rect 1562 3 1565 7
rect 1570 3 1573 7
rect 1573 3 1575 7
rect 1560 2 1565 3
rect 1570 2 1575 3
<< metal6 >>
rect 544 2407 560 2430
rect 549 2402 554 2407
rect 559 2402 560 2407
rect 544 2207 560 2402
rect 549 2202 554 2207
rect 559 2202 560 2207
rect 544 2007 560 2202
rect 549 2002 554 2007
rect 559 2002 560 2007
rect 544 1807 560 2002
rect 549 1802 554 1807
rect 559 1802 560 1807
rect 544 1607 560 1802
rect 549 1602 554 1607
rect 559 1602 560 1607
rect 544 1407 560 1602
rect 549 1402 554 1407
rect 559 1402 560 1407
rect 544 1207 560 1402
rect 549 1202 554 1207
rect 559 1202 560 1207
rect 544 1007 560 1202
rect 549 1002 554 1007
rect 559 1002 560 1007
rect 544 807 560 1002
rect 549 802 554 807
rect 559 802 560 807
rect 544 607 560 802
rect 549 602 554 607
rect 559 602 560 607
rect 544 407 560 602
rect 549 402 554 407
rect 559 402 560 407
rect 544 207 560 402
rect 549 202 554 207
rect 559 202 560 207
rect 544 7 560 202
rect 549 2 554 7
rect 559 2 560 7
rect 544 -30 560 2
rect 1056 2307 1072 2430
rect 1061 2302 1066 2307
rect 1071 2302 1072 2307
rect 1056 2107 1072 2302
rect 1061 2102 1066 2107
rect 1071 2102 1072 2107
rect 1056 1907 1072 2102
rect 1061 1902 1066 1907
rect 1071 1902 1072 1907
rect 1056 1707 1072 1902
rect 1061 1702 1066 1707
rect 1071 1702 1072 1707
rect 1056 1507 1072 1702
rect 1061 1502 1066 1507
rect 1071 1502 1072 1507
rect 1056 1307 1072 1502
rect 1061 1302 1066 1307
rect 1071 1302 1072 1307
rect 1056 1107 1072 1302
rect 1061 1102 1066 1107
rect 1071 1102 1072 1107
rect 1056 907 1072 1102
rect 1061 902 1066 907
rect 1071 902 1072 907
rect 1056 707 1072 902
rect 1061 702 1066 707
rect 1071 702 1072 707
rect 1056 507 1072 702
rect 1061 502 1066 507
rect 1071 502 1072 507
rect 1056 307 1072 502
rect 1061 302 1066 307
rect 1071 302 1072 307
rect 1056 107 1072 302
rect 1061 102 1066 107
rect 1071 102 1072 107
rect 1056 -30 1072 102
rect 1560 2407 1576 2430
rect 1565 2402 1570 2407
rect 1575 2402 1576 2407
rect 1560 2207 1576 2402
rect 1565 2202 1570 2207
rect 1575 2202 1576 2207
rect 1560 2007 1576 2202
rect 1565 2002 1570 2007
rect 1575 2002 1576 2007
rect 1560 1807 1576 2002
rect 1565 1802 1570 1807
rect 1575 1802 1576 1807
rect 1560 1607 1576 1802
rect 1565 1602 1570 1607
rect 1575 1602 1576 1607
rect 1560 1407 1576 1602
rect 1565 1402 1570 1407
rect 1575 1402 1576 1407
rect 1560 1207 1576 1402
rect 1565 1202 1570 1207
rect 1575 1202 1576 1207
rect 1560 1007 1576 1202
rect 1565 1002 1570 1007
rect 1575 1002 1576 1007
rect 1560 807 1576 1002
rect 1565 802 1570 807
rect 1575 802 1576 807
rect 1560 607 1576 802
rect 1565 602 1570 607
rect 1575 602 1576 607
rect 1560 407 1576 602
rect 1565 402 1570 407
rect 1575 402 1576 407
rect 1560 207 1576 402
rect 1565 202 1570 207
rect 1575 202 1576 207
rect 1560 7 1576 202
rect 1565 2 1570 7
rect 1575 2 1576 7
rect 1560 -30 1576 2
rect 2080 2307 2096 2430
rect 2085 2302 2090 2307
rect 2095 2302 2096 2307
rect 2080 2107 2096 2302
rect 2085 2102 2090 2107
rect 2095 2102 2096 2107
rect 2080 1907 2096 2102
rect 2085 1902 2090 1907
rect 2095 1902 2096 1907
rect 2080 1707 2096 1902
rect 2085 1702 2090 1707
rect 2095 1702 2096 1707
rect 2080 1507 2096 1702
rect 2085 1502 2090 1507
rect 2095 1502 2096 1507
rect 2080 1307 2096 1502
rect 2085 1302 2090 1307
rect 2095 1302 2096 1307
rect 2080 1107 2096 1302
rect 2085 1102 2090 1107
rect 2095 1102 2096 1107
rect 2080 907 2096 1102
rect 2085 902 2090 907
rect 2095 902 2096 907
rect 2080 707 2096 902
rect 2085 702 2090 707
rect 2095 702 2096 707
rect 2080 507 2096 702
rect 2085 502 2090 507
rect 2095 502 2096 507
rect 2080 307 2096 502
rect 2085 302 2090 307
rect 2095 302 2096 307
rect 2080 107 2096 302
rect 2085 102 2090 107
rect 2095 102 2096 107
rect 2080 -30 2096 102
use CLKBUF1  CLKBUF1_57
timestamp 1732942776
transform 1 0 4 0 -1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_168
timestamp 1732942776
transform 1 0 76 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1732942776
transform 1 0 100 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1732942776
transform -1 0 100 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_162
timestamp 1732942776
transform -1 0 132 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1732942776
transform -1 0 292 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_2
timestamp 1732942776
transform 1 0 132 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1732942776
transform -1 0 188 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_102
timestamp 1732942776
transform 1 0 188 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_93
timestamp 1732942776
transform 1 0 292 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1732942776
transform -1 0 332 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_98
timestamp 1732942776
transform -1 0 348 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_28
timestamp 1732942776
transform -1 0 420 0 -1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_3
timestamp 1732942776
transform 1 0 332 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1732942776
transform -1 0 388 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_51
timestamp 1732942776
transform -1 0 420 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_59
timestamp 1732942776
transform 1 0 420 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_24
timestamp 1732942776
transform -1 0 564 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_35
timestamp 1732942776
transform 1 0 420 0 1 105
box -2 -3 74 103
use INVX8  INVX8_4
timestamp 1732942776
transform -1 0 532 0 1 105
box -2 -3 42 103
use FILL  FILL_0_0_0
timestamp 1732942776
transform 1 0 564 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1732942776
transform 1 0 572 0 -1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_34
timestamp 1732942776
transform 1 0 580 0 -1 105
box -2 -3 74 103
use FILL  FILL_1_0_0
timestamp 1732942776
transform -1 0 540 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1732942776
transform -1 0 548 0 1 105
box -2 -3 10 103
use BUFX4  BUFX4_54
timestamp 1732942776
transform -1 0 580 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_165
timestamp 1732942776
transform 1 0 580 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_26
timestamp 1732942776
transform 1 0 652 0 -1 105
box -2 -3 50 103
use INVX1  INVX1_26
timestamp 1732942776
transform -1 0 716 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_171
timestamp 1732942776
transform -1 0 636 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1732942776
transform 1 0 636 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1732942776
transform 1 0 716 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_175
timestamp 1732942776
transform 1 0 732 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1732942776
transform 1 0 780 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1732942776
transform -1 0 908 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_96
timestamp 1732942776
transform 1 0 908 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_29
timestamp 1732942776
transform 1 0 876 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_29
timestamp 1732942776
transform -1 0 940 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_101
timestamp 1732942776
transform -1 0 964 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1732942776
transform 1 0 964 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1732942776
transform -1 0 1036 0 1 105
box -2 -3 98 103
use FILL  FILL_0_1_0
timestamp 1732942776
transform 1 0 1060 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1732942776
transform 1 0 1068 0 -1 105
box -2 -3 10 103
use INVX1  INVX1_63
timestamp 1732942776
transform 1 0 1076 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_253
timestamp 1732942776
transform -1 0 1140 0 -1 105
box -2 -3 50 103
use BUFX4  BUFX4_49
timestamp 1732942776
transform -1 0 1068 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1732942776
transform 1 0 1068 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1732942776
transform 1 0 1076 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_7
timestamp 1732942776
transform 1 0 1084 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_7
timestamp 1732942776
transform 1 0 1140 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1732942776
transform -1 0 1196 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1732942776
transform -1 0 1292 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_8
timestamp 1732942776
transform -1 0 1140 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_222
timestamp 1732942776
transform -1 0 1188 0 1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_223
timestamp 1732942776
transform -1 0 1236 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_173
timestamp 1732942776
transform 1 0 1292 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_167
timestamp 1732942776
transform -1 0 1348 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1732942776
transform -1 0 1332 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1732942776
transform -1 0 1444 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_45
timestamp 1732942776
transform 1 0 1332 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_61
timestamp 1732942776
transform -1 0 1476 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_27
timestamp 1732942776
transform 1 0 1444 0 -1 105
box -2 -3 74 103
use BUFX4  BUFX4_21
timestamp 1732942776
transform -1 0 1548 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1732942776
transform 1 0 1476 0 1 105
box -2 -3 98 103
use FILL  FILL_0_2_0
timestamp 1732942776
transform 1 0 1548 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1732942776
transform 1 0 1556 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1732942776
transform 1 0 1564 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_2_0
timestamp 1732942776
transform 1 0 1572 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1732942776
transform 1 0 1580 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_15
timestamp 1732942776
transform 1 0 1588 0 1 105
box -2 -3 50 103
use INVX1  INVX1_65
timestamp 1732942776
transform 1 0 1660 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_255
timestamp 1732942776
transform -1 0 1724 0 -1 105
box -2 -3 50 103
use INVX1  INVX1_15
timestamp 1732942776
transform -1 0 1652 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_207
timestamp 1732942776
transform 1 0 1652 0 1 105
box -2 -3 50 103
use INVX8  INVX8_7
timestamp 1732942776
transform 1 0 1700 0 1 105
box -2 -3 42 103
use INVX8  INVX8_9
timestamp 1732942776
transform -1 0 1764 0 -1 105
box -2 -3 42 103
use MUX2X1  MUX2X1_31
timestamp 1732942776
transform 1 0 1764 0 -1 105
box -2 -3 50 103
use INVX1  INVX1_31
timestamp 1732942776
transform -1 0 1828 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_63
timestamp 1732942776
transform 1 0 1740 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1732942776
transform -1 0 1796 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_208
timestamp 1732942776
transform -1 0 1844 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1732942776
transform -1 0 1924 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1732942776
transform 1 0 1844 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1732942776
transform 1 0 1924 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1732942776
transform 1 0 2020 0 -1 105
box -2 -3 98 103
use BUFX4  BUFX4_20
timestamp 1732942776
transform 1 0 1940 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_1
timestamp 1732942776
transform -1 0 2044 0 1 105
box -2 -3 74 103
use FILL  FILL_0_3_0
timestamp 1732942776
transform 1 0 2116 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1732942776
transform 1 0 2124 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_93
timestamp 1732942776
transform 1 0 2044 0 1 105
box -2 -3 34 103
use FILL  FILL_1_3_0
timestamp 1732942776
transform -1 0 2084 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1732942776
transform -1 0 2092 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_94
timestamp 1732942776
transform -1 0 2124 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1732942776
transform -1 0 2220 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_55
timestamp 1732942776
transform 1 0 2132 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1732942776
transform -1 0 2188 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_16
timestamp 1732942776
transform -1 0 2260 0 -1 105
box -2 -3 74 103
use BUFX4  BUFX4_50
timestamp 1732942776
transform 1 0 2220 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_39
timestamp 1732942776
transform -1 0 2292 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1732942776
transform -1 0 2388 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_44
timestamp 1732942776
transform 1 0 2252 0 1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_7
timestamp 1732942776
transform 1 0 2276 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1732942776
transform -1 0 2420 0 1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_55
timestamp 1732942776
transform 1 0 2388 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_46
timestamp 1732942776
transform 1 0 2420 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_36
timestamp 1732942776
transform 1 0 2460 0 -1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_50
timestamp 1732942776
transform 1 0 2492 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1732942776
transform 1 0 2524 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1732942776
transform -1 0 2628 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_1
timestamp 1732942776
transform -1 0 2636 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1732942776
transform -1 0 2644 0 1 105
box -2 -3 98 103
use FILL  FILL_1_2
timestamp 1732942776
transform -1 0 2644 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_3
timestamp 1732942776
transform -1 0 2652 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_1
timestamp 1732942776
transform 1 0 2644 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1732942776
transform 1 0 4 0 -1 305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_47
timestamp 1732942776
transform 1 0 100 0 -1 305
box -2 -3 74 103
use MUX2X1  MUX2X1_103
timestamp 1732942776
transform 1 0 172 0 -1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_104
timestamp 1732942776
transform -1 0 268 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1732942776
transform 1 0 268 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1732942776
transform 1 0 364 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_5
timestamp 1732942776
transform -1 0 492 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1732942776
transform 1 0 492 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1732942776
transform 1 0 588 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1732942776
transform 1 0 596 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_5
timestamp 1732942776
transform 1 0 604 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1732942776
transform 1 0 636 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_61
timestamp 1732942776
transform 1 0 668 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1732942776
transform -1 0 724 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1732942776
transform -1 0 820 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_160
timestamp 1732942776
transform -1 0 868 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_13
timestamp 1732942776
transform 1 0 868 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_13
timestamp 1732942776
transform -1 0 932 0 -1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_159
timestamp 1732942776
transform 1 0 932 0 -1 305
box -2 -3 50 103
use BUFX4  BUFX4_52
timestamp 1732942776
transform -1 0 1012 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1732942776
transform 1 0 1012 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_98
timestamp 1732942776
transform -1 0 1068 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_1_0
timestamp 1732942776
transform -1 0 1076 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1732942776
transform -1 0 1084 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1732942776
transform -1 0 1180 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_224
timestamp 1732942776
transform 1 0 1180 0 -1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_21
timestamp 1732942776
transform 1 0 1228 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_21
timestamp 1732942776
transform -1 0 1292 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1732942776
transform -1 0 1388 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1732942776
transform -1 0 1484 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_119
timestamp 1732942776
transform 1 0 1484 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1732942776
transform -1 0 1540 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_2_0
timestamp 1732942776
transform 1 0 1540 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1732942776
transform 1 0 1548 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1732942776
transform 1 0 1556 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_117
timestamp 1732942776
transform 1 0 1652 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_116
timestamp 1732942776
transform -1 0 1708 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1732942776
transform -1 0 1804 0 -1 305
box -2 -3 98 103
use BUFX4  BUFX4_53
timestamp 1732942776
transform -1 0 1836 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_18
timestamp 1732942776
transform 1 0 1836 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_18
timestamp 1732942776
transform -1 0 1900 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1732942776
transform -1 0 1996 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_84
timestamp 1732942776
transform 1 0 1996 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1732942776
transform -1 0 2060 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_3_0
timestamp 1732942776
transform 1 0 2060 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1732942776
transform 1 0 2068 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1732942776
transform 1 0 2076 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_202
timestamp 1732942776
transform 1 0 2172 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1732942776
transform -1 0 2316 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_7
timestamp 1732942776
transform -1 0 2332 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1732942776
transform -1 0 2428 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_113
timestamp 1732942776
transform 1 0 2428 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_114
timestamp 1732942776
transform -1 0 2484 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_91
timestamp 1732942776
transform 1 0 2484 0 -1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1732942776
transform -1 0 2628 0 -1 305
box -2 -3 98 103
use FILL  FILL_3_1
timestamp 1732942776
transform -1 0 2636 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1732942776
transform -1 0 2644 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_3
timestamp 1732942776
transform -1 0 2652 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_26
timestamp 1732942776
transform 1 0 4 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1732942776
transform -1 0 60 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_94
timestamp 1732942776
transform 1 0 60 0 1 305
box -2 -3 50 103
use INVX1  INVX1_51
timestamp 1732942776
transform 1 0 108 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1732942776
transform -1 0 220 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_50
timestamp 1732942776
transform -1 0 268 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_125
timestamp 1732942776
transform 1 0 268 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_124
timestamp 1732942776
transform -1 0 324 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1732942776
transform 1 0 324 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_76
timestamp 1732942776
transform -1 0 380 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_169
timestamp 1732942776
transform 1 0 380 0 1 305
box -2 -3 50 103
use NOR2X1  NOR2X1_6
timestamp 1732942776
transform -1 0 452 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1732942776
transform 1 0 452 0 1 305
box -2 -3 98 103
use FILL  FILL_3_0_0
timestamp 1732942776
transform -1 0 556 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1732942776
transform -1 0 564 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_174
timestamp 1732942776
transform -1 0 612 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_5
timestamp 1732942776
transform 1 0 612 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_176
timestamp 1732942776
transform 1 0 636 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_58
timestamp 1732942776
transform 1 0 684 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1732942776
transform -1 0 740 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1732942776
transform 1 0 740 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_88
timestamp 1732942776
transform 1 0 836 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_161
timestamp 1732942776
transform -1 0 932 0 1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1732942776
transform 1 0 932 0 1 305
box -2 -3 98 103
use INVX1  INVX1_5
timestamp 1732942776
transform 1 0 1028 0 1 305
box -2 -3 18 103
use FILL  FILL_3_1_0
timestamp 1732942776
transform -1 0 1052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1732942776
transform -1 0 1060 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_5
timestamp 1732942776
transform -1 0 1108 0 1 305
box -2 -3 50 103
use CLKBUF1  CLKBUF1_13
timestamp 1732942776
transform -1 0 1180 0 1 305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_2
timestamp 1732942776
transform -1 0 1252 0 1 305
box -2 -3 74 103
use MUX2X1  MUX2X1_157
timestamp 1732942776
transform 1 0 1252 0 1 305
box -2 -3 50 103
use BUFX4  BUFX4_46
timestamp 1732942776
transform 1 0 1300 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_156
timestamp 1732942776
transform 1 0 1332 0 1 305
box -2 -3 50 103
use NOR2X1  NOR2X1_26
timestamp 1732942776
transform 1 0 1380 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1732942776
transform -1 0 1436 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1732942776
transform 1 0 1436 0 1 305
box -2 -3 98 103
use OR2X2  OR2X2_1
timestamp 1732942776
transform 1 0 1532 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1732942776
transform 1 0 1564 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1732942776
transform 1 0 1572 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1732942776
transform 1 0 1580 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_209
timestamp 1732942776
transform 1 0 1676 0 1 305
box -2 -3 50 103
use NOR2X1  NOR2X1_28
timestamp 1732942776
transform 1 0 1724 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1732942776
transform -1 0 1780 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1732942776
transform 1 0 1780 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_23
timestamp 1732942776
transform 1 0 1876 0 1 305
box -2 -3 50 103
use INVX1  INVX1_23
timestamp 1732942776
transform -1 0 1940 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_85
timestamp 1732942776
transform 1 0 1940 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_205
timestamp 1732942776
transform -1 0 2036 0 1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_10
timestamp 1732942776
transform 1 0 2036 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1732942776
transform -1 0 2092 0 1 305
box -2 -3 26 103
use FILL  FILL_3_3_0
timestamp 1732942776
transform -1 0 2100 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1732942776
transform -1 0 2108 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_204
timestamp 1732942776
transform -1 0 2156 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_90
timestamp 1732942776
transform -1 0 2204 0 1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_15
timestamp 1732942776
transform 1 0 2204 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1732942776
transform 1 0 2236 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_82
timestamp 1732942776
transform 1 0 2260 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_39
timestamp 1732942776
transform 1 0 2308 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_34
timestamp 1732942776
transform -1 0 2364 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1732942776
transform -1 0 2460 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_42
timestamp 1732942776
transform 1 0 2460 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1732942776
transform -1 0 2516 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1732942776
transform -1 0 2612 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_26
timestamp 1732942776
transform 1 0 2612 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1732942776
transform 1 0 2644 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1732942776
transform 1 0 4 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_34
timestamp 1732942776
transform 1 0 100 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_34
timestamp 1732942776
transform -1 0 164 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1732942776
transform -1 0 260 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_42
timestamp 1732942776
transform 1 0 260 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_42
timestamp 1732942776
transform -1 0 324 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1732942776
transform -1 0 420 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1732942776
transform -1 0 516 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_73
timestamp 1732942776
transform 1 0 516 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1732942776
transform -1 0 548 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1732942776
transform -1 0 556 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_66
timestamp 1732942776
transform -1 0 588 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1732942776
transform -1 0 620 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1732942776
transform -1 0 716 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1732942776
transform -1 0 812 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_10
timestamp 1732942776
transform 1 0 812 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1732942776
transform -1 0 868 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1732942776
transform 1 0 868 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_21
timestamp 1732942776
transform 1 0 964 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_18
timestamp 1732942776
transform -1 0 1020 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1732942776
transform -1 0 1028 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1732942776
transform -1 0 1036 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1732942776
transform -1 0 1132 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1732942776
transform 1 0 1132 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_90
timestamp 1732942776
transform -1 0 1260 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1732942776
transform -1 0 1292 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1732942776
transform 1 0 1292 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_88
timestamp 1732942776
transform 1 0 1388 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1732942776
transform -1 0 1452 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_20
timestamp 1732942776
transform 1 0 1452 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_20
timestamp 1732942776
transform -1 0 1516 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_14
timestamp 1732942776
transform 1 0 1516 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_13
timestamp 1732942776
transform -1 0 1572 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1732942776
transform -1 0 1580 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1732942776
transform -1 0 1588 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1732942776
transform -1 0 1684 0 -1 505
box -2 -3 98 103
use BUFX4  BUFX4_45
timestamp 1732942776
transform 1 0 1684 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1732942776
transform 1 0 1716 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1732942776
transform -1 0 1772 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1732942776
transform -1 0 1868 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1732942776
transform 1 0 1868 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1732942776
transform 1 0 1964 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_23
timestamp 1732942776
transform 1 0 2060 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_3_0
timestamp 1732942776
transform -1 0 2092 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1732942776
transform -1 0 2100 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_18
timestamp 1732942776
transform -1 0 2132 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_206
timestamp 1732942776
transform 1 0 2132 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_52
timestamp 1732942776
transform -1 0 2204 0 -1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_210
timestamp 1732942776
transform 1 0 2204 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_92
timestamp 1732942776
transform 1 0 2252 0 -1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_79
timestamp 1732942776
transform 1 0 2300 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1732942776
transform -1 0 2356 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_36
timestamp 1732942776
transform 1 0 2356 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1732942776
transform -1 0 2476 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_16
timestamp 1732942776
transform -1 0 2500 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1732942776
transform 1 0 2500 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_34
timestamp 1732942776
transform 1 0 2596 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_29
timestamp 1732942776
transform 1 0 2620 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_48
timestamp 1732942776
transform 1 0 4 0 1 505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_25
timestamp 1732942776
transform 1 0 76 0 1 505
box -2 -3 74 103
use MUX2X1  MUX2X1_93
timestamp 1732942776
transform 1 0 148 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1732942776
transform 1 0 196 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_37
timestamp 1732942776
transform 1 0 292 0 1 505
box -2 -3 50 103
use INVX1  INVX1_37
timestamp 1732942776
transform -1 0 356 0 1 505
box -2 -3 18 103
use INVX1  INVX1_54
timestamp 1732942776
transform 1 0 356 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_53
timestamp 1732942776
transform -1 0 420 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_165
timestamp 1732942776
transform 1 0 420 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1732942776
transform 1 0 468 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1732942776
transform 1 0 564 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1732942776
transform 1 0 572 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_50
timestamp 1732942776
transform 1 0 580 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_54
timestamp 1732942776
transform 1 0 612 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_168
timestamp 1732942776
transform -1 0 684 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_109
timestamp 1732942776
transform 1 0 684 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_107
timestamp 1732942776
transform 1 0 716 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1732942776
transform -1 0 836 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_154
timestamp 1732942776
transform 1 0 836 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1732942776
transform 1 0 868 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_100
timestamp 1732942776
transform 1 0 892 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_99
timestamp 1732942776
transform 1 0 940 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1732942776
transform 1 0 988 0 1 505
box -2 -3 98 103
use FILL  FILL_5_1_0
timestamp 1732942776
transform -1 0 1092 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1732942776
transform -1 0 1100 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_15
timestamp 1732942776
transform -1 0 1132 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1732942776
transform 1 0 1132 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_55
timestamp 1732942776
transform -1 0 1188 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1732942776
transform 1 0 1188 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_163
timestamp 1732942776
transform 1 0 1284 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_157
timestamp 1732942776
transform -1 0 1340 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_158
timestamp 1732942776
transform -1 0 1388 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_172
timestamp 1732942776
transform 1 0 1388 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_133
timestamp 1732942776
transform 1 0 1436 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1732942776
transform 1 0 1484 0 1 505
box -2 -3 98 103
use FILL  FILL_5_2_0
timestamp 1732942776
transform 1 0 1580 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1732942776
transform 1 0 1588 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_37
timestamp 1732942776
transform 1 0 1596 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1732942776
transform -1 0 1652 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_154
timestamp 1732942776
transform -1 0 1700 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_171
timestamp 1732942776
transform -1 0 1748 0 1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_65
timestamp 1732942776
transform 1 0 1748 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_58
timestamp 1732942776
transform -1 0 1804 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1732942776
transform -1 0 1900 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_2
timestamp 1732942776
transform 1 0 1900 0 1 505
box -2 -3 50 103
use INVX1  INVX1_2
timestamp 1732942776
transform -1 0 1964 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_84
timestamp 1732942776
transform 1 0 1964 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_86
timestamp 1732942776
transform 1 0 2012 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_47
timestamp 1732942776
transform 1 0 2060 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1732942776
transform 1 0 2092 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1732942776
transform 1 0 2100 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1732942776
transform 1 0 2108 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_201
timestamp 1732942776
transform -1 0 2252 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_212
timestamp 1732942776
transform 1 0 2252 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_211
timestamp 1732942776
transform 1 0 2300 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_31
timestamp 1732942776
transform 1 0 2348 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1732942776
transform 1 0 2380 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_74
timestamp 1732942776
transform 1 0 2476 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1732942776
transform -1 0 2532 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_163
timestamp 1732942776
transform 1 0 2532 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_50
timestamp 1732942776
transform 1 0 2580 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_45
timestamp 1732942776
transform 1 0 2604 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1732942776
transform 1 0 2636 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1732942776
transform 1 0 2644 0 1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_62
timestamp 1732942776
transform -1 0 76 0 -1 705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_14
timestamp 1732942776
transform 1 0 76 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1732942776
transform 1 0 148 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_47
timestamp 1732942776
transform 1 0 244 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1732942776
transform -1 0 300 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_95
timestamp 1732942776
transform -1 0 348 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_250
timestamp 1732942776
transform 1 0 348 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_60
timestamp 1732942776
transform -1 0 412 0 -1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_166
timestamp 1732942776
transform -1 0 460 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_96
timestamp 1732942776
transform -1 0 508 0 -1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_7
timestamp 1732942776
transform 1 0 508 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_0_0
timestamp 1732942776
transform 1 0 548 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1732942776
transform 1 0 556 0 -1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_98
timestamp 1732942776
transform 1 0 564 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_97
timestamp 1732942776
transform -1 0 660 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_170
timestamp 1732942776
transform 1 0 660 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_167
timestamp 1732942776
transform 1 0 708 0 -1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_19
timestamp 1732942776
transform 1 0 756 0 -1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1732942776
transform 1 0 796 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_10
timestamp 1732942776
transform 1 0 892 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_10
timestamp 1732942776
transform -1 0 956 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_8
timestamp 1732942776
transform -1 0 996 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_101
timestamp 1732942776
transform -1 0 1044 0 -1 705
box -2 -3 50 103
use FILL  FILL_6_1_0
timestamp 1732942776
transform 1 0 1044 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1732942776
transform 1 0 1052 0 -1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_87
timestamp 1732942776
transform 1 0 1060 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_16
timestamp 1732942776
transform -1 0 1132 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_89
timestamp 1732942776
transform 1 0 1132 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_220
timestamp 1732942776
transform 1 0 1180 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_142
timestamp 1732942776
transform 1 0 1228 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_20
timestamp 1732942776
transform -1 0 1292 0 -1 705
box -2 -3 42 103
use AOI22X1  AOI22X1_28
timestamp 1732942776
transform -1 0 1332 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_221
timestamp 1732942776
transform -1 0 1380 0 -1 705
box -2 -3 50 103
use AOI21X1  AOI21X1_20
timestamp 1732942776
transform 1 0 1380 0 -1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_58
timestamp 1732942776
transform -1 0 1484 0 -1 705
box -2 -3 74 103
use OAI21X1  OAI21X1_28
timestamp 1732942776
transform 1 0 1484 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_173
timestamp 1732942776
transform -1 0 1564 0 -1 705
box -2 -3 50 103
use FILL  FILL_6_2_0
timestamp 1732942776
transform -1 0 1572 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1732942776
transform -1 0 1580 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_33
timestamp 1732942776
transform -1 0 1604 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_17
timestamp 1732942776
transform -1 0 1644 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_141
timestamp 1732942776
transform 1 0 1644 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_18
timestamp 1732942776
transform 1 0 1668 0 -1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1732942776
transform -1 0 1804 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_26
timestamp 1732942776
transform 1 0 1804 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_23
timestamp 1732942776
transform -1 0 1860 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1732942776
transform -1 0 1892 0 -1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_15
timestamp 1732942776
transform 1 0 1892 0 -1 705
box -2 -3 74 103
use AOI22X1  AOI22X1_6
timestamp 1732942776
transform 1 0 1964 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_132
timestamp 1732942776
transform -1 0 2028 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_5
timestamp 1732942776
transform -1 0 2068 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_3_0
timestamp 1732942776
transform 1 0 2068 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1732942776
transform 1 0 2076 0 -1 705
box -2 -3 10 103
use AOI22X1  AOI22X1_26
timestamp 1732942776
transform 1 0 2084 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_147
timestamp 1732942776
transform -1 0 2148 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_25
timestamp 1732942776
transform -1 0 2188 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_203
timestamp 1732942776
transform -1 0 2236 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_83
timestamp 1732942776
transform 1 0 2236 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1732942776
transform 1 0 2284 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_81
timestamp 1732942776
transform -1 0 2428 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_164
timestamp 1732942776
transform 1 0 2428 0 -1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_162
timestamp 1732942776
transform 1 0 2476 0 -1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_53
timestamp 1732942776
transform -1 0 2556 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1732942776
transform -1 0 2652 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1732942776
transform 1 0 4 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_104
timestamp 1732942776
transform 1 0 100 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_106
timestamp 1732942776
transform -1 0 156 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1732942776
transform 1 0 156 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_36
timestamp 1732942776
transform -1 0 276 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_29
timestamp 1732942776
transform -1 0 308 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1732942776
transform 1 0 308 0 1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_45
timestamp 1732942776
transform 1 0 404 0 1 705
box -2 -3 50 103
use INVX1  INVX1_45
timestamp 1732942776
transform -1 0 468 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1732942776
transform -1 0 564 0 1 705
box -2 -3 98 103
use FILL  FILL_7_0_0
timestamp 1732942776
transform -1 0 572 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1732942776
transform -1 0 580 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1732942776
transform -1 0 676 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_121
timestamp 1732942776
transform 1 0 676 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_122
timestamp 1732942776
transform -1 0 732 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1732942776
transform 1 0 732 0 1 705
box -2 -3 50 103
use INVX1  INVX1_47
timestamp 1732942776
transform -1 0 796 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1732942776
transform -1 0 892 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_101
timestamp 1732942776
transform 1 0 892 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1732942776
transform -1 0 948 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_133
timestamp 1732942776
transform 1 0 948 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_19
timestamp 1732942776
transform -1 0 1004 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1732942776
transform 1 0 1004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1732942776
transform 1 0 1036 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1732942776
transform -1 0 1076 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1732942776
transform -1 0 1084 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_165
timestamp 1732942776
transform -1 0 1108 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1732942776
transform 1 0 1108 0 1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_8
timestamp 1732942776
transform -1 0 1276 0 1 705
box -2 -3 74 103
use NAND2X1  NAND2X1_148
timestamp 1732942776
transform 1 0 1276 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1732942776
transform 1 0 1300 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_25
timestamp 1732942776
transform 1 0 1396 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_134
timestamp 1732942776
transform 1 0 1420 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1732942776
transform 1 0 1468 0 1 705
box -2 -3 98 103
use FILL  FILL_7_2_0
timestamp 1732942776
transform 1 0 1564 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1732942776
transform 1 0 1572 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_156
timestamp 1732942776
transform 1 0 1580 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1732942776
transform 1 0 1604 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_133
timestamp 1732942776
transform -1 0 1668 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_155
timestamp 1732942776
transform -1 0 1716 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_219
timestamp 1732942776
transform 1 0 1716 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1732942776
transform -1 0 1860 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_67
timestamp 1732942776
transform 1 0 1860 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_60
timestamp 1732942776
transform -1 0 1916 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_153
timestamp 1732942776
transform -1 0 1964 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_130
timestamp 1732942776
transform -1 0 1996 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_68
timestamp 1732942776
transform -1 0 2068 0 1 705
box -2 -3 74 103
use FILL  FILL_7_3_0
timestamp 1732942776
transform -1 0 2076 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1732942776
transform -1 0 2084 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_135
timestamp 1732942776
transform -1 0 2116 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1732942776
transform 1 0 2116 0 1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_150
timestamp 1732942776
transform -1 0 2244 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1732942776
transform 1 0 2244 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_140
timestamp 1732942776
transform 1 0 2268 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_77
timestamp 1732942776
transform -1 0 2332 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1732942776
transform -1 0 2428 0 1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_13
timestamp 1732942776
transform 1 0 2428 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1732942776
transform -1 0 2556 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1732942776
transform -1 0 2652 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1732942776
transform 1 0 4 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_35
timestamp 1732942776
transform 1 0 100 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_35
timestamp 1732942776
transform -1 0 164 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1732942776
transform -1 0 260 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_99
timestamp 1732942776
transform -1 0 292 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1732942776
transform 1 0 292 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_52
timestamp 1732942776
transform -1 0 420 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_216
timestamp 1732942776
transform -1 0 468 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_218
timestamp 1732942776
transform 1 0 468 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_217
timestamp 1732942776
transform -1 0 564 0 -1 905
box -2 -3 50 103
use FILL  FILL_8_0_0
timestamp 1732942776
transform 1 0 564 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1732942776
transform 1 0 572 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_126
timestamp 1732942776
transform 1 0 580 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1732942776
transform -1 0 700 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_78
timestamp 1732942776
transform -1 0 724 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_71
timestamp 1732942776
transform -1 0 756 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_27
timestamp 1732942776
transform -1 0 796 0 -1 905
box -2 -3 42 103
use MUX2X1  MUX2X1_213
timestamp 1732942776
transform -1 0 844 0 -1 905
box -2 -3 50 103
use CLKBUF1  CLKBUF1_66
timestamp 1732942776
transform 1 0 844 0 -1 905
box -2 -3 74 103
use INVX1  INVX1_39
timestamp 1732942776
transform 1 0 916 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1732942776
transform -1 0 1028 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_39
timestamp 1732942776
transform 1 0 1028 0 -1 905
box -2 -3 50 103
use FILL  FILL_8_1_0
timestamp 1732942776
transform 1 0 1076 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1732942776
transform 1 0 1084 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1732942776
transform 1 0 1092 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_28
timestamp 1732942776
transform 1 0 1188 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_28
timestamp 1732942776
transform -1 0 1252 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1732942776
transform 1 0 1252 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_4
timestamp 1732942776
transform 1 0 1348 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_4
timestamp 1732942776
transform -1 0 1412 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_132
timestamp 1732942776
transform -1 0 1460 0 -1 905
box -2 -3 50 103
use AND2X2  AND2X2_4
timestamp 1732942776
transform 1 0 1460 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_5
timestamp 1732942776
transform 1 0 1492 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1732942776
transform -1 0 1604 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_2_0
timestamp 1732942776
transform -1 0 1612 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1732942776
transform -1 0 1620 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_20
timestamp 1732942776
transform -1 0 1652 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_139
timestamp 1732942776
transform -1 0 1700 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1732942776
transform 1 0 1700 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_143
timestamp 1732942776
transform -1 0 1828 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_144
timestamp 1732942776
transform -1 0 1860 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1732942776
transform 1 0 1860 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1732942776
transform -1 0 1988 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_26
timestamp 1732942776
transform -1 0 2060 0 -1 905
box -2 -3 74 103
use INVX8  INVX8_11
timestamp 1732942776
transform 1 0 2060 0 -1 905
box -2 -3 42 103
use FILL  FILL_8_3_0
timestamp 1732942776
transform -1 0 2108 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1732942776
transform -1 0 2116 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_145
timestamp 1732942776
transform -1 0 2148 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_146
timestamp 1732942776
transform -1 0 2180 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1732942776
transform 1 0 2180 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1732942776
transform -1 0 2244 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1732942776
transform -1 0 2276 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_139
timestamp 1732942776
transform 1 0 2276 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1732942776
transform 1 0 2308 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1732942776
transform -1 0 2476 0 -1 905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_53
timestamp 1732942776
transform 1 0 2476 0 -1 905
box -2 -3 74 103
use AOI21X1  AOI21X1_44
timestamp 1732942776
transform -1 0 2580 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_21
timestamp 1732942776
transform 1 0 2580 0 -1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1732942776
transform 1 0 4 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_169
timestamp 1732942776
transform 1 0 100 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_163
timestamp 1732942776
transform -1 0 156 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_127
timestamp 1732942776
transform 1 0 156 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_94
timestamp 1732942776
transform 1 0 204 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1732942776
transform 1 0 228 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_75
timestamp 1732942776
transform 1 0 324 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_68
timestamp 1732942776
transform -1 0 380 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_56
timestamp 1732942776
transform 1 0 380 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_117
timestamp 1732942776
transform -1 0 452 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_111
timestamp 1732942776
transform 1 0 452 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_109
timestamp 1732942776
transform -1 0 508 0 1 905
box -2 -3 26 103
use FILL  FILL_9_0_0
timestamp 1732942776
transform -1 0 516 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1732942776
transform -1 0 524 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1732942776
transform -1 0 620 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_127
timestamp 1732942776
transform -1 0 652 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1732942776
transform -1 0 748 0 1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_39
timestamp 1732942776
transform -1 0 820 0 1 905
box -2 -3 74 103
use MUX2X1  MUX2X1_215
timestamp 1732942776
transform 1 0 820 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_214
timestamp 1732942776
transform -1 0 916 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_55
timestamp 1732942776
transform 1 0 916 0 1 905
box -2 -3 50 103
use INVX1  INVX1_56
timestamp 1732942776
transform -1 0 980 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1732942776
transform -1 0 1076 0 1 905
box -2 -3 98 103
use FILL  FILL_9_1_0
timestamp 1732942776
transform 1 0 1076 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1732942776
transform 1 0 1084 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_12
timestamp 1732942776
transform 1 0 1092 0 1 905
box -2 -3 50 103
use INVX1  INVX1_12
timestamp 1732942776
transform -1 0 1156 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1732942776
transform 1 0 1156 0 1 905
box -2 -3 98 103
use INVX1  INVX1_49
timestamp 1732942776
transform 1 0 1252 0 1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_31
timestamp 1732942776
transform 1 0 1268 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_136
timestamp 1732942776
transform 1 0 1292 0 1 905
box -2 -3 50 103
use BUFX4  BUFX4_27
timestamp 1732942776
transform 1 0 1340 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1732942776
transform 1 0 1372 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1732942776
transform 1 0 1404 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_64
timestamp 1732942776
transform 1 0 1500 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_147
timestamp 1732942776
transform -1 0 1572 0 1 905
box -2 -3 50 103
use FILL  FILL_9_2_0
timestamp 1732942776
transform 1 0 1572 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1732942776
transform 1 0 1580 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_23
timestamp 1732942776
transform 1 0 1588 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1732942776
transform 1 0 1612 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_49
timestamp 1732942776
transform 1 0 1708 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1732942776
transform -1 0 1764 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_129
timestamp 1732942776
transform -1 0 1812 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_140
timestamp 1732942776
transform -1 0 1860 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_138
timestamp 1732942776
transform -1 0 1908 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_58
timestamp 1732942776
transform 1 0 1908 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_32
timestamp 1732942776
transform -1 0 1964 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1732942776
transform -1 0 1996 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1732942776
transform -1 0 2028 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1732942776
transform 1 0 2028 0 1 905
box -2 -3 34 103
use FILL  FILL_9_3_0
timestamp 1732942776
transform -1 0 2068 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1732942776
transform -1 0 2076 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1732942776
transform -1 0 2172 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_140
timestamp 1732942776
transform 1 0 2172 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_266
timestamp 1732942776
transform 1 0 2196 0 1 905
box -2 -3 98 103
use BUFX4  BUFX4_37
timestamp 1732942776
transform -1 0 2324 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1732942776
transform -1 0 2356 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1732942776
transform 1 0 2356 0 1 905
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1732942776
transform -1 0 2396 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1732942776
transform -1 0 2492 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_59
timestamp 1732942776
transform 1 0 2492 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1732942776
transform 1 0 2516 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_5
timestamp 1732942776
transform 1 0 2548 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_41
timestamp 1732942776
transform 1 0 2572 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_146
timestamp 1732942776
transform 1 0 2596 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1732942776
transform 1 0 2620 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1732942776
transform 1 0 2644 0 1 905
box -2 -3 10 103
use INVX8  INVX8_6
timestamp 1732942776
transform 1 0 4 0 -1 1105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1732942776
transform 1 0 44 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_27
timestamp 1732942776
transform 1 0 140 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_34
timestamp 1732942776
transform -1 0 196 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1732942776
transform 1 0 196 0 -1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_118
timestamp 1732942776
transform 1 0 292 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_52
timestamp 1732942776
transform 1 0 340 0 -1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_51
timestamp 1732942776
transform -1 0 404 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_119
timestamp 1732942776
transform -1 0 452 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1732942776
transform -1 0 548 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_0_0
timestamp 1732942776
transform -1 0 556 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1732942776
transform -1 0 564 0 -1 1105
box -2 -3 10 103
use BUFX4  BUFX4_26
timestamp 1732942776
transform -1 0 596 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1732942776
transform 1 0 596 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_104
timestamp 1732942776
transform 1 0 692 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_99
timestamp 1732942776
transform -1 0 748 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1732942776
transform 1 0 748 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_5
timestamp 1732942776
transform 1 0 844 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1732942776
transform -1 0 900 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1732942776
transform 1 0 900 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_28
timestamp 1732942776
transform -1 0 1028 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1732942776
transform 1 0 1028 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1732942776
transform 1 0 1060 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1732942776
transform 1 0 1068 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_38
timestamp 1732942776
transform 1 0 1076 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_252
timestamp 1732942776
transform 1 0 1100 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_62
timestamp 1732942776
transform -1 0 1164 0 -1 1105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_38
timestamp 1732942776
transform -1 0 1236 0 -1 1105
box -2 -3 74 103
use BUFX4  BUFX4_24
timestamp 1732942776
transform -1 0 1268 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_67
timestamp 1732942776
transform -1 0 1292 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_135
timestamp 1732942776
transform 1 0 1292 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_137
timestamp 1732942776
transform 1 0 1340 0 -1 1105
box -2 -3 50 103
use INVX8  INVX8_2
timestamp 1732942776
transform -1 0 1428 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_49
timestamp 1732942776
transform 1 0 1428 0 -1 1105
box -2 -3 26 103
use OR2X2  OR2X2_2
timestamp 1732942776
transform -1 0 1484 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1732942776
transform -1 0 1508 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_25
timestamp 1732942776
transform 1 0 1508 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_131
timestamp 1732942776
transform -1 0 1588 0 -1 1105
box -2 -3 50 103
use FILL  FILL_10_2_0
timestamp 1732942776
transform 1 0 1588 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1732942776
transform 1 0 1596 0 -1 1105
box -2 -3 10 103
use AOI22X1  AOI22X1_13
timestamp 1732942776
transform 1 0 1604 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_138
timestamp 1732942776
transform 1 0 1644 0 -1 1105
box -2 -3 26 103
use AOI22X1  AOI22X1_14
timestamp 1732942776
transform 1 0 1668 0 -1 1105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1732942776
transform -1 0 1804 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_86
timestamp 1732942776
transform 1 0 1804 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_76
timestamp 1732942776
transform -1 0 1860 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1732942776
transform 1 0 1860 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1732942776
transform -1 0 1916 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1732942776
transform -1 0 2012 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_33
timestamp 1732942776
transform 1 0 2012 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1732942776
transform 1 0 2044 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_47
timestamp 1732942776
transform 1 0 2068 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_3_0
timestamp 1732942776
transform 1 0 2092 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1732942776
transform 1 0 2100 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_10
timestamp 1732942776
transform 1 0 2108 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1732942776
transform -1 0 2228 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_157
timestamp 1732942776
transform -1 0 2252 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_48
timestamp 1732942776
transform 1 0 2252 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_152
timestamp 1732942776
transform 1 0 2276 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_158
timestamp 1732942776
transform 1 0 2300 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1732942776
transform -1 0 2420 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_35
timestamp 1732942776
transform 1 0 2420 0 -1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_6
timestamp 1732942776
transform -1 0 2524 0 -1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_268
timestamp 1732942776
transform 1 0 2524 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_42
timestamp 1732942776
transform 1 0 2620 0 -1 1105
box -2 -3 26 103
use FILL  FILL_11_1
timestamp 1732942776
transform -1 0 2652 0 -1 1105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_60
timestamp 1732942776
transform 1 0 4 0 1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1732942776
transform 1 0 76 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_107
timestamp 1732942776
transform 1 0 172 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_105
timestamp 1732942776
transform -1 0 228 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_120
timestamp 1732942776
transform 1 0 228 0 1 1105
box -2 -3 50 103
use AOI21X1  AOI21X1_48
timestamp 1732942776
transform 1 0 276 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1732942776
transform 1 0 308 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_8
timestamp 1732942776
transform -1 0 364 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_43
timestamp 1732942776
transform 1 0 364 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_43
timestamp 1732942776
transform -1 0 428 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1732942776
transform -1 0 524 0 1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_49
timestamp 1732942776
transform 1 0 524 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1732942776
transform -1 0 564 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1732942776
transform -1 0 572 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_53
timestamp 1732942776
transform -1 0 596 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1732942776
transform 1 0 596 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_168
timestamp 1732942776
transform 1 0 692 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_174
timestamp 1732942776
transform 1 0 724 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_247
timestamp 1732942776
transform 1 0 748 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_150
timestamp 1732942776
transform 1 0 796 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_100
timestamp 1732942776
transform 1 0 844 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_95
timestamp 1732942776
transform -1 0 900 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_152
timestamp 1732942776
transform 1 0 900 0 1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1732942776
transform -1 0 1044 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_1_0
timestamp 1732942776
transform 1 0 1044 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1732942776
transform 1 0 1052 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1732942776
transform 1 0 1060 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1732942776
transform 1 0 1156 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_60
timestamp 1732942776
transform 1 0 1252 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_156
timestamp 1732942776
transform 1 0 1284 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_162
timestamp 1732942776
transform -1 0 1340 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1732942776
transform 1 0 1340 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_21
timestamp 1732942776
transform 1 0 1436 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_60
timestamp 1732942776
transform 1 0 1460 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_59
timestamp 1732942776
transform -1 0 1508 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_148
timestamp 1732942776
transform 1 0 1508 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_13
timestamp 1732942776
transform 1 0 1556 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_2_0
timestamp 1732942776
transform -1 0 1588 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1732942776
transform -1 0 1596 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_12
timestamp 1732942776
transform -1 0 1628 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1732942776
transform -1 0 1724 0 1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_5
timestamp 1732942776
transform -1 0 1796 0 1 1105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_42
timestamp 1732942776
transform 1 0 1796 0 1 1105
box -2 -3 74 103
use INVX2  INVX2_4
timestamp 1732942776
transform 1 0 1868 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1732942776
transform -1 0 1980 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_30
timestamp 1732942776
transform -1 0 2012 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_36
timestamp 1732942776
transform -1 0 2044 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_108
timestamp 1732942776
transform -1 0 2092 0 1 1105
box -2 -3 50 103
use FILL  FILL_11_3_0
timestamp 1732942776
transform 1 0 2092 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1732942776
transform 1 0 2100 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_154
timestamp 1732942776
transform 1 0 2108 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1732942776
transform 1 0 2132 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1732942776
transform -1 0 2188 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1732942776
transform 1 0 2188 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_40
timestamp 1732942776
transform 1 0 2284 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_35
timestamp 1732942776
transform -1 0 2340 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_33
timestamp 1732942776
transform 1 0 2340 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1732942776
transform 1 0 2372 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_40
timestamp 1732942776
transform 1 0 2404 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_40
timestamp 1732942776
transform 1 0 2428 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1732942776
transform -1 0 2556 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_267
timestamp 1732942776
transform 1 0 2556 0 1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_41
timestamp 1732942776
transform -1 0 76 0 -1 1305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1732942776
transform 1 0 76 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_122
timestamp 1732942776
transform 1 0 172 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_123
timestamp 1732942776
transform -1 0 228 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_122
timestamp 1732942776
transform -1 0 276 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1732942776
transform 1 0 276 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_124
timestamp 1732942776
transform 1 0 372 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1732942776
transform -1 0 428 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_11
timestamp 1732942776
transform 1 0 428 0 -1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_145
timestamp 1732942776
transform -1 0 516 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_146
timestamp 1732942776
transform -1 0 564 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_0_0
timestamp 1732942776
transform -1 0 572 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1732942776
transform -1 0 580 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_106
timestamp 1732942776
transform -1 0 604 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_144
timestamp 1732942776
transform 1 0 604 0 -1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_15
timestamp 1732942776
transform -1 0 692 0 -1 1305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1732942776
transform 1 0 692 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_4
timestamp 1732942776
transform 1 0 788 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1732942776
transform 1 0 820 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_170
timestamp 1732942776
transform 1 0 844 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_151
timestamp 1732942776
transform 1 0 868 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1732942776
transform -1 0 1012 0 -1 1305
box -2 -3 98 103
use BUFX4  BUFX4_11
timestamp 1732942776
transform 1 0 1012 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_136
timestamp 1732942776
transform 1 0 1044 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_1_0
timestamp 1732942776
transform 1 0 1068 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1732942776
transform 1 0 1076 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_8
timestamp 1732942776
transform 1 0 1084 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1732942776
transform 1 0 1116 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1732942776
transform -1 0 1180 0 -1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_1
timestamp 1732942776
transform -1 0 1212 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_19
timestamp 1732942776
transform 1 0 1212 0 -1 1305
box -2 -3 74 103
use NAND3X1  NAND3X1_3
timestamp 1732942776
transform 1 0 1284 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1732942776
transform 1 0 1316 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_116
timestamp 1732942776
transform 1 0 1412 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_115
timestamp 1732942776
transform -1 0 1468 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_130
timestamp 1732942776
transform 1 0 1468 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_149
timestamp 1732942776
transform -1 0 1564 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_2_0
timestamp 1732942776
transform 1 0 1564 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1732942776
transform 1 0 1572 0 -1 1305
box -2 -3 10 103
use INVX2  INVX2_7
timestamp 1732942776
transform 1 0 1580 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_28
timestamp 1732942776
transform 1 0 1596 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1732942776
transform -1 0 1652 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_46
timestamp 1732942776
transform 1 0 1652 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_132
timestamp 1732942776
transform 1 0 1676 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1732942776
transform -1 0 1740 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_15
timestamp 1732942776
transform 1 0 1740 0 -1 1305
box -2 -3 34 103
use INVX4  INVX4_1
timestamp 1732942776
transform -1 0 1796 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_41
timestamp 1732942776
transform 1 0 1796 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_137
timestamp 1732942776
transform 1 0 1828 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_265
timestamp 1732942776
transform 1 0 1852 0 -1 1305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_18
timestamp 1732942776
transform -1 0 2020 0 -1 1305
box -2 -3 74 103
use BUFX2  BUFX2_4
timestamp 1732942776
transform 1 0 2020 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_131
timestamp 1732942776
transform 1 0 2044 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1732942776
transform 1 0 2076 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1732942776
transform 1 0 2084 0 -1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_3
timestamp 1732942776
transform 1 0 2092 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_3
timestamp 1732942776
transform -1 0 2156 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1732942776
transform 1 0 2156 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_106
timestamp 1732942776
transform 1 0 2252 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_59
timestamp 1732942776
transform 1 0 2300 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1732942776
transform -1 0 2412 0 -1 1305
box -2 -3 98 103
use BUFX4  BUFX4_34
timestamp 1732942776
transform -1 0 2444 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1732942776
transform 1 0 2444 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1732942776
transform -1 0 2500 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1732942776
transform -1 0 2596 0 -1 1305
box -2 -3 98 103
use BUFX2  BUFX2_3
timestamp 1732942776
transform 1 0 2596 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_10
timestamp 1732942776
transform 1 0 2620 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1732942776
transform 1 0 4 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_4
timestamp 1732942776
transform 1 0 100 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1732942776
transform -1 0 156 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_121
timestamp 1732942776
transform -1 0 204 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_128
timestamp 1732942776
transform -1 0 252 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_9
timestamp 1732942776
transform -1 0 284 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_44
timestamp 1732942776
transform -1 0 332 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_44
timestamp 1732942776
transform -1 0 348 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1732942776
transform -1 0 444 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1732942776
transform 1 0 444 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_0_0
timestamp 1732942776
transform 1 0 540 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1732942776
transform 1 0 548 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_108
timestamp 1732942776
transform 1 0 556 0 1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_37
timestamp 1732942776
transform -1 0 660 0 1 1305
box -2 -3 74 103
use BUFX4  BUFX4_17
timestamp 1732942776
transform -1 0 692 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_16
timestamp 1732942776
transform -1 0 724 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_248
timestamp 1732942776
transform 1 0 724 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1732942776
transform 1 0 772 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_164
timestamp 1732942776
transform -1 0 900 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1732942776
transform -1 0 996 0 1 1305
box -2 -3 98 103
use NAND3X1  NAND3X1_12
timestamp 1732942776
transform -1 0 1028 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_100
timestamp 1732942776
transform 1 0 1028 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_1_0
timestamp 1732942776
transform -1 0 1060 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1732942776
transform -1 0 1068 0 1 1305
box -2 -3 10 103
use AOI22X1  AOI22X1_12
timestamp 1732942776
transform -1 0 1108 0 1 1305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1732942776
transform 1 0 1108 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_36
timestamp 1732942776
transform 1 0 1204 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1732942776
transform -1 0 1260 0 1 1305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_49
timestamp 1732942776
transform 1 0 1260 0 1 1305
box -2 -3 74 103
use BUFX4  BUFX4_14
timestamp 1732942776
transform -1 0 1364 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1732942776
transform 1 0 1364 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_19
timestamp 1732942776
transform -1 0 1404 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1732942776
transform 1 0 1404 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_82
timestamp 1732942776
transform -1 0 1452 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_91
timestamp 1732942776
transform 1 0 1452 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_20
timestamp 1732942776
transform -1 0 1500 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1732942776
transform -1 0 1524 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_54
timestamp 1732942776
transform -1 0 1548 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_155
timestamp 1732942776
transform -1 0 1572 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_2_0
timestamp 1732942776
transform -1 0 1580 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1732942776
transform -1 0 1588 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_153
timestamp 1732942776
transform -1 0 1612 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_58
timestamp 1732942776
transform 1 0 1612 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_175
timestamp 1732942776
transform -1 0 1660 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_45
timestamp 1732942776
transform 1 0 1660 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1732942776
transform -1 0 1780 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_19
timestamp 1732942776
transform 1 0 1780 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_19
timestamp 1732942776
transform -1 0 1844 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1732942776
transform 1 0 1844 0 1 1305
box -2 -3 98 103
use INVX2  INVX2_6
timestamp 1732942776
transform 1 0 1940 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_110
timestamp 1732942776
transform -1 0 2004 0 1 1305
box -2 -3 50 103
use AOI22X1  AOI22X1_9
timestamp 1732942776
transform -1 0 2044 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_135
timestamp 1732942776
transform 1 0 2044 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1732942776
transform -1 0 2084 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_3_0
timestamp 1732942776
transform 1 0 2084 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1732942776
transform 1 0 2092 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_6
timestamp 1732942776
transform 1 0 2100 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_107
timestamp 1732942776
transform -1 0 2180 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_9
timestamp 1732942776
transform -1 0 2212 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_12
timestamp 1732942776
transform -1 0 2236 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1732942776
transform -1 0 2332 0 1 1305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_32
timestamp 1732942776
transform -1 0 2404 0 1 1305
box -2 -3 74 103
use AOI21X1  AOI21X1_37
timestamp 1732942776
transform 1 0 2404 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1732942776
transform -1 0 2532 0 1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_36
timestamp 1732942776
transform 1 0 2532 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1732942776
transform 1 0 2564 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_43
timestamp 1732942776
transform 1 0 2588 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1732942776
transform 1 0 2612 0 1 1305
box -2 -3 26 103
use FILL  FILL_14_1
timestamp 1732942776
transform 1 0 2636 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1732942776
transform 1 0 2644 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1732942776
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_67
timestamp 1732942776
transform -1 0 132 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_3
timestamp 1732942776
transform 1 0 132 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1732942776
transform -1 0 188 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_126
timestamp 1732942776
transform 1 0 188 0 -1 1505
box -2 -3 50 103
use CLKBUF1  CLKBUF1_51
timestamp 1732942776
transform 1 0 236 0 -1 1505
box -2 -3 74 103
use MUX2X1  MUX2X1_36
timestamp 1732942776
transform 1 0 308 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_36
timestamp 1732942776
transform -1 0 372 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_141
timestamp 1732942776
transform 1 0 372 0 -1 1505
box -2 -3 50 103
use CLKBUF1  CLKBUF1_23
timestamp 1732942776
transform 1 0 420 0 -1 1505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1732942776
transform 1 0 492 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_0_0
timestamp 1732942776
transform 1 0 588 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1732942776
transform 1 0 596 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_8
timestamp 1732942776
transform 1 0 604 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1732942776
transform -1 0 660 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_143
timestamp 1732942776
transform 1 0 660 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_246
timestamp 1732942776
transform 1 0 708 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1732942776
transform -1 0 852 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_16
timestamp 1732942776
transform 1 0 852 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_16
timestamp 1732942776
transform -1 0 916 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_30
timestamp 1732942776
transform 1 0 916 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_30
timestamp 1732942776
transform -1 0 980 0 -1 1505
box -2 -3 50 103
use NAND3X1  NAND3X1_9
timestamp 1732942776
transform -1 0 1012 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1732942776
transform 1 0 1012 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_1_0
timestamp 1732942776
transform 1 0 1044 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1732942776
transform 1 0 1052 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_7
timestamp 1732942776
transform 1 0 1060 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1732942776
transform 1 0 1092 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_59
timestamp 1732942776
transform -1 0 1220 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1732942776
transform -1 0 1316 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_9
timestamp 1732942776
transform -1 0 1340 0 -1 1505
box -2 -3 26 103
use INVX2  INVX2_1
timestamp 1732942776
transform -1 0 1356 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_11
timestamp 1732942776
transform 1 0 1356 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1732942776
transform 1 0 1380 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1732942776
transform -1 0 1444 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1732942776
transform 1 0 1444 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1732942776
transform 1 0 1476 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1732942776
transform 1 0 1508 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_63
timestamp 1732942776
transform 1 0 1540 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_2_0
timestamp 1732942776
transform 1 0 1564 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1732942776
transform 1 0 1572 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_81
timestamp 1732942776
transform 1 0 1580 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1732942776
transform -1 0 1636 0 -1 1505
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1732942776
transform -1 0 1676 0 -1 1505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1732942776
transform -1 0 1772 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_251
timestamp 1732942776
transform 1 0 1772 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_61
timestamp 1732942776
transform -1 0 1836 0 -1 1505
box -2 -3 18 103
use BUFX4  BUFX4_10
timestamp 1732942776
transform 1 0 1836 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1732942776
transform -1 0 1964 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_109
timestamp 1732942776
transform -1 0 2012 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_85
timestamp 1732942776
transform 1 0 2012 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1732942776
transform -1 0 2076 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1732942776
transform -1 0 2084 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1732942776
transform -1 0 2092 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1732942776
transform -1 0 2188 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_7
timestamp 1732942776
transform 1 0 2188 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_66
timestamp 1732942776
transform -1 0 2268 0 -1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_48
timestamp 1732942776
transform 1 0 2268 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1732942776
transform -1 0 2324 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1732942776
transform 1 0 2324 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_49
timestamp 1732942776
transform 1 0 2420 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1732942776
transform -1 0 2476 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_134
timestamp 1732942776
transform 1 0 2476 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1732942776
transform -1 0 2596 0 -1 1505
box -2 -3 98 103
use INVX8  INVX8_5
timestamp 1732942776
transform -1 0 2636 0 -1 1505
box -2 -3 42 103
use FILL  FILL_15_1
timestamp 1732942776
transform -1 0 2644 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1732942776
transform -1 0 2652 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1732942776
transform 1 0 4 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_74
timestamp 1732942776
transform 1 0 100 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1732942776
transform 1 0 4 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_125
timestamp 1732942776
transform 1 0 100 0 -1 1705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_22
timestamp 1732942776
transform 1 0 124 0 1 1505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1732942776
transform 1 0 196 0 1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_126
timestamp 1732942776
transform -1 0 156 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1732942776
transform 1 0 156 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1732942776
transform 1 0 292 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_64
timestamp 1732942776
transform 1 0 252 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_254
timestamp 1732942776
transform -1 0 316 0 -1 1705
box -2 -3 50 103
use NOR2X1  NOR2X1_9
timestamp 1732942776
transform 1 0 388 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_120
timestamp 1732942776
transform 1 0 316 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_121
timestamp 1732942776
transform -1 0 372 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1732942776
transform -1 0 404 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1732942776
transform -1 0 500 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_8
timestamp 1732942776
transform -1 0 444 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1732942776
transform -1 0 476 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_256
timestamp 1732942776
transform 1 0 476 0 1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_53
timestamp 1732942776
transform -1 0 532 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1732942776
transform -1 0 540 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_0_0
timestamp 1732942776
transform 1 0 540 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1732942776
transform 1 0 548 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1732942776
transform 1 0 556 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_0_0
timestamp 1732942776
transform -1 0 540 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1732942776
transform -1 0 548 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1732942776
transform -1 0 644 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1732942776
transform 1 0 652 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_127
timestamp 1732942776
transform 1 0 644 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_128
timestamp 1732942776
transform -1 0 700 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1732942776
transform -1 0 796 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_231
timestamp 1732942776
transform -1 0 796 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_69
timestamp 1732942776
transform 1 0 796 0 1 1505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_11
timestamp 1732942776
transform 1 0 796 0 -1 1705
box -2 -3 74 103
use OAI21X1  OAI21X1_62
timestamp 1732942776
transform -1 0 852 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_184
timestamp 1732942776
transform -1 0 900 0 1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1732942776
transform 1 0 900 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_183
timestamp 1732942776
transform -1 0 916 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_195
timestamp 1732942776
transform 1 0 996 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_233
timestamp 1732942776
transform -1 0 964 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_145
timestamp 1732942776
transform 1 0 964 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_185
timestamp 1732942776
transform 1 0 988 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_25
timestamp 1732942776
transform 1 0 1044 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_1_0
timestamp 1732942776
transform -1 0 1076 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1732942776
transform -1 0 1084 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_22
timestamp 1732942776
transform -1 0 1116 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1_0
timestamp 1732942776
transform 1 0 1036 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1732942776
transform 1 0 1044 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1732942776
transform 1 0 1052 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_102
timestamp 1732942776
transform 1 0 1116 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_66
timestamp 1732942776
transform 1 0 1140 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1732942776
transform 1 0 1164 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_8
timestamp 1732942776
transform 1 0 1148 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_8
timestamp 1732942776
transform -1 0 1212 0 -1 1705
box -2 -3 50 103
use BUFX4  BUFX4_41
timestamp 1732942776
transform 1 0 1212 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1732942776
transform 1 0 1260 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1732942776
transform -1 0 1324 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_228
timestamp 1732942776
transform 1 0 1244 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_229
timestamp 1732942776
transform 1 0 1292 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1732942776
transform 1 0 1324 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_230
timestamp 1732942776
transform -1 0 1388 0 -1 1705
box -2 -3 50 103
use AOI22X1  AOI22X1_29
timestamp 1732942776
transform -1 0 1428 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_80
timestamp 1732942776
transform -1 0 1444 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_37
timestamp 1732942776
transform 1 0 1444 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_32
timestamp 1732942776
transform -1 0 1500 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1732942776
transform -1 0 1524 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_150
timestamp 1732942776
transform 1 0 1428 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_136
timestamp 1732942776
transform 1 0 1452 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_30
timestamp 1732942776
transform 1 0 1484 0 -1 1705
box -2 -3 42 103
use FILL  FILL_15_2_0
timestamp 1732942776
transform -1 0 1532 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1732942776
transform -1 0 1540 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1732942776
transform -1 0 1636 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_235
timestamp 1732942776
transform -1 0 1572 0 -1 1705
box -2 -3 50 103
use FILL  FILL_16_2_0
timestamp 1732942776
transform -1 0 1580 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1732942776
transform -1 0 1588 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_236
timestamp 1732942776
transform -1 0 1636 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_35
timestamp 1732942776
transform -1 0 1660 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_30
timestamp 1732942776
transform -1 0 1692 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_19
timestamp 1732942776
transform 1 0 1692 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1732942776
transform 1 0 1716 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_234
timestamp 1732942776
transform 1 0 1636 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_82
timestamp 1732942776
transform 1 0 1684 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_65
timestamp 1732942776
transform 1 0 1716 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_81
timestamp 1732942776
transform 1 0 1748 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_187
timestamp 1732942776
transform -1 0 1828 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_188
timestamp 1732942776
transform 1 0 1764 0 -1 1705
box -2 -3 50 103
use AOI21X1  AOI21X1_14
timestamp 1732942776
transform 1 0 1812 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1732942776
transform 1 0 1828 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_17
timestamp 1732942776
transform 1 0 1844 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_22
timestamp 1732942776
transform 1 0 1868 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_144
timestamp 1732942776
transform -1 0 1932 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_92
timestamp 1732942776
transform 1 0 1924 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1732942776
transform 1 0 1956 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1732942776
transform 1 0 1988 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_91
timestamp 1732942776
transform -1 0 2044 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_134
timestamp 1732942776
transform 1 0 1932 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1732942776
transform 1 0 1964 0 -1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_129
timestamp 1732942776
transform -1 0 2036 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_111
timestamp 1732942776
transform -1 0 2092 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_3_0
timestamp 1732942776
transform -1 0 2100 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1732942776
transform -1 0 2108 0 1 1505
box -2 -3 10 103
use AOI22X1  AOI22X1_10
timestamp 1732942776
transform -1 0 2148 0 1 1505
box -2 -3 42 103
use FILL  FILL_16_3_0
timestamp 1732942776
transform -1 0 2044 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1732942776
transform -1 0 2052 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1732942776
transform -1 0 2148 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_113
timestamp 1732942776
transform 1 0 2148 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_68
timestamp 1732942776
transform -1 0 2244 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_11
timestamp 1732942776
transform 1 0 2148 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_11
timestamp 1732942776
transform -1 0 2212 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_116
timestamp 1732942776
transform -1 0 2260 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_115
timestamp 1732942776
transform 1 0 2244 0 1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_38
timestamp 1732942776
transform -1 0 2324 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1732942776
transform 1 0 2324 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_67
timestamp 1732942776
transform -1 0 2308 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_114
timestamp 1732942776
transform -1 0 2356 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_128
timestamp 1732942776
transform -1 0 2444 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_33
timestamp 1732942776
transform -1 0 2388 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1732942776
transform -1 0 2412 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1732942776
transform -1 0 2444 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1732942776
transform 1 0 2444 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_27
timestamp 1732942776
transform -1 0 2500 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1732942776
transform 1 0 2500 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_25
timestamp 1732942776
transform -1 0 2556 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1732942776
transform 1 0 2444 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1732942776
transform -1 0 2564 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1732942776
transform -1 0 2652 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_43
timestamp 1732942776
transform -1 0 2596 0 -1 1705
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1732942776
transform 1 0 2596 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1732942776
transform 1 0 2620 0 -1 1705
box -2 -3 26 103
use FILL  FILL_17_1
timestamp 1732942776
transform -1 0 2652 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1732942776
transform -1 0 100 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_49
timestamp 1732942776
transform -1 0 148 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_193
timestamp 1732942776
transform 1 0 148 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_194
timestamp 1732942776
transform -1 0 244 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_73
timestamp 1732942776
transform -1 0 292 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_74
timestamp 1732942776
transform -1 0 340 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_72
timestamp 1732942776
transform -1 0 364 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_23
timestamp 1732942776
transform 1 0 364 0 1 1705
box -2 -3 42 103
use AOI22X1  AOI22X1_3
timestamp 1732942776
transform 1 0 404 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_42
timestamp 1732942776
transform -1 0 476 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_57
timestamp 1732942776
transform -1 0 500 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_240
timestamp 1732942776
transform -1 0 548 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_0_0
timestamp 1732942776
transform 1 0 548 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1732942776
transform 1 0 556 0 1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_242
timestamp 1732942776
transform 1 0 564 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_241
timestamp 1732942776
transform -1 0 660 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_79
timestamp 1732942776
transform 1 0 660 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1732942776
transform -1 0 716 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1732942776
transform -1 0 812 0 1 1705
box -2 -3 98 103
use AOI22X1  AOI22X1_31
timestamp 1732942776
transform -1 0 852 0 1 1705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1732942776
transform -1 0 948 0 1 1705
box -2 -3 98 103
use AOI22X1  AOI22X1_24
timestamp 1732942776
transform -1 0 988 0 1 1705
box -2 -3 42 103
use MUX2X1  MUX2X1_197
timestamp 1732942776
transform -1 0 1036 0 1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_130
timestamp 1732942776
transform 1 0 1036 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_1_0
timestamp 1732942776
transform -1 0 1068 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1732942776
transform -1 0 1076 0 1 1705
box -2 -3 10 103
use AOI22X1  AOI22X1_4
timestamp 1732942776
transform -1 0 1116 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_151
timestamp 1732942776
transform 1 0 1116 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_32
timestamp 1732942776
transform -1 0 1180 0 1 1705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1732942776
transform -1 0 1276 0 1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_29
timestamp 1732942776
transform 1 0 1276 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1732942776
transform -1 0 1332 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1732942776
transform 1 0 1332 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_24
timestamp 1732942776
transform 1 0 1428 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_24
timestamp 1732942776
transform -1 0 1492 0 1 1705
box -2 -3 50 103
use AOI21X1  AOI21X1_45
timestamp 1732942776
transform 1 0 1492 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_149
timestamp 1732942776
transform -1 0 1548 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_2_0
timestamp 1732942776
transform 1 0 1548 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1732942776
transform 1 0 1556 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1732942776
transform 1 0 1564 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_25
timestamp 1732942776
transform 1 0 1660 0 1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_25
timestamp 1732942776
transform -1 0 1724 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1732942776
transform 1 0 1724 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1732942776
transform -1 0 1916 0 1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_22
timestamp 1732942776
transform 1 0 1916 0 1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1732942776
transform 1 0 1964 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_22
timestamp 1732942776
transform -1 0 2076 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_3_0
timestamp 1732942776
transform -1 0 2084 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1732942776
transform -1 0 2092 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_129
timestamp 1732942776
transform -1 0 2116 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_1
timestamp 1732942776
transform 1 0 2116 0 1 1705
box -2 -3 42 103
use AOI22X1  AOI22X1_21
timestamp 1732942776
transform -1 0 2196 0 1 1705
box -2 -3 42 103
use MUX2X1  MUX2X1_181
timestamp 1732942776
transform -1 0 2244 0 1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_105
timestamp 1732942776
transform 1 0 2244 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_141
timestamp 1732942776
transform -1 0 2324 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1732942776
transform -1 0 2356 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1732942776
transform -1 0 2380 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1732942776
transform -1 0 2476 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_51
timestamp 1732942776
transform -1 0 2508 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1732942776
transform -1 0 2604 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_143
timestamp 1732942776
transform -1 0 2628 0 1 1705
box -2 -3 26 103
use FILL  FILL_18_1
timestamp 1732942776
transform 1 0 2628 0 1 1705
box -2 -3 10 103
use FILL  FILL_18_2
timestamp 1732942776
transform 1 0 2636 0 1 1705
box -2 -3 10 103
use FILL  FILL_18_3
timestamp 1732942776
transform 1 0 2644 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1732942776
transform 1 0 4 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_50
timestamp 1732942776
transform 1 0 100 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_70
timestamp 1732942776
transform -1 0 164 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1732942776
transform 1 0 164 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_33
timestamp 1732942776
transform 1 0 260 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_33
timestamp 1732942776
transform -1 0 324 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_191
timestamp 1732942776
transform -1 0 372 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_71
timestamp 1732942776
transform -1 0 420 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_69
timestamp 1732942776
transform 1 0 420 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_6
timestamp 1732942776
transform 1 0 468 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_198
timestamp 1732942776
transform 1 0 492 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_0_0
timestamp 1732942776
transform 1 0 540 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1732942776
transform 1 0 548 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_200
timestamp 1732942776
transform 1 0 556 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_199
timestamp 1732942776
transform 1 0 604 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_110
timestamp 1732942776
transform 1 0 652 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_32
timestamp 1732942776
transform 1 0 676 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_32
timestamp 1732942776
transform -1 0 740 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1732942776
transform 1 0 740 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_232
timestamp 1732942776
transform 1 0 836 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_14
timestamp 1732942776
transform 1 0 884 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_14
timestamp 1732942776
transform -1 0 948 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_80
timestamp 1732942776
transform -1 0 996 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_196
timestamp 1732942776
transform -1 0 1044 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_1_0
timestamp 1732942776
transform -1 0 1052 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1732942776
transform -1 0 1060 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1732942776
transform -1 0 1156 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_15
timestamp 1732942776
transform 1 0 1156 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_14
timestamp 1732942776
transform -1 0 1212 0 -1 1905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_44
timestamp 1732942776
transform 1 0 1212 0 -1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1732942776
transform 1 0 1284 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_120
timestamp 1732942776
transform 1 0 1380 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1732942776
transform -1 0 1436 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_269
timestamp 1732942776
transform 1 0 1436 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_2_0
timestamp 1732942776
transform 1 0 1532 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1732942776
transform 1 0 1540 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1732942776
transform 1 0 1548 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_58
timestamp 1732942776
transform 1 0 1644 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_249
timestamp 1732942776
transform -1 0 1708 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_63
timestamp 1732942776
transform -1 0 1756 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_64
timestamp 1732942776
transform 1 0 1756 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_186
timestamp 1732942776
transform 1 0 1804 0 -1 1905
box -2 -3 50 103
use BUFX4  BUFX4_4
timestamp 1732942776
transform 1 0 1852 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_61
timestamp 1732942776
transform 1 0 1884 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_62
timestamp 1732942776
transform -1 0 1980 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_57
timestamp 1732942776
transform -1 0 2028 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_59
timestamp 1732942776
transform 1 0 2028 0 -1 1905
box -2 -3 50 103
use FILL  FILL_18_3_0
timestamp 1732942776
transform 1 0 2076 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1732942776
transform 1 0 2084 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_180
timestamp 1732942776
transform 1 0 2092 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_182
timestamp 1732942776
transform 1 0 2140 0 -1 1905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1732942776
transform 1 0 2188 0 -1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_112
timestamp 1732942776
transform -1 0 2332 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_58
timestamp 1732942776
transform -1 0 2380 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_112
timestamp 1732942776
transform 1 0 2380 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_113
timestamp 1732942776
transform -1 0 2436 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1732942776
transform -1 0 2532 0 -1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_31
timestamp 1732942776
transform 1 0 2532 0 -1 1905
box -2 -3 74 103
use NAND2X1  NAND2X1_46
timestamp 1732942776
transform -1 0 2628 0 -1 1905
box -2 -3 26 103
use FILL  FILL_19_1
timestamp 1732942776
transform -1 0 2636 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_2
timestamp 1732942776
transform -1 0 2644 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_3
timestamp 1732942776
transform -1 0 2652 0 -1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_30
timestamp 1732942776
transform 1 0 4 0 1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1732942776
transform 1 0 76 0 1 1905
box -2 -3 98 103
use NOR2X1  NOR2X1_32
timestamp 1732942776
transform 1 0 172 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1732942776
transform -1 0 228 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_77
timestamp 1732942776
transform 1 0 228 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_70
timestamp 1732942776
transform -1 0 284 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1732942776
transform -1 0 380 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1732942776
transform 1 0 380 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_6
timestamp 1732942776
transform -1 0 508 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_0_0
timestamp 1732942776
transform -1 0 516 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1732942776
transform -1 0 524 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1732942776
transform -1 0 620 0 1 1905
box -2 -3 98 103
use AOI21X1  AOI21X1_6
timestamp 1732942776
transform 1 0 620 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1732942776
transform 1 0 652 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_112
timestamp 1732942776
transform -1 0 708 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1732942776
transform -1 0 804 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_239
timestamp 1732942776
transform 1 0 804 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_71
timestamp 1732942776
transform -1 0 876 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_48
timestamp 1732942776
transform 1 0 876 0 1 1905
box -2 -3 50 103
use INVX1  INVX1_48
timestamp 1732942776
transform -1 0 940 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1732942776
transform -1 0 1036 0 1 1905
box -2 -3 98 103
use BUFX4  BUFX4_56
timestamp 1732942776
transform -1 0 1068 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_1_0
timestamp 1732942776
transform -1 0 1076 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1732942776
transform -1 0 1084 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1732942776
transform -1 0 1180 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_164
timestamp 1732942776
transform 1 0 1180 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_158
timestamp 1732942776
transform -1 0 1236 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1732942776
transform -1 0 1268 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1732942776
transform -1 0 1292 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_40
timestamp 1732942776
transform -1 0 1324 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1732942776
transform 1 0 1324 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_226
timestamp 1732942776
transform 1 0 1420 0 1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_227
timestamp 1732942776
transform -1 0 1516 0 1 1905
box -2 -3 50 103
use BUFX2  BUFX2_8
timestamp 1732942776
transform 1 0 1516 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_56
timestamp 1732942776
transform 1 0 1540 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1732942776
transform -1 0 1580 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1732942776
transform -1 0 1588 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_62
timestamp 1732942776
transform -1 0 1612 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1732942776
transform -1 0 1708 0 1 1905
box -2 -3 98 103
use BUFX4  BUFX4_59
timestamp 1732942776
transform -1 0 1740 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1732942776
transform 1 0 1740 0 1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_9
timestamp 1732942776
transform -1 0 1804 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_60
timestamp 1732942776
transform 1 0 1804 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_54
timestamp 1732942776
transform -1 0 1860 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_17
timestamp 1732942776
transform 1 0 1860 0 1 1905
box -2 -3 50 103
use INVX1  INVX1_17
timestamp 1732942776
transform -1 0 1924 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1732942776
transform -1 0 2020 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1732942776
transform -1 0 2116 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_3_0
timestamp 1732942776
transform 1 0 2116 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1732942776
transform 1 0 2124 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_83
timestamp 1732942776
transform 1 0 2132 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_73
timestamp 1732942776
transform -1 0 2188 0 1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_179
timestamp 1732942776
transform 1 0 2188 0 1 1905
box -2 -3 50 103
use BUFX4  BUFX4_58
timestamp 1732942776
transform 1 0 2236 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_59
timestamp 1732942776
transform 1 0 2268 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1732942776
transform -1 0 2324 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1732942776
transform -1 0 2420 0 1 1905
box -2 -3 98 103
use MUX2X1  MUX2X1_27
timestamp 1732942776
transform 1 0 2420 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_78
timestamp 1732942776
transform 1 0 2468 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_27
timestamp 1732942776
transform -1 0 2516 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1732942776
transform -1 0 2612 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_41
timestamp 1732942776
transform 1 0 2612 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1732942776
transform 1 0 2644 0 1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1732942776
transform 1 0 4 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_105
timestamp 1732942776
transform -1 0 132 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1732942776
transform -1 0 156 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_55
timestamp 1732942776
transform -1 0 172 0 -1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_54
timestamp 1732942776
transform -1 0 220 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_192
timestamp 1732942776
transform -1 0 268 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_190
timestamp 1732942776
transform -1 0 316 0 -1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1732942776
transform 1 0 316 0 -1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_41
timestamp 1732942776
transform 1 0 412 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_41
timestamp 1732942776
transform -1 0 476 0 -1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_72
timestamp 1732942776
transform 1 0 476 0 -1 2105
box -2 -3 50 103
use FILL  FILL_20_0_0
timestamp 1732942776
transform 1 0 524 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1732942776
transform 1 0 532 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1732942776
transform 1 0 540 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_53
timestamp 1732942776
transform 1 0 636 0 -1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_52
timestamp 1732942776
transform -1 0 700 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_142
timestamp 1732942776
transform -1 0 748 0 -1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_35
timestamp 1732942776
transform 1 0 748 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_28
timestamp 1732942776
transform -1 0 804 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1732942776
transform 1 0 804 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_64
timestamp 1732942776
transform -1 0 932 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_237
timestamp 1732942776
transform 1 0 932 0 -1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_2
timestamp 1732942776
transform 1 0 980 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_78
timestamp 1732942776
transform -1 0 1052 0 -1 2105
box -2 -3 50 103
use FILL  FILL_20_1_0
timestamp 1732942776
transform 1 0 1052 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1732942776
transform 1 0 1060 0 -1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_238
timestamp 1732942776
transform 1 0 1068 0 -1 2105
box -2 -3 50 103
use MUX2X1  MUX2X1_56
timestamp 1732942776
transform 1 0 1116 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_1
timestamp 1732942776
transform 1 0 1164 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1732942776
transform -1 0 1220 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1732942776
transform -1 0 1316 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1732942776
transform 1 0 1316 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_80
timestamp 1732942776
transform 1 0 1412 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_90
timestamp 1732942776
transform -1 0 1468 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_225
timestamp 1732942776
transform 1 0 1468 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_151
timestamp 1732942776
transform -1 0 1548 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1732942776
transform -1 0 1580 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_2_0
timestamp 1732942776
transform 1 0 1580 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1732942776
transform 1 0 1588 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_48
timestamp 1732942776
transform 1 0 1596 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_53
timestamp 1732942776
transform -1 0 1652 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1732942776
transform -1 0 1748 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1732942776
transform -1 0 1844 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1732942776
transform -1 0 1940 0 -1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_138
timestamp 1732942776
transform 1 0 1940 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1732942776
transform -1 0 2004 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_60
timestamp 1732942776
transform 1 0 2004 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_1
timestamp 1732942776
transform 1 0 2052 0 -1 2105
box -2 -3 18 103
use FILL  FILL_20_3_0
timestamp 1732942776
transform -1 0 2076 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1732942776
transform -1 0 2084 0 -1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_1
timestamp 1732942776
transform -1 0 2132 0 -1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_27
timestamp 1732942776
transform 1 0 2132 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1732942776
transform -1 0 2188 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_177
timestamp 1732942776
transform 1 0 2188 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_147
timestamp 1732942776
transform 1 0 2236 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_148
timestamp 1732942776
transform -1 0 2300 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1732942776
transform -1 0 2396 0 -1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_6
timestamp 1732942776
transform 1 0 2396 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_6
timestamp 1732942776
transform -1 0 2460 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1732942776
transform -1 0 2556 0 -1 2105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_40
timestamp 1732942776
transform 1 0 2556 0 -1 2105
box -2 -3 74 103
use FILL  FILL_21_1
timestamp 1732942776
transform -1 0 2636 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_2
timestamp 1732942776
transform -1 0 2644 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_3
timestamp 1732942776
transform -1 0 2652 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1732942776
transform -1 0 100 0 1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_37
timestamp 1732942776
transform 1 0 100 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1732942776
transform -1 0 156 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1732942776
transform -1 0 252 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1732942776
transform -1 0 348 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_108
timestamp 1732942776
transform 1 0 348 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_110
timestamp 1732942776
transform -1 0 404 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1732942776
transform -1 0 436 0 1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_46
timestamp 1732942776
transform 1 0 436 0 1 2105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1732942776
transform 1 0 484 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_0_0
timestamp 1732942776
transform 1 0 580 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1732942776
transform 1 0 588 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_172
timestamp 1732942776
transform 1 0 596 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_166
timestamp 1732942776
transform -1 0 652 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1732942776
transform 1 0 652 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_97
timestamp 1732942776
transform -1 0 708 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1732942776
transform -1 0 804 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1732942776
transform -1 0 900 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1732942776
transform 1 0 900 0 1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_1
timestamp 1732942776
transform -1 0 1028 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_1_0
timestamp 1732942776
transform -1 0 1036 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1732942776
transform -1 0 1044 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1732942776
transform -1 0 1140 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_57
timestamp 1732942776
transform 1 0 1140 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_39
timestamp 1732942776
transform 1 0 1156 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_32
timestamp 1732942776
transform -1 0 1212 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1732942776
transform -1 0 1308 0 1 2105
box -2 -3 98 103
use MUX2X1  MUX2X1_245
timestamp 1732942776
transform -1 0 1356 0 1 2105
box -2 -3 50 103
use BUFX4  BUFX4_43
timestamp 1732942776
transform -1 0 1388 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1732942776
transform 1 0 1388 0 1 2105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_3
timestamp 1732942776
transform -1 0 1492 0 1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1732942776
transform -1 0 1588 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_2_0
timestamp 1732942776
transform -1 0 1596 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1732942776
transform -1 0 1604 0 1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_64
timestamp 1732942776
transform -1 0 1676 0 1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1732942776
transform -1 0 1772 0 1 2105
box -2 -3 98 103
use NAND2X1  NAND2X1_22
timestamp 1732942776
transform 1 0 1772 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_19
timestamp 1732942776
transform -1 0 1828 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1732942776
transform -1 0 1860 0 1 2105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_12
timestamp 1732942776
transform -1 0 1932 0 1 2105
box -2 -3 74 103
use OAI21X1  OAI21X1_57
timestamp 1732942776
transform 1 0 1932 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_64
timestamp 1732942776
transform -1 0 1988 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1732942776
transform -1 0 2084 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_3_0
timestamp 1732942776
transform 1 0 2084 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1732942776
transform 1 0 2092 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1732942776
transform 1 0 2100 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_5
timestamp 1732942776
transform 1 0 2196 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1732942776
transform -1 0 2260 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1732942776
transform -1 0 2356 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1732942776
transform -1 0 2452 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1732942776
transform 1 0 2452 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1732942776
transform 1 0 2548 0 1 2105
box -2 -3 98 103
use FILL  FILL_22_1
timestamp 1732942776
transform 1 0 2644 0 1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_29
timestamp 1732942776
transform 1 0 4 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1732942776
transform 1 0 76 0 -1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_51
timestamp 1732942776
transform 1 0 172 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_55
timestamp 1732942776
transform -1 0 228 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1732942776
transform 1 0 228 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_38
timestamp 1732942776
transform 1 0 324 0 -1 2305
box -2 -3 50 103
use INVX1  INVX1_38
timestamp 1732942776
transform -1 0 388 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_189
timestamp 1732942776
transform 1 0 388 0 -1 2305
box -2 -3 50 103
use BUFX4  BUFX4_1
timestamp 1732942776
transform -1 0 468 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_46
timestamp 1732942776
transform -1 0 484 0 -1 2305
box -2 -3 18 103
use INVX8  INVX8_8
timestamp 1732942776
transform 1 0 484 0 -1 2305
box -2 -3 42 103
use FILL  FILL_22_0_0
timestamp 1732942776
transform 1 0 524 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1732942776
transform 1 0 532 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1732942776
transform 1 0 540 0 -1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_97
timestamp 1732942776
transform 1 0 636 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1732942776
transform -1 0 692 0 -1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_79
timestamp 1732942776
transform -1 0 740 0 -1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1732942776
transform -1 0 836 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_50
timestamp 1732942776
transform 1 0 836 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_46
timestamp 1732942776
transform -1 0 892 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_33
timestamp 1732942776
transform 1 0 892 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1732942776
transform 1 0 964 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_1_0
timestamp 1732942776
transform 1 0 1060 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1732942776
transform 1 0 1068 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_76
timestamp 1732942776
transform 1 0 1076 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_10
timestamp 1732942776
transform 1 0 1124 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_55
timestamp 1732942776
transform 1 0 1148 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_10
timestamp 1732942776
transform 1 0 1180 0 -1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_77
timestamp 1732942776
transform -1 0 1268 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_244
timestamp 1732942776
transform 1 0 1268 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_243
timestamp 1732942776
transform 1 0 1316 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_27
timestamp 1732942776
transform 1 0 1364 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_24
timestamp 1732942776
transform -1 0 1420 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1732942776
transform -1 0 1516 0 -1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_125
timestamp 1732942776
transform 1 0 1516 0 -1 2305
box -2 -3 50 103
use FILL  FILL_22_2_0
timestamp 1732942776
transform -1 0 1572 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1732942776
transform -1 0 1580 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_123
timestamp 1732942776
transform -1 0 1628 0 -1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1732942776
transform -1 0 1724 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_63
timestamp 1732942776
transform 1 0 1724 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_56
timestamp 1732942776
transform -1 0 1780 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_75
timestamp 1732942776
transform -1 0 1828 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_20
timestamp 1732942776
transform -1 0 1852 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1732942776
transform -1 0 1948 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_61
timestamp 1732942776
transform 1 0 1948 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_54
timestamp 1732942776
transform -1 0 2004 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1732942776
transform -1 0 2100 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_3_0
timestamp 1732942776
transform 1 0 2100 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1732942776
transform 1 0 2108 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_22
timestamp 1732942776
transform 1 0 2116 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1732942776
transform -1 0 2172 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1732942776
transform 1 0 2172 0 -1 2305
box -2 -3 98 103
use INVX8  INVX8_3
timestamp 1732942776
transform -1 0 2308 0 -1 2305
box -2 -3 42 103
use MUX2X1  MUX2X1_178
timestamp 1732942776
transform -1 0 2356 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_38
timestamp 1732942776
transform 1 0 2356 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1732942776
transform -1 0 2412 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_117
timestamp 1732942776
transform 1 0 2412 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_118
timestamp 1732942776
transform -1 0 2468 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_52
timestamp 1732942776
transform -1 0 2540 0 -1 2305
box -2 -3 74 103
use NAND2X1  NAND2X1_56
timestamp 1732942776
transform -1 0 2564 0 -1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_10
timestamp 1732942776
transform 1 0 2564 0 -1 2305
box -2 -3 74 103
use FILL  FILL_23_1
timestamp 1732942776
transform -1 0 2644 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_2
timestamp 1732942776
transform -1 0 2652 0 -1 2305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_65
timestamp 1732942776
transform 1 0 4 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_67
timestamp 1732942776
transform 1 0 76 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_43
timestamp 1732942776
transform -1 0 220 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_63
timestamp 1732942776
transform 1 0 220 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_9
timestamp 1732942776
transform 1 0 292 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_20
timestamp 1732942776
transform 1 0 364 0 1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1732942776
transform 1 0 436 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_0_0
timestamp 1732942776
transform 1 0 532 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1732942776
transform 1 0 540 0 1 2305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_50
timestamp 1732942776
transform 1 0 548 0 1 2305
box -2 -3 74 103
use OAI21X1  OAI21X1_161
timestamp 1732942776
transform 1 0 620 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1732942776
transform -1 0 676 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1732942776
transform 1 0 676 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1732942776
transform 1 0 772 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_40
timestamp 1732942776
transform 1 0 868 0 1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_40
timestamp 1732942776
transform -1 0 932 0 1 2305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1732942776
transform 1 0 932 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_153
timestamp 1732942776
transform -1 0 1060 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_1_0
timestamp 1732942776
transform -1 0 1068 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1732942776
transform -1 0 1076 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_159
timestamp 1732942776
transform -1 0 1100 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1732942776
transform 1 0 1100 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1732942776
transform 1 0 1132 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_160
timestamp 1732942776
transform 1 0 1228 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_166
timestamp 1732942776
transform -1 0 1284 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1732942776
transform 1 0 1284 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_17
timestamp 1732942776
transform 1 0 1380 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_16
timestamp 1732942776
transform -1 0 1436 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1732942776
transform 1 0 1436 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1732942776
transform 1 0 1468 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1732942776
transform -1 0 1588 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_2_0
timestamp 1732942776
transform -1 0 1596 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1732942776
transform -1 0 1604 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_161
timestamp 1732942776
transform -1 0 1628 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_155
timestamp 1732942776
transform -1 0 1660 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1732942776
transform 1 0 1660 0 1 2305
box -2 -3 98 103
use MUX2X1  MUX2X1_124
timestamp 1732942776
transform 1 0 1756 0 1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_12
timestamp 1732942776
transform 1 0 1804 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_11
timestamp 1732942776
transform -1 0 1860 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1732942776
transform 1 0 1860 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1732942776
transform -1 0 2052 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_3_0
timestamp 1732942776
transform -1 0 2060 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1732942776
transform -1 0 2068 0 1 2305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_17
timestamp 1732942776
transform -1 0 2140 0 1 2305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_7
timestamp 1732942776
transform -1 0 2212 0 1 2305
box -2 -3 74 103
use OAI21X1  OAI21X1_75
timestamp 1732942776
transform 1 0 2212 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1732942776
transform -1 0 2268 0 1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_54
timestamp 1732942776
transform -1 0 2340 0 1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1732942776
transform 1 0 2340 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1732942776
transform -1 0 2532 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_88
timestamp 1732942776
transform -1 0 2556 0 1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_56
timestamp 1732942776
transform 1 0 2556 0 1 2305
box -2 -3 74 103
use FILL  FILL_24_1
timestamp 1732942776
transform 1 0 2628 0 1 2305
box -2 -3 10 103
use FILL  FILL_24_2
timestamp 1732942776
transform 1 0 2636 0 1 2305
box -2 -3 10 103
use FILL  FILL_24_3
timestamp 1732942776
transform 1 0 2644 0 1 2305
box -2 -3 10 103
<< labels >>
flabel metal6 s 544 -30 560 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1056 -30 1072 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s 2678 1318 2682 1322 3 FreeSans 24 0 0 0 en
port 2 nsew
flabel metal3 s 2678 1738 2682 1742 3 FreeSans 24 0 0 0 rw
port 3 nsew
flabel metal3 s -26 2338 -22 2342 7 FreeSans 24 90 0 0 clk
port 4 nsew
flabel metal3 s 2678 1168 2682 1172 3 FreeSans 24 0 0 0 ras
port 5 nsew
flabel metal3 s 2678 1278 2682 1282 3 FreeSans 24 0 0 0 cas
port 6 nsew
flabel metal2 s 2286 2428 2290 2432 3 FreeSans 24 90 0 0 datain[0]
port 7 nsew
flabel metal2 s 510 -22 514 -18 7 FreeSans 24 270 0 0 datain[1]
port 8 nsew
flabel metal3 s 2678 1448 2682 1452 3 FreeSans 24 0 0 0 datain[2]
port 9 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 datain[3]
port 10 nsew
flabel metal2 s 1718 -22 1722 -18 7 FreeSans 24 270 0 0 datain[4]
port 11 nsew
flabel metal2 s 502 2428 506 2432 3 FreeSans 24 90 0 0 datain[5]
port 12 nsew
flabel metal2 s 1742 -22 1746 -18 7 FreeSans 24 270 0 0 datain[6]
port 13 nsew
flabel metal2 s 1198 2428 1202 2432 3 FreeSans 24 90 0 0 datain[7]
port 14 nsew
flabel metal3 s 2678 1348 2682 1352 3 FreeSans 24 0 0 0 address[0]
port 15 nsew
flabel metal3 s 2678 1368 2682 1372 3 FreeSans 24 0 0 0 address[1]
port 16 nsew
flabel metal3 s 2678 1148 2682 1152 3 FreeSans 24 0 0 0 address[2]
port 17 nsew
flabel metal3 s 2678 948 2682 952 3 FreeSans 24 0 0 0 address[3]
port 18 nsew
flabel metal3 s 2678 1048 2682 1052 3 FreeSans 24 0 0 0 address[4]
port 19 nsew
flabel metal3 s 2678 1648 2682 1652 3 FreeSans 24 0 0 0 dataout[0]
port 20 nsew
flabel metal3 s 2678 968 2682 972 3 FreeSans 24 0 0 0 dataout[1]
port 21 nsew
flabel metal3 s 2678 1248 2682 1252 3 FreeSans 24 0 0 0 dataout[2]
port 22 nsew
flabel metal3 s 2678 1298 2682 1302 3 FreeSans 24 0 0 0 dataout[3]
port 23 nsew
flabel metal3 s 2678 988 2682 992 3 FreeSans 24 0 0 0 dataout[4]
port 24 nsew
flabel metal3 s 2678 1668 2682 1672 3 FreeSans 24 0 0 0 dataout[5]
port 25 nsew
flabel metal3 s 2678 1388 2682 1392 3 FreeSans 24 0 0 0 dataout[6]
port 26 nsew
flabel metal2 s 1526 2428 1530 2432 3 FreeSans 24 90 0 0 dataout[7]
port 27 nsew
<< end >>
