* NGSPICE file created from ram32_sdram_3split.ext - technology: scmos

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt ram32_sdram_3split vdd gnd en rw clk ras cas vas datain[0] datain[1] datain[2]
+ datain[3] datain[4] datain[5] datain[6] datain[7] address[0] address[1] address[2]
+ address[3] address[4] dataout[0] dataout[1] dataout[2] dataout[3] dataout[4] dataout[5]
+ dataout[6] dataout[7]
XMUX2X1_17 MUX2X1_17/A MUX2X1_17/B BUFX4_17/Y gnd MUX2X1_18/B vdd MUX2X1
XFILL_14_3_0 gnd vdd FILL
XMUX2X1_39 MUX2X1_39/A MUX2X1_39/B INVX4_8/A gnd MUX2X1_39/Y vdd MUX2X1
XMUX2X1_28 MUX2X1_28/A MUX2X1_28/B BUFX4_16/Y gnd MUX2X1_30/A vdd MUX2X1
XNAND2X1_54 MUX2X1_61/A NAND3X1_6/Y gnd OAI21X1_55/C vdd NAND2X1
XOAI21X1_190 INVX4_5/Y INVX4_6/Y OAI21X1_190/C gnd OAI21X1_191/B vdd OAI21X1
XNAND2X1_65 NAND2X1_65/A NAND3X1_8/Y gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_32 INVX1_4/A NAND3X1_4/Y gnd OAI21X1_33/C vdd NAND2X1
XNAND2X1_98 NAND2X1_98/A NAND2X1_98/B gnd AOI21X1_7/B vdd NAND2X1
XNAND2X1_87 INVX1_36/A NAND2X1_83/B gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_10 MUX2X1_19/B NAND2X1_8/B gnd OAI21X1_11/C vdd NAND2X1
XNAND2X1_21 MUX2X1_53/B NAND3X1_2/Y gnd NAND2X1_21/Y vdd NAND2X1
XNAND2X1_76 MUX2X1_44/B NAND3X1_9/Y gnd OAI21X1_77/C vdd NAND2X1
XNAND2X1_43 NAND2X1_43/A NAND3X1_5/Y gnd OAI21X1_44/C vdd NAND2X1
XOAI22X1_3 INVX1_13/Y OR2X2_3/B INVX4_3/A INVX1_12/Y gnd OAI22X1_3/Y vdd OAI22X1
XFILL_20_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XOAI21X1_19 BUFX4_3/Y NAND3X1_2/Y NAND2X1_18/Y gnd OAI21X1_19/Y vdd OAI21X1
XFILL_3_2_0 gnd vdd FILL
XDFFPOSX1_169 MUX2X1_35/B CLKBUF1_4/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 MUX2X1_69/B CLKBUF1_10/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 INVX1_12/A CLKBUF1_5/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XNAND2X1_217 NAND2X1_147/B NAND3X1_29/Y gnd NAND2X1_217/Y vdd NAND2X1
XDFFPOSX1_125 NAND2X1_44/A CLKBUF1_7/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 MUX2X1_73/A CLKBUF1_5/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XNAND2X1_206 MUX2X1_48/A NAND3X1_28/Y gnd OAI21X1_264/C vdd NAND2X1
XDFFPOSX1_147 NAND2X1_66/A CLKBUF1_14/Y OAI21X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 INVX1_37/A CLKBUF1_2/Y OAI21X1_78/Y gnd vdd DFFPOSX1
XBUFX4_52 BUFX4_50/A gnd BUFX4_52/Y vdd BUFX4
XBUFX4_63 INVX8_3/Y gnd BUFX4_63/Y vdd BUFX4
XBUFX4_41 BUFX4_42/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 INVX8_6/Y gnd BUFX4_30/Y vdd BUFX4
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XINVX8_11 BUFX4_35/Y gnd NOR2X1_1/B vdd INVX8
XFILL_0_0_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XMUX2X1_18 MUX2X1_16/Y MUX2X1_18/B OR2X2_4/B gnd MUX2X1_18/Y vdd MUX2X1
XMUX2X1_29 MUX2X1_29/A MUX2X1_29/B BUFX4_17/Y gnd MUX2X1_29/Y vdd MUX2X1
XNAND2X1_22 MUX2X1_69/B NAND3X1_2/Y gnd OAI21X1_23/C vdd NAND2X1
XNAND2X1_99 BUFX4_17/Y NAND2X1_99/B gnd NAND2X1_99/Y vdd NAND2X1
XNAND2X1_88 MUX2X1_67/B NAND2X1_83/B gnd NAND2X1_88/Y vdd NAND2X1
XFILL_14_3_1 gnd vdd FILL
XOAI21X1_191 NAND3X1_20/Y OAI21X1_191/B NAND3X1_19/Y gnd AOI21X1_24/B vdd OAI21X1
XNAND2X1_33 INVX1_12/A NAND3X1_4/Y gnd OAI21X1_34/C vdd NAND2X1
XAOI22X1_1 AOI22X1_1/A NOR2X1_9/Y INVX4_10/Y AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_44 NAND2X1_44/A NAND3X1_5/Y gnd OAI21X1_45/C vdd NAND2X1
XNAND2X1_55 MUX2X1_73/A NAND3X1_6/Y gnd OAI21X1_56/C vdd NAND2X1
XOAI21X1_180 INVX1_37/Y MUX2X1_7/S OAI21X1_180/C gnd OAI21X1_180/Y vdd OAI21X1
XNAND2X1_11 MUX2X1_28/B NAND2X1_8/B gnd OAI21X1_12/C vdd NAND2X1
XNAND2X1_66 NAND2X1_66/A NAND3X1_8/Y gnd NAND2X1_66/Y vdd NAND2X1
XNAND2X1_77 INVX1_37/A NAND3X1_9/Y gnd NAND2X1_77/Y vdd NAND2X1
XOAI22X1_4 INVX1_16/Y OR2X2_3/B INVX4_3/A INVX1_15/Y gnd OAI22X1_4/Y vdd OAI22X1
XFILL_20_1_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XDFFPOSX1_137 MUX2X1_2/B CLKBUF1_13/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_159 MUX2X1_66/B CLKBUF1_13/Y OAI21X1_79/Y gnd vdd DFFPOSX1
XNAND2X1_218 INVX4_9/Y INVX8_12/A gnd OAI21X1_291/A vdd NAND2X1
XDFFPOSX1_148 NAND2X1_67/A CLKBUF1_3/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 INVX1_41/A CLKBUF1_5/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XNAND2X1_207 MUX2X1_54/A NAND3X1_28/Y gnd NAND2X1_207/Y vdd NAND2X1
XDFFPOSX1_104 MUX2X1_75/B CLKBUF1_7/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 INVX1_20/A CLKBUF1_14/Y OAI21X1_35/Y gnd vdd DFFPOSX1
XBUFX4_64 INVX8_3/Y gnd BUFX4_64/Y vdd BUFX4
XBUFX4_42 BUFX4_42/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_20 BUFX4_20/A gnd MUX2X1_2/S vdd BUFX4
XBUFX4_53 INVX8_7/Y gnd BUFX4_53/Y vdd BUFX4
XBUFX4_31 INVX8_6/Y gnd BUFX4_31/Y vdd BUFX4
XINVX8_12 INVX8_12/A gnd BUFX4_50/A vdd INVX8
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_56 MUX2X1_2/B NAND3X1_7/Y gnd OAI21X1_57/C vdd NAND2X1
XAOI22X1_2 AOI22X1_2/A NOR2X1_9/Y INVX4_4/Y AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_78 MUX2X1_66/B NAND3X1_9/Y gnd NAND2X1_78/Y vdd NAND2X1
XOAI21X1_192 INVX8_1/Y BUFX2_7/A NOR2X1_12/Y gnd AOI21X1_24/C vdd OAI21X1
XNAND2X1_89 INVX1_48/A NAND2X1_83/B gnd NAND2X1_89/Y vdd NAND2X1
XNAND2X1_45 INVX1_41/A NAND3X1_5/Y gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_67 NAND2X1_67/A NAND3X1_8/Y gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_23 MUX2X1_75/B NAND3X1_2/Y gnd OAI21X1_24/C vdd NAND2X1
XOAI21X1_181 BUFX4_32/Y BUFX4_12/Y OAI21X1_180/Y gnd AOI21X1_20/A vdd OAI21X1
XNAND2X1_12 MUX2X1_38/B NAND2X1_8/B gnd OAI21X1_13/C vdd NAND2X1
XMUX2X1_19 MUX2X1_19/A MUX2X1_19/B MUX2X1_7/S gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_34 INVX1_20/A NAND3X1_4/Y gnd NAND2X1_34/Y vdd NAND2X1
XOAI21X1_170 INVX1_30/Y OR2X2_2/B NAND2X1_124/Y gnd OAI21X1_170/Y vdd OAI21X1
XOAI22X1_5 INVX1_21/Y OR2X2_3/B INVX4_3/A INVX1_20/Y gnd OAI22X1_5/Y vdd OAI22X1
XDFFPOSX1_138 MUX2X1_11/B CLKBUF1_8/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NAND2X1_46/A CLKBUF1_8/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 INVX1_7/A CLKBUF1_3/Y OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 INVX1_28/A CLKBUF1_3/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 INVX1_34/A CLKBUF1_7/Y OAI21X1_69/Y gnd vdd DFFPOSX1
XNAND2X1_208 MUX2X1_70/A NAND3X1_28/Y gnd OAI21X1_266/C vdd NAND2X1
XNAND2X1_219 NOR2X1_20/Y BUFX4_61/Y gnd BUFX4_44/A vdd NAND2X1
XINVX8_1 rw gnd INVX8_1/Y vdd INVX8
XBUFX4_32 BUFX4_33/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_10 BUFX4_9/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_43 BUFX4_42/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 BUFX4_20/A gnd MUX2X1_4/S vdd BUFX4
XBUFX4_65 BUFX4_67/A gnd BUFX4_65/Y vdd BUFX4
XFILL_10_2 gnd vdd FILL
XBUFX4_54 INVX8_7/Y gnd BUFX4_54/Y vdd BUFX4
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_9_1 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_193 INVX1_48/Y MUX2X1_2/S OAI21X1_193/C gnd NAND2X1_148/A vdd OAI21X1
XOAI21X1_182 NAND3X1_17/Y AOI21X1_20/Y NOR2X1_1/B gnd AOI21X1_22/B vdd OAI21X1
XOAI21X1_171 OAI21X1_170/Y OAI22X1_8/Y INVX4_8/A gnd OAI21X1_171/Y vdd OAI21X1
XOAI21X1_160 OAI21X1_159/Y OAI22X1_5/Y INVX4_8/Y gnd OAI21X1_160/Y vdd OAI21X1
XNAND2X1_57 MUX2X1_11/B NAND3X1_7/Y gnd OAI21X1_58/C vdd NAND2X1
XNAND2X1_24 INVX1_7/A NAND3X1_3/Y gnd OAI21X1_25/C vdd NAND2X1
XNAND2X1_46 NAND2X1_46/A NAND3X1_5/Y gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_35 INVX1_28/A NAND3X1_4/Y gnd NAND2X1_35/Y vdd NAND2X1
XNAND2X1_79 INVX1_49/A NAND3X1_9/Y gnd OAI21X1_80/C vdd NAND2X1
XNAND2X1_13 MUX2X1_50/B NAND2X1_8/B gnd OAI21X1_14/C vdd NAND2X1
XNAND2X1_68 INVX1_34/A NAND3X1_8/Y gnd NAND2X1_68/Y vdd NAND2X1
XOAI22X1_6 INVX1_24/Y OR2X2_3/B INVX4_3/A INVX1_23/Y gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_106 INVX1_15/A CLKBUF1_11/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 INVX1_53/A CLKBUF1_5/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 MUX2X1_20/B CLKBUF1_9/Y OAI21X1_59/Y gnd vdd DFFPOSX1
XNAND2X1_209 MUX2X1_76/A NAND3X1_28/Y gnd NAND2X1_209/Y vdd NAND2X1
XDFFPOSX1_117 INVX1_33/A CLKBUF1_7/Y OAI21X1_37/Y gnd vdd DFFPOSX1
XINVX8_2 datain[0] gnd INVX8_2/Y vdd INVX8
XFILL_3_0_0 gnd vdd FILL
XFILL_19_0_0 gnd vdd FILL
XBUFX4_66 BUFX4_67/A gnd INVX4_7/A vdd BUFX4
XBUFX4_44 BUFX4_44/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_11 BUFX4_9/A gnd OR2X2_4/B vdd BUFX4
XBUFX4_33 BUFX4_33/A gnd OR2X2_4/A vdd BUFX4
XBUFX4_55 INVX8_7/Y gnd BUFX4_55/Y vdd BUFX4
XBUFX4_22 BUFX4_20/A gnd INVX4_8/A vdd BUFX4
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_1_3_1 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_150 INVX1_11/Y OR2X2_2/B NAND2X1_105/Y gnd OAI21X1_151/A vdd OAI21X1
XOAI21X1_183 NOR2X1_2/A INVX1_38/Y NAND3X1_18/Y gnd OAI21X1_183/Y vdd OAI21X1
XOAI21X1_172 INVX8_1/Y BUFX2_4/A NOR2X1_12/Y gnd AOI21X1_17/C vdd OAI21X1
XOAI21X1_194 INVX1_49/Y INVX4_8/A OAI21X1_194/C gnd OAI21X1_194/Y vdd OAI21X1
XOAI21X1_161 INVX1_22/Y OR2X2_2/B NAND2X1_115/Y gnd OAI21X1_161/Y vdd OAI21X1
XNAND2X1_14 MUX2X1_60/B NAND2X1_8/B gnd OAI21X1_15/C vdd NAND2X1
XNAND2X1_25 INVX1_15/A NAND3X1_3/Y gnd OAI21X1_26/C vdd NAND2X1
XNAND2X1_69 INVX1_38/A NAND3X1_8/Y gnd OAI21X1_70/C vdd NAND2X1
XNAND2X1_47 INVX1_53/A NAND3X1_5/Y gnd NAND2X1_47/Y vdd NAND2X1
XNAND2X1_58 MUX2X1_20/B NAND3X1_7/Y gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_36 INVX1_33/A NAND3X1_4/Y gnd NAND2X1_36/Y vdd NAND2X1
XOAI22X1_7 INVX1_29/Y OR2X2_3/B INVX4_3/A INVX1_28/Y gnd OAI22X1_7/Y vdd OAI22X1
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XDFFPOSX1_129 MUX2X1_2/A CLKBUF1_13/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 INVX1_23/A CLKBUF1_3/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_118 INVX1_39/A CLKBUF1_11/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XFILL_3_0_1 gnd vdd FILL
XFILL_19_0_1 gnd vdd FILL
XBUFX4_67 BUFX4_67/A gnd BUFX4_67/Y vdd BUFX4
XBUFX4_45 BUFX4_44/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_12 BUFX4_9/A gnd BUFX4_12/Y vdd BUFX4
XBUFX4_34 BUFX4_33/A gnd NOR2X1_8/B vdd BUFX4
XBUFX4_56 INVX8_7/Y gnd BUFX4_56/Y vdd BUFX4
XBUFX4_23 BUFX4_20/A gnd MUX2X1_7/S vdd BUFX4
XNAND2X1_48 MUX2X1_2/A NAND3X1_6/Y gnd OAI21X1_49/C vdd NAND2X1
XNAND2X1_26 INVX1_23/A NAND3X1_3/Y gnd OAI21X1_27/C vdd NAND2X1
XOAI21X1_151 OAI21X1_151/A OAI22X1_3/Y INVX4_8/Y gnd NAND2X1_107/A vdd OAI21X1
XNAND2X1_37 INVX1_39/A NAND3X1_4/Y gnd NAND2X1_37/Y vdd NAND2X1
XOAI21X1_140 NAND3X1_11/Y AOI21X1_6/Y NOR2X1_1/B gnd AOI21X1_8/B vdd OAI21X1
XOAI21X1_184 OAI22X1_9/Y OAI21X1_183/Y INVX4_8/Y gnd OAI21X1_184/Y vdd OAI21X1
XOAI21X1_162 OAI21X1_161/Y OAI22X1_6/Y MUX2X1_2/S gnd NAND2X1_116/B vdd OAI21X1
XNAND2X1_15 MUX2X1_72/B NAND2X1_8/B gnd OAI21X1_16/C vdd NAND2X1
XNAND2X1_59 MUX2X1_29/B NAND3X1_7/Y gnd NAND2X1_59/Y vdd NAND2X1
XNAND2X1_190 MUX2X1_44/A NAND3X1_26/Y gnd NAND2X1_190/Y vdd NAND2X1
XOAI21X1_173 INVX1_33/Y MUX2X1_8/S NAND2X1_126/Y gnd AOI21X1_18/B vdd OAI21X1
XOAI21X1_195 NOR2X1_8/B BUFX4_10/Y OAI21X1_194/Y gnd AOI21X1_25/A vdd OAI21X1
XOAI22X1_8 INVX1_32/Y OR2X2_3/B INVX4_3/A INVX1_31/Y gnd OAI22X1_8/Y vdd OAI22X1
XFILL_19_1 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_3/A vdd MUX2X1
XDFFPOSX1_119 INVX1_45/A CLKBUF1_8/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_108 INVX1_31/A CLKBUF1_1/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XINVX8_4 datain[1] gnd INVX8_4/Y vdd INVX8
XDFFPOSX1_90 MUX2X1_10/B CLKBUF1_13/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XBUFX4_24 INVX8_9/Y gnd BUFX4_24/Y vdd BUFX4
XBUFX4_57 INVX8_4/Y gnd BUFX4_57/Y vdd BUFX4
XBUFX4_68 BUFX4_67/A gnd BUFX4_68/Y vdd BUFX4
XBUFX4_13 BUFX4_9/A gnd MUX2X1_3/S vdd BUFX4
XBUFX4_46 BUFX4_44/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_35 BUFX4_33/A gnd BUFX4_35/Y vdd BUFX4
XFILL_12_2_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XOAI21X1_300 BUFX4_45/Y BUFX4_65/Y NAND2X1_128/B gnd OAI21X1_301/C vdd OAI21X1
XNAND3X1_1 BUFX4_61/Y NAND3X1_7/B INVX4_9/Y gnd NAND2X1_8/B vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XNAND2X1_49 MUX2X1_11/A NAND3X1_6/Y gnd OAI21X1_50/C vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XOAI21X1_130 BUFX4_58/Y NAND2X1_83/B NAND2X1_83/Y gnd OAI21X1_130/Y vdd OAI21X1
XNAND2X1_180 INVX1_40/A NAND3X1_25/Y gnd OAI21X1_224/C vdd NAND2X1
XNAND2X1_38 INVX1_45/A NAND3X1_4/Y gnd OAI21X1_39/C vdd NAND2X1
XOAI21X1_152 INVX1_14/Y OR2X2_2/B NAND2X1_106/Y gnd OAI21X1_152/Y vdd OAI21X1
XOAI21X1_185 OAI22X1_11/Y OAI22X1_10/Y MUX2X1_4/S gnd OAI21X1_185/Y vdd OAI21X1
XFILL_9_2_0 gnd vdd FILL
XOAI21X1_174 INVX1_34/Y BUFX4_18/Y NAND2X1_127/Y gnd AOI22X1_1/A vdd OAI21X1
XOAI21X1_141 INVX1_3/Y OR2X2_2/B NAND2X1_96/Y gnd OAI21X1_141/Y vdd OAI21X1
XNAND2X1_16 MUX2X1_4/B NAND3X1_2/Y gnd OAI21X1_17/C vdd NAND2X1
XNAND2X1_191 DFFPOSX1_38/Q NAND3X1_26/Y gnd OAI21X1_249/C vdd NAND2X1
XNAND2X1_27 INVX1_31/A NAND3X1_3/Y gnd OAI21X1_28/C vdd NAND2X1
XOAI21X1_163 INVX8_1/Y BUFX2_3/A NOR2X1_12/Y gnd AOI21X1_14/C vdd OAI21X1
XOAI21X1_196 NAND3X1_21/Y AOI21X1_25/Y NOR2X1_1/B gnd AOI21X1_27/B vdd OAI21X1
XOAI22X1_9 INVX4_3/A INVX1_39/Y INVX1_40/Y OR2X2_2/B gnd OAI22X1_9/Y vdd OAI22X1
XFILL_19_2 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XDFFPOSX1_109 NAND2X1_28/A CLKBUF1_6/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XFILL_6_0_0 gnd vdd FILL
XBUFX4_25 INVX8_9/Y gnd BUFX4_25/Y vdd BUFX4
XBUFX4_58 INVX8_4/Y gnd BUFX4_58/Y vdd BUFX4
XBUFX4_36 INVX8_2/Y gnd BUFX4_36/Y vdd BUFX4
XBUFX4_14 BUFX4_9/A gnd MUX2X1_9/S vdd BUFX4
XBUFX4_47 BUFX4_44/A gnd OR2X2_1/A vdd BUFX4
XDFFPOSX1_80 INVX1_54/A CLKBUF1_5/Y OAI21X1_307/Y gnd vdd DFFPOSX1
XDFFPOSX1_91 MUX2X1_19/B CLKBUF1_9/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XINVX8_5 datain[2] gnd BUFX4_1/A vdd INVX8
XBUFX4_69 INVX8_8/Y gnd BUFX4_69/Y vdd BUFX4
XFILL_12_2_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XOAI21X1_301 BUFX4_53/Y NAND3X1_30/Y OAI21X1_301/C gnd DFFPOSX1_77/D vdd OAI21X1
XNAND3X1_2 BUFX4_62/Y NAND3X1_2/B INVX4_9/Y gnd NAND3X1_2/Y vdd NAND3X1
XNAND2X1_181 INVX1_47/A NAND3X1_25/Y gnd OAI21X1_225/C vdd NAND2X1
XNAND2X1_17 MUX2X1_13/B NAND3X1_2/Y gnd OAI21X1_18/C vdd NAND2X1
XNAND2X1_192 MUX2X1_66/A NAND3X1_26/Y gnd OAI21X1_250/C vdd NAND2X1
XOAI21X1_153 OAI21X1_152/Y OAI22X1_4/Y BUFX4_18/Y gnd NAND2X1_107/B vdd OAI21X1
XOAI21X1_120 OR2X2_1/Y BUFX4_30/Y OAI21X1_120/C gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_186 INVX8_1/Y BUFX2_6/A NOR2X1_12/Y gnd AOI21X1_22/C vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_175 INVX1_35/Y MUX2X1_2/S NAND2X1_128/Y gnd AOI22X1_1/D vdd OAI21X1
XOAI21X1_142 OAI21X1_141/Y OAI22X1_1/Y INVX4_8/Y gnd NAND2X1_98/A vdd OAI21X1
XOAI21X1_164 INVX1_25/Y INVX4_8/A NAND2X1_117/Y gnd OAI21X1_164/Y vdd OAI21X1
XOAI21X1_131 BUFX4_4/Y NAND2X1_83/B NAND2X1_84/Y gnd OAI21X1_131/Y vdd OAI21X1
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_39 INVX1_51/A NAND3X1_4/Y gnd OAI21X1_40/C vdd NAND2X1
XNAND2X1_170 INVX1_30/A NAND3X1_24/Y gnd NAND2X1_170/Y vdd NAND2X1
XOAI21X1_197 NOR2X1_2/A INVX1_50/Y NAND3X1_22/Y gnd OAI21X1_198/B vdd OAI21X1
XNAND2X1_28 NAND2X1_28/A NAND3X1_3/Y gnd NAND2X1_28/Y vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XFILL_19_3 gnd vdd FILL
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XMUX2X1_3 MUX2X1_3/A MUX2X1_2/Y MUX2X1_3/S gnd MUX2X1_3/Y vdd MUX2X1
XFILL_6_0_1 gnd vdd FILL
XBUFX4_59 INVX8_4/Y gnd BUFX4_59/Y vdd BUFX4
XDFFPOSX1_70 MUX2X1_56/B CLKBUF1_12/Y OAI21X1_287/Y gnd vdd DFFPOSX1
XBUFX4_48 BUFX4_50/A gnd BUFX4_48/Y vdd BUFX4
XBUFX4_26 INVX8_9/Y gnd BUFX4_26/Y vdd BUFX4
XBUFX4_37 INVX8_2/Y gnd BUFX4_37/Y vdd BUFX4
XDFFPOSX1_81 MUX2X1_4/A CLKBUF1_11/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_92 MUX2X1_28/B CLKBUF1_5/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XBUFX4_15 BUFX4_20/A gnd MUX2X1_8/S vdd BUFX4
XINVX8_6 datain[3] gnd INVX8_6/Y vdd INVX8
XOAI21X1_302 BUFX4_44/Y INVX4_7/A INVX1_42/A gnd OAI21X1_303/C vdd OAI21X1
XOAI21X1_110 OAI21X1_98/A BUFX4_25/Y OAI21X1_110/C gnd OAI21X1_110/Y vdd OAI21X1
XOAI21X1_187 INVX1_45/Y MUX2X1_7/S OAI21X1_187/C gnd AOI21X1_23/B vdd OAI21X1
XOAI21X1_132 BUFX4_29/Y NAND2X1_83/B NAND2X1_85/Y gnd OAI21X1_132/Y vdd OAI21X1
XOAI21X1_143 INVX1_6/Y OR2X2_2/B NAND2X1_97/Y gnd OAI21X1_144/A vdd OAI21X1
XNAND3X1_3 BUFX4_64/Y NOR2X1_1/Y INVX4_7/Y gnd NAND3X1_3/Y vdd NAND3X1
XOAI21X1_154 INVX8_1/Y BUFX2_2/A NOR2X1_12/Y gnd AOI21X1_11/C vdd OAI21X1
XOAI21X1_121 BUFX4_46/Y OR2X2_1/B INVX1_35/A gnd OAI21X1_122/C vdd OAI21X1
XOAI21X1_165 INVX1_26/Y MUX2X1_8/S NAND2X1_119/Y gnd OAI21X1_165/Y vdd OAI21X1
XOAI21X1_198 OAI22X1_12/Y OAI21X1_198/B INVX4_8/Y gnd OAI21X1_198/Y vdd OAI21X1
XOAI21X1_176 INVX4_5/Y INVX4_6/Y NAND2X1_129/Y gnd OAI21X1_176/Y vdd OAI21X1
XNAND2X1_160 MUX2X1_19/A NAND3X1_23/Y gnd OAI21X1_204/C vdd NAND2X1
XNAND2X1_29 INVX1_43/A NAND3X1_3/Y gnd OAI21X1_30/C vdd NAND2X1
XNAND2X1_182 INVX1_52/A NAND3X1_25/Y gnd OAI21X1_226/C vdd NAND2X1
XNAND2X1_18 MUX2X1_22/B NAND3X1_2/Y gnd NAND2X1_18/Y vdd NAND2X1
XNAND2X1_171 MUX2X1_37/A NAND3X1_24/Y gnd OAI21X1_214/C vdd NAND2X1
XNAND2X1_193 NAND2X1_149/B NAND3X1_26/Y gnd OAI21X1_251/C vdd NAND2X1
XFILL_10_3_0 gnd vdd FILL
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_4/S gnd MUX2X1_6/A vdd MUX2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XDFFPOSX1_71 MUX2X1_63/B CLKBUF1_12/Y OAI21X1_289/Y gnd vdd DFFPOSX1
XDFFPOSX1_82 NAND2X1_1/A CLKBUF1_10/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 MUX2X1_38/B CLKBUF1_9/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XINVX8_7 datain[4] gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_60 DFFPOSX1_60/Q CLKBUF1_6/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XBUFX4_49 BUFX4_50/A gnd BUFX4_49/Y vdd BUFX4
XFILL_15_2_0 gnd vdd FILL
XBUFX4_27 INVX8_9/Y gnd BUFX4_27/Y vdd BUFX4
XBUFX4_38 INVX8_2/Y gnd BUFX4_38/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XBUFX4_16 BUFX4_20/A gnd BUFX4_16/Y vdd BUFX4
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XOAI21X1_303 BUFX4_72/Y NAND3X1_30/Y OAI21X1_303/C gnd DFFPOSX1_78/D vdd OAI21X1
XFILL_12_0_0 gnd vdd FILL
XBUFX4_1 BUFX4_1/A gnd BUFX4_1/Y vdd BUFX4
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_100 OAI21X1_98/A BUFX4_59/Y OAI21X1_99/Y gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_111 INVX4_2/Y BUFX4_49/Y MUX2X1_79/A gnd OAI21X1_112/C vdd OAI21X1
XOAI21X1_188 INVX1_46/Y BUFX4_17/Y NAND2X1_141/Y gnd AOI22X1_2/A vdd OAI21X1
XOAI21X1_144 OAI21X1_144/A OAI22X1_2/Y BUFX4_16/Y gnd NAND2X1_98/B vdd OAI21X1
XNAND3X1_4 BUFX4_64/Y NOR2X1_1/Y INVX4_9/Y gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_166 NOR2X1_8/B BUFX4_10/Y OAI21X1_165/Y gnd AOI21X1_15/A vdd OAI21X1
XOAI21X1_122 OR2X2_1/Y BUFX4_53/Y OAI21X1_122/C gnd OAI21X1_122/Y vdd OAI21X1
XOAI21X1_199 OAI22X1_14/Y OAI22X1_13/Y MUX2X1_2/S gnd NAND2X1_153/B vdd OAI21X1
XOAI21X1_155 INVX1_17/Y MUX2X1_2/S NAND2X1_108/Y gnd OAI21X1_155/Y vdd OAI21X1
XOAI21X1_133 BUFX4_53/Y NAND2X1_83/B NAND2X1_86/Y gnd OAI21X1_133/Y vdd OAI21X1
XOAI21X1_177 NAND3X1_16/Y OAI21X1_176/Y NAND3X1_15/Y gnd AOI21X1_19/B vdd OAI21X1
XNAND2X1_183 INVX2_2/A INVX2_1/A gnd OR2X2_3/B vdd NAND2X1
XNAND2X1_172 INVX1_44/A NAND3X1_24/Y gnd NAND2X1_172/Y vdd NAND2X1
XNAND2X1_19 MUX2X1_31/B NAND3X1_2/Y gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_194 MUX2X1_5/B NAND3X1_27/Y gnd NAND2X1_194/Y vdd NAND2X1
XNAND2X1_161 MUX2X1_28/A NAND3X1_23/Y gnd OAI21X1_205/C vdd NAND2X1
XNAND2X1_150 INVX4_3/Y MUX2X1_74/Y gnd NAND3X1_21/A vdd NAND2X1
XFILL_5_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XOAI21X1_1 BUFX4_38/Y NAND2X1_5/B OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B INVX4_8/A gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XINVX8_8 datain[5] gnd INVX8_8/Y vdd INVX8
XDFFPOSX1_72 MUX2X1_78/B CLKBUF1_4/Y OAI21X1_291/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 MUX2X1_14/A CLKBUF1_13/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XFILL_15_2_1 gnd vdd FILL
XBUFX4_39 INVX8_2/Y gnd BUFX4_39/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XDFFPOSX1_61 MUX2X1_45/A CLKBUF1_5/Y OAI21X1_272/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 MUX2X1_50/B CLKBUF1_2/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_83 MUX2X1_22/A CLKBUF1_7/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XBUFX4_17 BUFX4_20/A gnd BUFX4_17/Y vdd BUFX4
XBUFX4_28 INVX8_6/Y gnd BUFX4_28/Y vdd BUFX4
XOAI21X1_304 BUFX4_44/Y INVX4_7/A MUX2X1_59/A gnd OAI21X1_305/C vdd OAI21X1
XBUFX4_2 BUFX4_1/A gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XOAI21X1_112 OAI21X1_98/A BUFX4_40/Y OAI21X1_112/C gnd OAI21X1_112/Y vdd OAI21X1
XOAI21X1_101 INVX4_2/Y BUFX4_49/Y MUX2X1_26/A gnd OAI21X1_102/C vdd OAI21X1
XNAND3X1_5 BUFX4_64/Y NOR2X1_2/Y INVX4_7/Y gnd NAND3X1_5/Y vdd NAND3X1
XNAND2X1_173 NAND2X1_173/A NAND3X1_24/Y gnd NAND2X1_173/Y vdd NAND2X1
XNAND2X1_195 MUX2X1_14/B NAND3X1_27/Y gnd OAI21X1_253/C vdd NAND2X1
XOAI21X1_189 INVX1_47/Y MUX2X1_1/S OAI21X1_189/C gnd AOI22X1_2/D vdd OAI21X1
XNAND2X1_140 INVX4_8/A NAND2X1_30/A gnd OAI21X1_187/C vdd NAND2X1
XNAND2X1_184 INVX4_7/Y INVX8_12/A gnd OAI21X1_231/A vdd NAND2X1
XOAI21X1_123 OR2X2_1/A INVX4_9/A NAND3X1_18/C gnd OAI21X1_123/Y vdd OAI21X1
XOAI21X1_178 INVX8_1/Y BUFX2_5/A NOR2X1_12/Y gnd AOI21X1_19/C vdd OAI21X1
XOAI21X1_145 INVX8_1/Y BUFX2_1/A NOR2X1_12/Y gnd AOI21X1_8/C vdd OAI21X1
XOAI21X1_167 NAND3X1_14/Y AOI21X1_15/Y NOR2X1_1/B gnd AOI21X1_17/B vdd OAI21X1
XOAI21X1_134 BUFX4_70/Y NAND2X1_83/B NAND2X1_87/Y gnd OAI21X1_134/Y vdd OAI21X1
XNAND2X1_151 INVX4_4/Y MUX2X1_77/Y gnd NAND3X1_21/B vdd NAND2X1
XNAND2X1_162 MUX2X1_38/A NAND3X1_23/Y gnd NAND2X1_162/Y vdd NAND2X1
XOAI21X1_156 INVX1_18/Y INVX4_8/A NAND2X1_110/Y gnd OAI21X1_156/Y vdd OAI21X1
XFILL_5_2 gnd vdd FILL
XOAI21X1_2 BUFX4_58/Y NAND2X1_5/B NAND2X1_1/Y gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XMUX2X1_6 MUX2X1_6/A MUX2X1_5/Y BUFX4_12/Y gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XINVX8_9 datain[6] gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_95 MUX2X1_60/B CLKBUF1_13/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_73 INVX1_8/A CLKBUF1_3/Y DFFPOSX1_73/D gnd vdd DFFPOSX1
XDFFPOSX1_62 NAND2X1_133/B CLKBUF1_11/Y OAI21X1_273/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 MUX2X1_23/A CLKBUF1_6/Y OAI21X1_262/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 MUX2X1_31/A CLKBUF1_2/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 NAND2X1_149/B CLKBUF1_6/Y OAI21X1_251/Y gnd vdd DFFPOSX1
XBUFX4_18 BUFX4_20/A gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 INVX8_6/Y gnd BUFX4_29/Y vdd BUFX4
XOAI21X1_305 BUFX4_27/Y NAND3X1_30/Y OAI21X1_305/C gnd DFFPOSX1_79/D vdd OAI21X1
XBUFX4_3 BUFX4_1/A gnd BUFX4_3/Y vdd BUFX4
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 BUFX4_61/Y NAND3X1_7/B INVX4_2/A gnd NAND3X1_6/Y vdd NAND3X1
XOAI21X1_102 OAI21X1_98/A BUFX4_1/Y OAI21X1_102/C gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_135 BUFX4_24/Y NAND2X1_83/B NAND2X1_88/Y gnd OAI21X1_135/Y vdd OAI21X1
XNAND2X1_141 BUFX4_16/Y NAND2X1_46/A gnd NAND2X1_141/Y vdd NAND2X1
XOAI21X1_146 INVX1_9/Y BUFX4_18/Y NAND2X1_99/Y gnd NAND2X1_100/A vdd OAI21X1
XFILL_13_3_0 gnd vdd FILL
XNAND2X1_130 INVX4_10/Y MUX2X1_43/Y gnd NAND3X1_16/A vdd NAND2X1
XOAI21X1_124 OR2X2_1/Y BUFX4_71/Y OAI21X1_123/Y gnd OAI21X1_124/Y vdd OAI21X1
XOAI21X1_168 INVX1_27/Y OR2X2_2/B NAND2X1_123/Y gnd OAI21X1_168/Y vdd OAI21X1
XNAND2X1_152 INVX4_10/Y MUX2X1_80/Y gnd NAND3X1_21/C vdd NAND2X1
XOAI21X1_113 BUFX4_46/Y OR2X2_1/B INVX1_5/A gnd OAI21X1_114/C vdd OAI21X1
XOAI21X1_179 INVX1_36/Y MUX2X1_4/S OAI21X1_179/C gnd NAND2X1_134/A vdd OAI21X1
XOAI21X1_157 NOR2X1_8/B BUFX4_9/Y OAI21X1_156/Y gnd AOI21X1_12/A vdd OAI21X1
XNAND2X1_174 INVX1_56/A NAND3X1_24/Y gnd OAI21X1_217/C vdd NAND2X1
XNAND2X1_163 MUX2X1_50/A NAND3X1_23/Y gnd NAND2X1_163/Y vdd NAND2X1
XNAND2X1_185 INVX2_2/Y INVX2_1/Y gnd NOR2X1_2/A vdd NAND2X1
XNAND2X1_196 MUX2X1_23/B NAND3X1_27/Y gnd OAI21X1_254/C vdd NAND2X1
XOAI21X1_3 BUFX4_3/Y NAND2X1_5/B NAND2X1_2/Y gnd OAI21X1_3/Y vdd OAI21X1
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_7/S gnd MUX2X1_9/A vdd MUX2X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_30 MUX2X1_56/A CLKBUF1_12/Y OAI21X1_239/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 MUX2X1_67/A CLKBUF1_10/Y OAI21X1_274/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX1_16/A CLKBUF1_3/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XBUFX4_19 BUFX4_20/A gnd MUX2X1_1/S vdd BUFX4
XDFFPOSX1_96 MUX2X1_72/B CLKBUF1_14/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 NAND2X1_4/A CLKBUF1_7/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 MUX2X1_5/B CLKBUF1_2/Y DFFPOSX1_41/D gnd vdd DFFPOSX1
XDFFPOSX1_52 MUX2X1_32/A CLKBUF1_2/Y OAI21X1_263/Y gnd vdd DFFPOSX1
XFILL_15_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XOAI21X1_306 BUFX4_45/Y BUFX4_65/Y INVX1_54/A gnd OAI21X1_306/Y vdd OAI21X1
XBUFX4_4 BUFX4_1/A gnd BUFX4_4/Y vdd BUFX4
XINVX4_4 OR2X2_2/B gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 BUFX4_62/Y NAND3X1_7/B INVX4_1/A gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_103 INVX4_2/Y BUFX4_50/Y MUX2X1_35/A gnd OAI21X1_104/C vdd OAI21X1
XNAND2X1_164 MUX2X1_60/A NAND3X1_23/Y gnd NAND2X1_164/Y vdd NAND2X1
XNAND2X1_142 BUFX4_18/Y NAND2X1_173/A gnd OAI21X1_189/C vdd NAND2X1
XOAI21X1_125 BUFX4_44/Y BUFX4_8/Y MUX2X1_59/B gnd OAI21X1_126/C vdd OAI21X1
XOAI21X1_147 INVX1_10/Y MUX2X1_2/S OAI21X1_147/C gnd OAI21X1_148/C vdd OAI21X1
XNAND2X1_186 NAND2X1_92/A NAND3X1_26/Y gnd OAI21X1_244/C vdd NAND2X1
XOAI21X1_136 BUFX4_40/Y NAND2X1_83/B NAND2X1_89/Y gnd OAI21X1_136/Y vdd OAI21X1
XOAI21X1_169 OAI21X1_168/Y OAI22X1_7/Y INVX4_8/Y gnd NAND2X1_125/A vdd OAI21X1
XOAI21X1_114 OR2X2_1/Y BUFX4_37/Y OAI21X1_114/C gnd OAI21X1_114/Y vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd dataout[0] vdd BUFX2
XNAND2X1_175 INVX1_3/A NAND3X1_25/Y gnd OAI21X1_219/C vdd NAND2X1
XOAI21X1_158 NAND3X1_13/Y AOI21X1_12/Y NOR2X1_1/B gnd AOI21X1_14/B vdd OAI21X1
XNAND2X1_197 MUX2X1_32/B NAND3X1_27/Y gnd NAND2X1_197/Y vdd NAND2X1
XNAND2X1_131 NOR2X1_9/Y MUX2X1_46/Y gnd NAND3X1_16/B vdd NAND2X1
XNAND2X1_153 OAI21X1_198/Y NAND2X1_153/B gnd AOI21X1_26/B vdd NAND2X1
XNAND2X1_120 INVX4_3/Y MUX2X1_30/Y gnd NAND3X1_14/A vdd NAND2X1
XFILL_13_3_1 gnd vdd FILL
XAOI21X1_1 cas INVX4_5/Y NOR2X1_3/Y gnd AOI21X1_1/Y vdd AOI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_20 AOI21X1_20/A AOI21X1_20/B NOR2X1_2/A gnd AOI21X1_20/Y vdd AOI21X1
XOAI21X1_4 BUFX4_28/Y NAND2X1_5/B OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B MUX2X1_8/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_2_2_1 gnd vdd FILL
XFILL_18_2_1 gnd vdd FILL
XDFFPOSX1_31 MUX2X1_63/A CLKBUF1_8/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_42 MUX2X1_14/B CLKBUF1_10/Y DFFPOSX1_42/D gnd vdd DFFPOSX1
XDFFPOSX1_75 INVX1_24/A CLKBUF1_3/Y DFFPOSX1_75/D gnd vdd DFFPOSX1
XDFFPOSX1_64 NAND2X1_147/B CLKBUF1_1/Y DFFPOSX1_64/D gnd vdd DFFPOSX1
XDFFPOSX1_20 INVX1_27/A CLKBUF1_1/Y DFFPOSX1_20/D gnd vdd DFFPOSX1
XDFFPOSX1_97 MUX2X1_4/B CLKBUF1_11/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_53 MUX2X1_48/A CLKBUF1_11/Y OAI21X1_264/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 NAND2X1_5/A CLKBUF1_2/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XOAI21X1_307 BUFX4_40/Y NAND3X1_30/Y OAI21X1_306/Y gnd OAI21X1_307/Y vdd OAI21X1
XBUFX4_5 BUFX4_6/A gnd OR2X2_1/B vdd BUFX4
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XOAI21X1_104 OAI21X1_98/A BUFX4_29/Y OAI21X1_104/C gnd OAI21X1_104/Y vdd OAI21X1
XNAND2X1_143 INVX4_3/Y MUX2X1_62/Y gnd OAI21X1_190/C vdd NAND2X1
XOAI21X1_126 OR2X2_1/Y BUFX4_27/Y OAI21X1_126/C gnd OAI21X1_126/Y vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd dataout[1] vdd BUFX2
XOAI21X1_148 BUFX4_32/Y BUFX4_12/Y OAI21X1_148/C gnd AOI21X1_9/A vdd OAI21X1
XOAI21X1_137 INVX1_1/Y BUFX4_16/Y NAND2X1_90/Y gnd NAND2X1_91/A vdd OAI21X1
XNAND3X1_8 BUFX4_64/Y NOR2X1_2/Y INVX4_9/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_115 OR2X2_1/A INVX4_9/A INVX1_13/A gnd OAI21X1_116/C vdd OAI21X1
XNAND2X1_121 INVX4_4/Y MUX2X1_33/Y gnd NAND3X1_14/B vdd NAND2X1
XNAND2X1_110 MUX2X1_4/S DFFPOSX1_35/Q gnd NAND2X1_110/Y vdd NAND2X1
XNAND2X1_132 INVX4_4/Y MUX2X1_49/Y gnd NAND3X1_16/C vdd NAND2X1
XOAI21X1_159 INVX1_19/Y OR2X2_2/B NAND2X1_114/Y gnd OAI21X1_159/Y vdd OAI21X1
XNAND2X1_187 DFFPOSX1_34/Q NAND3X1_26/Y gnd OAI21X1_245/C vdd NAND2X1
XNAND2X1_176 INVX1_11/A NAND3X1_25/Y gnd OAI21X1_220/C vdd NAND2X1
XNAND2X1_198 MUX2X1_48/B NAND3X1_27/Y gnd OAI21X1_256/C vdd NAND2X1
XNAND2X1_154 ras en gnd NOR2X1_12/A vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 ras INVX2_2/Y NOR2X1_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XNAND2X1_165 MUX2X1_72/A NAND3X1_23/Y gnd NAND2X1_165/Y vdd NAND2X1
XAOI21X1_21 BUFX4_32/Y AOI21X1_21/B rw gnd AOI21X1_22/A vdd AOI21X1
XAOI21X1_10 BUFX4_32/Y AOI21X1_10/B rw gnd AOI21X1_10/Y vdd AOI21X1
XOAI21X1_5 BUFX4_56/Y NAND2X1_5/B OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XMUX2X1_9 MUX2X1_9/A MUX2X1_8/Y MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XDFFPOSX1_10 INVX1_14/A CLKBUF1_8/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XDFFPOSX1_65 MUX2X1_7/B CLKBUF1_12/Y DFFPOSX1_65/D gnd vdd DFFPOSX1
XDFFPOSX1_32 MUX2X1_78/A CLKBUF1_4/Y OAI21X1_243/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 MUX2X1_13/B CLKBUF1_10/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 INVX1_32/A CLKBUF1_3/Y DFFPOSX1_76/D gnd vdd DFFPOSX1
XDFFPOSX1_87 MUX2X1_69/A CLKBUF1_10/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 MUX2X1_54/A CLKBUF1_11/Y DFFPOSX1_54/D gnd vdd DFFPOSX1
XDFFPOSX1_43 MUX2X1_23/B CLKBUF1_6/Y DFFPOSX1_43/D gnd vdd DFFPOSX1
XDFFPOSX1_21 MUX2X1_37/B CLKBUF1_9/Y DFFPOSX1_21/D gnd vdd DFFPOSX1
XBUFX4_6 BUFX4_6/A gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_200 BUFX2_3/A CLKBUF1_7/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XFILL_0_3_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XOAI21X1_105 INVX4_2/Y BUFX4_52/Y MUX2X1_42/A gnd OAI21X1_106/C vdd OAI21X1
XNAND3X1_9 BUFX4_64/Y NOR2X1_16/Y INVX4_9/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_149 NAND3X1_12/Y AOI21X1_9/Y NOR2X1_1/B gnd AOI21X1_11/B vdd OAI21X1
XOAI21X1_116 OR2X2_1/Y BUFX4_57/Y OAI21X1_116/C gnd OAI21X1_116/Y vdd OAI21X1
XOAI21X1_138 INVX1_2/Y BUFX4_18/Y NAND2X1_92/Y gnd OAI21X1_138/Y vdd OAI21X1
XOAI21X1_127 OR2X2_1/A INVX4_9/A NAND3X1_22/C gnd OAI21X1_128/C vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd dataout[2] vdd BUFX2
XNAND2X1_144 INVX4_10/Y MUX2X1_65/Y gnd NAND3X1_20/A vdd NAND2X1
XNAND2X1_100 NAND2X1_100/A NOR2X1_8/Y gnd AOI21X1_9/B vdd NAND2X1
XNAND2X1_133 MUX2X1_2/S NAND2X1_133/B gnd OAI21X1_179/C vdd NAND2X1
XNAND2X1_122 INVX4_10/Y MUX2X1_36/Y gnd NAND3X1_14/C vdd NAND2X1
XNAND2X1_199 MUX2X1_54/B NAND3X1_27/Y gnd NAND2X1_199/Y vdd NAND2X1
XNAND2X1_155 cas vas gnd NOR2X1_12/B vdd NAND2X1
XAOI21X1_3 ras INVX2_1/Y NOR2X1_5/Y gnd AOI21X1_3/Y vdd AOI21X1
XNAND2X1_166 INVX2_1/A INVX2_2/Y gnd OR2X2_2/B vdd NAND2X1
XNAND2X1_188 DFFPOSX1_35/Q NAND3X1_26/Y gnd OAI21X1_246/C vdd NAND2X1
XNAND2X1_111 INVX4_3/Y MUX2X1_21/Y gnd NAND3X1_13/A vdd NAND2X1
XNAND2X1_177 INVX1_19/A NAND3X1_25/Y gnd NAND2X1_177/Y vdd NAND2X1
XNOR2X1_1 INVX4_3/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XAOI21X1_11 AOI21X1_10/Y AOI21X1_11/B AOI21X1_11/C gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_22 AOI21X1_22/A AOI21X1_22/B AOI21X1_22/C gnd AOI21X1_22/Y vdd AOI21X1
XOAI21X1_6 BUFX4_70/Y NAND2X1_5/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 INVX1_22/A CLKBUF1_14/Y OAI21X1_212/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 MUX2X1_16/B CLKBUF1_4/Y DFFPOSX1_66/D gnd vdd DFFPOSX1
XDFFPOSX1_22 INVX1_40/A CLKBUF1_13/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XDFFPOSX1_33 NAND2X1_92/A CLKBUF1_5/Y OAI21X1_244/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 MUX2X1_70/A CLKBUF1_10/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XDFFPOSX1_88 MUX2X1_75/A CLKBUF1_5/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 NAND2X1_128/B CLKBUF1_1/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_99 MUX2X1_22/B CLKBUF1_9/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 MUX2X1_32/B CLKBUF1_2/Y DFFPOSX1_44/D gnd vdd DFFPOSX1
XFILL_18_0_0 gnd vdd FILL
XBUFX4_7 BUFX4_6/A gnd INVX4_9/A vdd BUFX4
XDFFPOSX1_201 BUFX2_4/A CLKBUF1_11/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XFILL_16_3_1 gnd vdd FILL
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XFILL_0_3_1 gnd vdd FILL
XOAI21X1_106 OAI21X1_98/A BUFX4_54/Y OAI21X1_106/C gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_128 OR2X2_1/Y BUFX4_42/Y OAI21X1_128/C gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_117 BUFX4_46/Y OR2X2_1/B INVX1_21/A gnd OAI21X1_117/Y vdd OAI21X1
XNAND2X1_167 INVX1_6/A NAND3X1_24/Y gnd NAND2X1_167/Y vdd NAND2X1
XNAND2X1_101 MUX2X1_1/S DFFPOSX1_34/Q gnd OAI21X1_147/C vdd NAND2X1
XNAND2X1_145 NOR2X1_9/Y MUX2X1_68/Y gnd NAND3X1_20/B vdd NAND2X1
XNAND2X1_156 rw NOR2X1_12/Y gnd INVX8_3/A vdd NAND2X1
XOAI21X1_139 BUFX4_32/Y OR2X2_4/B OAI21X1_138/Y gnd AOI21X1_6/A vdd OAI21X1
XNAND2X1_123 NAND2X1_67/A NOR2X1_9/Y gnd NAND2X1_123/Y vdd NAND2X1
XNAND2X1_178 INVX1_27/A NAND3X1_25/Y gnd NAND2X1_178/Y vdd NAND2X1
XNAND2X1_134 NAND2X1_134/A NOR2X1_8/Y gnd AOI21X1_20/B vdd NAND2X1
XBUFX2_4 BUFX2_4/A gnd dataout[3] vdd BUFX2
XNAND2X1_189 DFFPOSX1_36/Q NAND3X1_26/Y gnd NAND2X1_189/Y vdd NAND2X1
XAOI21X1_4 vas INVX4_8/Y NOR2X1_6/Y gnd AOI21X1_4/Y vdd AOI21X1
XNAND2X1_112 INVX4_4/Y MUX2X1_24/Y gnd NAND3X1_13/B vdd NAND2X1
XNOR2X1_2 NOR2X1_2/A NOR2X1_1/B gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_23 INVX4_3/Y AOI21X1_23/B NOR2X1_1/B gnd NAND3X1_19/C vdd AOI21X1
XOAI21X1_7 BUFX4_26/Y NAND2X1_5/B NAND2X1_6/Y gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_12 AOI21X1_12/A AOI21X1_12/B NOR2X1_2/A gnd AOI21X1_12/Y vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XDFFPOSX1_89 MUX2X1_1/B CLKBUF1_13/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 INVX1_47/A CLKBUF1_8/Y OAI21X1_225/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 MUX2X1_25/B CLKBUF1_4/Y DFFPOSX1_67/D gnd vdd DFFPOSX1
XDFFPOSX1_34 DFFPOSX1_34/Q CLKBUF1_10/Y OAI21X1_245/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 INVX1_42/A CLKBUF1_4/Y DFFPOSX1_78/D gnd vdd DFFPOSX1
XDFFPOSX1_45 MUX2X1_48/B CLKBUF1_7/Y DFFPOSX1_45/D gnd vdd DFFPOSX1
XDFFPOSX1_56 MUX2X1_76/A CLKBUF1_14/Y DFFPOSX1_56/D gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_12 INVX1_30/A CLKBUF1_14/Y DFFPOSX1_12/D gnd vdd DFFPOSX1
XFILL_18_0_1 gnd vdd FILL
XBUFX4_8 BUFX4_6/A gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_202 BUFX2_5/A CLKBUF1_11/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XOAI21X1_107 INVX4_2/Y BUFX4_50/Y MUX2X1_57/A gnd OAI21X1_107/Y vdd OAI21X1
XNAND2X1_168 INVX1_14/A NAND3X1_24/Y gnd NAND2X1_168/Y vdd NAND2X1
XNAND2X1_102 INVX4_3/Y MUX2X1_12/Y gnd NAND3X1_12/A vdd NAND2X1
XNAND2X1_146 INVX4_4/Y MUX2X1_71/Y gnd NAND3X1_20/C vdd NAND2X1
XNAND2X1_113 INVX4_10/Y MUX2X1_27/Y gnd NAND3X1_13/C vdd NAND2X1
XOAI21X1_129 BUFX4_38/Y NAND2X1_83/B NAND2X1_82/Y gnd OAI21X1_129/Y vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd dataout[4] vdd BUFX2
XNAND2X1_135 INVX4_8/A DFFPOSX1_38/Q gnd OAI21X1_180/C vdd NAND2X1
XOAI21X1_118 OR2X2_1/Y BUFX4_4/Y OAI21X1_117/Y gnd OAI21X1_118/Y vdd OAI21X1
XNAND2X1_157 INVX2_2/A INVX2_1/Y gnd INVX4_3/A vdd NAND2X1
XNAND2X1_179 MUX2X1_37/B NAND3X1_25/Y gnd NAND2X1_179/Y vdd NAND2X1
XNAND2X1_124 NAND2X1_43/A NOR2X1_9/Y gnd NAND2X1_124/Y vdd NAND2X1
XAOI21X1_5 vas INVX4_6/Y NOR2X1_7/Y gnd AOI21X1_5/Y vdd AOI21X1
XAOI21X1_24 INVX8_1/Y AOI21X1_24/B AOI21X1_24/C gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_13 BUFX4_35/Y AOI21X1_13/B rw gnd AOI21X1_13/Y vdd AOI21X1
XNOR2X1_3 cas address[0] gnd NOR2X1_3/Y vdd NOR2X1
XOAI22X1_10 INVX1_42/Y OR2X2_3/B NOR2X1_2/A INVX1_41/Y gnd OAI22X1_10/Y vdd OAI22X1
XOAI21X1_8 BUFX4_42/Y NAND2X1_5/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XOAI21X1_290 BUFX4_51/Y BUFX4_8/Y MUX2X1_78/B gnd OAI21X1_290/Y vdd OAI21X1
XDFFPOSX1_68 MUX2X1_34/B CLKBUF1_12/Y DFFPOSX1_68/D gnd vdd DFFPOSX1
XDFFPOSX1_79 MUX2X1_59/A CLKBUF1_4/Y DFFPOSX1_79/D gnd vdd DFFPOSX1
XDFFPOSX1_57 NAND2X1_90/B CLKBUF1_5/Y OAI21X1_268/Y gnd vdd DFFPOSX1
XDFFPOSX1_46 MUX2X1_54/B CLKBUF1_11/Y DFFPOSX1_46/D gnd vdd DFFPOSX1
XDFFPOSX1_13 MUX2X1_37/A CLKBUF1_9/Y DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_24 INVX1_52/A CLKBUF1_14/Y DFFPOSX1_24/D gnd vdd DFFPOSX1
XDFFPOSX1_35 DFFPOSX1_35/Q CLKBUF1_9/Y OAI21X1_246/Y gnd vdd DFFPOSX1
XFILL_20_2_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_203 BUFX2_6/A CLKBUF1_11/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XINVX4_9 INVX4_9/A gnd INVX4_9/Y vdd INVX4
XNAND2X1_158 MUX2X1_1/A NAND3X1_23/Y gnd OAI21X1_202/C vdd NAND2X1
XOAI21X1_108 OAI21X1_98/A BUFX4_72/Y OAI21X1_107/Y gnd OAI21X1_108/Y vdd OAI21X1
XNAND2X1_103 INVX4_4/Y MUX2X1_15/Y gnd NAND3X1_12/B vdd NAND2X1
XNAND2X1_147 MUX2X1_1/S NAND2X1_147/B gnd OAI21X1_193/C vdd NAND2X1
XOAI21X1_119 BUFX4_46/Y OR2X2_1/B INVX1_29/A gnd OAI21X1_120/C vdd OAI21X1
XBUFX2_6 BUFX2_6/A gnd dataout[5] vdd BUFX2
XNAND2X1_125 NAND2X1_125/A OAI21X1_171/Y gnd AOI21X1_16/B vdd NAND2X1
XNAND2X1_136 INVX4_3/Y MUX2X1_52/Y gnd NAND3X1_17/A vdd NAND2X1
XNAND2X1_169 INVX1_22/A NAND3X1_24/Y gnd OAI21X1_212/C vdd NAND2X1
XNAND2X1_1 NAND2X1_1/A NAND2X1_5/B gnd NAND2X1_1/Y vdd NAND2X1
XNAND2X1_114 NAND2X1_66/A NOR2X1_9/Y gnd NAND2X1_114/Y vdd NAND2X1
XDFFPOSX1_1 MUX2X1_1/A CLKBUF1_13/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_16_1_0 gnd vdd FILL
XAOI21X1_6 AOI21X1_6/A AOI21X1_6/B NOR2X1_2/A gnd AOI21X1_6/Y vdd AOI21X1
XFILL_8_2_0 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_4 ras address[1] gnd NOR2X1_4/Y vdd NOR2X1
XOAI21X1_9 BUFX4_36/Y NAND2X1_8/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_14 AOI21X1_13/Y AOI21X1_14/B AOI21X1_14/C gnd AOI21X1_14/Y vdd AOI21X1
XOAI22X1_11 INVX4_3/A INVX1_43/Y INVX1_44/Y OR2X2_2/B gnd OAI22X1_11/Y vdd OAI22X1
XAOI21X1_25 AOI21X1_25/A AOI21X1_25/B NOR2X1_2/A gnd AOI21X1_25/Y vdd AOI21X1
XOAI21X1_291 OAI21X1_291/A BUFX4_40/Y OAI21X1_290/Y gnd OAI21X1_291/Y vdd OAI21X1
XOAI21X1_280 BUFX4_51/Y BUFX4_8/Y MUX2X1_25/B gnd OAI21X1_281/C vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_25 MUX2X1_7/A CLKBUF1_12/Y OAI21X1_229/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 NAND2X1_99/B CLKBUF1_13/Y OAI21X1_269/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 MUX2X1_41/B CLKBUF1_8/Y DFFPOSX1_69/D gnd vdd DFFPOSX1
XDFFPOSX1_47 MUX2X1_70/B CLKBUF1_10/Y OAI21X1_258/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 DFFPOSX1_36/Q CLKBUF1_7/Y OAI21X1_247/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_44/A CLKBUF1_9/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XFILL_20_2_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XDFFPOSX1_204 BUFX2_7/A CLKBUF1_10/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XOAI21X1_109 INVX4_2/Y BUFX4_48/Y MUX2X1_64/A gnd OAI21X1_110/C vdd OAI21X1
XNAND2X1_159 MUX2X1_10/A NAND3X1_23/Y gnd NAND2X1_159/Y vdd NAND2X1
XNAND2X1_104 INVX4_10/Y MUX2X1_18/Y gnd NAND3X1_12/C vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd dataout[6] vdd BUFX2
XFILL_11_1 gnd vdd FILL
XNAND2X1_148 NAND2X1_148/A NOR2X1_8/Y gnd AOI21X1_25/B vdd NAND2X1
XNAND2X1_137 INVX4_4/Y MUX2X1_55/Y gnd NAND3X1_17/B vdd NAND2X1
XNAND2X1_115 NAND2X1_42/A NOR2X1_9/Y gnd NAND2X1_115/Y vdd NAND2X1
XNAND2X1_126 MUX2X1_7/S NAND2X1_28/A gnd NAND2X1_126/Y vdd NAND2X1
XAOI21X1_7 BUFX4_35/Y AOI21X1_7/B rw gnd AOI21X1_7/Y vdd AOI21X1
XFILL_8_2_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNAND2X1_2 MUX2X1_22/A NAND2X1_5/B gnd NAND2X1_2/Y vdd NAND2X1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XDFFPOSX1_2 MUX2X1_10/A CLKBUF1_13/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 ras address[2] gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_15 AOI21X1_15/A AOI21X1_15/B NOR2X1_2/A gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 BUFX4_35/Y AOI21X1_26/B rw gnd AOI21X1_26/Y vdd AOI21X1
XOAI22X1_12 INVX4_3/A INVX1_51/Y INVX1_52/Y OR2X2_2/B gnd OAI22X1_12/Y vdd OAI22X1
XOAI21X1_281 OAI21X1_291/A BUFX4_1/Y OAI21X1_281/C gnd DFFPOSX1_67/D vdd OAI21X1
XOAI21X1_292 BUFX4_44/Y BUFX4_65/Y INVX1_8/A gnd OAI21X1_293/C vdd OAI21X1
XFILL_5_0_1 gnd vdd FILL
XOAI21X1_270 BUFX4_4/Y NAND3X1_29/Y OAI21X1_270/C gnd DFFPOSX1_59/D vdd OAI21X1
XDFFPOSX1_15 NAND2X1_173/A CLKBUF1_8/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XDFFPOSX1_26 MUX2X1_16/A CLKBUF1_8/Y DFFPOSX1_26/D gnd vdd DFFPOSX1
XDFFPOSX1_48 MUX2X1_76/B CLKBUF1_14/Y DFFPOSX1_48/D gnd vdd DFFPOSX1
XDFFPOSX1_37 MUX2X1_44/A CLKBUF1_7/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XDFFPOSX1_59 NAND2X1_108/B CLKBUF1_1/Y DFFPOSX1_59/D gnd vdd DFFPOSX1
XDFFPOSX1_205 BUFX2_8/A CLKBUF1_7/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XFILL_11_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd dataout[7] vdd BUFX2
XNAND2X1_105 NAND2X1_65/A NOR2X1_9/Y gnd NAND2X1_105/Y vdd NAND2X1
XNAND2X1_138 INVX4_10/Y MUX2X1_58/Y gnd NAND3X1_17/C vdd NAND2X1
XNAND2X1_127 BUFX4_17/Y NAND2X1_44/A gnd NAND2X1_127/Y vdd NAND2X1
XAOI21X1_8 AOI21X1_7/Y AOI21X1_8/B AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XNAND2X1_149 MUX2X1_4/S NAND2X1_149/B gnd OAI21X1_194/C vdd NAND2X1
XNAND2X1_3 MUX2X1_31/A NAND2X1_5/B gnd OAI21X1_4/C vdd NAND2X1
XNAND2X1_116 OAI21X1_160/Y NAND2X1_116/B gnd AOI21X1_13/B vdd NAND2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XNOR2X1_6 vas address[3] gnd NOR2X1_6/Y vdd NOR2X1
XDFFPOSX1_3 MUX2X1_19/A CLKBUF1_9/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XAOI21X1_16 BUFX4_35/Y AOI21X1_16/B rw gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_27 AOI21X1_26/Y AOI21X1_27/B AOI21X1_27/C gnd AOI21X1_27/Y vdd AOI21X1
XOAI22X1_13 INVX1_54/Y OR2X2_3/B NOR2X1_2/A INVX1_53/Y gnd OAI22X1_13/Y vdd OAI22X1
XOAI21X1_90 OAI21X1_94/A BUFX4_54/Y OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XOAI21X1_282 BUFX4_51/Y BUFX4_8/Y MUX2X1_34/B gnd OAI21X1_282/Y vdd OAI21X1
XDFFPOSX1_27 MUX2X1_25/A CLKBUF1_4/Y DFFPOSX1_27/D gnd vdd DFFPOSX1
XOAI21X1_293 BUFX4_39/Y NAND3X1_30/Y OAI21X1_293/C gnd DFFPOSX1_73/D vdd OAI21X1
XOAI21X1_260 BUFX4_38/Y NAND3X1_28/Y OAI21X1_260/C gnd DFFPOSX1_49/D vdd OAI21X1
XDFFPOSX1_16 INVX1_56/A CLKBUF1_14/Y OAI21X1_217/Y gnd vdd DFFPOSX1
XOAI21X1_271 BUFX4_31/Y NAND3X1_29/Y OAI21X1_271/C gnd OAI21X1_271/Y vdd OAI21X1
XDFFPOSX1_38 DFFPOSX1_38/Q CLKBUF1_11/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 MUX2X1_5/A CLKBUF1_2/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNAND2X1_106 NAND2X1_41/A NOR2X1_9/Y gnd NAND2X1_106/Y vdd NAND2X1
XAOI21X1_9 AOI21X1_9/A AOI21X1_9/B NOR2X1_2/A gnd AOI21X1_9/Y vdd AOI21X1
XNAND2X1_139 OAI21X1_184/Y OAI21X1_185/Y gnd AOI21X1_21/B vdd NAND2X1
XNAND2X1_128 MUX2X1_1/S NAND2X1_128/B gnd NAND2X1_128/Y vdd NAND2X1
XNAND2X1_4 NAND2X1_4/A NAND2X1_5/B gnd OAI21X1_5/C vdd NAND2X1
XNAND2X1_117 MUX2X1_4/S DFFPOSX1_60/Q gnd NAND2X1_117/Y vdd NAND2X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNOR2X1_7 vas address[4] gnd NOR2X1_7/Y vdd NOR2X1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XDFFPOSX1_4 MUX2X1_28/A CLKBUF1_6/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XAOI21X1_17 AOI21X1_16/Y AOI21X1_17/B AOI21X1_17/C gnd AOI21X1_17/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI22X1_14 INVX4_3/A INVX1_55/Y INVX1_56/Y OR2X2_2/B gnd OAI22X1_14/Y vdd OAI22X1
XOAI21X1_91 INVX4_1/Y BUFX4_50/Y MUX2X1_57/B gnd OAI21X1_92/C vdd OAI21X1
XOAI21X1_80 BUFX4_41/Y NAND3X1_9/Y OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_283 OAI21X1_291/A BUFX4_29/Y OAI21X1_282/Y gnd DFFPOSX1_68/D vdd OAI21X1
XOAI21X1_261 BUFX4_58/Y NAND3X1_28/Y NAND2X1_203/Y gnd DFFPOSX1_50/D vdd OAI21X1
XOAI21X1_250 BUFX4_27/Y NAND3X1_26/Y OAI21X1_250/C gnd OAI21X1_250/Y vdd OAI21X1
XOAI21X1_294 BUFX4_44/Y INVX4_7/A INVX1_16/A gnd OAI21X1_295/C vdd OAI21X1
XOAI21X1_272 BUFX4_53/Y NAND3X1_29/Y OAI21X1_272/C gnd OAI21X1_272/Y vdd OAI21X1
XDFFPOSX1_28 MUX2X1_34/A CLKBUF1_4/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XDFFPOSX1_39 MUX2X1_66/A CLKBUF1_8/Y OAI21X1_250/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 INVX1_3/A CLKBUF1_1/Y OAI21X1_219/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_19_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND2X1_5 NAND2X1_5/A NAND2X1_5/B gnd OAI21X1_6/C vdd NAND2X1
XNAND2X1_107 NAND2X1_107/A NAND2X1_107/B gnd AOI21X1_10/B vdd NAND2X1
XNAND2X1_118 OAI21X1_164/Y NOR2X1_8/Y gnd AOI21X1_15/B vdd NAND2X1
XNAND2X1_129 INVX4_3/Y MUX2X1_40/Y gnd NAND2X1_129/Y vdd NAND2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XDFFPOSX1_5 MUX2X1_38/A CLKBUF1_9/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XNOR2X1_8 OR2X2_4/B NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 INVX4_3/Y AOI21X1_18/B NOR2X1_1/B gnd AOI21X1_18/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_92 OAI21X1_94/A BUFX4_72/Y OAI21X1_92/C gnd OAI21X1_92/Y vdd OAI21X1
XOAI21X1_81 INVX4_1/Y BUFX4_49/Y MUX2X1_8/B gnd OAI21X1_82/C vdd OAI21X1
XOAI21X1_70 BUFX4_71/Y NAND3X1_8/Y OAI21X1_70/C gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_240 BUFX4_52/Y BUFX4_67/Y MUX2X1_63/A gnd OAI21X1_240/Y vdd OAI21X1
XOAI21X1_284 BUFX4_52/Y BUFX4_6/Y MUX2X1_41/B gnd OAI21X1_285/C vdd OAI21X1
XOAI21X1_295 BUFX4_57/Y NAND3X1_30/Y OAI21X1_295/C gnd DFFPOSX1_74/D vdd OAI21X1
XOAI21X1_273 BUFX4_71/Y NAND3X1_29/Y OAI21X1_273/C gnd OAI21X1_273/Y vdd OAI21X1
XOAI21X1_262 BUFX4_2/Y NAND3X1_28/Y OAI21X1_262/C gnd OAI21X1_262/Y vdd OAI21X1
XOAI21X1_251 BUFX4_41/Y NAND3X1_26/Y OAI21X1_251/C gnd OAI21X1_251/Y vdd OAI21X1
XDFFPOSX1_29 MUX2X1_41/A CLKBUF1_12/Y OAI21X1_237/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 INVX1_11/A CLKBUF1_10/Y OAI21X1_220/Y gnd vdd DFFPOSX1
XNAND2X1_6 MUX2X1_69/A NAND2X1_5/B gnd NAND2X1_6/Y vdd NAND2X1
XNAND2X1_108 MUX2X1_1/S NAND2X1_108/B gnd NAND2X1_108/Y vdd NAND2X1
XNAND2X1_119 MUX2X1_7/S DFFPOSX1_36/Q gnd NAND2X1_119/Y vdd NAND2X1
XMUX2X1_80 MUX2X1_80/A MUX2X1_80/B MUX2X1_9/S gnd MUX2X1_80/Y vdd MUX2X1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XDFFPOSX1_6 MUX2X1_50/A CLKBUF1_2/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 INVX2_2/A INVX2_1/A gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 INVX8_1/Y AOI21X1_19/B AOI21X1_19/C gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_93 INVX4_1/Y BUFX4_48/Y MUX2X1_64/B gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_82 OAI21X1_94/A BUFX4_39/Y OAI21X1_82/C gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_71 BUFX4_27/Y NAND3X1_8/Y OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_60 BUFX4_31/Y NAND3X1_7/Y NAND2X1_59/Y gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_241 OAI21X1_231/A BUFX4_25/Y OAI21X1_240/Y gnd DFFPOSX1_31/D vdd OAI21X1
XOAI21X1_274 BUFX4_24/Y NAND3X1_29/Y OAI21X1_274/C gnd OAI21X1_274/Y vdd OAI21X1
XOAI21X1_230 BUFX4_52/Y BUFX4_67/Y MUX2X1_16/A gnd OAI21X1_231/C vdd OAI21X1
XOAI21X1_285 OAI21X1_291/A BUFX4_54/Y OAI21X1_285/C gnd DFFPOSX1_69/D vdd OAI21X1
XOAI21X1_296 BUFX4_45/Y BUFX4_65/Y INVX1_24/A gnd OAI21X1_297/C vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_263 BUFX4_28/Y NAND3X1_28/Y NAND2X1_205/Y gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_252 BUFX4_38/Y NAND3X1_27/Y NAND2X1_194/Y gnd DFFPOSX1_41/D vdd OAI21X1
XFILL_17_2_0 gnd vdd FILL
XDFFPOSX1_19 INVX1_19/A CLKBUF1_1/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XFILL_14_0_0 gnd vdd FILL
XINVX4_10 OR2X2_3/B gnd INVX4_10/Y vdd INVX4
XFILL_6_1_0 gnd vdd FILL
XNAND3X1_30 BUFX4_61/Y NOR2X1_20/Y INVX4_7/Y gnd NAND3X1_30/Y vdd NAND3X1
XNAND2X1_7 MUX2X1_75/A NAND2X1_5/B gnd OAI21X1_8/C vdd NAND2X1
XNAND2X1_109 OAI21X1_155/Y NOR2X1_8/Y gnd AOI21X1_12/B vdd NAND2X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XMUX2X1_70 MUX2X1_70/A MUX2X1_70/B BUFX4_18/Y gnd MUX2X1_70/Y vdd MUX2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XDFFPOSX1_7 MUX2X1_60/A CLKBUF1_13/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XFILL_12_3_1 gnd vdd FILL
XOAI21X1_94 OAI21X1_94/A BUFX4_25/Y OAI21X1_93/Y gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_83 INVX4_1/Y BUFX4_48/Y MUX2X1_17/B gnd OAI21X1_84/C vdd OAI21X1
XOAI21X1_50 BUFX4_59/Y NAND3X1_6/Y OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 BUFX4_55/Y NAND3X1_7/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_72 BUFX4_41/Y NAND3X1_8/Y OAI21X1_72/C gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_286 BUFX4_52/Y BUFX4_6/Y MUX2X1_56/B gnd OAI21X1_286/Y vdd OAI21X1
XOAI21X1_253 BUFX4_60/Y NAND3X1_27/Y OAI21X1_253/C gnd DFFPOSX1_42/D vdd OAI21X1
XOAI21X1_231 OAI21X1_231/A BUFX4_57/Y OAI21X1_231/C gnd DFFPOSX1_26/D vdd OAI21X1
XOAI21X1_242 BUFX4_51/Y BUFX4_68/Y MUX2X1_78/A gnd OAI21X1_242/Y vdd OAI21X1
XOAI21X1_220 BUFX4_60/Y NAND3X1_25/Y OAI21X1_220/C gnd OAI21X1_220/Y vdd OAI21X1
XOAI21X1_297 BUFX4_1/Y NAND3X1_30/Y OAI21X1_297/C gnd DFFPOSX1_75/D vdd OAI21X1
XOAI21X1_275 BUFX4_42/Y NAND3X1_29/Y NAND2X1_217/Y gnd DFFPOSX1_64/D vdd OAI21X1
XOAI21X1_264 BUFX4_54/Y NAND3X1_28/Y OAI21X1_264/C gnd OAI21X1_264/Y vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XFILL_9_3_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNAND3X1_20 NAND3X1_20/A NAND3X1_20/B NAND3X1_20/C gnd NAND3X1_20/Y vdd NAND3X1
XNOR2X1_20 OR2X2_3/B NOR2X1_1/B gnd NOR2X1_20/Y vdd NOR2X1
XNAND3X1_31 BUFX4_62/Y NAND3X1_2/B INVX4_7/Y gnd NAND2X1_5/B vdd NAND3X1
XNAND2X1_8 MUX2X1_1/B NAND2X1_8/B gnd OAI21X1_9/C vdd NAND2X1
XMUX2X1_60 MUX2X1_60/A MUX2X1_60/B MUX2X1_2/S gnd MUX2X1_60/Y vdd MUX2X1
XMUX2X1_71 MUX2X1_71/A MUX2X1_70/Y MUX2X1_3/S gnd MUX2X1_71/Y vdd MUX2X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XDFFPOSX1_8 MUX2X1_72/A CLKBUF1_6/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XOAI21X1_95 INVX4_1/Y BUFX4_49/Y MUX2X1_79/B gnd OAI21X1_96/C vdd OAI21X1
XOAI21X1_84 OAI21X1_94/A BUFX4_59/Y OAI21X1_84/C gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_210 BUFX4_39/Y NAND3X1_24/Y NAND2X1_167/Y gnd DFFPOSX1_9/D vdd OAI21X1
XOAI21X1_73 BUFX4_38/Y NAND3X1_9/Y NAND2X1_72/Y gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_62 BUFX4_69/Y NAND3X1_7/Y NAND2X1_61/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_51 BUFX4_3/Y NAND3X1_6/Y OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_40 BUFX4_43/Y NAND3X1_4/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_221 BUFX4_4/Y NAND3X1_25/Y NAND2X1_177/Y gnd DFFPOSX1_19/D vdd OAI21X1
XOAI21X1_287 OAI21X1_291/A BUFX4_72/Y OAI21X1_286/Y gnd OAI21X1_287/Y vdd OAI21X1
XOAI21X1_276 BUFX4_50/Y BUFX4_6/Y MUX2X1_7/B gnd OAI21X1_276/Y vdd OAI21X1
XOAI21X1_243 OAI21X1_231/A BUFX4_40/Y OAI21X1_242/Y gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_232 BUFX4_51/Y BUFX4_68/Y MUX2X1_25/A gnd OAI21X1_233/C vdd OAI21X1
XOAI21X1_298 BUFX4_45/Y BUFX4_65/Y INVX1_32/A gnd OAI21X1_299/C vdd OAI21X1
XDFFPOSX1_190 INVX1_1/A CLKBUF1_11/Y OAI21X1_129/Y gnd vdd DFFPOSX1
XOAI21X1_265 BUFX4_70/Y NAND3X1_28/Y NAND2X1_207/Y gnd DFFPOSX1_54/D vdd OAI21X1
XOAI21X1_254 BUFX4_2/Y NAND3X1_27/Y OAI21X1_254/C gnd DFFPOSX1_43/D vdd OAI21X1
XFILL_15_3_0 gnd vdd FILL
XNAND3X1_10 BUFX4_63/Y NOR2X1_16/Y INVX4_1/A gnd NAND2X1_83/B vdd NAND3X1
XNOR2X1_10 INVX4_5/Y INVX4_6/Y gnd BUFX4_33/A vdd NOR2X1
XNAND3X1_21 NAND3X1_21/A NAND3X1_21/B NAND3X1_21/C gnd NAND3X1_21/Y vdd NAND3X1
XMUX2X1_61 MUX2X1_61/A MUX2X1_61/B MUX2X1_4/S gnd MUX2X1_62/B vdd MUX2X1
XNAND2X1_9 MUX2X1_10/B NAND2X1_8/B gnd NAND2X1_9/Y vdd NAND2X1
XMUX2X1_72 MUX2X1_72/A MUX2X1_72/B MUX2X1_7/S gnd MUX2X1_72/Y vdd MUX2X1
XMUX2X1_50 MUX2X1_50/A MUX2X1_50/B MUX2X1_8/S gnd MUX2X1_50/Y vdd MUX2X1
XDFFPOSX1_9 INVX1_6/A CLKBUF1_3/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_63 BUFX4_24/Y NAND3X1_7/Y OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_96 OAI21X1_94/A BUFX4_40/Y OAI21X1_96/C gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_85 INVX4_1/Y BUFX4_49/Y MUX2X1_26/B gnd OAI21X1_86/C vdd OAI21X1
XOAI21X1_41 BUFX4_37/Y NAND3X1_5/Y OAI21X1_41/C gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_74 BUFX4_60/Y NAND3X1_9/Y NAND2X1_73/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_30 BUFX4_69/Y NAND3X1_3/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 BUFX4_31/Y NAND3X1_6/Y OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XDFFPOSX1_180 MUX2X1_64/A CLKBUF1_12/Y OAI21X1_110/Y gnd vdd DFFPOSX1
XOAI21X1_266 BUFX4_26/Y NAND3X1_28/Y OAI21X1_266/C gnd DFFPOSX1_55/D vdd OAI21X1
XOAI21X1_211 BUFX4_59/Y NAND3X1_24/Y NAND2X1_168/Y gnd DFFPOSX1_10/D vdd OAI21X1
XOAI21X1_288 BUFX4_48/Y BUFX4_6/Y MUX2X1_63/B gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_277 OAI21X1_291/A BUFX4_36/Y OAI21X1_276/Y gnd DFFPOSX1_65/D vdd OAI21X1
XDFFPOSX1_191 INVX1_9/A CLKBUF1_10/Y OAI21X1_130/Y gnd vdd DFFPOSX1
XOAI21X1_233 OAI21X1_231/A BUFX4_1/Y OAI21X1_233/C gnd DFFPOSX1_27/D vdd OAI21X1
XOAI21X1_244 BUFX4_39/Y NAND3X1_26/Y OAI21X1_244/C gnd OAI21X1_244/Y vdd OAI21X1
XOAI21X1_299 BUFX4_29/Y NAND3X1_30/Y OAI21X1_299/C gnd DFFPOSX1_76/D vdd OAI21X1
XOAI21X1_222 BUFX4_30/Y NAND3X1_25/Y NAND2X1_178/Y gnd DFFPOSX1_20/D vdd OAI21X1
XOAI21X1_200 INVX8_1/Y BUFX2_8/A NOR2X1_12/Y gnd AOI21X1_27/C vdd OAI21X1
XOAI21X1_255 BUFX4_28/Y NAND3X1_27/Y NAND2X1_197/Y gnd DFFPOSX1_44/D vdd OAI21X1
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XFILL_15_3_1 gnd vdd FILL
XNAND3X1_11 NAND3X1_11/A NAND2X1_94/Y NAND3X1_11/C gnd NAND3X1_11/Y vdd NAND3X1
XNAND3X1_22 INVX2_2/A INVX2_1/A NAND3X1_22/C gnd NAND3X1_22/Y vdd NAND3X1
XNOR2X1_11 INVX4_5/A INVX4_6/A gnd BUFX4_9/A vdd NOR2X1
XMUX2X1_62 MUX2X1_60/Y MUX2X1_62/B MUX2X1_3/S gnd MUX2X1_62/Y vdd MUX2X1
XMUX2X1_40 MUX2X1_38/Y MUX2X1_39/Y BUFX4_9/Y gnd MUX2X1_40/Y vdd MUX2X1
XMUX2X1_51 MUX2X1_51/A MUX2X1_51/B BUFX4_16/Y gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_73 MUX2X1_73/A MUX2X1_73/B MUX2X1_8/S gnd MUX2X1_73/Y vdd MUX2X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XOAI21X1_97 INVX4_2/Y BUFX4_49/Y MUX2X1_8/A gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_86 OAI21X1_94/A BUFX4_1/Y OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_31 BUFX4_24/Y NAND3X1_3/Y NAND2X1_30/Y gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_42 BUFX4_57/Y NAND3X1_5/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_75 BUFX4_2/Y NAND3X1_9/Y NAND2X1_74/Y gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_53 BUFX4_55/Y NAND3X1_6/Y NAND2X1_52/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_20 BUFX4_28/Y NAND3X1_2/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_64 BUFX4_41/Y NAND3X1_7/Y OAI21X1_64/C gnd OAI21X1_64/Y vdd OAI21X1
XDFFPOSX1_170 MUX2X1_42/B CLKBUF1_8/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_181 MUX2X1_79/A CLKBUF1_12/Y OAI21X1_112/Y gnd vdd DFFPOSX1
XOAI21X1_289 OAI21X1_291/A BUFX4_25/Y OAI21X1_288/Y gnd OAI21X1_289/Y vdd OAI21X1
XOAI21X1_278 BUFX4_52/Y BUFX4_6/Y MUX2X1_16/B gnd OAI21X1_279/C vdd OAI21X1
XOAI21X1_234 BUFX4_51/Y BUFX4_68/Y MUX2X1_34/A gnd OAI21X1_235/C vdd OAI21X1
XOAI21X1_201 OR2X2_4/A MUX2X1_9/S MUX2X1_4/S gnd BUFX4_67/A vdd OAI21X1
XOAI21X1_245 BUFX4_60/Y NAND3X1_26/Y OAI21X1_245/C gnd OAI21X1_245/Y vdd OAI21X1
XDFFPOSX1_192 INVX1_17/A CLKBUF1_1/Y OAI21X1_131/Y gnd vdd DFFPOSX1
XOAI21X1_256 BUFX4_54/Y NAND3X1_27/Y OAI21X1_256/C gnd DFFPOSX1_45/D vdd OAI21X1
XOAI21X1_212 BUFX4_2/Y NAND3X1_24/Y OAI21X1_212/C gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_267 BUFX4_41/Y NAND3X1_28/Y NAND2X1_209/Y gnd DFFPOSX1_56/D vdd OAI21X1
XOAI21X1_223 BUFX4_56/Y NAND3X1_25/Y NAND2X1_179/Y gnd DFFPOSX1_21/D vdd OAI21X1
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XNAND3X1_12 NAND3X1_12/A NAND3X1_12/B NAND3X1_12/C gnd NAND3X1_12/Y vdd NAND3X1
XNAND3X1_23 BUFX4_61/Y NAND3X1_7/B INVX4_7/Y gnd NAND3X1_23/Y vdd NAND3X1
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XMUX2X1_63 MUX2X1_63/A MUX2X1_63/B INVX4_8/A gnd MUX2X1_63/Y vdd MUX2X1
XMUX2X1_41 MUX2X1_41/A MUX2X1_41/B MUX2X1_7/S gnd MUX2X1_41/Y vdd MUX2X1
XMUX2X1_52 MUX2X1_50/Y MUX2X1_51/Y BUFX4_12/Y gnd MUX2X1_52/Y vdd MUX2X1
XMUX2X1_30 MUX2X1_30/A MUX2X1_29/Y BUFX4_10/Y gnd MUX2X1_30/Y vdd MUX2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XMUX2X1_74 MUX2X1_72/Y MUX2X1_73/Y BUFX4_10/Y gnd MUX2X1_74/Y vdd MUX2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XOAI21X1_98 OAI21X1_98/A BUFX4_39/Y OAI21X1_97/Y gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_87 INVX4_1/Y BUFX4_49/Y MUX2X1_35/B gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_10 BUFX4_58/Y NAND2X1_8/B NAND2X1_9/Y gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_65 BUFX4_37/Y NAND3X1_8/Y OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_32 BUFX4_43/Y NAND3X1_3/Y OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_54 BUFX4_69/Y NAND3X1_6/Y NAND2X1_53/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_43 BUFX4_4/Y NAND3X1_5/Y NAND2X1_42/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_76 BUFX4_28/Y NAND3X1_9/Y OAI21X1_76/C gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_21 BUFX4_56/Y NAND3X1_2/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_257 BUFX4_70/Y NAND3X1_27/Y NAND2X1_199/Y gnd DFFPOSX1_46/D vdd OAI21X1
XOAI21X1_202 BUFX4_36/Y NAND3X1_23/Y OAI21X1_202/C gnd DFFPOSX1_1/D vdd OAI21X1
XDFFPOSX1_171 MUX2X1_57/B CLKBUF1_12/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XOAI21X1_279 OAI21X1_291/A BUFX4_59/Y OAI21X1_279/C gnd DFFPOSX1_66/D vdd OAI21X1
XOAI21X1_235 OAI21X1_231/A BUFX4_29/Y OAI21X1_235/C gnd DFFPOSX1_28/D vdd OAI21X1
XDFFPOSX1_193 INVX1_25/A CLKBUF1_3/Y OAI21X1_132/Y gnd vdd DFFPOSX1
XOAI21X1_224 BUFX4_72/Y NAND3X1_25/Y OAI21X1_224/C gnd DFFPOSX1_22/D vdd OAI21X1
XOAI21X1_268 BUFX4_39/Y NAND3X1_29/Y OAI21X1_268/C gnd OAI21X1_268/Y vdd OAI21X1
XDFFPOSX1_182 INVX1_5/A CLKBUF1_1/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XDFFPOSX1_160 INVX1_49/A CLKBUF1_6/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XOAI21X1_246 BUFX4_3/Y NAND3X1_26/Y OAI21X1_246/C gnd OAI21X1_246/Y vdd OAI21X1
XOAI21X1_213 BUFX4_31/Y NAND3X1_24/Y NAND2X1_170/Y gnd DFFPOSX1_12/D vdd OAI21X1
XCLKBUF1_11 clk gnd CLKBUF1_11/Y vdd CLKBUF1
XFILL_10_2_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_18_3_0 gnd vdd FILL
XNOR2X1_13 INVX4_3/A OR2X2_4/A gnd NAND3X1_7/B vdd NOR2X1
XNAND3X1_24 BUFX4_63/Y NOR2X1_14/Y INVX4_7/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND3X1_13 NAND3X1_13/A NAND3X1_13/B NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XMUX2X1_64 MUX2X1_64/A MUX2X1_64/B MUX2X1_7/S gnd MUX2X1_65/B vdd MUX2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_42/B MUX2X1_8/S gnd MUX2X1_43/B vdd MUX2X1
XFILL_16_1 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XMUX2X1_75 MUX2X1_75/A MUX2X1_75/B BUFX4_16/Y gnd MUX2X1_77/A vdd MUX2X1
XMUX2X1_53 NAND2X1_5/A MUX2X1_53/B BUFX4_17/Y gnd MUX2X1_55/A vdd MUX2X1
XMUX2X1_20 MUX2X1_20/A MUX2X1_20/B MUX2X1_8/S gnd MUX2X1_20/Y vdd MUX2X1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XMUX2X1_31 MUX2X1_31/A MUX2X1_31/B BUFX4_18/Y gnd MUX2X1_31/Y vdd MUX2X1
XNAND2X1_90 MUX2X1_8/S NAND2X1_90/B gnd NAND2X1_90/Y vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_55 BUFX4_25/Y NAND3X1_6/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_99 INVX4_2/Y BUFX4_48/Y MUX2X1_17/A gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_88 OAI21X1_94/A BUFX4_29/Y OAI21X1_87/Y gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_66 BUFX4_57/Y NAND3X1_8/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_33 BUFX4_37/Y NAND3X1_4/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_11 BUFX4_2/Y NAND2X1_8/B OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_22 BUFX4_70/Y NAND3X1_2/Y NAND2X1_21/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_77 BUFX4_55/Y NAND3X1_9/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_44 BUFX4_30/Y NAND3X1_5/Y OAI21X1_44/C gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_225 BUFX4_25/Y NAND3X1_25/Y OAI21X1_225/C gnd OAI21X1_225/Y vdd OAI21X1
XOAI21X1_236 BUFX4_48/Y BUFX4_67/Y MUX2X1_41/A gnd OAI21X1_237/C vdd OAI21X1
XOAI21X1_203 BUFX4_58/Y NAND3X1_23/Y NAND2X1_159/Y gnd DFFPOSX1_2/D vdd OAI21X1
XOAI21X1_269 BUFX4_58/Y NAND3X1_29/Y NAND2X1_211/Y gnd OAI21X1_269/Y vdd OAI21X1
XOAI21X1_258 BUFX4_26/Y NAND3X1_27/Y OAI21X1_258/C gnd OAI21X1_258/Y vdd OAI21X1
XOAI21X1_247 BUFX4_28/Y NAND3X1_26/Y NAND2X1_189/Y gnd OAI21X1_247/Y vdd OAI21X1
XOAI21X1_214 BUFX4_55/Y NAND3X1_24/Y OAI21X1_214/C gnd DFFPOSX1_13/D vdd OAI21X1
XDFFPOSX1_172 MUX2X1_64/B CLKBUF1_12/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_183 INVX1_13/A CLKBUF1_5/Y OAI21X1_116/Y gnd vdd DFFPOSX1
XDFFPOSX1_150 INVX1_38/A CLKBUF1_5/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XNAND2X1_220 MUX2X1_4/A NAND2X1_5/B gnd OAI21X1_1/C vdd NAND2X1
XDFFPOSX1_161 INVX4_5/A CLKBUF1_9/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XFILL_4_0_0 gnd vdd FILL
XDFFPOSX1_194 MUX2X1_45/B CLKBUF1_6/Y OAI21X1_133/Y gnd vdd DFFPOSX1
XCLKBUF1_12 clk gnd CLKBUF1_12/Y vdd CLKBUF1
XFILL_4_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_14 OR2X2_2/B NOR2X1_1/B gnd NOR2X1_14/Y vdd NOR2X1
XNAND3X1_25 BUFX4_63/Y NOR2X1_14/Y INVX4_9/Y gnd NAND3X1_25/Y vdd NAND3X1
XNAND3X1_14 NAND3X1_14/A NAND3X1_14/B NAND3X1_14/C gnd NAND3X1_14/Y vdd NAND3X1
XMUX2X1_10 MUX2X1_10/A MUX2X1_10/B MUX2X1_4/S gnd MUX2X1_12/A vdd MUX2X1
XFILL_16_2 gnd vdd FILL
XMUX2X1_65 MUX2X1_63/Y MUX2X1_65/B OR2X2_4/B gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_43 MUX2X1_41/Y MUX2X1_43/B OR2X2_4/B gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_54 MUX2X1_54/A MUX2X1_54/B BUFX4_18/Y gnd MUX2X1_55/B vdd MUX2X1
XMUX2X1_76 MUX2X1_76/A MUX2X1_76/B BUFX4_17/Y gnd MUX2X1_76/Y vdd MUX2X1
XMUX2X1_21 MUX2X1_19/Y MUX2X1_20/Y BUFX4_9/Y gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_32 MUX2X1_32/A MUX2X1_32/B MUX2X1_1/S gnd MUX2X1_33/B vdd MUX2X1
XNAND2X1_80 INVX8_12/A INVX4_1/A gnd OAI21X1_94/A vdd NAND2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XNAND2X1_91 NAND2X1_91/A NOR2X1_8/Y gnd AOI21X1_6/B vdd NAND2X1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_23 BUFX4_26/Y NAND3X1_2/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_34 BUFX4_57/Y NAND3X1_4/Y OAI21X1_34/C gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 BUFX4_53/Y NAND3X1_5/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_12 BUFX4_31/Y NAND2X1_8/B OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_89 INVX4_1/Y BUFX4_48/Y MUX2X1_42/B gnd OAI21X1_90/C vdd OAI21X1
XOAI21X1_237 OAI21X1_231/A BUFX4_54/Y OAI21X1_237/C gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_56 BUFX4_42/Y NAND3X1_6/Y OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_204 BUFX4_3/Y NAND3X1_23/Y OAI21X1_204/C gnd DFFPOSX1_3/D vdd OAI21X1
XOAI21X1_226 BUFX4_43/Y NAND3X1_25/Y OAI21X1_226/C gnd DFFPOSX1_24/D vdd OAI21X1
XOAI21X1_215 BUFX4_69/Y NAND3X1_24/Y NAND2X1_172/Y gnd DFFPOSX1_14/D vdd OAI21X1
XOAI21X1_67 BUFX4_4/Y NAND3X1_8/Y NAND2X1_66/Y gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_78 BUFX4_70/Y NAND3X1_9/Y NAND2X1_77/Y gnd OAI21X1_78/Y vdd OAI21X1
XDFFPOSX1_173 MUX2X1_79/B CLKBUF1_4/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_151 INVX1_46/A CLKBUF1_4/Y OAI21X1_71/Y gnd vdd DFFPOSX1
XNAND2X1_210 NAND2X1_90/B NAND3X1_29/Y gnd OAI21X1_268/C vdd NAND2X1
XDFFPOSX1_195 INVX1_36/A CLKBUF1_11/Y OAI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 INVX2_2/A CLKBUF1_6/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_140 MUX2X1_29/B CLKBUF1_6/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XFILL_4_0_1 gnd vdd FILL
XOAI21X1_259 BUFX4_41/Y NAND3X1_27/Y NAND2X1_201/Y gnd DFFPOSX1_48/D vdd OAI21X1
XOAI21X1_248 BUFX4_56/Y NAND3X1_26/Y NAND2X1_190/Y gnd DFFPOSX1_37/D vdd OAI21X1
XDFFPOSX1_184 INVX1_21/A CLKBUF1_1/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XCLKBUF1_13 clk gnd CLKBUF1_13/Y vdd CLKBUF1
XNOR2X1_15 NOR2X1_15/A INVX8_3/A gnd INVX8_12/A vdd NOR2X1
XNAND3X1_26 BUFX4_63/Y NOR2X1_16/Y INVX4_7/Y gnd NAND3X1_26/Y vdd NAND3X1
XNAND3X1_15 OR2X2_2/Y AOI22X1_1/Y AOI21X1_18/Y gnd NAND3X1_15/Y vdd NAND3X1
XMUX2X1_11 MUX2X1_11/A MUX2X1_11/B INVX4_8/A gnd MUX2X1_11/Y vdd MUX2X1
XMUX2X1_66 MUX2X1_66/A MUX2X1_66/B MUX2X1_8/S gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B BUFX4_12/Y gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_77 MUX2X1_77/A MUX2X1_76/Y BUFX4_10/Y gnd MUX2X1_77/Y vdd MUX2X1
XMUX2X1_22 MUX2X1_22/A MUX2X1_22/B BUFX4_16/Y gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_44 MUX2X1_44/A MUX2X1_44/B BUFX4_16/Y gnd MUX2X1_44/Y vdd MUX2X1
XMUX2X1_33 MUX2X1_31/Y MUX2X1_33/B BUFX4_12/Y gnd MUX2X1_33/Y vdd MUX2X1
XNAND2X1_81 INVX8_12/A INVX4_2/A gnd OAI21X1_98/A vdd NAND2X1
XNAND2X1_70 INVX1_46/A NAND3X1_8/Y gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_92 NAND2X1_92/A BUFX4_17/Y gnd NAND2X1_92/Y vdd NAND2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XFILL_21_1 gnd vdd FILL
XOAI21X1_57 BUFX4_36/Y NAND3X1_7/Y OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_79 BUFX4_26/Y NAND3X1_9/Y NAND2X1_78/Y gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_68 BUFX4_30/Y NAND3X1_8/Y NAND2X1_67/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_46 BUFX4_71/Y NAND3X1_5/Y NAND2X1_45/Y gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_24 BUFX4_42/Y NAND3X1_2/Y OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_13 BUFX4_55/Y NAND2X1_8/B OAI21X1_13/C gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_35 BUFX4_2/Y NAND3X1_4/Y NAND2X1_34/Y gnd OAI21X1_35/Y vdd OAI21X1
XDFFPOSX1_174 MUX2X1_8/A CLKBUF1_4/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XOAI21X1_238 BUFX4_50/Y BUFX4_67/Y MUX2X1_56/A gnd OAI21X1_239/C vdd OAI21X1
XOAI21X1_216 BUFX4_24/Y NAND3X1_24/Y NAND2X1_173/Y gnd DFFPOSX1_15/D vdd OAI21X1
XNAND2X1_211 NAND2X1_99/B NAND3X1_29/Y gnd NAND2X1_211/Y vdd NAND2X1
XDFFPOSX1_130 MUX2X1_11/A CLKBUF1_8/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_196 MUX2X1_67/B CLKBUF1_8/Y OAI21X1_135/Y gnd vdd DFFPOSX1
XOAI21X1_227 INVX4_5/Y INVX4_6/Y INVX4_10/Y gnd NOR2X1_15/A vdd OAI21X1
XNAND2X1_200 MUX2X1_70/B NAND3X1_27/Y gnd OAI21X1_258/C vdd NAND2X1
XDFFPOSX1_185 INVX1_29/A CLKBUF1_1/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XOAI21X1_249 BUFX4_71/Y NAND3X1_26/Y OAI21X1_249/C gnd DFFPOSX1_38/D vdd OAI21X1
XDFFPOSX1_141 MUX2X1_39/B CLKBUF1_9/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_163 INVX2_1/A CLKBUF1_6/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 INVX1_50/A CLKBUF1_14/Y OAI21X1_72/Y gnd vdd DFFPOSX1
XOAI21X1_205 BUFX4_31/Y NAND3X1_23/Y OAI21X1_205/C gnd DFFPOSX1_4/D vdd OAI21X1
XCLKBUF1_14 clk gnd CLKBUF1_14/Y vdd CLKBUF1
XFILL_13_2_0 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XNAND3X1_27 BUFX4_62/Y NAND3X1_2/B INVX4_1/A gnd NAND3X1_27/Y vdd NAND3X1
XNOR2X1_16 NOR2X1_2/A OR2X2_4/A gnd NOR2X1_16/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNAND3X1_16 NAND3X1_16/A NAND3X1_16/B NAND3X1_16/C gnd NAND3X1_16/Y vdd NAND3X1
XMUX2X1_12 MUX2X1_12/A MUX2X1_11/Y MUX2X1_3/S gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_56 MUX2X1_56/A MUX2X1_56/B MUX2X1_1/S gnd MUX2X1_58/A vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B MUX2X1_2/S gnd MUX2X1_34/Y vdd MUX2X1
XMUX2X1_67 MUX2X1_67/A MUX2X1_67/B BUFX4_16/Y gnd MUX2X1_68/B vdd MUX2X1
XMUX2X1_78 MUX2X1_78/A MUX2X1_78/B BUFX4_18/Y gnd MUX2X1_80/A vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XMUX2X1_23 MUX2X1_23/A MUX2X1_23/B BUFX4_17/Y gnd MUX2X1_23/Y vdd MUX2X1
XMUX2X1_45 MUX2X1_45/A MUX2X1_45/B BUFX4_17/Y gnd MUX2X1_46/B vdd MUX2X1
XNAND2X1_93 INVX4_3/Y MUX2X1_3/Y gnd NAND3X1_11/A vdd NAND2X1
XNAND2X1_82 INVX1_1/A NAND2X1_83/B gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_60 MUX2X1_39/B NAND3X1_7/Y gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_71 INVX1_50/A NAND3X1_8/Y gnd OAI21X1_72/C vdd NAND2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_58 BUFX4_59/Y NAND3X1_7/Y OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_25 BUFX4_37/Y NAND3X1_3/Y OAI21X1_25/C gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_47 BUFX4_27/Y NAND3X1_5/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_36 BUFX4_30/Y NAND3X1_4/Y NAND2X1_35/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_14 BUFX4_69/Y NAND2X1_8/B OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_69 BUFX4_56/Y NAND3X1_8/Y NAND2X1_68/Y gnd OAI21X1_69/Y vdd OAI21X1
XDFFPOSX1_175 MUX2X1_17/A CLKBUF1_12/Y OAI21X1_100/Y gnd vdd DFFPOSX1
XOAI21X1_239 OAI21X1_231/A BUFX4_72/Y OAI21X1_239/C gnd OAI21X1_239/Y vdd OAI21X1
XOAI21X1_228 BUFX4_50/Y BUFX4_68/Y MUX2X1_7/A gnd OAI21X1_228/Y vdd OAI21X1
XDFFPOSX1_197 INVX1_48/A CLKBUF1_4/Y OAI21X1_136/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 INVX1_2/A CLKBUF1_7/Y OAI21X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_186 INVX1_35/A CLKBUF1_1/Y OAI21X1_122/Y gnd vdd DFFPOSX1
XDFFPOSX1_142 MUX2X1_51/B CLKBUF1_9/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XOAI21X1_206 BUFX4_55/Y NAND3X1_23/Y NAND2X1_162/Y gnd DFFPOSX1_5/D vdd OAI21X1
XDFFPOSX1_131 MUX2X1_20/A CLKBUF1_9/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XOAI21X1_217 BUFX4_43/Y NAND3X1_24/Y OAI21X1_217/C gnd OAI21X1_217/Y vdd OAI21X1
XDFFPOSX1_164 BUFX4_20/A CLKBUF1_2/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 INVX1_51/A CLKBUF1_14/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XNAND2X1_201 MUX2X1_76/B NAND3X1_27/Y gnd NAND2X1_201/Y vdd NAND2X1
XNAND2X1_212 NAND2X1_108/B NAND3X1_29/Y gnd OAI21X1_270/C vdd NAND2X1
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_5_3_1 gnd vdd FILL
XFILL_2_1 gnd vdd FILL
XNOR2X1_17 MUX2X1_7/S OR2X2_4/Y gnd INVX4_1/A vdd NOR2X1
XNAND3X1_28 BUFX4_62/Y NAND3X1_2/B INVX4_2/A gnd NAND3X1_28/Y vdd NAND3X1
XNAND3X1_17 NAND3X1_17/A NAND3X1_17/B NAND3X1_17/C gnd NAND3X1_17/Y vdd NAND3X1
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B MUX2X1_4/S gnd MUX2X1_36/B vdd MUX2X1
XMUX2X1_57 MUX2X1_57/A MUX2X1_57/B MUX2X1_2/S gnd MUX2X1_57/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_79 MUX2X1_79/A MUX2X1_79/B MUX2X1_1/S gnd MUX2X1_80/B vdd MUX2X1
XMUX2X1_13 NAND2X1_1/A MUX2X1_13/B MUX2X1_7/S gnd MUX2X1_13/Y vdd MUX2X1
XMUX2X1_68 MUX2X1_66/Y MUX2X1_68/B MUX2X1_3/S gnd MUX2X1_68/Y vdd MUX2X1
XFILL_10_0_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XMUX2X1_24 MUX2X1_22/Y MUX2X1_23/Y BUFX4_9/Y gnd MUX2X1_24/Y vdd MUX2X1
XMUX2X1_46 MUX2X1_44/Y MUX2X1_46/B BUFX4_9/Y gnd MUX2X1_46/Y vdd MUX2X1
XNAND2X1_83 INVX1_9/A NAND2X1_83/B gnd NAND2X1_83/Y vdd NAND2X1
XNAND2X1_94 INVX4_4/Y MUX2X1_6/Y gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_72 INVX1_2/A NAND3X1_9/Y gnd NAND2X1_72/Y vdd NAND2X1
XNAND2X1_61 MUX2X1_51/B NAND3X1_7/Y gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_50 MUX2X1_20/A NAND3X1_6/Y gnd OAI21X1_51/C vdd NAND2X1
XOAI21X1_15 BUFX4_24/Y NAND2X1_8/B OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_26 BUFX4_60/Y NAND3X1_3/Y OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_48 BUFX4_42/Y NAND3X1_5/Y NAND2X1_47/Y gnd OAI21X1_48/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_59 BUFX4_3/Y NAND3X1_7/Y NAND2X1_58/Y gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_37 BUFX4_56/Y NAND3X1_4/Y NAND2X1_36/Y gnd OAI21X1_37/Y vdd OAI21X1
XDFFPOSX1_143 MUX2X1_61/B CLKBUF1_13/Y OAI21X1_63/Y gnd vdd DFFPOSX1
XOAI21X1_229 OAI21X1_231/A BUFX4_36/Y OAI21X1_228/Y gnd OAI21X1_229/Y vdd OAI21X1
XDFFPOSX1_176 MUX2X1_26/A CLKBUF1_3/Y OAI21X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 NAND2X1_40/A CLKBUF1_3/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 INVX1_10/A CLKBUF1_10/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_187 NAND3X1_18/C CLKBUF1_5/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XOAI21X1_218 NOR2X1_8/B BUFX4_10/Y INVX4_8/Y gnd BUFX4_6/A vdd OAI21X1
XDFFPOSX1_198 BUFX2_1/A CLKBUF1_7/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XNAND2X1_202 MUX2X1_5/A NAND3X1_28/Y gnd OAI21X1_260/C vdd NAND2X1
XDFFPOSX1_165 INVX4_6/A CLKBUF1_2/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XOAI21X1_207 BUFX4_69/Y NAND3X1_23/Y NAND2X1_163/Y gnd DFFPOSX1_6/D vdd OAI21X1
XDFFPOSX1_132 MUX2X1_29/A CLKBUF1_14/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_110 INVX1_43/A CLKBUF1_2/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XNAND2X1_213 DFFPOSX1_60/Q NAND3X1_29/Y gnd OAI21X1_271/C vdd NAND2X1
XBUFX4_70 INVX8_8/Y gnd BUFX4_70/Y vdd BUFX4
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XNAND3X1_29 BUFX4_63/Y NOR2X1_16/Y INVX4_2/A gnd NAND3X1_29/Y vdd NAND3X1
XNOR2X1_18 OR2X2_2/B OR2X2_4/A gnd NAND3X1_2/B vdd NOR2X1
XNAND3X1_18 INVX2_2/A INVX2_1/A NAND3X1_18/C gnd NAND3X1_18/Y vdd NAND3X1
XNAND2X1_62 MUX2X1_61/B NAND3X1_7/Y gnd OAI21X1_63/C vdd NAND2X1
XMUX2X1_58 MUX2X1_58/A MUX2X1_57/Y MUX2X1_9/S gnd MUX2X1_58/Y vdd MUX2X1
XMUX2X1_36 MUX2X1_34/Y MUX2X1_36/B MUX2X1_9/S gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_14 MUX2X1_14/A MUX2X1_14/B MUX2X1_8/S gnd MUX2X1_15/B vdd MUX2X1
XNAND2X1_95 INVX4_10/Y MUX2X1_9/Y gnd NAND3X1_11/C vdd NAND2X1
XMUX2X1_25 MUX2X1_25/A MUX2X1_25/B BUFX4_18/Y gnd MUX2X1_27/A vdd MUX2X1
XNAND2X1_40 NAND2X1_40/A NAND3X1_5/Y gnd OAI21X1_41/C vdd NAND2X1
XNAND2X1_73 INVX1_10/A NAND3X1_9/Y gnd NAND2X1_73/Y vdd NAND2X1
XMUX2X1_69 MUX2X1_69/A MUX2X1_69/B BUFX4_17/Y gnd MUX2X1_71/A vdd MUX2X1
XNAND2X1_84 INVX1_17/A NAND2X1_83/B gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_51 MUX2X1_29/A NAND3X1_6/Y gnd OAI21X1_52/C vdd NAND2X1
XMUX2X1_47 NAND2X1_4/A MUX2X1_47/B BUFX4_18/Y gnd MUX2X1_49/A vdd MUX2X1
XFILL_20_3_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XOAI21X1_49 BUFX4_36/Y NAND3X1_6/Y OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_27 BUFX4_1/Y NAND3X1_3/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_38 BUFX4_71/Y NAND3X1_4/Y NAND2X1_37/Y gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_16 BUFX4_43/Y NAND2X1_8/B OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_208 BUFX4_26/Y NAND3X1_23/Y NAND2X1_164/Y gnd DFFPOSX1_7/D vdd OAI21X1
XDFFPOSX1_111 NAND2X1_30/A CLKBUF1_13/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 NAND2X1_41/A CLKBUF1_3/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XOAI21X1_219 BUFX4_37/Y NAND3X1_25/Y OAI21X1_219/C gnd OAI21X1_219/Y vdd OAI21X1
XDFFPOSX1_155 INVX1_18/A CLKBUF1_6/Y OAI21X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 MUX2X1_39/A CLKBUF1_9/Y OAI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 MUX2X1_31/B CLKBUF1_2/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_144 MUX2X1_73/B CLKBUF1_6/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_177 MUX2X1_35/A CLKBUF1_4/Y OAI21X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_166 MUX2X1_8/B CLKBUF1_3/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XNAND2X1_203 MUX2X1_14/A NAND3X1_28/Y gnd NAND2X1_203/Y vdd NAND2X1
XDFFPOSX1_188 MUX2X1_59/B CLKBUF1_4/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_199 BUFX2_2/A CLKBUF1_10/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XFILL_8_3_0 gnd vdd FILL
XNAND2X1_214 MUX2X1_45/A NAND3X1_29/Y gnd OAI21X1_272/C vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XBUFX4_60 INVX8_4/Y gnd BUFX4_60/Y vdd BUFX4
XBUFX4_71 INVX8_8/Y gnd BUFX4_71/Y vdd BUFX4
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XNAND3X1_19 OR2X2_3/Y AOI22X1_2/Y NAND3X1_19/C gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_19 INVX4_8/Y OR2X2_4/Y gnd INVX4_2/A vdd NOR2X1
XMUX2X1_26 MUX2X1_26/A MUX2X1_26/B MUX2X1_1/S gnd MUX2X1_27/B vdd MUX2X1
XMUX2X1_15 MUX2X1_13/Y MUX2X1_15/B MUX2X1_3/S gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_59 MUX2X1_59/A MUX2X1_59/B MUX2X1_8/S gnd OR2X2_3/A vdd MUX2X1
XMUX2X1_48 MUX2X1_48/A MUX2X1_48/B MUX2X1_1/S gnd MUX2X1_49/B vdd MUX2X1
XMUX2X1_37 MUX2X1_37/A MUX2X1_37/B BUFX4_16/Y gnd OR2X2_2/A vdd MUX2X1
XFILL_20_3_1 gnd vdd FILL
XNAND2X1_30 NAND2X1_30/A NAND3X1_3/Y gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_85 INVX1_25/A NAND2X1_83/B gnd NAND2X1_85/Y vdd NAND2X1
XNAND2X1_41 NAND2X1_41/A NAND3X1_5/Y gnd OAI21X1_42/C vdd NAND2X1
XNAND2X1_96 NAND2X1_96/A NOR2X1_9/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_74 INVX1_18/A NAND3X1_9/Y gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_52 MUX2X1_39/A NAND3X1_6/Y gnd NAND2X1_52/Y vdd NAND2X1
XNAND2X1_63 MUX2X1_73/B NAND3X1_7/Y gnd OAI21X1_64/C vdd NAND2X1
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 INVX1_5/Y OR2X2_3/B INVX4_3/A INVX1_4/Y gnd OAI22X1_1/Y vdd OAI22X1
XOAI21X1_39 BUFX4_27/Y NAND3X1_4/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_17 BUFX4_38/Y NAND3X1_2/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 BUFX4_30/Y NAND3X1_3/Y OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XOAI21X1_209 BUFX4_43/Y NAND3X1_23/Y NAND2X1_165/Y gnd DFFPOSX1_8/D vdd OAI21X1
XDFFPOSX1_167 MUX2X1_17/B CLKBUF1_8/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_178 MUX2X1_42/A CLKBUF1_8/Y OAI21X1_106/Y gnd vdd DFFPOSX1
XNAND2X1_215 NAND2X1_133/B NAND3X1_29/Y gnd OAI21X1_273/C vdd NAND2X1
XDFFPOSX1_189 NAND3X1_22/C CLKBUF1_5/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 NAND2X1_96/A CLKBUF1_1/Y OAI21X1_65/Y gnd vdd DFFPOSX1
XFILL_0_2_1 gnd vdd FILL
XNAND2X1_204 MUX2X1_23/A NAND3X1_28/Y gnd OAI21X1_262/C vdd NAND2X1
XDFFPOSX1_112 INVX1_55/A CLKBUF1_14/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 MUX2X1_51/A CLKBUF1_2/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 NAND2X1_42/A CLKBUF1_14/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 INVX1_26/A CLKBUF1_6/Y OAI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 MUX2X1_47/B CLKBUF1_7/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XFILL_16_2_1 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XBUFX4_50 BUFX4_50/A gnd BUFX4_50/Y vdd BUFX4
XBUFX4_61 INVX8_3/Y gnd BUFX4_61/Y vdd BUFX4
XBUFX4_72 INVX8_8/Y gnd BUFX4_72/Y vdd BUFX4
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XMUX2X1_16 MUX2X1_16/A MUX2X1_16/B BUFX4_16/Y gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_27 MUX2X1_27/A MUX2X1_27/B MUX2X1_9/S gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B MUX2X1_4/S gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B BUFX4_9/Y gnd MUX2X1_49/Y vdd MUX2X1
XNAND2X1_97 NAND2X1_40/A NOR2X1_9/Y gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_64 NAND2X1_96/A NAND3X1_8/Y gnd OAI21X1_65/C vdd NAND2X1
XNAND2X1_86 MUX2X1_45/B NAND2X1_83/B gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_31 INVX1_55/A NAND3X1_3/Y gnd OAI21X1_32/C vdd NAND2X1
XNAND2X1_53 MUX2X1_51/A NAND3X1_6/Y gnd NAND2X1_53/Y vdd NAND2X1
XNAND2X1_42 NAND2X1_42/A NAND3X1_5/Y gnd NAND2X1_42/Y vdd NAND2X1
XNAND2X1_75 INVX1_26/A NAND3X1_9/Y gnd OAI21X1_76/C vdd NAND2X1
XNAND2X1_20 MUX2X1_47/B NAND3X1_2/Y gnd OAI21X1_21/C vdd NAND2X1
XOAI22X1_2 INVX1_8/Y OR2X2_3/B INVX4_3/A INVX1_7/Y gnd OAI22X1_2/Y vdd OAI22X1
XOAI21X1_18 BUFX4_60/Y NAND3X1_2/Y OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 BUFX4_53/Y NAND3X1_3/Y NAND2X1_28/Y gnd OAI21X1_29/Y vdd OAI21X1
XDFFPOSX1_135 MUX2X1_61/A CLKBUF1_12/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_179 MUX2X1_57/A CLKBUF1_12/Y OAI21X1_108/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 MUX2X1_26/B CLKBUF1_3/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XNAND2X1_216 MUX2X1_67/A NAND3X1_29/Y gnd OAI21X1_274/C vdd NAND2X1
XDFFPOSX1_146 NAND2X1_65/A CLKBUF1_5/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_113 INVX1_4/A CLKBUF1_1/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_102 MUX2X1_53/B CLKBUF1_2/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 MUX2X1_44/B CLKBUF1_7/Y OAI21X1_77/Y gnd vdd DFFPOSX1
XNAND2X1_205 MUX2X1_32/A NAND3X1_28/Y gnd NAND2X1_205/Y vdd NAND2X1
XDFFPOSX1_124 NAND2X1_43/A CLKBUF1_1/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XBUFX4_51 BUFX4_50/A gnd BUFX4_51/Y vdd BUFX4
XBUFX4_62 INVX8_3/Y gnd BUFX4_62/Y vdd BUFX4
XBUFX4_40 BUFX4_42/A gnd BUFX4_40/Y vdd BUFX4
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XINVX8_10 datain[7] gnd BUFX4_42/A vdd INVX8
.ends

