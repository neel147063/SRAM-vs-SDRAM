* NGSPICE file created from ram32_sram.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt ram32_sram vdd gnd enable clk r_w datain[0] datain[1] datain[2] datain[3]
+ datain[4] datain[5] datain[6] datain[7] address[0] address[1] address[2] address[3]
+ address[4] dataout[0] dataout[1] dataout[2] dataout[3] dataout[4] dataout[5] dataout[6]
+ dataout[7]
XFILL_23_3_0 gnd vdd FILL
XMUX2X1_17 NOR2X1_35/A MUX2X1_17/B MUX2X1_1/S gnd MUX2X1_18/A vdd MUX2X1
XFILL_14_3_0 gnd vdd FILL
XMUX2X1_39 MUX2X1_38/Y MUX2X1_39/B BUFX4_11/Y gnd AOI22X1_7/A vdd MUX2X1
XMUX2X1_28 MUX2X1_28/A MUX2X1_28/B BUFX4_36/Y gnd MUX2X1_28/Y vdd MUX2X1
XNAND2X1_43 NAND2X1_43/A OAI21X1_38/B gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_54 MUX2X1_5/B OAI21X1_52/B gnd NAND2X1_54/Y vdd NAND2X1
XNAND2X1_65 MUX2X1_59/B NAND2X1_65/B gnd OAI21X1_57/C vdd NAND2X1
XOAI21X1_190 BUFX4_57/Y OAI21X1_183/B OAI21X1_190/C gnd DFFPOSX1_8/D vdd OAI21X1
XAOI22X1_30 AOI22X1_30/A AOI22X1_2/B AOI22X1_2/C MUX2X1_180/Y gnd AOI22X1_30/Y vdd
+ AOI22X1
XNAND2X1_10 MUX2X1_32/B OAI21X1_7/B gnd OAI21X1_8/C vdd NAND2X1
XNAND2X1_21 MUX2X1_73/B OAI21X1_18/B gnd OAI21X1_18/C vdd NAND2X1
XNAND2X1_87 MUX2X1_163/A NAND2X1_88/B gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_76 NAND2X1_76/A NAND2X1_79/B gnd NAND2X1_76/Y vdd NAND2X1
XNAND2X1_98 AND2X2_2/B NOR2X1_2/Y gnd OAI21X1_90/B vdd NAND2X1
XNAND2X1_32 MUX2X1_127/B NAND2X1_27/B gnd OAI21X1_28/C vdd NAND2X1
XFILL_20_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 BUFX4_3/Y OAI21X1_18/B NAND2X1_22/Y gnd OAI21X1_19/Y vdd OAI21X1
XDFFPOSX1_169 MUX2X1_22/B CLKBUF1_23/A OAI21X1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_147 MUX2X1_67/A CLKBUF1_22/Y OAI21X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 MUX2X1_179/B CLKBUF1_4/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XNAND2X1_228 MUX2X1_79/A OAI21X1_183/B gnd OAI21X1_186/C vdd NAND2X1
XFILL_12_3 gnd vdd FILL
XDFFPOSX1_114 MUX2X1_28/A CLKBUF1_25/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XNAND2X1_206 r_w BUFX2_4/A gnd AOI21X1_28/A vdd NAND2X1
XDFFPOSX1_158 MUX2X1_140/B CLKBUF1_43/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XNAND2X1_239 MUX2X1_130/A OAI21X1_193/B gnd OAI21X1_196/C vdd NAND2X1
XNAND2X1_217 AOI22X1_27/Y AOI22X1_28/Y gnd OAI21X1_181/B vdd NAND2X1
XDFFPOSX1_125 NAND2X1_58/A CLKBUF1_35/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 NOR2X1_17/A CLKBUF1_6/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XBUFX4_52 INVX8_2/Y gnd BUFX4_52/Y vdd BUFX4
XBUFX4_41 INVX8_7/Y gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 address[0] gnd MUX2X1_2/S vdd BUFX4
XFILL_0_0_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XMUX2X1_18 MUX2X1_18/A MUX2X1_16/Y BUFX4_12/Y gnd AOI22X1_3/D vdd MUX2X1
XMUX2X1_29 MUX2X1_29/A MUX2X1_29/B BUFX4_37/Y gnd MUX2X1_30/A vdd MUX2X1
XNAND2X1_88 MUX2X1_187/A NAND2X1_88/B gnd OAI21X1_78/C vdd NAND2X1
XNAND2X1_11 MUX2X1_56/B OAI21X1_7/B gnd OAI21X1_9/C vdd NAND2X1
XAOI22X1_1 MUX2X1_3/Y NOR2X1_2/Y AOI22X1_9/C MUX2X1_6/Y gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_99 MUX2X1_1/A OAI21X1_90/B gnd OAI21X1_87/C vdd NAND2X1
XOAI21X1_191 BUFX4_19/Y OAI21X1_193/B OAI21X1_191/C gnd DFFPOSX1_9/D vdd OAI21X1
XFILL_14_3_1 gnd vdd FILL
XNAND2X1_55 MUX2X1_29/B OAI21X1_52/B gnd OAI21X1_48/C vdd NAND2X1
XNAND2X1_77 NAND2X1_77/A NAND2X1_79/B gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_44 AND2X2_2/B AOI22X1_9/C gnd NAND2X1_50/B vdd NAND2X1
XNAND2X1_66 MUX2X1_83/B NAND2X1_65/B gnd OAI21X1_58/C vdd NAND2X1
XOAI21X1_180 NAND2X1_213/Y OAI21X1_180/B INVX4_2/Y gnd AOI21X1_30/B vdd OAI21X1
XNAND2X1_33 NAND2X1_33/A NAND2X1_27/B gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_22 MUX2X1_97/B OAI21X1_18/B gnd NAND2X1_22/Y vdd NAND2X1
XAOI22X1_31 AOI22X1_31/A AOI22X1_3/B INVX8_9/Y AOI22X1_31/D gnd AOI22X1_31/Y vdd AOI22X1
XAOI22X1_20 AOI22X1_20/A AOI22X1_4/B AOI22X1_4/C MUX2X1_120/Y gnd AOI22X1_20/Y vdd
+ AOI22X1
XFILL_20_1_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XDFFPOSX1_137 MUX2X1_19/B CLKBUF1_32/A OAI21X1_63/Y gnd vdd DFFPOSX1
XNAND2X1_218 r_w BUFX2_8/A gnd AOI21X1_32/A vdd NAND2X1
XDFFPOSX1_104 NOR2X1_18/A CLKBUF1_2/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_115 MUX2X1_52/A CLKBUF1_21/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 MUX2X1_91/A CLKBUF1_17/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XNAND2X1_207 AOI22X1_13/Y AOI22X1_14/Y gnd NAND2X1_207/Y vdd NAND2X1
XNAND2X1_229 MUX2X1_103/A OAI21X1_183/B gnd NAND2X1_229/Y vdd NAND2X1
XDFFPOSX1_126 MUX2X1_125/B CLKBUF1_9/A OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_159 MUX2X1_164/B CLKBUF1_7/A OAI21X1_85/Y gnd vdd DFFPOSX1
XBUFX4_20 INVX8_1/Y gnd BUFX4_20/Y vdd BUFX4
XBUFX4_53 INVX8_2/Y gnd BUFX4_53/Y vdd BUFX4
XBUFX4_42 INVX8_7/Y gnd BUFX4_42/Y vdd BUFX4
XBUFX4_31 address[0] gnd MUX2X1_4/S vdd BUFX4
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XMUX2X1_19 MUX2X1_19/A MUX2X1_19/B MUX2X1_2/S gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_56 MUX2X1_53/B OAI21X1_52/B gnd OAI21X1_49/C vdd NAND2X1
XOAI21X1_170 BUFX4_49/Y OAI21X1_174/B NAND2X1_192/Y gnd OAI21X1_170/Y vdd OAI21X1
XNAND2X1_45 MUX2X1_4/A NAND2X1_50/B gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_34 MUX2X1_175/B NAND2X1_27/B gnd OAI21X1_30/C vdd NAND2X1
XAOI22X1_2 MUX2X1_9/Y AOI22X1_2/B AOI22X1_2/C MUX2X1_12/Y gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_12 MUX2X1_80/B OAI21X1_7/B gnd OAI21X1_10/C vdd NAND2X1
XOAI21X1_192 BUFX4_54/Y OAI21X1_193/B NAND2X1_235/Y gnd DFFPOSX1_10/D vdd OAI21X1
XNAND2X1_78 MUX2X1_163/B NAND2X1_79/B gnd NAND2X1_78/Y vdd NAND2X1
XNAND2X1_89 AOI22X1_4/B NOR2X1_1/Y gnd NAND2X1_97/B vdd NAND2X1
XNAND2X1_23 MUX2X1_121/B OAI21X1_18/B gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_67 MUX2X1_107/B NAND2X1_65/B gnd NAND2X1_67/Y vdd NAND2X1
XOAI21X1_181 OAI21X1_181/A OAI21X1_181/B INVX4_2/Y gnd AOI21X1_31/B vdd OAI21X1
XAOI22X1_32 AOI22X1_32/A AOI22X1_4/B AOI22X1_4/C AOI22X1_32/D gnd AOI22X1_32/Y vdd
+ AOI22X1
XAOI22X1_10 MUX2X1_57/Y AOI22X1_2/B AOI22X1_2/C MUX2X1_60/Y gnd AOI22X1_10/Y vdd AOI22X1
XAOI22X1_21 MUX2X1_123/Y NOR2X1_2/Y AOI22X1_9/C AOI22X1_21/D gnd AOI22X1_21/Y vdd
+ AOI22X1
XDFFPOSX1_116 MUX2X1_76/A CLKBUF1_19/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 MUX2X1_5/A CLKBUF1_23/A OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 MUX2X1_43/B CLKBUF1_6/A OAI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 MUX2X1_115/A CLKBUF1_15/Y OAI21X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NAND2X1_60/A CLKBUF1_7/A OAI21X1_53/Y gnd vdd DFFPOSX1
XNAND2X1_219 AOI22X1_29/Y AOI22X1_30/Y gnd NAND2X1_219/Y vdd NAND2X1
XNAND2X1_208 AOI22X1_15/Y AOI22X1_16/Y gnd OAI21X1_178/B vdd NAND2X1
XINVX8_1 datain[0] gnd INVX8_1/Y vdd INVX8
XBUFX4_21 INVX8_1/Y gnd BUFX4_21/Y vdd BUFX4
XBUFX4_10 address[1] gnd BUFX4_10/Y vdd BUFX4
XBUFX4_43 INVX8_7/Y gnd BUFX4_43/Y vdd BUFX4
XBUFX4_32 address[0] gnd MUX2X1_5/S vdd BUFX4
XBUFX4_54 INVX8_2/Y gnd BUFX4_54/Y vdd BUFX4
XFILL_9_1 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_193 BUFX4_14/Y OAI21X1_193/B NAND2X1_236/Y gnd DFFPOSX1_11/D vdd OAI21X1
XOAI21X1_182 NAND2X1_219/Y OAI21X1_182/B INVX4_2/Y gnd AOI21X1_32/B vdd OAI21X1
XAOI22X1_3 MUX2X1_15/Y AOI22X1_3/B INVX8_9/Y AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_160 BUFX4_50/Y OAI21X1_162/B OAI21X1_160/C gnd OAI21X1_160/Y vdd OAI21X1
XOAI21X1_171 BUFX4_3/Y OAI21X1_174/B NAND2X1_193/Y gnd OAI21X1_171/Y vdd OAI21X1
XNAND2X1_79 MUX2X1_187/B NAND2X1_79/B gnd OAI21X1_70/C vdd NAND2X1
XAOI22X1_11 MUX2X1_63/Y AOI22X1_3/B INVX8_9/Y MUX2X1_66/Y gnd AOI22X1_11/Y vdd AOI22X1
XNAND2X1_57 MUX2X1_77/B OAI21X1_52/B gnd OAI21X1_50/C vdd NAND2X1
XNAND2X1_46 MUX2X1_28/A NAND2X1_50/B gnd OAI21X1_40/C vdd NAND2X1
XNAND2X1_35 AND2X2_4/B AOI22X1_9/C gnd OAI21X1_38/B vdd NAND2X1
XNAND2X1_68 MUX2X1_131/B NAND2X1_65/B gnd NAND2X1_68/Y vdd NAND2X1
XAOI22X1_22 AOI22X1_22/A AOI22X1_2/B AOI22X1_2/C AOI22X1_22/D gnd AOI22X1_22/Y vdd
+ AOI22X1
XNAND2X1_24 MUX2X1_145/B OAI21X1_18/B gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_13 MUX2X1_104/B OAI21X1_7/B gnd OAI21X1_11/C vdd NAND2X1
XFILL_23_1_0 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_128 MUX2X1_173/B CLKBUF1_1/A OAI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 MUX2X1_67/B CLKBUF1_32/A OAI21X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 MUX2X1_29/A CLKBUF1_31/A OAI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 MUX2X1_100/A CLKBUF1_13/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XNAND2X1_209 r_w BUFX2_5/A gnd AOI21X1_29/A vdd NAND2X1
XINVX8_2 datain[1] gnd INVX8_2/Y vdd INVX8
XFILL_3_0_0 gnd vdd FILL
XBUFX4_55 INVX8_8/Y gnd BUFX4_55/Y vdd BUFX4
XBUFX4_22 INVX8_1/Y gnd BUFX4_22/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_11 address[1] gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 INVX8_7/Y gnd BUFX4_44/Y vdd BUFX4
XBUFX4_33 address[0] gnd MUX2X1_7/S vdd BUFX4
XFILL_1_3_1 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_183 BUFX4_20/Y OAI21X1_183/B NAND2X1_225/Y gnd DFFPOSX1_1/D vdd OAI21X1
XOAI21X1_161 BUFX4_15/Y OAI21X1_162/B NAND2X1_182/Y gnd OAI21X1_161/Y vdd OAI21X1
XAOI22X1_4 AOI22X1_4/A AOI22X1_4/B AOI22X1_4/C AOI22X1_4/D gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_150 BUFX4_57/Y NAND2X1_169/B OAI21X1_150/C gnd OAI21X1_150/Y vdd OAI21X1
XOAI21X1_194 BUFX4_48/Y OAI21X1_193/B NAND2X1_237/Y gnd DFFPOSX1_12/D vdd OAI21X1
XOAI21X1_172 BUFX4_24/Y OAI21X1_174/B OAI21X1_172/C gnd OAI21X1_172/Y vdd OAI21X1
XAOI22X1_12 MUX2X1_69/Y AOI22X1_4/B AOI22X1_4/C MUX2X1_72/Y gnd AOI22X1_12/Y vdd AOI22X1
XNAND2X1_36 MUX2X1_5/A OAI21X1_38/B gnd OAI21X1_31/C vdd NAND2X1
XNAND2X1_47 MUX2X1_52/A NAND2X1_50/B gnd NAND2X1_47/Y vdd NAND2X1
XNAND2X1_14 MUX2X1_128/B OAI21X1_7/B gnd OAI21X1_12/C vdd NAND2X1
XAOI22X1_23 MUX2X1_135/Y AOI22X1_3/B INVX8_9/Y MUX2X1_138/Y gnd AOI22X1_23/Y vdd AOI22X1
XNAND2X1_25 NAND2X1_25/A OAI21X1_18/B gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_58 NAND2X1_58/A OAI21X1_52/B gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_69 MUX2X1_155/B NAND2X1_65/B gnd NAND2X1_69/Y vdd NAND2X1
XFILL_23_1_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XCLKBUF1_1 CLKBUF1_1/A gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_107 MUX2X1_53/A CLKBUF1_2/A OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_129 MUX2X1_11/B CLKBUF1_29/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_118 MUX2X1_124/A CLKBUF1_9/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XINVX8_3 datain[2] gnd INVX8_3/Y vdd INVX8
XFILL_3_0_1 gnd vdd FILL
XBUFX4_56 INVX8_8/Y gnd BUFX4_56/Y vdd BUFX4
XBUFX4_23 INVX8_1/Y gnd BUFX4_23/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_45 INVX8_4/Y gnd BUFX4_45/Y vdd BUFX4
XBUFX4_12 address[1] gnd BUFX4_12/Y vdd BUFX4
XBUFX4_34 address[0] gnd MUX2X1_8/S vdd BUFX4
XOAI21X1_151 BUFX4_23/Y NAND2X1_173/B OAI21X1_151/C gnd OAI21X1_151/Y vdd OAI21X1
XOAI21X1_184 BUFX4_52/Y OAI21X1_183/B NAND2X1_226/Y gnd DFFPOSX1_2/D vdd OAI21X1
XAOI22X1_5 MUX2X1_27/Y NOR2X1_2/Y AOI22X1_9/C MUX2X1_30/Y gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_190 MUX2X1_26/B OAI21X1_174/B gnd OAI21X1_168/C vdd NAND2X1
XNAND2X1_37 MUX2X1_29/A OAI21X1_38/B gnd OAI21X1_32/C vdd NAND2X1
XNAND2X1_48 MUX2X1_76/A NAND2X1_50/B gnd NAND2X1_48/Y vdd NAND2X1
XAOI22X1_13 MUX2X1_75/Y NOR2X1_2/Y AOI22X1_9/C MUX2X1_78/Y gnd AOI22X1_13/Y vdd AOI22X1
XNAND2X1_26 AOI22X1_2/B NOR2X1_33/Y gnd NAND2X1_27/B vdd NAND2X1
XOAI21X1_195 BUFX4_2/Y OAI21X1_193/B NAND2X1_238/Y gnd DFFPOSX1_13/D vdd OAI21X1
XOAI21X1_162 BUFX4_49/Y OAI21X1_162/B OAI21X1_162/C gnd OAI21X1_162/Y vdd OAI21X1
XAOI22X1_24 AOI22X1_24/A AOI22X1_4/B AOI22X1_4/C MUX2X1_144/Y gnd AOI22X1_24/Y vdd
+ AOI22X1
XOAI21X1_173 BUFX4_41/Y OAI21X1_174/B NAND2X1_195/Y gnd OAI21X1_173/Y vdd OAI21X1
XOAI21X1_140 BUFX4_28/Y NAND2X1_160/B NAND2X1_158/Y gnd OAI21X1_140/Y vdd OAI21X1
XNAND2X1_59 MUX2X1_125/B OAI21X1_52/B gnd OAI21X1_52/C vdd NAND2X1
XNAND2X1_15 MUX2X1_152/B OAI21X1_7/B gnd NAND2X1_15/Y vdd NAND2X1
XFILL_19_1 gnd vdd FILL
XCLKBUF1_2 CLKBUF1_2/A gnd CLKBUF1_2/Y vdd CLKBUF1
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_3/B vdd MUX2X1
XDFFPOSX1_108 MUX2X1_77/A CLKBUF1_43/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_119 MUX2X1_148/A CLKBUF1_5/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XBUFX4_57 INVX8_8/Y gnd BUFX4_57/Y vdd BUFX4
XBUFX4_24 INVX8_6/Y gnd BUFX4_24/Y vdd BUFX4
XDFFPOSX1_90 MUX2X1_31/B CLKBUF1_32/A OAI21X1_24/Y gnd vdd DFFPOSX1
XBUFX4_46 INVX8_4/Y gnd BUFX4_46/Y vdd BUFX4
XBUFX4_13 address[1] gnd BUFX4_13/Y vdd BUFX4
XINVX8_4 datain[3] gnd INVX8_4/Y vdd INVX8
XBUFX4_35 address[0] gnd BUFX4_35/Y vdd BUFX4
XFILL_21_2_0 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XNAND2X1_27 MUX2X1_7/B NAND2X1_27/B gnd OAI21X1_23/C vdd NAND2X1
XOAI21X1_174 BUFX4_55/Y OAI21X1_174/B NAND2X1_196/Y gnd OAI21X1_174/Y vdd OAI21X1
XNAND2X1_191 MUX2X1_50/B OAI21X1_174/B gnd OAI21X1_169/C vdd NAND2X1
XOAI21X1_185 BUFX4_14/Y OAI21X1_183/B OAI21X1_185/C gnd DFFPOSX1_3/D vdd OAI21X1
XNAND2X1_180 MUX2X1_16/B OAI21X1_162/B gnd NAND2X1_180/Y vdd NAND2X1
XNAND2X1_38 MUX2X1_53/A OAI21X1_38/B gnd OAI21X1_33/C vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XNAND2X1_16 NAND2X1_16/A OAI21X1_7/B gnd OAI21X1_14/C vdd NAND2X1
XOAI21X1_130 BUFX4_46/Y OAI21X1_134/B NAND2X1_147/Y gnd OAI21X1_130/Y vdd OAI21X1
XOAI21X1_152 BUFX4_50/Y NAND2X1_173/B OAI21X1_152/C gnd OAI21X1_152/Y vdd OAI21X1
XAOI22X1_6 AOI22X1_6/A AOI22X1_2/B AOI22X1_2/C MUX2X1_36/Y gnd AOI22X1_6/Y vdd AOI22X1
XFILL_9_2_0 gnd vdd FILL
XOAI21X1_196 BUFX4_25/Y OAI21X1_193/B OAI21X1_196/C gnd OAI21X1_196/Y vdd OAI21X1
XOAI21X1_163 BUFX4_1/Y OAI21X1_162/B OAI21X1_163/C gnd OAI21X1_163/Y vdd OAI21X1
XNAND2X1_49 MUX2X1_100/A NAND2X1_50/B gnd NAND2X1_49/Y vdd NAND2X1
XOAI21X1_141 BUFX4_44/Y NAND2X1_160/B NAND2X1_159/Y gnd OAI21X1_141/Y vdd OAI21X1
XAOI22X1_14 MUX2X1_81/Y AOI22X1_2/B AOI22X1_2/C MUX2X1_84/Y gnd AOI22X1_14/Y vdd AOI22X1
XAOI22X1_25 MUX2X1_147/Y NOR2X1_2/Y AOI22X1_9/C AOI22X1_25/D gnd AOI22X1_25/Y vdd
+ AOI22X1
XFILL_19_2 gnd vdd FILL
XMUX2X1_2 NOR2X1_3/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_3/A vdd MUX2X1
XCLKBUF1_3 CLKBUF1_2/A gnd CLKBUF1_3/Y vdd CLKBUF1
XDFFPOSX1_109 NAND2X1_40/A CLKBUF1_35/Y OAI21X1_35/Y gnd vdd DFFPOSX1
XFILL_6_0_0 gnd vdd FILL
XDFFPOSX1_80 NOR2X1_10/A CLKBUF1_33/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_91 MUX2X1_55/B CLKBUF1_23/A OAI21X1_25/Y gnd vdd DFFPOSX1
XBUFX4_14 INVX8_3/Y gnd BUFX4_14/Y vdd BUFX4
XBUFX4_58 INVX8_8/Y gnd BUFX4_58/Y vdd BUFX4
XBUFX4_47 INVX8_4/Y gnd BUFX4_47/Y vdd BUFX4
XBUFX4_25 INVX8_6/Y gnd BUFX4_25/Y vdd BUFX4
XINVX8_5 datain[4] gnd BUFX4_2/A vdd INVX8
XBUFX4_36 address[0] gnd BUFX4_36/Y vdd BUFX4
XFILL_21_2_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XOAI21X1_142 BUFX4_59/Y NAND2X1_160/B OAI21X1_142/C gnd OAI21X1_142/Y vdd OAI21X1
XOAI21X1_175 NAND2X1_198/Y OAI21X1_175/B INVX4_2/Y gnd AOI21X1_25/B vdd OAI21X1
XNAND2X1_28 MUX2X1_31/B NAND2X1_27/B gnd OAI21X1_24/C vdd NAND2X1
XOAI21X1_153 BUFX4_18/Y NAND2X1_173/B OAI21X1_153/C gnd OAI21X1_153/Y vdd OAI21X1
XNAND2X1_181 MUX2X1_40/B OAI21X1_162/B gnd OAI21X1_160/C vdd NAND2X1
XOAI21X1_120 BUFX4_50/Y OAI21X1_126/B NAND2X1_136/Y gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_186 BUFX4_45/Y OAI21X1_183/B OAI21X1_186/C gnd DFFPOSX1_4/D vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AOI22X1_3/B INVX8_9/Y AOI22X1_7/D gnd AOI22X1_7/Y vdd AOI22X1
XNAND2X1_192 MUX2X1_74/B OAI21X1_174/B gnd NAND2X1_192/Y vdd NAND2X1
XNAND2X1_170 AOI22X1_3/B AND2X2_4/B gnd NAND2X1_173/B vdd NAND2X1
XNAND2X1_39 MUX2X1_77/A OAI21X1_38/B gnd NAND2X1_39/Y vdd NAND2X1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_197 BUFX4_40/Y OAI21X1_193/B OAI21X1_197/C gnd OAI21X1_197/Y vdd OAI21X1
XNAND2X1_17 NOR2X1_33/Y NOR2X1_2/Y gnd OAI21X1_18/B vdd NAND2X1
XOAI21X1_131 BUFX4_4/Y OAI21X1_134/B NAND2X1_148/Y gnd OAI21X1_131/Y vdd OAI21X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_164 BUFX4_24/Y OAI21X1_162/B NAND2X1_185/Y gnd OAI21X1_164/Y vdd OAI21X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 MUX2X1_87/Y AOI22X1_3/B INVX8_9/Y MUX2X1_90/Y gnd AOI22X1_15/Y vdd AOI22X1
XAOI22X1_26 MUX2X1_153/Y AOI22X1_2/B AOI22X1_2/C AOI22X1_26/D gnd AOI22X1_26/Y vdd
+ AOI22X1
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B BUFX4_7/Y gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 CLKBUF1_4/A gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XFILL_24_1 gnd vdd FILL
XBUFX4_59 INVX8_8/Y gnd BUFX4_59/Y vdd BUFX4
XBUFX4_15 INVX8_3/Y gnd BUFX4_15/Y vdd BUFX4
XDFFPOSX1_81 MUX2X1_1/B CLKBUF1_29/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_92 MUX2X1_79/B CLKBUF1_38/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XBUFX4_48 INVX8_4/Y gnd BUFX4_48/Y vdd BUFX4
XBUFX4_26 INVX8_6/Y gnd BUFX4_26/Y vdd BUFX4
XDFFPOSX1_70 MUX2X1_128/B CLKBUF1_10/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XINVX8_6 datain[5] gnd INVX8_6/Y vdd INVX8
XBUFX4_37 address[0] gnd BUFX4_37/Y vdd BUFX4
XDFFPOSX1_260 BUFX2_4/A CLKBUF1_19/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XOAI21X1_121 BUFX4_17/Y OAI21X1_126/B OAI21X1_121/C gnd OAI21X1_121/Y vdd OAI21X1
XOAI21X1_110 BUFX4_59/Y OAI21X1_105/B NAND2X1_124/Y gnd OAI21X1_110/Y vdd OAI21X1
XOAI21X1_143 BUFX4_23/Y NAND2X1_169/B OAI21X1_143/C gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_198 BUFX4_57/Y OAI21X1_193/B OAI21X1_198/C gnd DFFPOSX1_16/D vdd OAI21X1
XOAI21X1_176 NAND2X1_201/Y NAND2X1_202/Y INVX4_2/Y gnd AOI21X1_26/B vdd OAI21X1
XAOI22X1_8 MUX2X1_45/Y AOI22X1_4/B AOI22X1_4/C MUX2X1_48/Y gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_154 BUFX4_48/Y NAND2X1_173/B NAND2X1_174/Y gnd OAI21X1_154/Y vdd OAI21X1
XOAI21X1_132 BUFX4_27/Y OAI21X1_134/B NAND2X1_149/Y gnd OAI21X1_132/Y vdd OAI21X1
XOAI21X1_187 BUFX4_3/Y OAI21X1_183/B NAND2X1_229/Y gnd DFFPOSX1_5/D vdd OAI21X1
XOAI21X1_165 BUFX4_42/Y OAI21X1_162/B NAND2X1_186/Y gnd OAI21X1_165/Y vdd OAI21X1
XNAND2X1_29 MUX2X1_55/B NAND2X1_27/B gnd NAND2X1_29/Y vdd NAND2X1
XNAND2X1_160 MUX2X1_181/A NAND2X1_160/B gnd OAI21X1_142/C vdd NAND2X1
XNAND2X1_182 MUX2X1_64/B OAI21X1_162/B gnd NAND2X1_182/Y vdd NAND2X1
XNAND2X1_18 MUX2X1_1/B OAI21X1_18/B gnd OAI21X1_15/C vdd NAND2X1
XNAND2X1_171 MUX2X1_14/A NAND2X1_173/B gnd OAI21X1_151/C vdd NAND2X1
XAOI22X1_16 MUX2X1_93/Y AOI22X1_4/B AOI22X1_4/C MUX2X1_96/Y gnd AOI22X1_16/Y vdd AOI22X1
XAOI22X1_27 MUX2X1_159/Y AOI22X1_3/B INVX8_9/Y AOI22X1_27/D gnd AOI22X1_27/Y vdd AOI22X1
XNAND2X1_193 MUX2X1_98/B OAI21X1_174/B gnd NAND2X1_193/Y vdd NAND2X1
XFILL_10_3_0 gnd vdd FILL
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_4/S gnd MUX2X1_4/Y vdd MUX2X1
XFILL_17_1 gnd vdd FILL
XCLKBUF1_5 CLKBUF1_7/A gnd CLKBUF1_5/Y vdd CLKBUF1
XDFFPOSX1_82 MUX2X1_25/B CLKBUF1_28/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_60 NAND2X1_2/A CLKBUF1_43/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XINVX8_7 datain[6] gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_93 MUX2X1_103/B CLKBUF1_8/A OAI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 MUX2X1_152/B CLKBUF1_6/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XBUFX4_16 INVX8_3/Y gnd BUFX4_16/Y vdd BUFX4
XFILL_15_2_0 gnd vdd FILL
XBUFX4_49 INVX8_4/Y gnd BUFX4_49/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XBUFX4_27 INVX8_6/Y gnd BUFX4_27/Y vdd BUFX4
XBUFX4_38 address[0] gnd INVX1_3/A vdd BUFX4
XFILL_21_0_0 gnd vdd FILL
XDFFPOSX1_250 MUX2X1_41/B CLKBUF1_31/A AOI21X1_18/Y gnd vdd DFFPOSX1
XFILL_12_0_0 gnd vdd FILL
XBUFX4_1 BUFX4_2/A gnd BUFX4_1/Y vdd BUFX4
XINVX4_1 enable gnd INVX4_1/Y vdd INVX4
XDFFPOSX1_261 BUFX2_5/A CLKBUF1_14/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_111 BUFX4_22/Y OAI21X1_118/B OAI21X1_111/C gnd OAI21X1_111/Y vdd OAI21X1
XOAI21X1_177 NAND2X1_204/Y OAI21X1_177/B INVX4_2/Y gnd AOI21X1_27/B vdd OAI21X1
XAOI22X1_9 MUX2X1_51/Y NOR2X1_2/Y AOI22X1_9/C AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_199 BUFX4_19/Y OAI21X1_201/B NAND2X1_244/Y gnd DFFPOSX1_17/D vdd OAI21X1
XOAI21X1_122 BUFX4_46/Y OAI21X1_126/B NAND2X1_138/Y gnd OAI21X1_122/Y vdd OAI21X1
XOAI21X1_144 BUFX4_53/Y NAND2X1_169/B NAND2X1_163/Y gnd OAI21X1_144/Y vdd OAI21X1
XOAI21X1_188 BUFX4_28/Y OAI21X1_183/B NAND2X1_230/Y gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_133 BUFX4_44/Y OAI21X1_134/B OAI21X1_133/C gnd OAI21X1_133/Y vdd OAI21X1
XOAI21X1_155 BUFX4_5/Y NAND2X1_173/B OAI21X1_155/C gnd OAI21X1_155/Y vdd OAI21X1
XOAI21X1_100 BUFX4_28/Y OAI21X1_97/B NAND2X1_113/Y gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_166 BUFX4_55/Y OAI21X1_162/B OAI21X1_166/C gnd OAI21X1_166/Y vdd OAI21X1
XNAND2X1_183 MUX2X1_88/B OAI21X1_162/B gnd OAI21X1_162/C vdd NAND2X1
XNAND2X1_19 MUX2X1_25/B OAI21X1_18/B gnd NAND2X1_19/Y vdd NAND2X1
XNAND2X1_172 MUX2X1_38/A NAND2X1_173/B gnd OAI21X1_152/C vdd NAND2X1
XAOI22X1_28 AOI22X1_28/A AOI22X1_4/B AOI22X1_4/C MUX2X1_168/Y gnd AOI22X1_28/Y vdd
+ AOI22X1
XNAND2X1_161 AOI22X1_3/B NOR2X1_1/Y gnd NAND2X1_169/B vdd NAND2X1
XNAND2X1_150 MUX2X1_157/B OAI21X1_134/B gnd OAI21X1_133/C vdd NAND2X1
XNAND2X1_194 MUX2X1_122/B OAI21X1_174/B gnd OAI21X1_172/C vdd NAND2X1
XAOI22X1_17 MUX2X1_99/Y NOR2X1_2/Y AOI22X1_9/C MUX2X1_102/Y gnd AOI22X1_17/Y vdd AOI22X1
XFILL_5_1 gnd vdd FILL
XOAI21X1_1 BUFX4_15/Y NAND2X1_1/B NAND2X1_1/Y gnd OAI21X1_1/Y vdd OAI21X1
XFILL_10_3_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B MUX2X1_5/S gnd MUX2X1_6/A vdd MUX2X1
XFILL_17_2 gnd vdd FILL
XCLKBUF1_6 CLKBUF1_6/A gnd CLKBUF1_6/Y vdd CLKBUF1
XINVX8_8 datain[7] gnd INVX8_8/Y vdd INVX8
XBUFX4_17 INVX8_3/Y gnd BUFX4_17/Y vdd BUFX4
XDFFPOSX1_72 NAND2X1_16/A CLKBUF1_3/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XFILL_15_2_1 gnd vdd FILL
XDFFPOSX1_83 MUX2X1_49/B CLKBUF1_24/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 MUX2X1_32/A CLKBUF1_28/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XFILL_7_3_1 gnd vdd FILL
XDFFPOSX1_61 NAND2X1_3/A CLKBUF1_6/A OAI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 MUX2X1_127/B CLKBUF1_9/A OAI21X1_28/Y gnd vdd DFFPOSX1
XBUFX4_28 INVX8_6/Y gnd BUFX4_28/Y vdd BUFX4
XBUFX4_39 address[0] gnd BUFX4_39/Y vdd BUFX4
XDFFPOSX1_240 MUX2X1_184/B CLKBUF1_33/Y OAI21X1_166/Y gnd vdd DFFPOSX1
XFILL_21_0_1 gnd vdd FILL
XDFFPOSX1_251 NOR2X1_23/A CLKBUF1_23/A AOI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_262 BUFX2_6/A CLKBUF1_10/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XBUFX4_2 BUFX4_2/A gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 r_w gnd INVX4_2/Y vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XOAI21X1_112 BUFX4_53/Y OAI21X1_118/B NAND2X1_127/Y gnd OAI21X1_112/Y vdd OAI21X1
XOAI21X1_101 BUFX4_43/Y OAI21X1_97/B NAND2X1_114/Y gnd OAI21X1_101/Y vdd OAI21X1
XOAI21X1_134 BUFX4_55/Y OAI21X1_134/B NAND2X1_151/Y gnd OAI21X1_134/Y vdd OAI21X1
XAOI22X1_29 AOI22X1_29/A NOR2X1_2/Y AOI22X1_9/C AOI22X1_29/D gnd AOI22X1_29/Y vdd
+ AOI22X1
XOAI21X1_167 BUFX4_23/Y OAI21X1_174/B NAND2X1_189/Y gnd OAI21X1_167/Y vdd OAI21X1
XOAI21X1_145 BUFX4_18/Y NAND2X1_169/B NAND2X1_164/Y gnd OAI21X1_145/Y vdd OAI21X1
XNAND2X1_173 MUX2X1_62/A NAND2X1_173/B gnd OAI21X1_153/C vdd NAND2X1
XNAND2X1_162 MUX2X1_14/B NAND2X1_169/B gnd OAI21X1_143/C vdd NAND2X1
XOAI21X1_178 NAND2X1_207/Y OAI21X1_178/B INVX4_2/Y gnd AOI21X1_28/B vdd OAI21X1
XNAND2X1_184 MUX2X1_112/B OAI21X1_162/B gnd OAI21X1_163/C vdd NAND2X1
XOAI21X1_156 BUFX4_27/Y NAND2X1_173/B OAI21X1_156/C gnd OAI21X1_156/Y vdd OAI21X1
XOAI21X1_189 BUFX4_41/Y OAI21X1_183/B OAI21X1_189/C gnd DFFPOSX1_7/D vdd OAI21X1
XNAND2X1_140 MUX2X1_143/A OAI21X1_126/B gnd OAI21X1_124/C vdd NAND2X1
XNAND2X1_195 MUX2X1_146/B OAI21X1_174/B gnd NAND2X1_195/Y vdd NAND2X1
XOAI21X1_123 BUFX4_4/Y OAI21X1_126/B OAI21X1_123/C gnd OAI21X1_123/Y vdd OAI21X1
XNAND2X1_151 MUX2X1_181/B OAI21X1_134/B gnd NAND2X1_151/Y vdd NAND2X1
XAOI22X1_18 MUX2X1_105/Y AOI22X1_2/B AOI22X1_2/C MUX2X1_108/Y gnd AOI22X1_18/Y vdd
+ AOI22X1
XMUX2X1_190 MUX2X1_190/A MUX2X1_190/B MUX2X1_8/S gnd MUX2X1_192/B vdd MUX2X1
XFILL_5_2 gnd vdd FILL
XAOI21X1_40 BUFX4_56/Y AND2X2_4/Y NOR2X1_42/Y gnd AOI21X1_40/Y vdd AOI21X1
XOAI21X1_2 BUFX4_47/Y NAND2X1_1/B NAND2X1_2/Y gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XMUX2X1_6 MUX2X1_6/A MUX2X1_4/Y BUFX4_8/Y gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 CLKBUF1_7/A gnd CLKBUF1_7/Y vdd CLKBUF1
XFILL_17_3 gnd vdd FILL
XDFFPOSX1_84 MUX2X1_73/B CLKBUF1_20/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 MUX2X1_188/A CLKBUF1_1/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_73 NOR2X1_3/A CLKBUF1_32/A AOI21X1_1/Y gnd vdd DFFPOSX1
XBUFX4_18 INVX8_3/Y gnd BUFX4_18/Y vdd BUFX4
XDFFPOSX1_51 MUX2X1_56/A CLKBUF1_24/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XINVX8_9 OR2X2_1/Y gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_62 NAND2X1_4/A CLKBUF1_43/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_95 NAND2X1_33/A CLKBUF1_6/A OAI21X1_29/Y gnd vdd DFFPOSX1
XBUFX4_29 address[0] gnd MUX2X1_1/S vdd BUFX4
XFILL_22_1 gnd vdd FILL
XDFFPOSX1_241 MUX2X1_2/B CLKBUF1_31/Y OAI21X1_167/Y gnd vdd DFFPOSX1
XDFFPOSX1_230 MUX2X1_134/A CLKBUF1_12/Y OAI21X1_156/Y gnd vdd DFFPOSX1
XBUFX4_3 BUFX4_2/A gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_263 BUFX2_7/A CLKBUF1_6/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_252 NOR2X1_24/A CLKBUF1_9/A AOI21X1_20/Y gnd vdd DFFPOSX1
XFILL_22_3_0 gnd vdd FILL
XNAND2X1_196 MUX2X1_170/B OAI21X1_174/B gnd NAND2X1_196/Y vdd NAND2X1
XOAI21X1_113 BUFX4_17/Y OAI21X1_118/B OAI21X1_113/C gnd OAI21X1_113/Y vdd OAI21X1
XOAI21X1_102 BUFX4_56/Y OAI21X1_97/B NAND2X1_115/Y gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_135 BUFX4_23/Y NAND2X1_160/B OAI21X1_135/C gnd OAI21X1_135/Y vdd OAI21X1
XFILL_13_3_0 gnd vdd FILL
XOAI21X1_168 BUFX4_52/Y OAI21X1_174/B OAI21X1_168/C gnd OAI21X1_168/Y vdd OAI21X1
XOAI21X1_146 BUFX4_48/Y NAND2X1_169/B OAI21X1_146/C gnd OAI21X1_146/Y vdd OAI21X1
XNAND2X1_174 MUX2X1_86/A NAND2X1_173/B gnd NAND2X1_174/Y vdd NAND2X1
XNAND2X1_163 MUX2X1_38/B NAND2X1_169/B gnd NAND2X1_163/Y vdd NAND2X1
XNAND2X1_152 AOI22X1_3/B AND2X2_2/B gnd NAND2X1_160/B vdd NAND2X1
XNAND2X1_141 MUX2X1_167/A OAI21X1_126/B gnd NAND2X1_141/Y vdd NAND2X1
XOAI21X1_157 BUFX4_44/Y NAND2X1_173/B OAI21X1_157/C gnd OAI21X1_157/Y vdd OAI21X1
XOAI21X1_124 BUFX4_27/Y OAI21X1_126/B OAI21X1_124/C gnd OAI21X1_124/Y vdd OAI21X1
XNAND2X1_130 MUX2X1_119/B OAI21X1_118/B gnd OAI21X1_115/C vdd NAND2X1
XNAND2X1_185 MUX2X1_136/B OAI21X1_162/B gnd NAND2X1_185/Y vdd NAND2X1
XOAI21X1_179 NAND2X1_210/Y OAI21X1_179/B INVX4_2/Y gnd AOI21X1_29/B vdd OAI21X1
XMUX2X1_191 MUX2X1_191/A MUX2X1_191/B BUFX4_35/Y gnd MUX2X1_192/A vdd MUX2X1
XMUX2X1_180 MUX2X1_180/A MUX2X1_178/Y BUFX4_10/Y gnd MUX2X1_180/Y vdd MUX2X1
XAOI22X1_19 MUX2X1_111/Y AOI22X1_3/B INVX8_9/Y MUX2X1_114/Y gnd AOI22X1_19/Y vdd AOI22X1
XAOI21X1_30 AOI21X1_30/A AOI21X1_30/B INVX4_1/Y gnd AOI21X1_30/Y vdd AOI21X1
XOAI21X1_3 BUFX4_5/Y NAND2X1_1/B NAND2X1_3/Y gnd OAI21X1_3/Y vdd OAI21X1
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_7/S gnd MUX2X1_9/B vdd MUX2X1
XFILL_10_1_0 gnd vdd FILL
XCLKBUF1_8 CLKBUF1_8/A gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_2_2_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_41 NOR2X1_35/A CLKBUF1_32/A AOI21X1_33/Y gnd vdd DFFPOSX1
XBUFX4_19 INVX8_1/Y gnd BUFX4_19/Y vdd BUFX4
XDFFPOSX1_96 MUX2X1_175/B CLKBUF1_43/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 NOR2X1_4/A CLKBUF1_31/A AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 MUX2X1_80/A CLKBUF1_17/Y OAI21X1_226/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 MUX2X1_130/B CLKBUF1_7/A DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_63 NAND2X1_5/A CLKBUF1_7/A OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 MUX2X1_97/B CLKBUF1_14/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XFILL_22_2 gnd vdd FILL
XFILL_15_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XDFFPOSX1_264 BUFX2_8/A CLKBUF1_1/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_242 MUX2X1_26/B CLKBUF1_28/Y OAI21X1_168/Y gnd vdd DFFPOSX1
XDFFPOSX1_220 MUX2X1_86/B CLKBUF1_43/Y OAI21X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_231 MUX2X1_158/A CLKBUF1_7/Y OAI21X1_157/Y gnd vdd DFFPOSX1
XBUFX4_4 BUFX4_2/A gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_253 NOR2X1_25/A CLKBUF1_6/A AOI21X1_21/Y gnd vdd DFFPOSX1
XOAI21X1_103 BUFX4_20/Y OAI21X1_105/B NAND2X1_117/Y gnd OAI21X1_103/Y vdd OAI21X1
XFILL_22_3_1 gnd vdd FILL
XNAND2X1_142 MUX2X1_191/A OAI21X1_126/B gnd NAND2X1_142/Y vdd NAND2X1
XOAI21X1_169 BUFX4_17/Y OAI21X1_174/B OAI21X1_169/C gnd OAI21X1_169/Y vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd dataout[0] vdd BUFX2
XNAND2X1_197 r_w BUFX2_1/A gnd AOI21X1_25/A vdd NAND2X1
XOAI21X1_158 BUFX4_58/Y NAND2X1_173/B OAI21X1_158/C gnd OAI21X1_158/Y vdd OAI21X1
XNAND2X1_164 MUX2X1_62/B NAND2X1_169/B gnd NAND2X1_164/Y vdd NAND2X1
XNAND2X1_153 MUX2X1_13/A NAND2X1_160/B gnd OAI21X1_135/C vdd NAND2X1
XNAND2X1_120 MUX2X1_94/A OAI21X1_105/B gnd NAND2X1_120/Y vdd NAND2X1
XOAI21X1_114 BUFX4_46/Y OAI21X1_118/B NAND2X1_129/Y gnd OAI21X1_114/Y vdd OAI21X1
XOAI21X1_136 BUFX4_53/Y NAND2X1_160/B OAI21X1_136/C gnd OAI21X1_136/Y vdd OAI21X1
XOAI21X1_125 BUFX4_44/Y OAI21X1_126/B NAND2X1_141/Y gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_147 BUFX4_5/Y NAND2X1_169/B NAND2X1_166/Y gnd OAI21X1_147/Y vdd OAI21X1
XNAND2X1_131 MUX2X1_143/B OAI21X1_118/B gnd OAI21X1_116/C vdd NAND2X1
XNAND2X1_175 MUX2X1_110/A NAND2X1_173/B gnd OAI21X1_155/C vdd NAND2X1
XNAND2X1_186 MUX2X1_160/B OAI21X1_162/B gnd NAND2X1_186/Y vdd NAND2X1
XAOI21X1_1 BUFX4_20/Y NOR2X1_5/B NOR2X1_3/Y gnd AOI21X1_1/Y vdd AOI21X1
XMUX2X1_170 NOR2X1_10/A MUX2X1_170/B MUX2X1_5/S gnd MUX2X1_171/A vdd MUX2X1
XMUX2X1_192 MUX2X1_192/A MUX2X1_192/B BUFX4_6/Y gnd AOI22X1_32/D vdd MUX2X1
XMUX2X1_181 MUX2X1_181/A MUX2X1_181/B BUFX4_39/Y gnd MUX2X1_183/B vdd MUX2X1
XINVX2_1 address[2] gnd OR2X2_1/B vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XOAI21X1_4 BUFX4_26/Y NAND2X1_1/B OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_31 AOI21X1_31/A AOI21X1_31/B INVX4_1/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_20 BUFX4_47/Y AND2X2_3/Y NOR2X1_24/Y gnd AOI21X1_20/Y vdd AOI21X1
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B MUX2X1_8/S gnd MUX2X1_9/A vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XCLKBUF1_9 CLKBUF1_9/A gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_18_2_1 gnd vdd FILL
XDFFPOSX1_75 NOR2X1_5/A CLKBUF1_2/A AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_97 MUX2X1_16/A CLKBUF1_30/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 NAND2X1_6/A CLKBUF1_4/A OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 MUX2X1_41/A CLKBUF1_31/A AOI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 MUX2X1_83/A CLKBUF1_18/Y DFFPOSX1_20/D gnd vdd DFFPOSX1
XDFFPOSX1_31 MUX2X1_154/B CLKBUF1_31/A DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_53 MUX2X1_104/A CLKBUF1_15/Y OAI21X1_227/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 MUX2X1_121/B CLKBUF1_11/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XFILL_15_2 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XDFFPOSX1_243 MUX2X1_50/B CLKBUF1_23/Y OAI21X1_169/Y gnd vdd DFFPOSX1
XDFFPOSX1_232 MUX2X1_182/A CLKBUF1_3/Y OAI21X1_158/Y gnd vdd DFFPOSX1
XDFFPOSX1_210 MUX2X1_37/A CLKBUF1_25/Y OAI21X1_136/Y gnd vdd DFFPOSX1
XDFFPOSX1_254 NOR2X1_26/A CLKBUF1_43/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_221 MUX2X1_110/B CLKBUF1_6/A OAI21X1_147/Y gnd vdd DFFPOSX1
XBUFX4_5 BUFX4_2/A gnd BUFX4_5/Y vdd BUFX4
XNAND2X1_110 MUX2X1_70/B OAI21X1_97/B gnd OAI21X1_97/C vdd NAND2X1
XOAI21X1_126 BUFX4_59/Y OAI21X1_126/B NAND2X1_142/Y gnd OAI21X1_126/Y vdd OAI21X1
XOAI21X1_137 BUFX4_15/Y NAND2X1_160/B OAI21X1_137/C gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_159 BUFX4_19/Y OAI21X1_162/B NAND2X1_180/Y gnd OAI21X1_159/Y vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd dataout[1] vdd BUFX2
XNAND2X1_143 AOI22X1_3/B NOR2X1_33/Y gnd OAI21X1_134/B vdd NAND2X1
XOAI21X1_104 BUFX4_51/Y OAI21X1_105/B OAI21X1_104/C gnd OAI21X1_104/Y vdd OAI21X1
XOAI21X1_148 BUFX4_27/Y NAND2X1_169/B OAI21X1_148/C gnd OAI21X1_148/Y vdd OAI21X1
XNAND2X1_132 MUX2X1_167/B OAI21X1_118/B gnd OAI21X1_117/C vdd NAND2X1
XNAND2X1_121 MUX2X1_118/A OAI21X1_105/B gnd NAND2X1_121/Y vdd NAND2X1
XOAI21X1_115 BUFX4_4/Y OAI21X1_118/B OAI21X1_115/C gnd OAI21X1_115/Y vdd OAI21X1
XNAND2X1_187 MUX2X1_184/B OAI21X1_162/B gnd OAI21X1_166/C vdd NAND2X1
XMUX2X1_171 MUX2X1_171/A MUX2X1_171/B BUFX4_7/Y gnd AOI22X1_29/A vdd MUX2X1
XNAND2X1_198 AOI22X1_1/Y AOI22X1_2/Y gnd NAND2X1_198/Y vdd NAND2X1
XMUX2X1_182 MUX2X1_182/A MUX2X1_182/B MUX2X1_1/S gnd MUX2X1_182/Y vdd MUX2X1
XNAND2X1_165 MUX2X1_86/B NAND2X1_169/B gnd OAI21X1_146/C vdd NAND2X1
XAOI21X1_2 BUFX4_51/Y NOR2X1_5/B NOR2X1_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XNAND2X1_154 MUX2X1_37/A NAND2X1_160/B gnd OAI21X1_136/C vdd NAND2X1
XNAND2X1_176 MUX2X1_134/A NAND2X1_173/B gnd OAI21X1_156/C vdd NAND2X1
XMUX2X1_160 NOR2X1_17/A MUX2X1_160/B BUFX4_36/Y gnd MUX2X1_160/Y vdd MUX2X1
XAOI21X1_32 AOI21X1_32/A AOI21X1_32/B INVX4_1/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_10 BUFX4_50/Y AND2X2_2/Y NOR2X1_12/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_21 BUFX4_1/Y AND2X2_3/Y NOR2X1_25/Y gnd AOI21X1_21/Y vdd AOI21X1
XOAI21X1_5 BUFX4_43/Y NAND2X1_1/B OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B BUFX4_9/Y gnd MUX2X1_9/Y vdd MUX2X1
XDFFPOSX1_43 MUX2X1_65/A CLKBUF1_23/A AOI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_65 MUX2X1_8/B CLKBUF1_31/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 MUX2X1_178/B CLKBUF1_2/A OAI21X1_214/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 MUX2X1_40/A CLKBUF1_27/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 NOR2X1_6/A CLKBUF1_4/A AOI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 MUX2X1_34/A CLKBUF1_40/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XDFFPOSX1_54 MUX2X1_128/A CLKBUF1_9/Y OAI21X1_228/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 MUX2X1_107/A CLKBUF1_16/Y OAI21X1_203/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 MUX2X1_145/B CLKBUF1_8/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XFILL_20_1 gnd vdd FILL
XDFFPOSX1_200 MUX2X1_191/A CLKBUF1_1/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_211 MUX2X1_61/A CLKBUF1_21/Y OAI21X1_137/Y gnd vdd DFFPOSX1
XDFFPOSX1_233 MUX2X1_16/B CLKBUF1_32/A OAI21X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_244 MUX2X1_74/B CLKBUF1_19/Y OAI21X1_170/Y gnd vdd DFFPOSX1
XDFFPOSX1_222 MUX2X1_134/B CLKBUF1_9/A OAI21X1_148/Y gnd vdd DFFPOSX1
XFILL_0_3_0 gnd vdd FILL
XBUFX4_6 address[1] gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_255 NOR2X1_27/A CLKBUF1_7/A AOI21X1_23/Y gnd vdd DFFPOSX1
XFILL_16_3_0 gnd vdd FILL
XOAI21X1_105 BUFX4_16/Y OAI21X1_105/B NAND2X1_119/Y gnd OAI21X1_105/Y vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd dataout[2] vdd BUFX2
XOAI21X1_127 BUFX4_22/Y OAI21X1_134/B NAND2X1_144/Y gnd OAI21X1_127/Y vdd OAI21X1
XOAI21X1_138 BUFX4_46/Y NAND2X1_160/B NAND2X1_156/Y gnd OAI21X1_138/Y vdd OAI21X1
XOAI21X1_116 BUFX4_27/Y OAI21X1_118/B OAI21X1_116/C gnd OAI21X1_116/Y vdd OAI21X1
XOAI21X1_149 BUFX4_43/Y NAND2X1_169/B OAI21X1_149/C gnd OAI21X1_149/Y vdd OAI21X1
XNAND2X1_133 MUX2X1_191/B OAI21X1_118/B gnd NAND2X1_133/Y vdd NAND2X1
XAOI21X1_3 BUFX4_17/Y NOR2X1_5/B NOR2X1_5/Y gnd AOI21X1_3/Y vdd AOI21X1
XNAND2X1_199 AOI22X1_3/Y AOI22X1_4/Y gnd OAI21X1_175/B vdd NAND2X1
XNAND2X1_155 MUX2X1_61/A NAND2X1_160/B gnd OAI21X1_137/C vdd NAND2X1
XMUX2X1_172 NAND2X1_52/A NAND2X1_6/A MUX2X1_7/S gnd MUX2X1_172/Y vdd MUX2X1
XMUX2X1_183 MUX2X1_182/Y MUX2X1_183/B BUFX4_11/Y gnd AOI22X1_31/A vdd MUX2X1
XNAND2X1_144 MUX2X1_13/B OAI21X1_134/B gnd NAND2X1_144/Y vdd NAND2X1
XNAND2X1_111 MUX2X1_94/B OAI21X1_97/B gnd OAI21X1_98/C vdd NAND2X1
XNAND2X1_100 MUX2X1_25/A OAI21X1_90/B gnd OAI21X1_88/C vdd NAND2X1
XNAND2X1_188 NOR2X1_1/Y NOR2X1_2/Y gnd OAI21X1_174/B vdd NAND2X1
XNAND2X1_177 MUX2X1_158/A NAND2X1_173/B gnd OAI21X1_157/C vdd NAND2X1
XNAND2X1_166 MUX2X1_110/B NAND2X1_169/B gnd NAND2X1_166/Y vdd NAND2X1
XNAND2X1_122 MUX2X1_142/A OAI21X1_105/B gnd NAND2X1_122/Y vdd NAND2X1
XMUX2X1_150 MUX2X1_149/Y MUX2X1_148/Y BUFX4_8/Y gnd AOI22X1_25/D vdd MUX2X1
XMUX2X1_161 NOR2X1_41/A NOR2X1_27/A BUFX4_37/Y gnd MUX2X1_162/A vdd MUX2X1
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XAOI21X1_33 BUFX4_21/Y AND2X2_4/Y NOR2X1_35/Y gnd AOI21X1_33/Y vdd AOI21X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_11 BUFX4_17/Y AND2X2_2/Y NOR2X1_13/Y gnd AOI21X1_11/Y vdd AOI21X1
XOAI21X1_6 BUFX4_58/Y NAND2X1_1/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_22 BUFX4_25/Y AND2X2_3/Y NOR2X1_26/Y gnd AOI21X1_22/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 MUX2X1_58/A CLKBUF1_32/A DFFPOSX1_11/D gnd vdd DFFPOSX1
XDFFPOSX1_33 MUX2X1_20/A CLKBUF1_32/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_99 MUX2X1_64/A CLKBUF1_21/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 NAND2X1_25/A CLKBUF1_4/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 MUX2X1_32/B CLKBUF1_25/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 MUX2X1_131/A CLKBUF1_10/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XDFFPOSX1_77 NOR2X1_7/A CLKBUF1_8/A AOI21X1_5/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_44 MUX2X1_89/A CLKBUF1_9/A AOI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 MUX2X1_152/A CLKBUF1_5/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_256 NOR2X1_28/A CLKBUF1_23/A AOI21X1_24/Y gnd vdd DFFPOSX1
XFILL_20_2 gnd vdd FILL
XDFFPOSX1_201 MUX2X1_13/B CLKBUF1_23/A OAI21X1_127/Y gnd vdd DFFPOSX1
XDFFPOSX1_234 MUX2X1_40/B CLKBUF1_38/Y OAI21X1_160/Y gnd vdd DFFPOSX1
XFILL_13_1 gnd vdd FILL
XDFFPOSX1_212 MUX2X1_85/A CLKBUF1_17/Y OAI21X1_138/Y gnd vdd DFFPOSX1
XBUFX4_7 address[1] gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_245 MUX2X1_98/B CLKBUF1_14/Y OAI21X1_171/Y gnd vdd DFFPOSX1
XDFFPOSX1_223 MUX2X1_158/B CLKBUF1_7/A OAI21X1_149/Y gnd vdd DFFPOSX1
XFILL_16_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XOAI21X1_106 BUFX4_45/Y OAI21X1_105/B NAND2X1_120/Y gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_128 BUFX4_50/Y OAI21X1_134/B NAND2X1_145/Y gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_117 BUFX4_44/Y OAI21X1_118/B OAI21X1_117/C gnd OAI21X1_117/Y vdd OAI21X1
XNAND2X1_189 MUX2X1_2/B OAI21X1_174/B gnd NAND2X1_189/Y vdd NAND2X1
XNAND2X1_178 MUX2X1_182/A NAND2X1_173/B gnd OAI21X1_158/C vdd NAND2X1
XNAND2X1_101 MUX2X1_49/A OAI21X1_90/B gnd OAI21X1_89/C vdd NAND2X1
XNAND2X1_145 MUX2X1_37/B OAI21X1_134/B gnd NAND2X1_145/Y vdd NAND2X1
XAOI21X1_4 BUFX4_46/Y NOR2X1_5/B NOR2X1_6/Y gnd AOI21X1_4/Y vdd AOI21X1
XNAND2X1_156 MUX2X1_85/A NAND2X1_160/B gnd NAND2X1_156/Y vdd NAND2X1
XBUFX2_4 BUFX2_4/A gnd dataout[3] vdd BUFX2
XNAND2X1_134 AND2X2_4/B AOI22X1_4/C gnd OAI21X1_126/B vdd NAND2X1
XNAND2X1_167 MUX2X1_134/B NAND2X1_169/B gnd OAI21X1_148/C vdd NAND2X1
XNAND2X1_112 MUX2X1_118/B OAI21X1_97/B gnd OAI21X1_99/C vdd NAND2X1
XNAND2X1_123 MUX2X1_166/A OAI21X1_105/B gnd NAND2X1_123/Y vdd NAND2X1
XOAI21X1_139 BUFX4_5/Y NAND2X1_160/B NAND2X1_157/Y gnd OAI21X1_139/Y vdd OAI21X1
XMUX2X1_173 NAND2X1_43/A MUX2X1_173/B MUX2X1_8/S gnd MUX2X1_174/A vdd MUX2X1
XMUX2X1_184 NOR2X1_18/A MUX2X1_184/B MUX2X1_2/S gnd MUX2X1_186/B vdd MUX2X1
XNOR2X1_2 address[2] NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XMUX2X1_140 MUX2X1_140/A MUX2X1_140/B MUX2X1_8/S gnd MUX2X1_141/A vdd MUX2X1
XMUX2X1_151 MUX2X1_151/A NAND2X1_33/A MUX2X1_2/S gnd MUX2X1_151/Y vdd MUX2X1
XMUX2X1_162 MUX2X1_162/A MUX2X1_160/Y BUFX4_12/Y gnd AOI22X1_27/D vdd MUX2X1
XFILL_22_1_1 gnd vdd FILL
XOAI21X1_7 BUFX4_22/Y OAI21X1_7/B NAND2X1_9/Y gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_34 BUFX4_50/Y AND2X2_4/Y NOR2X1_36/Y gnd AOI21X1_34/Y vdd AOI21X1
XAOI21X1_12 BUFX4_49/Y AND2X2_2/Y NOR2X1_14/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_23 BUFX4_42/Y AND2X2_3/Y NOR2X1_27/Y gnd AOI21X1_23/Y vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_89 MUX2X1_7/B CLKBUF1_32/A OAI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 MUX2X1_56/B CLKBUF1_24/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 MUX2X1_176/A CLKBUF1_3/Y OAI21X1_230/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 MUX2X1_82/A CLKBUF1_18/A DFFPOSX1_12/D gnd vdd DFFPOSX1
XDFFPOSX1_34 MUX2X1_44/A CLKBUF1_25/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XDFFPOSX1_23 MUX2X1_155/A CLKBUF1_5/Y DFFPOSX1_23/D gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_78 NOR2X1_8/A CLKBUF1_9/A AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_45 NOR2X1_39/A CLKBUF1_6/A AOI21X1_37/Y gnd vdd DFFPOSX1
XFILL_18_0_1 gnd vdd FILL
XDFFPOSX1_257 BUFX2_1/A CLKBUF1_30/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XFILL_20_3 gnd vdd FILL
XDFFPOSX1_235 MUX2X1_64/B CLKBUF1_2/A OAI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_224 MUX2X1_182/B CLKBUF1_2/A OAI21X1_150/Y gnd vdd DFFPOSX1
XDFFPOSX1_202 MUX2X1_37/B CLKBUF1_38/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XFILL_13_2 gnd vdd FILL
XBUFX4_8 address[1] gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_213 MUX2X1_109/A CLKBUF1_13/Y OAI21X1_139/Y gnd vdd DFFPOSX1
XDFFPOSX1_246 MUX2X1_122/B CLKBUF1_11/Y OAI21X1_172/Y gnd vdd DFFPOSX1
XNAND2X1_102 MUX2X1_73/A OAI21X1_90/B gnd OAI21X1_90/C vdd NAND2X1
XOAI21X1_118 BUFX4_55/Y OAI21X1_118/B NAND2X1_133/Y gnd OAI21X1_118/Y vdd OAI21X1
XNAND2X1_135 MUX2X1_23/A OAI21X1_126/B gnd OAI21X1_119/C vdd NAND2X1
XNAND2X1_124 MUX2X1_190/A OAI21X1_105/B gnd NAND2X1_124/Y vdd NAND2X1
XOAI21X1_129 BUFX4_15/Y OAI21X1_134/B NAND2X1_146/Y gnd OAI21X1_129/Y vdd OAI21X1
XNAND2X1_146 MUX2X1_61/B OAI21X1_134/B gnd NAND2X1_146/Y vdd NAND2X1
XNAND2X1_179 NOR2X1_33/Y INVX8_9/Y gnd OAI21X1_162/B vdd NAND2X1
XOAI21X1_107 BUFX4_4/Y OAI21X1_105/B NAND2X1_121/Y gnd OAI21X1_107/Y vdd OAI21X1
XNAND2X1_157 MUX2X1_109/A NAND2X1_160/B gnd NAND2X1_157/Y vdd NAND2X1
XNAND2X1_168 MUX2X1_158/B NAND2X1_169/B gnd OAI21X1_149/C vdd NAND2X1
XNAND2X1_113 MUX2X1_142/B OAI21X1_97/B gnd NAND2X1_113/Y vdd NAND2X1
XBUFX2_5 BUFX2_5/A gnd dataout[4] vdd BUFX2
XMUX2X1_185 NOR2X1_42/A NOR2X1_28/A MUX2X1_4/S gnd MUX2X1_186/A vdd MUX2X1
XMUX2X1_174 MUX2X1_174/A MUX2X1_172/Y BUFX4_8/Y gnd AOI22X1_29/D vdd MUX2X1
XMUX2X1_163 MUX2X1_163/A MUX2X1_163/B INVX1_3/A gnd MUX2X1_165/B vdd MUX2X1
XMUX2X1_141 MUX2X1_141/A MUX2X1_139/Y BUFX4_13/Y gnd AOI22X1_24/A vdd MUX2X1
XMUX2X1_130 MUX2X1_130/A MUX2X1_130/B INVX1_3/A gnd MUX2X1_130/Y vdd MUX2X1
XAOI21X1_5 BUFX4_3/Y NOR2X1_5/B NOR2X1_7/Y gnd AOI21X1_5/Y vdd AOI21X1
XMUX2X1_152 MUX2X1_152/A MUX2X1_152/B MUX2X1_4/S gnd MUX2X1_153/A vdd MUX2X1
XAOI21X1_24 BUFX4_56/Y AND2X2_3/Y NOR2X1_28/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_35 BUFX4_16/Y AND2X2_4/Y NOR2X1_37/Y gnd AOI21X1_35/Y vdd AOI21X1
XNOR2X1_3 NOR2X1_3/A NOR2X1_5/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_13 BUFX4_2/Y AND2X2_2/Y NOR2X1_15/Y gnd AOI21X1_13/Y vdd AOI21X1
XOAI21X1_8 BUFX4_51/Y OAI21X1_7/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XDFFPOSX1_35 MUX2X1_68/A CLKBUF1_23/Y DFFPOSX1_35/D gnd vdd DFFPOSX1
XDFFPOSX1_57 MUX2X1_4/B CLKBUF1_23/A DFFPOSX1_57/D gnd vdd DFFPOSX1
XDFFPOSX1_24 MUX2X1_179/A CLKBUF1_4/Y OAI21X1_206/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 MUX2X1_80/B CLKBUF1_18/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_46 NOR2X1_40/A CLKBUF1_43/Y AOI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 MUX2X1_106/A CLKBUF1_6/A DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_79 NOR2X1_9/A CLKBUF1_8/A AOI21X1_7/Y gnd vdd DFFPOSX1
XFILL_20_2_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_203 MUX2X1_61/B CLKBUF1_2/A OAI21X1_129/Y gnd vdd DFFPOSX1
XDFFPOSX1_225 MUX2X1_14/A CLKBUF1_29/Y OAI21X1_151/Y gnd vdd DFFPOSX1
XDFFPOSX1_258 BUFX2_2/A CLKBUF1_27/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XBUFX4_9 address[1] gnd BUFX4_9/Y vdd BUFX4
XDFFPOSX1_247 MUX2X1_146/B CLKBUF1_8/Y OAI21X1_173/Y gnd vdd DFFPOSX1
XDFFPOSX1_214 MUX2X1_133/A CLKBUF1_12/Y OAI21X1_140/Y gnd vdd DFFPOSX1
XDFFPOSX1_236 MUX2X1_88/B CLKBUF1_9/A OAI21X1_162/Y gnd vdd DFFPOSX1
XOAI21X1_119 BUFX4_20/Y OAI21X1_126/B OAI21X1_119/C gnd OAI21X1_119/Y vdd OAI21X1
XNAND2X1_1 MUX2X1_52/B NAND2X1_1/B gnd NAND2X1_1/Y vdd NAND2X1
XNAND2X1_169 MUX2X1_182/B NAND2X1_169/B gnd OAI21X1_150/C vdd NAND2X1
XNAND2X1_136 MUX2X1_47/A OAI21X1_126/B gnd NAND2X1_136/Y vdd NAND2X1
XNAND2X1_147 MUX2X1_85/B OAI21X1_134/B gnd NAND2X1_147/Y vdd NAND2X1
XNAND2X1_125 NOR2X1_1/Y AOI22X1_4/C gnd OAI21X1_118/B vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd dataout[5] vdd BUFX2
XNAND2X1_114 MUX2X1_166/B OAI21X1_97/B gnd NAND2X1_114/Y vdd NAND2X1
XNAND2X1_158 MUX2X1_133/A NAND2X1_160/B gnd NAND2X1_158/Y vdd NAND2X1
XNAND2X1_103 MUX2X1_97/A OAI21X1_90/B gnd OAI21X1_91/C vdd NAND2X1
XOAI21X1_108 BUFX4_28/Y OAI21X1_105/B NAND2X1_122/Y gnd OAI21X1_108/Y vdd OAI21X1
XDFFPOSX1_1 MUX2X1_7/A CLKBUF1_32/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XMUX2X1_186 MUX2X1_186/A MUX2X1_186/B BUFX4_12/Y gnd AOI22X1_31/D vdd MUX2X1
XMUX2X1_175 DFFPOSX1_8/Q MUX2X1_175/B BUFX4_35/Y gnd MUX2X1_175/Y vdd MUX2X1
XFILL_16_1_0 gnd vdd FILL
XMUX2X1_131 MUX2X1_131/A MUX2X1_131/B BUFX4_39/Y gnd MUX2X1_132/A vdd MUX2X1
XFILL_8_2_0 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XMUX2X1_120 MUX2X1_120/A MUX2X1_118/Y BUFX4_6/Y gnd MUX2X1_120/Y vdd MUX2X1
XMUX2X1_142 MUX2X1_142/A MUX2X1_142/B BUFX4_35/Y gnd MUX2X1_142/Y vdd MUX2X1
XAOI21X1_6 BUFX4_24/Y NOR2X1_5/B NOR2X1_8/Y gnd AOI21X1_6/Y vdd AOI21X1
XMUX2X1_164 MUX2X1_164/A MUX2X1_164/B BUFX4_39/Y gnd MUX2X1_164/Y vdd MUX2X1
XMUX2X1_153 MUX2X1_153/A MUX2X1_151/Y BUFX4_9/Y gnd MUX2X1_153/Y vdd MUX2X1
XNOR2X1_4 NOR2X1_4/A NOR2X1_5/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_25 AOI21X1_25/A AOI21X1_25/B INVX4_1/Y gnd AOI21X1_25/Y vdd AOI21X1
XOAI21X1_9 BUFX4_18/Y OAI21X1_7/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_36 BUFX4_47/Y AND2X2_4/Y NOR2X1_38/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_14 BUFX4_24/Y AND2X2_2/Y NOR2X1_16/Y gnd AOI21X1_14/Y vdd AOI21X1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_25 MUX2X1_10/B CLKBUF1_31/A DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_36 MUX2X1_92/A CLKBUF1_17/Y OAI21X1_218/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 MUX2X1_28/B CLKBUF1_6/A OAI21X1_232/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 MUX2X1_130/A CLKBUF1_7/A OAI21X1_196/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 NOR2X1_41/A CLKBUF1_7/A AOI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 MUX2X1_104/B CLKBUF1_14/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XFILL_20_2_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XDFFPOSX1_248 MUX2X1_170/B CLKBUF1_1/Y OAI21X1_174/Y gnd vdd DFFPOSX1
XDFFPOSX1_259 BUFX2_3/A CLKBUF1_23/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_204 MUX2X1_85/B CLKBUF1_43/Y OAI21X1_130/Y gnd vdd DFFPOSX1
XDFFPOSX1_226 MUX2X1_38/A CLKBUF1_27/Y OAI21X1_152/Y gnd vdd DFFPOSX1
XDFFPOSX1_237 MUX2X1_112/B CLKBUF1_6/A OAI21X1_163/Y gnd vdd DFFPOSX1
XDFFPOSX1_215 MUX2X1_157/A CLKBUF1_7/Y OAI21X1_141/Y gnd vdd DFFPOSX1
XNAND2X1_137 MUX2X1_71/A OAI21X1_126/B gnd OAI21X1_121/C vdd NAND2X1
XNAND2X1_126 MUX2X1_23/B OAI21X1_118/B gnd OAI21X1_111/C vdd NAND2X1
XNAND2X1_115 MUX2X1_190/B OAI21X1_97/B gnd NAND2X1_115/Y vdd NAND2X1
XFILL_11_1 gnd vdd FILL
XNAND2X1_148 MUX2X1_109/B OAI21X1_134/B gnd NAND2X1_148/Y vdd NAND2X1
XOAI21X1_109 BUFX4_43/Y OAI21X1_105/B NAND2X1_123/Y gnd OAI21X1_109/Y vdd OAI21X1
XBUFX2_7 BUFX2_7/A gnd dataout[6] vdd BUFX2
XNAND2X1_159 MUX2X1_157/A NAND2X1_160/B gnd NAND2X1_159/Y vdd NAND2X1
XNAND2X1_104 MUX2X1_121/A OAI21X1_90/B gnd OAI21X1_92/C vdd NAND2X1
XMUX2X1_187 MUX2X1_187/A MUX2X1_187/B MUX2X1_5/S gnd MUX2X1_187/Y vdd MUX2X1
XMUX2X1_176 MUX2X1_176/A NAND2X1_16/A BUFX4_36/Y gnd MUX2X1_176/Y vdd MUX2X1
XNAND2X1_2 NAND2X1_2/A NAND2X1_1/B gnd NAND2X1_2/Y vdd NAND2X1
XFILL_8_2_1 gnd vdd FILL
XMUX2X1_154 MUX2X1_154/A MUX2X1_154/B MUX2X1_5/S gnd MUX2X1_156/B vdd MUX2X1
XMUX2X1_132 MUX2X1_132/A MUX2X1_130/Y BUFX4_10/Y gnd AOI22X1_22/D vdd MUX2X1
XMUX2X1_165 MUX2X1_164/Y MUX2X1_165/B BUFX4_13/Y gnd AOI22X1_28/A vdd MUX2X1
XFILL_0_1_1 gnd vdd FILL
XMUX2X1_110 MUX2X1_110/A MUX2X1_110/B BUFX4_36/Y gnd MUX2X1_110/Y vdd MUX2X1
XAOI21X1_7 BUFX4_41/Y NOR2X1_5/B NOR2X1_9/Y gnd AOI21X1_7/Y vdd AOI21X1
XMUX2X1_143 MUX2X1_143/A MUX2X1_143/B BUFX4_36/Y gnd MUX2X1_143/Y vdd MUX2X1
XMUX2X1_121 MUX2X1_121/A MUX2X1_121/B MUX2X1_5/S gnd MUX2X1_121/Y vdd MUX2X1
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XFILL_16_1_1 gnd vdd FILL
XDFFPOSX1_2 MUX2X1_31/A CLKBUF1_28/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XAOI21X1_26 AOI21X1_26/A AOI21X1_26/B INVX4_1/Y gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_37 BUFX4_1/Y AND2X2_4/Y NOR2X1_39/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_15 BUFX4_43/Y AND2X2_2/Y NOR2X1_17/Y gnd AOI21X1_15/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_48 NOR2X1_42/A CLKBUF1_23/A AOI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 MUX2X1_52/B CLKBUF1_2/A OAI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 MUX2X1_34/B CLKBUF1_40/Y OAI21X1_208/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 MUX2X1_154/A CLKBUF1_7/A OAI21X1_197/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 MUX2X1_116/A CLKBUF1_15/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XDFFPOSX1_249 MUX2X1_17/B CLKBUF1_32/A AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_216 MUX2X1_181/A CLKBUF1_2/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_227 MUX2X1_62/A CLKBUF1_24/Y OAI21X1_153/Y gnd vdd DFFPOSX1
XDFFPOSX1_205 MUX2X1_109/B CLKBUF1_35/Y OAI21X1_131/Y gnd vdd DFFPOSX1
XDFFPOSX1_238 MUX2X1_136/B CLKBUF1_9/A OAI21X1_164/Y gnd vdd DFFPOSX1
XBUFX2_8 BUFX2_8/A gnd dataout[7] vdd BUFX2
XMUX2X1_188 MUX2X1_188/A MUX2X1_188/B MUX2X1_7/S gnd MUX2X1_189/A vdd MUX2X1
XAOI21X1_8 BUFX4_55/Y NOR2X1_5/B NOR2X1_10/Y gnd AOI21X1_8/Y vdd AOI21X1
XMUX2X1_177 MUX2X1_176/Y MUX2X1_175/Y BUFX4_9/Y gnd AOI22X1_30/A vdd MUX2X1
XNAND2X1_138 MUX2X1_95/A OAI21X1_126/B gnd NAND2X1_138/Y vdd NAND2X1
XNAND2X1_127 MUX2X1_47/B OAI21X1_118/B gnd NAND2X1_127/Y vdd NAND2X1
XMUX2X1_155 MUX2X1_155/A MUX2X1_155/B MUX2X1_7/S gnd MUX2X1_156/A vdd MUX2X1
XNAND2X1_116 AND2X2_2/B AOI22X1_4/C gnd OAI21X1_105/B vdd NAND2X1
XNAND2X1_149 MUX2X1_133/B OAI21X1_134/B gnd NAND2X1_149/Y vdd NAND2X1
XMUX2X1_166 MUX2X1_166/A MUX2X1_166/B MUX2X1_1/S gnd MUX2X1_166/Y vdd MUX2X1
XMUX2X1_100 MUX2X1_100/A NAND2X1_3/A MUX2X1_1/S gnd MUX2X1_100/Y vdd MUX2X1
XMUX2X1_133 MUX2X1_133/A MUX2X1_133/B MUX2X1_1/S gnd MUX2X1_135/B vdd MUX2X1
XNAND2X1_3 NAND2X1_3/A NAND2X1_1/B gnd NAND2X1_3/Y vdd NAND2X1
XMUX2X1_111 MUX2X1_110/Y MUX2X1_109/Y BUFX4_11/Y gnd MUX2X1_111/Y vdd MUX2X1
XMUX2X1_144 MUX2X1_143/Y MUX2X1_142/Y BUFX4_6/Y gnd MUX2X1_144/Y vdd MUX2X1
XMUX2X1_122 NOR2X1_8/A MUX2X1_122/B MUX2X1_7/S gnd MUX2X1_123/A vdd MUX2X1
XNAND2X1_105 MUX2X1_145/A OAI21X1_90/B gnd OAI21X1_93/C vdd NAND2X1
XDFFPOSX1_3 MUX2X1_55/A CLKBUF1_22/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_5/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 BUFX4_56/Y AND2X2_2/Y NOR2X1_18/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_27 AOI21X1_27/A AOI21X1_27/B INVX4_1/Y gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_38 BUFX4_25/Y AND2X2_4/Y NOR2X1_40/Y gnd AOI21X1_38/Y vdd AOI21X1
XOAI21X1_90 BUFX4_49/Y OAI21X1_90/B OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XDFFPOSX1_27 MUX2X1_58/B CLKBUF1_32/A DFFPOSX1_27/D gnd vdd DFFPOSX1
XDFFPOSX1_16 MUX2X1_178/A CLKBUF1_2/A DFFPOSX1_16/D gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XDFFPOSX1_49 MUX2X1_8/A CLKBUF1_31/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XDFFPOSX1_38 MUX2X1_140/A CLKBUF1_9/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XDFFPOSX1_217 MUX2X1_14/B CLKBUF1_31/A OAI21X1_143/Y gnd vdd DFFPOSX1
XDFFPOSX1_228 MUX2X1_86/A CLKBUF1_19/Y OAI21X1_154/Y gnd vdd DFFPOSX1
XDFFPOSX1_206 MUX2X1_133/B CLKBUF1_9/A OAI21X1_132/Y gnd vdd DFFPOSX1
XDFFPOSX1_239 MUX2X1_160/B CLKBUF1_7/A OAI21X1_165/Y gnd vdd DFFPOSX1
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNAND2X1_117 MUX2X1_22/A OAI21X1_105/B gnd NAND2X1_117/Y vdd NAND2X1
XNAND2X1_128 MUX2X1_71/B OAI21X1_118/B gnd OAI21X1_113/C vdd NAND2X1
XNAND2X1_106 MUX2X1_169/A OAI21X1_90/B gnd OAI21X1_94/C vdd NAND2X1
XAOI21X1_9 BUFX4_19/Y AND2X2_2/Y NOR2X1_11/Y gnd AOI21X1_9/Y vdd AOI21X1
XNAND2X1_4 NAND2X1_4/A NAND2X1_1/B gnd OAI21X1_4/C vdd NAND2X1
XNAND2X1_139 MUX2X1_119/A OAI21X1_126/B gnd OAI21X1_123/C vdd NAND2X1
XMUX2X1_189 MUX2X1_189/A MUX2X1_187/Y BUFX4_13/Y gnd AOI22X1_32/A vdd MUX2X1
XMUX2X1_178 MUX2X1_178/A MUX2X1_178/B BUFX4_37/Y gnd MUX2X1_178/Y vdd MUX2X1
XDFFPOSX1_4 MUX2X1_79/A CLKBUF1_18/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XMUX2X1_156 MUX2X1_156/A MUX2X1_156/B BUFX4_10/Y gnd AOI22X1_26/D vdd MUX2X1
XMUX2X1_112 NOR2X1_15/A MUX2X1_112/B BUFX4_37/Y gnd MUX2X1_114/B vdd MUX2X1
XMUX2X1_134 MUX2X1_134/A MUX2X1_134/B MUX2X1_2/S gnd MUX2X1_134/Y vdd MUX2X1
XMUX2X1_167 MUX2X1_167/A MUX2X1_167/B MUX2X1_2/S gnd MUX2X1_168/A vdd MUX2X1
XNOR2X1_7 NOR2X1_7/A NOR2X1_5/B gnd NOR2X1_7/Y vdd NOR2X1
XMUX2X1_101 NAND2X1_40/A NAND2X1_58/A MUX2X1_2/S gnd MUX2X1_102/A vdd MUX2X1
XMUX2X1_123 MUX2X1_123/A MUX2X1_121/Y BUFX4_7/Y gnd MUX2X1_123/Y vdd MUX2X1
XMUX2X1_145 MUX2X1_145/A MUX2X1_145/B BUFX4_37/Y gnd MUX2X1_145/Y vdd MUX2X1
XAOI21X1_17 BUFX4_21/Y AND2X2_3/Y NOR2X1_21/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 AOI21X1_28/A AOI21X1_28/B INVX4_1/Y gnd AOI21X1_28/Y vdd AOI21X1
XAOI21X1_39 BUFX4_40/Y AND2X2_4/Y NOR2X1_41/Y gnd AOI21X1_39/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_80 BUFX4_51/Y NAND2X1_97/B NAND2X1_91/Y gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 BUFX4_3/Y OAI21X1_90/B OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XFILL_23_2_1 gnd vdd FILL
XDFFPOSX1_17 MUX2X1_11/A CLKBUF1_29/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XDFFPOSX1_28 MUX2X1_82/B CLKBUF1_38/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XDFFPOSX1_39 MUX2X1_164/A CLKBUF1_7/Y OAI21X1_221/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XDFFPOSX1_218 MUX2X1_38/B CLKBUF1_31/A OAI21X1_144/Y gnd vdd DFFPOSX1
XDFFPOSX1_207 MUX2X1_157/B CLKBUF1_7/A OAI21X1_133/Y gnd vdd DFFPOSX1
XDFFPOSX1_229 MUX2X1_110/A CLKBUF1_13/Y OAI21X1_155/Y gnd vdd DFFPOSX1
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_19_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND2X1_129 MUX2X1_95/B OAI21X1_118/B gnd NAND2X1_129/Y vdd NAND2X1
XNAND2X1_107 AOI22X1_4/C NOR2X1_33/Y gnd OAI21X1_97/B vdd NAND2X1
XNAND2X1_118 MUX2X1_46/A OAI21X1_105/B gnd OAI21X1_104/C vdd NAND2X1
XMUX2X1_90 MUX2X1_89/Y MUX2X1_90/B BUFX4_12/Y gnd MUX2X1_90/Y vdd MUX2X1
XNAND2X1_5 NAND2X1_5/A NAND2X1_1/B gnd OAI21X1_5/C vdd NAND2X1
XMUX2X1_179 MUX2X1_179/A MUX2X1_179/B INVX1_3/A gnd MUX2X1_180/A vdd MUX2X1
XMUX2X1_124 MUX2X1_124/A NAND2X1_4/A MUX2X1_8/S gnd MUX2X1_126/B vdd MUX2X1
XMUX2X1_168 MUX2X1_168/A MUX2X1_166/Y BUFX4_6/Y gnd MUX2X1_168/Y vdd MUX2X1
XMUX2X1_157 MUX2X1_157/A MUX2X1_157/B MUX2X1_8/S gnd MUX2X1_159/B vdd MUX2X1
XDFFPOSX1_5 MUX2X1_103/A CLKBUF1_16/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XMUX2X1_146 NOR2X1_9/A MUX2X1_146/B INVX1_3/A gnd MUX2X1_146/Y vdd MUX2X1
XMUX2X1_102 MUX2X1_102/A MUX2X1_100/Y BUFX4_8/Y gnd MUX2X1_102/Y vdd MUX2X1
XMUX2X1_135 MUX2X1_134/Y MUX2X1_135/B BUFX4_11/Y gnd MUX2X1_135/Y vdd MUX2X1
XMUX2X1_113 NOR2X1_39/A NOR2X1_25/A INVX1_3/A gnd MUX2X1_113/Y vdd MUX2X1
XAOI21X1_18 BUFX4_50/Y AND2X2_3/Y NOR2X1_22/Y gnd AOI21X1_18/Y vdd AOI21X1
XNOR2X1_8 NOR2X1_8/A NOR2X1_5/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_29 AOI21X1_29/A AOI21X1_29/B INVX4_1/Y gnd AOI21X1_29/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_70 BUFX4_56/Y NAND2X1_79/B OAI21X1_70/C gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_81 BUFX4_16/Y NAND2X1_97/B OAI21X1_81/C gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_92 BUFX4_24/Y OAI21X1_90/B OAI21X1_92/C gnd OAI21X1_92/Y vdd OAI21X1
XDFFPOSX1_18 MUX2X1_35/A CLKBUF1_26/Y DFFPOSX1_18/D gnd vdd DFFPOSX1
XDFFPOSX1_29 MUX2X1_106/B CLKBUF1_6/A OAI21X1_211/Y gnd vdd DFFPOSX1
XDFFPOSX1_208 MUX2X1_181/B CLKBUF1_2/A OAI21X1_134/Y gnd vdd DFFPOSX1
XDFFPOSX1_219 MUX2X1_62/B CLKBUF1_2/A OAI21X1_145/Y gnd vdd DFFPOSX1
XNAND2X1_119 MUX2X1_70/A OAI21X1_105/B gnd NAND2X1_119/Y vdd NAND2X1
XNAND2X1_108 MUX2X1_22/B OAI21X1_97/B gnd OAI21X1_95/C vdd NAND2X1
XNAND2X1_6 NAND2X1_6/A NAND2X1_1/B gnd OAI21X1_6/C vdd NAND2X1
XNOR2X1_40 NOR2X1_40/A AND2X2_4/Y gnd NOR2X1_40/Y vdd NOR2X1
XFILL_21_3_0 gnd vdd FILL
XMUX2X1_169 MUX2X1_169/A NAND2X1_25/A MUX2X1_4/S gnd MUX2X1_171/B vdd MUX2X1
XMUX2X1_91 MUX2X1_91/A MUX2X1_91/B MUX2X1_8/S gnd MUX2X1_93/B vdd MUX2X1
XMUX2X1_80 MUX2X1_80/A MUX2X1_80/B INVX1_3/A gnd MUX2X1_81/A vdd MUX2X1
XDFFPOSX1_6 MUX2X1_127/A CLKBUF1_12/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XMUX2X1_158 MUX2X1_158/A MUX2X1_158/B BUFX4_35/Y gnd MUX2X1_158/Y vdd MUX2X1
XMUX2X1_103 MUX2X1_103/A MUX2X1_103/B MUX2X1_4/S gnd MUX2X1_103/Y vdd MUX2X1
XMUX2X1_125 MUX2X1_125/A MUX2X1_125/B BUFX4_35/Y gnd MUX2X1_125/Y vdd MUX2X1
XMUX2X1_136 NOR2X1_16/A MUX2X1_136/B MUX2X1_4/S gnd MUX2X1_136/Y vdd MUX2X1
XMUX2X1_147 MUX2X1_146/Y MUX2X1_145/Y BUFX4_7/Y gnd MUX2X1_147/Y vdd MUX2X1
XMUX2X1_114 MUX2X1_113/Y MUX2X1_114/B BUFX4_12/Y gnd MUX2X1_114/Y vdd MUX2X1
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_5/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 BUFX4_15/Y AND2X2_3/Y NOR2X1_23/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_71 BUFX4_21/Y NAND2X1_88/B OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_82 BUFX4_46/Y NAND2X1_97/B NAND2X1_93/Y gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_60 BUFX4_26/Y NAND2X1_65/B NAND2X1_68/Y gnd OAI21X1_60/Y vdd OAI21X1
XFILL_8_1 gnd vdd FILL
XOAI21X1_93 BUFX4_41/Y OAI21X1_90/B OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_230 BUFX4_58/Y NAND2X1_279/B NAND2X1_281/Y gnd OAI21X1_230/Y vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XDFFPOSX1_19 MUX2X1_59/A CLKBUF1_22/Y OAI21X1_201/Y gnd vdd DFFPOSX1
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_280 MUX2X1_152/A NAND2X1_279/B gnd NAND2X1_280/Y vdd NAND2X1
XFILL_23_0_0 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XDFFPOSX1_209 MUX2X1_13/A CLKBUF1_31/Y OAI21X1_135/Y gnd vdd DFFPOSX1
XNAND2X1_109 MUX2X1_46/B OAI21X1_97/B gnd OAI21X1_96/C vdd NAND2X1
XNOR2X1_41 NOR2X1_41/A AND2X2_4/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_30 NOR2X1_1/A NOR2X1_30/B gnd AND2X2_2/B vdd NOR2X1
XNAND2X1_7 BUFX4_6/Y INVX1_3/Y gnd NOR2X1_1/B vdd NAND2X1
XMUX2X1_70 MUX2X1_70/A MUX2X1_70/B MUX2X1_4/S gnd MUX2X1_72/B vdd MUX2X1
XFILL_21_3_1 gnd vdd FILL
XMUX2X1_92 MUX2X1_92/A MUX2X1_92/B BUFX4_35/Y gnd MUX2X1_93/A vdd MUX2X1
XMUX2X1_81 MUX2X1_81/A MUX2X1_81/B BUFX4_9/Y gnd MUX2X1_81/Y vdd MUX2X1
XMUX2X1_115 MUX2X1_115/A NAND2X1_76/A BUFX4_39/Y gnd MUX2X1_117/B vdd MUX2X1
XMUX2X1_137 NOR2X1_40/A NOR2X1_26/A MUX2X1_5/S gnd MUX2X1_138/A vdd MUX2X1
XMUX2X1_126 MUX2X1_125/Y MUX2X1_126/B BUFX4_8/Y gnd AOI22X1_21/D vdd MUX2X1
XMUX2X1_148 MUX2X1_148/A NAND2X1_5/A BUFX4_39/Y gnd MUX2X1_148/Y vdd MUX2X1
XMUX2X1_159 MUX2X1_158/Y MUX2X1_159/B BUFX4_11/Y gnd MUX2X1_159/Y vdd MUX2X1
XMUX2X1_104 MUX2X1_104/A MUX2X1_104/B MUX2X1_5/S gnd MUX2X1_105/A vdd MUX2X1
XFILL_12_3_1 gnd vdd FILL
XDFFPOSX1_7 MUX2X1_151/A CLKBUF1_8/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XOAI21X1_94 BUFX4_59/Y OAI21X1_90/B OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_50 BUFX4_47/Y OAI21X1_52/B OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_72 BUFX4_54/Y NAND2X1_88/B NAND2X1_82/Y gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_83 BUFX4_2/Y NAND2X1_97/B NAND2X1_94/Y gnd OAI21X1_83/Y vdd OAI21X1
XFILL_8_2 gnd vdd FILL
XOAI21X1_61 BUFX4_42/Y NAND2X1_65/B NAND2X1_69/Y gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_231 BUFX4_22/Y NAND2X1_1/B NAND2X1_284/Y gnd DFFPOSX1_57/D vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_220 BUFX4_24/Y NAND2X1_267/B OAI21X1_220/C gnd DFFPOSX1_38/D vdd OAI21X1
XFILL_17_2_1 gnd vdd FILL
XNAND2X1_281 MUX2X1_176/A NAND2X1_279/B gnd NAND2X1_281/Y vdd NAND2X1
XFILL_9_3_1 gnd vdd FILL
XNAND2X1_270 MUX2X1_164/A NAND2X1_267/B gnd OAI21X1_221/C vdd NAND2X1
XCLKBUF1_40 clk gnd CLKBUF1_40/Y vdd CLKBUF1
XFILL_23_0_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_42 NOR2X1_42/A AND2X2_4/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_31 OR2X2_1/B NOR2X1_31/B gnd AOI22X1_2/C vdd NOR2X1
XNOR2X1_20 address[2] OR2X2_1/A gnd AOI22X1_3/B vdd NOR2X1
XMUX2X1_71 MUX2X1_71/A MUX2X1_71/B MUX2X1_5/S gnd MUX2X1_72/A vdd MUX2X1
XMUX2X1_60 MUX2X1_59/Y MUX2X1_60/B BUFX4_10/Y gnd MUX2X1_60/Y vdd MUX2X1
XMUX2X1_93 MUX2X1_93/A MUX2X1_93/B BUFX4_13/Y gnd MUX2X1_93/Y vdd MUX2X1
XMUX2X1_82 MUX2X1_82/A MUX2X1_82/B BUFX4_39/Y gnd MUX2X1_84/B vdd MUX2X1
XNAND2X1_8 AOI22X1_2/B NOR2X1_1/Y gnd OAI21X1_7/B vdd NAND2X1
XMUX2X1_116 MUX2X1_116/A NAND2X1_94/A MUX2X1_1/S gnd MUX2X1_116/Y vdd MUX2X1
XMUX2X1_138 MUX2X1_138/A MUX2X1_136/Y BUFX4_12/Y gnd MUX2X1_138/Y vdd MUX2X1
XMUX2X1_127 MUX2X1_127/A MUX2X1_127/B BUFX4_36/Y gnd MUX2X1_127/Y vdd MUX2X1
XMUX2X1_105 MUX2X1_105/A MUX2X1_103/Y BUFX4_9/Y gnd MUX2X1_105/Y vdd MUX2X1
XMUX2X1_149 MUX2X1_149/A NAND2X1_60/A MUX2X1_1/S gnd MUX2X1_149/Y vdd MUX2X1
XDFFPOSX1_8 DFFPOSX1_8/Q CLKBUF1_3/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XOAI21X1_95 BUFX4_20/Y OAI21X1_97/B OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_73 BUFX4_14/Y NAND2X1_88/B OAI21X1_73/C gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_62 BUFX4_59/Y NAND2X1_65/B NAND2X1_70/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_210 BUFX4_45/Y NAND2X1_256/B NAND2X1_257/Y gnd DFFPOSX1_28/D vdd OAI21X1
XOAI21X1_40 BUFX4_51/Y NAND2X1_50/B OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_84 BUFX4_26/Y NAND2X1_97/B NAND2X1_95/Y gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_51 BUFX4_4/Y OAI21X1_52/B NAND2X1_58/Y gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_221 BUFX4_42/Y NAND2X1_267/B OAI21X1_221/C gnd OAI21X1_221/Y vdd OAI21X1
XNAND2X1_271 MUX2X1_188/A NAND2X1_267/B gnd NAND2X1_271/Y vdd NAND2X1
XNAND2X1_282 INVX1_4/Y INVX1_1/Y gnd NOR2X1_2/B vdd NAND2X1
XOAI21X1_232 BUFX4_51/Y NAND2X1_1/B OAI21X1_232/C gnd OAI21X1_232/Y vdd OAI21X1
XNAND2X1_260 MUX2X1_154/B NAND2X1_256/B gnd OAI21X1_213/C vdd NAND2X1
XDFFPOSX1_190 MUX2X1_143/B CLKBUF1_9/A OAI21X1_116/Y gnd vdd DFFPOSX1
XCLKBUF1_41 clk gnd CLKBUF1_32/A vdd CLKBUF1
XCLKBUF1_30 CLKBUF1_32/A gnd CLKBUF1_30/Y vdd CLKBUF1
XFILL_18_1 gnd vdd FILL
XNOR2X1_21 MUX2X1_17/B AND2X2_3/Y gnd NOR2X1_21/Y vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_5/B gnd NOR2X1_10/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNOR2X1_43 OR2X2_1/B NOR2X1_2/B gnd AOI22X1_9/C vdd NOR2X1
XNOR2X1_32 NOR2X1_1/A NOR2X1_32/B gnd AND2X2_4/B vdd NOR2X1
XMUX2X1_50 NOR2X1_5/A MUX2X1_50/B MUX2X1_1/S gnd MUX2X1_51/A vdd MUX2X1
XMUX2X1_72 MUX2X1_72/A MUX2X1_72/B BUFX4_6/Y gnd MUX2X1_72/Y vdd MUX2X1
XNAND2X1_9 MUX2X1_8/B OAI21X1_7/B gnd NAND2X1_9/Y vdd NAND2X1
XMUX2X1_61 MUX2X1_61/A MUX2X1_61/B BUFX4_36/Y gnd MUX2X1_63/B vdd MUX2X1
XMUX2X1_94 MUX2X1_94/A MUX2X1_94/B BUFX4_36/Y gnd MUX2X1_94/Y vdd MUX2X1
XMUX2X1_83 MUX2X1_83/A MUX2X1_83/B MUX2X1_1/S gnd MUX2X1_83/Y vdd MUX2X1
XDFFPOSX1_9 MUX2X1_10/A CLKBUF1_31/A DFFPOSX1_9/D gnd vdd DFFPOSX1
XMUX2X1_139 NAND2X1_86/A NAND2X1_77/A MUX2X1_7/S gnd MUX2X1_139/Y vdd MUX2X1
XMUX2X1_117 MUX2X1_116/Y MUX2X1_117/B BUFX4_13/Y gnd AOI22X1_20/A vdd MUX2X1
XMUX2X1_106 MUX2X1_106/A MUX2X1_106/B MUX2X1_7/S gnd MUX2X1_108/B vdd MUX2X1
XMUX2X1_128 MUX2X1_128/A MUX2X1_128/B BUFX4_37/Y gnd MUX2X1_129/A vdd MUX2X1
XFILL_21_1_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_63 BUFX4_21/Y NAND2X1_79/B OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_41 BUFX4_15/Y NAND2X1_50/B NAND2X1_47/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_30 BUFX4_57/Y NAND2X1_27/B OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_74 BUFX4_45/Y NAND2X1_88/B OAI21X1_74/C gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 BUFX4_53/Y OAI21X1_97/B OAI21X1_96/C gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_52 BUFX4_28/Y OAI21X1_52/B OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_85 BUFX4_44/Y NAND2X1_97/B NAND2X1_96/Y gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_222 BUFX4_55/Y NAND2X1_267/B NAND2X1_271/Y gnd DFFPOSX1_40/D vdd OAI21X1
XNAND2X1_261 MUX2X1_178/B NAND2X1_256/B gnd OAI21X1_214/C vdd NAND2X1
XNAND2X1_272 address[3] address[4] gnd OR2X2_1/A vdd NAND2X1
XDFFPOSX1_180 MUX2X1_94/A CLKBUF1_18/Y OAI21X1_106/Y gnd vdd DFFPOSX1
XOAI21X1_200 BUFX4_54/Y OAI21X1_201/B NAND2X1_245/Y gnd DFFPOSX1_18/D vdd OAI21X1
XNAND2X1_283 NOR2X1_33/Y AOI22X1_9/C gnd NAND2X1_1/B vdd NAND2X1
XOAI21X1_211 BUFX4_1/Y NAND2X1_256/B OAI21X1_211/C gnd OAI21X1_211/Y vdd OAI21X1
XNAND2X1_250 MUX2X1_155/A OAI21X1_201/B gnd NAND2X1_250/Y vdd NAND2X1
XDFFPOSX1_191 MUX2X1_167/B CLKBUF1_9/A OAI21X1_117/Y gnd vdd DFFPOSX1
XFILL_6_1 gnd vdd FILL
XCLKBUF1_31 CLKBUF1_31/A gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_42 clk gnd CLKBUF1_31/A vdd CLKBUF1
XCLKBUF1_20 CLKBUF1_43/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XFILL_1_0_0 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XFILL_18_2 gnd vdd FILL
XNOR2X1_11 MUX2X1_16/A AND2X2_2/Y gnd NOR2X1_11/Y vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_22 MUX2X1_41/B AND2X2_3/Y gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_33 NOR2X1_1/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XMUX2X1_51 MUX2X1_51/A MUX2X1_49/Y BUFX4_7/Y gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_62 MUX2X1_62/A MUX2X1_62/B BUFX4_37/Y gnd MUX2X1_62/Y vdd MUX2X1
XMUX2X1_40 MUX2X1_40/A MUX2X1_40/B MUX2X1_7/S gnd MUX2X1_42/B vdd MUX2X1
XMUX2X1_95 MUX2X1_95/A MUX2X1_95/B BUFX4_37/Y gnd MUX2X1_96/A vdd MUX2X1
XMUX2X1_84 MUX2X1_83/Y MUX2X1_84/B BUFX4_10/Y gnd MUX2X1_84/Y vdd MUX2X1
XMUX2X1_73 MUX2X1_73/A MUX2X1_73/B MUX2X1_7/S gnd MUX2X1_73/Y vdd MUX2X1
XMUX2X1_129 MUX2X1_129/A MUX2X1_127/Y BUFX4_9/Y gnd AOI22X1_22/A vdd MUX2X1
XMUX2X1_118 MUX2X1_118/A MUX2X1_118/B MUX2X1_2/S gnd MUX2X1_118/Y vdd MUX2X1
XMUX2X1_107 MUX2X1_107/A MUX2X1_107/B MUX2X1_8/S gnd MUX2X1_107/Y vdd MUX2X1
XFILL_21_1_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XOAI21X1_97 BUFX4_16/Y OAI21X1_97/B OAI21X1_97/C gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_86 BUFX4_55/Y NAND2X1_97/B OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_31 BUFX4_22/Y OAI21X1_38/B OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_42 BUFX4_49/Y NAND2X1_50/B NAND2X1_48/Y gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_64 BUFX4_54/Y NAND2X1_79/B NAND2X1_73/Y gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_75 BUFX4_2/Y NAND2X1_88/B OAI21X1_75/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_20 BUFX4_24/Y OAI21X1_18/B OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_53 BUFX4_42/Y OAI21X1_52/B NAND2X1_60/Y gnd OAI21X1_53/Y vdd OAI21X1
XDFFPOSX1_192 MUX2X1_191/B CLKBUF1_33/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XNAND2X1_284 MUX2X1_4/B NAND2X1_1/B gnd NAND2X1_284/Y vdd NAND2X1
XOAI21X1_223 BUFX4_22/Y NAND2X1_279/B NAND2X1_274/Y gnd DFFPOSX1_49/D vdd OAI21X1
XOAI21X1_201 BUFX4_14/Y OAI21X1_201/B NAND2X1_246/Y gnd OAI21X1_201/Y vdd OAI21X1
XNAND2X1_251 MUX2X1_179/A OAI21X1_201/B gnd NAND2X1_251/Y vdd NAND2X1
XNAND2X1_262 address[4] INVX1_4/Y gnd NOR2X1_19/B vdd NAND2X1
XDFFPOSX1_170 MUX2X1_46/B CLKBUF1_31/A OAI21X1_96/Y gnd vdd DFFPOSX1
XNAND2X1_273 AND2X2_4/B AOI22X1_2/B gnd NAND2X1_279/B vdd NAND2X1
XNAND2X1_240 MUX2X1_154/A OAI21X1_193/B gnd OAI21X1_197/C vdd NAND2X1
XOAI21X1_212 BUFX4_25/Y NAND2X1_256/B NAND2X1_259/Y gnd DFFPOSX1_30/D vdd OAI21X1
XDFFPOSX1_181 MUX2X1_118/A CLKBUF1_13/Y OAI21X1_107/Y gnd vdd DFFPOSX1
XFILL_6_2 gnd vdd FILL
XCLKBUF1_21 CLKBUF1_23/A gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_32 CLKBUF1_32/A gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_43 clk gnd CLKBUF1_43/Y vdd CLKBUF1
XCLKBUF1_10 CLKBUF1_18/A gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XNOR2X1_12 MUX2X1_40/A AND2X2_2/Y gnd NOR2X1_12/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A AND2X2_3/Y gnd NOR2X1_23/Y vdd NOR2X1
XMUX2X1_52 MUX2X1_52/A MUX2X1_52/B MUX2X1_2/S gnd MUX2X1_54/B vdd MUX2X1
XMUX2X1_63 MUX2X1_62/Y MUX2X1_63/B BUFX4_11/Y gnd MUX2X1_63/Y vdd MUX2X1
XMUX2X1_41 MUX2X1_41/A MUX2X1_41/B MUX2X1_8/S gnd MUX2X1_42/A vdd MUX2X1
XNOR2X1_34 address[2] NOR2X1_19/B gnd AOI22X1_4/B vdd NOR2X1
XMUX2X1_30 MUX2X1_30/A MUX2X1_28/Y BUFX4_8/Y gnd MUX2X1_30/Y vdd MUX2X1
XFILL_23_1 gnd vdd FILL
XMUX2X1_96 MUX2X1_96/A MUX2X1_94/Y BUFX4_6/Y gnd MUX2X1_96/Y vdd MUX2X1
XMUX2X1_85 MUX2X1_85/A MUX2X1_85/B MUX2X1_2/S gnd MUX2X1_87/B vdd MUX2X1
XMUX2X1_74 NOR2X1_6/A MUX2X1_74/B MUX2X1_8/S gnd MUX2X1_75/A vdd MUX2X1
XMUX2X1_119 MUX2X1_119/A MUX2X1_119/B MUX2X1_4/S gnd MUX2X1_120/A vdd MUX2X1
XMUX2X1_108 MUX2X1_107/Y MUX2X1_108/B BUFX4_10/Y gnd MUX2X1_108/Y vdd MUX2X1
XOAI21X1_54 BUFX4_59/Y OAI21X1_52/B OAI21X1_54/C gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_65 BUFX4_14/Y NAND2X1_79/B NAND2X1_74/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_87 BUFX4_19/Y OAI21X1_90/B OAI21X1_87/C gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_98 BUFX4_45/Y OAI21X1_97/B OAI21X1_98/C gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_10 BUFX4_48/Y OAI21X1_7/B OAI21X1_10/C gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_32 BUFX4_53/Y OAI21X1_38/B OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_76 BUFX4_25/Y NAND2X1_88/B NAND2X1_86/Y gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_43 BUFX4_5/Y NAND2X1_50/B NAND2X1_49/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_21 BUFX4_41/Y OAI21X1_18/B NAND2X1_24/Y gnd OAI21X1_21/Y vdd OAI21X1
XDFFPOSX1_160 MUX2X1_188/B CLKBUF1_33/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_171 MUX2X1_70/B CLKBUF1_23/A OAI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_193 MUX2X1_23/A CLKBUF1_32/Y OAI21X1_119/Y gnd vdd DFFPOSX1
XNAND2X1_241 MUX2X1_178/A OAI21X1_193/B gnd OAI21X1_198/C vdd NAND2X1
XOAI21X1_224 BUFX4_52/Y NAND2X1_279/B OAI21X1_224/C gnd DFFPOSX1_50/D vdd OAI21X1
XOAI21X1_202 BUFX4_48/Y OAI21X1_201/B NAND2X1_247/Y gnd DFFPOSX1_20/D vdd OAI21X1
XOAI21X1_213 BUFX4_40/Y NAND2X1_256/B OAI21X1_213/C gnd DFFPOSX1_31/D vdd OAI21X1
XNAND2X1_230 MUX2X1_127/A OAI21X1_183/B gnd NAND2X1_230/Y vdd NAND2X1
XDFFPOSX1_182 MUX2X1_142/A CLKBUF1_12/Y OAI21X1_108/Y gnd vdd DFFPOSX1
XNAND2X1_252 INVX1_3/Y INVX1_2/Y gnd NOR2X1_33/B vdd NAND2X1
XNAND2X1_274 MUX2X1_8/A NAND2X1_279/B gnd NAND2X1_274/Y vdd NAND2X1
XNAND2X1_285 MUX2X1_28/B NAND2X1_1/B gnd OAI21X1_232/C vdd NAND2X1
XNAND2X1_263 AND2X2_4/B AOI22X1_4/B gnd NAND2X1_267/B vdd NAND2X1
XFILL_6_3 gnd vdd FILL
XCLKBUF1_22 CLKBUF1_32/A gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_44 clk gnd CLKBUF1_2/A vdd CLKBUF1
XCLKBUF1_33 clk gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_11 CLKBUF1_9/A gnd CLKBUF1_11/Y vdd CLKBUF1
XFILL_10_2_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_18_3_0 gnd vdd FILL
XNOR2X1_35 NOR2X1_35/A AND2X2_4/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_13 MUX2X1_64/A AND2X2_2/Y gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A AND2X2_3/Y gnd NOR2X1_24/Y vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XMUX2X1_20 MUX2X1_20/A MUX2X1_20/B MUX2X1_4/S gnd MUX2X1_20/Y vdd MUX2X1
XMUX2X1_64 MUX2X1_64/A MUX2X1_64/B INVX1_3/A gnd MUX2X1_66/B vdd MUX2X1
XMUX2X1_53 MUX2X1_53/A MUX2X1_53/B MUX2X1_4/S gnd MUX2X1_54/A vdd MUX2X1
XFILL_16_1 gnd vdd FILL
XMUX2X1_31 MUX2X1_31/A MUX2X1_31/B INVX1_3/A gnd MUX2X1_33/B vdd MUX2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_42/B BUFX4_12/Y gnd AOI22X1_7/D vdd MUX2X1
XMUX2X1_86 MUX2X1_86/A MUX2X1_86/B MUX2X1_4/S gnd MUX2X1_86/Y vdd MUX2X1
XMUX2X1_75 MUX2X1_75/A MUX2X1_73/Y BUFX4_7/Y gnd MUX2X1_75/Y vdd MUX2X1
XMUX2X1_109 MUX2X1_109/A MUX2X1_109/B BUFX4_35/Y gnd MUX2X1_109/Y vdd MUX2X1
XMUX2X1_97 MUX2X1_97/A MUX2X1_97/B INVX1_3/A gnd MUX2X1_97/Y vdd MUX2X1
XNAND2X1_90 MUX2X1_20/B NAND2X1_97/B gnd OAI21X1_79/C vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_33 BUFX4_15/Y OAI21X1_38/B OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_22 BUFX4_58/Y OAI21X1_18/B NAND2X1_25/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_55 BUFX4_19/Y NAND2X1_65/B NAND2X1_63/Y gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_66 BUFX4_45/Y NAND2X1_79/B OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_88 BUFX4_52/Y OAI21X1_90/B OAI21X1_88/C gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_77 BUFX4_40/Y NAND2X1_88/B NAND2X1_87/Y gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_44 BUFX4_26/Y NAND2X1_50/B NAND2X1_50/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_99 BUFX4_4/Y OAI21X1_97/B OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_11 BUFX4_1/Y OAI21X1_7/B OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_225 BUFX4_18/Y NAND2X1_279/B NAND2X1_276/Y gnd DFFPOSX1_51/D vdd OAI21X1
XOAI21X1_214 BUFX4_57/Y NAND2X1_256/B OAI21X1_214/C gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_203 BUFX4_1/Y OAI21X1_201/B NAND2X1_248/Y gnd OAI21X1_203/Y vdd OAI21X1
XNAND2X1_264 MUX2X1_20/A NAND2X1_267/B gnd NAND2X1_264/Y vdd NAND2X1
XNAND2X1_220 AOI22X1_31/Y AOI22X1_32/Y gnd OAI21X1_182/B vdd NAND2X1
XDFFPOSX1_161 MUX2X1_1/A CLKBUF1_29/Y OAI21X1_87/Y gnd vdd DFFPOSX1
XDFFPOSX1_172 MUX2X1_94/B CLKBUF1_2/A OAI21X1_98/Y gnd vdd DFFPOSX1
XNAND2X1_275 MUX2X1_32/A NAND2X1_279/B gnd OAI21X1_224/C vdd NAND2X1
XDFFPOSX1_194 MUX2X1_47/A CLKBUF1_27/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XNAND2X1_253 AOI22X1_2/C NOR2X1_33/Y gnd NAND2X1_256/B vdd NAND2X1
XDFFPOSX1_150 NAND2X1_86/A CLKBUF1_10/Y OAI21X1_76/Y gnd vdd DFFPOSX1
XNAND2X1_242 BUFX4_37/Y BUFX4_8/Y gnd NOR2X1_32/B vdd NAND2X1
XDFFPOSX1_183 MUX2X1_166/A CLKBUF1_6/Y OAI21X1_109/Y gnd vdd DFFPOSX1
XNAND2X1_231 MUX2X1_151/A OAI21X1_183/B gnd OAI21X1_189/C vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XCLKBUF1_23 CLKBUF1_23/A gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_34 clk gnd CLKBUF1_1/A vdd CLKBUF1
XCLKBUF1_45 clk gnd CLKBUF1_9/A vdd CLKBUF1
XCLKBUF1_12 CLKBUF1_9/A gnd CLKBUF1_12/Y vdd CLKBUF1
XFILL_4_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_36 MUX2X1_41/A AND2X2_4/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_14 NOR2X1_14/A AND2X2_2/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A AND2X2_3/Y gnd NOR2X1_25/Y vdd NOR2X1
XFILL_23_3 gnd vdd FILL
XMUX2X1_21 MUX2X1_20/Y MUX2X1_19/Y BUFX4_13/Y gnd AOI22X1_4/A vdd MUX2X1
XMUX2X1_65 MUX2X1_65/A NOR2X1_23/A BUFX4_39/Y gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_54 MUX2X1_54/A MUX2X1_54/B BUFX4_8/Y gnd AOI22X1_9/D vdd MUX2X1
XMUX2X1_10 MUX2X1_10/A MUX2X1_10/B BUFX4_35/Y gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_32 MUX2X1_32/A MUX2X1_32/B BUFX4_39/Y gnd MUX2X1_32/Y vdd MUX2X1
XMUX2X1_87 MUX2X1_86/Y MUX2X1_87/B BUFX4_11/Y gnd MUX2X1_87/Y vdd MUX2X1
XMUX2X1_76 MUX2X1_76/A NAND2X1_2/A BUFX4_35/Y gnd MUX2X1_78/B vdd MUX2X1
XMUX2X1_43 MUX2X1_43/A MUX2X1_43/B BUFX4_35/Y gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_98 NOR2X1_7/A MUX2X1_98/B BUFX4_39/Y gnd MUX2X1_98/Y vdd MUX2X1
XNAND2X1_91 MUX2X1_44/B NAND2X1_97/B gnd NAND2X1_91/Y vdd NAND2X1
XNAND2X1_80 AND2X2_2/B AOI22X1_4/B gnd NAND2X1_88/B vdd NAND2X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_23 BUFX4_21/Y NAND2X1_27/B OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_34 BUFX4_47/Y OAI21X1_38/B NAND2X1_39/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_12 BUFX4_25/Y OAI21X1_7/B OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_45 BUFX4_42/Y NAND2X1_50/B OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_78 BUFX4_56/Y NAND2X1_88/B OAI21X1_78/C gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_215 BUFX4_20/Y NAND2X1_267/B NAND2X1_264/Y gnd DFFPOSX1_33/D vdd OAI21X1
XOAI21X1_89 BUFX4_18/Y OAI21X1_90/B OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XOAI21X1_226 BUFX4_48/Y NAND2X1_279/B OAI21X1_226/C gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_204 BUFX4_26/Y OAI21X1_201/B NAND2X1_249/Y gnd DFFPOSX1_22/D vdd OAI21X1
XOAI21X1_67 BUFX4_2/Y NAND2X1_79/B NAND2X1_76/Y gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_56 BUFX4_54/Y NAND2X1_65/B NAND2X1_64/Y gnd OAI21X1_56/Y vdd OAI21X1
XDFFPOSX1_195 MUX2X1_71/A CLKBUF1_21/Y OAI21X1_121/Y gnd vdd DFFPOSX1
XDFFPOSX1_184 MUX2X1_190/A CLKBUF1_2/Y OAI21X1_110/Y gnd vdd DFFPOSX1
XNAND2X1_232 DFFPOSX1_8/Q OAI21X1_183/B gnd OAI21X1_190/C vdd NAND2X1
XNAND2X1_276 MUX2X1_56/A NAND2X1_279/B gnd NAND2X1_276/Y vdd NAND2X1
XNAND2X1_254 MUX2X1_10/B NAND2X1_256/B gnd NAND2X1_254/Y vdd NAND2X1
XNAND2X1_221 address[3] INVX1_1/Y gnd NOR2X1_31/B vdd NAND2X1
XDFFPOSX1_140 MUX2X1_91/B CLKBUF1_43/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 MUX2X1_25/A CLKBUF1_26/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XNAND2X1_265 MUX2X1_44/A NAND2X1_267/B gnd NAND2X1_265/Y vdd NAND2X1
XDFFPOSX1_151 MUX2X1_163/A CLKBUF1_5/Y OAI21X1_77/Y gnd vdd DFFPOSX1
XNAND2X1_243 AND2X2_4/B AOI22X1_2/C gnd OAI21X1_201/B vdd NAND2X1
XDFFPOSX1_173 MUX2X1_118/B CLKBUF1_7/A OAI21X1_99/Y gnd vdd DFFPOSX1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_210 AOI22X1_17/Y AOI22X1_18/Y gnd NAND2X1_210/Y vdd NAND2X1
XCLKBUF1_24 CLKBUF1_23/A gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_46 clk gnd CLKBUF1_6/A vdd CLKBUF1
XCLKBUF1_13 CLKBUF1_35/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_35 clk gnd CLKBUF1_35/Y vdd CLKBUF1
XNOR2X1_37 MUX2X1_65/A AND2X2_4/Y gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A AND2X2_3/Y gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_15 NOR2X1_15/A AND2X2_2/Y gnd NOR2X1_15/Y vdd NOR2X1
XMUX2X1_22 MUX2X1_22/A MUX2X1_22/B MUX2X1_5/S gnd MUX2X1_24/B vdd MUX2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B MUX2X1_5/S gnd MUX2X1_57/B vdd MUX2X1
XMUX2X1_66 MUX2X1_65/Y MUX2X1_66/B BUFX4_12/Y gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_11 MUX2X1_11/A MUX2X1_11/B BUFX4_36/Y gnd MUX2X1_11/Y vdd MUX2X1
XMUX2X1_33 MUX2X1_32/Y MUX2X1_33/B BUFX4_9/Y gnd AOI22X1_6/A vdd MUX2X1
XMUX2X1_44 MUX2X1_44/A MUX2X1_44/B BUFX4_36/Y gnd MUX2X1_45/A vdd MUX2X1
XMUX2X1_77 MUX2X1_77/A MUX2X1_77/B BUFX4_36/Y gnd MUX2X1_78/A vdd MUX2X1
XMUX2X1_88 NOR2X1_14/A MUX2X1_88/B MUX2X1_5/S gnd MUX2X1_90/B vdd MUX2X1
XMUX2X1_99 MUX2X1_98/Y MUX2X1_97/Y BUFX4_7/Y gnd MUX2X1_99/Y vdd MUX2X1
XNAND2X1_81 MUX2X1_19/A NAND2X1_88/B gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_92 MUX2X1_68/B NAND2X1_97/B gnd OAI21X1_81/C vdd NAND2X1
XNAND2X1_70 MUX2X1_179/B NAND2X1_65/B gnd NAND2X1_70/Y vdd NAND2X1
XFILL_21_1 gnd vdd FILL
XOAI21X1_79 BUFX4_21/Y NAND2X1_97/B OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_57 BUFX4_14/Y NAND2X1_65/B OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_46 BUFX4_58/Y NAND2X1_50/B OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_24 BUFX4_52/Y NAND2X1_27/B OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_68 BUFX4_26/Y NAND2X1_79/B NAND2X1_77/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_35 BUFX4_5/Y OAI21X1_38/B OAI21X1_35/C gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_13 BUFX4_43/Y OAI21X1_7/B NAND2X1_15/Y gnd OAI21X1_13/Y vdd OAI21X1
XDFFPOSX1_152 MUX2X1_187/A CLKBUF1_1/Y OAI21X1_78/Y gnd vdd DFFPOSX1
XNAND2X1_266 MUX2X1_68/A NAND2X1_267/B gnd OAI21X1_217/C vdd NAND2X1
XDFFPOSX1_185 MUX2X1_23/B CLKBUF1_23/A OAI21X1_111/Y gnd vdd DFFPOSX1
XDFFPOSX1_163 MUX2X1_49/A CLKBUF1_21/Y OAI21X1_89/Y gnd vdd DFFPOSX1
XNAND2X1_244 MUX2X1_11/A OAI21X1_201/B gnd NAND2X1_244/Y vdd NAND2X1
XNAND2X1_200 r_w BUFX2_2/A gnd AOI21X1_26/A vdd NAND2X1
XDFFPOSX1_196 MUX2X1_95/A CLKBUF1_17/Y OAI21X1_122/Y gnd vdd DFFPOSX1
XNAND2X1_277 MUX2X1_80/A NAND2X1_279/B gnd OAI21X1_226/C vdd NAND2X1
XNAND2X1_255 MUX2X1_34/B NAND2X1_256/B gnd NAND2X1_255/Y vdd NAND2X1
XOAI21X1_216 BUFX4_51/Y NAND2X1_267/B NAND2X1_265/Y gnd DFFPOSX1_34/D vdd OAI21X1
XDFFPOSX1_130 MUX2X1_35/B CLKBUF1_26/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_141 NAND2X1_76/A CLKBUF1_6/A OAI21X1_67/Y gnd vdd DFFPOSX1
XNAND2X1_233 AND2X2_2/B AOI22X1_2/C gnd OAI21X1_193/B vdd NAND2X1
XOAI21X1_227 BUFX4_2/Y NAND2X1_279/B OAI21X1_227/C gnd OAI21X1_227/Y vdd OAI21X1
XOAI21X1_205 BUFX4_40/Y OAI21X1_201/B NAND2X1_250/Y gnd DFFPOSX1_23/D vdd OAI21X1
XDFFPOSX1_174 MUX2X1_142/B CLKBUF1_9/A OAI21X1_100/Y gnd vdd DFFPOSX1
XNAND2X1_222 r_w enable gnd NOR2X1_1/A vdd NAND2X1
XNAND2X1_211 AOI22X1_19/Y AOI22X1_20/Y gnd OAI21X1_179/B vdd NAND2X1
XFILL_22_2_0 gnd vdd FILL
XCLKBUF1_25 CLKBUF1_31/A gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_47 clk gnd CLKBUF1_7/A vdd CLKBUF1
XCLKBUF1_14 CLKBUF1_6/A gnd CLKBUF1_14/Y vdd CLKBUF1
XCLKBUF1_36 clk gnd CLKBUF1_4/A vdd CLKBUF1
XFILL_13_2_0 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_16 NOR2X1_16/A AND2X2_2/Y gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A AND2X2_3/Y gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_38 MUX2X1_89/A AND2X2_4/Y gnd NOR2X1_38/Y vdd NOR2X1
XMUX2X1_23 MUX2X1_23/A MUX2X1_23/B MUX2X1_7/S gnd MUX2X1_24/A vdd MUX2X1
XMUX2X1_67 MUX2X1_67/A MUX2X1_67/B MUX2X1_1/S gnd MUX2X1_67/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_56 MUX2X1_56/A MUX2X1_56/B MUX2X1_7/S gnd MUX2X1_57/A vdd MUX2X1
XMUX2X1_12 MUX2X1_11/Y MUX2X1_10/Y BUFX4_10/Y gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B MUX2X1_1/S gnd MUX2X1_34/Y vdd MUX2X1
XMUX2X1_78 MUX2X1_78/A MUX2X1_78/B BUFX4_8/Y gnd MUX2X1_78/Y vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XMUX2X1_45 MUX2X1_45/A MUX2X1_43/Y BUFX4_13/Y gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_89 MUX2X1_89/A NOR2X1_24/A MUX2X1_7/S gnd MUX2X1_89/Y vdd MUX2X1
XNAND2X1_93 MUX2X1_92/B NAND2X1_97/B gnd NAND2X1_93/Y vdd NAND2X1
XNAND2X1_71 AOI22X1_4/B NOR2X1_33/Y gnd NAND2X1_79/B vdd NAND2X1
XNAND2X1_82 MUX2X1_43/A NAND2X1_88/B gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_60 NAND2X1_60/A OAI21X1_52/B gnd NAND2X1_60/Y vdd NAND2X1
XFILL_21_2 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_25 BUFX4_16/Y NAND2X1_27/B NAND2X1_29/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_47 BUFX4_20/Y OAI21X1_52/B NAND2X1_54/Y gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_14 BUFX4_57/Y OAI21X1_7/B OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_69 BUFX4_40/Y NAND2X1_79/B NAND2X1_78/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_58 BUFX4_47/Y NAND2X1_65/B OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_36 BUFX4_27/Y OAI21X1_38/B OAI21X1_36/C gnd OAI21X1_36/Y vdd OAI21X1
XNAND2X1_267 MUX2X1_92/A NAND2X1_267/B gnd OAI21X1_218/C vdd NAND2X1
XOAI21X1_217 BUFX4_16/Y NAND2X1_267/B OAI21X1_217/C gnd DFFPOSX1_35/D vdd OAI21X1
XDFFPOSX1_153 MUX2X1_20/B CLKBUF1_32/A OAI21X1_79/Y gnd vdd DFFPOSX1
XNAND2X1_256 MUX2X1_58/B NAND2X1_256/B gnd OAI21X1_209/C vdd NAND2X1
XDFFPOSX1_131 MUX2X1_59/B CLKBUF1_22/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 NAND2X1_52/A CLKBUF1_4/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XOAI21X1_206 BUFX4_58/Y OAI21X1_201/B NAND2X1_251/Y gnd OAI21X1_206/Y vdd OAI21X1
XNAND2X1_234 MUX2X1_10/A OAI21X1_193/B gnd OAI21X1_191/C vdd NAND2X1
XDFFPOSX1_186 MUX2X1_47/B CLKBUF1_31/A OAI21X1_112/Y gnd vdd DFFPOSX1
XNAND2X1_201 AOI22X1_5/Y AOI22X1_6/Y gnd NAND2X1_201/Y vdd NAND2X1
XNAND2X1_245 MUX2X1_35/A OAI21X1_201/B gnd NAND2X1_245/Y vdd NAND2X1
XDFFPOSX1_142 NAND2X1_77/A CLKBUF1_43/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XOAI21X1_228 BUFX4_25/Y NAND2X1_279/B NAND2X1_279/Y gnd OAI21X1_228/Y vdd OAI21X1
XNAND2X1_212 r_w BUFX2_6/A gnd AOI21X1_30/A vdd NAND2X1
XNAND2X1_278 MUX2X1_104/A NAND2X1_279/B gnd OAI21X1_227/C vdd NAND2X1
XDFFPOSX1_164 MUX2X1_73/A CLKBUF1_20/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_175 MUX2X1_166/B CLKBUF1_7/A OAI21X1_101/Y gnd vdd DFFPOSX1
XDFFPOSX1_197 MUX2X1_119/A CLKBUF1_13/Y OAI21X1_123/Y gnd vdd DFFPOSX1
XNAND2X1_223 BUFX4_36/Y INVX1_2/Y gnd NOR2X1_30/B vdd NAND2X1
XFILL_22_2_1 gnd vdd FILL
XCLKBUF1_48 clk gnd CLKBUF1_23/A vdd CLKBUF1
XCLKBUF1_26 CLKBUF1_40/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_15 CLKBUF1_31/A gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_37 clk gnd CLKBUF1_8/A vdd CLKBUF1
XINVX1_1 address[4] gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XAND2X2_1 NOR2X1_2/Y AND2X2_4/B gnd NOR2X1_5/B vdd AND2X2
XNOR2X1_28 NOR2X1_28/A AND2X2_3/Y gnd NOR2X1_28/Y vdd NOR2X1
XNOR2X1_17 NOR2X1_17/A AND2X2_2/Y gnd NOR2X1_17/Y vdd NOR2X1
XMUX2X1_68 MUX2X1_68/A MUX2X1_68/B MUX2X1_2/S gnd MUX2X1_69/A vdd MUX2X1
XMUX2X1_24 MUX2X1_24/A MUX2X1_24/B BUFX4_6/Y gnd AOI22X1_4/D vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_57 MUX2X1_57/A MUX2X1_57/B BUFX4_9/Y gnd MUX2X1_57/Y vdd MUX2X1
XMUX2X1_13 MUX2X1_13/A MUX2X1_13/B BUFX4_37/Y gnd MUX2X1_15/B vdd MUX2X1
XMUX2X1_79 MUX2X1_79/A MUX2X1_79/B BUFX4_37/Y gnd MUX2X1_81/B vdd MUX2X1
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B MUX2X1_2/S gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_46 MUX2X1_46/A MUX2X1_46/B BUFX4_37/Y gnd MUX2X1_46/Y vdd MUX2X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_39 NOR2X1_39/A AND2X2_4/Y gnd NOR2X1_39/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XNAND2X1_72 MUX2X1_19/B NAND2X1_79/B gnd OAI21X1_63/C vdd NAND2X1
XNAND2X1_61 MUX2X1_173/B OAI21X1_52/B gnd OAI21X1_54/C vdd NAND2X1
XNAND2X1_83 MUX2X1_67/A NAND2X1_88/B gnd OAI21X1_73/C vdd NAND2X1
XNAND2X1_50 MUX2X1_124/A NAND2X1_50/B gnd NAND2X1_50/Y vdd NAND2X1
XNAND2X1_94 NAND2X1_94/A NAND2X1_97/B gnd NAND2X1_94/Y vdd NAND2X1
XFILL_21_3 gnd vdd FILL
XFILL_14_2 gnd vdd FILL
XOAI21X1_15 BUFX4_19/Y OAI21X1_18/B OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_26 BUFX4_45/Y NAND2X1_27/B NAND2X1_30/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_48 BUFX4_53/Y OAI21X1_52/B OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_37 BUFX4_41/Y OAI21X1_38/B OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_59 BUFX4_1/Y NAND2X1_65/B NAND2X1_67/Y gnd OAI21X1_59/Y vdd OAI21X1
XDFFPOSX1_187 MUX2X1_71/B CLKBUF1_2/A OAI21X1_113/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 MUX2X1_5/B CLKBUF1_23/A OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_176 MUX2X1_190/B CLKBUF1_2/A OAI21X1_102/Y gnd vdd DFFPOSX1
XNAND2X1_246 MUX2X1_59/A OAI21X1_201/B gnd NAND2X1_246/Y vdd NAND2X1
XOAI21X1_207 BUFX4_23/Y NAND2X1_256/B NAND2X1_254/Y gnd DFFPOSX1_25/D vdd OAI21X1
XOAI21X1_218 BUFX4_46/Y NAND2X1_267/B OAI21X1_218/C gnd OAI21X1_218/Y vdd OAI21X1
XNAND2X1_257 MUX2X1_82/B NAND2X1_256/B gnd NAND2X1_257/Y vdd NAND2X1
XNAND2X1_202 AOI22X1_7/Y AOI22X1_8/Y gnd NAND2X1_202/Y vdd NAND2X1
XDFFPOSX1_143 MUX2X1_163/B CLKBUF1_18/A OAI21X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 MUX2X1_44/B CLKBUF1_40/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XNAND2X1_235 MUX2X1_34/A OAI21X1_193/B gnd NAND2X1_235/Y vdd NAND2X1
XNAND2X1_268 MUX2X1_116/A NAND2X1_267/B gnd NAND2X1_268/Y vdd NAND2X1
XOAI21X1_229 BUFX4_40/Y NAND2X1_279/B NAND2X1_280/Y gnd DFFPOSX1_55/D vdd OAI21X1
XDFFPOSX1_132 MUX2X1_83/B CLKBUF1_20/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XNAND2X1_213 AOI22X1_21/Y AOI22X1_22/Y gnd NAND2X1_213/Y vdd NAND2X1
XDFFPOSX1_110 MUX2X1_125/A CLKBUF1_9/A OAI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_198 MUX2X1_143/A CLKBUF1_11/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XDFFPOSX1_165 MUX2X1_97/A CLKBUF1_16/Y OAI21X1_91/Y gnd vdd DFFPOSX1
XNAND2X1_224 AOI22X1_2/B AND2X2_2/B gnd OAI21X1_183/B vdd NAND2X1
XNAND2X1_279 MUX2X1_128/A NAND2X1_279/B gnd NAND2X1_279/Y vdd NAND2X1
XCLKBUF1_38 clk gnd CLKBUF1_38/Y vdd CLKBUF1
XCLKBUF1_27 CLKBUF1_31/A gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_16 CLKBUF1_6/A gnd CLKBUF1_16/Y vdd CLKBUF1
XINVX1_2 BUFX4_7/Y gnd INVX1_2/Y vdd INVX1
XAND2X2_2 INVX8_9/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 NOR2X1_18/A AND2X2_2/Y gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 address[2] NOR2X1_31/B gnd AOI22X1_2/B vdd NOR2X1
XMUX2X1_69 MUX2X1_69/A MUX2X1_67/Y BUFX4_13/Y gnd MUX2X1_69/Y vdd MUX2X1
XMUX2X1_58 MUX2X1_58/A MUX2X1_58/B MUX2X1_8/S gnd MUX2X1_60/B vdd MUX2X1
XMUX2X1_14 MUX2X1_14/A MUX2X1_14/B INVX1_3/A gnd MUX2X1_14/Y vdd MUX2X1
XNAND2X1_84 MUX2X1_91/A NAND2X1_88/B gnd OAI21X1_74/C vdd NAND2X1
XMUX2X1_47 MUX2X1_47/A MUX2X1_47/B INVX1_3/A gnd MUX2X1_48/A vdd MUX2X1
XMUX2X1_25 MUX2X1_25/A MUX2X1_25/B MUX2X1_8/S gnd MUX2X1_25/Y vdd MUX2X1
XMUX2X1_36 MUX2X1_35/Y MUX2X1_34/Y BUFX4_10/Y gnd MUX2X1_36/Y vdd MUX2X1
XNAND2X1_62 AOI22X1_2/C NOR2X1_1/Y gnd NAND2X1_65/B vdd NAND2X1
XNAND2X1_73 MUX2X1_43/B NAND2X1_79/B gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_95 MUX2X1_140/B NAND2X1_97/B gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_40 NAND2X1_40/A OAI21X1_38/B gnd OAI21X1_35/C vdd NAND2X1
XNAND2X1_51 MUX2X1_148/A NAND2X1_50/B gnd OAI21X1_45/C vdd NAND2X1
XFILL_20_3_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_14_3 gnd vdd FILL
XOAI21X1_38 BUFX4_56/Y OAI21X1_38/B OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_49 BUFX4_17/Y OAI21X1_52/B OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_16 BUFX4_52/Y OAI21X1_18/B NAND2X1_19/Y gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_27 BUFX4_3/Y NAND2X1_27/B NAND2X1_31/Y gnd OAI21X1_27/Y vdd OAI21X1
XDFFPOSX1_144 MUX2X1_187/B CLKBUF1_1/A OAI21X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_155 MUX2X1_68/B CLKBUF1_23/A OAI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 MUX2X1_29/B CLKBUF1_31/A OAI21X1_48/Y gnd vdd DFFPOSX1
XOAI21X1_208 BUFX4_54/Y NAND2X1_256/B NAND2X1_255/Y gnd OAI21X1_208/Y vdd OAI21X1
XOAI21X1_219 BUFX4_2/Y NAND2X1_267/B NAND2X1_268/Y gnd DFFPOSX1_37/D vdd OAI21X1
XDFFPOSX1_100 NOR2X1_14/A CLKBUF1_20/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 MUX2X1_149/A CLKBUF1_6/A OAI21X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 MUX2X1_107/B CLKBUF1_16/Y OAI21X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_177 MUX2X1_22/A CLKBUF1_32/Y OAI21X1_103/Y gnd vdd DFFPOSX1
XNAND2X1_225 MUX2X1_7/A OAI21X1_183/B gnd NAND2X1_225/Y vdd NAND2X1
XNAND2X1_203 r_w BUFX2_3/A gnd AOI21X1_27/A vdd NAND2X1
XNAND2X1_236 MUX2X1_58/A OAI21X1_193/B gnd NAND2X1_236/Y vdd NAND2X1
XDFFPOSX1_188 MUX2X1_95/B CLKBUF1_43/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XNAND2X1_247 MUX2X1_83/A OAI21X1_201/B gnd NAND2X1_247/Y vdd NAND2X1
XFILL_8_3_0 gnd vdd FILL
XNAND2X1_214 AOI22X1_23/Y AOI22X1_24/Y gnd OAI21X1_180/B vdd NAND2X1
XNAND2X1_258 MUX2X1_106/B NAND2X1_256/B gnd OAI21X1_211/C vdd NAND2X1
XNAND2X1_269 MUX2X1_140/A NAND2X1_267/B gnd OAI21X1_220/C vdd NAND2X1
XDFFPOSX1_199 MUX2X1_167/A CLKBUF1_7/Y OAI21X1_125/Y gnd vdd DFFPOSX1
XFILL_0_2_0 gnd vdd FILL
XDFFPOSX1_166 MUX2X1_121/A CLKBUF1_11/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XFILL_16_2_0 gnd vdd FILL
XCLKBUF1_28 CLKBUF1_32/A gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_17 CLKBUF1_4/A gnd CLKBUF1_17/Y vdd CLKBUF1
XCLKBUF1_39 clk gnd CLKBUF1_18/A vdd CLKBUF1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_22_0_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 INVX8_9/Y NOR2X1_1/Y gnd AND2X2_3/Y vdd AND2X2
XNOR2X1_19 OR2X2_1/B NOR2X1_19/B gnd AOI22X1_4/C vdd NOR2X1
XMUX2X1_59 MUX2X1_59/A MUX2X1_59/B BUFX4_35/Y gnd MUX2X1_59/Y vdd MUX2X1
XMUX2X1_15 MUX2X1_14/Y MUX2X1_15/B BUFX4_11/Y gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_37 MUX2X1_37/A MUX2X1_37/B MUX2X1_4/S gnd MUX2X1_39/B vdd MUX2X1
XMUX2X1_48 MUX2X1_48/A MUX2X1_46/Y BUFX4_6/Y gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_26 NOR2X1_4/A MUX2X1_26/B BUFX4_35/Y gnd MUX2X1_26/Y vdd MUX2X1
XFILL_20_3_1 gnd vdd FILL
XNAND2X1_74 MUX2X1_67/B NAND2X1_79/B gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_52 NAND2X1_52/A NAND2X1_50/B gnd OAI21X1_46/C vdd NAND2X1
XNAND2X1_63 MUX2X1_11/B NAND2X1_65/B gnd NAND2X1_63/Y vdd NAND2X1
XNAND2X1_30 MUX2X1_79/B NAND2X1_27/B gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_85 MUX2X1_115/A NAND2X1_88/B gnd OAI21X1_75/C vdd NAND2X1
XNAND2X1_41 MUX2X1_125/A OAI21X1_38/B gnd OAI21X1_36/C vdd NAND2X1
XNAND2X1_96 MUX2X1_164/B NAND2X1_97/B gnd NAND2X1_96/Y vdd NAND2X1
XFILL_11_3_1 gnd vdd FILL
XOAI21X1_39 BUFX4_23/Y NAND2X1_50/B NAND2X1_45/Y gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_17 BUFX4_18/Y OAI21X1_18/B NAND2X1_20/Y gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 BUFX4_28/Y NAND2X1_27/B OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_209 BUFX4_14/Y NAND2X1_256/B OAI21X1_209/C gnd DFFPOSX1_27/D vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_112 NAND2X1_43/A CLKBUF1_1/A OAI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 MUX2X1_19/A CLKBUF1_30/Y OAI21X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 MUX2X1_53/B CLKBUF1_2/A OAI21X1_49/Y gnd vdd DFFPOSX1
XNAND2X1_204 AOI22X1_9/Y AOI22X1_10/Y gnd NAND2X1_204/Y vdd NAND2X1
XNAND2X1_226 MUX2X1_31/A OAI21X1_183/B gnd NAND2X1_226/Y vdd NAND2X1
XDFFPOSX1_156 MUX2X1_92/B CLKBUF1_43/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XNAND2X1_237 MUX2X1_82/A OAI21X1_193/B gnd NAND2X1_237/Y vdd NAND2X1
XDFFPOSX1_178 MUX2X1_46/A CLKBUF1_25/Y OAI21X1_104/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 MUX2X1_131/B CLKBUF1_9/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 NOR2X1_15/A CLKBUF1_15/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XNAND2X1_259 MUX2X1_130/B NAND2X1_256/B gnd NAND2X1_259/Y vdd NAND2X1
XFILL_0_2_1 gnd vdd FILL
XDFFPOSX1_189 MUX2X1_119/B CLKBUF1_7/A OAI21X1_115/Y gnd vdd DFFPOSX1
XNAND2X1_215 r_w BUFX2_7/A gnd AOI21X1_31/A vdd NAND2X1
XDFFPOSX1_167 MUX2X1_145/A CLKBUF1_8/Y OAI21X1_93/Y gnd vdd DFFPOSX1
XNAND2X1_248 MUX2X1_107/A OAI21X1_201/B gnd NAND2X1_248/Y vdd NAND2X1
XFILL_16_2_1 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XCLKBUF1_29 CLKBUF1_32/A gnd CLKBUF1_29/Y vdd CLKBUF1
XBUFX4_50 INVX8_2/Y gnd BUFX4_50/Y vdd BUFX4
XCLKBUF1_18 CLKBUF1_18/A gnd CLKBUF1_18/Y vdd CLKBUF1
XINVX1_4 address[3] gnd INVX1_4/Y vdd INVX1
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XAND2X2_4 INVX8_9/Y AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XMUX2X1_16 MUX2X1_16/A MUX2X1_16/B BUFX4_39/Y gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B BUFX4_39/Y gnd MUX2X1_49/Y vdd MUX2X1
XMUX2X1_27 MUX2X1_26/Y MUX2X1_25/Y BUFX4_7/Y gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B MUX2X1_5/S gnd MUX2X1_38/Y vdd MUX2X1
XNAND2X1_97 MUX2X1_188/B NAND2X1_97/B gnd OAI21X1_86/C vdd NAND2X1
XNAND2X1_20 MUX2X1_49/B OAI21X1_18/B gnd NAND2X1_20/Y vdd NAND2X1
XNAND2X1_75 MUX2X1_91/B NAND2X1_79/B gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_86 NAND2X1_86/A NAND2X1_88/B gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_53 NOR2X1_1/Y AOI22X1_9/C gnd OAI21X1_52/B vdd NAND2X1
XNAND2X1_64 MUX2X1_35/B NAND2X1_65/B gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_31 MUX2X1_103/B NAND2X1_27/B gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_42 MUX2X1_149/A OAI21X1_38/B gnd OAI21X1_37/C vdd NAND2X1
XOAI21X1_18 BUFX4_49/Y OAI21X1_18/B OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 BUFX4_41/Y NAND2X1_27/B OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XDFFPOSX1_179 MUX2X1_70/A CLKBUF1_23/Y OAI21X1_105/Y gnd vdd DFFPOSX1
XNAND2X1_227 MUX2X1_55/A OAI21X1_183/B gnd OAI21X1_185/C vdd NAND2X1
XDFFPOSX1_113 MUX2X1_4/A CLKBUF1_30/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 MUX2X1_169/A CLKBUF1_2/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XNAND2X1_205 AOI22X1_11/Y AOI22X1_12/Y gnd OAI21X1_177/B vdd NAND2X1
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_146 MUX2X1_43/A CLKBUF1_26/Y OAI21X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 MUX2X1_77/B CLKBUF1_43/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 NAND2X1_94/A CLKBUF1_6/A OAI21X1_83/Y gnd vdd DFFPOSX1
XNAND2X1_238 MUX2X1_106/A OAI21X1_193/B gnd NAND2X1_238/Y vdd NAND2X1
XNAND2X1_249 MUX2X1_131/A OAI21X1_201/B gnd NAND2X1_249/Y vdd NAND2X1
XDFFPOSX1_135 MUX2X1_155/B CLKBUF1_5/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_102 NOR2X1_16/A CLKBUF1_9/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XNAND2X1_216 AOI22X1_25/Y AOI22X1_26/Y gnd OAI21X1_181/A vdd NAND2X1
XBUFX4_51 INVX8_2/Y gnd BUFX4_51/Y vdd BUFX4
XCLKBUF1_19 CLKBUF1_43/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_40 INVX8_7/Y gnd BUFX4_40/Y vdd BUFX4
.ends

