VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram32_sdram_2split
  CLASS BLOCK ;
  FOREIGN ram32_sdram_2split ;
  ORIGIN 2.600 3.000 ;
  SIZE 270.800 BY 246.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 240.200 265.400 240.800 ;
        RECT 0.600 235.900 1.000 240.200 ;
        RECT 2.200 235.900 2.600 240.200 ;
        RECT 3.800 235.900 4.200 240.200 ;
        RECT 5.400 235.900 5.800 240.200 ;
        RECT 7.000 235.900 7.400 240.200 ;
        RECT 7.800 235.900 8.200 240.200 ;
        RECT 9.400 235.900 9.800 240.200 ;
        RECT 11.000 235.900 11.400 240.200 ;
        RECT 12.600 235.900 13.000 240.200 ;
        RECT 14.200 235.900 14.600 240.200 ;
        RECT 15.000 235.900 15.400 240.200 ;
        RECT 16.600 235.900 17.000 240.200 ;
        RECT 18.200 235.900 18.600 240.200 ;
        RECT 19.800 235.900 20.200 240.200 ;
        RECT 21.400 235.900 21.800 240.200 ;
        RECT 22.200 235.900 22.600 240.200 ;
        RECT 23.800 235.900 24.200 240.200 ;
        RECT 25.400 235.900 25.800 240.200 ;
        RECT 27.000 235.900 27.400 240.200 ;
        RECT 28.600 235.900 29.000 240.200 ;
        RECT 29.400 235.900 29.800 240.200 ;
        RECT 31.000 235.900 31.400 240.200 ;
        RECT 32.600 235.900 33.000 240.200 ;
        RECT 34.200 235.900 34.600 240.200 ;
        RECT 35.800 235.900 36.200 240.200 ;
        RECT 36.600 235.900 37.000 240.200 ;
        RECT 38.200 235.900 38.600 240.200 ;
        RECT 39.800 235.900 40.200 240.200 ;
        RECT 41.400 235.900 41.800 240.200 ;
        RECT 43.000 235.900 43.400 240.200 ;
        RECT 44.600 236.000 45.000 240.200 ;
        RECT 47.400 237.900 47.800 240.200 ;
        RECT 49.000 237.900 49.400 240.200 ;
        RECT 51.800 235.900 52.200 240.200 ;
        RECT 55.000 235.900 55.400 240.200 ;
        RECT 56.600 235.900 57.000 240.200 ;
        RECT 58.200 235.900 58.600 240.200 ;
        RECT 59.800 235.900 60.200 240.200 ;
        RECT 61.400 235.900 61.800 240.200 ;
        RECT 62.200 235.900 62.600 240.200 ;
        RECT 64.300 237.900 64.700 240.200 ;
        RECT 65.400 237.900 65.800 240.200 ;
        RECT 67.000 237.900 67.400 240.200 ;
        RECT 68.600 236.000 69.000 240.200 ;
        RECT 71.400 237.900 71.800 240.200 ;
        RECT 73.000 237.900 73.400 240.200 ;
        RECT 75.800 235.900 76.200 240.200 ;
        RECT 78.200 236.000 78.600 240.200 ;
        RECT 81.000 237.900 81.400 240.200 ;
        RECT 82.600 237.900 83.000 240.200 ;
        RECT 85.400 235.900 85.800 240.200 ;
        RECT 87.000 237.900 87.400 240.200 ;
        RECT 89.200 235.900 89.600 240.200 ;
        RECT 91.800 236.100 92.200 240.200 ;
        RECT 94.200 236.000 94.600 240.200 ;
        RECT 97.000 237.900 97.400 240.200 ;
        RECT 98.600 237.900 99.000 240.200 ;
        RECT 101.400 235.900 101.800 240.200 ;
        RECT 103.300 237.900 103.700 240.200 ;
        RECT 105.400 235.900 105.800 240.200 ;
        RECT 107.800 237.900 108.200 240.200 ;
        RECT 109.400 237.900 109.800 240.200 ;
        RECT 110.200 235.900 110.600 240.200 ;
        RECT 112.300 237.900 112.700 240.200 ;
        RECT 114.200 236.000 114.600 240.200 ;
        RECT 117.000 237.900 117.400 240.200 ;
        RECT 118.600 237.900 119.000 240.200 ;
        RECT 121.400 235.900 121.800 240.200 ;
        RECT 123.000 235.900 123.400 240.200 ;
        RECT 125.100 237.900 125.500 240.200 ;
        RECT 126.200 237.900 126.600 240.200 ;
        RECT 127.800 237.900 128.200 240.200 ;
        RECT 129.400 236.000 129.800 240.200 ;
        RECT 132.200 237.900 132.600 240.200 ;
        RECT 133.800 237.900 134.200 240.200 ;
        RECT 136.600 235.900 137.000 240.200 ;
        RECT 138.200 237.900 138.600 240.200 ;
        RECT 139.800 237.900 140.200 240.200 ;
        RECT 140.900 237.900 141.300 240.200 ;
        RECT 143.000 235.900 143.400 240.200 ;
        RECT 144.600 236.500 145.000 240.200 ;
        RECT 147.000 235.900 147.400 240.200 ;
        RECT 150.200 235.900 150.600 240.200 ;
        RECT 153.000 237.900 153.400 240.200 ;
        RECT 154.600 237.900 155.000 240.200 ;
        RECT 157.400 236.000 157.800 240.200 ;
        RECT 160.600 237.900 161.000 240.200 ;
        RECT 162.200 237.900 162.600 240.200 ;
        RECT 163.300 237.900 163.700 240.200 ;
        RECT 165.400 235.900 165.800 240.200 ;
        RECT 167.000 236.000 167.400 240.200 ;
        RECT 169.800 237.900 170.200 240.200 ;
        RECT 171.400 237.900 171.800 240.200 ;
        RECT 174.200 235.900 174.600 240.200 ;
        RECT 176.600 236.100 177.000 240.200 ;
        RECT 179.200 235.900 179.600 240.200 ;
        RECT 180.600 237.900 181.000 240.200 ;
        RECT 182.200 237.900 182.600 240.200 ;
        RECT 183.300 237.900 183.700 240.200 ;
        RECT 185.400 235.900 185.800 240.200 ;
        RECT 187.000 236.000 187.400 240.200 ;
        RECT 189.800 237.900 190.200 240.200 ;
        RECT 191.400 237.900 191.800 240.200 ;
        RECT 194.200 235.900 194.600 240.200 ;
        RECT 196.600 235.900 197.000 240.200 ;
        RECT 199.400 237.900 199.800 240.200 ;
        RECT 201.000 237.900 201.400 240.200 ;
        RECT 203.800 236.000 204.200 240.200 ;
        RECT 207.000 235.900 207.400 240.200 ;
        RECT 208.600 235.900 209.000 240.200 ;
        RECT 210.200 235.900 210.600 240.200 ;
        RECT 211.800 235.900 212.200 240.200 ;
        RECT 213.400 235.900 213.800 240.200 ;
        RECT 214.200 235.900 214.600 240.200 ;
        RECT 215.800 235.900 216.200 240.200 ;
        RECT 217.400 235.900 217.800 240.200 ;
        RECT 219.000 235.900 219.400 240.200 ;
        RECT 220.600 235.900 221.000 240.200 ;
        RECT 221.400 235.900 221.800 240.200 ;
        RECT 223.500 237.900 223.900 240.200 ;
        RECT 224.600 237.900 225.000 240.200 ;
        RECT 226.200 237.900 226.600 240.200 ;
        RECT 227.000 235.900 227.400 240.200 ;
        RECT 228.600 235.900 229.000 240.200 ;
        RECT 230.200 235.900 230.600 240.200 ;
        RECT 231.800 235.900 232.200 240.200 ;
        RECT 233.400 235.900 233.800 240.200 ;
        RECT 235.000 236.000 235.400 240.200 ;
        RECT 237.800 237.900 238.200 240.200 ;
        RECT 239.400 237.900 239.800 240.200 ;
        RECT 242.200 235.900 242.600 240.200 ;
        RECT 244.600 235.900 245.000 240.200 ;
        RECT 247.400 237.900 247.800 240.200 ;
        RECT 249.000 237.900 249.400 240.200 ;
        RECT 251.800 236.000 252.200 240.200 ;
        RECT 253.400 237.900 253.800 240.200 ;
        RECT 255.000 237.900 255.400 240.200 ;
        RECT 255.800 235.900 256.200 240.200 ;
        RECT 257.400 235.900 257.800 240.200 ;
        RECT 259.000 235.900 259.400 240.200 ;
        RECT 260.600 235.900 261.000 240.200 ;
        RECT 262.200 235.900 262.600 240.200 ;
        RECT 0.600 220.800 1.000 225.100 ;
        RECT 2.200 220.800 2.600 225.100 ;
        RECT 3.800 220.800 4.200 225.100 ;
        RECT 5.400 220.800 5.800 225.100 ;
        RECT 7.000 220.800 7.400 225.100 ;
        RECT 8.600 220.800 9.000 225.000 ;
        RECT 11.400 220.800 11.800 223.100 ;
        RECT 13.000 220.800 13.400 223.100 ;
        RECT 15.800 220.800 16.200 225.100 ;
        RECT 18.200 220.800 18.600 224.500 ;
        RECT 22.200 220.800 22.600 225.100 ;
        RECT 23.800 220.800 24.200 225.000 ;
        RECT 26.600 220.800 27.000 223.100 ;
        RECT 28.200 220.800 28.600 223.100 ;
        RECT 31.000 220.800 31.400 225.100 ;
        RECT 33.400 220.800 33.800 224.900 ;
        RECT 36.000 220.800 36.400 225.100 ;
        RECT 38.200 220.800 38.600 223.100 ;
        RECT 39.800 220.800 40.200 224.900 ;
        RECT 42.400 220.800 42.800 225.100 ;
        RECT 43.800 220.800 44.200 225.100 ;
        RECT 45.400 220.800 45.800 224.500 ;
        RECT 47.800 220.800 48.200 223.100 ;
        RECT 48.600 220.800 49.000 225.100 ;
        RECT 50.200 220.800 50.600 225.100 ;
        RECT 51.800 220.800 52.200 225.100 ;
        RECT 55.000 220.800 55.400 225.000 ;
        RECT 57.800 220.800 58.200 223.100 ;
        RECT 59.400 220.800 59.800 223.100 ;
        RECT 62.200 220.800 62.600 225.100 ;
        RECT 63.800 220.800 64.200 225.100 ;
        RECT 65.900 220.800 66.300 223.100 ;
        RECT 67.000 220.800 67.400 223.100 ;
        RECT 68.600 220.800 69.000 223.100 ;
        RECT 70.000 220.800 70.400 225.100 ;
        RECT 72.600 220.800 73.000 224.900 ;
        RECT 75.000 220.800 75.400 225.100 ;
        RECT 77.800 220.800 78.200 223.100 ;
        RECT 79.400 220.800 79.800 223.100 ;
        RECT 82.200 220.800 82.600 225.000 ;
        RECT 83.800 220.800 84.200 225.100 ;
        RECT 87.800 220.800 88.200 224.500 ;
        RECT 89.400 220.800 89.800 225.100 ;
        RECT 91.000 220.800 91.400 225.100 ;
        RECT 92.600 220.800 93.000 225.100 ;
        RECT 94.200 220.800 94.600 225.100 ;
        RECT 95.800 220.800 96.200 225.100 ;
        RECT 97.400 220.800 97.800 225.000 ;
        RECT 100.200 220.800 100.600 223.100 ;
        RECT 101.800 220.800 102.200 223.100 ;
        RECT 104.600 220.800 105.000 225.100 ;
        RECT 108.600 220.800 109.000 224.900 ;
        RECT 111.200 220.800 111.600 225.100 ;
        RECT 112.600 220.800 113.000 223.100 ;
        RECT 114.200 220.800 114.600 223.100 ;
        RECT 115.800 220.800 116.200 224.500 ;
        RECT 117.400 220.800 117.800 225.100 ;
        RECT 118.200 220.800 118.600 225.100 ;
        RECT 119.800 220.800 120.200 225.100 ;
        RECT 121.400 220.800 121.800 225.100 ;
        RECT 122.800 220.800 123.200 225.100 ;
        RECT 125.400 220.800 125.800 224.900 ;
        RECT 127.800 220.800 128.200 224.900 ;
        RECT 130.400 220.800 130.800 225.100 ;
        RECT 132.600 220.800 133.000 224.900 ;
        RECT 135.200 220.800 135.600 225.100 ;
        RECT 136.600 220.800 137.000 223.100 ;
        RECT 138.200 220.800 138.600 223.100 ;
        RECT 139.300 220.800 139.700 223.100 ;
        RECT 141.400 220.800 141.800 225.100 ;
        RECT 143.000 220.800 143.400 225.100 ;
        RECT 145.800 220.800 146.200 223.100 ;
        RECT 147.400 220.800 147.800 223.100 ;
        RECT 150.200 220.800 150.600 225.000 ;
        RECT 152.600 220.800 153.000 224.900 ;
        RECT 155.200 220.800 155.600 225.100 ;
        RECT 158.800 220.800 159.200 225.100 ;
        RECT 161.400 220.800 161.800 224.900 ;
        RECT 163.800 220.800 164.200 225.100 ;
        RECT 166.600 220.800 167.000 223.100 ;
        RECT 168.200 220.800 168.600 223.100 ;
        RECT 171.000 220.800 171.400 225.000 ;
        RECT 172.600 220.800 173.000 225.100 ;
        RECT 176.600 220.800 177.000 224.500 ;
        RECT 178.800 220.800 179.200 225.100 ;
        RECT 181.400 220.800 181.800 224.900 ;
        RECT 183.000 220.800 183.400 223.100 ;
        RECT 184.600 220.800 185.000 223.100 ;
        RECT 186.200 220.800 186.600 225.100 ;
        RECT 189.000 220.800 189.400 223.100 ;
        RECT 190.600 220.800 191.000 223.100 ;
        RECT 193.400 220.800 193.800 225.000 ;
        RECT 195.000 220.800 195.400 225.100 ;
        RECT 199.000 220.800 199.400 224.500 ;
        RECT 201.400 220.800 201.800 225.100 ;
        RECT 204.200 220.800 204.600 223.100 ;
        RECT 205.800 220.800 206.200 223.100 ;
        RECT 208.600 220.800 209.000 225.000 ;
        RECT 211.800 220.800 212.200 225.100 ;
        RECT 215.800 220.800 216.200 224.500 ;
        RECT 218.200 220.800 218.600 225.000 ;
        RECT 221.000 220.800 221.400 223.100 ;
        RECT 222.600 220.800 223.000 223.100 ;
        RECT 225.400 220.800 225.800 225.100 ;
        RECT 227.000 220.800 227.400 225.100 ;
        RECT 228.600 220.800 229.000 225.100 ;
        RECT 230.200 220.800 230.600 225.100 ;
        RECT 231.600 220.800 232.000 225.100 ;
        RECT 234.200 220.800 234.600 224.900 ;
        RECT 235.800 220.800 236.200 225.100 ;
        RECT 237.900 220.800 238.300 223.100 ;
        RECT 239.000 220.800 239.400 223.100 ;
        RECT 240.600 220.800 241.000 223.100 ;
        RECT 241.400 220.800 241.800 223.100 ;
        RECT 243.000 220.800 243.400 223.100 ;
        RECT 244.100 220.800 244.500 223.100 ;
        RECT 246.200 220.800 246.600 225.100 ;
        RECT 247.000 220.800 247.400 225.100 ;
        RECT 248.600 220.800 249.000 225.100 ;
        RECT 250.200 220.800 250.600 225.100 ;
        RECT 251.800 220.800 252.200 225.100 ;
        RECT 253.400 220.800 253.800 225.100 ;
        RECT 254.200 220.800 254.600 223.100 ;
        RECT 255.800 220.800 256.200 223.100 ;
        RECT 256.600 220.800 257.000 225.100 ;
        RECT 258.200 220.800 258.600 225.100 ;
        RECT 259.800 220.800 260.200 225.100 ;
        RECT 261.400 220.800 261.800 225.100 ;
        RECT 263.000 220.800 263.400 225.100 ;
        RECT 0.200 220.200 265.400 220.800 ;
        RECT 1.400 215.900 1.800 220.200 ;
        RECT 4.200 217.900 4.600 220.200 ;
        RECT 5.800 217.900 6.200 220.200 ;
        RECT 8.600 216.000 9.000 220.200 ;
        RECT 10.200 215.900 10.600 220.200 ;
        RECT 14.200 216.500 14.600 220.200 ;
        RECT 16.600 215.900 17.000 220.200 ;
        RECT 19.400 217.900 19.800 220.200 ;
        RECT 21.000 217.900 21.400 220.200 ;
        RECT 23.800 216.000 24.200 220.200 ;
        RECT 26.200 215.900 26.600 220.200 ;
        RECT 29.000 217.900 29.400 220.200 ;
        RECT 30.600 217.900 31.000 220.200 ;
        RECT 33.400 216.000 33.800 220.200 ;
        RECT 35.000 217.900 35.400 220.200 ;
        RECT 36.600 217.900 37.000 220.200 ;
        RECT 37.700 217.900 38.100 220.200 ;
        RECT 39.800 215.900 40.200 220.200 ;
        RECT 40.600 215.900 41.000 220.200 ;
        RECT 42.200 216.500 42.600 220.200 ;
        RECT 44.600 216.100 45.000 220.200 ;
        RECT 47.200 215.900 47.600 220.200 ;
        RECT 49.400 216.000 49.800 220.200 ;
        RECT 52.200 217.900 52.600 220.200 ;
        RECT 53.800 217.900 54.200 220.200 ;
        RECT 56.600 215.900 57.000 220.200 ;
        RECT 59.800 217.900 60.200 220.200 ;
        RECT 61.400 217.900 61.800 220.200 ;
        RECT 62.500 217.900 62.900 220.200 ;
        RECT 64.600 215.900 65.000 220.200 ;
        RECT 65.400 215.900 65.800 220.200 ;
        RECT 67.500 217.900 67.900 220.200 ;
        RECT 68.600 217.900 69.000 220.200 ;
        RECT 70.200 217.900 70.600 220.200 ;
        RECT 71.800 215.900 72.200 220.200 ;
        RECT 74.600 217.900 75.000 220.200 ;
        RECT 76.200 217.900 76.600 220.200 ;
        RECT 79.000 216.000 79.400 220.200 ;
        RECT 81.400 215.900 81.800 220.200 ;
        RECT 84.200 217.900 84.600 220.200 ;
        RECT 85.800 217.900 86.200 220.200 ;
        RECT 88.600 216.000 89.000 220.200 ;
        RECT 91.000 216.000 91.400 220.200 ;
        RECT 93.800 217.900 94.200 220.200 ;
        RECT 95.400 217.900 95.800 220.200 ;
        RECT 98.200 215.900 98.600 220.200 ;
        RECT 101.400 216.500 101.800 220.200 ;
        RECT 105.400 215.900 105.800 220.200 ;
        RECT 108.200 217.900 108.600 220.200 ;
        RECT 109.800 217.900 110.200 220.200 ;
        RECT 112.600 216.000 113.000 220.200 ;
        RECT 114.200 217.900 114.600 220.200 ;
        RECT 115.800 215.900 116.200 220.200 ;
        RECT 119.800 216.500 120.200 220.200 ;
        RECT 122.200 215.900 122.600 220.200 ;
        RECT 125.000 217.900 125.400 220.200 ;
        RECT 126.600 217.900 127.000 220.200 ;
        RECT 129.400 216.000 129.800 220.200 ;
        RECT 131.600 215.900 132.000 220.200 ;
        RECT 134.200 216.100 134.600 220.200 ;
        RECT 135.800 215.900 136.200 220.200 ;
        RECT 137.400 216.500 137.800 220.200 ;
        RECT 139.800 216.500 140.200 220.200 ;
        RECT 141.400 215.900 141.800 220.200 ;
        RECT 142.200 215.900 142.600 220.200 ;
        RECT 143.800 215.900 144.200 220.200 ;
        RECT 145.400 215.900 145.800 220.200 ;
        RECT 147.000 215.900 147.400 220.200 ;
        RECT 148.600 215.900 149.000 220.200 ;
        RECT 150.200 215.900 150.600 220.200 ;
        RECT 153.000 217.900 153.400 220.200 ;
        RECT 154.600 217.900 155.000 220.200 ;
        RECT 157.400 216.000 157.800 220.200 ;
        RECT 160.600 215.900 161.000 220.200 ;
        RECT 162.200 215.900 162.600 220.200 ;
        RECT 163.800 215.900 164.200 220.200 ;
        RECT 165.400 215.900 165.800 220.200 ;
        RECT 167.000 215.900 167.400 220.200 ;
        RECT 168.600 215.900 169.000 220.200 ;
        RECT 171.400 217.900 171.800 220.200 ;
        RECT 173.000 217.900 173.400 220.200 ;
        RECT 175.800 216.000 176.200 220.200 ;
        RECT 177.400 217.900 177.800 220.200 ;
        RECT 179.000 217.900 179.400 220.200 ;
        RECT 180.100 217.900 180.500 220.200 ;
        RECT 182.200 215.900 182.600 220.200 ;
        RECT 183.300 217.900 183.700 220.200 ;
        RECT 185.400 215.900 185.800 220.200 ;
        RECT 186.200 215.900 186.600 220.200 ;
        RECT 187.800 215.900 188.200 220.200 ;
        RECT 189.400 215.900 189.800 220.200 ;
        RECT 191.000 215.900 191.400 220.200 ;
        RECT 192.600 215.900 193.000 220.200 ;
        RECT 193.400 215.900 193.800 220.200 ;
        RECT 195.500 217.900 195.900 220.200 ;
        RECT 196.600 217.900 197.000 220.200 ;
        RECT 198.200 217.900 198.600 220.200 ;
        RECT 199.800 215.900 200.200 220.200 ;
        RECT 202.600 217.900 203.000 220.200 ;
        RECT 204.200 217.900 204.600 220.200 ;
        RECT 207.000 216.000 207.400 220.200 ;
        RECT 211.000 216.000 211.400 220.200 ;
        RECT 213.800 217.900 214.200 220.200 ;
        RECT 215.400 217.900 215.800 220.200 ;
        RECT 218.200 215.900 218.600 220.200 ;
        RECT 220.600 216.500 221.000 220.200 ;
        RECT 222.200 215.900 222.600 220.200 ;
        RECT 223.000 215.900 223.400 220.200 ;
        RECT 224.600 216.500 225.000 220.200 ;
        RECT 227.000 215.900 227.400 220.200 ;
        RECT 229.800 217.900 230.200 220.200 ;
        RECT 231.400 217.900 231.800 220.200 ;
        RECT 234.200 216.000 234.600 220.200 ;
        RECT 236.600 215.900 237.000 220.200 ;
        RECT 239.400 217.900 239.800 220.200 ;
        RECT 241.000 217.900 241.400 220.200 ;
        RECT 243.800 216.000 244.200 220.200 ;
        RECT 246.200 216.000 246.600 220.200 ;
        RECT 249.000 217.900 249.400 220.200 ;
        RECT 250.600 217.900 251.000 220.200 ;
        RECT 253.400 215.900 253.800 220.200 ;
        RECT 255.800 216.000 256.200 220.200 ;
        RECT 258.600 217.900 259.000 220.200 ;
        RECT 260.200 217.900 260.600 220.200 ;
        RECT 263.000 215.900 263.400 220.200 ;
        RECT 1.400 200.800 1.800 205.000 ;
        RECT 4.200 200.800 4.600 203.100 ;
        RECT 5.800 200.800 6.200 203.100 ;
        RECT 8.600 200.800 9.000 205.100 ;
        RECT 10.500 200.800 10.900 203.100 ;
        RECT 12.600 200.800 13.000 205.100 ;
        RECT 13.400 200.800 13.800 203.100 ;
        RECT 15.000 200.800 15.400 203.100 ;
        RECT 16.600 200.800 17.000 203.100 ;
        RECT 18.000 200.800 18.400 205.100 ;
        RECT 20.600 200.800 21.000 204.900 ;
        RECT 22.800 200.800 23.200 205.100 ;
        RECT 25.400 200.800 25.800 204.900 ;
        RECT 27.600 200.800 28.000 205.100 ;
        RECT 30.200 200.800 30.600 204.900 ;
        RECT 32.600 200.800 33.000 205.000 ;
        RECT 35.400 200.800 35.800 203.100 ;
        RECT 37.000 200.800 37.400 203.100 ;
        RECT 39.800 200.800 40.200 205.100 ;
        RECT 42.200 200.800 42.600 204.900 ;
        RECT 44.800 200.800 45.200 205.100 ;
        RECT 47.000 200.800 47.400 203.100 ;
        RECT 48.600 200.800 49.000 204.900 ;
        RECT 51.200 200.800 51.600 205.100 ;
        RECT 55.000 200.800 55.400 205.000 ;
        RECT 57.800 200.800 58.200 203.100 ;
        RECT 59.400 200.800 59.800 203.100 ;
        RECT 62.200 200.800 62.600 205.100 ;
        RECT 63.800 200.800 64.200 203.100 ;
        RECT 66.000 200.800 66.400 205.100 ;
        RECT 68.600 200.800 69.000 204.900 ;
        RECT 70.800 200.800 71.200 205.100 ;
        RECT 73.400 200.800 73.800 204.900 ;
        RECT 75.000 200.800 75.400 205.100 ;
        RECT 79.000 200.800 79.400 204.500 ;
        RECT 81.400 200.800 81.800 205.000 ;
        RECT 84.200 200.800 84.600 203.100 ;
        RECT 85.800 200.800 86.200 203.100 ;
        RECT 88.600 200.800 89.000 205.100 ;
        RECT 90.500 200.800 90.900 203.100 ;
        RECT 92.600 200.800 93.000 205.100 ;
        RECT 94.200 200.800 94.600 204.900 ;
        RECT 96.800 200.800 97.200 205.100 ;
        RECT 98.200 200.800 98.600 205.100 ;
        RECT 101.200 200.800 101.600 205.100 ;
        RECT 103.800 200.800 104.200 204.900 ;
        RECT 107.800 200.800 108.200 204.900 ;
        RECT 110.400 200.800 110.800 205.100 ;
        RECT 112.600 200.800 113.000 204.900 ;
        RECT 115.200 200.800 115.600 205.100 ;
        RECT 116.600 200.800 117.000 205.100 ;
        RECT 118.700 200.800 119.100 203.100 ;
        RECT 119.800 200.800 120.200 203.100 ;
        RECT 121.400 200.800 121.800 203.100 ;
        RECT 123.000 200.800 123.400 205.100 ;
        RECT 125.800 200.800 126.200 203.100 ;
        RECT 127.400 200.800 127.800 203.100 ;
        RECT 130.200 200.800 130.600 205.000 ;
        RECT 132.600 200.800 133.000 205.000 ;
        RECT 135.400 200.800 135.800 203.100 ;
        RECT 137.000 200.800 137.400 203.100 ;
        RECT 139.800 200.800 140.200 205.100 ;
        RECT 141.400 200.800 141.800 205.100 ;
        RECT 143.500 200.800 143.900 203.100 ;
        RECT 144.600 200.800 145.000 203.100 ;
        RECT 146.200 200.800 146.600 203.100 ;
        RECT 147.800 200.800 148.200 204.900 ;
        RECT 150.400 200.800 150.800 205.100 ;
        RECT 152.100 200.800 152.500 203.100 ;
        RECT 154.200 200.800 154.600 205.100 ;
        RECT 155.300 200.800 155.700 203.100 ;
        RECT 157.400 200.800 157.800 205.100 ;
        RECT 159.800 200.800 160.200 205.100 ;
        RECT 161.900 200.800 162.300 203.100 ;
        RECT 163.000 200.800 163.400 203.100 ;
        RECT 164.600 200.800 165.000 203.100 ;
        RECT 166.200 200.800 166.600 205.100 ;
        RECT 169.000 200.800 169.400 203.100 ;
        RECT 170.600 200.800 171.000 203.100 ;
        RECT 173.400 200.800 173.800 205.000 ;
        RECT 175.800 200.800 176.200 205.100 ;
        RECT 178.600 200.800 179.000 203.100 ;
        RECT 180.200 200.800 180.600 203.100 ;
        RECT 183.000 200.800 183.400 205.000 ;
        RECT 185.400 200.800 185.800 205.100 ;
        RECT 188.200 200.800 188.600 203.100 ;
        RECT 189.800 200.800 190.200 203.100 ;
        RECT 192.600 200.800 193.000 205.000 ;
        RECT 194.200 200.800 194.600 205.100 ;
        RECT 196.300 200.800 196.700 203.100 ;
        RECT 197.700 200.800 198.100 203.100 ;
        RECT 199.800 200.800 200.200 205.100 ;
        RECT 201.400 200.800 201.800 204.900 ;
        RECT 204.000 200.800 204.400 205.100 ;
        RECT 205.400 200.800 205.800 203.100 ;
        RECT 209.200 200.800 209.600 205.100 ;
        RECT 211.800 200.800 212.200 204.900 ;
        RECT 213.400 200.800 213.800 205.100 ;
        RECT 217.400 200.800 217.800 204.500 ;
        RECT 219.800 200.800 220.200 204.900 ;
        RECT 222.400 200.800 222.800 205.100 ;
        RECT 223.800 200.800 224.200 205.100 ;
        RECT 225.900 200.800 226.300 203.100 ;
        RECT 227.300 200.800 227.700 203.100 ;
        RECT 229.400 200.800 229.800 205.100 ;
        RECT 231.000 200.800 231.400 205.100 ;
        RECT 233.800 200.800 234.200 203.100 ;
        RECT 235.400 200.800 235.800 203.100 ;
        RECT 238.200 200.800 238.600 205.000 ;
        RECT 240.600 200.800 241.000 204.900 ;
        RECT 243.200 200.800 243.600 205.100 ;
        RECT 245.400 200.800 245.800 203.100 ;
        RECT 247.000 200.800 247.400 205.100 ;
        RECT 249.800 200.800 250.200 203.100 ;
        RECT 251.400 200.800 251.800 203.100 ;
        RECT 254.200 200.800 254.600 205.000 ;
        RECT 255.800 200.800 256.200 205.100 ;
        RECT 257.400 200.800 257.800 205.100 ;
        RECT 259.000 200.800 259.400 205.100 ;
        RECT 260.600 200.800 261.000 205.100 ;
        RECT 262.200 200.800 262.600 205.100 ;
        RECT 0.200 200.200 265.400 200.800 ;
        RECT 0.600 195.900 1.000 200.200 ;
        RECT 2.200 195.900 2.600 200.200 ;
        RECT 3.800 195.900 4.200 200.200 ;
        RECT 5.400 195.900 5.800 200.200 ;
        RECT 7.000 195.900 7.400 200.200 ;
        RECT 8.600 196.000 9.000 200.200 ;
        RECT 11.400 197.900 11.800 200.200 ;
        RECT 13.000 197.900 13.400 200.200 ;
        RECT 15.800 195.900 16.200 200.200 ;
        RECT 17.400 195.900 17.800 200.200 ;
        RECT 21.400 196.500 21.800 200.200 ;
        RECT 23.000 197.900 23.400 200.200 ;
        RECT 24.600 197.900 25.000 200.200 ;
        RECT 25.700 197.900 26.100 200.200 ;
        RECT 27.800 195.900 28.200 200.200 ;
        RECT 29.400 195.900 29.800 200.200 ;
        RECT 32.200 197.900 32.600 200.200 ;
        RECT 33.800 197.900 34.200 200.200 ;
        RECT 36.600 196.000 37.000 200.200 ;
        RECT 39.000 196.000 39.400 200.200 ;
        RECT 41.800 197.900 42.200 200.200 ;
        RECT 43.400 197.900 43.800 200.200 ;
        RECT 46.200 195.900 46.600 200.200 ;
        RECT 48.100 197.900 48.500 200.200 ;
        RECT 50.200 195.900 50.600 200.200 ;
        RECT 53.400 195.900 53.800 200.200 ;
        RECT 56.200 197.900 56.600 200.200 ;
        RECT 57.800 197.900 58.200 200.200 ;
        RECT 60.600 196.000 61.000 200.200 ;
        RECT 63.000 196.500 63.400 200.200 ;
        RECT 65.400 195.900 65.800 200.200 ;
        RECT 68.100 197.900 68.500 200.200 ;
        RECT 70.200 195.900 70.600 200.200 ;
        RECT 71.800 195.900 72.200 200.200 ;
        RECT 74.600 197.900 75.000 200.200 ;
        RECT 76.200 197.900 76.600 200.200 ;
        RECT 79.000 196.000 79.400 200.200 ;
        RECT 81.400 196.100 81.800 200.200 ;
        RECT 84.000 195.900 84.400 200.200 ;
        RECT 85.400 197.900 85.800 200.200 ;
        RECT 87.000 197.900 87.400 200.200 ;
        RECT 88.600 196.100 89.000 200.200 ;
        RECT 91.200 195.900 91.600 200.200 ;
        RECT 93.400 197.900 93.800 200.200 ;
        RECT 95.000 195.900 95.400 200.200 ;
        RECT 97.800 197.900 98.200 200.200 ;
        RECT 99.400 197.900 99.800 200.200 ;
        RECT 102.200 196.000 102.600 200.200 ;
        RECT 103.800 195.900 104.200 200.200 ;
        RECT 105.400 196.500 105.800 200.200 ;
        RECT 109.400 195.900 109.800 200.200 ;
        RECT 112.200 197.900 112.600 200.200 ;
        RECT 113.800 197.900 114.200 200.200 ;
        RECT 116.600 196.000 117.000 200.200 ;
        RECT 118.200 197.900 118.600 200.200 ;
        RECT 119.800 197.900 120.200 200.200 ;
        RECT 120.900 197.900 121.300 200.200 ;
        RECT 123.000 195.900 123.400 200.200 ;
        RECT 123.800 195.900 124.200 200.200 ;
        RECT 125.400 196.500 125.800 200.200 ;
        RECT 127.000 197.900 127.400 200.200 ;
        RECT 128.600 197.900 129.000 200.200 ;
        RECT 129.700 197.900 130.100 200.200 ;
        RECT 131.800 195.900 132.200 200.200 ;
        RECT 133.400 196.000 133.800 200.200 ;
        RECT 136.200 197.900 136.600 200.200 ;
        RECT 137.800 197.900 138.200 200.200 ;
        RECT 140.600 195.900 141.000 200.200 ;
        RECT 143.000 196.100 143.400 200.200 ;
        RECT 145.600 195.900 146.000 200.200 ;
        RECT 147.600 195.900 148.000 200.200 ;
        RECT 150.200 196.100 150.600 200.200 ;
        RECT 152.600 196.500 153.000 200.200 ;
        RECT 154.200 195.900 154.600 200.200 ;
        RECT 156.300 197.900 156.700 200.200 ;
        RECT 159.000 197.900 159.400 200.200 ;
        RECT 160.600 197.900 161.000 200.200 ;
        RECT 162.200 195.900 162.600 200.200 ;
        RECT 165.000 197.900 165.400 200.200 ;
        RECT 166.600 197.900 167.000 200.200 ;
        RECT 169.400 196.000 169.800 200.200 ;
        RECT 171.000 195.900 171.400 200.200 ;
        RECT 172.600 196.500 173.000 200.200 ;
        RECT 174.200 197.900 174.600 200.200 ;
        RECT 176.400 195.900 176.800 200.200 ;
        RECT 179.000 196.100 179.400 200.200 ;
        RECT 180.600 197.900 181.000 200.200 ;
        RECT 182.200 197.900 182.600 200.200 ;
        RECT 183.300 197.900 183.700 200.200 ;
        RECT 185.400 195.900 185.800 200.200 ;
        RECT 187.000 196.100 187.400 200.200 ;
        RECT 189.600 195.900 190.000 200.200 ;
        RECT 191.800 197.900 192.200 200.200 ;
        RECT 193.400 195.900 193.800 200.200 ;
        RECT 196.200 197.900 196.600 200.200 ;
        RECT 197.800 197.900 198.200 200.200 ;
        RECT 200.600 196.000 201.000 200.200 ;
        RECT 203.000 195.900 203.400 200.200 ;
        RECT 205.800 197.900 206.200 200.200 ;
        RECT 207.400 197.900 207.800 200.200 ;
        RECT 210.200 196.000 210.600 200.200 ;
        RECT 213.400 197.900 213.800 200.200 ;
        RECT 215.000 197.900 215.400 200.200 ;
        RECT 216.100 197.900 216.500 200.200 ;
        RECT 218.200 195.900 218.600 200.200 ;
        RECT 219.800 196.100 220.200 200.200 ;
        RECT 222.400 195.900 222.800 200.200 ;
        RECT 224.600 196.500 225.000 200.200 ;
        RECT 226.200 195.900 226.600 200.200 ;
        RECT 227.000 195.900 227.400 200.200 ;
        RECT 229.100 197.900 229.500 200.200 ;
        RECT 230.200 197.900 230.600 200.200 ;
        RECT 231.800 197.900 232.200 200.200 ;
        RECT 233.400 195.900 233.800 200.200 ;
        RECT 236.200 197.900 236.600 200.200 ;
        RECT 237.800 197.900 238.200 200.200 ;
        RECT 240.600 196.000 241.000 200.200 ;
        RECT 243.000 196.100 243.400 200.200 ;
        RECT 245.600 195.900 246.000 200.200 ;
        RECT 247.000 195.900 247.400 200.200 ;
        RECT 249.100 197.900 249.500 200.200 ;
        RECT 251.000 197.900 251.400 200.200 ;
        RECT 252.600 195.900 253.000 200.200 ;
        RECT 255.400 197.900 255.800 200.200 ;
        RECT 257.000 197.900 257.400 200.200 ;
        RECT 259.800 196.000 260.200 200.200 ;
        RECT 261.400 195.900 261.800 200.200 ;
        RECT 263.500 197.900 263.900 200.200 ;
        RECT 1.400 180.800 1.800 185.000 ;
        RECT 4.200 180.800 4.600 183.100 ;
        RECT 5.800 180.800 6.200 183.100 ;
        RECT 8.600 180.800 9.000 185.100 ;
        RECT 10.200 180.800 10.600 183.100 ;
        RECT 12.400 180.800 12.800 185.100 ;
        RECT 15.000 180.800 15.400 184.900 ;
        RECT 17.400 180.800 17.800 185.000 ;
        RECT 20.200 180.800 20.600 183.100 ;
        RECT 21.800 180.800 22.200 183.100 ;
        RECT 24.600 180.800 25.000 185.100 ;
        RECT 27.000 180.800 27.400 184.900 ;
        RECT 29.600 180.800 30.000 185.100 ;
        RECT 31.800 180.800 32.200 183.100 ;
        RECT 33.200 180.800 33.600 185.100 ;
        RECT 35.800 180.800 36.200 184.900 ;
        RECT 38.000 180.800 38.400 185.100 ;
        RECT 40.600 180.800 41.000 184.900 ;
        RECT 43.000 180.800 43.400 184.900 ;
        RECT 45.600 180.800 46.000 185.100 ;
        RECT 47.000 180.800 47.400 183.100 ;
        RECT 48.600 180.800 49.000 183.100 ;
        RECT 50.200 180.800 50.600 184.900 ;
        RECT 52.800 180.800 53.200 185.100 ;
        RECT 56.600 180.800 57.000 184.900 ;
        RECT 59.200 180.800 59.600 185.100 ;
        RECT 61.400 180.800 61.800 184.900 ;
        RECT 64.000 180.800 64.400 185.100 ;
        RECT 65.400 180.800 65.800 183.100 ;
        RECT 67.000 180.800 67.400 183.100 ;
        RECT 68.600 180.800 69.000 184.900 ;
        RECT 71.200 180.800 71.600 185.100 ;
        RECT 73.400 180.800 73.800 183.100 ;
        RECT 75.000 180.800 75.400 185.000 ;
        RECT 77.800 180.800 78.200 183.100 ;
        RECT 79.400 180.800 79.800 183.100 ;
        RECT 82.200 180.800 82.600 185.100 ;
        RECT 84.600 180.800 85.000 184.900 ;
        RECT 87.200 180.800 87.600 185.100 ;
        RECT 88.600 180.800 89.000 183.100 ;
        RECT 90.800 180.800 91.200 185.100 ;
        RECT 93.400 180.800 93.800 184.900 ;
        RECT 95.600 180.800 96.000 185.100 ;
        RECT 98.200 180.800 98.600 184.900 ;
        RECT 100.400 180.800 100.800 185.100 ;
        RECT 103.000 180.800 103.400 184.900 ;
        RECT 107.000 180.800 107.400 185.100 ;
        RECT 109.800 180.800 110.200 183.100 ;
        RECT 111.400 180.800 111.800 183.100 ;
        RECT 114.200 180.800 114.600 185.000 ;
        RECT 115.800 180.800 116.200 183.100 ;
        RECT 117.400 180.800 117.800 183.100 ;
        RECT 118.500 180.800 118.900 183.100 ;
        RECT 120.600 180.800 121.000 185.100 ;
        RECT 121.400 180.800 121.800 185.100 ;
        RECT 123.000 180.800 123.400 185.100 ;
        RECT 124.600 180.800 125.000 185.100 ;
        RECT 126.200 180.800 126.600 185.100 ;
        RECT 127.800 180.800 128.200 185.100 ;
        RECT 129.400 180.800 129.800 185.000 ;
        RECT 132.200 180.800 132.600 183.100 ;
        RECT 133.800 180.800 134.200 183.100 ;
        RECT 136.600 180.800 137.000 185.100 ;
        RECT 138.200 180.800 138.600 185.100 ;
        RECT 140.300 180.800 140.700 183.100 ;
        RECT 141.400 180.800 141.800 183.100 ;
        RECT 143.000 180.800 143.400 183.100 ;
        RECT 144.600 180.800 145.000 185.000 ;
        RECT 147.400 180.800 147.800 183.100 ;
        RECT 149.000 180.800 149.400 183.100 ;
        RECT 151.800 180.800 152.200 185.100 ;
        RECT 155.800 180.800 156.200 185.000 ;
        RECT 158.600 180.800 159.000 183.100 ;
        RECT 160.200 180.800 160.600 183.100 ;
        RECT 163.000 180.800 163.400 185.100 ;
        RECT 164.600 180.800 165.000 183.100 ;
        RECT 166.800 180.800 167.200 185.100 ;
        RECT 169.400 180.800 169.800 184.900 ;
        RECT 171.600 180.800 172.000 185.100 ;
        RECT 174.200 180.800 174.600 184.900 ;
        RECT 176.600 180.800 177.000 184.900 ;
        RECT 179.200 180.800 179.600 185.100 ;
        RECT 181.400 180.800 181.800 184.900 ;
        RECT 184.000 180.800 184.400 185.100 ;
        RECT 186.200 180.800 186.600 184.500 ;
        RECT 187.800 180.800 188.200 185.100 ;
        RECT 189.400 180.800 189.800 184.900 ;
        RECT 192.000 180.800 192.400 185.100 ;
        RECT 194.000 180.800 194.400 185.100 ;
        RECT 196.600 180.800 197.000 184.900 ;
        RECT 198.800 180.800 199.200 185.100 ;
        RECT 201.400 180.800 201.800 184.900 ;
        RECT 203.800 180.800 204.200 184.900 ;
        RECT 206.400 180.800 206.800 185.100 ;
        RECT 210.200 180.800 210.600 184.900 ;
        RECT 212.800 180.800 213.200 185.100 ;
        RECT 215.000 180.800 215.400 184.900 ;
        RECT 217.600 180.800 218.000 185.100 ;
        RECT 219.800 180.800 220.200 185.000 ;
        RECT 222.600 180.800 223.000 183.100 ;
        RECT 224.200 180.800 224.600 183.100 ;
        RECT 227.000 180.800 227.400 185.100 ;
        RECT 229.200 180.800 229.600 185.100 ;
        RECT 231.800 180.800 232.200 184.900 ;
        RECT 234.000 180.800 234.400 185.100 ;
        RECT 236.600 180.800 237.000 184.900 ;
        RECT 238.200 180.800 238.600 183.100 ;
        RECT 239.800 180.800 240.200 183.100 ;
        RECT 240.900 180.800 241.300 183.100 ;
        RECT 243.000 180.800 243.400 185.100 ;
        RECT 244.600 180.800 245.000 185.100 ;
        RECT 247.400 180.800 247.800 183.100 ;
        RECT 249.000 180.800 249.400 183.100 ;
        RECT 251.800 180.800 252.200 185.000 ;
        RECT 253.400 180.800 253.800 185.100 ;
        RECT 255.000 180.800 255.400 185.100 ;
        RECT 256.600 180.800 257.000 185.100 ;
        RECT 258.200 180.800 258.600 185.100 ;
        RECT 259.800 180.800 260.200 185.100 ;
        RECT 260.600 180.800 261.000 183.100 ;
        RECT 262.200 180.800 262.600 183.100 ;
        RECT 0.200 180.200 265.400 180.800 ;
        RECT 1.400 175.900 1.800 180.200 ;
        RECT 4.200 177.900 4.600 180.200 ;
        RECT 5.800 177.900 6.200 180.200 ;
        RECT 8.600 176.000 9.000 180.200 ;
        RECT 10.800 175.900 11.200 180.200 ;
        RECT 13.400 176.100 13.800 180.200 ;
        RECT 15.800 176.100 16.200 180.200 ;
        RECT 18.400 175.900 18.800 180.200 ;
        RECT 20.400 175.900 20.800 180.200 ;
        RECT 23.000 176.100 23.400 180.200 ;
        RECT 25.200 175.900 25.600 180.200 ;
        RECT 27.800 176.100 28.200 180.200 ;
        RECT 30.000 175.900 30.400 180.200 ;
        RECT 32.600 176.100 33.000 180.200 ;
        RECT 34.200 177.900 34.600 180.200 ;
        RECT 35.800 177.900 36.200 180.200 ;
        RECT 37.400 176.500 37.800 180.200 ;
        RECT 41.400 176.500 41.800 180.200 ;
        RECT 44.600 175.900 45.000 180.200 ;
        RECT 46.200 176.500 46.600 180.200 ;
        RECT 49.400 175.900 49.800 180.200 ;
        RECT 50.800 175.900 51.200 180.200 ;
        RECT 53.400 176.100 53.800 180.200 ;
        RECT 57.400 176.100 57.800 180.200 ;
        RECT 60.000 175.900 60.400 180.200 ;
        RECT 62.000 175.900 62.400 180.200 ;
        RECT 64.600 176.100 65.000 180.200 ;
        RECT 66.200 177.900 66.600 180.200 ;
        RECT 67.800 177.900 68.200 180.200 ;
        RECT 68.900 177.900 69.300 180.200 ;
        RECT 71.000 175.900 71.400 180.200 ;
        RECT 72.600 175.900 73.000 180.200 ;
        RECT 75.400 177.900 75.800 180.200 ;
        RECT 77.000 177.900 77.400 180.200 ;
        RECT 79.800 176.000 80.200 180.200 ;
        RECT 83.800 176.500 84.200 180.200 ;
        RECT 86.200 175.900 86.600 180.200 ;
        RECT 89.000 177.900 89.400 180.200 ;
        RECT 90.600 177.900 91.000 180.200 ;
        RECT 93.400 176.000 93.800 180.200 ;
        RECT 97.400 176.500 97.800 180.200 ;
        RECT 99.600 175.900 100.000 180.200 ;
        RECT 102.200 176.100 102.600 180.200 ;
        RECT 103.800 177.900 104.200 180.200 ;
        RECT 105.400 177.900 105.800 180.200 ;
        RECT 110.200 176.500 110.600 180.200 ;
        RECT 111.800 177.900 112.200 180.200 ;
        RECT 113.400 177.900 113.800 180.200 ;
        RECT 116.600 176.500 117.000 180.200 ;
        RECT 119.000 175.900 119.400 180.200 ;
        RECT 121.800 177.900 122.200 180.200 ;
        RECT 123.400 177.900 123.800 180.200 ;
        RECT 126.200 176.000 126.600 180.200 ;
        RECT 127.800 175.900 128.200 180.200 ;
        RECT 131.800 176.500 132.200 180.200 ;
        RECT 134.200 176.000 134.600 180.200 ;
        RECT 137.000 177.900 137.400 180.200 ;
        RECT 138.600 177.900 139.000 180.200 ;
        RECT 141.400 175.900 141.800 180.200 ;
        RECT 143.000 177.900 143.400 180.200 ;
        RECT 145.200 175.900 145.600 180.200 ;
        RECT 147.800 176.100 148.200 180.200 ;
        RECT 150.200 176.500 150.600 180.200 ;
        RECT 152.600 177.900 153.000 180.200 ;
        RECT 154.200 177.900 154.600 180.200 ;
        RECT 157.400 176.000 157.800 180.200 ;
        RECT 160.200 177.900 160.600 180.200 ;
        RECT 161.800 177.900 162.200 180.200 ;
        RECT 164.600 175.900 165.000 180.200 ;
        RECT 166.200 177.900 166.600 180.200 ;
        RECT 168.400 175.900 168.800 180.200 ;
        RECT 171.000 176.100 171.400 180.200 ;
        RECT 173.400 176.000 173.800 180.200 ;
        RECT 176.200 177.900 176.600 180.200 ;
        RECT 177.800 177.900 178.200 180.200 ;
        RECT 180.600 175.900 181.000 180.200 ;
        RECT 183.000 175.900 183.400 180.200 ;
        RECT 185.800 177.900 186.200 180.200 ;
        RECT 187.400 177.900 187.800 180.200 ;
        RECT 190.200 176.000 190.600 180.200 ;
        RECT 192.600 176.100 193.000 180.200 ;
        RECT 195.200 175.900 195.600 180.200 ;
        RECT 197.400 176.000 197.800 180.200 ;
        RECT 200.200 177.900 200.600 180.200 ;
        RECT 201.800 177.900 202.200 180.200 ;
        RECT 204.600 175.900 205.000 180.200 ;
        RECT 207.000 177.900 207.400 180.200 ;
        RECT 209.400 177.900 209.800 180.200 ;
        RECT 211.000 177.900 211.400 180.200 ;
        RECT 212.600 176.500 213.000 180.200 ;
        RECT 218.200 176.500 218.600 180.200 ;
        RECT 220.400 175.900 220.800 180.200 ;
        RECT 223.000 176.100 223.400 180.200 ;
        RECT 225.400 176.100 225.800 180.200 ;
        RECT 228.000 175.900 228.400 180.200 ;
        RECT 229.700 177.900 230.100 180.200 ;
        RECT 231.800 175.900 232.200 180.200 ;
        RECT 232.900 177.900 233.300 180.200 ;
        RECT 235.000 175.900 235.400 180.200 ;
        RECT 235.800 177.900 236.200 180.200 ;
        RECT 237.400 177.900 237.800 180.200 ;
        RECT 239.000 175.900 239.400 180.200 ;
        RECT 241.800 177.900 242.200 180.200 ;
        RECT 243.400 177.900 243.800 180.200 ;
        RECT 246.200 176.000 246.600 180.200 ;
        RECT 248.100 177.900 248.500 180.200 ;
        RECT 250.200 175.900 250.600 180.200 ;
        RECT 251.800 175.900 252.200 180.200 ;
        RECT 254.600 177.900 255.000 180.200 ;
        RECT 256.200 177.900 256.600 180.200 ;
        RECT 259.000 176.000 259.400 180.200 ;
        RECT 260.600 177.900 261.000 180.200 ;
        RECT 262.200 177.900 262.600 180.200 ;
        RECT 1.400 160.800 1.800 165.000 ;
        RECT 4.200 160.800 4.600 163.100 ;
        RECT 5.800 160.800 6.200 163.100 ;
        RECT 8.600 160.800 9.000 165.100 ;
        RECT 10.200 160.800 10.600 163.100 ;
        RECT 11.800 160.800 12.200 163.100 ;
        RECT 12.900 160.800 13.300 163.100 ;
        RECT 15.000 160.800 15.400 165.100 ;
        RECT 16.600 160.800 17.000 165.000 ;
        RECT 19.400 160.800 19.800 163.100 ;
        RECT 21.000 160.800 21.400 163.100 ;
        RECT 23.800 160.800 24.200 165.100 ;
        RECT 25.400 160.800 25.800 163.100 ;
        RECT 27.600 160.800 28.000 165.100 ;
        RECT 30.200 160.800 30.600 164.900 ;
        RECT 31.800 160.800 32.200 163.100 ;
        RECT 33.400 160.800 33.800 163.100 ;
        RECT 34.500 160.800 34.900 163.100 ;
        RECT 36.600 160.800 37.000 165.100 ;
        RECT 37.700 160.800 38.100 163.100 ;
        RECT 39.800 160.800 40.200 165.100 ;
        RECT 41.400 160.800 41.800 165.100 ;
        RECT 44.200 160.800 44.600 163.100 ;
        RECT 45.800 160.800 46.200 163.100 ;
        RECT 48.600 160.800 49.000 165.000 ;
        RECT 51.800 160.800 52.200 164.500 ;
        RECT 55.800 160.800 56.200 165.100 ;
        RECT 58.600 160.800 59.000 163.100 ;
        RECT 60.200 160.800 60.600 163.100 ;
        RECT 63.000 160.800 63.400 165.000 ;
        RECT 64.600 160.800 65.000 163.100 ;
        RECT 66.200 160.800 66.600 163.100 ;
        RECT 67.300 160.800 67.700 163.100 ;
        RECT 69.400 160.800 69.800 165.100 ;
        RECT 71.000 160.800 71.400 165.100 ;
        RECT 73.800 160.800 74.200 163.100 ;
        RECT 75.400 160.800 75.800 163.100 ;
        RECT 78.200 160.800 78.600 165.000 ;
        RECT 79.800 160.800 80.200 165.100 ;
        RECT 81.400 160.800 81.800 165.100 ;
        RECT 83.000 160.800 83.400 165.100 ;
        RECT 84.600 160.800 85.000 165.100 ;
        RECT 86.200 160.800 86.600 165.100 ;
        RECT 87.600 160.800 88.000 165.100 ;
        RECT 90.200 160.800 90.600 164.900 ;
        RECT 92.400 160.800 92.800 165.100 ;
        RECT 95.000 160.800 95.400 164.900 ;
        RECT 96.600 160.800 97.000 163.100 ;
        RECT 98.200 160.800 98.600 163.100 ;
        RECT 99.800 160.800 100.200 164.900 ;
        RECT 102.400 160.800 102.800 165.100 ;
        RECT 106.200 160.800 106.600 165.000 ;
        RECT 109.000 160.800 109.400 163.100 ;
        RECT 110.600 160.800 111.000 163.100 ;
        RECT 113.400 160.800 113.800 165.100 ;
        RECT 115.000 160.800 115.400 163.100 ;
        RECT 117.200 160.800 117.600 165.100 ;
        RECT 119.800 160.800 120.200 164.900 ;
        RECT 122.200 160.800 122.600 164.500 ;
        RECT 123.800 160.800 124.200 165.100 ;
        RECT 125.400 160.800 125.800 164.900 ;
        RECT 128.000 160.800 128.400 165.100 ;
        RECT 130.200 160.800 130.600 164.900 ;
        RECT 132.800 160.800 133.200 165.100 ;
        RECT 134.800 160.800 135.200 165.100 ;
        RECT 137.400 160.800 137.800 164.900 ;
        RECT 141.400 160.800 141.800 164.500 ;
        RECT 143.000 160.800 143.400 163.100 ;
        RECT 144.600 160.800 145.000 163.100 ;
        RECT 145.400 160.800 145.800 165.100 ;
        RECT 147.500 160.800 147.900 163.100 ;
        RECT 149.400 160.800 149.800 164.500 ;
        RECT 153.200 160.800 153.600 165.100 ;
        RECT 155.800 160.800 156.200 164.900 ;
        RECT 159.600 160.800 160.000 165.100 ;
        RECT 162.200 160.800 162.600 164.900 ;
        RECT 164.600 160.800 165.000 164.900 ;
        RECT 167.200 160.800 167.600 165.100 ;
        RECT 168.600 160.800 169.000 165.100 ;
        RECT 170.700 160.800 171.100 163.100 ;
        RECT 172.600 160.800 173.000 164.900 ;
        RECT 175.200 160.800 175.600 165.100 ;
        RECT 177.400 160.800 177.800 164.900 ;
        RECT 180.000 160.800 180.400 165.100 ;
        RECT 182.200 160.800 182.600 164.500 ;
        RECT 184.600 160.800 185.000 165.100 ;
        RECT 187.800 160.800 188.200 164.500 ;
        RECT 191.000 160.800 191.400 163.100 ;
        RECT 192.600 160.800 193.000 163.100 ;
        RECT 193.400 160.800 193.800 165.100 ;
        RECT 195.500 160.800 195.900 163.100 ;
        RECT 197.400 160.800 197.800 164.500 ;
        RECT 200.900 160.800 201.300 163.100 ;
        RECT 203.000 160.800 203.400 165.100 ;
        RECT 206.200 160.800 206.600 165.100 ;
        RECT 209.000 160.800 209.400 163.100 ;
        RECT 210.600 160.800 211.000 163.100 ;
        RECT 213.400 160.800 213.800 165.000 ;
        RECT 215.000 160.800 215.400 163.100 ;
        RECT 217.200 160.800 217.600 165.100 ;
        RECT 219.800 160.800 220.200 164.900 ;
        RECT 222.000 160.800 222.400 165.100 ;
        RECT 224.600 160.800 225.000 164.900 ;
        RECT 226.800 160.800 227.200 165.100 ;
        RECT 229.400 160.800 229.800 164.900 ;
        RECT 231.600 160.800 232.000 165.100 ;
        RECT 234.200 160.800 234.600 164.900 ;
        RECT 236.100 160.800 236.500 163.100 ;
        RECT 238.200 160.800 238.600 165.100 ;
        RECT 240.600 160.800 241.000 165.100 ;
        RECT 243.000 160.800 243.400 164.500 ;
        RECT 244.600 160.800 245.000 163.100 ;
        RECT 246.200 160.800 246.600 163.100 ;
        RECT 247.800 160.800 248.200 165.100 ;
        RECT 250.600 160.800 251.000 163.100 ;
        RECT 252.200 160.800 252.600 163.100 ;
        RECT 255.000 160.800 255.400 165.000 ;
        RECT 258.200 160.800 258.600 164.500 ;
        RECT 260.600 160.800 261.000 164.500 ;
        RECT 263.000 160.800 263.400 164.500 ;
        RECT 0.200 160.200 265.400 160.800 ;
        RECT 1.400 156.000 1.800 160.200 ;
        RECT 4.200 157.900 4.600 160.200 ;
        RECT 5.800 157.900 6.200 160.200 ;
        RECT 8.600 155.900 9.000 160.200 ;
        RECT 10.200 157.900 10.600 160.200 ;
        RECT 11.800 157.900 12.200 160.200 ;
        RECT 12.600 155.900 13.000 160.200 ;
        RECT 14.200 155.900 14.600 160.200 ;
        RECT 15.800 155.900 16.200 160.200 ;
        RECT 17.400 155.900 17.800 160.200 ;
        RECT 19.000 155.900 19.400 160.200 ;
        RECT 20.600 156.000 21.000 160.200 ;
        RECT 23.400 157.900 23.800 160.200 ;
        RECT 25.000 157.900 25.400 160.200 ;
        RECT 27.800 155.900 28.200 160.200 ;
        RECT 30.200 156.000 30.600 160.200 ;
        RECT 33.000 157.900 33.400 160.200 ;
        RECT 34.600 157.900 35.000 160.200 ;
        RECT 37.400 155.900 37.800 160.200 ;
        RECT 39.000 155.900 39.400 160.200 ;
        RECT 43.000 156.500 43.400 160.200 ;
        RECT 44.600 155.900 45.000 160.200 ;
        RECT 46.200 156.500 46.600 160.200 ;
        RECT 48.600 156.100 49.000 160.200 ;
        RECT 51.200 155.900 51.600 160.200 ;
        RECT 53.400 157.900 53.800 160.200 ;
        RECT 56.600 156.000 57.000 160.200 ;
        RECT 59.400 157.900 59.800 160.200 ;
        RECT 61.000 157.900 61.400 160.200 ;
        RECT 63.800 155.900 64.200 160.200 ;
        RECT 66.200 156.000 66.600 160.200 ;
        RECT 69.000 157.900 69.400 160.200 ;
        RECT 70.600 157.900 71.000 160.200 ;
        RECT 73.400 155.900 73.800 160.200 ;
        RECT 75.600 155.900 76.000 160.200 ;
        RECT 78.200 156.100 78.600 160.200 ;
        RECT 79.800 157.900 80.200 160.200 ;
        RECT 81.400 157.900 81.800 160.200 ;
        RECT 82.500 157.900 82.900 160.200 ;
        RECT 84.600 155.900 85.000 160.200 ;
        RECT 86.000 155.900 86.400 160.200 ;
        RECT 88.600 156.100 89.000 160.200 ;
        RECT 91.000 156.000 91.400 160.200 ;
        RECT 93.800 157.900 94.200 160.200 ;
        RECT 95.400 157.900 95.800 160.200 ;
        RECT 98.200 155.900 98.600 160.200 ;
        RECT 100.600 156.100 101.000 160.200 ;
        RECT 103.200 155.900 103.600 160.200 ;
        RECT 104.600 157.900 105.000 160.200 ;
        RECT 106.200 157.900 106.600 160.200 ;
        RECT 108.900 157.900 109.300 160.200 ;
        RECT 111.000 155.900 111.400 160.200 ;
        RECT 111.800 157.900 112.200 160.200 ;
        RECT 113.400 157.900 113.800 160.200 ;
        RECT 114.200 155.900 114.600 160.200 ;
        RECT 117.400 156.000 117.800 160.200 ;
        RECT 120.200 157.900 120.600 160.200 ;
        RECT 121.800 157.900 122.200 160.200 ;
        RECT 124.600 155.900 125.000 160.200 ;
        RECT 126.200 155.900 126.600 160.200 ;
        RECT 128.300 157.900 128.700 160.200 ;
        RECT 129.700 157.900 130.100 160.200 ;
        RECT 131.800 155.900 132.200 160.200 ;
        RECT 133.400 156.000 133.800 160.200 ;
        RECT 136.200 157.900 136.600 160.200 ;
        RECT 137.800 157.900 138.200 160.200 ;
        RECT 140.600 155.900 141.000 160.200 ;
        RECT 142.200 157.900 142.600 160.200 ;
        RECT 143.800 157.900 144.200 160.200 ;
        RECT 144.600 157.900 145.000 160.200 ;
        RECT 146.200 157.900 146.600 160.200 ;
        RECT 147.300 157.900 147.700 160.200 ;
        RECT 149.400 155.900 149.800 160.200 ;
        RECT 150.200 157.900 150.600 160.200 ;
        RECT 151.800 157.900 152.200 160.200 ;
        RECT 155.000 155.900 155.400 160.200 ;
        RECT 157.800 157.900 158.200 160.200 ;
        RECT 159.400 157.900 159.800 160.200 ;
        RECT 162.200 156.000 162.600 160.200 ;
        RECT 163.800 157.900 164.200 160.200 ;
        RECT 165.400 157.900 165.800 160.200 ;
        RECT 166.500 157.900 166.900 160.200 ;
        RECT 168.600 155.900 169.000 160.200 ;
        RECT 169.400 155.900 169.800 160.200 ;
        RECT 172.600 156.500 173.000 160.200 ;
        RECT 175.000 155.900 175.400 160.200 ;
        RECT 177.100 157.900 177.500 160.200 ;
        RECT 178.800 155.900 179.200 160.200 ;
        RECT 181.400 156.100 181.800 160.200 ;
        RECT 183.800 156.000 184.200 160.200 ;
        RECT 186.600 157.900 187.000 160.200 ;
        RECT 188.200 157.900 188.600 160.200 ;
        RECT 191.000 155.900 191.400 160.200 ;
        RECT 192.600 155.900 193.000 160.200 ;
        RECT 194.700 157.900 195.100 160.200 ;
        RECT 195.800 155.900 196.200 160.200 ;
        RECT 197.900 157.900 198.300 160.200 ;
        RECT 199.000 157.900 199.400 160.200 ;
        RECT 200.600 157.900 201.000 160.200 ;
        RECT 201.700 157.900 202.100 160.200 ;
        RECT 203.800 155.900 204.200 160.200 ;
        RECT 205.200 155.900 205.600 160.200 ;
        RECT 207.800 156.100 208.200 160.200 ;
        RECT 213.400 156.500 213.800 160.200 ;
        RECT 215.800 156.100 216.200 160.200 ;
        RECT 218.400 155.900 218.800 160.200 ;
        RECT 220.400 155.900 220.800 160.200 ;
        RECT 223.000 156.100 223.400 160.200 ;
        RECT 225.400 156.100 225.800 160.200 ;
        RECT 228.000 155.900 228.400 160.200 ;
        RECT 231.000 156.500 231.400 160.200 ;
        RECT 233.400 156.000 233.800 160.200 ;
        RECT 236.200 157.900 236.600 160.200 ;
        RECT 237.800 157.900 238.200 160.200 ;
        RECT 240.600 155.900 241.000 160.200 ;
        RECT 242.200 157.900 242.600 160.200 ;
        RECT 243.800 157.900 244.200 160.200 ;
        RECT 244.600 157.900 245.000 160.200 ;
        RECT 246.200 157.900 246.600 160.200 ;
        RECT 247.300 157.900 247.700 160.200 ;
        RECT 249.400 155.900 249.800 160.200 ;
        RECT 250.200 157.900 250.600 160.200 ;
        RECT 251.800 157.900 252.200 160.200 ;
        RECT 252.900 157.900 253.300 160.200 ;
        RECT 255.000 155.900 255.400 160.200 ;
        RECT 256.600 155.900 257.000 160.200 ;
        RECT 259.400 157.900 259.800 160.200 ;
        RECT 261.000 157.900 261.400 160.200 ;
        RECT 263.800 156.000 264.200 160.200 ;
        RECT 1.400 140.800 1.800 145.000 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.100 ;
        RECT 10.500 140.800 10.900 143.100 ;
        RECT 12.600 140.800 13.000 145.100 ;
        RECT 13.400 140.800 13.800 145.100 ;
        RECT 15.500 140.800 15.900 143.100 ;
        RECT 16.600 140.800 17.000 143.100 ;
        RECT 18.200 140.800 18.600 143.100 ;
        RECT 19.800 140.800 20.200 144.900 ;
        RECT 22.400 140.800 22.800 145.100 ;
        RECT 23.800 140.800 24.200 145.100 ;
        RECT 25.400 140.800 25.800 145.100 ;
        RECT 27.000 140.800 27.400 145.100 ;
        RECT 28.600 140.800 29.000 145.100 ;
        RECT 30.200 140.800 30.600 145.100 ;
        RECT 31.800 140.800 32.200 144.900 ;
        RECT 34.400 140.800 34.800 145.100 ;
        RECT 36.600 140.800 37.000 143.100 ;
        RECT 38.200 140.800 38.600 144.900 ;
        RECT 40.800 140.800 41.200 145.100 ;
        RECT 42.200 140.800 42.600 145.100 ;
        RECT 43.800 140.800 44.200 145.100 ;
        RECT 45.400 140.800 45.800 145.100 ;
        RECT 47.000 140.800 47.400 145.100 ;
        RECT 48.600 140.800 49.000 145.100 ;
        RECT 50.200 140.800 50.600 145.000 ;
        RECT 53.000 140.800 53.400 143.100 ;
        RECT 54.600 140.800 55.000 143.100 ;
        RECT 57.400 140.800 57.800 145.100 ;
        RECT 60.600 140.800 61.000 145.100 ;
        RECT 62.700 140.800 63.100 143.100 ;
        RECT 63.800 140.800 64.200 143.100 ;
        RECT 65.400 140.800 65.800 143.100 ;
        RECT 67.000 140.800 67.400 144.900 ;
        RECT 69.600 140.800 70.000 145.100 ;
        RECT 71.800 140.800 72.200 144.900 ;
        RECT 74.400 140.800 74.800 145.100 ;
        RECT 76.600 140.800 77.000 145.100 ;
        RECT 79.400 140.800 79.800 143.100 ;
        RECT 81.000 140.800 81.400 143.100 ;
        RECT 83.800 140.800 84.200 145.000 ;
        RECT 85.400 140.800 85.800 143.100 ;
        RECT 87.600 140.800 88.000 145.100 ;
        RECT 90.200 140.800 90.600 144.900 ;
        RECT 91.800 140.800 92.200 143.100 ;
        RECT 94.000 140.800 94.400 145.100 ;
        RECT 96.600 140.800 97.000 144.900 ;
        RECT 99.000 140.800 99.400 142.900 ;
        RECT 100.600 140.800 101.000 143.100 ;
        RECT 101.400 140.800 101.800 143.100 ;
        RECT 103.000 140.800 103.400 142.900 ;
        RECT 106.200 140.800 106.600 143.100 ;
        RECT 107.800 140.800 108.200 142.900 ;
        RECT 110.200 140.800 110.600 145.000 ;
        RECT 113.000 140.800 113.400 143.100 ;
        RECT 114.600 140.800 115.000 143.100 ;
        RECT 117.400 140.800 117.800 145.100 ;
        RECT 120.600 140.800 121.000 144.500 ;
        RECT 123.000 140.800 123.400 145.100 ;
        RECT 125.800 140.800 126.200 143.100 ;
        RECT 127.400 140.800 127.800 143.100 ;
        RECT 130.200 140.800 130.600 145.000 ;
        RECT 131.800 140.800 132.200 143.100 ;
        RECT 133.400 140.800 133.800 143.100 ;
        RECT 135.000 140.800 135.400 145.100 ;
        RECT 135.800 140.800 136.200 145.100 ;
        RECT 139.000 140.800 139.400 144.500 ;
        RECT 140.600 140.800 141.000 145.100 ;
        RECT 142.200 140.800 142.600 142.900 ;
        RECT 143.800 140.800 144.200 143.100 ;
        RECT 144.600 140.800 145.000 143.100 ;
        RECT 146.200 140.800 146.600 142.900 ;
        RECT 147.800 140.800 148.200 143.100 ;
        RECT 149.400 140.800 149.800 142.900 ;
        RECT 151.800 140.800 152.200 144.500 ;
        RECT 153.400 140.800 153.800 145.100 ;
        RECT 154.200 140.800 154.600 143.100 ;
        RECT 155.800 140.800 156.200 143.100 ;
        RECT 158.200 140.800 158.600 143.100 ;
        RECT 159.800 140.800 160.200 143.100 ;
        RECT 161.400 140.800 161.800 142.900 ;
        RECT 163.000 140.800 163.400 143.100 ;
        RECT 163.800 140.800 164.200 145.100 ;
        RECT 165.400 140.800 165.800 145.100 ;
        RECT 167.000 140.800 167.400 145.100 ;
        RECT 168.600 140.800 169.000 145.100 ;
        RECT 171.400 140.800 171.800 143.100 ;
        RECT 173.000 140.800 173.400 143.100 ;
        RECT 175.800 140.800 176.200 145.000 ;
        RECT 178.200 140.800 178.600 144.900 ;
        RECT 180.800 140.800 181.200 145.100 ;
        RECT 183.000 140.800 183.400 143.100 ;
        RECT 184.600 140.800 185.000 144.500 ;
        RECT 186.200 140.800 186.600 145.100 ;
        RECT 187.800 140.800 188.200 145.100 ;
        RECT 190.600 140.800 191.000 143.100 ;
        RECT 192.200 140.800 192.600 143.100 ;
        RECT 195.000 140.800 195.400 145.000 ;
        RECT 197.200 140.800 197.600 145.100 ;
        RECT 199.800 140.800 200.200 144.900 ;
        RECT 201.400 140.800 201.800 145.100 ;
        RECT 203.500 140.800 203.900 143.100 ;
        RECT 204.900 140.800 205.300 143.100 ;
        RECT 207.000 140.800 207.400 145.100 ;
        RECT 210.200 140.800 210.600 145.100 ;
        RECT 213.000 140.800 213.400 143.100 ;
        RECT 214.600 140.800 215.000 143.100 ;
        RECT 217.400 140.800 217.800 145.000 ;
        RECT 219.800 140.800 220.200 144.500 ;
        RECT 221.400 140.800 221.800 145.100 ;
        RECT 222.800 140.800 223.200 145.100 ;
        RECT 225.400 140.800 225.800 144.900 ;
        RECT 227.000 140.800 227.400 143.100 ;
        RECT 228.600 140.800 229.000 143.100 ;
        RECT 229.700 140.800 230.100 143.100 ;
        RECT 231.800 140.800 232.200 145.100 ;
        RECT 233.400 140.800 233.800 145.000 ;
        RECT 236.200 140.800 236.600 143.100 ;
        RECT 237.800 140.800 238.200 143.100 ;
        RECT 240.600 140.800 241.000 145.100 ;
        RECT 242.200 140.800 242.600 145.100 ;
        RECT 244.300 140.800 244.700 143.100 ;
        RECT 245.400 140.800 245.800 143.100 ;
        RECT 247.000 140.800 247.400 143.100 ;
        RECT 247.800 140.800 248.200 143.100 ;
        RECT 249.400 140.800 249.800 143.100 ;
        RECT 251.000 140.800 251.400 145.100 ;
        RECT 253.800 140.800 254.200 143.100 ;
        RECT 255.400 140.800 255.800 143.100 ;
        RECT 258.200 140.800 258.600 145.000 ;
        RECT 259.800 140.800 260.200 145.100 ;
        RECT 261.400 140.800 261.800 145.100 ;
        RECT 263.000 140.800 263.400 145.100 ;
        RECT 0.200 140.200 265.400 140.800 ;
        RECT 1.400 136.000 1.800 140.200 ;
        RECT 4.200 137.900 4.600 140.200 ;
        RECT 5.800 137.900 6.200 140.200 ;
        RECT 8.600 135.900 9.000 140.200 ;
        RECT 10.200 135.900 10.600 140.200 ;
        RECT 14.200 136.500 14.600 140.200 ;
        RECT 16.400 135.900 16.800 140.200 ;
        RECT 19.000 136.100 19.400 140.200 ;
        RECT 21.200 135.900 21.600 140.200 ;
        RECT 23.800 136.100 24.200 140.200 ;
        RECT 25.400 135.900 25.800 140.200 ;
        RECT 27.000 136.500 27.400 140.200 ;
        RECT 29.200 135.900 29.600 140.200 ;
        RECT 31.800 136.100 32.200 140.200 ;
        RECT 34.200 137.900 34.600 140.200 ;
        RECT 35.800 135.900 36.200 140.200 ;
        RECT 38.600 137.900 39.000 140.200 ;
        RECT 40.200 137.900 40.600 140.200 ;
        RECT 43.000 136.000 43.400 140.200 ;
        RECT 45.400 136.000 45.800 140.200 ;
        RECT 48.200 137.900 48.600 140.200 ;
        RECT 49.800 137.900 50.200 140.200 ;
        RECT 52.600 135.900 53.000 140.200 ;
        RECT 55.800 135.900 56.200 140.200 ;
        RECT 57.900 137.900 58.300 140.200 ;
        RECT 59.000 135.900 59.400 140.200 ;
        RECT 60.600 135.900 61.000 140.200 ;
        RECT 62.200 135.900 62.600 140.200 ;
        RECT 63.800 135.900 64.200 140.200 ;
        RECT 65.400 135.900 65.800 140.200 ;
        RECT 66.200 135.900 66.600 140.200 ;
        RECT 67.800 136.500 68.200 140.200 ;
        RECT 69.400 135.900 69.800 140.200 ;
        RECT 71.000 136.500 71.400 140.200 ;
        RECT 73.400 136.100 73.800 140.200 ;
        RECT 76.000 135.900 76.400 140.200 ;
        RECT 78.200 136.000 78.600 140.200 ;
        RECT 81.000 137.900 81.400 140.200 ;
        RECT 82.600 137.900 83.000 140.200 ;
        RECT 85.400 135.900 85.800 140.200 ;
        RECT 87.300 137.900 87.700 140.200 ;
        RECT 89.400 135.900 89.800 140.200 ;
        RECT 91.000 135.900 91.400 140.200 ;
        RECT 93.800 137.900 94.200 140.200 ;
        RECT 95.400 137.900 95.800 140.200 ;
        RECT 98.200 136.000 98.600 140.200 ;
        RECT 100.600 138.100 101.000 140.200 ;
        RECT 102.200 137.900 102.600 140.200 ;
        RECT 103.000 137.900 103.400 140.200 ;
        RECT 104.600 137.900 105.000 140.200 ;
        RECT 109.400 136.500 109.800 140.200 ;
        RECT 111.800 136.000 112.200 140.200 ;
        RECT 114.600 137.900 115.000 140.200 ;
        RECT 116.200 137.900 116.600 140.200 ;
        RECT 119.000 135.900 119.400 140.200 ;
        RECT 120.600 135.900 121.000 140.200 ;
        RECT 122.700 137.900 123.100 140.200 ;
        RECT 123.800 137.900 124.200 140.200 ;
        RECT 125.400 137.900 125.800 140.200 ;
        RECT 126.200 135.900 126.600 140.200 ;
        RECT 127.800 135.900 128.200 140.200 ;
        RECT 129.400 135.900 129.800 140.200 ;
        RECT 131.000 135.900 131.400 140.200 ;
        RECT 132.600 135.900 133.000 140.200 ;
        RECT 133.400 135.900 133.800 140.200 ;
        RECT 135.000 136.500 135.400 140.200 ;
        RECT 136.600 135.900 137.000 140.200 ;
        RECT 138.200 137.900 138.600 140.200 ;
        RECT 139.800 137.900 140.200 140.200 ;
        RECT 140.600 137.900 141.000 140.200 ;
        RECT 142.200 137.900 142.600 140.200 ;
        RECT 143.000 137.900 143.400 140.200 ;
        RECT 144.600 137.900 145.000 140.200 ;
        RECT 145.400 137.900 145.800 140.200 ;
        RECT 147.000 137.900 147.400 140.200 ;
        RECT 149.400 135.900 149.800 140.200 ;
        RECT 151.800 135.900 152.200 140.200 ;
        RECT 152.600 137.900 153.000 140.200 ;
        RECT 154.200 137.900 154.600 140.200 ;
        RECT 155.000 137.900 155.400 140.200 ;
        RECT 156.600 137.900 157.000 140.200 ;
        RECT 159.000 137.900 159.400 140.200 ;
        RECT 160.600 137.900 161.000 140.200 ;
        RECT 161.400 135.900 161.800 140.200 ;
        RECT 163.800 137.900 164.200 140.200 ;
        RECT 165.400 137.900 165.800 140.200 ;
        RECT 166.200 135.900 166.600 140.200 ;
        RECT 169.400 135.900 169.800 140.200 ;
        RECT 172.200 137.900 172.600 140.200 ;
        RECT 173.800 137.900 174.200 140.200 ;
        RECT 176.600 136.000 177.000 140.200 ;
        RECT 179.000 136.100 179.400 140.200 ;
        RECT 181.600 135.900 182.000 140.200 ;
        RECT 183.800 137.900 184.200 140.200 ;
        RECT 185.400 136.000 185.800 140.200 ;
        RECT 188.200 137.900 188.600 140.200 ;
        RECT 189.800 137.900 190.200 140.200 ;
        RECT 192.600 135.900 193.000 140.200 ;
        RECT 194.200 135.900 194.600 140.200 ;
        RECT 196.400 135.900 196.800 140.200 ;
        RECT 199.000 136.100 199.400 140.200 ;
        RECT 203.000 136.500 203.400 140.200 ;
        RECT 204.600 137.900 205.000 140.200 ;
        RECT 206.200 137.900 206.600 140.200 ;
        RECT 207.800 135.900 208.200 140.200 ;
        RECT 211.000 136.500 211.400 140.200 ;
        RECT 212.600 135.900 213.000 140.200 ;
        RECT 214.000 135.900 214.400 140.200 ;
        RECT 216.600 136.100 217.000 140.200 ;
        RECT 219.800 136.500 220.200 140.200 ;
        RECT 223.000 135.900 223.400 140.200 ;
        RECT 224.600 135.900 225.000 140.200 ;
        RECT 227.400 137.900 227.800 140.200 ;
        RECT 229.000 137.900 229.400 140.200 ;
        RECT 231.800 136.000 232.200 140.200 ;
        RECT 233.400 135.900 233.800 140.200 ;
        RECT 235.000 135.900 235.400 140.200 ;
        RECT 236.600 135.900 237.000 140.200 ;
        RECT 238.200 135.900 238.600 140.200 ;
        RECT 239.800 135.900 240.200 140.200 ;
        RECT 241.400 136.500 241.800 140.200 ;
        RECT 244.600 135.900 245.000 140.200 ;
        RECT 247.400 137.900 247.800 140.200 ;
        RECT 249.000 137.900 249.400 140.200 ;
        RECT 251.800 136.000 252.200 140.200 ;
        RECT 254.200 136.500 254.600 140.200 ;
        RECT 256.600 135.900 257.000 140.200 ;
        RECT 259.000 135.900 259.400 140.200 ;
        RECT 262.200 136.500 262.600 140.200 ;
        RECT 0.600 120.800 1.000 125.100 ;
        RECT 2.200 120.800 2.600 125.100 ;
        RECT 3.800 120.800 4.200 125.100 ;
        RECT 5.400 120.800 5.800 125.100 ;
        RECT 7.000 120.800 7.400 125.100 ;
        RECT 8.600 120.800 9.000 125.000 ;
        RECT 11.400 120.800 11.800 123.100 ;
        RECT 13.000 120.800 13.400 123.100 ;
        RECT 15.800 120.800 16.200 125.100 ;
        RECT 17.400 120.800 17.800 123.100 ;
        RECT 19.000 120.800 19.400 123.100 ;
        RECT 20.100 120.800 20.500 123.100 ;
        RECT 22.200 120.800 22.600 125.100 ;
        RECT 23.600 120.800 24.000 125.100 ;
        RECT 26.200 120.800 26.600 124.900 ;
        RECT 28.600 120.800 29.000 125.000 ;
        RECT 31.400 120.800 31.800 123.100 ;
        RECT 33.000 120.800 33.400 123.100 ;
        RECT 35.800 120.800 36.200 125.100 ;
        RECT 37.400 120.800 37.800 125.100 ;
        RECT 39.500 120.800 39.900 123.100 ;
        RECT 40.600 120.800 41.000 123.100 ;
        RECT 42.200 120.800 42.600 123.100 ;
        RECT 43.800 120.800 44.200 124.500 ;
        RECT 47.600 120.800 48.000 125.100 ;
        RECT 50.200 120.800 50.600 124.900 ;
        RECT 52.400 120.800 52.800 125.100 ;
        RECT 55.000 120.800 55.400 124.900 ;
        RECT 58.200 120.800 58.600 123.100 ;
        RECT 59.800 120.800 60.200 123.100 ;
        RECT 61.400 120.800 61.800 124.900 ;
        RECT 64.000 120.800 64.400 125.100 ;
        RECT 67.800 120.800 68.200 124.500 ;
        RECT 70.200 120.800 70.600 125.000 ;
        RECT 73.000 120.800 73.400 123.100 ;
        RECT 74.600 120.800 75.000 123.100 ;
        RECT 77.400 120.800 77.800 125.100 ;
        RECT 79.000 120.800 79.400 125.100 ;
        RECT 81.100 120.800 81.500 123.100 ;
        RECT 82.200 120.800 82.600 123.100 ;
        RECT 83.800 120.800 84.200 123.100 ;
        RECT 84.600 120.800 85.000 123.100 ;
        RECT 86.200 120.800 86.600 123.100 ;
        RECT 87.800 120.800 88.200 124.900 ;
        RECT 90.400 120.800 90.800 125.100 ;
        RECT 92.600 120.800 93.000 125.100 ;
        RECT 95.400 120.800 95.800 123.100 ;
        RECT 97.000 120.800 97.400 123.100 ;
        RECT 99.800 120.800 100.200 125.000 ;
        RECT 102.200 120.800 102.600 124.500 ;
        RECT 103.800 120.800 104.200 125.100 ;
        RECT 104.600 120.800 105.000 123.100 ;
        RECT 106.200 120.800 106.600 123.100 ;
        RECT 108.600 120.800 109.000 123.100 ;
        RECT 110.200 120.800 110.600 122.900 ;
        RECT 111.800 120.800 112.200 123.100 ;
        RECT 113.400 120.800 113.800 123.100 ;
        RECT 116.600 120.800 117.000 124.500 ;
        RECT 119.000 120.800 119.400 122.900 ;
        RECT 120.600 120.800 121.000 123.100 ;
        RECT 121.400 120.800 121.800 125.100 ;
        RECT 123.000 120.800 123.400 125.100 ;
        RECT 124.600 120.800 125.000 125.100 ;
        RECT 126.200 120.800 126.600 125.100 ;
        RECT 127.800 120.800 128.200 125.100 ;
        RECT 128.600 120.800 129.000 123.100 ;
        RECT 130.200 120.800 130.600 122.900 ;
        RECT 132.600 120.800 133.000 125.000 ;
        RECT 135.400 120.800 135.800 123.100 ;
        RECT 137.000 120.800 137.400 123.100 ;
        RECT 139.800 120.800 140.200 125.100 ;
        RECT 141.400 120.800 141.800 125.100 ;
        RECT 143.500 120.800 143.900 123.100 ;
        RECT 144.600 120.800 145.000 123.100 ;
        RECT 146.200 120.800 146.600 123.100 ;
        RECT 147.800 120.800 148.200 124.900 ;
        RECT 150.400 120.800 150.800 125.100 ;
        RECT 152.400 120.800 152.800 125.100 ;
        RECT 155.000 120.800 155.400 124.900 ;
        RECT 158.200 120.800 158.600 125.100 ;
        RECT 159.800 120.800 160.200 123.100 ;
        RECT 161.400 120.800 161.800 123.100 ;
        RECT 163.000 120.800 163.400 124.900 ;
        RECT 164.600 120.800 165.000 123.100 ;
        RECT 165.400 120.800 165.800 125.100 ;
        RECT 167.800 120.800 168.200 125.100 ;
        RECT 169.900 120.800 170.300 123.100 ;
        RECT 171.000 120.800 171.400 125.100 ;
        RECT 172.600 120.800 173.000 124.500 ;
        RECT 175.000 120.800 175.400 124.500 ;
        RECT 176.600 120.800 177.000 125.100 ;
        RECT 177.400 120.800 177.800 125.100 ;
        RECT 179.000 120.800 179.400 125.100 ;
        RECT 180.600 120.800 181.000 124.500 ;
        RECT 183.000 120.800 183.400 123.100 ;
        RECT 184.600 120.800 185.000 123.100 ;
        RECT 186.200 120.800 186.600 125.000 ;
        RECT 189.000 120.800 189.400 123.100 ;
        RECT 190.600 120.800 191.000 123.100 ;
        RECT 193.400 120.800 193.800 125.100 ;
        RECT 195.000 120.800 195.400 125.100 ;
        RECT 196.600 120.800 197.000 125.100 ;
        RECT 198.200 120.800 198.600 125.100 ;
        RECT 199.800 120.800 200.200 125.100 ;
        RECT 201.400 120.800 201.800 125.100 ;
        RECT 203.000 120.800 203.400 124.500 ;
        RECT 204.600 120.800 205.000 125.100 ;
        RECT 206.700 120.800 207.100 123.100 ;
        RECT 210.200 120.800 210.600 124.900 ;
        RECT 212.800 120.800 213.200 125.100 ;
        RECT 215.000 120.800 215.400 123.100 ;
        RECT 216.600 120.800 217.000 125.000 ;
        RECT 219.400 120.800 219.800 123.100 ;
        RECT 221.000 120.800 221.400 123.100 ;
        RECT 223.800 120.800 224.200 125.100 ;
        RECT 226.200 120.800 226.600 124.900 ;
        RECT 228.800 120.800 229.200 125.100 ;
        RECT 230.200 120.800 230.600 123.100 ;
        RECT 232.600 120.800 233.000 125.100 ;
        RECT 235.400 120.800 235.800 123.100 ;
        RECT 237.000 120.800 237.400 123.100 ;
        RECT 239.800 120.800 240.200 125.000 ;
        RECT 241.400 120.800 241.800 125.100 ;
        RECT 243.000 120.800 243.400 124.500 ;
        RECT 244.600 120.800 245.000 125.100 ;
        RECT 246.700 120.800 247.100 123.100 ;
        RECT 247.800 120.800 248.200 123.100 ;
        RECT 249.400 120.800 249.800 123.100 ;
        RECT 251.000 120.800 251.400 125.100 ;
        RECT 253.800 120.800 254.200 123.100 ;
        RECT 255.400 120.800 255.800 123.100 ;
        RECT 258.200 120.800 258.600 125.000 ;
        RECT 260.600 120.800 261.000 124.500 ;
        RECT 262.200 120.800 262.600 123.100 ;
        RECT 263.800 120.800 264.200 122.900 ;
        RECT 0.200 120.200 265.400 120.800 ;
        RECT 0.600 115.900 1.000 120.200 ;
        RECT 2.200 115.900 2.600 120.200 ;
        RECT 3.800 115.900 4.200 120.200 ;
        RECT 5.400 115.900 5.800 120.200 ;
        RECT 7.000 115.900 7.400 120.200 ;
        RECT 8.600 116.000 9.000 120.200 ;
        RECT 11.400 117.900 11.800 120.200 ;
        RECT 13.000 117.900 13.400 120.200 ;
        RECT 15.800 115.900 16.200 120.200 ;
        RECT 17.400 115.900 17.800 120.200 ;
        RECT 19.500 117.900 19.900 120.200 ;
        RECT 20.600 117.900 21.000 120.200 ;
        RECT 22.200 117.900 22.600 120.200 ;
        RECT 23.800 116.100 24.200 120.200 ;
        RECT 26.400 115.900 26.800 120.200 ;
        RECT 28.600 116.500 29.000 120.200 ;
        RECT 31.000 115.900 31.400 120.200 ;
        RECT 33.400 115.900 33.800 120.200 ;
        RECT 35.000 116.500 35.400 120.200 ;
        RECT 37.400 116.100 37.800 120.200 ;
        RECT 40.000 115.900 40.400 120.200 ;
        RECT 42.200 117.900 42.600 120.200 ;
        RECT 43.800 115.900 44.200 120.200 ;
        RECT 46.600 117.900 47.000 120.200 ;
        RECT 48.200 117.900 48.600 120.200 ;
        RECT 51.000 116.000 51.400 120.200 ;
        RECT 53.400 116.500 53.800 120.200 ;
        RECT 59.000 115.900 59.400 120.200 ;
        RECT 60.600 116.000 61.000 120.200 ;
        RECT 63.400 117.900 63.800 120.200 ;
        RECT 65.000 117.900 65.400 120.200 ;
        RECT 67.800 115.900 68.200 120.200 ;
        RECT 69.400 115.900 69.800 120.200 ;
        RECT 71.500 117.900 71.900 120.200 ;
        RECT 72.600 117.900 73.000 120.200 ;
        RECT 74.200 117.900 74.600 120.200 ;
        RECT 75.800 116.100 76.200 120.200 ;
        RECT 78.400 115.900 78.800 120.200 ;
        RECT 80.600 116.100 81.000 120.200 ;
        RECT 83.200 115.900 83.600 120.200 ;
        RECT 84.600 115.900 85.000 120.200 ;
        RECT 86.700 117.900 87.100 120.200 ;
        RECT 87.800 117.900 88.200 120.200 ;
        RECT 89.400 117.900 89.800 120.200 ;
        RECT 91.000 116.100 91.400 120.200 ;
        RECT 93.600 115.900 94.000 120.200 ;
        RECT 95.800 115.900 96.200 120.200 ;
        RECT 98.600 117.900 99.000 120.200 ;
        RECT 100.200 117.900 100.600 120.200 ;
        RECT 103.000 116.000 103.400 120.200 ;
        RECT 107.000 116.000 107.400 120.200 ;
        RECT 109.800 117.900 110.200 120.200 ;
        RECT 111.400 117.900 111.800 120.200 ;
        RECT 114.200 115.900 114.600 120.200 ;
        RECT 116.600 116.000 117.000 120.200 ;
        RECT 119.400 117.900 119.800 120.200 ;
        RECT 121.000 117.900 121.400 120.200 ;
        RECT 123.800 115.900 124.200 120.200 ;
        RECT 125.400 115.900 125.800 120.200 ;
        RECT 127.500 117.900 127.900 120.200 ;
        RECT 128.600 115.900 129.000 120.200 ;
        RECT 130.700 117.900 131.100 120.200 ;
        RECT 131.800 117.900 132.200 120.200 ;
        RECT 133.400 117.900 133.800 120.200 ;
        RECT 135.000 116.000 135.400 120.200 ;
        RECT 137.800 117.900 138.200 120.200 ;
        RECT 139.400 117.900 139.800 120.200 ;
        RECT 142.200 115.900 142.600 120.200 ;
        RECT 143.800 115.900 144.200 120.200 ;
        RECT 146.200 115.900 146.600 120.200 ;
        RECT 150.200 115.900 150.600 120.200 ;
        RECT 151.800 116.100 152.200 120.200 ;
        RECT 154.400 115.900 154.800 120.200 ;
        RECT 155.800 117.900 156.200 120.200 ;
        RECT 157.400 117.900 157.800 120.200 ;
        RECT 160.100 117.900 160.500 120.200 ;
        RECT 162.200 115.900 162.600 120.200 ;
        RECT 163.800 115.900 164.200 120.200 ;
        RECT 166.600 117.900 167.000 120.200 ;
        RECT 168.200 117.900 168.600 120.200 ;
        RECT 171.000 116.000 171.400 120.200 ;
        RECT 172.600 115.900 173.000 120.200 ;
        RECT 174.200 115.900 174.600 120.200 ;
        RECT 175.800 115.900 176.200 120.200 ;
        RECT 177.400 115.900 177.800 120.200 ;
        RECT 179.000 115.900 179.400 120.200 ;
        RECT 179.800 115.900 180.200 120.200 ;
        RECT 181.400 115.900 181.800 120.200 ;
        RECT 183.000 115.900 183.400 120.200 ;
        RECT 184.600 115.900 185.000 120.200 ;
        RECT 186.200 115.900 186.600 120.200 ;
        RECT 187.000 115.900 187.400 120.200 ;
        RECT 189.400 115.900 189.800 120.200 ;
        RECT 192.200 117.900 192.600 120.200 ;
        RECT 193.800 117.900 194.200 120.200 ;
        RECT 196.600 116.000 197.000 120.200 ;
        RECT 198.200 115.900 198.600 120.200 ;
        RECT 199.800 116.500 200.200 120.200 ;
        RECT 201.400 115.900 201.800 120.200 ;
        RECT 203.000 116.500 203.400 120.200 ;
        RECT 205.200 115.900 205.600 120.200 ;
        RECT 207.800 116.100 208.200 120.200 ;
        RECT 211.000 117.900 211.400 120.200 ;
        RECT 212.600 117.900 213.000 120.200 ;
        RECT 213.400 115.900 213.800 120.200 ;
        RECT 217.400 116.500 217.800 120.200 ;
        RECT 219.800 116.000 220.200 120.200 ;
        RECT 222.600 117.900 223.000 120.200 ;
        RECT 224.200 117.900 224.600 120.200 ;
        RECT 227.000 115.900 227.400 120.200 ;
        RECT 228.600 117.900 229.000 120.200 ;
        RECT 230.200 117.900 230.600 120.200 ;
        RECT 231.300 117.900 231.700 120.200 ;
        RECT 233.400 115.900 233.800 120.200 ;
        RECT 235.000 116.500 235.400 120.200 ;
        RECT 238.200 116.500 238.600 120.200 ;
        RECT 239.800 115.900 240.200 120.200 ;
        RECT 240.600 115.900 241.000 120.200 ;
        RECT 243.800 116.500 244.200 120.200 ;
        RECT 247.000 115.900 247.400 120.200 ;
        RECT 249.800 117.900 250.200 120.200 ;
        RECT 251.400 117.900 251.800 120.200 ;
        RECT 254.200 116.000 254.600 120.200 ;
        RECT 256.600 116.000 257.000 120.200 ;
        RECT 259.400 117.900 259.800 120.200 ;
        RECT 261.000 117.900 261.400 120.200 ;
        RECT 263.800 115.900 264.200 120.200 ;
        RECT 0.600 100.800 1.000 105.100 ;
        RECT 2.200 100.800 2.600 105.100 ;
        RECT 3.800 100.800 4.200 105.100 ;
        RECT 5.400 100.800 5.800 105.000 ;
        RECT 8.200 100.800 8.600 103.100 ;
        RECT 9.800 100.800 10.200 103.100 ;
        RECT 12.600 100.800 13.000 105.100 ;
        RECT 15.000 100.800 15.400 104.500 ;
        RECT 19.000 100.800 19.400 105.100 ;
        RECT 20.600 100.800 21.000 105.000 ;
        RECT 23.400 100.800 23.800 103.100 ;
        RECT 25.000 100.800 25.400 103.100 ;
        RECT 27.800 100.800 28.200 105.100 ;
        RECT 30.200 100.800 30.600 104.900 ;
        RECT 32.800 100.800 33.200 105.100 ;
        RECT 34.200 100.800 34.600 103.100 ;
        RECT 36.400 100.800 36.800 105.100 ;
        RECT 39.000 100.800 39.400 104.900 ;
        RECT 41.200 100.800 41.600 105.100 ;
        RECT 43.800 100.800 44.200 104.900 ;
        RECT 46.200 100.800 46.600 105.100 ;
        RECT 49.000 100.800 49.400 103.100 ;
        RECT 50.600 100.800 51.000 103.100 ;
        RECT 53.400 100.800 53.800 105.000 ;
        RECT 56.600 100.800 57.000 105.100 ;
        RECT 58.200 100.800 58.600 104.500 ;
        RECT 60.600 100.800 61.000 105.000 ;
        RECT 63.400 100.800 63.800 103.100 ;
        RECT 65.000 100.800 65.400 103.100 ;
        RECT 67.800 100.800 68.200 105.100 ;
        RECT 69.400 100.800 69.800 105.100 ;
        RECT 71.500 100.800 71.900 103.100 ;
        RECT 72.600 100.800 73.000 103.100 ;
        RECT 74.200 100.800 74.600 103.100 ;
        RECT 75.800 100.800 76.200 105.000 ;
        RECT 78.600 100.800 79.000 103.100 ;
        RECT 80.200 100.800 80.600 103.100 ;
        RECT 83.000 100.800 83.400 105.100 ;
        RECT 84.600 100.800 85.000 105.100 ;
        RECT 88.600 100.800 89.000 104.500 ;
        RECT 91.000 100.800 91.400 105.000 ;
        RECT 93.800 100.800 94.200 103.100 ;
        RECT 95.400 100.800 95.800 103.100 ;
        RECT 98.200 100.800 98.600 105.100 ;
        RECT 99.800 100.800 100.200 105.100 ;
        RECT 101.400 100.800 101.800 104.500 ;
        RECT 103.800 100.800 104.200 104.500 ;
        RECT 107.800 100.800 108.200 105.100 ;
        RECT 111.000 100.800 111.400 104.900 ;
        RECT 113.600 100.800 114.000 105.100 ;
        RECT 115.800 100.800 116.200 103.100 ;
        RECT 116.600 100.800 117.000 105.100 ;
        RECT 118.200 100.800 118.600 105.100 ;
        RECT 119.800 100.800 120.200 105.100 ;
        RECT 121.400 100.800 121.800 105.100 ;
        RECT 123.000 100.800 123.400 105.100 ;
        RECT 123.800 100.800 124.200 105.100 ;
        RECT 125.400 100.800 125.800 104.500 ;
        RECT 127.000 100.800 127.400 103.100 ;
        RECT 128.600 100.800 129.000 103.100 ;
        RECT 130.200 100.800 130.600 104.900 ;
        RECT 132.800 100.800 133.200 105.100 ;
        RECT 135.000 100.800 135.400 104.900 ;
        RECT 137.600 100.800 138.000 105.100 ;
        RECT 139.000 100.800 139.400 105.100 ;
        RECT 140.600 100.800 141.000 105.100 ;
        RECT 142.200 100.800 142.600 105.100 ;
        RECT 143.000 100.800 143.400 105.100 ;
        RECT 146.500 100.800 146.900 105.100 ;
        RECT 150.200 100.800 150.600 105.100 ;
        RECT 151.800 100.800 152.200 104.500 ;
        RECT 153.400 100.800 153.800 105.100 ;
        RECT 154.800 100.800 155.200 105.100 ;
        RECT 157.400 100.800 157.800 104.900 ;
        RECT 161.400 100.800 161.800 104.500 ;
        RECT 164.600 100.800 165.000 103.100 ;
        RECT 166.200 100.800 166.600 103.100 ;
        RECT 167.800 100.800 168.200 104.500 ;
        RECT 171.800 100.800 172.200 105.100 ;
        RECT 174.600 100.800 175.000 103.100 ;
        RECT 176.200 100.800 176.600 103.100 ;
        RECT 179.000 100.800 179.400 105.000 ;
        RECT 180.600 100.800 181.000 103.100 ;
        RECT 182.200 100.800 182.600 103.100 ;
        RECT 183.300 100.800 183.700 103.100 ;
        RECT 185.400 100.800 185.800 105.100 ;
        RECT 187.000 100.800 187.400 104.500 ;
        RECT 191.000 100.800 191.400 105.100 ;
        RECT 192.600 100.800 193.000 105.100 ;
        RECT 195.400 100.800 195.800 103.100 ;
        RECT 197.000 100.800 197.400 103.100 ;
        RECT 199.800 100.800 200.200 105.000 ;
        RECT 202.200 100.800 202.600 104.500 ;
        RECT 203.800 100.800 204.200 105.100 ;
        RECT 204.600 100.800 205.000 103.100 ;
        RECT 206.200 100.800 206.600 103.100 ;
        RECT 207.000 100.800 207.400 105.100 ;
        RECT 211.000 100.800 211.400 105.100 ;
        RECT 214.200 100.800 214.600 105.100 ;
        RECT 217.000 100.800 217.400 103.100 ;
        RECT 218.600 100.800 219.000 103.100 ;
        RECT 221.400 100.800 221.800 105.000 ;
        RECT 223.000 100.800 223.400 103.100 ;
        RECT 224.600 100.800 225.000 103.100 ;
        RECT 225.400 100.800 225.800 105.100 ;
        RECT 227.800 100.800 228.200 103.100 ;
        RECT 229.400 100.800 229.800 103.100 ;
        RECT 230.200 100.800 230.600 103.100 ;
        RECT 231.800 100.800 232.200 103.100 ;
        RECT 233.400 100.800 233.800 105.100 ;
        RECT 236.200 100.800 236.600 103.100 ;
        RECT 237.800 100.800 238.200 103.100 ;
        RECT 240.600 100.800 241.000 105.000 ;
        RECT 243.000 100.800 243.400 104.500 ;
        RECT 245.400 100.800 245.800 105.100 ;
        RECT 247.000 100.800 247.400 105.100 ;
        RECT 248.600 100.800 249.000 105.100 ;
        RECT 250.200 100.800 250.600 105.100 ;
        RECT 251.800 100.800 252.200 105.100 ;
        RECT 253.400 100.800 253.800 105.000 ;
        RECT 256.200 100.800 256.600 103.100 ;
        RECT 257.800 100.800 258.200 103.100 ;
        RECT 260.600 100.800 261.000 105.100 ;
        RECT 262.200 100.800 262.600 105.100 ;
        RECT 0.200 100.200 265.400 100.800 ;
        RECT 1.400 96.000 1.800 100.200 ;
        RECT 4.200 97.900 4.600 100.200 ;
        RECT 5.800 97.900 6.200 100.200 ;
        RECT 8.600 95.900 9.000 100.200 ;
        RECT 10.200 97.900 10.600 100.200 ;
        RECT 11.800 97.900 12.200 100.200 ;
        RECT 12.900 97.900 13.300 100.200 ;
        RECT 15.000 95.900 15.400 100.200 ;
        RECT 16.600 96.100 17.000 100.200 ;
        RECT 19.200 95.900 19.600 100.200 ;
        RECT 20.600 97.900 21.000 100.200 ;
        RECT 22.200 97.900 22.600 100.200 ;
        RECT 23.800 96.000 24.200 100.200 ;
        RECT 26.600 97.900 27.000 100.200 ;
        RECT 28.200 97.900 28.600 100.200 ;
        RECT 31.000 95.900 31.400 100.200 ;
        RECT 32.600 97.900 33.000 100.200 ;
        RECT 34.200 97.900 34.600 100.200 ;
        RECT 35.300 97.900 35.700 100.200 ;
        RECT 37.400 95.900 37.800 100.200 ;
        RECT 38.200 95.900 38.600 100.200 ;
        RECT 41.200 95.900 41.600 100.200 ;
        RECT 43.800 96.100 44.200 100.200 ;
        RECT 45.400 95.900 45.800 100.200 ;
        RECT 47.500 97.900 47.900 100.200 ;
        RECT 48.600 97.900 49.000 100.200 ;
        RECT 50.200 97.900 50.600 100.200 ;
        RECT 53.400 95.900 53.800 100.200 ;
        RECT 56.200 97.900 56.600 100.200 ;
        RECT 57.800 97.900 58.200 100.200 ;
        RECT 60.600 96.000 61.000 100.200 ;
        RECT 62.500 97.900 62.900 100.200 ;
        RECT 64.600 95.900 65.000 100.200 ;
        RECT 66.200 95.900 66.600 100.200 ;
        RECT 69.000 97.900 69.400 100.200 ;
        RECT 70.600 97.900 71.000 100.200 ;
        RECT 73.400 96.000 73.800 100.200 ;
        RECT 75.000 95.900 75.400 100.200 ;
        RECT 76.600 95.900 77.000 100.200 ;
        RECT 78.200 95.900 78.600 100.200 ;
        RECT 79.800 95.900 80.200 100.200 ;
        RECT 81.400 95.900 81.800 100.200 ;
        RECT 83.000 96.100 83.400 100.200 ;
        RECT 85.600 95.900 86.000 100.200 ;
        RECT 87.600 95.900 88.000 100.200 ;
        RECT 90.200 96.100 90.600 100.200 ;
        RECT 92.600 96.100 93.000 100.200 ;
        RECT 95.200 95.900 95.600 100.200 ;
        RECT 97.400 97.900 97.800 100.200 ;
        RECT 99.000 95.900 99.400 100.200 ;
        RECT 101.800 97.900 102.200 100.200 ;
        RECT 103.400 97.900 103.800 100.200 ;
        RECT 106.200 96.000 106.600 100.200 ;
        RECT 110.200 96.100 110.600 100.200 ;
        RECT 112.800 95.900 113.200 100.200 ;
        RECT 115.000 97.900 115.400 100.200 ;
        RECT 116.600 96.000 117.000 100.200 ;
        RECT 119.400 97.900 119.800 100.200 ;
        RECT 121.000 97.900 121.400 100.200 ;
        RECT 123.800 95.900 124.200 100.200 ;
        RECT 125.400 97.900 125.800 100.200 ;
        RECT 127.000 95.900 127.400 100.200 ;
        RECT 130.200 96.100 130.600 100.200 ;
        RECT 132.800 95.900 133.200 100.200 ;
        RECT 135.000 96.500 135.400 100.200 ;
        RECT 136.600 95.900 137.000 100.200 ;
        RECT 138.200 96.500 138.600 100.200 ;
        RECT 141.400 96.000 141.800 100.200 ;
        RECT 144.200 97.900 144.600 100.200 ;
        RECT 145.800 97.900 146.200 100.200 ;
        RECT 148.600 95.900 149.000 100.200 ;
        RECT 150.200 95.900 150.600 100.200 ;
        RECT 153.200 95.900 153.600 100.200 ;
        RECT 155.800 96.100 156.200 100.200 ;
        RECT 159.000 97.900 159.400 100.200 ;
        RECT 160.600 97.900 161.000 100.200 ;
        RECT 162.200 96.000 162.600 100.200 ;
        RECT 165.000 97.900 165.400 100.200 ;
        RECT 166.600 97.900 167.000 100.200 ;
        RECT 169.400 95.900 169.800 100.200 ;
        RECT 171.000 97.900 171.400 100.200 ;
        RECT 172.600 97.900 173.000 100.200 ;
        RECT 173.700 97.900 174.100 100.200 ;
        RECT 175.800 95.900 176.200 100.200 ;
        RECT 177.200 95.900 177.600 100.200 ;
        RECT 179.800 96.100 180.200 100.200 ;
        RECT 182.000 95.900 182.400 100.200 ;
        RECT 184.600 96.100 185.000 100.200 ;
        RECT 186.800 95.900 187.200 100.200 ;
        RECT 189.400 96.100 189.800 100.200 ;
        RECT 191.000 97.900 191.400 100.200 ;
        RECT 192.600 97.900 193.000 100.200 ;
        RECT 193.400 95.900 193.800 100.200 ;
        RECT 195.000 96.500 195.400 100.200 ;
        RECT 196.600 95.900 197.000 100.200 ;
        RECT 198.200 96.500 198.600 100.200 ;
        RECT 199.800 95.900 200.200 100.200 ;
        RECT 201.400 96.500 201.800 100.200 ;
        RECT 203.800 96.500 204.200 100.200 ;
        RECT 205.400 95.900 205.800 100.200 ;
        RECT 208.600 95.900 209.000 100.200 ;
        RECT 211.400 97.900 211.800 100.200 ;
        RECT 213.000 97.900 213.400 100.200 ;
        RECT 215.800 96.000 216.200 100.200 ;
        RECT 217.400 97.900 217.800 100.200 ;
        RECT 219.000 97.900 219.400 100.200 ;
        RECT 220.600 96.000 221.000 100.200 ;
        RECT 223.400 97.900 223.800 100.200 ;
        RECT 225.000 97.900 225.400 100.200 ;
        RECT 227.800 95.900 228.200 100.200 ;
        RECT 229.400 95.900 229.800 100.200 ;
        RECT 231.000 96.500 231.400 100.200 ;
        RECT 234.200 96.500 234.600 100.200 ;
        RECT 235.800 97.900 236.200 100.200 ;
        RECT 237.400 97.900 237.800 100.200 ;
        RECT 239.000 97.900 239.400 100.200 ;
        RECT 240.600 95.900 241.000 100.200 ;
        RECT 243.400 97.900 243.800 100.200 ;
        RECT 245.000 97.900 245.400 100.200 ;
        RECT 247.800 96.000 248.200 100.200 ;
        RECT 249.400 97.900 249.800 100.200 ;
        RECT 251.000 97.900 251.400 100.200 ;
        RECT 252.600 96.500 253.000 100.200 ;
        RECT 255.800 96.500 256.200 100.200 ;
        RECT 257.400 95.900 257.800 100.200 ;
        RECT 259.800 97.900 260.200 100.200 ;
        RECT 261.400 97.900 261.800 100.200 ;
        RECT 263.000 96.500 263.400 100.200 ;
        RECT 1.400 80.800 1.800 85.000 ;
        RECT 4.200 80.800 4.600 83.100 ;
        RECT 5.800 80.800 6.200 83.100 ;
        RECT 8.600 80.800 9.000 85.100 ;
        RECT 10.200 80.800 10.600 83.100 ;
        RECT 12.400 80.800 12.800 85.100 ;
        RECT 15.000 80.800 15.400 84.900 ;
        RECT 17.400 80.800 17.800 85.100 ;
        RECT 20.200 80.800 20.600 83.100 ;
        RECT 21.800 80.800 22.200 83.100 ;
        RECT 24.600 80.800 25.000 85.000 ;
        RECT 26.500 80.800 26.900 83.100 ;
        RECT 28.600 80.800 29.000 85.100 ;
        RECT 30.200 80.800 30.600 85.000 ;
        RECT 33.000 80.800 33.400 83.100 ;
        RECT 34.600 80.800 35.000 83.100 ;
        RECT 37.400 80.800 37.800 85.100 ;
        RECT 40.600 80.800 41.000 84.500 ;
        RECT 42.800 80.800 43.200 85.100 ;
        RECT 45.400 80.800 45.800 84.900 ;
        RECT 47.800 80.800 48.200 84.900 ;
        RECT 50.400 80.800 50.800 85.100 ;
        RECT 52.400 80.800 52.800 85.100 ;
        RECT 55.000 80.800 55.400 84.900 ;
        RECT 58.200 80.800 58.600 83.100 ;
        RECT 59.800 80.800 60.200 83.100 ;
        RECT 61.400 80.800 61.800 85.100 ;
        RECT 64.200 80.800 64.600 83.100 ;
        RECT 65.800 80.800 66.200 83.100 ;
        RECT 68.600 80.800 69.000 85.000 ;
        RECT 70.200 80.800 70.600 83.100 ;
        RECT 71.800 80.800 72.200 83.100 ;
        RECT 72.900 80.800 73.300 83.100 ;
        RECT 75.000 80.800 75.400 85.100 ;
        RECT 78.200 80.800 78.600 84.500 ;
        RECT 80.400 80.800 80.800 85.100 ;
        RECT 83.000 80.800 83.400 84.900 ;
        RECT 84.600 80.800 85.000 85.100 ;
        RECT 86.200 80.800 86.600 85.100 ;
        RECT 87.800 80.800 88.200 85.100 ;
        RECT 89.400 80.800 89.800 85.100 ;
        RECT 91.000 80.800 91.400 85.100 ;
        RECT 91.800 80.800 92.200 83.100 ;
        RECT 94.200 80.800 94.600 85.100 ;
        RECT 97.000 80.800 97.400 83.100 ;
        RECT 98.600 80.800 99.000 83.100 ;
        RECT 101.400 80.800 101.800 85.000 ;
        RECT 103.800 80.800 104.200 84.900 ;
        RECT 106.400 80.800 106.800 85.100 ;
        RECT 110.200 80.800 110.600 85.000 ;
        RECT 113.000 80.800 113.400 83.100 ;
        RECT 114.600 80.800 115.000 83.100 ;
        RECT 117.400 80.800 117.800 85.100 ;
        RECT 119.000 80.800 119.400 83.100 ;
        RECT 121.200 80.800 121.600 85.100 ;
        RECT 123.800 80.800 124.200 84.900 ;
        RECT 126.200 80.800 126.600 85.000 ;
        RECT 129.000 80.800 129.400 83.100 ;
        RECT 130.600 80.800 131.000 83.100 ;
        RECT 133.400 80.800 133.800 85.100 ;
        RECT 135.000 80.800 135.400 83.100 ;
        RECT 137.200 80.800 137.600 85.100 ;
        RECT 139.800 80.800 140.200 84.900 ;
        RECT 142.000 80.800 142.400 85.100 ;
        RECT 144.600 80.800 145.000 84.900 ;
        RECT 146.200 80.800 146.600 83.100 ;
        RECT 147.800 80.800 148.200 84.900 ;
        RECT 149.400 80.800 149.800 85.100 ;
        RECT 151.800 80.800 152.200 85.100 ;
        RECT 154.600 80.800 155.000 83.100 ;
        RECT 156.200 80.800 156.600 83.100 ;
        RECT 159.000 80.800 159.400 85.000 ;
        RECT 162.500 80.800 162.900 83.100 ;
        RECT 164.600 80.800 165.000 85.100 ;
        RECT 166.000 80.800 166.400 85.100 ;
        RECT 168.600 80.800 169.000 84.900 ;
        RECT 171.000 80.800 171.400 85.000 ;
        RECT 173.800 80.800 174.200 83.100 ;
        RECT 175.400 80.800 175.800 83.100 ;
        RECT 178.200 80.800 178.600 85.100 ;
        RECT 180.100 80.800 180.500 83.100 ;
        RECT 182.200 80.800 182.600 85.100 ;
        RECT 183.300 80.800 183.700 83.100 ;
        RECT 185.400 80.800 185.800 85.100 ;
        RECT 186.200 80.800 186.600 85.100 ;
        RECT 188.300 80.800 188.700 83.100 ;
        RECT 190.200 80.800 190.600 85.100 ;
        RECT 193.000 80.800 193.400 83.100 ;
        RECT 194.600 80.800 195.000 83.100 ;
        RECT 197.400 80.800 197.800 85.000 ;
        RECT 199.000 80.800 199.400 85.100 ;
        RECT 200.600 80.800 201.000 85.100 ;
        RECT 202.200 80.800 202.600 85.100 ;
        RECT 203.800 80.800 204.200 85.100 ;
        RECT 205.400 80.800 205.800 85.100 ;
        RECT 206.200 80.800 206.600 85.100 ;
        RECT 207.800 80.800 208.200 85.100 ;
        RECT 209.400 80.800 209.800 85.100 ;
        RECT 212.100 80.800 212.500 83.100 ;
        RECT 214.200 80.800 214.600 85.100 ;
        RECT 215.300 80.800 215.700 83.100 ;
        RECT 217.400 80.800 217.800 85.100 ;
        RECT 219.000 80.800 219.400 84.500 ;
        RECT 221.700 80.800 222.100 83.100 ;
        RECT 223.800 80.800 224.200 85.100 ;
        RECT 224.600 80.800 225.000 85.100 ;
        RECT 226.200 80.800 226.600 84.500 ;
        RECT 227.800 80.800 228.200 85.100 ;
        RECT 229.900 80.800 230.300 83.100 ;
        RECT 231.800 80.800 232.200 85.000 ;
        RECT 234.600 80.800 235.000 83.100 ;
        RECT 236.200 80.800 236.600 83.100 ;
        RECT 239.000 80.800 239.400 85.100 ;
        RECT 240.600 80.800 241.000 85.100 ;
        RECT 242.200 80.800 242.600 85.100 ;
        RECT 243.800 80.800 244.200 85.100 ;
        RECT 245.400 80.800 245.800 85.100 ;
        RECT 247.000 80.800 247.400 85.100 ;
        RECT 247.800 80.800 248.200 85.100 ;
        RECT 249.400 80.800 249.800 85.100 ;
        RECT 251.000 80.800 251.400 85.100 ;
        RECT 252.600 80.800 253.000 85.100 ;
        RECT 254.200 80.800 254.600 85.100 ;
        RECT 256.600 80.800 257.000 84.500 ;
        RECT 258.200 80.800 258.600 85.100 ;
        RECT 259.800 80.800 260.200 85.100 ;
        RECT 261.400 80.800 261.800 85.100 ;
        RECT 263.000 80.800 263.400 85.100 ;
        RECT 264.600 80.800 265.000 85.100 ;
        RECT 0.200 80.200 265.400 80.800 ;
        RECT 1.400 76.000 1.800 80.200 ;
        RECT 4.200 77.900 4.600 80.200 ;
        RECT 5.800 77.900 6.200 80.200 ;
        RECT 8.600 75.900 9.000 80.200 ;
        RECT 10.200 77.900 10.600 80.200 ;
        RECT 11.800 77.900 12.200 80.200 ;
        RECT 12.900 77.900 13.300 80.200 ;
        RECT 15.000 75.900 15.400 80.200 ;
        RECT 16.600 76.000 17.000 80.200 ;
        RECT 19.400 77.900 19.800 80.200 ;
        RECT 21.000 77.900 21.400 80.200 ;
        RECT 23.800 75.900 24.200 80.200 ;
        RECT 27.000 75.900 27.400 80.200 ;
        RECT 29.400 76.500 29.800 80.200 ;
        RECT 31.800 76.000 32.200 80.200 ;
        RECT 34.600 77.900 35.000 80.200 ;
        RECT 36.200 77.900 36.600 80.200 ;
        RECT 39.000 75.900 39.400 80.200 ;
        RECT 41.400 76.100 41.800 80.200 ;
        RECT 44.000 75.900 44.400 80.200 ;
        RECT 46.200 77.900 46.600 80.200 ;
        RECT 47.800 75.900 48.200 80.200 ;
        RECT 50.600 77.900 51.000 80.200 ;
        RECT 52.200 77.900 52.600 80.200 ;
        RECT 55.000 76.000 55.400 80.200 ;
        RECT 59.000 75.900 59.400 80.200 ;
        RECT 61.800 77.900 62.200 80.200 ;
        RECT 63.400 77.900 63.800 80.200 ;
        RECT 66.200 76.000 66.600 80.200 ;
        RECT 67.800 77.900 68.200 80.200 ;
        RECT 69.400 77.900 69.800 80.200 ;
        RECT 70.500 77.900 70.900 80.200 ;
        RECT 72.600 75.900 73.000 80.200 ;
        RECT 74.200 76.100 74.600 80.200 ;
        RECT 76.800 75.900 77.200 80.200 ;
        RECT 79.000 77.900 79.400 80.200 ;
        RECT 80.600 75.900 81.000 80.200 ;
        RECT 83.400 77.900 83.800 80.200 ;
        RECT 85.000 77.900 85.400 80.200 ;
        RECT 87.800 76.000 88.200 80.200 ;
        RECT 89.400 77.900 89.800 80.200 ;
        RECT 91.000 77.900 91.400 80.200 ;
        RECT 92.600 76.100 93.000 80.200 ;
        RECT 94.200 77.900 94.600 80.200 ;
        RECT 95.000 77.900 95.400 80.200 ;
        RECT 96.600 77.900 97.000 80.200 ;
        RECT 97.400 75.900 97.800 80.200 ;
        RECT 99.000 76.500 99.400 80.200 ;
        RECT 101.400 76.500 101.800 80.200 ;
        RECT 103.000 75.900 103.400 80.200 ;
        RECT 103.800 75.900 104.200 80.200 ;
        RECT 105.900 77.900 106.300 80.200 ;
        RECT 108.600 77.900 109.000 80.200 ;
        RECT 110.200 77.900 110.600 80.200 ;
        RECT 111.800 76.000 112.200 80.200 ;
        RECT 114.600 77.900 115.000 80.200 ;
        RECT 116.200 77.900 116.600 80.200 ;
        RECT 119.000 75.900 119.400 80.200 ;
        RECT 120.600 75.900 121.000 80.200 ;
        RECT 122.200 75.900 122.600 80.200 ;
        RECT 123.800 75.900 124.200 80.200 ;
        RECT 125.400 75.900 125.800 80.200 ;
        RECT 127.000 75.900 127.400 80.200 ;
        RECT 127.800 77.900 128.200 80.200 ;
        RECT 129.400 77.900 129.800 80.200 ;
        RECT 131.000 76.000 131.400 80.200 ;
        RECT 133.800 77.900 134.200 80.200 ;
        RECT 135.400 77.900 135.800 80.200 ;
        RECT 138.200 75.900 138.600 80.200 ;
        RECT 139.800 75.900 140.200 80.200 ;
        RECT 143.000 76.100 143.400 80.200 ;
        RECT 145.600 75.900 146.000 80.200 ;
        RECT 147.800 76.000 148.200 80.200 ;
        RECT 150.600 77.900 151.000 80.200 ;
        RECT 152.200 77.900 152.600 80.200 ;
        RECT 155.000 75.900 155.400 80.200 ;
        RECT 158.200 77.900 158.600 80.200 ;
        RECT 159.800 77.900 160.200 80.200 ;
        RECT 160.600 77.900 161.000 80.200 ;
        RECT 162.200 76.100 162.600 80.200 ;
        RECT 164.100 77.900 164.500 80.200 ;
        RECT 166.200 75.900 166.600 80.200 ;
        RECT 167.600 75.900 168.000 80.200 ;
        RECT 170.200 76.100 170.600 80.200 ;
        RECT 172.600 76.100 173.000 80.200 ;
        RECT 175.200 75.900 175.600 80.200 ;
        RECT 177.400 75.900 177.800 80.200 ;
        RECT 180.200 77.900 180.600 80.200 ;
        RECT 181.800 77.900 182.200 80.200 ;
        RECT 184.600 76.000 185.000 80.200 ;
        RECT 186.200 75.900 186.600 80.200 ;
        RECT 190.200 76.500 190.600 80.200 ;
        RECT 192.400 75.900 192.800 80.200 ;
        RECT 195.000 76.100 195.400 80.200 ;
        RECT 196.900 77.900 197.300 80.200 ;
        RECT 199.000 75.900 199.400 80.200 ;
        RECT 199.800 75.900 200.200 80.200 ;
        RECT 201.400 75.900 201.800 80.200 ;
        RECT 203.000 75.900 203.400 80.200 ;
        RECT 204.600 75.900 205.000 80.200 ;
        RECT 206.200 75.900 206.600 80.200 ;
        RECT 208.900 77.900 209.300 80.200 ;
        RECT 211.000 75.900 211.400 80.200 ;
        RECT 212.600 76.000 213.000 80.200 ;
        RECT 215.400 77.900 215.800 80.200 ;
        RECT 217.000 77.900 217.400 80.200 ;
        RECT 219.800 75.900 220.200 80.200 ;
        RECT 221.700 77.900 222.100 80.200 ;
        RECT 223.800 75.900 224.200 80.200 ;
        RECT 224.600 77.900 225.000 80.200 ;
        RECT 226.200 77.900 226.600 80.200 ;
        RECT 227.000 75.900 227.400 80.200 ;
        RECT 229.100 77.900 229.500 80.200 ;
        RECT 230.500 77.900 230.900 80.200 ;
        RECT 232.600 75.900 233.000 80.200 ;
        RECT 234.200 75.900 234.600 80.200 ;
        RECT 237.000 77.900 237.400 80.200 ;
        RECT 238.600 77.900 239.000 80.200 ;
        RECT 241.400 76.000 241.800 80.200 ;
        RECT 243.800 76.500 244.200 80.200 ;
        RECT 247.000 75.900 247.400 80.200 ;
        RECT 249.800 77.900 250.200 80.200 ;
        RECT 251.400 77.900 251.800 80.200 ;
        RECT 254.200 76.000 254.600 80.200 ;
        RECT 256.600 75.900 257.000 80.200 ;
        RECT 259.400 77.900 259.800 80.200 ;
        RECT 261.000 77.900 261.400 80.200 ;
        RECT 263.800 76.000 264.200 80.200 ;
        RECT 0.600 60.800 1.000 65.100 ;
        RECT 2.200 60.800 2.600 65.100 ;
        RECT 3.800 60.800 4.200 65.100 ;
        RECT 5.400 60.800 5.800 65.100 ;
        RECT 7.000 60.800 7.400 65.100 ;
        RECT 7.800 60.800 8.200 65.100 ;
        RECT 9.400 60.800 9.800 65.100 ;
        RECT 11.000 60.800 11.400 65.100 ;
        RECT 12.600 60.800 13.000 65.100 ;
        RECT 14.200 60.800 14.600 65.100 ;
        RECT 15.800 60.800 16.200 65.000 ;
        RECT 18.600 60.800 19.000 63.100 ;
        RECT 20.200 60.800 20.600 63.100 ;
        RECT 23.000 60.800 23.400 65.100 ;
        RECT 25.400 60.800 25.800 64.500 ;
        RECT 29.400 60.800 29.800 65.100 ;
        RECT 30.800 60.800 31.200 65.100 ;
        RECT 33.400 60.800 33.800 64.900 ;
        RECT 35.800 60.800 36.200 64.900 ;
        RECT 38.400 60.800 38.800 65.100 ;
        RECT 40.600 60.800 41.000 63.100 ;
        RECT 42.000 60.800 42.400 65.100 ;
        RECT 44.600 60.800 45.000 64.900 ;
        RECT 46.800 60.800 47.200 65.100 ;
        RECT 49.400 60.800 49.800 64.900 ;
        RECT 51.800 60.800 52.200 64.500 ;
        RECT 57.400 60.800 57.800 64.900 ;
        RECT 60.000 60.800 60.400 65.100 ;
        RECT 62.000 60.800 62.400 65.100 ;
        RECT 64.600 60.800 65.000 64.900 ;
        RECT 67.000 60.800 67.400 64.900 ;
        RECT 69.600 60.800 70.000 65.100 ;
        RECT 71.800 60.800 72.200 64.900 ;
        RECT 74.400 60.800 74.800 65.100 ;
        RECT 76.600 60.800 77.000 64.500 ;
        RECT 80.600 60.800 81.000 65.000 ;
        RECT 83.400 60.800 83.800 63.100 ;
        RECT 85.000 60.800 85.400 63.100 ;
        RECT 87.800 60.800 88.200 65.100 ;
        RECT 90.200 60.800 90.600 64.900 ;
        RECT 92.800 60.800 93.200 65.100 ;
        RECT 95.000 60.800 95.400 63.100 ;
        RECT 98.200 60.800 98.600 64.500 ;
        RECT 100.400 60.800 100.800 65.100 ;
        RECT 103.000 60.800 103.400 64.900 ;
        RECT 107.000 60.800 107.400 64.900 ;
        RECT 109.600 60.800 110.000 65.100 ;
        RECT 111.000 60.800 111.400 63.100 ;
        RECT 112.600 60.800 113.000 63.100 ;
        RECT 114.200 60.800 114.600 64.900 ;
        RECT 116.800 60.800 117.200 65.100 ;
        RECT 119.000 60.800 119.400 64.900 ;
        RECT 121.600 60.800 122.000 65.100 ;
        RECT 123.000 60.800 123.400 63.100 ;
        RECT 124.600 60.800 125.000 63.100 ;
        RECT 127.800 60.800 128.200 64.500 ;
        RECT 131.800 60.800 132.200 64.500 ;
        RECT 134.000 60.800 134.400 65.100 ;
        RECT 136.600 60.800 137.000 64.900 ;
        RECT 139.000 60.800 139.400 64.500 ;
        RECT 141.400 60.800 141.800 65.100 ;
        RECT 143.000 60.800 143.400 65.100 ;
        RECT 144.600 60.800 145.000 65.100 ;
        RECT 146.200 60.800 146.600 65.100 ;
        RECT 147.800 60.800 148.200 65.100 ;
        RECT 148.600 60.800 149.000 65.100 ;
        RECT 150.700 60.800 151.100 63.100 ;
        RECT 152.400 60.800 152.800 65.100 ;
        RECT 155.000 60.800 155.400 64.900 ;
        RECT 158.200 60.800 158.600 63.100 ;
        RECT 159.800 60.800 160.200 63.100 ;
        RECT 163.000 60.800 163.400 64.500 ;
        RECT 164.600 60.800 165.000 63.100 ;
        RECT 166.200 60.800 166.600 63.100 ;
        RECT 167.800 60.800 168.200 64.500 ;
        RECT 171.800 60.800 172.200 65.100 ;
        RECT 174.600 60.800 175.000 63.100 ;
        RECT 176.200 60.800 176.600 63.100 ;
        RECT 179.000 60.800 179.400 65.000 ;
        RECT 180.600 60.800 181.000 63.100 ;
        RECT 182.200 60.800 182.600 63.100 ;
        RECT 183.300 60.800 183.700 63.100 ;
        RECT 185.400 60.800 185.800 65.100 ;
        RECT 186.200 60.800 186.600 65.100 ;
        RECT 187.800 60.800 188.200 64.500 ;
        RECT 189.400 60.800 189.800 65.100 ;
        RECT 191.000 60.800 191.400 65.100 ;
        RECT 192.600 60.800 193.000 65.100 ;
        RECT 194.200 60.800 194.600 65.100 ;
        RECT 195.800 60.800 196.200 65.100 ;
        RECT 197.400 60.800 197.800 64.500 ;
        RECT 200.600 60.800 201.000 63.100 ;
        RECT 202.200 60.800 202.600 63.100 ;
        RECT 205.400 60.800 205.800 64.500 ;
        RECT 209.400 60.800 209.800 64.500 ;
        RECT 212.600 60.800 213.000 63.100 ;
        RECT 214.200 60.800 214.600 63.100 ;
        RECT 217.400 60.800 217.800 64.500 ;
        RECT 219.600 60.800 220.000 65.100 ;
        RECT 222.200 60.800 222.600 64.900 ;
        RECT 224.600 60.800 225.000 64.900 ;
        RECT 227.200 60.800 227.600 65.100 ;
        RECT 229.400 60.800 229.800 65.000 ;
        RECT 232.200 60.800 232.600 63.100 ;
        RECT 233.800 60.800 234.200 63.100 ;
        RECT 236.600 60.800 237.000 65.100 ;
        RECT 238.800 60.800 239.200 65.100 ;
        RECT 241.400 60.800 241.800 64.900 ;
        RECT 243.800 60.800 244.200 64.900 ;
        RECT 246.400 60.800 246.800 65.100 ;
        RECT 248.600 60.800 249.000 64.900 ;
        RECT 251.200 60.800 251.600 65.100 ;
        RECT 252.900 60.800 253.300 63.100 ;
        RECT 255.000 60.800 255.400 65.100 ;
        RECT 256.600 60.800 257.000 65.100 ;
        RECT 259.400 60.800 259.800 63.100 ;
        RECT 261.000 60.800 261.400 63.100 ;
        RECT 263.800 60.800 264.200 65.000 ;
        RECT 0.200 60.200 265.400 60.800 ;
        RECT 0.600 55.900 1.000 60.200 ;
        RECT 2.200 55.900 2.600 60.200 ;
        RECT 3.800 55.900 4.200 60.200 ;
        RECT 5.400 55.900 5.800 60.200 ;
        RECT 7.000 55.900 7.400 60.200 ;
        RECT 7.800 55.900 8.200 60.200 ;
        RECT 9.400 55.900 9.800 60.200 ;
        RECT 11.000 55.900 11.400 60.200 ;
        RECT 12.600 55.900 13.000 60.200 ;
        RECT 14.200 55.900 14.600 60.200 ;
        RECT 15.800 56.100 16.200 60.200 ;
        RECT 18.400 55.900 18.800 60.200 ;
        RECT 20.600 56.000 21.000 60.200 ;
        RECT 23.400 57.900 23.800 60.200 ;
        RECT 25.000 57.900 25.400 60.200 ;
        RECT 27.800 55.900 28.200 60.200 ;
        RECT 30.200 56.100 30.600 60.200 ;
        RECT 32.800 55.900 33.200 60.200 ;
        RECT 35.000 57.900 35.400 60.200 ;
        RECT 35.800 57.900 36.200 60.200 ;
        RECT 38.000 55.900 38.400 60.200 ;
        RECT 40.600 56.100 41.000 60.200 ;
        RECT 43.000 56.100 43.400 60.200 ;
        RECT 45.600 55.900 46.000 60.200 ;
        RECT 47.800 56.000 48.200 60.200 ;
        RECT 50.600 57.900 51.000 60.200 ;
        RECT 52.200 57.900 52.600 60.200 ;
        RECT 55.000 55.900 55.400 60.200 ;
        RECT 59.000 56.500 59.400 60.200 ;
        RECT 61.400 55.900 61.800 60.200 ;
        RECT 64.400 55.900 64.800 60.200 ;
        RECT 67.000 56.100 67.400 60.200 ;
        RECT 68.600 55.900 69.000 60.200 ;
        RECT 70.700 57.900 71.100 60.200 ;
        RECT 71.800 57.900 72.200 60.200 ;
        RECT 73.400 57.900 73.800 60.200 ;
        RECT 75.000 55.900 75.400 60.200 ;
        RECT 77.800 57.900 78.200 60.200 ;
        RECT 79.400 57.900 79.800 60.200 ;
        RECT 82.200 56.000 82.600 60.200 ;
        RECT 83.800 55.900 84.200 60.200 ;
        RECT 85.900 57.900 86.300 60.200 ;
        RECT 87.000 57.900 87.400 60.200 ;
        RECT 88.600 57.900 89.000 60.200 ;
        RECT 90.200 56.100 90.600 60.200 ;
        RECT 92.800 55.900 93.200 60.200 ;
        RECT 95.000 56.100 95.400 60.200 ;
        RECT 97.600 55.900 98.000 60.200 ;
        RECT 99.800 56.000 100.200 60.200 ;
        RECT 102.600 57.900 103.000 60.200 ;
        RECT 104.200 57.900 104.600 60.200 ;
        RECT 107.000 55.900 107.400 60.200 ;
        RECT 110.500 57.900 110.900 60.200 ;
        RECT 112.600 55.900 113.000 60.200 ;
        RECT 113.400 55.900 113.800 60.200 ;
        RECT 117.400 56.500 117.800 60.200 ;
        RECT 119.800 56.000 120.200 60.200 ;
        RECT 122.600 57.900 123.000 60.200 ;
        RECT 124.200 57.900 124.600 60.200 ;
        RECT 127.000 55.900 127.400 60.200 ;
        RECT 128.600 57.900 129.000 60.200 ;
        RECT 130.200 57.900 130.600 60.200 ;
        RECT 131.300 57.900 131.700 60.200 ;
        RECT 133.400 55.900 133.800 60.200 ;
        RECT 134.800 55.900 135.200 60.200 ;
        RECT 137.400 56.100 137.800 60.200 ;
        RECT 139.800 56.100 140.200 60.200 ;
        RECT 142.400 55.900 142.800 60.200 ;
        RECT 144.600 56.100 145.000 60.200 ;
        RECT 147.200 55.900 147.600 60.200 ;
        RECT 149.400 56.000 149.800 60.200 ;
        RECT 152.200 57.900 152.600 60.200 ;
        RECT 153.800 57.900 154.200 60.200 ;
        RECT 156.600 55.900 157.000 60.200 ;
        RECT 159.800 55.900 160.200 60.200 ;
        RECT 161.900 57.900 162.300 60.200 ;
        RECT 163.000 57.900 163.400 60.200 ;
        RECT 164.600 57.900 165.000 60.200 ;
        RECT 166.000 55.900 166.400 60.200 ;
        RECT 168.600 56.100 169.000 60.200 ;
        RECT 170.800 55.900 171.200 60.200 ;
        RECT 173.400 56.100 173.800 60.200 ;
        RECT 175.000 55.900 175.400 60.200 ;
        RECT 179.000 56.500 179.400 60.200 ;
        RECT 181.400 55.900 181.800 60.200 ;
        RECT 184.200 57.900 184.600 60.200 ;
        RECT 185.800 57.900 186.200 60.200 ;
        RECT 188.600 56.000 189.000 60.200 ;
        RECT 191.000 56.100 191.400 60.200 ;
        RECT 193.600 55.900 194.000 60.200 ;
        RECT 195.800 57.900 196.200 60.200 ;
        RECT 197.400 56.100 197.800 60.200 ;
        RECT 200.000 55.900 200.400 60.200 ;
        RECT 202.200 56.100 202.600 60.200 ;
        RECT 204.800 55.900 205.200 60.200 ;
        RECT 206.200 55.900 206.600 60.200 ;
        RECT 208.300 57.900 208.700 60.200 ;
        RECT 211.800 56.000 212.200 60.200 ;
        RECT 214.600 57.900 215.000 60.200 ;
        RECT 216.200 57.900 216.600 60.200 ;
        RECT 219.000 55.900 219.400 60.200 ;
        RECT 221.200 55.900 221.600 60.200 ;
        RECT 223.800 56.100 224.200 60.200 ;
        RECT 226.200 56.100 226.600 60.200 ;
        RECT 228.800 55.900 229.200 60.200 ;
        RECT 231.000 56.100 231.400 60.200 ;
        RECT 233.600 55.900 234.000 60.200 ;
        RECT 235.000 55.900 235.400 60.200 ;
        RECT 237.100 57.900 237.500 60.200 ;
        RECT 239.000 56.000 239.400 60.200 ;
        RECT 241.800 57.900 242.200 60.200 ;
        RECT 243.400 57.900 243.800 60.200 ;
        RECT 246.200 55.900 246.600 60.200 ;
        RECT 247.800 55.900 248.200 60.200 ;
        RECT 249.900 57.900 250.300 60.200 ;
        RECT 251.000 57.900 251.400 60.200 ;
        RECT 252.600 57.900 253.000 60.200 ;
        RECT 254.200 56.100 254.600 60.200 ;
        RECT 256.800 55.900 257.200 60.200 ;
        RECT 258.200 57.900 258.600 60.200 ;
        RECT 259.800 57.900 260.200 60.200 ;
        RECT 260.600 55.900 261.000 60.200 ;
        RECT 262.700 57.900 263.100 60.200 ;
        RECT 1.400 40.800 1.800 45.000 ;
        RECT 4.200 40.800 4.600 43.100 ;
        RECT 5.800 40.800 6.200 43.100 ;
        RECT 8.600 40.800 9.000 45.100 ;
        RECT 10.200 40.800 10.600 43.100 ;
        RECT 12.400 40.800 12.800 45.100 ;
        RECT 15.000 40.800 15.400 44.900 ;
        RECT 17.400 40.800 17.800 45.100 ;
        RECT 20.200 40.800 20.600 43.100 ;
        RECT 21.800 40.800 22.200 43.100 ;
        RECT 24.600 40.800 25.000 45.000 ;
        RECT 26.200 40.800 26.600 43.100 ;
        RECT 28.400 40.800 28.800 45.100 ;
        RECT 31.000 40.800 31.400 44.900 ;
        RECT 33.400 40.800 33.800 45.100 ;
        RECT 36.200 40.800 36.600 43.100 ;
        RECT 37.800 40.800 38.200 43.100 ;
        RECT 40.600 40.800 41.000 45.000 ;
        RECT 43.000 40.800 43.400 45.100 ;
        RECT 45.800 40.800 46.200 43.100 ;
        RECT 47.400 40.800 47.800 43.100 ;
        RECT 50.200 40.800 50.600 45.000 ;
        RECT 51.800 40.800 52.200 43.100 ;
        RECT 53.400 40.800 53.800 43.100 ;
        RECT 56.100 40.800 56.500 43.100 ;
        RECT 58.200 40.800 58.600 45.100 ;
        RECT 59.000 40.800 59.400 45.100 ;
        RECT 60.600 40.800 61.000 44.500 ;
        RECT 63.000 40.800 63.400 45.100 ;
        RECT 65.800 40.800 66.200 43.100 ;
        RECT 67.400 40.800 67.800 43.100 ;
        RECT 70.200 40.800 70.600 45.000 ;
        RECT 72.600 40.800 73.000 45.100 ;
        RECT 75.400 40.800 75.800 43.100 ;
        RECT 77.000 40.800 77.400 43.100 ;
        RECT 79.800 40.800 80.200 45.000 ;
        RECT 81.400 40.800 81.800 45.100 ;
        RECT 83.500 40.800 83.900 43.100 ;
        RECT 84.600 40.800 85.000 43.100 ;
        RECT 86.200 40.800 86.600 43.100 ;
        RECT 87.800 40.800 88.200 45.000 ;
        RECT 90.600 40.800 91.000 43.100 ;
        RECT 92.200 40.800 92.600 43.100 ;
        RECT 95.000 40.800 95.400 45.100 ;
        RECT 96.600 40.800 97.000 43.100 ;
        RECT 98.200 40.800 98.600 43.100 ;
        RECT 99.300 40.800 99.700 43.100 ;
        RECT 101.400 40.800 101.800 45.100 ;
        RECT 104.600 40.800 105.000 45.100 ;
        RECT 107.400 40.800 107.800 43.100 ;
        RECT 109.000 40.800 109.400 43.100 ;
        RECT 111.800 40.800 112.200 45.000 ;
        RECT 114.200 40.800 114.600 45.000 ;
        RECT 117.000 40.800 117.400 43.100 ;
        RECT 118.600 40.800 119.000 43.100 ;
        RECT 121.400 40.800 121.800 45.100 ;
        RECT 123.300 40.800 123.700 43.100 ;
        RECT 125.400 40.800 125.800 45.100 ;
        RECT 126.500 40.800 126.900 43.100 ;
        RECT 128.600 40.800 129.000 45.100 ;
        RECT 130.200 40.800 130.600 45.000 ;
        RECT 133.000 40.800 133.400 43.100 ;
        RECT 134.600 40.800 135.000 43.100 ;
        RECT 137.400 40.800 137.800 45.100 ;
        RECT 139.000 40.800 139.400 45.100 ;
        RECT 141.100 40.800 141.500 43.100 ;
        RECT 142.500 40.800 142.900 43.100 ;
        RECT 144.600 40.800 145.000 45.100 ;
        RECT 146.200 40.800 146.600 44.900 ;
        RECT 148.800 40.800 149.200 45.100 ;
        RECT 151.000 40.800 151.400 43.100 ;
        RECT 151.800 40.800 152.200 43.100 ;
        RECT 153.400 40.800 153.800 43.100 ;
        RECT 154.500 40.800 154.900 43.100 ;
        RECT 156.600 40.800 157.000 45.100 ;
        RECT 159.800 40.800 160.200 45.100 ;
        RECT 162.600 40.800 163.000 43.100 ;
        RECT 164.200 40.800 164.600 43.100 ;
        RECT 167.000 40.800 167.400 45.000 ;
        RECT 169.400 40.800 169.800 44.500 ;
        RECT 171.000 40.800 171.400 45.100 ;
        RECT 171.800 40.800 172.200 45.100 ;
        RECT 173.900 40.800 174.300 43.100 ;
        RECT 175.000 40.800 175.400 43.100 ;
        RECT 176.600 40.800 177.000 43.100 ;
        RECT 178.200 40.800 178.600 45.100 ;
        RECT 181.000 40.800 181.400 43.100 ;
        RECT 182.600 40.800 183.000 43.100 ;
        RECT 185.400 40.800 185.800 45.000 ;
        RECT 187.800 40.800 188.200 45.000 ;
        RECT 190.600 40.800 191.000 43.100 ;
        RECT 192.200 40.800 192.600 43.100 ;
        RECT 195.000 40.800 195.400 45.100 ;
        RECT 197.400 40.800 197.800 45.000 ;
        RECT 200.200 40.800 200.600 43.100 ;
        RECT 201.800 40.800 202.200 43.100 ;
        RECT 204.600 40.800 205.000 45.100 ;
        RECT 206.200 40.800 206.600 45.100 ;
        RECT 211.800 40.800 212.200 44.500 ;
        RECT 214.200 40.800 214.600 44.900 ;
        RECT 216.800 40.800 217.200 45.100 ;
        RECT 218.200 40.800 218.600 43.100 ;
        RECT 219.800 40.800 220.200 43.100 ;
        RECT 221.400 40.800 221.800 44.900 ;
        RECT 224.000 40.800 224.400 45.100 ;
        RECT 226.200 40.800 226.600 44.900 ;
        RECT 228.800 40.800 229.200 45.100 ;
        RECT 230.200 40.800 230.600 45.100 ;
        RECT 232.300 40.800 232.700 43.100 ;
        RECT 233.400 40.800 233.800 43.100 ;
        RECT 235.000 40.800 235.400 43.100 ;
        RECT 235.800 40.800 236.200 43.100 ;
        RECT 237.400 40.800 237.800 43.100 ;
        RECT 239.000 40.800 239.400 45.100 ;
        RECT 241.800 40.800 242.200 43.100 ;
        RECT 243.400 40.800 243.800 43.100 ;
        RECT 246.200 40.800 246.600 45.000 ;
        RECT 249.400 40.800 249.800 45.100 ;
        RECT 251.000 40.800 251.400 45.000 ;
        RECT 253.800 40.800 254.200 43.100 ;
        RECT 255.400 40.800 255.800 43.100 ;
        RECT 258.200 40.800 258.600 45.100 ;
        RECT 259.800 40.800 260.200 43.100 ;
        RECT 261.400 40.800 261.800 43.100 ;
        RECT 262.200 40.800 262.600 45.100 ;
        RECT 264.300 40.800 264.700 43.100 ;
        RECT 0.200 40.200 265.400 40.800 ;
        RECT 1.400 36.500 1.800 40.200 ;
        RECT 5.400 35.900 5.800 40.200 ;
        RECT 7.000 36.100 7.400 40.200 ;
        RECT 9.600 35.900 10.000 40.200 ;
        RECT 11.000 37.900 11.400 40.200 ;
        RECT 13.400 35.900 13.800 40.200 ;
        RECT 16.200 37.900 16.600 40.200 ;
        RECT 17.800 37.900 18.200 40.200 ;
        RECT 20.600 36.000 21.000 40.200 ;
        RECT 22.800 35.900 23.200 40.200 ;
        RECT 25.400 36.100 25.800 40.200 ;
        RECT 27.000 35.900 27.400 40.200 ;
        RECT 29.100 37.900 29.500 40.200 ;
        RECT 30.200 37.900 30.600 40.200 ;
        RECT 31.800 37.900 32.200 40.200 ;
        RECT 32.600 35.900 33.000 40.200 ;
        RECT 34.700 37.900 35.100 40.200 ;
        RECT 35.800 37.900 36.200 40.200 ;
        RECT 37.400 37.900 37.800 40.200 ;
        RECT 39.000 36.100 39.400 40.200 ;
        RECT 41.600 35.900 42.000 40.200 ;
        RECT 44.600 35.900 45.000 40.200 ;
        RECT 46.200 36.000 46.600 40.200 ;
        RECT 49.000 37.900 49.400 40.200 ;
        RECT 50.600 37.900 51.000 40.200 ;
        RECT 53.400 35.900 53.800 40.200 ;
        RECT 57.200 35.900 57.600 40.200 ;
        RECT 59.800 36.100 60.200 40.200 ;
        RECT 61.400 37.900 61.800 40.200 ;
        RECT 63.000 37.900 63.400 40.200 ;
        RECT 64.600 36.100 65.000 40.200 ;
        RECT 67.200 35.900 67.600 40.200 ;
        RECT 68.600 35.900 69.000 40.200 ;
        RECT 70.700 37.900 71.100 40.200 ;
        RECT 71.800 37.900 72.200 40.200 ;
        RECT 73.400 37.900 73.800 40.200 ;
        RECT 75.000 36.000 75.400 40.200 ;
        RECT 77.800 37.900 78.200 40.200 ;
        RECT 79.400 37.900 79.800 40.200 ;
        RECT 82.200 35.900 82.600 40.200 ;
        RECT 84.600 36.100 85.000 40.200 ;
        RECT 87.200 35.900 87.600 40.200 ;
        RECT 89.200 35.900 89.600 40.200 ;
        RECT 91.800 36.100 92.200 40.200 ;
        RECT 94.200 36.000 94.600 40.200 ;
        RECT 97.000 37.900 97.400 40.200 ;
        RECT 98.600 37.900 99.000 40.200 ;
        RECT 101.400 35.900 101.800 40.200 ;
        RECT 103.000 37.900 103.400 40.200 ;
        RECT 106.800 35.900 107.200 40.200 ;
        RECT 109.400 36.100 109.800 40.200 ;
        RECT 111.000 35.900 111.400 40.200 ;
        RECT 112.600 35.900 113.000 40.200 ;
        RECT 114.200 35.900 114.600 40.200 ;
        RECT 115.800 35.900 116.200 40.200 ;
        RECT 117.400 35.900 117.800 40.200 ;
        RECT 118.200 35.900 118.600 40.200 ;
        RECT 119.800 35.900 120.200 40.200 ;
        RECT 121.400 35.900 121.800 40.200 ;
        RECT 123.000 35.900 123.400 40.200 ;
        RECT 124.600 35.900 125.000 40.200 ;
        RECT 126.200 36.100 126.600 40.200 ;
        RECT 128.800 35.900 129.200 40.200 ;
        RECT 131.000 36.500 131.400 40.200 ;
        RECT 132.600 35.900 133.000 40.200 ;
        RECT 134.200 36.100 134.600 40.200 ;
        RECT 136.800 35.900 137.200 40.200 ;
        RECT 138.200 35.900 138.600 40.200 ;
        RECT 142.200 36.500 142.600 40.200 ;
        RECT 144.600 36.000 145.000 40.200 ;
        RECT 147.400 37.900 147.800 40.200 ;
        RECT 149.000 37.900 149.400 40.200 ;
        RECT 151.800 35.900 152.200 40.200 ;
        RECT 154.700 35.900 155.100 40.200 ;
        RECT 159.000 36.000 159.400 40.200 ;
        RECT 161.800 37.900 162.200 40.200 ;
        RECT 163.400 37.900 163.800 40.200 ;
        RECT 166.200 35.900 166.600 40.200 ;
        RECT 168.600 36.100 169.000 40.200 ;
        RECT 171.200 35.900 171.600 40.200 ;
        RECT 172.600 35.900 173.000 40.200 ;
        RECT 176.600 36.500 177.000 40.200 ;
        RECT 179.000 36.000 179.400 40.200 ;
        RECT 181.800 37.900 182.200 40.200 ;
        RECT 183.400 37.900 183.800 40.200 ;
        RECT 186.200 35.900 186.600 40.200 ;
        RECT 188.600 36.100 189.000 40.200 ;
        RECT 191.200 35.900 191.600 40.200 ;
        RECT 193.400 37.900 193.800 40.200 ;
        RECT 195.000 36.100 195.400 40.200 ;
        RECT 197.600 35.900 198.000 40.200 ;
        RECT 199.600 35.900 200.000 40.200 ;
        RECT 202.200 36.100 202.600 40.200 ;
        RECT 204.600 36.500 205.000 40.200 ;
        RECT 208.600 35.900 209.000 40.200 ;
        RECT 211.600 35.900 212.000 40.200 ;
        RECT 214.200 36.100 214.600 40.200 ;
        RECT 216.400 35.900 216.800 40.200 ;
        RECT 219.000 36.100 219.400 40.200 ;
        RECT 221.400 36.500 221.800 40.200 ;
        RECT 223.800 35.900 224.200 40.200 ;
        RECT 227.000 36.100 227.400 40.200 ;
        RECT 229.600 35.900 230.000 40.200 ;
        RECT 231.000 37.900 231.400 40.200 ;
        RECT 232.600 37.900 233.000 40.200 ;
        RECT 233.700 37.900 234.100 40.200 ;
        RECT 235.800 35.900 236.200 40.200 ;
        RECT 237.400 35.900 237.800 40.200 ;
        RECT 240.200 37.900 240.600 40.200 ;
        RECT 241.800 37.900 242.200 40.200 ;
        RECT 244.600 36.000 245.000 40.200 ;
        RECT 246.200 35.900 246.600 40.200 ;
        RECT 248.300 37.900 248.700 40.200 ;
        RECT 249.400 37.900 249.800 40.200 ;
        RECT 251.000 37.900 251.400 40.200 ;
        RECT 252.600 35.900 253.000 40.200 ;
        RECT 255.400 37.900 255.800 40.200 ;
        RECT 257.000 37.900 257.400 40.200 ;
        RECT 259.800 36.000 260.200 40.200 ;
        RECT 261.400 35.900 261.800 40.200 ;
        RECT 263.500 37.900 263.900 40.200 ;
        RECT 1.400 20.800 1.800 25.000 ;
        RECT 4.200 20.800 4.600 23.100 ;
        RECT 5.800 20.800 6.200 23.100 ;
        RECT 8.600 20.800 9.000 25.100 ;
        RECT 10.200 20.800 10.600 25.100 ;
        RECT 11.800 20.800 12.200 25.100 ;
        RECT 13.400 20.800 13.800 25.100 ;
        RECT 15.000 20.800 15.400 25.100 ;
        RECT 16.600 20.800 17.000 25.100 ;
        RECT 18.200 20.800 18.600 24.900 ;
        RECT 20.800 20.800 21.200 25.100 ;
        RECT 22.800 20.800 23.200 25.100 ;
        RECT 25.400 20.800 25.800 24.900 ;
        RECT 27.800 20.800 28.200 25.000 ;
        RECT 30.600 20.800 31.000 23.100 ;
        RECT 32.200 20.800 32.600 23.100 ;
        RECT 35.000 20.800 35.400 25.100 ;
        RECT 37.400 20.800 37.800 25.000 ;
        RECT 40.200 20.800 40.600 23.100 ;
        RECT 41.800 20.800 42.200 23.100 ;
        RECT 44.600 20.800 45.000 25.100 ;
        RECT 47.800 20.800 48.200 24.500 ;
        RECT 50.200 20.800 50.600 25.000 ;
        RECT 53.000 20.800 53.400 23.100 ;
        RECT 54.600 20.800 55.000 23.100 ;
        RECT 57.400 20.800 57.800 25.100 ;
        RECT 60.600 20.800 61.000 25.100 ;
        RECT 62.700 20.800 63.100 23.100 ;
        RECT 64.600 20.800 65.000 24.500 ;
        RECT 66.200 20.800 66.600 25.100 ;
        RECT 67.000 20.800 67.400 25.100 ;
        RECT 69.100 20.800 69.500 23.100 ;
        RECT 70.200 20.800 70.600 23.100 ;
        RECT 71.800 20.800 72.200 23.100 ;
        RECT 73.400 20.800 73.800 25.100 ;
        RECT 76.200 20.800 76.600 23.100 ;
        RECT 77.800 20.800 78.200 23.100 ;
        RECT 80.600 20.800 81.000 25.000 ;
        RECT 82.800 20.800 83.200 25.100 ;
        RECT 85.400 20.800 85.800 24.900 ;
        RECT 87.000 20.800 87.400 23.100 ;
        RECT 89.200 20.800 89.600 25.100 ;
        RECT 91.800 20.800 92.200 24.900 ;
        RECT 94.200 20.800 94.600 24.900 ;
        RECT 96.800 20.800 97.200 25.100 ;
        RECT 98.200 20.800 98.600 25.100 ;
        RECT 99.800 20.800 100.200 24.500 ;
        RECT 101.400 20.800 101.800 25.100 ;
        RECT 103.500 20.800 103.900 23.100 ;
        RECT 104.600 20.800 105.000 23.100 ;
        RECT 106.200 20.800 106.600 23.100 ;
        RECT 109.400 20.800 109.800 25.100 ;
        RECT 112.200 20.800 112.600 23.100 ;
        RECT 113.800 20.800 114.200 23.100 ;
        RECT 116.600 20.800 117.000 25.000 ;
        RECT 119.000 20.800 119.400 24.900 ;
        RECT 121.600 20.800 122.000 25.100 ;
        RECT 123.800 20.800 124.200 24.900 ;
        RECT 126.400 20.800 126.800 25.100 ;
        RECT 128.600 20.800 129.000 23.100 ;
        RECT 130.200 20.800 130.600 25.100 ;
        RECT 133.000 20.800 133.400 23.100 ;
        RECT 134.600 20.800 135.000 23.100 ;
        RECT 137.400 20.800 137.800 25.000 ;
        RECT 139.800 20.800 140.200 25.100 ;
        RECT 142.600 20.800 143.000 23.100 ;
        RECT 144.200 20.800 144.600 23.100 ;
        RECT 147.000 20.800 147.400 25.000 ;
        RECT 148.600 20.800 149.000 25.100 ;
        RECT 150.700 20.800 151.100 23.100 ;
        RECT 151.800 20.800 152.200 23.100 ;
        RECT 153.400 20.800 153.800 23.100 ;
        RECT 156.600 20.800 157.000 25.000 ;
        RECT 159.400 20.800 159.800 23.100 ;
        RECT 161.000 20.800 161.400 23.100 ;
        RECT 163.800 20.800 164.200 25.100 ;
        RECT 165.400 20.800 165.800 25.100 ;
        RECT 167.500 20.800 167.900 23.100 ;
        RECT 168.600 20.800 169.000 23.100 ;
        RECT 170.200 20.800 170.600 23.100 ;
        RECT 171.800 20.800 172.200 25.100 ;
        RECT 174.600 20.800 175.000 23.100 ;
        RECT 176.200 20.800 176.600 23.100 ;
        RECT 179.000 20.800 179.400 25.000 ;
        RECT 180.600 20.800 181.000 25.100 ;
        RECT 182.200 20.800 182.600 24.500 ;
        RECT 184.600 20.800 185.000 24.900 ;
        RECT 187.200 20.800 187.600 25.100 ;
        RECT 189.400 20.800 189.800 23.100 ;
        RECT 191.000 20.800 191.400 25.100 ;
        RECT 193.800 20.800 194.200 23.100 ;
        RECT 195.400 20.800 195.800 23.100 ;
        RECT 198.200 20.800 198.600 25.000 ;
        RECT 199.800 20.800 200.200 25.100 ;
        RECT 201.900 20.800 202.300 23.100 ;
        RECT 203.300 20.800 203.700 23.100 ;
        RECT 205.400 20.800 205.800 25.100 ;
        RECT 208.600 20.800 209.000 25.000 ;
        RECT 211.400 20.800 211.800 23.100 ;
        RECT 213.000 20.800 213.400 23.100 ;
        RECT 215.800 20.800 216.200 25.100 ;
        RECT 218.200 20.800 218.600 24.900 ;
        RECT 220.800 20.800 221.200 25.100 ;
        RECT 223.000 20.800 223.400 25.100 ;
        RECT 225.800 20.800 226.200 23.100 ;
        RECT 227.400 20.800 227.800 23.100 ;
        RECT 230.200 20.800 230.600 25.000 ;
        RECT 232.600 20.800 233.000 23.100 ;
        RECT 234.200 20.800 234.600 25.100 ;
        RECT 237.000 20.800 237.400 23.100 ;
        RECT 238.600 20.800 239.000 23.100 ;
        RECT 241.400 20.800 241.800 25.000 ;
        RECT 243.000 20.800 243.400 23.100 ;
        RECT 244.600 20.800 245.000 23.100 ;
        RECT 245.700 20.800 246.100 23.100 ;
        RECT 247.800 20.800 248.200 25.100 ;
        RECT 249.400 20.800 249.800 24.900 ;
        RECT 252.000 20.800 252.400 25.100 ;
        RECT 254.200 20.800 254.600 25.100 ;
        RECT 257.000 20.800 257.400 23.100 ;
        RECT 258.600 20.800 259.000 23.100 ;
        RECT 261.400 20.800 261.800 25.000 ;
        RECT 0.200 20.200 265.400 20.800 ;
        RECT 1.400 15.900 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 16.000 9.000 20.200 ;
        RECT 10.500 17.900 10.900 20.200 ;
        RECT 12.600 15.900 13.000 20.200 ;
        RECT 13.400 15.900 13.800 20.200 ;
        RECT 15.500 17.900 15.900 20.200 ;
        RECT 16.600 17.900 17.000 20.200 ;
        RECT 18.200 17.900 18.600 20.200 ;
        RECT 19.800 16.100 20.200 20.200 ;
        RECT 22.400 15.900 22.800 20.200 ;
        RECT 24.600 15.900 25.000 20.200 ;
        RECT 27.400 17.900 27.800 20.200 ;
        RECT 29.000 17.900 29.400 20.200 ;
        RECT 31.800 16.000 32.200 20.200 ;
        RECT 33.400 15.900 33.800 20.200 ;
        RECT 37.400 16.500 37.800 20.200 ;
        RECT 39.000 15.900 39.400 20.200 ;
        RECT 40.600 16.500 41.000 20.200 ;
        RECT 42.200 15.900 42.600 20.200 ;
        RECT 43.800 15.900 44.200 20.200 ;
        RECT 45.400 15.900 45.800 20.200 ;
        RECT 47.000 15.900 47.400 20.200 ;
        RECT 48.600 15.900 49.000 20.200 ;
        RECT 49.400 15.900 49.800 20.200 ;
        RECT 51.000 15.900 51.400 20.200 ;
        RECT 52.600 15.900 53.000 20.200 ;
        RECT 55.000 15.900 55.400 20.200 ;
        RECT 56.600 16.500 57.000 20.200 ;
        RECT 58.200 15.900 58.600 20.200 ;
        RECT 60.300 17.900 60.700 20.200 ;
        RECT 61.400 17.900 61.800 20.200 ;
        RECT 63.000 17.900 63.400 20.200 ;
        RECT 64.600 16.000 65.000 20.200 ;
        RECT 67.400 17.900 67.800 20.200 ;
        RECT 69.000 17.900 69.400 20.200 ;
        RECT 71.800 15.900 72.200 20.200 ;
        RECT 74.200 16.100 74.600 20.200 ;
        RECT 76.800 15.900 77.200 20.200 ;
        RECT 79.000 16.000 79.400 20.200 ;
        RECT 81.800 17.900 82.200 20.200 ;
        RECT 83.400 17.900 83.800 20.200 ;
        RECT 86.200 15.900 86.600 20.200 ;
        RECT 87.800 17.900 88.200 20.200 ;
        RECT 90.000 15.900 90.400 20.200 ;
        RECT 92.600 16.100 93.000 20.200 ;
        RECT 95.000 15.900 95.400 20.200 ;
        RECT 97.800 17.900 98.200 20.200 ;
        RECT 99.400 17.900 99.800 20.200 ;
        RECT 102.200 16.000 102.600 20.200 ;
        RECT 103.800 15.900 104.200 20.200 ;
        RECT 105.400 16.500 105.800 20.200 ;
        RECT 109.400 16.500 109.800 20.200 ;
        RECT 113.400 15.900 113.800 20.200 ;
        RECT 114.800 15.900 115.200 20.200 ;
        RECT 117.400 16.100 117.800 20.200 ;
        RECT 119.600 15.900 120.000 20.200 ;
        RECT 122.200 16.100 122.600 20.200 ;
        RECT 124.600 15.900 125.000 20.200 ;
        RECT 127.400 17.900 127.800 20.200 ;
        RECT 129.000 17.900 129.400 20.200 ;
        RECT 131.800 16.000 132.200 20.200 ;
        RECT 133.400 15.900 133.800 20.200 ;
        RECT 135.000 15.900 135.400 20.200 ;
        RECT 136.600 15.900 137.000 20.200 ;
        RECT 138.200 15.900 138.600 20.200 ;
        RECT 139.800 15.900 140.200 20.200 ;
        RECT 140.600 15.900 141.000 20.200 ;
        RECT 142.200 15.900 142.600 20.200 ;
        RECT 143.800 15.900 144.200 20.200 ;
        RECT 145.400 15.900 145.800 20.200 ;
        RECT 147.000 15.900 147.400 20.200 ;
        RECT 148.600 16.000 149.000 20.200 ;
        RECT 151.400 17.900 151.800 20.200 ;
        RECT 153.000 17.900 153.400 20.200 ;
        RECT 155.800 15.900 156.200 20.200 ;
        RECT 159.800 16.100 160.200 20.200 ;
        RECT 162.400 15.900 162.800 20.200 ;
        RECT 164.600 17.900 165.000 20.200 ;
        RECT 166.200 16.100 166.600 20.200 ;
        RECT 168.800 15.900 169.200 20.200 ;
        RECT 170.200 15.900 170.600 20.200 ;
        RECT 171.800 15.900 172.200 20.200 ;
        RECT 173.400 15.900 173.800 20.200 ;
        RECT 174.200 15.900 174.600 20.200 ;
        RECT 176.300 17.900 176.700 20.200 ;
        RECT 177.400 17.900 177.800 20.200 ;
        RECT 179.000 17.900 179.400 20.200 ;
        RECT 180.400 15.900 180.800 20.200 ;
        RECT 183.000 16.100 183.400 20.200 ;
        RECT 185.400 16.000 185.800 20.200 ;
        RECT 188.200 17.900 188.600 20.200 ;
        RECT 189.800 17.900 190.200 20.200 ;
        RECT 192.600 15.900 193.000 20.200 ;
        RECT 195.000 16.500 195.400 20.200 ;
        RECT 196.600 15.900 197.000 20.200 ;
        RECT 197.400 15.900 197.800 20.200 ;
        RECT 199.000 15.900 199.400 20.200 ;
        RECT 200.600 15.900 201.000 20.200 ;
        RECT 202.200 15.900 202.600 20.200 ;
        RECT 203.800 15.900 204.200 20.200 ;
        RECT 204.600 15.900 205.000 20.200 ;
        RECT 206.700 17.900 207.100 20.200 ;
        RECT 209.700 17.900 210.100 20.200 ;
        RECT 211.800 15.900 212.200 20.200 ;
        RECT 213.400 15.900 213.800 20.200 ;
        RECT 216.200 17.900 216.600 20.200 ;
        RECT 217.800 17.900 218.200 20.200 ;
        RECT 220.600 16.000 221.000 20.200 ;
        RECT 223.000 16.500 223.400 20.200 ;
        RECT 224.600 15.900 225.000 20.200 ;
        RECT 225.400 17.900 225.800 20.200 ;
        RECT 227.000 17.900 227.400 20.200 ;
        RECT 228.600 16.100 229.000 20.200 ;
        RECT 231.200 15.900 231.600 20.200 ;
        RECT 233.400 15.900 233.800 20.200 ;
        RECT 236.200 17.900 236.600 20.200 ;
        RECT 237.800 17.900 238.200 20.200 ;
        RECT 240.600 16.000 241.000 20.200 ;
        RECT 242.200 15.900 242.600 20.200 ;
        RECT 243.800 15.900 244.200 20.200 ;
        RECT 245.400 15.900 245.800 20.200 ;
        RECT 247.000 15.900 247.400 20.200 ;
        RECT 248.600 15.900 249.000 20.200 ;
        RECT 249.400 15.900 249.800 20.200 ;
        RECT 251.500 17.900 251.900 20.200 ;
        RECT 252.600 17.900 253.000 20.200 ;
        RECT 254.200 17.900 254.600 20.200 ;
        RECT 255.800 15.900 256.200 20.200 ;
        RECT 258.600 17.900 259.000 20.200 ;
        RECT 260.200 17.900 260.600 20.200 ;
        RECT 263.000 16.000 263.400 20.200 ;
        RECT 0.600 0.800 1.000 5.100 ;
        RECT 2.200 0.800 2.600 5.100 ;
        RECT 3.800 0.800 4.200 5.100 ;
        RECT 5.400 0.800 5.800 5.100 ;
        RECT 7.000 0.800 7.400 5.100 ;
        RECT 7.800 0.800 8.200 3.100 ;
        RECT 9.400 0.800 9.800 3.100 ;
        RECT 11.000 0.800 11.400 5.000 ;
        RECT 13.800 0.800 14.200 3.100 ;
        RECT 15.400 0.800 15.800 3.100 ;
        RECT 18.200 0.800 18.600 5.100 ;
        RECT 20.600 0.800 21.000 5.100 ;
        RECT 23.400 0.800 23.800 3.100 ;
        RECT 25.000 0.800 25.400 3.100 ;
        RECT 27.800 0.800 28.200 5.000 ;
        RECT 29.400 0.800 29.800 3.100 ;
        RECT 31.000 0.800 31.400 3.100 ;
        RECT 32.100 0.800 32.500 3.100 ;
        RECT 34.200 0.800 34.600 5.100 ;
        RECT 35.000 0.800 35.400 5.100 ;
        RECT 36.600 0.800 37.000 5.100 ;
        RECT 38.200 0.800 38.600 5.100 ;
        RECT 39.800 0.800 40.200 5.100 ;
        RECT 41.400 0.800 41.800 5.100 ;
        RECT 42.200 0.800 42.600 5.100 ;
        RECT 43.800 0.800 44.200 5.100 ;
        RECT 45.400 0.800 45.800 5.100 ;
        RECT 47.000 0.800 47.400 5.100 ;
        RECT 48.600 0.800 49.000 5.100 ;
        RECT 49.400 0.800 49.800 5.100 ;
        RECT 51.000 0.800 51.400 5.100 ;
        RECT 52.600 0.800 53.000 5.100 ;
        RECT 54.200 0.800 54.600 5.100 ;
        RECT 55.800 0.800 56.200 5.100 ;
        RECT 58.200 0.800 58.600 5.100 ;
        RECT 59.800 0.800 60.200 5.100 ;
        RECT 61.400 0.800 61.800 5.100 ;
        RECT 63.000 0.800 63.400 5.100 ;
        RECT 64.600 0.800 65.000 5.100 ;
        RECT 66.200 0.800 66.600 4.900 ;
        RECT 68.800 0.800 69.200 5.100 ;
        RECT 71.000 0.800 71.400 3.100 ;
        RECT 72.600 0.800 73.000 5.000 ;
        RECT 75.400 0.800 75.800 3.100 ;
        RECT 77.000 0.800 77.400 3.100 ;
        RECT 79.800 0.800 80.200 5.100 ;
        RECT 82.200 0.800 82.600 5.100 ;
        RECT 85.000 0.800 85.400 3.100 ;
        RECT 86.600 0.800 87.000 3.100 ;
        RECT 89.400 0.800 89.800 5.000 ;
        RECT 91.000 0.800 91.400 3.100 ;
        RECT 92.600 0.800 93.000 3.100 ;
        RECT 93.700 0.800 94.100 3.100 ;
        RECT 95.800 0.800 96.200 5.100 ;
        RECT 97.400 0.800 97.800 5.000 ;
        RECT 100.200 0.800 100.600 3.100 ;
        RECT 101.800 0.800 102.200 3.100 ;
        RECT 104.600 0.800 105.000 5.100 ;
        RECT 107.800 0.800 108.200 3.100 ;
        RECT 110.000 0.800 110.400 5.100 ;
        RECT 112.600 0.800 113.000 4.900 ;
        RECT 114.200 0.800 114.600 5.100 ;
        RECT 116.300 0.800 116.700 3.100 ;
        RECT 117.400 0.800 117.800 3.100 ;
        RECT 119.000 0.800 119.400 3.100 ;
        RECT 120.600 0.800 121.000 5.100 ;
        RECT 123.400 0.800 123.800 3.100 ;
        RECT 125.000 0.800 125.400 3.100 ;
        RECT 127.800 0.800 128.200 5.000 ;
        RECT 129.400 0.800 129.800 3.100 ;
        RECT 131.000 0.800 131.400 3.100 ;
        RECT 132.100 0.800 132.500 3.100 ;
        RECT 134.200 0.800 134.600 5.100 ;
        RECT 135.800 0.800 136.200 5.100 ;
        RECT 138.600 0.800 139.000 3.100 ;
        RECT 140.200 0.800 140.600 3.100 ;
        RECT 143.000 0.800 143.400 5.000 ;
        RECT 144.600 0.800 145.000 5.100 ;
        RECT 146.200 0.800 146.600 5.100 ;
        RECT 147.800 0.800 148.200 5.100 ;
        RECT 149.400 0.800 149.800 5.100 ;
        RECT 151.000 0.800 151.400 5.100 ;
        RECT 151.800 0.800 152.200 5.100 ;
        RECT 153.400 0.800 153.800 4.500 ;
        RECT 157.400 0.800 157.800 5.000 ;
        RECT 160.200 0.800 160.600 3.100 ;
        RECT 161.800 0.800 162.200 3.100 ;
        RECT 164.600 0.800 165.000 5.100 ;
        RECT 166.200 0.800 166.600 3.100 ;
        RECT 168.400 0.800 168.800 5.100 ;
        RECT 171.000 0.800 171.400 4.900 ;
        RECT 172.600 0.800 173.000 5.100 ;
        RECT 174.200 0.800 174.600 5.100 ;
        RECT 175.800 0.800 176.200 5.100 ;
        RECT 177.400 0.800 177.800 4.900 ;
        RECT 180.000 0.800 180.400 5.100 ;
        RECT 182.200 0.800 182.600 3.100 ;
        RECT 183.800 0.800 184.200 5.100 ;
        RECT 186.600 0.800 187.000 3.100 ;
        RECT 188.200 0.800 188.600 3.100 ;
        RECT 191.000 0.800 191.400 5.000 ;
        RECT 193.400 0.800 193.800 5.000 ;
        RECT 196.200 0.800 196.600 3.100 ;
        RECT 197.800 0.800 198.200 3.100 ;
        RECT 200.600 0.800 201.000 5.100 ;
        RECT 203.000 0.800 203.400 5.000 ;
        RECT 205.800 0.800 206.200 3.100 ;
        RECT 207.400 0.800 207.800 3.100 ;
        RECT 210.200 0.800 210.600 5.100 ;
        RECT 213.400 0.800 213.800 5.100 ;
        RECT 215.500 0.800 215.900 3.100 ;
        RECT 216.600 0.800 217.000 3.100 ;
        RECT 218.200 0.800 218.600 3.100 ;
        RECT 219.000 0.800 219.400 5.100 ;
        RECT 220.600 0.800 221.000 5.100 ;
        RECT 222.200 0.800 222.600 5.100 ;
        RECT 223.800 0.800 224.200 5.100 ;
        RECT 225.400 0.800 225.800 5.100 ;
        RECT 226.500 0.800 226.900 3.100 ;
        RECT 228.600 0.800 229.000 5.100 ;
        RECT 230.200 0.800 230.600 5.100 ;
        RECT 233.000 0.800 233.400 3.100 ;
        RECT 234.600 0.800 235.000 3.100 ;
        RECT 237.400 0.800 237.800 5.000 ;
        RECT 239.000 0.800 239.400 5.100 ;
        RECT 240.600 0.800 241.000 5.100 ;
        RECT 242.200 0.800 242.600 5.100 ;
        RECT 243.800 0.800 244.200 5.100 ;
        RECT 245.400 0.800 245.800 5.100 ;
        RECT 246.200 0.800 246.600 5.100 ;
        RECT 247.800 0.800 248.200 5.100 ;
        RECT 249.400 0.800 249.800 5.100 ;
        RECT 251.000 0.800 251.400 5.100 ;
        RECT 252.600 0.800 253.000 5.100 ;
        RECT 254.200 0.800 254.600 5.100 ;
        RECT 257.000 0.800 257.400 3.100 ;
        RECT 258.600 0.800 259.000 3.100 ;
        RECT 261.400 0.800 261.800 5.000 ;
        RECT 0.200 0.200 265.400 0.800 ;
      LAYER via1 ;
        RECT 54.600 240.300 55.000 240.700 ;
        RECT 55.300 240.300 55.700 240.700 ;
        RECT 156.200 240.300 156.600 240.700 ;
        RECT 156.900 240.300 157.300 240.700 ;
        RECT 54.600 220.300 55.000 220.700 ;
        RECT 55.300 220.300 55.700 220.700 ;
        RECT 156.200 220.300 156.600 220.700 ;
        RECT 156.900 220.300 157.300 220.700 ;
        RECT 54.600 200.300 55.000 200.700 ;
        RECT 55.300 200.300 55.700 200.700 ;
        RECT 156.200 200.300 156.600 200.700 ;
        RECT 156.900 200.300 157.300 200.700 ;
        RECT 54.600 180.300 55.000 180.700 ;
        RECT 55.300 180.300 55.700 180.700 ;
        RECT 156.200 180.300 156.600 180.700 ;
        RECT 156.900 180.300 157.300 180.700 ;
        RECT 54.600 160.300 55.000 160.700 ;
        RECT 55.300 160.300 55.700 160.700 ;
        RECT 156.200 160.300 156.600 160.700 ;
        RECT 156.900 160.300 157.300 160.700 ;
        RECT 54.600 140.300 55.000 140.700 ;
        RECT 55.300 140.300 55.700 140.700 ;
        RECT 156.200 140.300 156.600 140.700 ;
        RECT 156.900 140.300 157.300 140.700 ;
        RECT 54.600 120.300 55.000 120.700 ;
        RECT 55.300 120.300 55.700 120.700 ;
        RECT 156.200 120.300 156.600 120.700 ;
        RECT 156.900 120.300 157.300 120.700 ;
        RECT 54.600 100.300 55.000 100.700 ;
        RECT 55.300 100.300 55.700 100.700 ;
        RECT 156.200 100.300 156.600 100.700 ;
        RECT 156.900 100.300 157.300 100.700 ;
        RECT 54.600 80.300 55.000 80.700 ;
        RECT 55.300 80.300 55.700 80.700 ;
        RECT 156.200 80.300 156.600 80.700 ;
        RECT 156.900 80.300 157.300 80.700 ;
        RECT 54.600 60.300 55.000 60.700 ;
        RECT 55.300 60.300 55.700 60.700 ;
        RECT 156.200 60.300 156.600 60.700 ;
        RECT 156.900 60.300 157.300 60.700 ;
        RECT 54.600 40.300 55.000 40.700 ;
        RECT 55.300 40.300 55.700 40.700 ;
        RECT 156.200 40.300 156.600 40.700 ;
        RECT 156.900 40.300 157.300 40.700 ;
        RECT 54.600 20.300 55.000 20.700 ;
        RECT 55.300 20.300 55.700 20.700 ;
        RECT 156.200 20.300 156.600 20.700 ;
        RECT 156.900 20.300 157.300 20.700 ;
        RECT 54.600 0.300 55.000 0.700 ;
        RECT 55.300 0.300 55.700 0.700 ;
        RECT 156.200 0.300 156.600 0.700 ;
        RECT 156.900 0.300 157.300 0.700 ;
      LAYER metal2 ;
        RECT 54.400 240.300 56.000 240.700 ;
        RECT 156.000 240.300 157.600 240.700 ;
        RECT 54.400 220.300 56.000 220.700 ;
        RECT 156.000 220.300 157.600 220.700 ;
        RECT 54.400 200.300 56.000 200.700 ;
        RECT 156.000 200.300 157.600 200.700 ;
        RECT 54.400 180.300 56.000 180.700 ;
        RECT 156.000 180.300 157.600 180.700 ;
        RECT 54.400 160.300 56.000 160.700 ;
        RECT 156.000 160.300 157.600 160.700 ;
        RECT 54.400 140.300 56.000 140.700 ;
        RECT 156.000 140.300 157.600 140.700 ;
        RECT 54.400 120.300 56.000 120.700 ;
        RECT 156.000 120.300 157.600 120.700 ;
        RECT 54.400 100.300 56.000 100.700 ;
        RECT 156.000 100.300 157.600 100.700 ;
        RECT 54.400 80.300 56.000 80.700 ;
        RECT 156.000 80.300 157.600 80.700 ;
        RECT 54.400 60.300 56.000 60.700 ;
        RECT 156.000 60.300 157.600 60.700 ;
        RECT 54.400 40.300 56.000 40.700 ;
        RECT 156.000 40.300 157.600 40.700 ;
        RECT 54.400 20.300 56.000 20.700 ;
        RECT 156.000 20.300 157.600 20.700 ;
        RECT 54.400 0.300 56.000 0.700 ;
        RECT 156.000 0.300 157.600 0.700 ;
      LAYER via2 ;
        RECT 54.600 240.300 55.000 240.700 ;
        RECT 55.300 240.300 55.700 240.700 ;
        RECT 156.200 240.300 156.600 240.700 ;
        RECT 156.900 240.300 157.300 240.700 ;
        RECT 54.600 220.300 55.000 220.700 ;
        RECT 55.300 220.300 55.700 220.700 ;
        RECT 156.200 220.300 156.600 220.700 ;
        RECT 156.900 220.300 157.300 220.700 ;
        RECT 54.600 200.300 55.000 200.700 ;
        RECT 55.300 200.300 55.700 200.700 ;
        RECT 156.200 200.300 156.600 200.700 ;
        RECT 156.900 200.300 157.300 200.700 ;
        RECT 54.600 180.300 55.000 180.700 ;
        RECT 55.300 180.300 55.700 180.700 ;
        RECT 156.200 180.300 156.600 180.700 ;
        RECT 156.900 180.300 157.300 180.700 ;
        RECT 54.600 160.300 55.000 160.700 ;
        RECT 55.300 160.300 55.700 160.700 ;
        RECT 156.200 160.300 156.600 160.700 ;
        RECT 156.900 160.300 157.300 160.700 ;
        RECT 54.600 140.300 55.000 140.700 ;
        RECT 55.300 140.300 55.700 140.700 ;
        RECT 156.200 140.300 156.600 140.700 ;
        RECT 156.900 140.300 157.300 140.700 ;
        RECT 54.600 120.300 55.000 120.700 ;
        RECT 55.300 120.300 55.700 120.700 ;
        RECT 156.200 120.300 156.600 120.700 ;
        RECT 156.900 120.300 157.300 120.700 ;
        RECT 54.600 100.300 55.000 100.700 ;
        RECT 55.300 100.300 55.700 100.700 ;
        RECT 156.200 100.300 156.600 100.700 ;
        RECT 156.900 100.300 157.300 100.700 ;
        RECT 54.600 80.300 55.000 80.700 ;
        RECT 55.300 80.300 55.700 80.700 ;
        RECT 156.200 80.300 156.600 80.700 ;
        RECT 156.900 80.300 157.300 80.700 ;
        RECT 54.600 60.300 55.000 60.700 ;
        RECT 55.300 60.300 55.700 60.700 ;
        RECT 156.200 60.300 156.600 60.700 ;
        RECT 156.900 60.300 157.300 60.700 ;
        RECT 54.600 40.300 55.000 40.700 ;
        RECT 55.300 40.300 55.700 40.700 ;
        RECT 156.200 40.300 156.600 40.700 ;
        RECT 156.900 40.300 157.300 40.700 ;
        RECT 54.600 20.300 55.000 20.700 ;
        RECT 55.300 20.300 55.700 20.700 ;
        RECT 156.200 20.300 156.600 20.700 ;
        RECT 156.900 20.300 157.300 20.700 ;
        RECT 54.600 0.300 55.000 0.700 ;
        RECT 55.300 0.300 55.700 0.700 ;
        RECT 156.200 0.300 156.600 0.700 ;
        RECT 156.900 0.300 157.300 0.700 ;
      LAYER metal3 ;
        RECT 54.400 240.300 56.000 240.700 ;
        RECT 156.000 240.300 157.600 240.700 ;
        RECT 54.400 220.300 56.000 220.700 ;
        RECT 156.000 220.300 157.600 220.700 ;
        RECT 54.400 200.300 56.000 200.700 ;
        RECT 156.000 200.300 157.600 200.700 ;
        RECT 54.400 180.300 56.000 180.700 ;
        RECT 156.000 180.300 157.600 180.700 ;
        RECT 54.400 160.300 56.000 160.700 ;
        RECT 156.000 160.300 157.600 160.700 ;
        RECT 54.400 140.300 56.000 140.700 ;
        RECT 156.000 140.300 157.600 140.700 ;
        RECT 54.400 120.300 56.000 120.700 ;
        RECT 156.000 120.300 157.600 120.700 ;
        RECT 54.400 100.300 56.000 100.700 ;
        RECT 156.000 100.300 157.600 100.700 ;
        RECT 54.400 80.300 56.000 80.700 ;
        RECT 156.000 80.300 157.600 80.700 ;
        RECT 54.400 60.300 56.000 60.700 ;
        RECT 156.000 60.300 157.600 60.700 ;
        RECT 54.400 40.300 56.000 40.700 ;
        RECT 156.000 40.300 157.600 40.700 ;
        RECT 54.400 20.300 56.000 20.700 ;
        RECT 156.000 20.300 157.600 20.700 ;
        RECT 54.400 0.300 56.000 0.700 ;
        RECT 156.000 0.300 157.600 0.700 ;
      LAYER via3 ;
        RECT 54.600 240.300 55.000 240.700 ;
        RECT 55.400 240.300 55.800 240.700 ;
        RECT 156.200 240.300 156.600 240.700 ;
        RECT 157.000 240.300 157.400 240.700 ;
        RECT 54.600 220.300 55.000 220.700 ;
        RECT 55.400 220.300 55.800 220.700 ;
        RECT 156.200 220.300 156.600 220.700 ;
        RECT 157.000 220.300 157.400 220.700 ;
        RECT 54.600 200.300 55.000 200.700 ;
        RECT 55.400 200.300 55.800 200.700 ;
        RECT 156.200 200.300 156.600 200.700 ;
        RECT 157.000 200.300 157.400 200.700 ;
        RECT 54.600 180.300 55.000 180.700 ;
        RECT 55.400 180.300 55.800 180.700 ;
        RECT 156.200 180.300 156.600 180.700 ;
        RECT 157.000 180.300 157.400 180.700 ;
        RECT 54.600 160.300 55.000 160.700 ;
        RECT 55.400 160.300 55.800 160.700 ;
        RECT 156.200 160.300 156.600 160.700 ;
        RECT 157.000 160.300 157.400 160.700 ;
        RECT 54.600 140.300 55.000 140.700 ;
        RECT 55.400 140.300 55.800 140.700 ;
        RECT 156.200 140.300 156.600 140.700 ;
        RECT 157.000 140.300 157.400 140.700 ;
        RECT 54.600 120.300 55.000 120.700 ;
        RECT 55.400 120.300 55.800 120.700 ;
        RECT 156.200 120.300 156.600 120.700 ;
        RECT 157.000 120.300 157.400 120.700 ;
        RECT 54.600 100.300 55.000 100.700 ;
        RECT 55.400 100.300 55.800 100.700 ;
        RECT 156.200 100.300 156.600 100.700 ;
        RECT 157.000 100.300 157.400 100.700 ;
        RECT 54.600 80.300 55.000 80.700 ;
        RECT 55.400 80.300 55.800 80.700 ;
        RECT 156.200 80.300 156.600 80.700 ;
        RECT 157.000 80.300 157.400 80.700 ;
        RECT 54.600 60.300 55.000 60.700 ;
        RECT 55.400 60.300 55.800 60.700 ;
        RECT 156.200 60.300 156.600 60.700 ;
        RECT 157.000 60.300 157.400 60.700 ;
        RECT 54.600 40.300 55.000 40.700 ;
        RECT 55.400 40.300 55.800 40.700 ;
        RECT 156.200 40.300 156.600 40.700 ;
        RECT 157.000 40.300 157.400 40.700 ;
        RECT 54.600 20.300 55.000 20.700 ;
        RECT 55.400 20.300 55.800 20.700 ;
        RECT 156.200 20.300 156.600 20.700 ;
        RECT 157.000 20.300 157.400 20.700 ;
        RECT 54.600 0.300 55.000 0.700 ;
        RECT 55.400 0.300 55.800 0.700 ;
        RECT 156.200 0.300 156.600 0.700 ;
        RECT 157.000 0.300 157.400 0.700 ;
      LAYER metal4 ;
        RECT 54.400 240.300 56.000 240.700 ;
        RECT 156.000 240.300 157.600 240.700 ;
        RECT 54.400 220.300 56.000 220.700 ;
        RECT 156.000 220.300 157.600 220.700 ;
        RECT 54.400 200.300 56.000 200.700 ;
        RECT 156.000 200.300 157.600 200.700 ;
        RECT 54.400 180.300 56.000 180.700 ;
        RECT 156.000 180.300 157.600 180.700 ;
        RECT 54.400 160.300 56.000 160.700 ;
        RECT 156.000 160.300 157.600 160.700 ;
        RECT 54.400 140.300 56.000 140.700 ;
        RECT 156.000 140.300 157.600 140.700 ;
        RECT 54.400 120.300 56.000 120.700 ;
        RECT 156.000 120.300 157.600 120.700 ;
        RECT 54.400 100.300 56.000 100.700 ;
        RECT 156.000 100.300 157.600 100.700 ;
        RECT 54.400 80.300 56.000 80.700 ;
        RECT 156.000 80.300 157.600 80.700 ;
        RECT 54.400 60.300 56.000 60.700 ;
        RECT 156.000 60.300 157.600 60.700 ;
        RECT 54.400 40.300 56.000 40.700 ;
        RECT 156.000 40.300 157.600 40.700 ;
        RECT 54.400 20.300 56.000 20.700 ;
        RECT 156.000 20.300 157.600 20.700 ;
        RECT 54.400 0.300 56.000 0.700 ;
        RECT 156.000 0.300 157.600 0.700 ;
      LAYER via4 ;
        RECT 54.600 240.300 55.000 240.700 ;
        RECT 55.300 240.300 55.700 240.700 ;
        RECT 156.200 240.300 156.600 240.700 ;
        RECT 156.900 240.300 157.300 240.700 ;
        RECT 54.600 220.300 55.000 220.700 ;
        RECT 55.300 220.300 55.700 220.700 ;
        RECT 156.200 220.300 156.600 220.700 ;
        RECT 156.900 220.300 157.300 220.700 ;
        RECT 54.600 200.300 55.000 200.700 ;
        RECT 55.300 200.300 55.700 200.700 ;
        RECT 156.200 200.300 156.600 200.700 ;
        RECT 156.900 200.300 157.300 200.700 ;
        RECT 54.600 180.300 55.000 180.700 ;
        RECT 55.300 180.300 55.700 180.700 ;
        RECT 156.200 180.300 156.600 180.700 ;
        RECT 156.900 180.300 157.300 180.700 ;
        RECT 54.600 160.300 55.000 160.700 ;
        RECT 55.300 160.300 55.700 160.700 ;
        RECT 156.200 160.300 156.600 160.700 ;
        RECT 156.900 160.300 157.300 160.700 ;
        RECT 54.600 140.300 55.000 140.700 ;
        RECT 55.300 140.300 55.700 140.700 ;
        RECT 156.200 140.300 156.600 140.700 ;
        RECT 156.900 140.300 157.300 140.700 ;
        RECT 54.600 120.300 55.000 120.700 ;
        RECT 55.300 120.300 55.700 120.700 ;
        RECT 156.200 120.300 156.600 120.700 ;
        RECT 156.900 120.300 157.300 120.700 ;
        RECT 54.600 100.300 55.000 100.700 ;
        RECT 55.300 100.300 55.700 100.700 ;
        RECT 156.200 100.300 156.600 100.700 ;
        RECT 156.900 100.300 157.300 100.700 ;
        RECT 54.600 80.300 55.000 80.700 ;
        RECT 55.300 80.300 55.700 80.700 ;
        RECT 156.200 80.300 156.600 80.700 ;
        RECT 156.900 80.300 157.300 80.700 ;
        RECT 54.600 60.300 55.000 60.700 ;
        RECT 55.300 60.300 55.700 60.700 ;
        RECT 156.200 60.300 156.600 60.700 ;
        RECT 156.900 60.300 157.300 60.700 ;
        RECT 54.600 40.300 55.000 40.700 ;
        RECT 55.300 40.300 55.700 40.700 ;
        RECT 156.200 40.300 156.600 40.700 ;
        RECT 156.900 40.300 157.300 40.700 ;
        RECT 54.600 20.300 55.000 20.700 ;
        RECT 55.300 20.300 55.700 20.700 ;
        RECT 156.200 20.300 156.600 20.700 ;
        RECT 156.900 20.300 157.300 20.700 ;
        RECT 54.600 0.300 55.000 0.700 ;
        RECT 55.300 0.300 55.700 0.700 ;
        RECT 156.200 0.300 156.600 0.700 ;
        RECT 156.900 0.300 157.300 0.700 ;
      LAYER metal5 ;
        RECT 54.400 240.200 56.000 240.700 ;
        RECT 156.000 240.200 157.600 240.700 ;
        RECT 54.400 220.200 56.000 220.700 ;
        RECT 156.000 220.200 157.600 220.700 ;
        RECT 54.400 200.200 56.000 200.700 ;
        RECT 156.000 200.200 157.600 200.700 ;
        RECT 54.400 180.200 56.000 180.700 ;
        RECT 156.000 180.200 157.600 180.700 ;
        RECT 54.400 160.200 56.000 160.700 ;
        RECT 156.000 160.200 157.600 160.700 ;
        RECT 54.400 140.200 56.000 140.700 ;
        RECT 156.000 140.200 157.600 140.700 ;
        RECT 54.400 120.200 56.000 120.700 ;
        RECT 156.000 120.200 157.600 120.700 ;
        RECT 54.400 100.200 56.000 100.700 ;
        RECT 156.000 100.200 157.600 100.700 ;
        RECT 54.400 80.200 56.000 80.700 ;
        RECT 156.000 80.200 157.600 80.700 ;
        RECT 54.400 60.200 56.000 60.700 ;
        RECT 156.000 60.200 157.600 60.700 ;
        RECT 54.400 40.200 56.000 40.700 ;
        RECT 156.000 40.200 157.600 40.700 ;
        RECT 54.400 20.200 56.000 20.700 ;
        RECT 156.000 20.200 157.600 20.700 ;
        RECT 54.400 0.200 56.000 0.700 ;
        RECT 156.000 0.200 157.600 0.700 ;
      LAYER via5 ;
        RECT 55.400 240.200 55.900 240.700 ;
        RECT 157.000 240.200 157.500 240.700 ;
        RECT 55.400 220.200 55.900 220.700 ;
        RECT 157.000 220.200 157.500 220.700 ;
        RECT 55.400 200.200 55.900 200.700 ;
        RECT 157.000 200.200 157.500 200.700 ;
        RECT 55.400 180.200 55.900 180.700 ;
        RECT 157.000 180.200 157.500 180.700 ;
        RECT 55.400 160.200 55.900 160.700 ;
        RECT 157.000 160.200 157.500 160.700 ;
        RECT 55.400 140.200 55.900 140.700 ;
        RECT 157.000 140.200 157.500 140.700 ;
        RECT 55.400 120.200 55.900 120.700 ;
        RECT 157.000 120.200 157.500 120.700 ;
        RECT 55.400 100.200 55.900 100.700 ;
        RECT 157.000 100.200 157.500 100.700 ;
        RECT 55.400 80.200 55.900 80.700 ;
        RECT 157.000 80.200 157.500 80.700 ;
        RECT 55.400 60.200 55.900 60.700 ;
        RECT 157.000 60.200 157.500 60.700 ;
        RECT 55.400 40.200 55.900 40.700 ;
        RECT 157.000 40.200 157.500 40.700 ;
        RECT 55.400 20.200 55.900 20.700 ;
        RECT 157.000 20.200 157.500 20.700 ;
        RECT 55.400 0.200 55.900 0.700 ;
        RECT 157.000 0.200 157.500 0.700 ;
      LAYER metal6 ;
        RECT 54.400 -3.000 56.000 243.000 ;
        RECT 156.000 -3.000 157.600 243.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 230.800 1.000 233.100 ;
        RECT 2.200 230.800 2.600 233.100 ;
        RECT 3.800 230.800 4.200 233.100 ;
        RECT 5.400 230.800 5.800 233.100 ;
        RECT 7.000 230.800 7.400 233.100 ;
        RECT 7.800 230.800 8.200 233.100 ;
        RECT 9.400 230.800 9.800 233.100 ;
        RECT 11.000 230.800 11.400 233.100 ;
        RECT 12.600 230.800 13.000 233.100 ;
        RECT 14.200 230.800 14.600 233.100 ;
        RECT 15.000 230.800 15.400 233.100 ;
        RECT 16.600 230.800 17.000 233.100 ;
        RECT 18.200 230.800 18.600 233.100 ;
        RECT 19.800 230.800 20.200 233.100 ;
        RECT 21.400 230.800 21.800 233.100 ;
        RECT 22.200 230.800 22.600 233.100 ;
        RECT 23.800 230.800 24.200 233.100 ;
        RECT 25.400 230.800 25.800 233.100 ;
        RECT 27.000 230.800 27.400 233.100 ;
        RECT 28.600 230.800 29.000 233.100 ;
        RECT 29.400 230.800 29.800 233.100 ;
        RECT 31.000 230.800 31.400 233.100 ;
        RECT 32.600 230.800 33.000 233.100 ;
        RECT 34.200 230.800 34.600 233.100 ;
        RECT 35.800 230.800 36.200 233.100 ;
        RECT 36.600 230.800 37.000 233.100 ;
        RECT 38.200 230.800 38.600 233.100 ;
        RECT 39.800 230.800 40.200 233.100 ;
        RECT 41.400 230.800 41.800 233.100 ;
        RECT 43.000 230.800 43.400 233.100 ;
        RECT 44.600 230.800 45.000 233.100 ;
        RECT 47.300 230.800 47.800 232.100 ;
        RECT 49.000 230.800 49.400 232.100 ;
        RECT 51.800 230.800 52.200 233.000 ;
        RECT 55.000 230.800 55.400 233.100 ;
        RECT 56.600 230.800 57.000 233.100 ;
        RECT 58.200 230.800 58.600 233.100 ;
        RECT 59.800 230.800 60.200 233.100 ;
        RECT 61.400 230.800 61.800 233.100 ;
        RECT 63.000 230.800 63.400 232.700 ;
        RECT 67.000 230.800 67.400 233.100 ;
        RECT 68.600 230.800 69.000 233.100 ;
        RECT 71.300 230.800 71.800 232.100 ;
        RECT 73.000 230.800 73.400 232.100 ;
        RECT 75.800 230.800 76.200 233.000 ;
        RECT 78.200 230.800 78.600 233.100 ;
        RECT 80.900 230.800 81.400 232.100 ;
        RECT 82.600 230.800 83.000 232.100 ;
        RECT 85.400 230.800 85.800 233.000 ;
        RECT 87.000 230.800 87.400 232.100 ;
        RECT 89.200 230.800 89.600 233.500 ;
        RECT 91.800 230.800 92.200 233.300 ;
        RECT 94.200 230.800 94.600 233.100 ;
        RECT 96.900 230.800 97.400 232.100 ;
        RECT 98.600 230.800 99.000 232.100 ;
        RECT 101.400 230.800 101.800 233.000 ;
        RECT 104.600 230.800 105.000 232.700 ;
        RECT 109.400 230.800 109.800 233.100 ;
        RECT 111.000 230.800 111.400 232.700 ;
        RECT 114.200 230.800 114.600 233.100 ;
        RECT 116.900 230.800 117.400 232.100 ;
        RECT 118.600 230.800 119.000 232.100 ;
        RECT 121.400 230.800 121.800 233.000 ;
        RECT 123.800 230.800 124.200 232.700 ;
        RECT 127.800 230.800 128.200 233.100 ;
        RECT 129.400 230.800 129.800 233.100 ;
        RECT 132.100 230.800 132.600 232.100 ;
        RECT 133.800 230.800 134.200 232.100 ;
        RECT 136.600 230.800 137.000 233.000 ;
        RECT 138.200 230.800 138.600 233.100 ;
        RECT 142.200 230.800 142.600 232.700 ;
        RECT 144.100 230.800 144.500 233.100 ;
        RECT 146.200 230.800 146.600 232.100 ;
        RECT 147.000 230.800 147.400 232.100 ;
        RECT 148.600 230.800 149.000 232.100 ;
        RECT 150.200 230.800 150.600 233.000 ;
        RECT 153.000 230.800 153.400 232.100 ;
        RECT 154.600 230.800 155.100 232.100 ;
        RECT 157.400 230.800 157.800 233.100 ;
        RECT 162.200 230.800 162.600 233.100 ;
        RECT 164.600 230.800 165.000 232.700 ;
        RECT 167.000 230.800 167.400 233.100 ;
        RECT 169.700 230.800 170.200 232.100 ;
        RECT 171.400 230.800 171.800 232.100 ;
        RECT 174.200 230.800 174.600 233.000 ;
        RECT 176.600 230.800 177.000 233.300 ;
        RECT 179.200 230.800 179.600 233.500 ;
        RECT 180.600 230.800 181.000 233.100 ;
        RECT 184.600 230.800 185.000 232.700 ;
        RECT 187.000 230.800 187.400 233.100 ;
        RECT 189.700 230.800 190.200 232.100 ;
        RECT 191.400 230.800 191.800 232.100 ;
        RECT 194.200 230.800 194.600 233.000 ;
        RECT 196.600 230.800 197.000 233.000 ;
        RECT 199.400 230.800 199.800 232.100 ;
        RECT 201.000 230.800 201.500 232.100 ;
        RECT 203.800 230.800 204.200 233.100 ;
        RECT 207.000 230.800 207.400 233.100 ;
        RECT 208.600 230.800 209.000 233.100 ;
        RECT 210.200 230.800 210.600 233.100 ;
        RECT 211.800 230.800 212.200 233.100 ;
        RECT 213.400 230.800 213.800 233.100 ;
        RECT 214.200 230.800 214.600 233.100 ;
        RECT 215.800 230.800 216.200 233.100 ;
        RECT 217.400 230.800 217.800 233.100 ;
        RECT 219.000 230.800 219.400 233.100 ;
        RECT 220.600 230.800 221.000 233.100 ;
        RECT 222.200 230.800 222.600 232.700 ;
        RECT 226.200 230.800 226.600 233.100 ;
        RECT 227.000 230.800 227.400 233.100 ;
        RECT 228.600 230.800 229.000 233.100 ;
        RECT 230.200 230.800 230.600 233.100 ;
        RECT 231.800 230.800 232.200 233.100 ;
        RECT 233.400 230.800 233.800 233.100 ;
        RECT 235.000 230.800 235.400 233.100 ;
        RECT 237.700 230.800 238.200 232.100 ;
        RECT 239.400 230.800 239.800 232.100 ;
        RECT 242.200 230.800 242.600 233.000 ;
        RECT 244.600 230.800 245.000 233.000 ;
        RECT 247.400 230.800 247.800 232.100 ;
        RECT 249.000 230.800 249.500 232.100 ;
        RECT 251.800 230.800 252.200 233.100 ;
        RECT 255.000 230.800 255.400 233.100 ;
        RECT 255.800 230.800 256.200 233.100 ;
        RECT 257.400 230.800 257.800 233.100 ;
        RECT 259.000 230.800 259.400 233.100 ;
        RECT 260.600 230.800 261.000 233.100 ;
        RECT 262.200 230.800 262.600 233.100 ;
        RECT 0.200 230.200 265.400 230.800 ;
        RECT 0.600 227.900 1.000 230.200 ;
        RECT 2.200 227.900 2.600 230.200 ;
        RECT 3.800 227.900 4.200 230.200 ;
        RECT 5.400 227.900 5.800 230.200 ;
        RECT 7.000 227.900 7.400 230.200 ;
        RECT 8.600 227.900 9.000 230.200 ;
        RECT 11.300 228.900 11.800 230.200 ;
        RECT 13.000 228.900 13.400 230.200 ;
        RECT 15.800 228.000 16.200 230.200 ;
        RECT 17.700 227.900 18.100 230.200 ;
        RECT 19.800 228.900 20.200 230.200 ;
        RECT 20.600 228.900 21.000 230.200 ;
        RECT 22.200 228.900 22.600 230.200 ;
        RECT 23.800 227.900 24.200 230.200 ;
        RECT 26.500 228.900 27.000 230.200 ;
        RECT 28.200 228.900 28.600 230.200 ;
        RECT 31.000 228.000 31.400 230.200 ;
        RECT 33.400 227.700 33.800 230.200 ;
        RECT 36.000 227.500 36.400 230.200 ;
        RECT 38.200 228.900 38.600 230.200 ;
        RECT 39.800 227.700 40.200 230.200 ;
        RECT 42.400 227.500 42.800 230.200 ;
        RECT 43.800 227.900 44.200 230.200 ;
        RECT 45.400 227.900 45.800 230.200 ;
        RECT 47.800 228.900 48.200 230.200 ;
        RECT 48.600 227.900 49.000 230.200 ;
        RECT 50.200 227.900 50.600 230.200 ;
        RECT 51.800 227.900 52.200 230.200 ;
        RECT 55.000 227.900 55.400 230.200 ;
        RECT 57.700 228.900 58.200 230.200 ;
        RECT 59.400 228.900 59.800 230.200 ;
        RECT 62.200 228.000 62.600 230.200 ;
        RECT 64.600 228.300 65.000 230.200 ;
        RECT 68.600 227.900 69.000 230.200 ;
        RECT 70.000 227.500 70.400 230.200 ;
        RECT 72.600 227.700 73.000 230.200 ;
        RECT 75.000 228.000 75.400 230.200 ;
        RECT 77.800 228.900 78.200 230.200 ;
        RECT 79.400 228.900 79.900 230.200 ;
        RECT 82.200 227.900 82.600 230.200 ;
        RECT 83.800 228.900 84.200 230.200 ;
        RECT 85.400 228.900 85.800 230.200 ;
        RECT 86.200 228.900 86.600 230.200 ;
        RECT 88.300 227.900 88.700 230.200 ;
        RECT 89.400 227.900 89.800 230.200 ;
        RECT 91.000 227.900 91.400 230.200 ;
        RECT 92.600 227.900 93.000 230.200 ;
        RECT 94.200 227.900 94.600 230.200 ;
        RECT 95.800 227.900 96.200 230.200 ;
        RECT 97.400 227.900 97.800 230.200 ;
        RECT 100.100 228.900 100.600 230.200 ;
        RECT 101.800 228.900 102.200 230.200 ;
        RECT 104.600 228.000 105.000 230.200 ;
        RECT 108.600 227.700 109.000 230.200 ;
        RECT 111.200 227.500 111.600 230.200 ;
        RECT 112.600 227.900 113.000 230.200 ;
        RECT 115.800 227.900 116.200 230.200 ;
        RECT 117.400 227.900 117.800 230.200 ;
        RECT 118.200 227.900 118.600 230.200 ;
        RECT 119.800 227.900 120.200 230.200 ;
        RECT 121.400 227.900 121.800 230.200 ;
        RECT 122.800 227.500 123.200 230.200 ;
        RECT 125.400 227.700 125.800 230.200 ;
        RECT 127.800 227.700 128.200 230.200 ;
        RECT 130.400 227.500 130.800 230.200 ;
        RECT 132.600 227.700 133.000 230.200 ;
        RECT 135.200 227.500 135.600 230.200 ;
        RECT 136.600 227.900 137.000 230.200 ;
        RECT 140.600 228.300 141.000 230.200 ;
        RECT 143.000 228.000 143.400 230.200 ;
        RECT 145.800 228.900 146.200 230.200 ;
        RECT 147.400 228.900 147.900 230.200 ;
        RECT 150.200 227.900 150.600 230.200 ;
        RECT 152.600 227.700 153.000 230.200 ;
        RECT 155.200 227.500 155.600 230.200 ;
        RECT 158.800 227.500 159.200 230.200 ;
        RECT 161.400 227.700 161.800 230.200 ;
        RECT 163.800 228.000 164.200 230.200 ;
        RECT 166.600 228.900 167.000 230.200 ;
        RECT 168.200 228.900 168.700 230.200 ;
        RECT 171.000 227.900 171.400 230.200 ;
        RECT 172.600 228.900 173.000 230.200 ;
        RECT 174.200 228.900 174.600 230.200 ;
        RECT 175.000 228.900 175.400 230.200 ;
        RECT 177.100 227.900 177.500 230.200 ;
        RECT 178.800 227.500 179.200 230.200 ;
        RECT 181.400 227.700 181.800 230.200 ;
        RECT 184.600 227.900 185.000 230.200 ;
        RECT 186.200 228.000 186.600 230.200 ;
        RECT 189.000 228.900 189.400 230.200 ;
        RECT 190.600 228.900 191.100 230.200 ;
        RECT 193.400 227.900 193.800 230.200 ;
        RECT 195.000 228.900 195.400 230.200 ;
        RECT 196.600 228.900 197.000 230.200 ;
        RECT 197.400 228.900 197.800 230.200 ;
        RECT 199.500 227.900 199.900 230.200 ;
        RECT 201.400 228.000 201.800 230.200 ;
        RECT 204.200 228.900 204.600 230.200 ;
        RECT 205.800 228.900 206.300 230.200 ;
        RECT 208.600 227.900 209.000 230.200 ;
        RECT 211.800 228.900 212.200 230.200 ;
        RECT 213.400 228.900 213.800 230.200 ;
        RECT 214.200 228.900 214.600 230.200 ;
        RECT 216.300 227.900 216.700 230.200 ;
        RECT 218.200 227.900 218.600 230.200 ;
        RECT 220.900 228.900 221.400 230.200 ;
        RECT 222.600 228.900 223.000 230.200 ;
        RECT 225.400 228.000 225.800 230.200 ;
        RECT 227.000 227.900 227.400 230.200 ;
        RECT 228.600 227.900 229.000 230.200 ;
        RECT 230.200 227.900 230.600 230.200 ;
        RECT 231.600 227.500 232.000 230.200 ;
        RECT 234.200 227.700 234.600 230.200 ;
        RECT 236.600 228.300 237.000 230.200 ;
        RECT 240.600 227.900 241.000 230.200 ;
        RECT 241.400 227.900 241.800 230.200 ;
        RECT 245.400 228.300 245.800 230.200 ;
        RECT 247.000 227.900 247.400 230.200 ;
        RECT 248.600 227.900 249.000 230.200 ;
        RECT 250.200 227.900 250.600 230.200 ;
        RECT 251.800 227.900 252.200 230.200 ;
        RECT 253.400 227.900 253.800 230.200 ;
        RECT 255.800 227.900 256.200 230.200 ;
        RECT 256.600 227.900 257.000 230.200 ;
        RECT 258.200 227.900 258.600 230.200 ;
        RECT 259.800 227.900 260.200 230.200 ;
        RECT 261.400 227.900 261.800 230.200 ;
        RECT 263.000 227.900 263.400 230.200 ;
        RECT 1.400 210.800 1.800 213.000 ;
        RECT 4.200 210.800 4.600 212.100 ;
        RECT 5.800 210.800 6.300 212.100 ;
        RECT 8.600 210.800 9.000 213.100 ;
        RECT 10.200 210.800 10.600 212.100 ;
        RECT 11.800 210.800 12.200 212.100 ;
        RECT 12.600 210.800 13.000 212.100 ;
        RECT 14.700 210.800 15.100 213.100 ;
        RECT 16.600 210.800 17.000 213.000 ;
        RECT 19.400 210.800 19.800 212.100 ;
        RECT 21.000 210.800 21.500 212.100 ;
        RECT 23.800 210.800 24.200 213.100 ;
        RECT 26.200 210.800 26.600 213.000 ;
        RECT 29.000 210.800 29.400 212.100 ;
        RECT 30.600 210.800 31.100 212.100 ;
        RECT 33.400 210.800 33.800 213.100 ;
        RECT 35.000 210.800 35.400 213.100 ;
        RECT 39.000 210.800 39.400 212.700 ;
        RECT 40.600 210.800 41.000 213.100 ;
        RECT 42.200 210.800 42.600 213.100 ;
        RECT 44.600 210.800 45.000 213.300 ;
        RECT 47.200 210.800 47.600 213.500 ;
        RECT 49.400 210.800 49.800 213.100 ;
        RECT 52.100 210.800 52.600 212.100 ;
        RECT 53.800 210.800 54.200 212.100 ;
        RECT 56.600 210.800 57.000 213.000 ;
        RECT 59.800 210.800 60.200 213.100 ;
        RECT 63.800 210.800 64.200 212.700 ;
        RECT 66.200 210.800 66.600 212.700 ;
        RECT 70.200 210.800 70.600 213.100 ;
        RECT 71.800 210.800 72.200 213.000 ;
        RECT 74.600 210.800 75.000 212.100 ;
        RECT 76.200 210.800 76.700 212.100 ;
        RECT 79.000 210.800 79.400 213.100 ;
        RECT 81.400 210.800 81.800 213.000 ;
        RECT 84.200 210.800 84.600 212.100 ;
        RECT 85.800 210.800 86.300 212.100 ;
        RECT 88.600 210.800 89.000 213.100 ;
        RECT 91.000 210.800 91.400 213.100 ;
        RECT 93.700 210.800 94.200 212.100 ;
        RECT 95.400 210.800 95.800 212.100 ;
        RECT 98.200 210.800 98.600 213.000 ;
        RECT 99.800 210.800 100.200 212.100 ;
        RECT 101.900 210.800 102.300 213.100 ;
        RECT 105.400 210.800 105.800 213.000 ;
        RECT 108.200 210.800 108.600 212.100 ;
        RECT 109.800 210.800 110.300 212.100 ;
        RECT 112.600 210.800 113.000 213.100 ;
        RECT 114.200 210.800 114.600 212.100 ;
        RECT 115.800 210.800 116.200 212.100 ;
        RECT 117.400 210.800 117.800 212.100 ;
        RECT 118.200 210.800 118.600 212.100 ;
        RECT 120.300 210.800 120.700 213.100 ;
        RECT 122.200 210.800 122.600 213.000 ;
        RECT 125.000 210.800 125.400 212.100 ;
        RECT 126.600 210.800 127.100 212.100 ;
        RECT 129.400 210.800 129.800 213.100 ;
        RECT 131.600 210.800 132.000 213.500 ;
        RECT 134.200 210.800 134.600 213.300 ;
        RECT 135.800 210.800 136.200 213.100 ;
        RECT 137.400 210.800 137.800 213.100 ;
        RECT 139.800 210.800 140.200 213.100 ;
        RECT 141.400 210.800 141.800 213.100 ;
        RECT 142.200 210.800 142.600 213.100 ;
        RECT 143.800 210.800 144.200 213.100 ;
        RECT 145.400 210.800 145.800 213.100 ;
        RECT 147.000 210.800 147.400 213.100 ;
        RECT 148.600 210.800 149.000 213.100 ;
        RECT 150.200 210.800 150.600 213.000 ;
        RECT 153.000 210.800 153.400 212.100 ;
        RECT 154.600 210.800 155.100 212.100 ;
        RECT 157.400 210.800 157.800 213.100 ;
        RECT 160.600 210.800 161.000 213.100 ;
        RECT 162.200 210.800 162.600 213.100 ;
        RECT 163.800 210.800 164.200 213.100 ;
        RECT 165.400 210.800 165.800 213.100 ;
        RECT 167.000 210.800 167.400 213.100 ;
        RECT 168.600 210.800 169.000 213.000 ;
        RECT 171.400 210.800 171.800 212.100 ;
        RECT 173.000 210.800 173.500 212.100 ;
        RECT 175.800 210.800 176.200 213.100 ;
        RECT 177.400 210.800 177.800 213.100 ;
        RECT 181.400 210.800 181.800 212.700 ;
        RECT 184.600 210.800 185.000 212.700 ;
        RECT 186.200 210.800 186.600 213.100 ;
        RECT 187.800 210.800 188.200 213.100 ;
        RECT 189.400 210.800 189.800 213.100 ;
        RECT 191.000 210.800 191.400 213.100 ;
        RECT 192.600 210.800 193.000 213.100 ;
        RECT 194.200 210.800 194.600 212.700 ;
        RECT 198.200 210.800 198.600 213.100 ;
        RECT 199.800 210.800 200.200 213.000 ;
        RECT 202.600 210.800 203.000 212.100 ;
        RECT 204.200 210.800 204.700 212.100 ;
        RECT 207.000 210.800 207.400 213.100 ;
        RECT 211.000 210.800 211.400 213.100 ;
        RECT 213.700 210.800 214.200 212.100 ;
        RECT 215.400 210.800 215.800 212.100 ;
        RECT 218.200 210.800 218.600 213.000 ;
        RECT 220.600 210.800 221.000 213.100 ;
        RECT 222.200 210.800 222.600 213.100 ;
        RECT 223.000 210.800 223.400 213.100 ;
        RECT 224.600 210.800 225.000 213.100 ;
        RECT 227.000 210.800 227.400 213.000 ;
        RECT 229.800 210.800 230.200 212.100 ;
        RECT 231.400 210.800 231.900 212.100 ;
        RECT 234.200 210.800 234.600 213.100 ;
        RECT 236.600 210.800 237.000 213.000 ;
        RECT 239.400 210.800 239.800 212.100 ;
        RECT 241.000 210.800 241.500 212.100 ;
        RECT 243.800 210.800 244.200 213.100 ;
        RECT 246.200 210.800 246.600 213.100 ;
        RECT 248.900 210.800 249.400 212.100 ;
        RECT 250.600 210.800 251.000 212.100 ;
        RECT 253.400 210.800 253.800 213.000 ;
        RECT 255.800 210.800 256.200 213.100 ;
        RECT 258.500 210.800 259.000 212.100 ;
        RECT 260.200 210.800 260.600 212.100 ;
        RECT 263.000 210.800 263.400 213.000 ;
        RECT 0.200 210.200 265.400 210.800 ;
        RECT 1.400 207.900 1.800 210.200 ;
        RECT 4.100 208.900 4.600 210.200 ;
        RECT 5.800 208.900 6.200 210.200 ;
        RECT 8.600 208.000 9.000 210.200 ;
        RECT 11.800 208.300 12.200 210.200 ;
        RECT 15.000 207.900 15.400 210.200 ;
        RECT 16.600 208.900 17.000 210.200 ;
        RECT 18.000 207.500 18.400 210.200 ;
        RECT 20.600 207.700 21.000 210.200 ;
        RECT 22.800 207.500 23.200 210.200 ;
        RECT 25.400 207.700 25.800 210.200 ;
        RECT 27.600 207.500 28.000 210.200 ;
        RECT 30.200 207.700 30.600 210.200 ;
        RECT 32.600 207.900 33.000 210.200 ;
        RECT 35.300 208.900 35.800 210.200 ;
        RECT 37.000 208.900 37.400 210.200 ;
        RECT 39.800 208.000 40.200 210.200 ;
        RECT 42.200 207.700 42.600 210.200 ;
        RECT 44.800 207.500 45.200 210.200 ;
        RECT 47.000 208.900 47.400 210.200 ;
        RECT 48.600 207.700 49.000 210.200 ;
        RECT 51.200 207.500 51.600 210.200 ;
        RECT 55.000 207.900 55.400 210.200 ;
        RECT 57.700 208.900 58.200 210.200 ;
        RECT 59.400 208.900 59.800 210.200 ;
        RECT 62.200 208.000 62.600 210.200 ;
        RECT 63.800 208.900 64.200 210.200 ;
        RECT 66.000 207.500 66.400 210.200 ;
        RECT 68.600 207.700 69.000 210.200 ;
        RECT 70.800 207.500 71.200 210.200 ;
        RECT 73.400 207.700 73.800 210.200 ;
        RECT 75.000 208.900 75.400 210.200 ;
        RECT 76.600 208.900 77.000 210.200 ;
        RECT 77.400 208.900 77.800 210.200 ;
        RECT 79.500 207.900 79.900 210.200 ;
        RECT 81.400 207.900 81.800 210.200 ;
        RECT 84.100 208.900 84.600 210.200 ;
        RECT 85.800 208.900 86.200 210.200 ;
        RECT 88.600 208.000 89.000 210.200 ;
        RECT 91.800 208.300 92.200 210.200 ;
        RECT 94.200 207.700 94.600 210.200 ;
        RECT 96.800 207.500 97.200 210.200 ;
        RECT 98.200 208.900 98.600 210.200 ;
        RECT 99.800 208.900 100.200 210.200 ;
        RECT 101.200 207.500 101.600 210.200 ;
        RECT 103.800 207.700 104.200 210.200 ;
        RECT 107.800 207.700 108.200 210.200 ;
        RECT 110.400 207.500 110.800 210.200 ;
        RECT 112.600 207.700 113.000 210.200 ;
        RECT 115.200 207.500 115.600 210.200 ;
        RECT 117.400 208.300 117.800 210.200 ;
        RECT 121.400 207.900 121.800 210.200 ;
        RECT 123.000 208.000 123.400 210.200 ;
        RECT 125.800 208.900 126.200 210.200 ;
        RECT 127.400 208.900 127.900 210.200 ;
        RECT 130.200 207.900 130.600 210.200 ;
        RECT 132.600 207.900 133.000 210.200 ;
        RECT 135.300 208.900 135.800 210.200 ;
        RECT 137.000 208.900 137.400 210.200 ;
        RECT 139.800 208.000 140.200 210.200 ;
        RECT 142.200 208.300 142.600 210.200 ;
        RECT 146.200 207.900 146.600 210.200 ;
        RECT 147.800 207.700 148.200 210.200 ;
        RECT 150.400 207.500 150.800 210.200 ;
        RECT 153.400 208.300 153.800 210.200 ;
        RECT 156.600 208.300 157.000 210.200 ;
        RECT 160.600 208.300 161.000 210.200 ;
        RECT 164.600 207.900 165.000 210.200 ;
        RECT 166.200 208.000 166.600 210.200 ;
        RECT 169.000 208.900 169.400 210.200 ;
        RECT 170.600 208.900 171.100 210.200 ;
        RECT 173.400 207.900 173.800 210.200 ;
        RECT 175.800 208.000 176.200 210.200 ;
        RECT 178.600 208.900 179.000 210.200 ;
        RECT 180.200 208.900 180.700 210.200 ;
        RECT 183.000 207.900 183.400 210.200 ;
        RECT 185.400 208.000 185.800 210.200 ;
        RECT 188.200 208.900 188.600 210.200 ;
        RECT 189.800 208.900 190.300 210.200 ;
        RECT 192.600 207.900 193.000 210.200 ;
        RECT 195.000 208.300 195.400 210.200 ;
        RECT 199.000 208.300 199.400 210.200 ;
        RECT 201.400 207.700 201.800 210.200 ;
        RECT 204.000 207.500 204.400 210.200 ;
        RECT 205.400 208.900 205.800 210.200 ;
        RECT 209.200 207.500 209.600 210.200 ;
        RECT 211.800 207.700 212.200 210.200 ;
        RECT 213.400 208.900 213.800 210.200 ;
        RECT 215.000 208.900 215.400 210.200 ;
        RECT 215.800 208.900 216.200 210.200 ;
        RECT 217.900 207.900 218.300 210.200 ;
        RECT 219.800 207.700 220.200 210.200 ;
        RECT 222.400 207.500 222.800 210.200 ;
        RECT 224.600 208.300 225.000 210.200 ;
        RECT 228.600 208.300 229.000 210.200 ;
        RECT 231.000 208.000 231.400 210.200 ;
        RECT 233.800 208.900 234.200 210.200 ;
        RECT 235.400 208.900 235.900 210.200 ;
        RECT 238.200 207.900 238.600 210.200 ;
        RECT 240.600 207.700 241.000 210.200 ;
        RECT 243.200 207.500 243.600 210.200 ;
        RECT 245.400 208.900 245.800 210.200 ;
        RECT 247.000 208.000 247.400 210.200 ;
        RECT 249.800 208.900 250.200 210.200 ;
        RECT 251.400 208.900 251.900 210.200 ;
        RECT 254.200 207.900 254.600 210.200 ;
        RECT 255.800 207.900 256.200 210.200 ;
        RECT 257.400 207.900 257.800 210.200 ;
        RECT 259.000 207.900 259.400 210.200 ;
        RECT 260.600 207.900 261.000 210.200 ;
        RECT 262.200 207.900 262.600 210.200 ;
        RECT 0.600 190.800 1.000 193.100 ;
        RECT 2.200 190.800 2.600 193.100 ;
        RECT 3.800 190.800 4.200 193.100 ;
        RECT 5.400 190.800 5.800 193.100 ;
        RECT 7.000 190.800 7.400 193.100 ;
        RECT 8.600 190.800 9.000 193.100 ;
        RECT 11.300 190.800 11.800 192.100 ;
        RECT 13.000 190.800 13.400 192.100 ;
        RECT 15.800 190.800 16.200 193.000 ;
        RECT 17.400 190.800 17.800 192.100 ;
        RECT 19.000 190.800 19.400 192.100 ;
        RECT 19.800 190.800 20.200 192.100 ;
        RECT 21.900 190.800 22.300 193.100 ;
        RECT 23.000 190.800 23.400 193.100 ;
        RECT 27.000 190.800 27.400 192.700 ;
        RECT 29.400 190.800 29.800 193.000 ;
        RECT 32.200 190.800 32.600 192.100 ;
        RECT 33.800 190.800 34.300 192.100 ;
        RECT 36.600 190.800 37.000 193.100 ;
        RECT 39.000 190.800 39.400 193.100 ;
        RECT 41.700 190.800 42.200 192.100 ;
        RECT 43.400 190.800 43.800 192.100 ;
        RECT 46.200 190.800 46.600 193.000 ;
        RECT 49.400 190.800 49.800 192.700 ;
        RECT 53.400 190.800 53.800 193.000 ;
        RECT 56.200 190.800 56.600 192.100 ;
        RECT 57.800 190.800 58.300 192.100 ;
        RECT 60.600 190.800 61.000 193.100 ;
        RECT 62.500 190.800 62.900 193.100 ;
        RECT 64.600 190.800 65.000 192.100 ;
        RECT 65.400 190.800 65.800 192.100 ;
        RECT 67.000 190.800 67.400 192.100 ;
        RECT 69.400 190.800 69.800 192.700 ;
        RECT 71.800 190.800 72.200 193.000 ;
        RECT 74.600 190.800 75.000 192.100 ;
        RECT 76.200 190.800 76.700 192.100 ;
        RECT 79.000 190.800 79.400 193.100 ;
        RECT 81.400 190.800 81.800 193.300 ;
        RECT 84.000 190.800 84.400 193.500 ;
        RECT 87.000 190.800 87.400 193.100 ;
        RECT 88.600 190.800 89.000 193.300 ;
        RECT 91.200 190.800 91.600 193.500 ;
        RECT 93.400 190.800 93.800 192.100 ;
        RECT 95.000 190.800 95.400 193.000 ;
        RECT 97.800 190.800 98.200 192.100 ;
        RECT 99.400 190.800 99.900 192.100 ;
        RECT 102.200 190.800 102.600 193.100 ;
        RECT 103.800 190.800 104.200 193.100 ;
        RECT 105.400 190.800 105.800 193.100 ;
        RECT 109.400 190.800 109.800 193.000 ;
        RECT 112.200 190.800 112.600 192.100 ;
        RECT 113.800 190.800 114.300 192.100 ;
        RECT 116.600 190.800 117.000 193.100 ;
        RECT 118.200 190.800 118.600 193.100 ;
        RECT 122.200 190.800 122.600 192.700 ;
        RECT 123.800 190.800 124.200 193.100 ;
        RECT 125.400 190.800 125.800 193.100 ;
        RECT 128.600 190.800 129.000 193.100 ;
        RECT 131.000 190.800 131.400 192.700 ;
        RECT 133.400 190.800 133.800 193.100 ;
        RECT 136.100 190.800 136.600 192.100 ;
        RECT 137.800 190.800 138.200 192.100 ;
        RECT 140.600 190.800 141.000 193.000 ;
        RECT 143.000 190.800 143.400 193.300 ;
        RECT 145.600 190.800 146.000 193.500 ;
        RECT 147.600 190.800 148.000 193.500 ;
        RECT 150.200 190.800 150.600 193.300 ;
        RECT 152.600 190.800 153.000 193.100 ;
        RECT 155.000 190.800 155.400 192.700 ;
        RECT 160.600 190.800 161.000 193.100 ;
        RECT 162.200 190.800 162.600 193.000 ;
        RECT 165.000 190.800 165.400 192.100 ;
        RECT 166.600 190.800 167.100 192.100 ;
        RECT 169.400 190.800 169.800 193.100 ;
        RECT 171.000 190.800 171.400 193.100 ;
        RECT 172.600 190.800 173.000 193.100 ;
        RECT 174.200 190.800 174.600 192.100 ;
        RECT 176.400 190.800 176.800 193.500 ;
        RECT 179.000 190.800 179.400 193.300 ;
        RECT 180.600 190.800 181.000 193.100 ;
        RECT 184.600 190.800 185.000 192.700 ;
        RECT 187.000 190.800 187.400 193.300 ;
        RECT 189.600 190.800 190.000 193.500 ;
        RECT 191.800 190.800 192.200 192.100 ;
        RECT 193.400 190.800 193.800 193.000 ;
        RECT 196.200 190.800 196.600 192.100 ;
        RECT 197.800 190.800 198.300 192.100 ;
        RECT 200.600 190.800 201.000 193.100 ;
        RECT 203.000 190.800 203.400 193.000 ;
        RECT 205.800 190.800 206.200 192.100 ;
        RECT 207.400 190.800 207.900 192.100 ;
        RECT 210.200 190.800 210.600 193.100 ;
        RECT 213.400 190.800 213.800 193.100 ;
        RECT 217.400 190.800 217.800 192.700 ;
        RECT 219.800 190.800 220.200 193.300 ;
        RECT 222.400 190.800 222.800 193.500 ;
        RECT 224.600 190.800 225.000 193.100 ;
        RECT 226.200 190.800 226.600 193.100 ;
        RECT 227.800 190.800 228.200 192.700 ;
        RECT 231.800 190.800 232.200 193.100 ;
        RECT 233.400 190.800 233.800 193.000 ;
        RECT 236.200 190.800 236.600 192.100 ;
        RECT 237.800 190.800 238.300 192.100 ;
        RECT 240.600 190.800 241.000 193.100 ;
        RECT 243.000 190.800 243.400 193.300 ;
        RECT 245.600 190.800 246.000 193.500 ;
        RECT 247.800 190.800 248.200 192.700 ;
        RECT 251.000 190.800 251.400 192.100 ;
        RECT 252.600 190.800 253.000 193.000 ;
        RECT 255.400 190.800 255.800 192.100 ;
        RECT 257.000 190.800 257.500 192.100 ;
        RECT 259.800 190.800 260.200 193.100 ;
        RECT 262.200 190.800 262.600 192.700 ;
        RECT 0.200 190.200 265.400 190.800 ;
        RECT 1.400 187.900 1.800 190.200 ;
        RECT 4.100 188.900 4.600 190.200 ;
        RECT 5.800 188.900 6.200 190.200 ;
        RECT 8.600 188.000 9.000 190.200 ;
        RECT 10.200 188.900 10.600 190.200 ;
        RECT 12.400 187.500 12.800 190.200 ;
        RECT 15.000 187.700 15.400 190.200 ;
        RECT 17.400 187.900 17.800 190.200 ;
        RECT 20.100 188.900 20.600 190.200 ;
        RECT 21.800 188.900 22.200 190.200 ;
        RECT 24.600 188.000 25.000 190.200 ;
        RECT 27.000 187.700 27.400 190.200 ;
        RECT 29.600 187.500 30.000 190.200 ;
        RECT 31.800 188.900 32.200 190.200 ;
        RECT 33.200 187.500 33.600 190.200 ;
        RECT 35.800 187.700 36.200 190.200 ;
        RECT 38.000 187.500 38.400 190.200 ;
        RECT 40.600 187.700 41.000 190.200 ;
        RECT 43.000 187.700 43.400 190.200 ;
        RECT 45.600 187.500 46.000 190.200 ;
        RECT 47.000 187.900 47.400 190.200 ;
        RECT 50.200 187.700 50.600 190.200 ;
        RECT 52.800 187.500 53.200 190.200 ;
        RECT 56.600 187.700 57.000 190.200 ;
        RECT 59.200 187.500 59.600 190.200 ;
        RECT 61.400 187.700 61.800 190.200 ;
        RECT 64.000 187.500 64.400 190.200 ;
        RECT 65.400 187.900 65.800 190.200 ;
        RECT 68.600 187.700 69.000 190.200 ;
        RECT 71.200 187.500 71.600 190.200 ;
        RECT 73.400 188.900 73.800 190.200 ;
        RECT 75.000 187.900 75.400 190.200 ;
        RECT 77.700 188.900 78.200 190.200 ;
        RECT 79.400 188.900 79.800 190.200 ;
        RECT 82.200 188.000 82.600 190.200 ;
        RECT 84.600 187.700 85.000 190.200 ;
        RECT 87.200 187.500 87.600 190.200 ;
        RECT 88.600 188.900 89.000 190.200 ;
        RECT 90.800 187.500 91.200 190.200 ;
        RECT 93.400 187.700 93.800 190.200 ;
        RECT 95.600 187.500 96.000 190.200 ;
        RECT 98.200 187.700 98.600 190.200 ;
        RECT 100.400 187.500 100.800 190.200 ;
        RECT 103.000 187.700 103.400 190.200 ;
        RECT 107.000 188.000 107.400 190.200 ;
        RECT 109.800 188.900 110.200 190.200 ;
        RECT 111.400 188.900 111.900 190.200 ;
        RECT 114.200 187.900 114.600 190.200 ;
        RECT 115.800 187.900 116.200 190.200 ;
        RECT 119.800 188.300 120.200 190.200 ;
        RECT 121.400 187.900 121.800 190.200 ;
        RECT 123.000 187.900 123.400 190.200 ;
        RECT 124.600 187.900 125.000 190.200 ;
        RECT 126.200 187.900 126.600 190.200 ;
        RECT 127.800 187.900 128.200 190.200 ;
        RECT 129.400 187.900 129.800 190.200 ;
        RECT 132.100 188.900 132.600 190.200 ;
        RECT 133.800 188.900 134.200 190.200 ;
        RECT 136.600 188.000 137.000 190.200 ;
        RECT 139.000 188.300 139.400 190.200 ;
        RECT 143.000 187.900 143.400 190.200 ;
        RECT 144.600 187.900 145.000 190.200 ;
        RECT 147.300 188.900 147.800 190.200 ;
        RECT 149.000 188.900 149.400 190.200 ;
        RECT 151.800 188.000 152.200 190.200 ;
        RECT 155.800 187.900 156.200 190.200 ;
        RECT 158.500 188.900 159.000 190.200 ;
        RECT 160.200 188.900 160.600 190.200 ;
        RECT 163.000 188.000 163.400 190.200 ;
        RECT 164.600 188.900 165.000 190.200 ;
        RECT 166.800 187.500 167.200 190.200 ;
        RECT 169.400 187.700 169.800 190.200 ;
        RECT 171.600 187.500 172.000 190.200 ;
        RECT 174.200 187.700 174.600 190.200 ;
        RECT 176.600 187.700 177.000 190.200 ;
        RECT 179.200 187.500 179.600 190.200 ;
        RECT 181.400 187.700 181.800 190.200 ;
        RECT 184.000 187.500 184.400 190.200 ;
        RECT 186.200 187.900 186.600 190.200 ;
        RECT 187.800 187.900 188.200 190.200 ;
        RECT 189.400 187.700 189.800 190.200 ;
        RECT 192.000 187.500 192.400 190.200 ;
        RECT 194.000 187.500 194.400 190.200 ;
        RECT 196.600 187.700 197.000 190.200 ;
        RECT 198.800 187.500 199.200 190.200 ;
        RECT 201.400 187.700 201.800 190.200 ;
        RECT 203.800 187.700 204.200 190.200 ;
        RECT 206.400 187.500 206.800 190.200 ;
        RECT 210.200 187.700 210.600 190.200 ;
        RECT 212.800 187.500 213.200 190.200 ;
        RECT 215.000 187.700 215.400 190.200 ;
        RECT 217.600 187.500 218.000 190.200 ;
        RECT 219.800 187.900 220.200 190.200 ;
        RECT 222.500 188.900 223.000 190.200 ;
        RECT 224.200 188.900 224.600 190.200 ;
        RECT 227.000 188.000 227.400 190.200 ;
        RECT 229.200 187.500 229.600 190.200 ;
        RECT 231.800 187.700 232.200 190.200 ;
        RECT 234.000 187.500 234.400 190.200 ;
        RECT 236.600 187.700 237.000 190.200 ;
        RECT 238.200 187.900 238.600 190.200 ;
        RECT 242.200 188.300 242.600 190.200 ;
        RECT 244.600 188.000 245.000 190.200 ;
        RECT 247.400 188.900 247.800 190.200 ;
        RECT 249.000 188.900 249.500 190.200 ;
        RECT 251.800 187.900 252.200 190.200 ;
        RECT 253.400 187.900 253.800 190.200 ;
        RECT 255.000 187.900 255.400 190.200 ;
        RECT 256.600 187.900 257.000 190.200 ;
        RECT 258.200 187.900 258.600 190.200 ;
        RECT 259.800 187.900 260.200 190.200 ;
        RECT 262.200 187.900 262.600 190.200 ;
        RECT 1.400 170.800 1.800 173.000 ;
        RECT 4.200 170.800 4.600 172.100 ;
        RECT 5.800 170.800 6.300 172.100 ;
        RECT 8.600 170.800 9.000 173.100 ;
        RECT 10.800 170.800 11.200 173.500 ;
        RECT 13.400 170.800 13.800 173.300 ;
        RECT 15.800 170.800 16.200 173.300 ;
        RECT 18.400 170.800 18.800 173.500 ;
        RECT 20.400 170.800 20.800 173.500 ;
        RECT 23.000 170.800 23.400 173.300 ;
        RECT 25.200 170.800 25.600 173.500 ;
        RECT 27.800 170.800 28.200 173.300 ;
        RECT 30.000 170.800 30.400 173.500 ;
        RECT 32.600 170.800 33.000 173.300 ;
        RECT 35.800 170.800 36.200 173.100 ;
        RECT 36.800 170.800 37.200 173.100 ;
        RECT 39.800 170.800 40.200 173.100 ;
        RECT 40.800 170.800 41.200 173.100 ;
        RECT 43.800 170.800 44.200 173.100 ;
        RECT 44.600 170.800 45.000 173.100 ;
        RECT 46.200 170.800 46.600 173.100 ;
        RECT 47.800 170.800 48.200 172.100 ;
        RECT 49.400 170.800 49.800 172.100 ;
        RECT 50.800 170.800 51.200 173.500 ;
        RECT 53.400 170.800 53.800 173.300 ;
        RECT 57.400 170.800 57.800 173.300 ;
        RECT 60.000 170.800 60.400 173.500 ;
        RECT 62.000 170.800 62.400 173.500 ;
        RECT 64.600 170.800 65.000 173.300 ;
        RECT 66.200 170.800 66.600 173.100 ;
        RECT 70.200 170.800 70.600 172.700 ;
        RECT 72.600 170.800 73.000 173.000 ;
        RECT 75.400 170.800 75.800 172.100 ;
        RECT 77.000 170.800 77.500 172.100 ;
        RECT 79.800 170.800 80.200 173.100 ;
        RECT 81.400 170.800 81.800 173.100 ;
        RECT 84.400 170.800 84.800 173.100 ;
        RECT 86.200 170.800 86.600 173.000 ;
        RECT 89.000 170.800 89.400 172.100 ;
        RECT 90.600 170.800 91.100 172.100 ;
        RECT 93.400 170.800 93.800 173.100 ;
        RECT 95.000 170.800 95.400 173.100 ;
        RECT 98.000 170.800 98.400 173.100 ;
        RECT 99.600 170.800 100.000 173.500 ;
        RECT 102.200 170.800 102.600 173.300 ;
        RECT 103.800 170.800 104.200 173.100 ;
        RECT 107.800 170.800 108.200 173.100 ;
        RECT 110.800 170.800 111.200 173.100 ;
        RECT 111.800 170.800 112.200 173.100 ;
        RECT 114.200 170.800 114.600 173.100 ;
        RECT 117.200 170.800 117.600 173.100 ;
        RECT 119.000 170.800 119.400 173.000 ;
        RECT 121.800 170.800 122.200 172.100 ;
        RECT 123.400 170.800 123.900 172.100 ;
        RECT 126.200 170.800 126.600 173.100 ;
        RECT 127.800 170.800 128.200 172.100 ;
        RECT 129.400 170.800 129.800 172.100 ;
        RECT 130.200 170.800 130.600 172.100 ;
        RECT 132.300 170.800 132.700 173.100 ;
        RECT 134.200 170.800 134.600 173.100 ;
        RECT 136.900 170.800 137.400 172.100 ;
        RECT 138.600 170.800 139.000 172.100 ;
        RECT 141.400 170.800 141.800 173.000 ;
        RECT 143.000 170.800 143.400 172.100 ;
        RECT 145.200 170.800 145.600 173.500 ;
        RECT 147.800 170.800 148.200 173.300 ;
        RECT 149.700 170.800 150.100 173.100 ;
        RECT 151.800 170.800 152.200 172.100 ;
        RECT 154.200 170.800 154.600 173.100 ;
        RECT 157.400 170.800 157.800 173.100 ;
        RECT 160.100 170.800 160.600 172.100 ;
        RECT 161.800 170.800 162.200 172.100 ;
        RECT 164.600 170.800 165.000 173.000 ;
        RECT 166.200 170.800 166.600 172.100 ;
        RECT 168.400 170.800 168.800 173.500 ;
        RECT 171.000 170.800 171.400 173.300 ;
        RECT 173.400 170.800 173.800 173.100 ;
        RECT 176.100 170.800 176.600 172.100 ;
        RECT 177.800 170.800 178.200 172.100 ;
        RECT 180.600 170.800 181.000 173.000 ;
        RECT 183.000 170.800 183.400 173.000 ;
        RECT 185.800 170.800 186.200 172.100 ;
        RECT 187.400 170.800 187.900 172.100 ;
        RECT 190.200 170.800 190.600 173.100 ;
        RECT 192.600 170.800 193.000 173.300 ;
        RECT 195.200 170.800 195.600 173.500 ;
        RECT 197.400 170.800 197.800 173.100 ;
        RECT 200.100 170.800 200.600 172.100 ;
        RECT 201.800 170.800 202.200 172.100 ;
        RECT 204.600 170.800 205.000 173.000 ;
        RECT 207.000 170.800 207.400 172.100 ;
        RECT 211.000 170.800 211.400 173.100 ;
        RECT 212.000 170.800 212.400 173.100 ;
        RECT 215.000 170.800 215.400 173.100 ;
        RECT 215.800 170.800 216.200 173.100 ;
        RECT 218.800 170.800 219.200 173.100 ;
        RECT 220.400 170.800 220.800 173.500 ;
        RECT 223.000 170.800 223.400 173.300 ;
        RECT 225.400 170.800 225.800 173.300 ;
        RECT 228.000 170.800 228.400 173.500 ;
        RECT 231.000 170.800 231.400 172.700 ;
        RECT 234.200 170.800 234.600 172.700 ;
        RECT 237.400 170.800 237.800 173.100 ;
        RECT 239.000 170.800 239.400 173.000 ;
        RECT 241.800 170.800 242.200 172.100 ;
        RECT 243.400 170.800 243.900 172.100 ;
        RECT 246.200 170.800 246.600 173.100 ;
        RECT 249.400 170.800 249.800 172.700 ;
        RECT 251.800 170.800 252.200 173.000 ;
        RECT 254.600 170.800 255.000 172.100 ;
        RECT 256.200 170.800 256.700 172.100 ;
        RECT 259.000 170.800 259.400 173.100 ;
        RECT 262.200 170.800 262.600 173.100 ;
        RECT 0.200 170.200 265.400 170.800 ;
        RECT 1.400 167.900 1.800 170.200 ;
        RECT 4.100 168.900 4.600 170.200 ;
        RECT 5.800 168.900 6.200 170.200 ;
        RECT 8.600 168.000 9.000 170.200 ;
        RECT 10.200 167.900 10.600 170.200 ;
        RECT 14.200 168.300 14.600 170.200 ;
        RECT 16.600 167.900 17.000 170.200 ;
        RECT 19.300 168.900 19.800 170.200 ;
        RECT 21.000 168.900 21.400 170.200 ;
        RECT 23.800 168.000 24.200 170.200 ;
        RECT 25.400 168.900 25.800 170.200 ;
        RECT 27.600 167.500 28.000 170.200 ;
        RECT 30.200 167.700 30.600 170.200 ;
        RECT 31.800 167.900 32.200 170.200 ;
        RECT 35.800 168.300 36.200 170.200 ;
        RECT 39.000 168.300 39.400 170.200 ;
        RECT 41.400 168.000 41.800 170.200 ;
        RECT 44.200 168.900 44.600 170.200 ;
        RECT 45.800 168.900 46.300 170.200 ;
        RECT 48.600 167.900 49.000 170.200 ;
        RECT 50.200 168.900 50.600 170.200 ;
        RECT 52.300 167.900 52.700 170.200 ;
        RECT 55.800 168.000 56.200 170.200 ;
        RECT 58.600 168.900 59.000 170.200 ;
        RECT 60.200 168.900 60.700 170.200 ;
        RECT 63.000 167.900 63.400 170.200 ;
        RECT 64.600 167.900 65.000 170.200 ;
        RECT 68.600 168.300 69.000 170.200 ;
        RECT 71.000 168.000 71.400 170.200 ;
        RECT 73.800 168.900 74.200 170.200 ;
        RECT 75.400 168.900 75.900 170.200 ;
        RECT 78.200 167.900 78.600 170.200 ;
        RECT 79.800 167.900 80.200 170.200 ;
        RECT 81.400 167.900 81.800 170.200 ;
        RECT 83.000 167.900 83.400 170.200 ;
        RECT 84.600 167.900 85.000 170.200 ;
        RECT 86.200 167.900 86.600 170.200 ;
        RECT 87.600 167.500 88.000 170.200 ;
        RECT 90.200 167.700 90.600 170.200 ;
        RECT 92.400 167.500 92.800 170.200 ;
        RECT 95.000 167.700 95.400 170.200 ;
        RECT 96.600 167.900 97.000 170.200 ;
        RECT 99.800 167.700 100.200 170.200 ;
        RECT 102.400 167.500 102.800 170.200 ;
        RECT 106.200 167.900 106.600 170.200 ;
        RECT 108.900 168.900 109.400 170.200 ;
        RECT 110.600 168.900 111.000 170.200 ;
        RECT 113.400 168.000 113.800 170.200 ;
        RECT 115.000 168.900 115.400 170.200 ;
        RECT 117.200 167.500 117.600 170.200 ;
        RECT 119.800 167.700 120.200 170.200 ;
        RECT 122.200 167.900 122.600 170.200 ;
        RECT 123.800 167.900 124.200 170.200 ;
        RECT 125.400 167.700 125.800 170.200 ;
        RECT 128.000 167.500 128.400 170.200 ;
        RECT 130.200 167.700 130.600 170.200 ;
        RECT 132.800 167.500 133.200 170.200 ;
        RECT 134.800 167.500 135.200 170.200 ;
        RECT 137.400 167.700 137.800 170.200 ;
        RECT 139.000 167.900 139.400 170.200 ;
        RECT 142.000 167.900 142.400 170.200 ;
        RECT 143.000 167.900 143.400 170.200 ;
        RECT 146.200 168.300 146.600 170.200 ;
        RECT 148.800 167.900 149.200 170.200 ;
        RECT 151.800 167.900 152.200 170.200 ;
        RECT 153.200 167.500 153.600 170.200 ;
        RECT 155.800 167.700 156.200 170.200 ;
        RECT 159.600 167.500 160.000 170.200 ;
        RECT 162.200 167.700 162.600 170.200 ;
        RECT 164.600 167.700 165.000 170.200 ;
        RECT 167.200 167.500 167.600 170.200 ;
        RECT 169.400 168.300 169.800 170.200 ;
        RECT 172.600 167.700 173.000 170.200 ;
        RECT 175.200 167.500 175.600 170.200 ;
        RECT 177.400 167.700 177.800 170.200 ;
        RECT 180.000 167.500 180.400 170.200 ;
        RECT 181.700 167.900 182.100 170.200 ;
        RECT 183.800 168.900 184.200 170.200 ;
        RECT 184.600 168.900 185.000 170.200 ;
        RECT 186.200 168.900 186.600 170.200 ;
        RECT 187.200 167.900 187.600 170.200 ;
        RECT 190.200 167.900 190.600 170.200 ;
        RECT 192.600 167.900 193.000 170.200 ;
        RECT 194.200 168.300 194.600 170.200 ;
        RECT 196.800 167.900 197.200 170.200 ;
        RECT 199.800 167.900 200.200 170.200 ;
        RECT 202.200 168.300 202.600 170.200 ;
        RECT 206.200 168.000 206.600 170.200 ;
        RECT 209.000 168.900 209.400 170.200 ;
        RECT 210.600 168.900 211.100 170.200 ;
        RECT 213.400 167.900 213.800 170.200 ;
        RECT 215.000 168.900 215.400 170.200 ;
        RECT 217.200 167.500 217.600 170.200 ;
        RECT 219.800 167.700 220.200 170.200 ;
        RECT 222.000 167.500 222.400 170.200 ;
        RECT 224.600 167.700 225.000 170.200 ;
        RECT 226.800 167.500 227.200 170.200 ;
        RECT 229.400 167.700 229.800 170.200 ;
        RECT 231.600 167.500 232.000 170.200 ;
        RECT 234.200 167.700 234.600 170.200 ;
        RECT 237.400 168.300 237.800 170.200 ;
        RECT 239.000 168.900 239.400 170.200 ;
        RECT 240.600 168.900 241.000 170.200 ;
        RECT 241.400 168.900 241.800 170.200 ;
        RECT 243.500 167.900 243.900 170.200 ;
        RECT 244.600 167.900 245.000 170.200 ;
        RECT 247.800 168.000 248.200 170.200 ;
        RECT 250.600 168.900 251.000 170.200 ;
        RECT 252.200 168.900 252.700 170.200 ;
        RECT 255.000 167.900 255.400 170.200 ;
        RECT 256.600 168.900 257.000 170.200 ;
        RECT 258.700 167.900 259.100 170.200 ;
        RECT 260.600 167.900 261.000 170.200 ;
        RECT 263.000 167.900 263.400 170.200 ;
        RECT 1.400 150.800 1.800 153.100 ;
        RECT 4.100 150.800 4.600 152.100 ;
        RECT 5.800 150.800 6.200 152.100 ;
        RECT 8.600 150.800 9.000 153.000 ;
        RECT 10.200 150.800 10.600 153.100 ;
        RECT 12.600 150.800 13.000 153.100 ;
        RECT 14.200 150.800 14.600 153.100 ;
        RECT 15.800 150.800 16.200 153.100 ;
        RECT 17.400 150.800 17.800 153.100 ;
        RECT 19.000 150.800 19.400 153.100 ;
        RECT 20.600 150.800 21.000 153.100 ;
        RECT 23.300 150.800 23.800 152.100 ;
        RECT 25.000 150.800 25.400 152.100 ;
        RECT 27.800 150.800 28.200 153.000 ;
        RECT 30.200 150.800 30.600 153.100 ;
        RECT 32.900 150.800 33.400 152.100 ;
        RECT 34.600 150.800 35.000 152.100 ;
        RECT 37.400 150.800 37.800 153.000 ;
        RECT 39.000 150.800 39.400 152.100 ;
        RECT 40.600 150.800 41.000 152.100 ;
        RECT 41.400 150.800 41.800 152.100 ;
        RECT 43.500 150.800 43.900 153.100 ;
        RECT 44.600 150.800 45.000 153.100 ;
        RECT 46.200 150.800 46.600 153.100 ;
        RECT 48.600 150.800 49.000 153.300 ;
        RECT 51.200 150.800 51.600 153.500 ;
        RECT 53.400 150.800 53.800 152.100 ;
        RECT 56.600 150.800 57.000 153.100 ;
        RECT 59.300 150.800 59.800 152.100 ;
        RECT 61.000 150.800 61.400 152.100 ;
        RECT 63.800 150.800 64.200 153.000 ;
        RECT 66.200 150.800 66.600 153.100 ;
        RECT 68.900 150.800 69.400 152.100 ;
        RECT 70.600 150.800 71.000 152.100 ;
        RECT 73.400 150.800 73.800 153.000 ;
        RECT 75.600 150.800 76.000 153.500 ;
        RECT 78.200 150.800 78.600 153.300 ;
        RECT 79.800 150.800 80.200 153.100 ;
        RECT 83.800 150.800 84.200 152.700 ;
        RECT 86.000 150.800 86.400 153.500 ;
        RECT 88.600 150.800 89.000 153.300 ;
        RECT 91.000 150.800 91.400 153.100 ;
        RECT 93.700 150.800 94.200 152.100 ;
        RECT 95.400 150.800 95.800 152.100 ;
        RECT 98.200 150.800 98.600 153.000 ;
        RECT 100.600 150.800 101.000 153.300 ;
        RECT 103.200 150.800 103.600 153.500 ;
        RECT 104.600 150.800 105.000 153.100 ;
        RECT 110.200 150.800 110.600 152.700 ;
        RECT 111.800 150.800 112.200 153.100 ;
        RECT 114.200 150.800 114.600 152.100 ;
        RECT 115.800 150.800 116.200 152.100 ;
        RECT 117.400 150.800 117.800 153.100 ;
        RECT 120.100 150.800 120.600 152.100 ;
        RECT 121.800 150.800 122.200 152.100 ;
        RECT 124.600 150.800 125.000 153.000 ;
        RECT 127.000 150.800 127.400 152.700 ;
        RECT 131.000 150.800 131.400 152.700 ;
        RECT 133.400 150.800 133.800 153.100 ;
        RECT 136.100 150.800 136.600 152.100 ;
        RECT 137.800 150.800 138.200 152.100 ;
        RECT 140.600 150.800 141.000 153.000 ;
        RECT 143.800 150.800 144.200 153.100 ;
        RECT 144.600 150.800 145.000 153.100 ;
        RECT 148.600 150.800 149.000 152.700 ;
        RECT 151.800 150.800 152.200 153.100 ;
        RECT 155.000 150.800 155.400 153.000 ;
        RECT 157.800 150.800 158.200 152.100 ;
        RECT 159.400 150.800 159.900 152.100 ;
        RECT 162.200 150.800 162.600 153.100 ;
        RECT 165.400 150.800 165.800 153.100 ;
        RECT 167.800 150.800 168.200 152.700 ;
        RECT 169.400 150.800 169.800 152.100 ;
        RECT 171.000 150.800 171.400 152.100 ;
        RECT 172.100 150.800 172.500 153.100 ;
        RECT 174.200 150.800 174.600 152.100 ;
        RECT 175.800 150.800 176.200 152.700 ;
        RECT 178.800 150.800 179.200 153.500 ;
        RECT 181.400 150.800 181.800 153.300 ;
        RECT 183.800 150.800 184.200 153.100 ;
        RECT 186.500 150.800 187.000 152.100 ;
        RECT 188.200 150.800 188.600 152.100 ;
        RECT 191.000 150.800 191.400 153.000 ;
        RECT 193.400 150.800 193.800 152.700 ;
        RECT 196.600 150.800 197.000 152.700 ;
        RECT 199.000 150.800 199.400 153.100 ;
        RECT 203.000 150.800 203.400 152.700 ;
        RECT 205.200 150.800 205.600 153.500 ;
        RECT 207.800 150.800 208.200 153.300 ;
        RECT 211.000 150.800 211.400 153.100 ;
        RECT 214.000 150.800 214.400 153.100 ;
        RECT 215.800 150.800 216.200 153.300 ;
        RECT 218.400 150.800 218.800 153.500 ;
        RECT 220.400 150.800 220.800 153.500 ;
        RECT 223.000 150.800 223.400 153.300 ;
        RECT 225.400 150.800 225.800 153.300 ;
        RECT 228.000 150.800 228.400 153.500 ;
        RECT 229.400 150.800 229.800 152.100 ;
        RECT 231.500 150.800 231.900 153.100 ;
        RECT 233.400 150.800 233.800 153.100 ;
        RECT 236.100 150.800 236.600 152.100 ;
        RECT 237.800 150.800 238.200 152.100 ;
        RECT 240.600 150.800 241.000 153.000 ;
        RECT 243.800 150.800 244.200 153.100 ;
        RECT 244.600 150.800 245.000 153.100 ;
        RECT 248.600 150.800 249.000 152.700 ;
        RECT 250.200 150.800 250.600 153.100 ;
        RECT 254.200 150.800 254.600 152.700 ;
        RECT 256.600 150.800 257.000 153.000 ;
        RECT 259.400 150.800 259.800 152.100 ;
        RECT 261.000 150.800 261.500 152.100 ;
        RECT 263.800 150.800 264.200 153.100 ;
        RECT 0.200 150.200 265.400 150.800 ;
        RECT 1.400 147.900 1.800 150.200 ;
        RECT 4.100 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.200 150.200 ;
        RECT 8.600 148.000 9.000 150.200 ;
        RECT 11.800 148.300 12.200 150.200 ;
        RECT 14.200 148.300 14.600 150.200 ;
        RECT 18.200 147.900 18.600 150.200 ;
        RECT 19.800 147.700 20.200 150.200 ;
        RECT 22.400 147.500 22.800 150.200 ;
        RECT 23.800 147.900 24.200 150.200 ;
        RECT 25.400 147.900 25.800 150.200 ;
        RECT 27.000 147.900 27.400 150.200 ;
        RECT 28.600 147.900 29.000 150.200 ;
        RECT 30.200 147.900 30.600 150.200 ;
        RECT 31.800 147.700 32.200 150.200 ;
        RECT 34.400 147.500 34.800 150.200 ;
        RECT 36.600 148.900 37.000 150.200 ;
        RECT 38.200 147.700 38.600 150.200 ;
        RECT 40.800 147.500 41.200 150.200 ;
        RECT 42.200 147.900 42.600 150.200 ;
        RECT 43.800 147.900 44.200 150.200 ;
        RECT 45.400 147.900 45.800 150.200 ;
        RECT 47.000 147.900 47.400 150.200 ;
        RECT 48.600 147.900 49.000 150.200 ;
        RECT 50.200 147.900 50.600 150.200 ;
        RECT 52.900 148.900 53.400 150.200 ;
        RECT 54.600 148.900 55.000 150.200 ;
        RECT 57.400 148.000 57.800 150.200 ;
        RECT 61.400 148.300 61.800 150.200 ;
        RECT 65.400 147.900 65.800 150.200 ;
        RECT 67.000 147.700 67.400 150.200 ;
        RECT 69.600 147.500 70.000 150.200 ;
        RECT 71.800 147.700 72.200 150.200 ;
        RECT 74.400 147.500 74.800 150.200 ;
        RECT 76.600 148.000 77.000 150.200 ;
        RECT 79.400 148.900 79.800 150.200 ;
        RECT 81.000 148.900 81.500 150.200 ;
        RECT 83.800 147.900 84.200 150.200 ;
        RECT 85.400 148.900 85.800 150.200 ;
        RECT 87.600 147.500 88.000 150.200 ;
        RECT 90.200 147.700 90.600 150.200 ;
        RECT 91.800 148.900 92.200 150.200 ;
        RECT 94.000 147.500 94.400 150.200 ;
        RECT 96.600 147.700 97.000 150.200 ;
        RECT 100.600 146.900 101.000 150.200 ;
        RECT 101.400 146.900 101.800 150.200 ;
        RECT 106.200 146.900 106.600 150.200 ;
        RECT 110.200 147.900 110.600 150.200 ;
        RECT 112.900 148.900 113.400 150.200 ;
        RECT 114.600 148.900 115.000 150.200 ;
        RECT 117.400 148.000 117.800 150.200 ;
        RECT 119.000 148.900 119.400 150.200 ;
        RECT 121.100 147.900 121.500 150.200 ;
        RECT 123.000 148.000 123.400 150.200 ;
        RECT 125.800 148.900 126.200 150.200 ;
        RECT 127.400 148.900 127.900 150.200 ;
        RECT 130.200 147.900 130.600 150.200 ;
        RECT 133.400 147.900 133.800 150.200 ;
        RECT 135.000 147.900 135.400 150.200 ;
        RECT 135.800 148.900 136.200 150.200 ;
        RECT 137.400 148.900 137.800 150.200 ;
        RECT 139.000 147.900 139.400 150.200 ;
        RECT 140.600 147.900 141.000 150.200 ;
        RECT 143.800 146.900 144.200 150.200 ;
        RECT 144.600 146.900 145.000 150.200 ;
        RECT 147.800 146.900 148.200 150.200 ;
        RECT 151.800 147.900 152.200 150.200 ;
        RECT 153.400 147.900 153.800 150.200 ;
        RECT 154.200 147.900 154.600 150.200 ;
        RECT 158.200 147.900 158.600 150.200 ;
        RECT 163.000 146.900 163.400 150.200 ;
        RECT 163.800 147.900 164.200 150.200 ;
        RECT 165.400 147.900 165.800 150.200 ;
        RECT 167.000 147.900 167.400 150.200 ;
        RECT 168.600 148.000 169.000 150.200 ;
        RECT 171.400 148.900 171.800 150.200 ;
        RECT 173.000 148.900 173.500 150.200 ;
        RECT 175.800 147.900 176.200 150.200 ;
        RECT 178.200 147.700 178.600 150.200 ;
        RECT 180.800 147.500 181.200 150.200 ;
        RECT 183.000 148.900 183.400 150.200 ;
        RECT 184.600 147.900 185.000 150.200 ;
        RECT 186.200 147.900 186.600 150.200 ;
        RECT 187.800 148.000 188.200 150.200 ;
        RECT 190.600 148.900 191.000 150.200 ;
        RECT 192.200 148.900 192.700 150.200 ;
        RECT 195.000 147.900 195.400 150.200 ;
        RECT 197.200 147.500 197.600 150.200 ;
        RECT 199.800 147.700 200.200 150.200 ;
        RECT 202.200 148.300 202.600 150.200 ;
        RECT 206.200 148.300 206.600 150.200 ;
        RECT 210.200 148.000 210.600 150.200 ;
        RECT 213.000 148.900 213.400 150.200 ;
        RECT 214.600 148.900 215.100 150.200 ;
        RECT 217.400 147.900 217.800 150.200 ;
        RECT 219.800 147.900 220.200 150.200 ;
        RECT 221.400 147.900 221.800 150.200 ;
        RECT 222.800 147.500 223.200 150.200 ;
        RECT 225.400 147.700 225.800 150.200 ;
        RECT 227.000 147.900 227.400 150.200 ;
        RECT 231.000 148.300 231.400 150.200 ;
        RECT 233.400 147.900 233.800 150.200 ;
        RECT 236.100 148.900 236.600 150.200 ;
        RECT 237.800 148.900 238.200 150.200 ;
        RECT 240.600 148.000 241.000 150.200 ;
        RECT 243.000 148.300 243.400 150.200 ;
        RECT 247.000 147.900 247.400 150.200 ;
        RECT 247.800 147.900 248.200 150.200 ;
        RECT 251.000 148.000 251.400 150.200 ;
        RECT 253.800 148.900 254.200 150.200 ;
        RECT 255.400 148.900 255.900 150.200 ;
        RECT 258.200 147.900 258.600 150.200 ;
        RECT 259.800 147.900 260.200 150.200 ;
        RECT 261.400 147.900 261.800 150.200 ;
        RECT 263.000 147.900 263.400 150.200 ;
        RECT 1.400 130.800 1.800 133.100 ;
        RECT 4.100 130.800 4.600 132.100 ;
        RECT 5.800 130.800 6.200 132.100 ;
        RECT 8.600 130.800 9.000 133.000 ;
        RECT 10.200 130.800 10.600 132.100 ;
        RECT 11.800 130.800 12.200 132.100 ;
        RECT 12.600 130.800 13.000 132.100 ;
        RECT 14.700 130.800 15.100 133.100 ;
        RECT 16.400 130.800 16.800 133.500 ;
        RECT 19.000 130.800 19.400 133.300 ;
        RECT 21.200 130.800 21.600 133.500 ;
        RECT 23.800 130.800 24.200 133.300 ;
        RECT 25.400 130.800 25.800 133.100 ;
        RECT 27.000 130.800 27.400 133.100 ;
        RECT 29.200 130.800 29.600 133.500 ;
        RECT 31.800 130.800 32.200 133.300 ;
        RECT 34.200 130.800 34.600 132.100 ;
        RECT 35.800 130.800 36.200 133.000 ;
        RECT 38.600 130.800 39.000 132.100 ;
        RECT 40.200 130.800 40.700 132.100 ;
        RECT 43.000 130.800 43.400 133.100 ;
        RECT 45.400 130.800 45.800 133.100 ;
        RECT 48.100 130.800 48.600 132.100 ;
        RECT 49.800 130.800 50.200 132.100 ;
        RECT 52.600 130.800 53.000 133.000 ;
        RECT 56.600 130.800 57.000 132.700 ;
        RECT 59.000 130.800 59.400 133.100 ;
        RECT 60.600 130.800 61.000 133.100 ;
        RECT 62.200 130.800 62.600 133.100 ;
        RECT 63.800 130.800 64.200 133.100 ;
        RECT 65.400 130.800 65.800 133.100 ;
        RECT 66.200 130.800 66.600 133.100 ;
        RECT 67.800 130.800 68.200 133.100 ;
        RECT 69.400 130.800 69.800 133.100 ;
        RECT 71.000 130.800 71.400 133.100 ;
        RECT 73.400 130.800 73.800 133.300 ;
        RECT 76.000 130.800 76.400 133.500 ;
        RECT 78.200 130.800 78.600 133.100 ;
        RECT 80.900 130.800 81.400 132.100 ;
        RECT 82.600 130.800 83.000 132.100 ;
        RECT 85.400 130.800 85.800 133.000 ;
        RECT 88.600 130.800 89.000 132.700 ;
        RECT 91.000 130.800 91.400 133.000 ;
        RECT 93.800 130.800 94.200 132.100 ;
        RECT 95.400 130.800 95.900 132.100 ;
        RECT 98.200 130.800 98.600 133.100 ;
        RECT 102.200 130.800 102.600 134.100 ;
        RECT 103.000 130.800 103.400 133.100 ;
        RECT 107.000 130.800 107.400 133.100 ;
        RECT 110.000 130.800 110.400 133.100 ;
        RECT 111.800 130.800 112.200 133.100 ;
        RECT 114.500 130.800 115.000 132.100 ;
        RECT 116.200 130.800 116.600 132.100 ;
        RECT 119.000 130.800 119.400 133.000 ;
        RECT 121.400 130.800 121.800 132.700 ;
        RECT 125.400 130.800 125.800 133.100 ;
        RECT 126.200 130.800 126.600 133.100 ;
        RECT 127.800 130.800 128.200 133.100 ;
        RECT 129.400 130.800 129.800 133.100 ;
        RECT 131.000 130.800 131.400 133.100 ;
        RECT 132.600 130.800 133.000 133.100 ;
        RECT 133.400 130.800 133.800 133.100 ;
        RECT 135.000 130.800 135.400 133.100 ;
        RECT 136.600 130.800 137.000 133.100 ;
        RECT 139.800 130.800 140.200 133.100 ;
        RECT 140.600 130.800 141.000 133.100 ;
        RECT 144.600 130.800 145.000 133.100 ;
        RECT 145.400 130.800 145.800 133.100 ;
        RECT 147.800 130.800 148.200 132.100 ;
        RECT 149.400 130.800 149.800 132.100 ;
        RECT 150.200 130.800 150.600 132.100 ;
        RECT 151.800 130.800 152.200 132.100 ;
        RECT 154.200 130.800 154.600 133.100 ;
        RECT 156.600 130.800 157.000 133.100 ;
        RECT 160.600 130.800 161.000 133.100 ;
        RECT 161.400 130.800 161.800 132.100 ;
        RECT 163.000 130.800 163.400 132.100 ;
        RECT 165.400 130.800 165.800 133.100 ;
        RECT 166.200 130.800 166.600 132.100 ;
        RECT 167.800 130.800 168.200 132.100 ;
        RECT 169.400 130.800 169.800 133.000 ;
        RECT 172.200 130.800 172.600 132.100 ;
        RECT 173.800 130.800 174.300 132.100 ;
        RECT 176.600 130.800 177.000 133.100 ;
        RECT 179.000 130.800 179.400 133.300 ;
        RECT 181.600 130.800 182.000 133.500 ;
        RECT 183.800 130.800 184.200 132.100 ;
        RECT 185.400 130.800 185.800 133.100 ;
        RECT 188.100 130.800 188.600 132.100 ;
        RECT 189.800 130.800 190.200 132.100 ;
        RECT 192.600 130.800 193.000 133.000 ;
        RECT 194.200 130.800 194.600 133.100 ;
        RECT 196.400 130.800 196.800 133.500 ;
        RECT 199.000 130.800 199.400 133.300 ;
        RECT 200.600 130.800 201.000 133.100 ;
        RECT 203.600 130.800 204.000 133.100 ;
        RECT 204.600 130.800 205.000 133.100 ;
        RECT 207.800 130.800 208.200 133.100 ;
        RECT 211.000 130.800 211.400 133.100 ;
        RECT 212.600 130.800 213.000 133.100 ;
        RECT 214.000 130.800 214.400 133.500 ;
        RECT 216.600 130.800 217.000 133.300 ;
        RECT 218.200 130.800 218.600 132.100 ;
        RECT 220.300 130.800 220.700 133.100 ;
        RECT 221.400 130.800 221.800 132.100 ;
        RECT 223.000 130.800 223.400 132.100 ;
        RECT 224.600 130.800 225.000 133.000 ;
        RECT 227.400 130.800 227.800 132.100 ;
        RECT 229.000 130.800 229.500 132.100 ;
        RECT 231.800 130.800 232.200 133.100 ;
        RECT 233.400 130.800 233.800 133.100 ;
        RECT 235.000 130.800 235.400 133.100 ;
        RECT 236.600 130.800 237.000 133.100 ;
        RECT 238.200 130.800 238.600 133.100 ;
        RECT 239.800 130.800 240.200 133.100 ;
        RECT 240.900 130.800 241.300 133.100 ;
        RECT 243.000 130.800 243.400 132.100 ;
        RECT 244.600 130.800 245.000 133.000 ;
        RECT 247.400 130.800 247.800 132.100 ;
        RECT 249.000 130.800 249.500 132.100 ;
        RECT 251.800 130.800 252.200 133.100 ;
        RECT 253.700 130.800 254.100 133.100 ;
        RECT 255.800 130.800 256.200 132.100 ;
        RECT 256.600 130.800 257.000 132.100 ;
        RECT 258.200 130.800 258.600 132.100 ;
        RECT 259.000 130.800 259.400 132.100 ;
        RECT 260.600 130.800 261.000 132.100 ;
        RECT 262.200 130.800 262.600 133.100 ;
        RECT 0.200 130.200 265.400 130.800 ;
        RECT 0.600 127.900 1.000 130.200 ;
        RECT 2.200 127.900 2.600 130.200 ;
        RECT 3.800 127.900 4.200 130.200 ;
        RECT 5.400 127.900 5.800 130.200 ;
        RECT 7.000 127.900 7.400 130.200 ;
        RECT 8.600 127.900 9.000 130.200 ;
        RECT 11.300 128.900 11.800 130.200 ;
        RECT 13.000 128.900 13.400 130.200 ;
        RECT 15.800 128.000 16.200 130.200 ;
        RECT 17.400 127.900 17.800 130.200 ;
        RECT 21.400 128.300 21.800 130.200 ;
        RECT 23.600 127.500 24.000 130.200 ;
        RECT 26.200 127.700 26.600 130.200 ;
        RECT 28.600 127.900 29.000 130.200 ;
        RECT 31.300 128.900 31.800 130.200 ;
        RECT 33.000 128.900 33.400 130.200 ;
        RECT 35.800 128.000 36.200 130.200 ;
        RECT 38.200 128.300 38.600 130.200 ;
        RECT 42.200 127.900 42.600 130.200 ;
        RECT 43.200 127.900 43.600 130.200 ;
        RECT 46.200 127.900 46.600 130.200 ;
        RECT 47.600 127.500 48.000 130.200 ;
        RECT 50.200 127.700 50.600 130.200 ;
        RECT 52.400 127.500 52.800 130.200 ;
        RECT 55.000 127.700 55.400 130.200 ;
        RECT 59.800 127.900 60.200 130.200 ;
        RECT 61.400 127.700 61.800 130.200 ;
        RECT 64.000 127.500 64.400 130.200 ;
        RECT 65.400 127.900 65.800 130.200 ;
        RECT 68.400 127.900 68.800 130.200 ;
        RECT 70.200 127.900 70.600 130.200 ;
        RECT 72.900 128.900 73.400 130.200 ;
        RECT 74.600 128.900 75.000 130.200 ;
        RECT 77.400 128.000 77.800 130.200 ;
        RECT 79.800 128.300 80.200 130.200 ;
        RECT 82.200 127.900 82.600 130.200 ;
        RECT 84.600 127.900 85.000 130.200 ;
        RECT 87.800 127.700 88.200 130.200 ;
        RECT 90.400 127.500 90.800 130.200 ;
        RECT 92.600 128.000 93.000 130.200 ;
        RECT 95.400 128.900 95.800 130.200 ;
        RECT 97.000 128.900 97.500 130.200 ;
        RECT 99.800 127.900 100.200 130.200 ;
        RECT 102.200 127.900 102.600 130.200 ;
        RECT 103.800 127.900 104.200 130.200 ;
        RECT 104.600 127.900 105.000 130.200 ;
        RECT 108.600 126.900 109.000 130.200 ;
        RECT 111.800 127.900 112.200 130.200 ;
        RECT 114.200 127.900 114.600 130.200 ;
        RECT 117.200 127.900 117.600 130.200 ;
        RECT 120.600 126.900 121.000 130.200 ;
        RECT 121.400 127.900 121.800 130.200 ;
        RECT 123.000 127.900 123.400 130.200 ;
        RECT 124.600 127.900 125.000 130.200 ;
        RECT 126.200 127.900 126.600 130.200 ;
        RECT 127.800 127.900 128.200 130.200 ;
        RECT 128.600 126.900 129.000 130.200 ;
        RECT 132.600 127.900 133.000 130.200 ;
        RECT 135.300 128.900 135.800 130.200 ;
        RECT 137.000 128.900 137.400 130.200 ;
        RECT 139.800 128.000 140.200 130.200 ;
        RECT 142.200 128.300 142.600 130.200 ;
        RECT 146.200 127.900 146.600 130.200 ;
        RECT 147.800 127.700 148.200 130.200 ;
        RECT 150.400 127.500 150.800 130.200 ;
        RECT 152.400 127.500 152.800 130.200 ;
        RECT 155.000 127.700 155.400 130.200 ;
        RECT 158.200 127.900 158.600 130.200 ;
        RECT 159.800 127.900 160.200 130.200 ;
        RECT 163.300 128.000 163.700 130.200 ;
        RECT 165.400 128.900 165.800 130.200 ;
        RECT 167.000 128.900 167.400 130.200 ;
        RECT 168.600 128.300 169.000 130.200 ;
        RECT 171.000 127.900 171.400 130.200 ;
        RECT 172.600 127.900 173.000 130.200 ;
        RECT 175.000 127.900 175.400 130.200 ;
        RECT 176.600 127.900 177.000 130.200 ;
        RECT 177.400 127.900 177.800 130.200 ;
        RECT 179.000 127.900 179.400 130.200 ;
        RECT 180.100 127.900 180.500 130.200 ;
        RECT 182.200 128.900 182.600 130.200 ;
        RECT 183.000 127.900 183.400 130.200 ;
        RECT 186.200 127.900 186.600 130.200 ;
        RECT 188.900 128.900 189.400 130.200 ;
        RECT 190.600 128.900 191.000 130.200 ;
        RECT 193.400 128.000 193.800 130.200 ;
        RECT 195.000 127.900 195.400 130.200 ;
        RECT 196.600 127.900 197.000 130.200 ;
        RECT 198.200 127.900 198.600 130.200 ;
        RECT 199.800 127.900 200.200 130.200 ;
        RECT 201.400 127.900 201.800 130.200 ;
        RECT 203.000 127.900 203.400 130.200 ;
        RECT 205.400 128.300 205.800 130.200 ;
        RECT 210.200 127.700 210.600 130.200 ;
        RECT 212.800 127.500 213.200 130.200 ;
        RECT 215.000 128.900 215.400 130.200 ;
        RECT 216.600 127.900 217.000 130.200 ;
        RECT 219.300 128.900 219.800 130.200 ;
        RECT 221.000 128.900 221.400 130.200 ;
        RECT 223.800 128.000 224.200 130.200 ;
        RECT 226.200 127.700 226.600 130.200 ;
        RECT 228.800 127.500 229.200 130.200 ;
        RECT 230.200 128.900 230.600 130.200 ;
        RECT 232.600 128.000 233.000 130.200 ;
        RECT 235.400 128.900 235.800 130.200 ;
        RECT 237.000 128.900 237.500 130.200 ;
        RECT 239.800 127.900 240.200 130.200 ;
        RECT 241.400 127.900 241.800 130.200 ;
        RECT 243.000 127.900 243.400 130.200 ;
        RECT 245.400 128.300 245.800 130.200 ;
        RECT 249.400 127.900 249.800 130.200 ;
        RECT 251.000 128.000 251.400 130.200 ;
        RECT 253.800 128.900 254.200 130.200 ;
        RECT 255.400 128.900 255.900 130.200 ;
        RECT 258.200 127.900 258.600 130.200 ;
        RECT 260.600 127.900 261.000 130.200 ;
        RECT 262.200 126.900 262.600 130.200 ;
        RECT 0.600 110.800 1.000 113.100 ;
        RECT 2.200 110.800 2.600 113.100 ;
        RECT 3.800 110.800 4.200 113.100 ;
        RECT 5.400 110.800 5.800 113.100 ;
        RECT 7.000 110.800 7.400 113.100 ;
        RECT 8.600 110.800 9.000 113.100 ;
        RECT 11.300 110.800 11.800 112.100 ;
        RECT 13.000 110.800 13.400 112.100 ;
        RECT 15.800 110.800 16.200 113.000 ;
        RECT 18.200 110.800 18.600 112.700 ;
        RECT 22.200 110.800 22.600 113.100 ;
        RECT 23.800 110.800 24.200 113.300 ;
        RECT 26.400 110.800 26.800 113.500 ;
        RECT 28.100 110.800 28.500 113.100 ;
        RECT 30.200 110.800 30.600 112.100 ;
        RECT 31.000 110.800 31.400 112.100 ;
        RECT 32.600 110.800 33.000 112.100 ;
        RECT 33.400 110.800 33.800 113.100 ;
        RECT 35.000 110.800 35.400 113.100 ;
        RECT 37.400 110.800 37.800 113.300 ;
        RECT 40.000 110.800 40.400 113.500 ;
        RECT 42.200 110.800 42.600 112.100 ;
        RECT 43.800 110.800 44.200 113.000 ;
        RECT 46.600 110.800 47.000 112.100 ;
        RECT 48.200 110.800 48.700 112.100 ;
        RECT 51.000 110.800 51.400 113.100 ;
        RECT 52.900 110.800 53.300 113.100 ;
        RECT 55.000 110.800 55.400 112.100 ;
        RECT 57.400 110.800 57.800 112.100 ;
        RECT 59.000 110.800 59.400 112.100 ;
        RECT 60.600 110.800 61.000 113.100 ;
        RECT 63.300 110.800 63.800 112.100 ;
        RECT 65.000 110.800 65.400 112.100 ;
        RECT 67.800 110.800 68.200 113.000 ;
        RECT 70.200 110.800 70.600 112.700 ;
        RECT 72.600 110.800 73.000 113.100 ;
        RECT 75.800 110.800 76.200 113.300 ;
        RECT 78.400 110.800 78.800 113.500 ;
        RECT 80.600 110.800 81.000 113.300 ;
        RECT 83.200 110.800 83.600 113.500 ;
        RECT 85.400 110.800 85.800 112.700 ;
        RECT 89.400 110.800 89.800 113.100 ;
        RECT 91.000 110.800 91.400 113.300 ;
        RECT 93.600 110.800 94.000 113.500 ;
        RECT 95.800 110.800 96.200 113.000 ;
        RECT 98.600 110.800 99.000 112.100 ;
        RECT 100.200 110.800 100.700 112.100 ;
        RECT 103.000 110.800 103.400 113.100 ;
        RECT 107.000 110.800 107.400 113.100 ;
        RECT 109.700 110.800 110.200 112.100 ;
        RECT 111.400 110.800 111.800 112.100 ;
        RECT 114.200 110.800 114.600 113.000 ;
        RECT 116.600 110.800 117.000 113.100 ;
        RECT 119.300 110.800 119.800 112.100 ;
        RECT 121.000 110.800 121.400 112.100 ;
        RECT 123.800 110.800 124.200 113.000 ;
        RECT 126.200 110.800 126.600 112.700 ;
        RECT 129.400 110.800 129.800 112.700 ;
        RECT 133.400 110.800 133.800 113.100 ;
        RECT 135.000 110.800 135.400 113.100 ;
        RECT 137.700 110.800 138.200 112.100 ;
        RECT 139.400 110.800 139.800 112.100 ;
        RECT 142.200 110.800 142.600 113.000 ;
        RECT 143.800 110.800 144.200 112.100 ;
        RECT 145.400 110.800 145.800 112.100 ;
        RECT 146.200 110.800 146.600 112.100 ;
        RECT 147.800 110.800 148.200 112.100 ;
        RECT 148.600 110.800 149.000 112.100 ;
        RECT 150.200 110.800 150.600 112.100 ;
        RECT 151.800 110.800 152.200 113.300 ;
        RECT 154.400 110.800 154.800 113.500 ;
        RECT 155.800 110.800 156.200 113.100 ;
        RECT 161.400 110.800 161.800 112.700 ;
        RECT 163.800 110.800 164.200 113.000 ;
        RECT 166.600 110.800 167.000 112.100 ;
        RECT 168.200 110.800 168.700 112.100 ;
        RECT 171.000 110.800 171.400 113.100 ;
        RECT 172.600 110.800 173.000 113.100 ;
        RECT 174.200 110.800 174.600 113.100 ;
        RECT 175.800 110.800 176.200 113.100 ;
        RECT 177.400 110.800 177.800 113.100 ;
        RECT 179.000 110.800 179.400 113.100 ;
        RECT 179.800 110.800 180.200 113.100 ;
        RECT 181.400 110.800 181.800 113.100 ;
        RECT 183.000 110.800 183.400 113.100 ;
        RECT 184.600 110.800 185.000 113.100 ;
        RECT 186.200 110.800 186.600 113.100 ;
        RECT 187.000 110.800 187.400 113.100 ;
        RECT 189.400 110.800 189.800 113.000 ;
        RECT 192.200 110.800 192.600 112.100 ;
        RECT 193.800 110.800 194.300 112.100 ;
        RECT 196.600 110.800 197.000 113.100 ;
        RECT 198.200 110.800 198.600 113.100 ;
        RECT 199.800 110.800 200.200 113.100 ;
        RECT 201.400 110.800 201.800 113.100 ;
        RECT 203.000 110.800 203.400 113.100 ;
        RECT 205.200 110.800 205.600 113.500 ;
        RECT 207.800 110.800 208.200 113.300 ;
        RECT 211.000 110.800 211.400 113.100 ;
        RECT 213.400 110.800 213.800 112.100 ;
        RECT 215.000 110.800 215.400 112.100 ;
        RECT 215.800 110.800 216.200 112.100 ;
        RECT 217.900 110.800 218.300 113.100 ;
        RECT 219.800 110.800 220.200 113.100 ;
        RECT 222.500 110.800 223.000 112.100 ;
        RECT 224.200 110.800 224.600 112.100 ;
        RECT 227.000 110.800 227.400 113.000 ;
        RECT 228.600 110.800 229.000 113.100 ;
        RECT 232.600 110.800 233.000 112.700 ;
        RECT 234.500 110.800 234.900 113.100 ;
        RECT 236.600 110.800 237.000 112.100 ;
        RECT 238.200 110.800 238.600 113.100 ;
        RECT 239.800 110.800 240.200 113.100 ;
        RECT 240.600 110.800 241.000 112.100 ;
        RECT 242.200 110.800 242.600 112.100 ;
        RECT 243.300 110.800 243.700 113.100 ;
        RECT 245.400 110.800 245.800 112.100 ;
        RECT 247.000 110.800 247.400 113.000 ;
        RECT 249.800 110.800 250.200 112.100 ;
        RECT 251.400 110.800 251.900 112.100 ;
        RECT 254.200 110.800 254.600 113.100 ;
        RECT 256.600 110.800 257.000 113.100 ;
        RECT 259.300 110.800 259.800 112.100 ;
        RECT 261.000 110.800 261.400 112.100 ;
        RECT 263.800 110.800 264.200 113.000 ;
        RECT 0.200 110.200 265.400 110.800 ;
        RECT 0.600 107.900 1.000 110.200 ;
        RECT 2.200 107.900 2.600 110.200 ;
        RECT 3.800 107.900 4.200 110.200 ;
        RECT 5.400 107.900 5.800 110.200 ;
        RECT 8.100 108.900 8.600 110.200 ;
        RECT 9.800 108.900 10.200 110.200 ;
        RECT 12.600 108.000 13.000 110.200 ;
        RECT 14.500 107.900 14.900 110.200 ;
        RECT 16.600 108.900 17.000 110.200 ;
        RECT 17.400 108.900 17.800 110.200 ;
        RECT 19.000 108.900 19.400 110.200 ;
        RECT 20.600 107.900 21.000 110.200 ;
        RECT 23.300 108.900 23.800 110.200 ;
        RECT 25.000 108.900 25.400 110.200 ;
        RECT 27.800 108.000 28.200 110.200 ;
        RECT 30.200 107.700 30.600 110.200 ;
        RECT 32.800 107.500 33.200 110.200 ;
        RECT 34.200 108.900 34.600 110.200 ;
        RECT 36.400 107.500 36.800 110.200 ;
        RECT 39.000 107.700 39.400 110.200 ;
        RECT 41.200 107.500 41.600 110.200 ;
        RECT 43.800 107.700 44.200 110.200 ;
        RECT 46.200 108.000 46.600 110.200 ;
        RECT 49.000 108.900 49.400 110.200 ;
        RECT 50.600 108.900 51.100 110.200 ;
        RECT 53.400 107.900 53.800 110.200 ;
        RECT 56.600 107.900 57.000 110.200 ;
        RECT 58.200 107.900 58.600 110.200 ;
        RECT 60.600 107.900 61.000 110.200 ;
        RECT 63.300 108.900 63.800 110.200 ;
        RECT 65.000 108.900 65.400 110.200 ;
        RECT 67.800 108.000 68.200 110.200 ;
        RECT 70.200 108.300 70.600 110.200 ;
        RECT 74.200 107.900 74.600 110.200 ;
        RECT 75.800 107.900 76.200 110.200 ;
        RECT 78.500 108.900 79.000 110.200 ;
        RECT 80.200 108.900 80.600 110.200 ;
        RECT 83.000 108.000 83.400 110.200 ;
        RECT 84.600 108.900 85.000 110.200 ;
        RECT 86.200 108.900 86.600 110.200 ;
        RECT 87.000 108.900 87.400 110.200 ;
        RECT 89.100 107.900 89.500 110.200 ;
        RECT 91.000 107.900 91.400 110.200 ;
        RECT 93.700 108.900 94.200 110.200 ;
        RECT 95.400 108.900 95.800 110.200 ;
        RECT 98.200 108.000 98.600 110.200 ;
        RECT 99.800 107.900 100.200 110.200 ;
        RECT 101.400 107.900 101.800 110.200 ;
        RECT 103.300 107.900 103.700 110.200 ;
        RECT 105.400 108.900 105.800 110.200 ;
        RECT 107.800 108.900 108.200 110.200 ;
        RECT 109.400 108.900 109.800 110.200 ;
        RECT 111.000 107.700 111.400 110.200 ;
        RECT 113.600 107.500 114.000 110.200 ;
        RECT 115.800 108.900 116.200 110.200 ;
        RECT 116.600 107.900 117.000 110.200 ;
        RECT 118.200 107.900 118.600 110.200 ;
        RECT 119.800 107.900 120.200 110.200 ;
        RECT 121.400 107.900 121.800 110.200 ;
        RECT 123.000 107.900 123.400 110.200 ;
        RECT 123.800 107.900 124.200 110.200 ;
        RECT 125.400 107.900 125.800 110.200 ;
        RECT 128.600 107.900 129.000 110.200 ;
        RECT 130.200 107.700 130.600 110.200 ;
        RECT 132.800 107.500 133.200 110.200 ;
        RECT 135.000 107.700 135.400 110.200 ;
        RECT 137.600 107.500 138.000 110.200 ;
        RECT 139.000 107.900 139.400 110.200 ;
        RECT 140.600 107.900 141.000 110.200 ;
        RECT 142.200 107.900 142.600 110.200 ;
        RECT 143.000 108.900 143.400 110.200 ;
        RECT 144.600 108.900 145.000 110.200 ;
        RECT 146.200 108.100 146.600 110.200 ;
        RECT 147.800 108.900 148.200 110.200 ;
        RECT 148.600 108.900 149.000 110.200 ;
        RECT 150.200 108.900 150.600 110.200 ;
        RECT 151.800 107.900 152.200 110.200 ;
        RECT 153.400 107.900 153.800 110.200 ;
        RECT 154.800 107.500 155.200 110.200 ;
        RECT 157.400 107.700 157.800 110.200 ;
        RECT 160.800 107.900 161.200 110.200 ;
        RECT 163.800 107.900 164.200 110.200 ;
        RECT 164.600 107.900 165.000 110.200 ;
        RECT 167.200 107.900 167.600 110.200 ;
        RECT 170.200 107.900 170.600 110.200 ;
        RECT 171.800 108.000 172.200 110.200 ;
        RECT 174.600 108.900 175.000 110.200 ;
        RECT 176.200 108.900 176.700 110.200 ;
        RECT 179.000 107.900 179.400 110.200 ;
        RECT 180.600 107.900 181.000 110.200 ;
        RECT 184.600 108.300 185.000 110.200 ;
        RECT 186.500 107.900 186.900 110.200 ;
        RECT 188.600 108.900 189.000 110.200 ;
        RECT 189.400 108.900 189.800 110.200 ;
        RECT 191.000 108.900 191.400 110.200 ;
        RECT 192.600 108.000 193.000 110.200 ;
        RECT 195.400 108.900 195.800 110.200 ;
        RECT 197.000 108.900 197.500 110.200 ;
        RECT 199.800 107.900 200.200 110.200 ;
        RECT 202.200 107.900 202.600 110.200 ;
        RECT 203.800 107.900 204.200 110.200 ;
        RECT 204.600 107.900 205.000 110.200 ;
        RECT 207.000 108.900 207.400 110.200 ;
        RECT 208.600 108.900 209.000 110.200 ;
        RECT 211.000 108.900 211.400 110.200 ;
        RECT 212.600 108.900 213.000 110.200 ;
        RECT 214.200 108.000 214.600 110.200 ;
        RECT 217.000 108.900 217.400 110.200 ;
        RECT 218.600 108.900 219.100 110.200 ;
        RECT 221.400 107.900 221.800 110.200 ;
        RECT 224.600 107.900 225.000 110.200 ;
        RECT 225.400 108.900 225.800 110.200 ;
        RECT 227.000 108.900 227.400 110.200 ;
        RECT 227.800 107.900 228.200 110.200 ;
        RECT 230.200 107.900 230.600 110.200 ;
        RECT 233.400 108.000 233.800 110.200 ;
        RECT 236.200 108.900 236.600 110.200 ;
        RECT 237.800 108.900 238.300 110.200 ;
        RECT 240.600 107.900 241.000 110.200 ;
        RECT 242.500 107.900 242.900 110.200 ;
        RECT 244.600 108.900 245.000 110.200 ;
        RECT 245.400 107.900 245.800 110.200 ;
        RECT 247.000 107.900 247.400 110.200 ;
        RECT 248.600 107.900 249.000 110.200 ;
        RECT 250.200 107.900 250.600 110.200 ;
        RECT 251.800 107.900 252.200 110.200 ;
        RECT 253.400 107.900 253.800 110.200 ;
        RECT 256.100 108.900 256.600 110.200 ;
        RECT 257.800 108.900 258.200 110.200 ;
        RECT 260.600 108.000 261.000 110.200 ;
        RECT 262.200 108.900 262.600 110.200 ;
        RECT 263.800 108.900 264.200 110.200 ;
        RECT 1.400 90.800 1.800 93.100 ;
        RECT 4.100 90.800 4.600 92.100 ;
        RECT 5.800 90.800 6.200 92.100 ;
        RECT 8.600 90.800 9.000 93.000 ;
        RECT 10.200 90.800 10.600 93.100 ;
        RECT 14.200 90.800 14.600 92.700 ;
        RECT 16.600 90.800 17.000 93.300 ;
        RECT 19.200 90.800 19.600 93.500 ;
        RECT 20.600 90.800 21.000 93.100 ;
        RECT 23.800 90.800 24.200 93.100 ;
        RECT 26.500 90.800 27.000 92.100 ;
        RECT 28.200 90.800 28.600 92.100 ;
        RECT 31.000 90.800 31.400 93.000 ;
        RECT 32.600 90.800 33.000 93.100 ;
        RECT 36.600 90.800 37.000 92.700 ;
        RECT 38.200 90.800 38.600 92.100 ;
        RECT 39.800 90.800 40.200 92.100 ;
        RECT 41.200 90.800 41.600 93.500 ;
        RECT 43.800 90.800 44.200 93.300 ;
        RECT 46.200 90.800 46.600 92.700 ;
        RECT 50.200 90.800 50.600 93.100 ;
        RECT 53.400 90.800 53.800 93.000 ;
        RECT 56.200 90.800 56.600 92.100 ;
        RECT 57.800 90.800 58.300 92.100 ;
        RECT 60.600 90.800 61.000 93.100 ;
        RECT 63.800 90.800 64.200 92.700 ;
        RECT 66.200 90.800 66.600 93.000 ;
        RECT 69.000 90.800 69.400 92.100 ;
        RECT 70.600 90.800 71.100 92.100 ;
        RECT 73.400 90.800 73.800 93.100 ;
        RECT 75.000 90.800 75.400 93.100 ;
        RECT 76.600 90.800 77.000 93.100 ;
        RECT 78.200 90.800 78.600 93.100 ;
        RECT 79.800 90.800 80.200 93.100 ;
        RECT 81.400 90.800 81.800 93.100 ;
        RECT 83.000 90.800 83.400 93.300 ;
        RECT 85.600 90.800 86.000 93.500 ;
        RECT 87.600 90.800 88.000 93.500 ;
        RECT 90.200 90.800 90.600 93.300 ;
        RECT 92.600 90.800 93.000 93.300 ;
        RECT 95.200 90.800 95.600 93.500 ;
        RECT 97.400 90.800 97.800 92.100 ;
        RECT 99.000 90.800 99.400 93.000 ;
        RECT 101.800 90.800 102.200 92.100 ;
        RECT 103.400 90.800 103.900 92.100 ;
        RECT 106.200 90.800 106.600 93.100 ;
        RECT 110.200 90.800 110.600 93.300 ;
        RECT 112.800 90.800 113.200 93.500 ;
        RECT 115.000 90.800 115.400 92.100 ;
        RECT 116.600 90.800 117.000 93.100 ;
        RECT 119.300 90.800 119.800 92.100 ;
        RECT 121.000 90.800 121.400 92.100 ;
        RECT 123.800 90.800 124.200 93.000 ;
        RECT 125.400 90.800 125.800 92.100 ;
        RECT 127.000 90.800 127.400 92.100 ;
        RECT 128.600 90.800 129.000 92.100 ;
        RECT 130.200 90.800 130.600 93.300 ;
        RECT 132.800 90.800 133.200 93.500 ;
        RECT 135.000 90.800 135.400 93.100 ;
        RECT 136.600 90.800 137.000 93.100 ;
        RECT 137.700 90.800 138.100 93.100 ;
        RECT 139.800 90.800 140.200 92.100 ;
        RECT 141.400 90.800 141.800 93.100 ;
        RECT 144.100 90.800 144.600 92.100 ;
        RECT 145.800 90.800 146.200 92.100 ;
        RECT 148.600 90.800 149.000 93.000 ;
        RECT 150.200 90.800 150.600 92.100 ;
        RECT 151.800 90.800 152.200 92.100 ;
        RECT 153.200 90.800 153.600 93.500 ;
        RECT 155.800 90.800 156.200 93.300 ;
        RECT 159.000 90.800 159.400 93.100 ;
        RECT 162.200 90.800 162.600 93.100 ;
        RECT 164.900 90.800 165.400 92.100 ;
        RECT 166.600 90.800 167.000 92.100 ;
        RECT 169.400 90.800 169.800 93.000 ;
        RECT 171.000 90.800 171.400 93.100 ;
        RECT 175.000 90.800 175.400 92.700 ;
        RECT 177.200 90.800 177.600 93.500 ;
        RECT 179.800 90.800 180.200 93.300 ;
        RECT 182.000 90.800 182.400 93.500 ;
        RECT 184.600 90.800 185.000 93.300 ;
        RECT 186.800 90.800 187.200 93.500 ;
        RECT 189.400 90.800 189.800 93.300 ;
        RECT 191.000 90.800 191.400 93.100 ;
        RECT 193.400 90.800 193.800 93.100 ;
        RECT 195.000 90.800 195.400 93.100 ;
        RECT 196.600 90.800 197.000 93.100 ;
        RECT 198.200 90.800 198.600 93.100 ;
        RECT 199.800 90.800 200.200 93.100 ;
        RECT 201.400 90.800 201.800 93.100 ;
        RECT 203.800 90.800 204.200 93.100 ;
        RECT 205.400 90.800 205.800 93.100 ;
        RECT 208.600 90.800 209.000 93.000 ;
        RECT 211.400 90.800 211.800 92.100 ;
        RECT 213.000 90.800 213.500 92.100 ;
        RECT 215.800 90.800 216.200 93.100 ;
        RECT 217.400 90.800 217.800 93.100 ;
        RECT 220.600 90.800 221.000 93.100 ;
        RECT 223.300 90.800 223.800 92.100 ;
        RECT 225.000 90.800 225.400 92.100 ;
        RECT 227.800 90.800 228.200 93.000 ;
        RECT 229.400 90.800 229.800 93.100 ;
        RECT 231.000 90.800 231.400 93.100 ;
        RECT 232.600 90.800 233.000 92.100 ;
        RECT 234.700 90.800 235.100 93.100 ;
        RECT 235.800 90.800 236.200 93.100 ;
        RECT 239.000 90.800 239.400 92.100 ;
        RECT 240.600 90.800 241.000 93.000 ;
        RECT 243.400 90.800 243.800 92.100 ;
        RECT 245.000 90.800 245.500 92.100 ;
        RECT 247.800 90.800 248.200 93.100 ;
        RECT 249.400 90.800 249.800 93.100 ;
        RECT 252.100 90.800 252.500 93.100 ;
        RECT 254.200 90.800 254.600 92.100 ;
        RECT 255.800 90.800 256.200 93.100 ;
        RECT 257.400 90.800 257.800 92.100 ;
        RECT 259.000 90.800 259.400 92.100 ;
        RECT 259.800 90.800 260.200 93.100 ;
        RECT 263.000 90.800 263.400 93.100 ;
        RECT 0.200 90.200 265.400 90.800 ;
        RECT 1.400 87.900 1.800 90.200 ;
        RECT 4.100 88.900 4.600 90.200 ;
        RECT 5.800 88.900 6.200 90.200 ;
        RECT 8.600 88.000 9.000 90.200 ;
        RECT 10.200 88.900 10.600 90.200 ;
        RECT 12.400 87.500 12.800 90.200 ;
        RECT 15.000 87.700 15.400 90.200 ;
        RECT 17.400 88.000 17.800 90.200 ;
        RECT 20.200 88.900 20.600 90.200 ;
        RECT 21.800 88.900 22.300 90.200 ;
        RECT 24.600 87.900 25.000 90.200 ;
        RECT 27.800 88.300 28.200 90.200 ;
        RECT 30.200 87.900 30.600 90.200 ;
        RECT 32.900 88.900 33.400 90.200 ;
        RECT 34.600 88.900 35.000 90.200 ;
        RECT 37.400 88.000 37.800 90.200 ;
        RECT 39.000 88.900 39.400 90.200 ;
        RECT 41.100 87.900 41.500 90.200 ;
        RECT 42.800 87.500 43.200 90.200 ;
        RECT 45.400 87.700 45.800 90.200 ;
        RECT 47.800 87.700 48.200 90.200 ;
        RECT 50.400 87.500 50.800 90.200 ;
        RECT 52.400 87.500 52.800 90.200 ;
        RECT 55.000 87.700 55.400 90.200 ;
        RECT 58.200 87.900 58.600 90.200 ;
        RECT 61.400 88.000 61.800 90.200 ;
        RECT 64.200 88.900 64.600 90.200 ;
        RECT 65.800 88.900 66.300 90.200 ;
        RECT 68.600 87.900 69.000 90.200 ;
        RECT 71.800 87.900 72.200 90.200 ;
        RECT 74.200 88.300 74.600 90.200 ;
        RECT 75.800 87.900 76.200 90.200 ;
        RECT 78.800 87.900 79.200 90.200 ;
        RECT 80.400 87.500 80.800 90.200 ;
        RECT 83.000 87.700 83.400 90.200 ;
        RECT 84.600 87.900 85.000 90.200 ;
        RECT 86.200 87.900 86.600 90.200 ;
        RECT 87.800 87.900 88.200 90.200 ;
        RECT 89.400 87.900 89.800 90.200 ;
        RECT 91.000 87.900 91.400 90.200 ;
        RECT 91.800 88.900 92.200 90.200 ;
        RECT 94.200 88.000 94.600 90.200 ;
        RECT 97.000 88.900 97.400 90.200 ;
        RECT 98.600 88.900 99.100 90.200 ;
        RECT 101.400 87.900 101.800 90.200 ;
        RECT 103.800 87.700 104.200 90.200 ;
        RECT 106.400 87.500 106.800 90.200 ;
        RECT 110.200 87.900 110.600 90.200 ;
        RECT 112.900 88.900 113.400 90.200 ;
        RECT 114.600 88.900 115.000 90.200 ;
        RECT 117.400 88.000 117.800 90.200 ;
        RECT 119.000 88.900 119.400 90.200 ;
        RECT 121.200 87.500 121.600 90.200 ;
        RECT 123.800 87.700 124.200 90.200 ;
        RECT 126.200 87.900 126.600 90.200 ;
        RECT 128.900 88.900 129.400 90.200 ;
        RECT 130.600 88.900 131.000 90.200 ;
        RECT 133.400 88.000 133.800 90.200 ;
        RECT 135.000 88.900 135.400 90.200 ;
        RECT 137.200 87.500 137.600 90.200 ;
        RECT 139.800 87.700 140.200 90.200 ;
        RECT 142.000 87.500 142.400 90.200 ;
        RECT 144.600 87.700 145.000 90.200 ;
        RECT 147.500 88.000 147.900 90.200 ;
        RECT 149.400 87.900 149.800 90.200 ;
        RECT 151.800 88.000 152.200 90.200 ;
        RECT 154.600 88.900 155.000 90.200 ;
        RECT 156.200 88.900 156.700 90.200 ;
        RECT 159.000 87.900 159.400 90.200 ;
        RECT 163.800 88.300 164.200 90.200 ;
        RECT 166.000 87.500 166.400 90.200 ;
        RECT 168.600 87.700 169.000 90.200 ;
        RECT 171.000 87.900 171.400 90.200 ;
        RECT 173.700 88.900 174.200 90.200 ;
        RECT 175.400 88.900 175.800 90.200 ;
        RECT 178.200 88.000 178.600 90.200 ;
        RECT 181.400 88.300 181.800 90.200 ;
        RECT 184.600 88.300 185.000 90.200 ;
        RECT 187.000 88.300 187.400 90.200 ;
        RECT 190.200 88.000 190.600 90.200 ;
        RECT 193.000 88.900 193.400 90.200 ;
        RECT 194.600 88.900 195.100 90.200 ;
        RECT 197.400 87.900 197.800 90.200 ;
        RECT 199.000 87.900 199.400 90.200 ;
        RECT 200.600 87.900 201.000 90.200 ;
        RECT 202.200 87.900 202.600 90.200 ;
        RECT 203.800 87.900 204.200 90.200 ;
        RECT 205.400 87.900 205.800 90.200 ;
        RECT 206.200 87.900 206.600 90.200 ;
        RECT 207.800 87.900 208.200 90.200 ;
        RECT 209.400 87.900 209.800 90.200 ;
        RECT 213.400 88.300 213.800 90.200 ;
        RECT 216.600 88.300 217.000 90.200 ;
        RECT 218.500 87.900 218.900 90.200 ;
        RECT 220.600 88.900 221.000 90.200 ;
        RECT 223.000 88.300 223.400 90.200 ;
        RECT 224.600 87.900 225.000 90.200 ;
        RECT 226.200 87.900 226.600 90.200 ;
        RECT 228.600 88.300 229.000 90.200 ;
        RECT 231.800 87.900 232.200 90.200 ;
        RECT 234.500 88.900 235.000 90.200 ;
        RECT 236.200 88.900 236.600 90.200 ;
        RECT 239.000 88.000 239.400 90.200 ;
        RECT 240.600 87.900 241.000 90.200 ;
        RECT 242.200 87.900 242.600 90.200 ;
        RECT 243.800 87.900 244.200 90.200 ;
        RECT 245.400 87.900 245.800 90.200 ;
        RECT 247.000 87.900 247.400 90.200 ;
        RECT 247.800 87.900 248.200 90.200 ;
        RECT 249.400 87.900 249.800 90.200 ;
        RECT 251.000 87.900 251.400 90.200 ;
        RECT 252.600 87.900 253.000 90.200 ;
        RECT 254.200 87.900 254.600 90.200 ;
        RECT 255.000 88.900 255.400 90.200 ;
        RECT 257.100 87.900 257.500 90.200 ;
        RECT 258.200 87.900 258.600 90.200 ;
        RECT 259.800 87.900 260.200 90.200 ;
        RECT 261.400 87.900 261.800 90.200 ;
        RECT 263.000 87.900 263.400 90.200 ;
        RECT 264.600 87.900 265.000 90.200 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 4.100 70.800 4.600 72.100 ;
        RECT 5.800 70.800 6.200 72.100 ;
        RECT 8.600 70.800 9.000 73.000 ;
        RECT 10.200 70.800 10.600 73.100 ;
        RECT 14.200 70.800 14.600 72.700 ;
        RECT 16.600 70.800 17.000 73.100 ;
        RECT 19.300 70.800 19.800 72.100 ;
        RECT 21.000 70.800 21.400 72.100 ;
        RECT 23.800 70.800 24.200 73.000 ;
        RECT 25.400 70.800 25.800 72.100 ;
        RECT 27.000 70.800 27.400 72.100 ;
        RECT 27.800 70.800 28.200 72.100 ;
        RECT 29.900 70.800 30.300 73.100 ;
        RECT 31.800 70.800 32.200 73.100 ;
        RECT 34.500 70.800 35.000 72.100 ;
        RECT 36.200 70.800 36.600 72.100 ;
        RECT 39.000 70.800 39.400 73.000 ;
        RECT 41.400 70.800 41.800 73.300 ;
        RECT 44.000 70.800 44.400 73.500 ;
        RECT 46.200 70.800 46.600 72.100 ;
        RECT 47.800 70.800 48.200 73.000 ;
        RECT 50.600 70.800 51.000 72.100 ;
        RECT 52.200 70.800 52.700 72.100 ;
        RECT 55.000 70.800 55.400 73.100 ;
        RECT 59.000 70.800 59.400 73.000 ;
        RECT 61.800 70.800 62.200 72.100 ;
        RECT 63.400 70.800 63.900 72.100 ;
        RECT 66.200 70.800 66.600 73.100 ;
        RECT 67.800 70.800 68.200 73.100 ;
        RECT 71.800 70.800 72.200 72.700 ;
        RECT 74.200 70.800 74.600 73.300 ;
        RECT 76.800 70.800 77.200 73.500 ;
        RECT 79.000 70.800 79.400 72.100 ;
        RECT 80.600 70.800 81.000 73.000 ;
        RECT 83.400 70.800 83.800 72.100 ;
        RECT 85.000 70.800 85.500 72.100 ;
        RECT 87.800 70.800 88.200 73.100 ;
        RECT 89.400 70.800 89.800 73.100 ;
        RECT 92.900 70.800 93.300 73.000 ;
        RECT 95.000 70.800 95.400 73.100 ;
        RECT 97.400 70.800 97.800 73.100 ;
        RECT 99.000 70.800 99.400 73.100 ;
        RECT 101.400 70.800 101.800 73.100 ;
        RECT 103.000 70.800 103.400 73.100 ;
        RECT 104.600 70.800 105.000 72.700 ;
        RECT 110.200 70.800 110.600 73.100 ;
        RECT 111.800 70.800 112.200 73.100 ;
        RECT 114.500 70.800 115.000 72.100 ;
        RECT 116.200 70.800 116.600 72.100 ;
        RECT 119.000 70.800 119.400 73.000 ;
        RECT 120.600 70.800 121.000 73.100 ;
        RECT 122.200 70.800 122.600 73.100 ;
        RECT 123.800 70.800 124.200 73.100 ;
        RECT 125.400 70.800 125.800 73.100 ;
        RECT 127.000 70.800 127.400 73.100 ;
        RECT 127.800 70.800 128.200 73.100 ;
        RECT 131.000 70.800 131.400 73.100 ;
        RECT 133.700 70.800 134.200 72.100 ;
        RECT 135.400 70.800 135.800 72.100 ;
        RECT 138.200 70.800 138.600 73.000 ;
        RECT 139.800 70.800 140.200 72.100 ;
        RECT 141.400 70.800 141.800 72.100 ;
        RECT 143.000 70.800 143.400 73.300 ;
        RECT 145.600 70.800 146.000 73.500 ;
        RECT 147.800 70.800 148.200 73.100 ;
        RECT 150.500 70.800 151.000 72.100 ;
        RECT 152.200 70.800 152.600 72.100 ;
        RECT 155.000 70.800 155.400 73.000 ;
        RECT 158.200 70.800 158.600 73.100 ;
        RECT 161.900 70.800 162.300 73.000 ;
        RECT 165.400 70.800 165.800 72.700 ;
        RECT 167.600 70.800 168.000 73.500 ;
        RECT 170.200 70.800 170.600 73.300 ;
        RECT 172.600 70.800 173.000 73.300 ;
        RECT 175.200 70.800 175.600 73.500 ;
        RECT 177.400 70.800 177.800 73.000 ;
        RECT 180.200 70.800 180.600 72.100 ;
        RECT 181.800 70.800 182.300 72.100 ;
        RECT 184.600 70.800 185.000 73.100 ;
        RECT 186.200 70.800 186.600 72.100 ;
        RECT 187.800 70.800 188.200 72.100 ;
        RECT 188.600 70.800 189.000 72.100 ;
        RECT 190.700 70.800 191.100 73.100 ;
        RECT 192.400 70.800 192.800 73.500 ;
        RECT 195.000 70.800 195.400 73.300 ;
        RECT 198.200 70.800 198.600 72.700 ;
        RECT 199.800 70.800 200.200 73.100 ;
        RECT 201.400 70.800 201.800 73.100 ;
        RECT 203.000 70.800 203.400 73.100 ;
        RECT 204.600 70.800 205.000 73.100 ;
        RECT 206.200 70.800 206.600 73.100 ;
        RECT 210.200 70.800 210.600 72.700 ;
        RECT 212.600 70.800 213.000 73.100 ;
        RECT 215.300 70.800 215.800 72.100 ;
        RECT 217.000 70.800 217.400 72.100 ;
        RECT 219.800 70.800 220.200 73.000 ;
        RECT 223.000 70.800 223.400 72.700 ;
        RECT 224.600 70.800 225.000 73.100 ;
        RECT 227.800 70.800 228.200 72.700 ;
        RECT 231.800 70.800 232.200 72.700 ;
        RECT 234.200 70.800 234.600 73.000 ;
        RECT 237.000 70.800 237.400 72.100 ;
        RECT 238.600 70.800 239.100 72.100 ;
        RECT 241.400 70.800 241.800 73.100 ;
        RECT 243.300 70.800 243.700 73.100 ;
        RECT 245.400 70.800 245.800 72.100 ;
        RECT 247.000 70.800 247.400 73.000 ;
        RECT 249.800 70.800 250.200 72.100 ;
        RECT 251.400 70.800 251.900 72.100 ;
        RECT 254.200 70.800 254.600 73.100 ;
        RECT 256.600 70.800 257.000 73.000 ;
        RECT 259.400 70.800 259.800 72.100 ;
        RECT 261.000 70.800 261.500 72.100 ;
        RECT 263.800 70.800 264.200 73.100 ;
        RECT 0.200 70.200 265.400 70.800 ;
        RECT 0.600 67.900 1.000 70.200 ;
        RECT 2.200 67.900 2.600 70.200 ;
        RECT 3.800 67.900 4.200 70.200 ;
        RECT 5.400 67.900 5.800 70.200 ;
        RECT 7.000 67.900 7.400 70.200 ;
        RECT 7.800 67.900 8.200 70.200 ;
        RECT 9.400 67.900 9.800 70.200 ;
        RECT 11.000 67.900 11.400 70.200 ;
        RECT 12.600 67.900 13.000 70.200 ;
        RECT 14.200 67.900 14.600 70.200 ;
        RECT 15.800 67.900 16.200 70.200 ;
        RECT 18.500 68.900 19.000 70.200 ;
        RECT 20.200 68.900 20.600 70.200 ;
        RECT 23.000 68.000 23.400 70.200 ;
        RECT 24.900 67.900 25.300 70.200 ;
        RECT 27.000 68.900 27.400 70.200 ;
        RECT 27.800 68.900 28.200 70.200 ;
        RECT 29.400 68.900 29.800 70.200 ;
        RECT 30.800 67.500 31.200 70.200 ;
        RECT 33.400 67.700 33.800 70.200 ;
        RECT 35.800 67.700 36.200 70.200 ;
        RECT 38.400 67.500 38.800 70.200 ;
        RECT 40.600 68.900 41.000 70.200 ;
        RECT 42.000 67.500 42.400 70.200 ;
        RECT 44.600 67.700 45.000 70.200 ;
        RECT 46.800 67.500 47.200 70.200 ;
        RECT 49.400 67.700 49.800 70.200 ;
        RECT 51.200 67.900 51.600 70.200 ;
        RECT 54.200 67.900 54.600 70.200 ;
        RECT 57.400 67.700 57.800 70.200 ;
        RECT 60.000 67.500 60.400 70.200 ;
        RECT 62.000 67.500 62.400 70.200 ;
        RECT 64.600 67.700 65.000 70.200 ;
        RECT 67.000 67.700 67.400 70.200 ;
        RECT 69.600 67.500 70.000 70.200 ;
        RECT 71.800 67.700 72.200 70.200 ;
        RECT 74.400 67.500 74.800 70.200 ;
        RECT 76.000 67.900 76.400 70.200 ;
        RECT 79.000 67.900 79.400 70.200 ;
        RECT 80.600 67.900 81.000 70.200 ;
        RECT 83.300 68.900 83.800 70.200 ;
        RECT 85.000 68.900 85.400 70.200 ;
        RECT 87.800 68.000 88.200 70.200 ;
        RECT 90.200 67.700 90.600 70.200 ;
        RECT 92.800 67.500 93.200 70.200 ;
        RECT 95.000 68.900 95.400 70.200 ;
        RECT 95.800 67.900 96.200 70.200 ;
        RECT 98.800 67.900 99.200 70.200 ;
        RECT 100.400 67.500 100.800 70.200 ;
        RECT 103.000 67.700 103.400 70.200 ;
        RECT 107.000 67.700 107.400 70.200 ;
        RECT 109.600 67.500 110.000 70.200 ;
        RECT 112.600 67.900 113.000 70.200 ;
        RECT 114.200 67.700 114.600 70.200 ;
        RECT 116.800 67.500 117.200 70.200 ;
        RECT 119.000 67.700 119.400 70.200 ;
        RECT 121.600 67.500 122.000 70.200 ;
        RECT 123.000 67.900 123.400 70.200 ;
        RECT 125.400 67.900 125.800 70.200 ;
        RECT 128.400 67.900 128.800 70.200 ;
        RECT 129.400 67.900 129.800 70.200 ;
        RECT 132.400 67.900 132.800 70.200 ;
        RECT 134.000 67.500 134.400 70.200 ;
        RECT 136.600 67.700 137.000 70.200 ;
        RECT 138.500 67.900 138.900 70.200 ;
        RECT 140.600 68.900 141.000 70.200 ;
        RECT 141.400 67.900 141.800 70.200 ;
        RECT 143.000 67.900 143.400 70.200 ;
        RECT 144.600 67.900 145.000 70.200 ;
        RECT 146.200 67.900 146.600 70.200 ;
        RECT 147.800 67.900 148.200 70.200 ;
        RECT 149.400 68.300 149.800 70.200 ;
        RECT 152.400 67.500 152.800 70.200 ;
        RECT 155.000 67.700 155.400 70.200 ;
        RECT 159.800 67.900 160.200 70.200 ;
        RECT 160.600 67.900 161.000 70.200 ;
        RECT 163.600 67.900 164.000 70.200 ;
        RECT 164.600 67.900 165.000 70.200 ;
        RECT 167.200 67.900 167.600 70.200 ;
        RECT 170.200 67.900 170.600 70.200 ;
        RECT 171.800 68.000 172.200 70.200 ;
        RECT 174.600 68.900 175.000 70.200 ;
        RECT 176.200 68.900 176.700 70.200 ;
        RECT 179.000 67.900 179.400 70.200 ;
        RECT 180.600 67.900 181.000 70.200 ;
        RECT 184.600 68.300 185.000 70.200 ;
        RECT 186.200 67.900 186.600 70.200 ;
        RECT 187.800 67.900 188.200 70.200 ;
        RECT 189.400 67.900 189.800 70.200 ;
        RECT 191.000 67.900 191.400 70.200 ;
        RECT 192.600 67.900 193.000 70.200 ;
        RECT 194.200 67.900 194.600 70.200 ;
        RECT 195.800 67.900 196.200 70.200 ;
        RECT 196.800 67.900 197.200 70.200 ;
        RECT 199.800 67.900 200.200 70.200 ;
        RECT 202.200 67.900 202.600 70.200 ;
        RECT 203.000 67.900 203.400 70.200 ;
        RECT 206.000 67.900 206.400 70.200 ;
        RECT 208.800 67.900 209.200 70.200 ;
        RECT 211.800 67.900 212.200 70.200 ;
        RECT 214.200 67.900 214.600 70.200 ;
        RECT 215.000 67.900 215.400 70.200 ;
        RECT 218.000 67.900 218.400 70.200 ;
        RECT 219.600 67.500 220.000 70.200 ;
        RECT 222.200 67.700 222.600 70.200 ;
        RECT 224.600 67.700 225.000 70.200 ;
        RECT 227.200 67.500 227.600 70.200 ;
        RECT 229.400 67.900 229.800 70.200 ;
        RECT 232.100 68.900 232.600 70.200 ;
        RECT 233.800 68.900 234.200 70.200 ;
        RECT 236.600 68.000 237.000 70.200 ;
        RECT 238.800 67.500 239.200 70.200 ;
        RECT 241.400 67.700 241.800 70.200 ;
        RECT 243.800 67.700 244.200 70.200 ;
        RECT 246.400 67.500 246.800 70.200 ;
        RECT 248.600 67.700 249.000 70.200 ;
        RECT 251.200 67.500 251.600 70.200 ;
        RECT 254.200 68.300 254.600 70.200 ;
        RECT 256.600 68.000 257.000 70.200 ;
        RECT 259.400 68.900 259.800 70.200 ;
        RECT 261.000 68.900 261.500 70.200 ;
        RECT 263.800 67.900 264.200 70.200 ;
        RECT 0.600 50.800 1.000 53.100 ;
        RECT 2.200 50.800 2.600 53.100 ;
        RECT 3.800 50.800 4.200 53.100 ;
        RECT 5.400 50.800 5.800 53.100 ;
        RECT 7.000 50.800 7.400 53.100 ;
        RECT 7.800 50.800 8.200 53.100 ;
        RECT 9.400 50.800 9.800 53.100 ;
        RECT 11.000 50.800 11.400 53.100 ;
        RECT 12.600 50.800 13.000 53.100 ;
        RECT 14.200 50.800 14.600 53.100 ;
        RECT 15.800 50.800 16.200 53.300 ;
        RECT 18.400 50.800 18.800 53.500 ;
        RECT 20.600 50.800 21.000 53.100 ;
        RECT 23.300 50.800 23.800 52.100 ;
        RECT 25.000 50.800 25.400 52.100 ;
        RECT 27.800 50.800 28.200 53.000 ;
        RECT 30.200 50.800 30.600 53.300 ;
        RECT 32.800 50.800 33.200 53.500 ;
        RECT 35.000 50.800 35.400 52.100 ;
        RECT 35.800 50.800 36.200 52.100 ;
        RECT 38.000 50.800 38.400 53.500 ;
        RECT 40.600 50.800 41.000 53.300 ;
        RECT 43.000 50.800 43.400 53.300 ;
        RECT 45.600 50.800 46.000 53.500 ;
        RECT 47.800 50.800 48.200 53.100 ;
        RECT 50.500 50.800 51.000 52.100 ;
        RECT 52.200 50.800 52.600 52.100 ;
        RECT 55.000 50.800 55.400 53.000 ;
        RECT 58.500 50.800 58.900 53.100 ;
        RECT 60.600 50.800 61.000 52.100 ;
        RECT 61.400 50.800 61.800 52.100 ;
        RECT 63.000 50.800 63.400 52.100 ;
        RECT 64.400 50.800 64.800 53.500 ;
        RECT 67.000 50.800 67.400 53.300 ;
        RECT 69.400 50.800 69.800 52.700 ;
        RECT 71.800 50.800 72.200 53.100 ;
        RECT 75.000 50.800 75.400 53.000 ;
        RECT 77.800 50.800 78.200 52.100 ;
        RECT 79.400 50.800 79.900 52.100 ;
        RECT 82.200 50.800 82.600 53.100 ;
        RECT 84.600 50.800 85.000 52.700 ;
        RECT 87.000 50.800 87.400 53.100 ;
        RECT 90.200 50.800 90.600 53.300 ;
        RECT 92.800 50.800 93.200 53.500 ;
        RECT 95.000 50.800 95.400 53.300 ;
        RECT 97.600 50.800 98.000 53.500 ;
        RECT 99.800 50.800 100.200 53.100 ;
        RECT 102.500 50.800 103.000 52.100 ;
        RECT 104.200 50.800 104.600 52.100 ;
        RECT 107.000 50.800 107.400 53.000 ;
        RECT 111.800 50.800 112.200 52.700 ;
        RECT 113.400 50.800 113.800 52.100 ;
        RECT 115.000 50.800 115.400 52.100 ;
        RECT 115.800 50.800 116.200 52.100 ;
        RECT 117.900 50.800 118.300 53.100 ;
        RECT 119.800 50.800 120.200 53.100 ;
        RECT 122.500 50.800 123.000 52.100 ;
        RECT 124.200 50.800 124.600 52.100 ;
        RECT 127.000 50.800 127.400 53.000 ;
        RECT 128.600 50.800 129.000 53.100 ;
        RECT 132.600 50.800 133.000 52.700 ;
        RECT 134.800 50.800 135.200 53.500 ;
        RECT 137.400 50.800 137.800 53.300 ;
        RECT 139.800 50.800 140.200 53.300 ;
        RECT 142.400 50.800 142.800 53.500 ;
        RECT 144.600 50.800 145.000 53.300 ;
        RECT 147.200 50.800 147.600 53.500 ;
        RECT 149.400 50.800 149.800 53.100 ;
        RECT 152.100 50.800 152.600 52.100 ;
        RECT 153.800 50.800 154.200 52.100 ;
        RECT 156.600 50.800 157.000 53.000 ;
        RECT 160.600 50.800 161.000 52.700 ;
        RECT 164.600 50.800 165.000 53.100 ;
        RECT 166.000 50.800 166.400 53.500 ;
        RECT 168.600 50.800 169.000 53.300 ;
        RECT 170.800 50.800 171.200 53.500 ;
        RECT 173.400 50.800 173.800 53.300 ;
        RECT 175.000 50.800 175.400 52.100 ;
        RECT 176.600 50.800 177.000 52.100 ;
        RECT 177.400 50.800 177.800 52.100 ;
        RECT 179.500 50.800 179.900 53.100 ;
        RECT 181.400 50.800 181.800 53.000 ;
        RECT 184.200 50.800 184.600 52.100 ;
        RECT 185.800 50.800 186.300 52.100 ;
        RECT 188.600 50.800 189.000 53.100 ;
        RECT 191.000 50.800 191.400 53.300 ;
        RECT 193.600 50.800 194.000 53.500 ;
        RECT 195.800 50.800 196.200 52.100 ;
        RECT 197.400 50.800 197.800 53.300 ;
        RECT 200.000 50.800 200.400 53.500 ;
        RECT 202.200 50.800 202.600 53.300 ;
        RECT 204.800 50.800 205.200 53.500 ;
        RECT 207.000 50.800 207.400 52.700 ;
        RECT 211.800 50.800 212.200 53.100 ;
        RECT 214.500 50.800 215.000 52.100 ;
        RECT 216.200 50.800 216.600 52.100 ;
        RECT 219.000 50.800 219.400 53.000 ;
        RECT 221.200 50.800 221.600 53.500 ;
        RECT 223.800 50.800 224.200 53.300 ;
        RECT 226.200 50.800 226.600 53.300 ;
        RECT 228.800 50.800 229.200 53.500 ;
        RECT 231.000 50.800 231.400 53.300 ;
        RECT 233.600 50.800 234.000 53.500 ;
        RECT 235.800 50.800 236.200 52.700 ;
        RECT 239.000 50.800 239.400 53.100 ;
        RECT 241.700 50.800 242.200 52.100 ;
        RECT 243.400 50.800 243.800 52.100 ;
        RECT 246.200 50.800 246.600 53.000 ;
        RECT 248.600 50.800 249.000 52.700 ;
        RECT 252.600 50.800 253.000 53.100 ;
        RECT 254.200 50.800 254.600 53.300 ;
        RECT 256.800 50.800 257.200 53.500 ;
        RECT 258.200 50.800 258.600 53.100 ;
        RECT 261.400 50.800 261.800 52.700 ;
        RECT 0.200 50.200 265.400 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 4.100 48.900 4.600 50.200 ;
        RECT 5.800 48.900 6.200 50.200 ;
        RECT 8.600 48.000 9.000 50.200 ;
        RECT 10.200 48.900 10.600 50.200 ;
        RECT 12.400 47.500 12.800 50.200 ;
        RECT 15.000 47.700 15.400 50.200 ;
        RECT 17.400 48.000 17.800 50.200 ;
        RECT 20.200 48.900 20.600 50.200 ;
        RECT 21.800 48.900 22.300 50.200 ;
        RECT 24.600 47.900 25.000 50.200 ;
        RECT 26.200 48.900 26.600 50.200 ;
        RECT 28.400 47.500 28.800 50.200 ;
        RECT 31.000 47.700 31.400 50.200 ;
        RECT 33.400 48.000 33.800 50.200 ;
        RECT 36.200 48.900 36.600 50.200 ;
        RECT 37.800 48.900 38.300 50.200 ;
        RECT 40.600 47.900 41.000 50.200 ;
        RECT 43.000 48.000 43.400 50.200 ;
        RECT 45.800 48.900 46.200 50.200 ;
        RECT 47.400 48.900 47.900 50.200 ;
        RECT 50.200 47.900 50.600 50.200 ;
        RECT 51.800 47.900 52.200 50.200 ;
        RECT 57.400 48.300 57.800 50.200 ;
        RECT 59.000 47.900 59.400 50.200 ;
        RECT 60.600 47.900 61.000 50.200 ;
        RECT 63.000 48.000 63.400 50.200 ;
        RECT 65.800 48.900 66.200 50.200 ;
        RECT 67.400 48.900 67.900 50.200 ;
        RECT 70.200 47.900 70.600 50.200 ;
        RECT 72.600 48.000 73.000 50.200 ;
        RECT 75.400 48.900 75.800 50.200 ;
        RECT 77.000 48.900 77.500 50.200 ;
        RECT 79.800 47.900 80.200 50.200 ;
        RECT 82.200 48.300 82.600 50.200 ;
        RECT 86.200 47.900 86.600 50.200 ;
        RECT 87.800 47.900 88.200 50.200 ;
        RECT 90.500 48.900 91.000 50.200 ;
        RECT 92.200 48.900 92.600 50.200 ;
        RECT 95.000 48.000 95.400 50.200 ;
        RECT 96.600 47.900 97.000 50.200 ;
        RECT 100.600 48.300 101.000 50.200 ;
        RECT 104.600 48.000 105.000 50.200 ;
        RECT 107.400 48.900 107.800 50.200 ;
        RECT 109.000 48.900 109.500 50.200 ;
        RECT 111.800 47.900 112.200 50.200 ;
        RECT 114.200 47.900 114.600 50.200 ;
        RECT 116.900 48.900 117.400 50.200 ;
        RECT 118.600 48.900 119.000 50.200 ;
        RECT 121.400 48.000 121.800 50.200 ;
        RECT 124.600 48.300 125.000 50.200 ;
        RECT 127.800 48.300 128.200 50.200 ;
        RECT 130.200 47.900 130.600 50.200 ;
        RECT 132.900 48.900 133.400 50.200 ;
        RECT 134.600 48.900 135.000 50.200 ;
        RECT 137.400 48.000 137.800 50.200 ;
        RECT 139.800 48.300 140.200 50.200 ;
        RECT 143.800 48.300 144.200 50.200 ;
        RECT 146.200 47.700 146.600 50.200 ;
        RECT 148.800 47.500 149.200 50.200 ;
        RECT 151.000 48.900 151.400 50.200 ;
        RECT 151.800 47.900 152.200 50.200 ;
        RECT 155.800 48.300 156.200 50.200 ;
        RECT 159.800 48.000 160.200 50.200 ;
        RECT 162.600 48.900 163.000 50.200 ;
        RECT 164.200 48.900 164.700 50.200 ;
        RECT 167.000 47.900 167.400 50.200 ;
        RECT 169.400 47.900 169.800 50.200 ;
        RECT 171.000 47.900 171.400 50.200 ;
        RECT 172.600 48.300 173.000 50.200 ;
        RECT 176.600 47.900 177.000 50.200 ;
        RECT 178.200 48.000 178.600 50.200 ;
        RECT 181.000 48.900 181.400 50.200 ;
        RECT 182.600 48.900 183.100 50.200 ;
        RECT 185.400 47.900 185.800 50.200 ;
        RECT 187.800 47.900 188.200 50.200 ;
        RECT 190.500 48.900 191.000 50.200 ;
        RECT 192.200 48.900 192.600 50.200 ;
        RECT 195.000 48.000 195.400 50.200 ;
        RECT 197.400 47.900 197.800 50.200 ;
        RECT 200.100 48.900 200.600 50.200 ;
        RECT 201.800 48.900 202.200 50.200 ;
        RECT 204.600 48.000 205.000 50.200 ;
        RECT 206.200 48.900 206.600 50.200 ;
        RECT 207.800 48.900 208.200 50.200 ;
        RECT 210.200 48.900 210.600 50.200 ;
        RECT 212.300 47.900 212.700 50.200 ;
        RECT 214.200 47.700 214.600 50.200 ;
        RECT 216.800 47.500 217.200 50.200 ;
        RECT 219.800 47.900 220.200 50.200 ;
        RECT 221.400 47.700 221.800 50.200 ;
        RECT 224.000 47.500 224.400 50.200 ;
        RECT 226.200 47.700 226.600 50.200 ;
        RECT 228.800 47.500 229.200 50.200 ;
        RECT 231.000 48.300 231.400 50.200 ;
        RECT 235.000 47.900 235.400 50.200 ;
        RECT 235.800 47.900 236.200 50.200 ;
        RECT 239.000 48.000 239.400 50.200 ;
        RECT 241.800 48.900 242.200 50.200 ;
        RECT 243.400 48.900 243.900 50.200 ;
        RECT 246.200 47.900 246.600 50.200 ;
        RECT 247.800 48.900 248.200 50.200 ;
        RECT 249.400 48.900 249.800 50.200 ;
        RECT 251.000 47.900 251.400 50.200 ;
        RECT 253.700 48.900 254.200 50.200 ;
        RECT 255.400 48.900 255.800 50.200 ;
        RECT 258.200 48.000 258.600 50.200 ;
        RECT 259.800 47.900 260.200 50.200 ;
        RECT 263.000 48.300 263.400 50.200 ;
        RECT 0.900 30.800 1.300 33.100 ;
        RECT 3.000 30.800 3.400 32.100 ;
        RECT 3.800 30.800 4.200 32.100 ;
        RECT 5.400 30.800 5.800 32.100 ;
        RECT 7.000 30.800 7.400 33.300 ;
        RECT 9.600 30.800 10.000 33.500 ;
        RECT 11.000 30.800 11.400 32.100 ;
        RECT 13.400 30.800 13.800 33.000 ;
        RECT 16.200 30.800 16.600 32.100 ;
        RECT 17.800 30.800 18.300 32.100 ;
        RECT 20.600 30.800 21.000 33.100 ;
        RECT 22.800 30.800 23.200 33.500 ;
        RECT 25.400 30.800 25.800 33.300 ;
        RECT 27.800 30.800 28.200 32.700 ;
        RECT 31.800 30.800 32.200 33.100 ;
        RECT 33.400 30.800 33.800 32.700 ;
        RECT 37.400 30.800 37.800 33.100 ;
        RECT 39.000 30.800 39.400 33.300 ;
        RECT 41.600 30.800 42.000 33.500 ;
        RECT 43.000 30.800 43.400 32.100 ;
        RECT 44.600 30.800 45.000 32.100 ;
        RECT 46.200 30.800 46.600 33.100 ;
        RECT 48.900 30.800 49.400 32.100 ;
        RECT 50.600 30.800 51.000 32.100 ;
        RECT 53.400 30.800 53.800 33.000 ;
        RECT 57.200 30.800 57.600 33.500 ;
        RECT 59.800 30.800 60.200 33.300 ;
        RECT 61.400 30.800 61.800 33.100 ;
        RECT 64.600 30.800 65.000 33.300 ;
        RECT 67.200 30.800 67.600 33.500 ;
        RECT 69.400 30.800 69.800 32.700 ;
        RECT 73.400 30.800 73.800 33.100 ;
        RECT 75.000 30.800 75.400 33.100 ;
        RECT 77.700 30.800 78.200 32.100 ;
        RECT 79.400 30.800 79.800 32.100 ;
        RECT 82.200 30.800 82.600 33.000 ;
        RECT 84.600 30.800 85.000 33.300 ;
        RECT 87.200 30.800 87.600 33.500 ;
        RECT 89.200 30.800 89.600 33.500 ;
        RECT 91.800 30.800 92.200 33.300 ;
        RECT 94.200 30.800 94.600 33.100 ;
        RECT 96.900 30.800 97.400 32.100 ;
        RECT 98.600 30.800 99.000 32.100 ;
        RECT 101.400 30.800 101.800 33.000 ;
        RECT 103.000 30.800 103.400 32.100 ;
        RECT 106.800 30.800 107.200 33.500 ;
        RECT 109.400 30.800 109.800 33.300 ;
        RECT 111.000 30.800 111.400 33.100 ;
        RECT 112.600 30.800 113.000 33.100 ;
        RECT 114.200 30.800 114.600 33.100 ;
        RECT 115.800 30.800 116.200 33.100 ;
        RECT 117.400 30.800 117.800 33.100 ;
        RECT 118.200 30.800 118.600 33.100 ;
        RECT 119.800 30.800 120.200 33.100 ;
        RECT 121.400 30.800 121.800 33.100 ;
        RECT 123.000 30.800 123.400 33.100 ;
        RECT 124.600 30.800 125.000 33.100 ;
        RECT 126.200 30.800 126.600 33.300 ;
        RECT 128.800 30.800 129.200 33.500 ;
        RECT 131.000 30.800 131.400 33.100 ;
        RECT 132.600 30.800 133.000 33.100 ;
        RECT 134.200 30.800 134.600 33.300 ;
        RECT 136.800 30.800 137.200 33.500 ;
        RECT 138.200 30.800 138.600 32.100 ;
        RECT 139.800 30.800 140.200 32.100 ;
        RECT 140.600 30.800 141.000 32.100 ;
        RECT 142.700 30.800 143.100 33.100 ;
        RECT 144.600 30.800 145.000 33.100 ;
        RECT 147.300 30.800 147.800 32.100 ;
        RECT 149.000 30.800 149.400 32.100 ;
        RECT 151.800 30.800 152.200 33.000 ;
        RECT 153.400 30.800 153.800 32.100 ;
        RECT 155.000 30.800 155.400 32.900 ;
        RECT 159.000 30.800 159.400 33.100 ;
        RECT 161.700 30.800 162.200 32.100 ;
        RECT 163.400 30.800 163.800 32.100 ;
        RECT 166.200 30.800 166.600 33.000 ;
        RECT 168.600 30.800 169.000 33.300 ;
        RECT 171.200 30.800 171.600 33.500 ;
        RECT 172.600 30.800 173.000 32.100 ;
        RECT 174.200 30.800 174.600 32.100 ;
        RECT 175.000 30.800 175.400 32.100 ;
        RECT 177.100 30.800 177.500 33.100 ;
        RECT 179.000 30.800 179.400 33.100 ;
        RECT 181.700 30.800 182.200 32.100 ;
        RECT 183.400 30.800 183.800 32.100 ;
        RECT 186.200 30.800 186.600 33.000 ;
        RECT 188.600 30.800 189.000 33.300 ;
        RECT 191.200 30.800 191.600 33.500 ;
        RECT 193.400 30.800 193.800 32.100 ;
        RECT 195.000 30.800 195.400 33.300 ;
        RECT 197.600 30.800 198.000 33.500 ;
        RECT 199.600 30.800 200.000 33.500 ;
        RECT 202.200 30.800 202.600 33.300 ;
        RECT 204.100 30.800 204.500 33.100 ;
        RECT 206.200 30.800 206.600 32.100 ;
        RECT 207.000 30.800 207.400 32.100 ;
        RECT 208.600 30.800 209.000 32.100 ;
        RECT 211.600 30.800 212.000 33.500 ;
        RECT 214.200 30.800 214.600 33.300 ;
        RECT 216.400 30.800 216.800 33.500 ;
        RECT 219.000 30.800 219.400 33.300 ;
        RECT 220.900 30.800 221.300 33.100 ;
        RECT 223.000 30.800 223.400 32.100 ;
        RECT 223.800 30.800 224.200 32.100 ;
        RECT 225.400 30.800 225.800 32.100 ;
        RECT 227.000 30.800 227.400 33.300 ;
        RECT 229.600 30.800 230.000 33.500 ;
        RECT 231.000 30.800 231.400 33.100 ;
        RECT 235.000 30.800 235.400 32.700 ;
        RECT 237.400 30.800 237.800 33.000 ;
        RECT 240.200 30.800 240.600 32.100 ;
        RECT 241.800 30.800 242.300 32.100 ;
        RECT 244.600 30.800 245.000 33.100 ;
        RECT 247.000 30.800 247.400 32.700 ;
        RECT 251.000 30.800 251.400 33.100 ;
        RECT 252.600 30.800 253.000 33.000 ;
        RECT 255.400 30.800 255.800 32.100 ;
        RECT 257.000 30.800 257.500 32.100 ;
        RECT 259.800 30.800 260.200 33.100 ;
        RECT 262.200 30.800 262.600 32.700 ;
        RECT 0.200 30.200 265.400 30.800 ;
        RECT 1.400 27.900 1.800 30.200 ;
        RECT 4.100 28.900 4.600 30.200 ;
        RECT 5.800 28.900 6.200 30.200 ;
        RECT 8.600 28.000 9.000 30.200 ;
        RECT 10.200 27.900 10.600 30.200 ;
        RECT 11.800 27.900 12.200 30.200 ;
        RECT 13.400 27.900 13.800 30.200 ;
        RECT 15.000 27.900 15.400 30.200 ;
        RECT 16.600 27.900 17.000 30.200 ;
        RECT 18.200 27.700 18.600 30.200 ;
        RECT 20.800 27.500 21.200 30.200 ;
        RECT 22.800 27.500 23.200 30.200 ;
        RECT 25.400 27.700 25.800 30.200 ;
        RECT 27.800 27.900 28.200 30.200 ;
        RECT 30.500 28.900 31.000 30.200 ;
        RECT 32.200 28.900 32.600 30.200 ;
        RECT 35.000 28.000 35.400 30.200 ;
        RECT 37.400 27.900 37.800 30.200 ;
        RECT 40.100 28.900 40.600 30.200 ;
        RECT 41.800 28.900 42.200 30.200 ;
        RECT 44.600 28.000 45.000 30.200 ;
        RECT 46.200 28.900 46.600 30.200 ;
        RECT 48.300 27.900 48.700 30.200 ;
        RECT 50.200 27.900 50.600 30.200 ;
        RECT 52.900 28.900 53.400 30.200 ;
        RECT 54.600 28.900 55.000 30.200 ;
        RECT 57.400 28.000 57.800 30.200 ;
        RECT 61.400 28.300 61.800 30.200 ;
        RECT 64.600 27.900 65.000 30.200 ;
        RECT 66.200 27.900 66.600 30.200 ;
        RECT 67.800 28.300 68.200 30.200 ;
        RECT 71.800 27.900 72.200 30.200 ;
        RECT 73.400 28.000 73.800 30.200 ;
        RECT 76.200 28.900 76.600 30.200 ;
        RECT 77.800 28.900 78.300 30.200 ;
        RECT 80.600 27.900 81.000 30.200 ;
        RECT 82.800 27.500 83.200 30.200 ;
        RECT 85.400 27.700 85.800 30.200 ;
        RECT 87.000 28.900 87.400 30.200 ;
        RECT 89.200 27.500 89.600 30.200 ;
        RECT 91.800 27.700 92.200 30.200 ;
        RECT 94.200 27.700 94.600 30.200 ;
        RECT 96.800 27.500 97.200 30.200 ;
        RECT 98.200 27.900 98.600 30.200 ;
        RECT 99.800 27.900 100.200 30.200 ;
        RECT 102.200 28.300 102.600 30.200 ;
        RECT 106.200 27.900 106.600 30.200 ;
        RECT 109.400 28.000 109.800 30.200 ;
        RECT 112.200 28.900 112.600 30.200 ;
        RECT 113.800 28.900 114.300 30.200 ;
        RECT 116.600 27.900 117.000 30.200 ;
        RECT 119.000 27.700 119.400 30.200 ;
        RECT 121.600 27.500 122.000 30.200 ;
        RECT 123.800 27.700 124.200 30.200 ;
        RECT 126.400 27.500 126.800 30.200 ;
        RECT 128.600 28.900 129.000 30.200 ;
        RECT 130.200 28.000 130.600 30.200 ;
        RECT 133.000 28.900 133.400 30.200 ;
        RECT 134.600 28.900 135.100 30.200 ;
        RECT 137.400 27.900 137.800 30.200 ;
        RECT 139.800 28.000 140.200 30.200 ;
        RECT 142.600 28.900 143.000 30.200 ;
        RECT 144.200 28.900 144.700 30.200 ;
        RECT 147.000 27.900 147.400 30.200 ;
        RECT 149.400 28.300 149.800 30.200 ;
        RECT 153.400 27.900 153.800 30.200 ;
        RECT 156.600 27.900 157.000 30.200 ;
        RECT 159.300 28.900 159.800 30.200 ;
        RECT 161.000 28.900 161.400 30.200 ;
        RECT 163.800 28.000 164.200 30.200 ;
        RECT 166.200 28.300 166.600 30.200 ;
        RECT 170.200 27.900 170.600 30.200 ;
        RECT 171.800 28.000 172.200 30.200 ;
        RECT 174.600 28.900 175.000 30.200 ;
        RECT 176.200 28.900 176.700 30.200 ;
        RECT 179.000 27.900 179.400 30.200 ;
        RECT 180.600 27.900 181.000 30.200 ;
        RECT 182.200 27.900 182.600 30.200 ;
        RECT 184.600 27.700 185.000 30.200 ;
        RECT 187.200 27.500 187.600 30.200 ;
        RECT 189.400 28.900 189.800 30.200 ;
        RECT 191.000 28.000 191.400 30.200 ;
        RECT 193.800 28.900 194.200 30.200 ;
        RECT 195.400 28.900 195.900 30.200 ;
        RECT 198.200 27.900 198.600 30.200 ;
        RECT 200.600 28.300 201.000 30.200 ;
        RECT 204.600 28.300 205.000 30.200 ;
        RECT 208.600 27.900 209.000 30.200 ;
        RECT 211.300 28.900 211.800 30.200 ;
        RECT 213.000 28.900 213.400 30.200 ;
        RECT 215.800 28.000 216.200 30.200 ;
        RECT 218.200 27.700 218.600 30.200 ;
        RECT 220.800 27.500 221.200 30.200 ;
        RECT 223.000 28.000 223.400 30.200 ;
        RECT 225.800 28.900 226.200 30.200 ;
        RECT 227.400 28.900 227.900 30.200 ;
        RECT 230.200 27.900 230.600 30.200 ;
        RECT 232.600 28.900 233.000 30.200 ;
        RECT 234.200 28.000 234.600 30.200 ;
        RECT 237.000 28.900 237.400 30.200 ;
        RECT 238.600 28.900 239.100 30.200 ;
        RECT 241.400 27.900 241.800 30.200 ;
        RECT 243.000 27.900 243.400 30.200 ;
        RECT 247.000 28.300 247.400 30.200 ;
        RECT 249.400 27.700 249.800 30.200 ;
        RECT 252.000 27.500 252.400 30.200 ;
        RECT 254.200 28.000 254.600 30.200 ;
        RECT 257.000 28.900 257.400 30.200 ;
        RECT 258.600 28.900 259.100 30.200 ;
        RECT 261.400 27.900 261.800 30.200 ;
        RECT 1.400 10.800 1.800 13.000 ;
        RECT 4.200 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.300 12.100 ;
        RECT 8.600 10.800 9.000 13.100 ;
        RECT 11.800 10.800 12.200 12.700 ;
        RECT 14.200 10.800 14.600 12.700 ;
        RECT 18.200 10.800 18.600 13.100 ;
        RECT 19.800 10.800 20.200 13.300 ;
        RECT 22.400 10.800 22.800 13.500 ;
        RECT 24.600 10.800 25.000 13.000 ;
        RECT 27.400 10.800 27.800 12.100 ;
        RECT 29.000 10.800 29.500 12.100 ;
        RECT 31.800 10.800 32.200 13.100 ;
        RECT 33.400 10.800 33.800 12.100 ;
        RECT 35.000 10.800 35.400 12.100 ;
        RECT 35.800 10.800 36.200 12.100 ;
        RECT 37.900 10.800 38.300 13.100 ;
        RECT 39.000 10.800 39.400 13.100 ;
        RECT 40.600 10.800 41.000 13.100 ;
        RECT 42.200 10.800 42.600 13.100 ;
        RECT 43.800 10.800 44.200 13.100 ;
        RECT 45.400 10.800 45.800 13.100 ;
        RECT 47.000 10.800 47.400 13.100 ;
        RECT 48.600 10.800 49.000 13.100 ;
        RECT 49.400 10.800 49.800 13.100 ;
        RECT 51.000 10.800 51.400 13.100 ;
        RECT 52.600 10.800 53.000 13.100 ;
        RECT 55.000 10.800 55.400 13.100 ;
        RECT 56.600 10.800 57.000 13.100 ;
        RECT 59.000 10.800 59.400 12.700 ;
        RECT 63.000 10.800 63.400 13.100 ;
        RECT 64.600 10.800 65.000 13.100 ;
        RECT 67.300 10.800 67.800 12.100 ;
        RECT 69.000 10.800 69.400 12.100 ;
        RECT 71.800 10.800 72.200 13.000 ;
        RECT 74.200 10.800 74.600 13.300 ;
        RECT 76.800 10.800 77.200 13.500 ;
        RECT 79.000 10.800 79.400 13.100 ;
        RECT 81.700 10.800 82.200 12.100 ;
        RECT 83.400 10.800 83.800 12.100 ;
        RECT 86.200 10.800 86.600 13.000 ;
        RECT 87.800 10.800 88.200 12.100 ;
        RECT 90.000 10.800 90.400 13.500 ;
        RECT 92.600 10.800 93.000 13.300 ;
        RECT 95.000 10.800 95.400 13.000 ;
        RECT 97.800 10.800 98.200 12.100 ;
        RECT 99.400 10.800 99.900 12.100 ;
        RECT 102.200 10.800 102.600 13.100 ;
        RECT 103.800 10.800 104.200 13.100 ;
        RECT 105.400 10.800 105.800 13.100 ;
        RECT 108.900 10.800 109.300 13.100 ;
        RECT 111.000 10.800 111.400 12.100 ;
        RECT 111.800 10.800 112.200 12.100 ;
        RECT 113.400 10.800 113.800 12.100 ;
        RECT 114.800 10.800 115.200 13.500 ;
        RECT 117.400 10.800 117.800 13.300 ;
        RECT 119.600 10.800 120.000 13.500 ;
        RECT 122.200 10.800 122.600 13.300 ;
        RECT 124.600 10.800 125.000 13.000 ;
        RECT 127.400 10.800 127.800 12.100 ;
        RECT 129.000 10.800 129.500 12.100 ;
        RECT 131.800 10.800 132.200 13.100 ;
        RECT 133.400 10.800 133.800 13.100 ;
        RECT 135.000 10.800 135.400 13.100 ;
        RECT 136.600 10.800 137.000 13.100 ;
        RECT 138.200 10.800 138.600 13.100 ;
        RECT 139.800 10.800 140.200 13.100 ;
        RECT 140.600 10.800 141.000 13.100 ;
        RECT 142.200 10.800 142.600 13.100 ;
        RECT 143.800 10.800 144.200 13.100 ;
        RECT 145.400 10.800 145.800 13.100 ;
        RECT 147.000 10.800 147.400 13.100 ;
        RECT 148.600 10.800 149.000 13.100 ;
        RECT 151.300 10.800 151.800 12.100 ;
        RECT 153.000 10.800 153.400 12.100 ;
        RECT 155.800 10.800 156.200 13.000 ;
        RECT 159.800 10.800 160.200 13.300 ;
        RECT 162.400 10.800 162.800 13.500 ;
        RECT 164.600 10.800 165.000 12.100 ;
        RECT 166.200 10.800 166.600 13.300 ;
        RECT 168.800 10.800 169.200 13.500 ;
        RECT 170.200 10.800 170.600 13.100 ;
        RECT 171.800 10.800 172.200 13.100 ;
        RECT 173.400 10.800 173.800 13.100 ;
        RECT 175.000 10.800 175.400 12.700 ;
        RECT 179.000 10.800 179.400 13.100 ;
        RECT 180.400 10.800 180.800 13.500 ;
        RECT 183.000 10.800 183.400 13.300 ;
        RECT 185.400 10.800 185.800 13.100 ;
        RECT 188.100 10.800 188.600 12.100 ;
        RECT 189.800 10.800 190.200 12.100 ;
        RECT 192.600 10.800 193.000 13.000 ;
        RECT 195.000 10.800 195.400 13.100 ;
        RECT 196.600 10.800 197.000 13.100 ;
        RECT 197.400 10.800 197.800 13.100 ;
        RECT 199.000 10.800 199.400 13.100 ;
        RECT 200.600 10.800 201.000 13.100 ;
        RECT 202.200 10.800 202.600 13.100 ;
        RECT 203.800 10.800 204.200 13.100 ;
        RECT 205.400 10.800 205.800 12.700 ;
        RECT 211.000 10.800 211.400 12.700 ;
        RECT 213.400 10.800 213.800 13.000 ;
        RECT 216.200 10.800 216.600 12.100 ;
        RECT 217.800 10.800 218.300 12.100 ;
        RECT 220.600 10.800 221.000 13.100 ;
        RECT 223.000 10.800 223.400 13.100 ;
        RECT 224.600 10.800 225.000 13.100 ;
        RECT 225.400 10.800 225.800 13.100 ;
        RECT 228.600 10.800 229.000 13.300 ;
        RECT 231.200 10.800 231.600 13.500 ;
        RECT 233.400 10.800 233.800 13.000 ;
        RECT 236.200 10.800 236.600 12.100 ;
        RECT 237.800 10.800 238.300 12.100 ;
        RECT 240.600 10.800 241.000 13.100 ;
        RECT 242.200 10.800 242.600 13.100 ;
        RECT 243.800 10.800 244.200 13.100 ;
        RECT 245.400 10.800 245.800 13.100 ;
        RECT 247.000 10.800 247.400 13.100 ;
        RECT 248.600 10.800 249.000 13.100 ;
        RECT 250.200 10.800 250.600 12.700 ;
        RECT 252.600 10.800 253.000 13.100 ;
        RECT 255.800 10.800 256.200 13.000 ;
        RECT 258.600 10.800 259.000 12.100 ;
        RECT 260.200 10.800 260.700 12.100 ;
        RECT 263.000 10.800 263.400 13.100 ;
        RECT 0.200 10.200 265.400 10.800 ;
        RECT 0.600 7.900 1.000 10.200 ;
        RECT 2.200 7.900 2.600 10.200 ;
        RECT 3.800 7.900 4.200 10.200 ;
        RECT 5.400 7.900 5.800 10.200 ;
        RECT 7.000 7.900 7.400 10.200 ;
        RECT 7.800 7.900 8.200 10.200 ;
        RECT 11.000 7.900 11.400 10.200 ;
        RECT 13.700 8.900 14.200 10.200 ;
        RECT 15.400 8.900 15.800 10.200 ;
        RECT 18.200 8.000 18.600 10.200 ;
        RECT 20.600 8.000 21.000 10.200 ;
        RECT 23.400 8.900 23.800 10.200 ;
        RECT 25.000 8.900 25.500 10.200 ;
        RECT 27.800 7.900 28.200 10.200 ;
        RECT 29.400 7.900 29.800 10.200 ;
        RECT 33.400 8.300 33.800 10.200 ;
        RECT 35.000 7.900 35.400 10.200 ;
        RECT 36.600 7.900 37.000 10.200 ;
        RECT 38.200 7.900 38.600 10.200 ;
        RECT 39.800 7.900 40.200 10.200 ;
        RECT 41.400 7.900 41.800 10.200 ;
        RECT 42.200 7.900 42.600 10.200 ;
        RECT 43.800 7.900 44.200 10.200 ;
        RECT 45.400 7.900 45.800 10.200 ;
        RECT 47.000 7.900 47.400 10.200 ;
        RECT 48.600 7.900 49.000 10.200 ;
        RECT 49.400 7.900 49.800 10.200 ;
        RECT 51.000 7.900 51.400 10.200 ;
        RECT 52.600 7.900 53.000 10.200 ;
        RECT 54.200 7.900 54.600 10.200 ;
        RECT 55.800 7.900 56.200 10.200 ;
        RECT 58.200 7.900 58.600 10.200 ;
        RECT 59.800 7.900 60.200 10.200 ;
        RECT 61.400 7.900 61.800 10.200 ;
        RECT 63.000 7.900 63.400 10.200 ;
        RECT 64.600 7.900 65.000 10.200 ;
        RECT 66.200 7.700 66.600 10.200 ;
        RECT 68.800 7.500 69.200 10.200 ;
        RECT 71.000 8.900 71.400 10.200 ;
        RECT 72.600 7.900 73.000 10.200 ;
        RECT 75.300 8.900 75.800 10.200 ;
        RECT 77.000 8.900 77.400 10.200 ;
        RECT 79.800 8.000 80.200 10.200 ;
        RECT 82.200 8.000 82.600 10.200 ;
        RECT 85.000 8.900 85.400 10.200 ;
        RECT 86.600 8.900 87.100 10.200 ;
        RECT 89.400 7.900 89.800 10.200 ;
        RECT 91.000 7.900 91.400 10.200 ;
        RECT 95.000 8.300 95.400 10.200 ;
        RECT 97.400 7.900 97.800 10.200 ;
        RECT 100.100 8.900 100.600 10.200 ;
        RECT 101.800 8.900 102.200 10.200 ;
        RECT 104.600 8.000 105.000 10.200 ;
        RECT 107.800 8.900 108.200 10.200 ;
        RECT 110.000 7.500 110.400 10.200 ;
        RECT 112.600 7.700 113.000 10.200 ;
        RECT 115.000 8.300 115.400 10.200 ;
        RECT 119.000 7.900 119.400 10.200 ;
        RECT 120.600 8.000 121.000 10.200 ;
        RECT 123.400 8.900 123.800 10.200 ;
        RECT 125.000 8.900 125.500 10.200 ;
        RECT 127.800 7.900 128.200 10.200 ;
        RECT 129.400 7.900 129.800 10.200 ;
        RECT 133.400 8.300 133.800 10.200 ;
        RECT 135.800 8.000 136.200 10.200 ;
        RECT 138.600 8.900 139.000 10.200 ;
        RECT 140.200 8.900 140.700 10.200 ;
        RECT 143.000 7.900 143.400 10.200 ;
        RECT 144.600 7.900 145.000 10.200 ;
        RECT 146.200 7.900 146.600 10.200 ;
        RECT 147.800 7.900 148.200 10.200 ;
        RECT 149.400 7.900 149.800 10.200 ;
        RECT 151.000 7.900 151.400 10.200 ;
        RECT 151.800 7.900 152.200 10.200 ;
        RECT 153.400 7.900 153.800 10.200 ;
        RECT 157.400 7.900 157.800 10.200 ;
        RECT 160.100 8.900 160.600 10.200 ;
        RECT 161.800 8.900 162.200 10.200 ;
        RECT 164.600 8.000 165.000 10.200 ;
        RECT 166.200 8.900 166.600 10.200 ;
        RECT 168.400 7.500 168.800 10.200 ;
        RECT 171.000 7.700 171.400 10.200 ;
        RECT 172.600 7.900 173.000 10.200 ;
        RECT 174.200 7.900 174.600 10.200 ;
        RECT 175.800 7.900 176.200 10.200 ;
        RECT 177.400 7.700 177.800 10.200 ;
        RECT 180.000 7.500 180.400 10.200 ;
        RECT 182.200 8.900 182.600 10.200 ;
        RECT 183.800 8.000 184.200 10.200 ;
        RECT 186.600 8.900 187.000 10.200 ;
        RECT 188.200 8.900 188.700 10.200 ;
        RECT 191.000 7.900 191.400 10.200 ;
        RECT 193.400 7.900 193.800 10.200 ;
        RECT 196.100 8.900 196.600 10.200 ;
        RECT 197.800 8.900 198.200 10.200 ;
        RECT 200.600 8.000 201.000 10.200 ;
        RECT 203.000 7.900 203.400 10.200 ;
        RECT 205.700 8.900 206.200 10.200 ;
        RECT 207.400 8.900 207.800 10.200 ;
        RECT 210.200 8.000 210.600 10.200 ;
        RECT 214.200 8.300 214.600 10.200 ;
        RECT 218.200 7.900 218.600 10.200 ;
        RECT 219.000 7.900 219.400 10.200 ;
        RECT 220.600 7.900 221.000 10.200 ;
        RECT 222.200 7.900 222.600 10.200 ;
        RECT 223.800 7.900 224.200 10.200 ;
        RECT 225.400 7.900 225.800 10.200 ;
        RECT 227.800 8.300 228.200 10.200 ;
        RECT 230.200 8.000 230.600 10.200 ;
        RECT 233.000 8.900 233.400 10.200 ;
        RECT 234.600 8.900 235.100 10.200 ;
        RECT 237.400 7.900 237.800 10.200 ;
        RECT 239.000 7.900 239.400 10.200 ;
        RECT 240.600 7.900 241.000 10.200 ;
        RECT 242.200 7.900 242.600 10.200 ;
        RECT 243.800 7.900 244.200 10.200 ;
        RECT 245.400 7.900 245.800 10.200 ;
        RECT 246.200 7.900 246.600 10.200 ;
        RECT 247.800 7.900 248.200 10.200 ;
        RECT 249.400 7.900 249.800 10.200 ;
        RECT 251.000 7.900 251.400 10.200 ;
        RECT 252.600 7.900 253.000 10.200 ;
        RECT 254.200 8.000 254.600 10.200 ;
        RECT 257.000 8.900 257.400 10.200 ;
        RECT 258.600 8.900 259.100 10.200 ;
        RECT 261.400 7.900 261.800 10.200 ;
      LAYER via1 ;
        RECT 105.800 230.300 106.200 230.700 ;
        RECT 106.500 230.300 106.900 230.700 ;
        RECT 208.200 230.300 208.600 230.700 ;
        RECT 208.900 230.300 209.300 230.700 ;
        RECT 105.800 210.300 106.200 210.700 ;
        RECT 106.500 210.300 106.900 210.700 ;
        RECT 208.200 210.300 208.600 210.700 ;
        RECT 208.900 210.300 209.300 210.700 ;
        RECT 105.800 190.300 106.200 190.700 ;
        RECT 106.500 190.300 106.900 190.700 ;
        RECT 208.200 190.300 208.600 190.700 ;
        RECT 208.900 190.300 209.300 190.700 ;
        RECT 105.800 170.300 106.200 170.700 ;
        RECT 106.500 170.300 106.900 170.700 ;
        RECT 208.200 170.300 208.600 170.700 ;
        RECT 208.900 170.300 209.300 170.700 ;
        RECT 105.800 150.300 106.200 150.700 ;
        RECT 106.500 150.300 106.900 150.700 ;
        RECT 208.200 150.300 208.600 150.700 ;
        RECT 208.900 150.300 209.300 150.700 ;
        RECT 105.800 130.300 106.200 130.700 ;
        RECT 106.500 130.300 106.900 130.700 ;
        RECT 208.200 130.300 208.600 130.700 ;
        RECT 208.900 130.300 209.300 130.700 ;
        RECT 105.800 110.300 106.200 110.700 ;
        RECT 106.500 110.300 106.900 110.700 ;
        RECT 208.200 110.300 208.600 110.700 ;
        RECT 208.900 110.300 209.300 110.700 ;
        RECT 105.800 90.300 106.200 90.700 ;
        RECT 106.500 90.300 106.900 90.700 ;
        RECT 208.200 90.300 208.600 90.700 ;
        RECT 208.900 90.300 209.300 90.700 ;
        RECT 105.800 70.300 106.200 70.700 ;
        RECT 106.500 70.300 106.900 70.700 ;
        RECT 208.200 70.300 208.600 70.700 ;
        RECT 208.900 70.300 209.300 70.700 ;
        RECT 105.800 50.300 106.200 50.700 ;
        RECT 106.500 50.300 106.900 50.700 ;
        RECT 208.200 50.300 208.600 50.700 ;
        RECT 208.900 50.300 209.300 50.700 ;
        RECT 105.800 30.300 106.200 30.700 ;
        RECT 106.500 30.300 106.900 30.700 ;
        RECT 208.200 30.300 208.600 30.700 ;
        RECT 208.900 30.300 209.300 30.700 ;
        RECT 105.800 10.300 106.200 10.700 ;
        RECT 106.500 10.300 106.900 10.700 ;
        RECT 208.200 10.300 208.600 10.700 ;
        RECT 208.900 10.300 209.300 10.700 ;
      LAYER metal2 ;
        RECT 105.600 230.300 107.200 230.700 ;
        RECT 208.000 230.300 209.600 230.700 ;
        RECT 105.600 210.300 107.200 210.700 ;
        RECT 208.000 210.300 209.600 210.700 ;
        RECT 105.600 190.300 107.200 190.700 ;
        RECT 208.000 190.300 209.600 190.700 ;
        RECT 105.600 170.300 107.200 170.700 ;
        RECT 208.000 170.300 209.600 170.700 ;
        RECT 105.600 150.300 107.200 150.700 ;
        RECT 208.000 150.300 209.600 150.700 ;
        RECT 105.600 130.300 107.200 130.700 ;
        RECT 208.000 130.300 209.600 130.700 ;
        RECT 105.600 110.300 107.200 110.700 ;
        RECT 208.000 110.300 209.600 110.700 ;
        RECT 105.600 90.300 107.200 90.700 ;
        RECT 208.000 90.300 209.600 90.700 ;
        RECT 105.600 70.300 107.200 70.700 ;
        RECT 208.000 70.300 209.600 70.700 ;
        RECT 105.600 50.300 107.200 50.700 ;
        RECT 208.000 50.300 209.600 50.700 ;
        RECT 105.600 30.300 107.200 30.700 ;
        RECT 208.000 30.300 209.600 30.700 ;
        RECT 105.600 10.300 107.200 10.700 ;
        RECT 208.000 10.300 209.600 10.700 ;
      LAYER via2 ;
        RECT 105.800 230.300 106.200 230.700 ;
        RECT 106.500 230.300 106.900 230.700 ;
        RECT 208.200 230.300 208.600 230.700 ;
        RECT 208.900 230.300 209.300 230.700 ;
        RECT 105.800 210.300 106.200 210.700 ;
        RECT 106.500 210.300 106.900 210.700 ;
        RECT 208.200 210.300 208.600 210.700 ;
        RECT 208.900 210.300 209.300 210.700 ;
        RECT 105.800 190.300 106.200 190.700 ;
        RECT 106.500 190.300 106.900 190.700 ;
        RECT 208.200 190.300 208.600 190.700 ;
        RECT 208.900 190.300 209.300 190.700 ;
        RECT 105.800 170.300 106.200 170.700 ;
        RECT 106.500 170.300 106.900 170.700 ;
        RECT 208.200 170.300 208.600 170.700 ;
        RECT 208.900 170.300 209.300 170.700 ;
        RECT 105.800 150.300 106.200 150.700 ;
        RECT 106.500 150.300 106.900 150.700 ;
        RECT 208.200 150.300 208.600 150.700 ;
        RECT 208.900 150.300 209.300 150.700 ;
        RECT 105.800 130.300 106.200 130.700 ;
        RECT 106.500 130.300 106.900 130.700 ;
        RECT 208.200 130.300 208.600 130.700 ;
        RECT 208.900 130.300 209.300 130.700 ;
        RECT 105.800 110.300 106.200 110.700 ;
        RECT 106.500 110.300 106.900 110.700 ;
        RECT 208.200 110.300 208.600 110.700 ;
        RECT 208.900 110.300 209.300 110.700 ;
        RECT 105.800 90.300 106.200 90.700 ;
        RECT 106.500 90.300 106.900 90.700 ;
        RECT 208.200 90.300 208.600 90.700 ;
        RECT 208.900 90.300 209.300 90.700 ;
        RECT 105.800 70.300 106.200 70.700 ;
        RECT 106.500 70.300 106.900 70.700 ;
        RECT 208.200 70.300 208.600 70.700 ;
        RECT 208.900 70.300 209.300 70.700 ;
        RECT 105.800 50.300 106.200 50.700 ;
        RECT 106.500 50.300 106.900 50.700 ;
        RECT 208.200 50.300 208.600 50.700 ;
        RECT 208.900 50.300 209.300 50.700 ;
        RECT 105.800 30.300 106.200 30.700 ;
        RECT 106.500 30.300 106.900 30.700 ;
        RECT 208.200 30.300 208.600 30.700 ;
        RECT 208.900 30.300 209.300 30.700 ;
        RECT 105.800 10.300 106.200 10.700 ;
        RECT 106.500 10.300 106.900 10.700 ;
        RECT 208.200 10.300 208.600 10.700 ;
        RECT 208.900 10.300 209.300 10.700 ;
      LAYER metal3 ;
        RECT 105.600 230.300 107.200 230.700 ;
        RECT 208.000 230.300 209.600 230.700 ;
        RECT 105.600 210.300 107.200 210.700 ;
        RECT 208.000 210.300 209.600 210.700 ;
        RECT 105.600 190.300 107.200 190.700 ;
        RECT 208.000 190.300 209.600 190.700 ;
        RECT 105.600 170.300 107.200 170.700 ;
        RECT 208.000 170.300 209.600 170.700 ;
        RECT 105.600 150.300 107.200 150.700 ;
        RECT 208.000 150.300 209.600 150.700 ;
        RECT 105.600 130.300 107.200 130.700 ;
        RECT 208.000 130.300 209.600 130.700 ;
        RECT 105.600 110.300 107.200 110.700 ;
        RECT 208.000 110.300 209.600 110.700 ;
        RECT 105.600 90.300 107.200 90.700 ;
        RECT 208.000 90.300 209.600 90.700 ;
        RECT 105.600 70.300 107.200 70.700 ;
        RECT 208.000 70.300 209.600 70.700 ;
        RECT 105.600 50.300 107.200 50.700 ;
        RECT 208.000 50.300 209.600 50.700 ;
        RECT 105.600 30.300 107.200 30.700 ;
        RECT 208.000 30.300 209.600 30.700 ;
        RECT 105.600 10.300 107.200 10.700 ;
        RECT 208.000 10.300 209.600 10.700 ;
      LAYER via3 ;
        RECT 105.800 230.300 106.200 230.700 ;
        RECT 106.600 230.300 107.000 230.700 ;
        RECT 208.200 230.300 208.600 230.700 ;
        RECT 209.000 230.300 209.400 230.700 ;
        RECT 105.800 210.300 106.200 210.700 ;
        RECT 106.600 210.300 107.000 210.700 ;
        RECT 208.200 210.300 208.600 210.700 ;
        RECT 209.000 210.300 209.400 210.700 ;
        RECT 105.800 190.300 106.200 190.700 ;
        RECT 106.600 190.300 107.000 190.700 ;
        RECT 208.200 190.300 208.600 190.700 ;
        RECT 209.000 190.300 209.400 190.700 ;
        RECT 105.800 170.300 106.200 170.700 ;
        RECT 106.600 170.300 107.000 170.700 ;
        RECT 208.200 170.300 208.600 170.700 ;
        RECT 209.000 170.300 209.400 170.700 ;
        RECT 105.800 150.300 106.200 150.700 ;
        RECT 106.600 150.300 107.000 150.700 ;
        RECT 208.200 150.300 208.600 150.700 ;
        RECT 209.000 150.300 209.400 150.700 ;
        RECT 105.800 130.300 106.200 130.700 ;
        RECT 106.600 130.300 107.000 130.700 ;
        RECT 208.200 130.300 208.600 130.700 ;
        RECT 209.000 130.300 209.400 130.700 ;
        RECT 105.800 110.300 106.200 110.700 ;
        RECT 106.600 110.300 107.000 110.700 ;
        RECT 208.200 110.300 208.600 110.700 ;
        RECT 209.000 110.300 209.400 110.700 ;
        RECT 105.800 90.300 106.200 90.700 ;
        RECT 106.600 90.300 107.000 90.700 ;
        RECT 208.200 90.300 208.600 90.700 ;
        RECT 209.000 90.300 209.400 90.700 ;
        RECT 105.800 70.300 106.200 70.700 ;
        RECT 106.600 70.300 107.000 70.700 ;
        RECT 208.200 70.300 208.600 70.700 ;
        RECT 209.000 70.300 209.400 70.700 ;
        RECT 105.800 50.300 106.200 50.700 ;
        RECT 106.600 50.300 107.000 50.700 ;
        RECT 208.200 50.300 208.600 50.700 ;
        RECT 209.000 50.300 209.400 50.700 ;
        RECT 105.800 30.300 106.200 30.700 ;
        RECT 106.600 30.300 107.000 30.700 ;
        RECT 208.200 30.300 208.600 30.700 ;
        RECT 209.000 30.300 209.400 30.700 ;
        RECT 105.800 10.300 106.200 10.700 ;
        RECT 106.600 10.300 107.000 10.700 ;
        RECT 208.200 10.300 208.600 10.700 ;
        RECT 209.000 10.300 209.400 10.700 ;
      LAYER metal4 ;
        RECT 105.600 230.300 107.200 230.700 ;
        RECT 208.000 230.300 209.600 230.700 ;
        RECT 105.600 210.300 107.200 210.700 ;
        RECT 208.000 210.300 209.600 210.700 ;
        RECT 105.600 190.300 107.200 190.700 ;
        RECT 208.000 190.300 209.600 190.700 ;
        RECT 105.600 170.300 107.200 170.700 ;
        RECT 208.000 170.300 209.600 170.700 ;
        RECT 105.600 150.300 107.200 150.700 ;
        RECT 208.000 150.300 209.600 150.700 ;
        RECT 105.600 130.300 107.200 130.700 ;
        RECT 208.000 130.300 209.600 130.700 ;
        RECT 105.600 110.300 107.200 110.700 ;
        RECT 208.000 110.300 209.600 110.700 ;
        RECT 105.600 90.300 107.200 90.700 ;
        RECT 208.000 90.300 209.600 90.700 ;
        RECT 105.600 70.300 107.200 70.700 ;
        RECT 208.000 70.300 209.600 70.700 ;
        RECT 105.600 50.300 107.200 50.700 ;
        RECT 208.000 50.300 209.600 50.700 ;
        RECT 105.600 30.300 107.200 30.700 ;
        RECT 208.000 30.300 209.600 30.700 ;
        RECT 105.600 10.300 107.200 10.700 ;
        RECT 208.000 10.300 209.600 10.700 ;
      LAYER via4 ;
        RECT 105.800 230.300 106.200 230.700 ;
        RECT 106.500 230.300 106.900 230.700 ;
        RECT 208.200 230.300 208.600 230.700 ;
        RECT 208.900 230.300 209.300 230.700 ;
        RECT 105.800 210.300 106.200 210.700 ;
        RECT 106.500 210.300 106.900 210.700 ;
        RECT 208.200 210.300 208.600 210.700 ;
        RECT 208.900 210.300 209.300 210.700 ;
        RECT 105.800 190.300 106.200 190.700 ;
        RECT 106.500 190.300 106.900 190.700 ;
        RECT 208.200 190.300 208.600 190.700 ;
        RECT 208.900 190.300 209.300 190.700 ;
        RECT 105.800 170.300 106.200 170.700 ;
        RECT 106.500 170.300 106.900 170.700 ;
        RECT 208.200 170.300 208.600 170.700 ;
        RECT 208.900 170.300 209.300 170.700 ;
        RECT 105.800 150.300 106.200 150.700 ;
        RECT 106.500 150.300 106.900 150.700 ;
        RECT 208.200 150.300 208.600 150.700 ;
        RECT 208.900 150.300 209.300 150.700 ;
        RECT 105.800 130.300 106.200 130.700 ;
        RECT 106.500 130.300 106.900 130.700 ;
        RECT 208.200 130.300 208.600 130.700 ;
        RECT 208.900 130.300 209.300 130.700 ;
        RECT 105.800 110.300 106.200 110.700 ;
        RECT 106.500 110.300 106.900 110.700 ;
        RECT 208.200 110.300 208.600 110.700 ;
        RECT 208.900 110.300 209.300 110.700 ;
        RECT 105.800 90.300 106.200 90.700 ;
        RECT 106.500 90.300 106.900 90.700 ;
        RECT 208.200 90.300 208.600 90.700 ;
        RECT 208.900 90.300 209.300 90.700 ;
        RECT 105.800 70.300 106.200 70.700 ;
        RECT 106.500 70.300 106.900 70.700 ;
        RECT 208.200 70.300 208.600 70.700 ;
        RECT 208.900 70.300 209.300 70.700 ;
        RECT 105.800 50.300 106.200 50.700 ;
        RECT 106.500 50.300 106.900 50.700 ;
        RECT 208.200 50.300 208.600 50.700 ;
        RECT 208.900 50.300 209.300 50.700 ;
        RECT 105.800 30.300 106.200 30.700 ;
        RECT 106.500 30.300 106.900 30.700 ;
        RECT 208.200 30.300 208.600 30.700 ;
        RECT 208.900 30.300 209.300 30.700 ;
        RECT 105.800 10.300 106.200 10.700 ;
        RECT 106.500 10.300 106.900 10.700 ;
        RECT 208.200 10.300 208.600 10.700 ;
        RECT 208.900 10.300 209.300 10.700 ;
      LAYER metal5 ;
        RECT 105.600 230.200 107.200 230.700 ;
        RECT 208.000 230.200 209.600 230.700 ;
        RECT 105.600 210.200 107.200 210.700 ;
        RECT 208.000 210.200 209.600 210.700 ;
        RECT 105.600 190.200 107.200 190.700 ;
        RECT 208.000 190.200 209.600 190.700 ;
        RECT 105.600 170.200 107.200 170.700 ;
        RECT 208.000 170.200 209.600 170.700 ;
        RECT 105.600 150.200 107.200 150.700 ;
        RECT 208.000 150.200 209.600 150.700 ;
        RECT 105.600 130.200 107.200 130.700 ;
        RECT 208.000 130.200 209.600 130.700 ;
        RECT 105.600 110.200 107.200 110.700 ;
        RECT 208.000 110.200 209.600 110.700 ;
        RECT 105.600 90.200 107.200 90.700 ;
        RECT 208.000 90.200 209.600 90.700 ;
        RECT 105.600 70.200 107.200 70.700 ;
        RECT 208.000 70.200 209.600 70.700 ;
        RECT 105.600 50.200 107.200 50.700 ;
        RECT 208.000 50.200 209.600 50.700 ;
        RECT 105.600 30.200 107.200 30.700 ;
        RECT 208.000 30.200 209.600 30.700 ;
        RECT 105.600 10.200 107.200 10.700 ;
        RECT 208.000 10.200 209.600 10.700 ;
      LAYER via5 ;
        RECT 106.600 230.200 107.100 230.700 ;
        RECT 209.000 230.200 209.500 230.700 ;
        RECT 106.600 210.200 107.100 210.700 ;
        RECT 209.000 210.200 209.500 210.700 ;
        RECT 106.600 190.200 107.100 190.700 ;
        RECT 209.000 190.200 209.500 190.700 ;
        RECT 106.600 170.200 107.100 170.700 ;
        RECT 209.000 170.200 209.500 170.700 ;
        RECT 106.600 150.200 107.100 150.700 ;
        RECT 209.000 150.200 209.500 150.700 ;
        RECT 106.600 130.200 107.100 130.700 ;
        RECT 209.000 130.200 209.500 130.700 ;
        RECT 106.600 110.200 107.100 110.700 ;
        RECT 209.000 110.200 209.500 110.700 ;
        RECT 106.600 90.200 107.100 90.700 ;
        RECT 209.000 90.200 209.500 90.700 ;
        RECT 106.600 70.200 107.100 70.700 ;
        RECT 209.000 70.200 209.500 70.700 ;
        RECT 106.600 50.200 107.100 50.700 ;
        RECT 209.000 50.200 209.500 50.700 ;
        RECT 106.600 30.200 107.100 30.700 ;
        RECT 209.000 30.200 209.500 30.700 ;
        RECT 106.600 10.200 107.100 10.700 ;
        RECT 209.000 10.200 209.500 10.700 ;
      LAYER metal6 ;
        RECT 105.600 -3.000 107.200 243.000 ;
        RECT 208.000 -3.000 209.600 243.000 ;
    END
  END gnd
  PIN en
    PORT
      LAYER metal1 ;
        RECT 263.000 125.800 264.200 126.200 ;
      LAYER via1 ;
        RECT 263.800 125.800 264.200 126.200 ;
      LAYER metal2 ;
        RECT 263.800 131.800 264.200 132.200 ;
        RECT 263.800 126.200 264.100 131.800 ;
        RECT 263.800 125.800 264.200 126.200 ;
      LAYER metal3 ;
        RECT 263.800 132.100 264.200 132.200 ;
        RECT 267.800 132.100 268.200 132.200 ;
        RECT 263.800 131.800 268.200 132.100 ;
    END
  END en
  PIN rw
    PORT
      LAYER metal1 ;
        RECT 154.200 173.400 154.600 174.200 ;
        RECT 262.200 174.100 262.600 174.200 ;
        RECT 263.800 174.100 264.200 174.200 ;
        RECT 262.200 173.800 264.200 174.100 ;
        RECT 262.200 173.400 262.600 173.800 ;
        RECT 243.800 153.400 244.200 154.200 ;
        RECT 247.800 146.800 248.200 147.600 ;
        RECT 179.000 127.100 179.400 127.600 ;
        RECT 179.800 127.100 180.200 127.200 ;
        RECT 179.000 126.800 180.200 127.100 ;
        RECT 183.000 126.800 183.400 127.600 ;
        RECT 217.400 93.400 217.800 94.200 ;
        RECT 235.800 93.400 236.200 94.200 ;
        RECT 259.800 93.400 260.200 94.200 ;
      LAYER via1 ;
        RECT 154.200 173.800 154.600 174.200 ;
        RECT 263.800 173.800 264.200 174.200 ;
        RECT 243.800 153.800 244.200 154.200 ;
        RECT 179.800 126.800 180.200 127.200 ;
        RECT 217.400 93.800 217.800 94.200 ;
        RECT 235.800 93.800 236.200 94.200 ;
        RECT 259.800 93.800 260.200 94.200 ;
      LAYER metal2 ;
        RECT 154.200 173.800 154.600 174.200 ;
        RECT 263.800 173.800 264.200 174.200 ;
        RECT 154.200 167.200 154.500 173.800 ;
        RECT 154.200 166.800 154.600 167.200 ;
        RECT 243.800 153.800 244.200 154.200 ;
        RECT 243.800 148.200 244.100 153.800 ;
        RECT 263.800 148.200 264.100 173.800 ;
        RECT 243.800 147.800 244.200 148.200 ;
        RECT 247.800 147.800 248.200 148.200 ;
        RECT 263.800 147.800 264.200 148.200 ;
        RECT 247.800 147.200 248.100 147.800 ;
        RECT 247.800 146.800 248.200 147.200 ;
        RECT 179.800 126.800 180.200 127.200 ;
        RECT 183.000 126.800 183.400 127.200 ;
        RECT 179.800 126.200 180.100 126.800 ;
        RECT 179.800 125.800 180.200 126.200 ;
        RECT 183.000 114.200 183.300 126.800 ;
        RECT 183.000 113.800 183.400 114.200 ;
        RECT 259.800 104.800 260.200 105.200 ;
        RECT 259.800 94.200 260.100 104.800 ;
        RECT 217.400 94.100 217.800 94.200 ;
        RECT 218.200 94.100 218.600 94.200 ;
        RECT 217.400 93.800 218.600 94.100 ;
        RECT 235.800 94.100 236.200 94.200 ;
        RECT 236.600 94.100 237.000 94.200 ;
        RECT 235.800 93.800 237.000 94.100 ;
        RECT 259.800 93.800 260.200 94.200 ;
      LAYER via2 ;
        RECT 218.200 93.800 218.600 94.200 ;
        RECT 236.600 93.800 237.000 94.200 ;
      LAYER metal3 ;
        RECT 263.800 174.100 264.200 174.200 ;
        RECT 267.800 174.100 268.200 174.200 ;
        RECT 263.800 173.800 268.200 174.100 ;
        RECT 154.200 167.100 154.600 167.200 ;
        RECT 179.800 167.100 180.200 167.200 ;
        RECT 154.200 166.800 180.200 167.100 ;
        RECT 243.800 148.100 244.200 148.200 ;
        RECT 247.800 148.100 248.200 148.200 ;
        RECT 259.800 148.100 260.200 148.200 ;
        RECT 263.800 148.100 264.200 148.200 ;
        RECT 243.800 147.800 264.200 148.100 ;
        RECT 179.800 127.100 180.200 127.200 ;
        RECT 183.000 127.100 183.400 127.200 ;
        RECT 179.800 126.800 183.400 127.100 ;
        RECT 179.800 126.200 180.100 126.800 ;
        RECT 179.800 125.800 180.200 126.200 ;
        RECT 183.000 114.100 183.400 114.200 ;
        RECT 192.600 114.100 193.000 114.200 ;
        RECT 183.000 113.800 193.000 114.100 ;
        RECT 259.800 105.100 260.200 105.200 ;
        RECT 260.600 105.100 261.000 105.200 ;
        RECT 259.800 104.800 261.000 105.100 ;
        RECT 192.600 94.100 193.000 94.200 ;
        RECT 218.200 94.100 218.600 94.200 ;
        RECT 236.600 94.100 237.000 94.200 ;
        RECT 259.800 94.100 260.200 94.200 ;
        RECT 192.600 93.800 260.200 94.100 ;
      LAYER via3 ;
        RECT 179.800 166.800 180.200 167.200 ;
        RECT 259.800 147.800 260.200 148.200 ;
        RECT 192.600 113.800 193.000 114.200 ;
        RECT 260.600 104.800 261.000 105.200 ;
      LAYER metal4 ;
        RECT 179.800 166.800 180.200 167.200 ;
        RECT 179.800 127.200 180.100 166.800 ;
        RECT 259.800 147.800 260.200 148.200 ;
        RECT 179.800 126.800 180.200 127.200 ;
        RECT 192.600 113.800 193.000 114.200 ;
        RECT 192.600 94.200 192.900 113.800 ;
        RECT 259.800 105.100 260.100 147.800 ;
        RECT 260.600 105.100 261.000 105.200 ;
        RECT 259.800 104.800 261.000 105.100 ;
        RECT 192.600 93.800 193.000 94.200 ;
    END
  END rw
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 0.600 234.100 1.500 234.500 ;
        RECT 7.800 234.100 8.700 234.500 ;
        RECT 22.200 234.100 23.100 234.500 ;
        RECT 232.900 234.100 233.800 234.500 ;
        RECT 0.600 233.800 1.000 234.100 ;
        RECT 7.800 233.800 8.200 234.100 ;
        RECT 22.200 233.800 22.600 234.100 ;
        RECT 233.400 233.800 233.800 234.100 ;
        RECT 255.800 234.100 256.700 234.500 ;
        RECT 255.800 233.800 256.200 234.100 ;
        RECT 166.500 214.100 167.400 214.500 ;
        RECT 167.000 213.800 167.400 214.100 ;
        RECT 0.600 114.100 1.500 114.500 ;
        RECT 0.600 113.800 1.000 114.100 ;
        RECT 84.600 86.900 85.000 87.200 ;
        RECT 247.800 86.900 248.200 87.200 ;
        RECT 84.600 86.500 85.500 86.900 ;
        RECT 247.800 86.500 248.700 86.900 ;
        RECT 205.700 74.100 206.600 74.500 ;
        RECT 206.200 73.800 206.600 74.100 ;
        RECT 7.000 66.900 7.400 67.200 ;
        RECT 147.800 66.900 148.200 67.200 ;
        RECT 6.500 66.500 7.400 66.900 ;
        RECT 147.300 66.500 148.200 66.900 ;
        RECT 146.500 14.100 147.400 14.500 ;
        RECT 147.000 13.800 147.400 14.100 ;
        RECT 0.600 6.900 1.000 7.200 ;
        RECT 42.200 6.900 42.600 7.200 ;
        RECT 239.000 6.900 239.400 7.200 ;
        RECT 0.600 6.500 1.500 6.900 ;
        RECT 42.200 6.500 43.100 6.900 ;
        RECT 239.000 6.500 239.900 6.900 ;
      LAYER via1 ;
        RECT 84.600 86.800 85.000 87.200 ;
        RECT 247.800 86.800 248.200 87.200 ;
        RECT 7.000 66.800 7.400 67.200 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 42.200 6.800 42.600 7.200 ;
        RECT 239.000 6.800 239.400 7.200 ;
      LAYER metal2 ;
        RECT 0.600 234.100 1.000 234.200 ;
        RECT 1.400 234.100 1.800 234.200 ;
        RECT 0.600 233.800 1.800 234.100 ;
        RECT 7.000 234.100 7.400 234.200 ;
        RECT 7.800 234.100 8.200 234.200 ;
        RECT 7.000 233.800 8.200 234.100 ;
        RECT 22.200 234.100 22.600 234.200 ;
        RECT 23.000 234.100 23.400 234.200 ;
        RECT 22.200 233.800 23.400 234.100 ;
        RECT 233.400 233.800 233.800 234.200 ;
        RECT 255.800 233.800 256.200 234.200 ;
        RECT 233.400 232.200 233.700 233.800 ;
        RECT 255.800 232.200 256.100 233.800 ;
        RECT 233.400 231.800 233.800 232.200 ;
        RECT 255.800 231.800 256.200 232.200 ;
        RECT 167.000 214.100 167.400 214.200 ;
        RECT 167.800 214.100 168.200 214.200 ;
        RECT 167.000 213.800 168.200 214.100 ;
        RECT 0.600 114.100 1.000 114.200 ;
        RECT 1.400 114.100 1.800 114.200 ;
        RECT 0.600 113.800 1.800 114.100 ;
        RECT 84.600 86.800 85.000 87.200 ;
        RECT 247.800 86.800 248.200 87.200 ;
        RECT 84.600 83.200 84.900 86.800 ;
        RECT 84.600 82.800 85.000 83.200 ;
        RECT 7.800 81.800 8.200 82.200 ;
        RECT 7.800 68.100 8.100 81.800 ;
        RECT 247.800 74.200 248.100 86.800 ;
        RECT 206.200 74.100 206.600 74.200 ;
        RECT 207.000 74.100 207.400 74.200 ;
        RECT 206.200 73.800 207.400 74.100 ;
        RECT 247.800 73.800 248.200 74.200 ;
        RECT 7.000 67.800 8.100 68.100 ;
        RECT 147.800 67.800 148.200 68.200 ;
        RECT 7.000 67.200 7.300 67.800 ;
        RECT 147.800 67.200 148.100 67.800 ;
        RECT 7.000 66.800 7.400 67.200 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 147.000 17.800 147.400 18.200 ;
        RECT 147.000 14.200 147.300 17.800 ;
        RECT 147.000 13.800 147.400 14.200 ;
        RECT 0.600 7.800 1.000 8.200 ;
        RECT 42.200 7.800 42.600 8.200 ;
        RECT 239.000 7.800 239.400 8.200 ;
        RECT 0.600 7.200 0.900 7.800 ;
        RECT 42.200 7.200 42.500 7.800 ;
        RECT 239.000 7.200 239.300 7.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 42.200 6.800 42.600 7.200 ;
        RECT 239.000 6.800 239.400 7.200 ;
      LAYER via2 ;
        RECT 1.400 233.800 1.800 234.200 ;
        RECT 23.000 233.800 23.400 234.200 ;
        RECT 167.800 213.800 168.200 214.200 ;
        RECT 1.400 113.800 1.800 114.200 ;
        RECT 207.000 73.800 207.400 74.200 ;
      LAYER metal3 ;
        RECT -2.600 234.100 -2.200 234.200 ;
        RECT 0.600 234.100 1.000 234.200 ;
        RECT 1.400 234.100 1.800 234.200 ;
        RECT 7.000 234.100 7.400 234.200 ;
        RECT 23.000 234.100 23.400 234.200 ;
        RECT -2.600 233.800 23.400 234.100 ;
        RECT 171.000 232.100 171.400 232.200 ;
        RECT 233.400 232.100 233.800 232.200 ;
        RECT 255.800 232.100 256.200 232.200 ;
        RECT 171.000 231.800 256.200 232.100 ;
        RECT 167.800 214.100 168.200 214.200 ;
        RECT 171.000 214.100 171.400 214.200 ;
        RECT 167.800 213.800 171.400 214.100 ;
        RECT 0.600 114.100 1.000 114.200 ;
        RECT 1.400 114.100 1.800 114.200 ;
        RECT 0.600 113.800 1.800 114.100 ;
        RECT 84.600 83.100 85.000 83.200 ;
        RECT 147.800 83.100 148.200 83.200 ;
        RECT 84.600 82.800 148.200 83.100 ;
        RECT 0.600 82.100 1.000 82.200 ;
        RECT 7.800 82.100 8.200 82.200 ;
        RECT 84.600 82.100 84.900 82.800 ;
        RECT 0.600 81.800 84.900 82.100 ;
        RECT 201.400 74.100 201.800 74.200 ;
        RECT 207.000 74.100 207.400 74.200 ;
        RECT 239.000 74.100 239.400 74.200 ;
        RECT 247.800 74.100 248.200 74.200 ;
        RECT 201.400 73.800 248.200 74.100 ;
        RECT 147.800 67.800 148.200 68.200 ;
        RECT 147.800 67.200 148.100 67.800 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 147.000 18.100 147.400 18.200 ;
        RECT 147.800 18.100 148.200 18.200 ;
        RECT 147.000 17.800 148.200 18.100 ;
        RECT 0.600 8.100 1.000 8.200 ;
        RECT 42.200 8.100 42.600 8.200 ;
        RECT 0.600 7.800 42.600 8.100 ;
        RECT 239.000 7.800 239.400 8.200 ;
        RECT 0.600 7.200 0.900 7.800 ;
        RECT 239.000 7.200 239.300 7.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 239.000 6.800 239.400 7.200 ;
      LAYER via3 ;
        RECT 0.600 233.800 1.000 234.200 ;
        RECT 171.000 213.800 171.400 214.200 ;
        RECT 147.800 82.800 148.200 83.200 ;
        RECT 239.000 73.800 239.400 74.200 ;
        RECT 147.800 17.800 148.200 18.200 ;
      LAYER metal4 ;
        RECT 0.600 233.800 1.000 234.200 ;
        RECT 0.600 114.200 0.900 233.800 ;
        RECT 171.000 231.800 171.400 232.200 ;
        RECT 171.000 214.200 171.300 231.800 ;
        RECT 171.000 213.800 171.400 214.200 ;
        RECT 0.600 113.800 1.000 114.200 ;
        RECT 0.600 82.200 0.900 113.800 ;
        RECT 147.800 82.800 148.200 83.200 ;
        RECT 0.600 81.800 1.000 82.200 ;
        RECT 0.600 7.200 0.900 81.800 ;
        RECT 147.800 69.200 148.100 82.800 ;
        RECT 171.000 69.200 171.300 213.800 ;
        RECT 201.400 73.800 201.800 74.200 ;
        RECT 239.000 73.800 239.400 74.200 ;
        RECT 201.400 69.200 201.700 73.800 ;
        RECT 147.800 68.800 148.200 69.200 ;
        RECT 171.000 68.800 171.400 69.200 ;
        RECT 201.400 68.800 201.800 69.200 ;
        RECT 147.800 67.200 148.100 68.800 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 147.800 18.200 148.100 66.800 ;
        RECT 147.800 17.800 148.200 18.200 ;
        RECT 239.000 7.200 239.300 73.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 239.000 6.800 239.400 7.200 ;
      LAYER metal5 ;
        RECT 147.800 69.100 148.200 69.200 ;
        RECT 171.000 69.100 171.400 69.200 ;
        RECT 201.400 69.100 201.800 69.200 ;
        RECT 147.800 68.800 201.800 69.100 ;
    END
  END clk
  PIN ras
    PORT
      LAYER metal1 ;
        RECT 262.200 124.800 262.600 125.600 ;
        RECT 234.600 115.200 235.000 115.400 ;
        RECT 234.200 114.900 235.000 115.200 ;
        RECT 234.200 114.800 234.600 114.900 ;
        RECT 240.600 112.400 241.000 113.200 ;
        RECT 262.200 107.800 262.600 108.600 ;
        RECT 242.200 106.100 242.600 106.200 ;
        RECT 242.200 105.800 243.000 106.100 ;
        RECT 242.600 105.600 243.000 105.800 ;
        RECT 252.200 95.200 252.600 95.400 ;
        RECT 251.800 94.900 252.600 95.200 ;
        RECT 251.800 94.800 252.200 94.900 ;
        RECT 257.400 92.400 257.800 93.200 ;
      LAYER via1 ;
        RECT 240.600 112.800 241.000 113.200 ;
        RECT 257.400 92.800 257.800 93.200 ;
      LAYER metal2 ;
        RECT 262.200 125.100 262.600 125.200 ;
        RECT 261.400 124.800 262.600 125.100 ;
        RECT 261.400 117.200 261.700 124.800 ;
        RECT 261.400 116.800 261.800 117.200 ;
        RECT 234.200 115.100 234.600 115.200 ;
        RECT 235.000 115.100 235.400 115.200 ;
        RECT 234.200 114.800 235.400 115.100 ;
        RECT 240.600 114.800 241.000 115.200 ;
        RECT 240.600 113.200 240.900 114.800 ;
        RECT 240.600 112.800 241.000 113.200 ;
        RECT 240.600 108.200 240.900 112.800 ;
        RECT 261.400 108.200 261.700 116.800 ;
        RECT 240.600 107.800 241.000 108.200 ;
        RECT 242.200 107.800 242.600 108.200 ;
        RECT 257.400 107.800 257.800 108.200 ;
        RECT 261.400 108.100 261.800 108.200 ;
        RECT 262.200 108.100 262.600 108.200 ;
        RECT 261.400 107.800 262.600 108.100 ;
        RECT 242.200 106.200 242.500 107.800 ;
        RECT 242.200 105.800 242.600 106.200 ;
        RECT 257.400 95.200 257.700 107.800 ;
        RECT 251.800 95.100 252.200 95.200 ;
        RECT 252.600 95.100 253.000 95.200 ;
        RECT 251.800 94.800 253.000 95.100 ;
        RECT 257.400 94.800 257.800 95.200 ;
        RECT 257.400 93.200 257.700 94.800 ;
        RECT 257.400 92.800 257.800 93.200 ;
      LAYER via2 ;
        RECT 235.000 114.800 235.400 115.200 ;
        RECT 252.600 94.800 253.000 95.200 ;
      LAYER metal3 ;
        RECT 261.400 117.100 261.800 117.200 ;
        RECT 267.800 117.100 268.200 117.200 ;
        RECT 261.400 116.800 268.200 117.100 ;
        RECT 235.000 115.100 235.400 115.200 ;
        RECT 240.600 115.100 241.000 115.200 ;
        RECT 235.000 114.800 241.000 115.100 ;
        RECT 240.600 108.100 241.000 108.200 ;
        RECT 242.200 108.100 242.600 108.200 ;
        RECT 257.400 108.100 257.800 108.200 ;
        RECT 261.400 108.100 261.800 108.200 ;
        RECT 240.600 107.800 261.800 108.100 ;
        RECT 252.600 95.100 253.000 95.200 ;
        RECT 257.400 95.100 257.800 95.200 ;
        RECT 252.600 94.800 257.800 95.100 ;
    END
  END ras
  PIN cas
    PORT
      LAYER metal1 ;
        RECT 241.000 135.200 241.400 135.400 ;
        RECT 253.800 135.200 254.200 135.400 ;
        RECT 240.600 134.900 241.400 135.200 ;
        RECT 253.400 134.900 254.200 135.200 ;
        RECT 240.600 134.800 241.000 134.900 ;
        RECT 253.400 134.800 253.800 134.900 ;
        RECT 258.200 133.800 258.600 134.200 ;
        RECT 256.600 132.400 257.000 133.200 ;
        RECT 258.200 133.100 258.500 133.800 ;
        RECT 259.000 133.100 259.400 133.200 ;
        RECT 258.200 132.800 259.400 133.100 ;
        RECT 259.000 132.400 259.400 132.800 ;
        RECT 263.800 123.800 264.200 124.600 ;
      LAYER via1 ;
        RECT 256.600 132.800 257.000 133.200 ;
      LAYER metal2 ;
        RECT 240.600 134.800 241.000 135.200 ;
        RECT 253.400 134.800 253.800 135.200 ;
        RECT 240.600 133.200 240.900 134.800 ;
        RECT 253.400 133.200 253.700 134.800 ;
        RECT 258.200 133.800 258.600 134.200 ;
        RECT 258.200 133.200 258.500 133.800 ;
        RECT 240.600 132.800 241.000 133.200 ;
        RECT 253.400 132.800 253.800 133.200 ;
        RECT 256.600 133.100 257.000 133.200 ;
        RECT 257.400 133.100 257.800 133.200 ;
        RECT 256.600 132.800 257.800 133.100 ;
        RECT 258.200 132.800 258.600 133.200 ;
        RECT 258.200 128.200 258.500 132.800 ;
        RECT 258.200 127.800 258.600 128.200 ;
        RECT 264.600 127.800 265.000 128.200 ;
        RECT 263.800 124.100 264.200 124.200 ;
        RECT 264.600 124.100 264.900 127.800 ;
        RECT 263.800 123.800 264.900 124.100 ;
      LAYER via2 ;
        RECT 257.400 132.800 257.800 133.200 ;
      LAYER metal3 ;
        RECT 240.600 133.100 241.000 133.200 ;
        RECT 253.400 133.100 253.800 133.200 ;
        RECT 257.400 133.100 257.800 133.200 ;
        RECT 258.200 133.100 258.600 133.200 ;
        RECT 240.600 132.800 258.600 133.100 ;
        RECT 258.200 128.100 258.600 128.200 ;
        RECT 264.600 128.100 265.000 128.200 ;
        RECT 267.800 128.100 268.200 128.200 ;
        RECT 258.200 127.800 268.200 128.100 ;
    END
  END cas
  PIN datain[0]
    PORT
      LAYER metal1 ;
        RECT 230.200 226.800 230.600 227.600 ;
      LAYER metal2 ;
        RECT 228.600 242.800 229.000 243.200 ;
        RECT 228.600 240.200 228.900 242.800 ;
        RECT 228.600 239.800 229.000 240.200 ;
        RECT 230.200 239.800 230.600 240.200 ;
        RECT 230.200 227.200 230.500 239.800 ;
        RECT 230.200 226.800 230.600 227.200 ;
      LAYER metal3 ;
        RECT 228.600 240.100 229.000 240.200 ;
        RECT 230.200 240.100 230.600 240.200 ;
        RECT 228.600 239.800 230.600 240.100 ;
    END
  END datain[0]
  PIN datain[1]
    PORT
      LAYER metal1 ;
        RECT 52.600 13.400 53.000 14.200 ;
      LAYER via1 ;
        RECT 52.600 13.800 53.000 14.200 ;
      LAYER metal2 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 52.600 1.200 52.900 13.800 ;
        RECT 51.000 0.800 51.400 1.200 ;
        RECT 52.600 0.800 53.000 1.200 ;
        RECT 51.000 -1.800 51.300 0.800 ;
        RECT 51.000 -2.200 51.400 -1.800 ;
      LAYER metal3 ;
        RECT 51.000 1.100 51.400 1.200 ;
        RECT 52.600 1.100 53.000 1.200 ;
        RECT 51.000 0.800 53.000 1.100 ;
    END
  END datain[1]
  PIN datain[2]
    PORT
      LAYER metal1 ;
        RECT 263.000 147.100 263.400 147.600 ;
        RECT 264.600 147.100 265.000 147.200 ;
        RECT 263.000 146.800 265.000 147.100 ;
      LAYER via1 ;
        RECT 264.600 146.800 265.000 147.200 ;
      LAYER metal2 ;
        RECT 264.600 146.800 265.000 147.200 ;
        RECT 264.600 145.200 264.900 146.800 ;
        RECT 264.600 144.800 265.000 145.200 ;
      LAYER metal3 ;
        RECT 264.600 145.100 265.000 145.200 ;
        RECT 267.800 145.100 268.200 145.200 ;
        RECT 264.600 144.800 268.200 145.100 ;
    END
  END datain[2]
  PIN datain[3]
    PORT
      LAYER metal1 ;
        RECT 0.600 106.800 1.000 107.600 ;
      LAYER metal2 ;
        RECT 0.600 106.800 1.000 107.200 ;
        RECT 0.600 105.200 0.900 106.800 ;
        RECT 0.600 104.800 1.000 105.200 ;
      LAYER metal3 ;
        RECT -2.600 105.100 -2.200 105.200 ;
        RECT 0.600 105.100 1.000 105.200 ;
        RECT -2.600 104.800 1.000 105.100 ;
    END
  END datain[3]
  PIN datain[4]
    PORT
      LAYER metal1 ;
        RECT 170.200 13.400 170.600 14.200 ;
      LAYER via1 ;
        RECT 170.200 13.800 170.600 14.200 ;
      LAYER metal2 ;
        RECT 170.200 13.800 170.600 14.200 ;
        RECT 170.200 -1.900 170.500 13.800 ;
        RECT 171.800 -1.900 172.200 -1.800 ;
        RECT 170.200 -2.200 172.200 -1.900 ;
    END
  END datain[4]
  PIN datain[5]
    PORT
      LAYER metal1 ;
        RECT 48.600 226.800 49.000 227.600 ;
      LAYER metal2 ;
        RECT 50.200 242.800 50.600 243.200 ;
        RECT 50.200 240.200 50.500 242.800 ;
        RECT 48.600 239.800 49.000 240.200 ;
        RECT 50.200 239.800 50.600 240.200 ;
        RECT 48.600 227.200 48.900 239.800 ;
        RECT 48.600 226.800 49.000 227.200 ;
      LAYER metal3 ;
        RECT 48.600 240.100 49.000 240.200 ;
        RECT 50.200 240.100 50.600 240.200 ;
        RECT 48.600 239.800 50.600 240.100 ;
    END
  END datain[5]
  PIN datain[6]
    PORT
      LAYER metal1 ;
        RECT 175.800 6.800 176.200 7.600 ;
      LAYER metal2 ;
        RECT 174.200 6.800 174.600 7.200 ;
        RECT 175.800 7.100 176.200 7.200 ;
        RECT 176.600 7.100 177.000 7.200 ;
        RECT 175.800 6.800 177.000 7.100 ;
        RECT 174.200 -1.800 174.500 6.800 ;
        RECT 174.200 -2.200 174.600 -1.800 ;
      LAYER via2 ;
        RECT 176.600 6.800 177.000 7.200 ;
      LAYER metal3 ;
        RECT 174.200 7.100 174.600 7.200 ;
        RECT 176.600 7.100 177.000 7.200 ;
        RECT 174.200 6.800 177.000 7.100 ;
    END
  END datain[6]
  PIN datain[7]
    PORT
      LAYER metal1 ;
        RECT 117.400 227.100 117.800 227.200 ;
        RECT 118.200 227.100 118.600 227.600 ;
        RECT 117.400 226.800 118.600 227.100 ;
      LAYER metal2 ;
        RECT 119.800 242.800 120.200 243.200 ;
        RECT 119.800 240.200 120.100 242.800 ;
        RECT 117.400 239.800 117.800 240.200 ;
        RECT 119.800 239.800 120.200 240.200 ;
        RECT 117.400 227.200 117.700 239.800 ;
        RECT 117.400 226.800 117.800 227.200 ;
      LAYER metal3 ;
        RECT 117.400 240.100 117.800 240.200 ;
        RECT 119.800 240.100 120.200 240.200 ;
        RECT 117.400 239.800 120.200 240.100 ;
    END
  END datain[7]
  PIN address[0]
    PORT
      LAYER metal1 ;
        RECT 260.600 134.800 261.000 135.600 ;
        RECT 260.600 134.200 260.900 134.800 ;
        RECT 260.600 133.800 261.000 134.200 ;
      LAYER metal2 ;
        RECT 260.600 134.800 261.000 135.200 ;
        RECT 260.600 134.200 260.900 134.800 ;
        RECT 260.600 133.800 261.000 134.200 ;
      LAYER metal3 ;
        RECT 260.600 135.100 261.000 135.200 ;
        RECT 267.800 135.100 268.200 135.200 ;
        RECT 260.600 134.800 268.200 135.100 ;
    END
  END address[0]
  PIN address[1]
    PORT
      LAYER metal1 ;
        RECT 258.200 135.100 258.600 135.600 ;
        RECT 259.000 135.100 259.400 135.200 ;
        RECT 258.200 134.800 259.400 135.100 ;
      LAYER via1 ;
        RECT 259.000 134.800 259.400 135.200 ;
      LAYER metal2 ;
        RECT 259.000 136.800 259.400 137.200 ;
        RECT 259.000 135.200 259.300 136.800 ;
        RECT 259.000 134.800 259.400 135.200 ;
      LAYER metal3 ;
        RECT 259.000 137.100 259.400 137.200 ;
        RECT 267.800 137.100 268.200 137.200 ;
        RECT 259.000 136.800 268.200 137.100 ;
    END
  END address[1]
  PIN address[2]
    PORT
      LAYER metal1 ;
        RECT 242.200 114.800 242.600 115.600 ;
        RECT 242.200 114.200 242.500 114.800 ;
        RECT 242.200 113.800 242.600 114.200 ;
      LAYER metal2 ;
        RECT 242.200 114.800 242.600 115.200 ;
        RECT 242.200 114.200 242.500 114.800 ;
        RECT 242.200 113.800 242.600 114.200 ;
      LAYER metal3 ;
        RECT 257.400 115.800 268.100 116.100 ;
        RECT 242.200 115.100 242.600 115.200 ;
        RECT 257.400 115.100 257.700 115.800 ;
        RECT 242.200 114.800 257.700 115.100 ;
        RECT 267.800 115.200 268.100 115.800 ;
        RECT 267.800 114.800 268.200 115.200 ;
    END
  END address[2]
  PIN address[3]
    PORT
      LAYER metal1 ;
        RECT 259.000 94.800 259.400 95.600 ;
        RECT 259.000 94.200 259.300 94.800 ;
        RECT 259.000 93.800 259.400 94.200 ;
      LAYER metal2 ;
        RECT 259.000 94.800 259.400 95.200 ;
        RECT 259.000 94.200 259.300 94.800 ;
        RECT 259.000 93.800 259.400 94.200 ;
      LAYER metal3 ;
        RECT 259.000 95.100 259.400 95.200 ;
        RECT 267.800 95.100 268.200 95.200 ;
        RECT 259.000 94.800 268.200 95.100 ;
    END
  END address[3]
  PIN address[4]
    PORT
      LAYER metal1 ;
        RECT 263.800 106.100 264.200 106.200 ;
        RECT 264.600 106.100 265.000 106.200 ;
        RECT 263.800 105.800 265.000 106.100 ;
        RECT 263.800 105.400 264.200 105.800 ;
      LAYER via1 ;
        RECT 264.600 105.800 265.000 106.200 ;
      LAYER metal2 ;
        RECT 264.600 105.800 265.000 106.200 ;
        RECT 264.600 105.200 264.900 105.800 ;
        RECT 264.600 104.800 265.000 105.200 ;
      LAYER metal3 ;
        RECT 264.600 105.100 265.000 105.200 ;
        RECT 267.800 105.100 268.200 105.200 ;
        RECT 264.600 104.800 268.200 105.100 ;
    END
  END address[4]
  PIN dataout[0]
    PORT
      LAYER metal1 ;
        RECT 263.800 166.200 264.200 169.900 ;
        RECT 263.900 165.100 264.200 166.200 ;
        RECT 263.800 164.100 264.200 165.100 ;
        RECT 264.600 164.100 265.000 164.200 ;
        RECT 263.800 163.800 265.000 164.100 ;
        RECT 263.800 161.100 264.200 163.800 ;
      LAYER via1 ;
        RECT 264.600 163.800 265.000 164.200 ;
      LAYER metal2 ;
        RECT 264.600 164.800 265.000 165.200 ;
        RECT 264.600 164.200 264.900 164.800 ;
        RECT 264.600 163.800 265.000 164.200 ;
      LAYER metal3 ;
        RECT 264.600 165.100 265.000 165.200 ;
        RECT 267.800 165.100 268.200 165.200 ;
        RECT 264.600 164.800 268.200 165.100 ;
    END
  END dataout[0]
  PIN dataout[1]
    PORT
      LAYER metal1 ;
        RECT 263.800 97.100 264.200 99.900 ;
        RECT 264.600 97.800 265.000 98.200 ;
        RECT 264.600 97.100 264.900 97.800 ;
        RECT 263.800 96.800 264.900 97.100 ;
        RECT 263.800 95.900 264.200 96.800 ;
        RECT 263.900 94.800 264.200 95.900 ;
        RECT 263.800 91.100 264.200 94.800 ;
      LAYER metal2 ;
        RECT 264.600 97.800 265.000 98.200 ;
        RECT 264.600 97.200 264.900 97.800 ;
        RECT 264.600 96.800 265.000 97.200 ;
      LAYER metal3 ;
        RECT 264.600 97.100 265.000 97.200 ;
        RECT 267.800 97.100 268.200 97.200 ;
        RECT 264.600 96.800 268.200 97.100 ;
    END
  END dataout[1]
  PIN dataout[2]
    PORT
      LAYER metal1 ;
        RECT 261.400 126.200 261.800 129.900 ;
        RECT 261.500 125.100 261.800 126.200 ;
        RECT 261.400 124.100 261.800 125.100 ;
        RECT 263.000 124.100 263.400 124.200 ;
        RECT 261.400 123.800 263.400 124.100 ;
        RECT 261.400 121.100 261.800 123.800 ;
      LAYER via1 ;
        RECT 263.000 123.800 263.400 124.200 ;
      LAYER metal2 ;
        RECT 263.000 124.800 263.400 125.200 ;
        RECT 263.000 124.200 263.300 124.800 ;
        RECT 263.000 123.800 263.400 124.200 ;
      LAYER metal3 ;
        RECT 263.000 125.100 263.400 125.200 ;
        RECT 267.800 125.100 268.200 125.200 ;
        RECT 263.000 124.800 268.200 125.100 ;
    END
  END dataout[2]
  PIN dataout[3]
    PORT
      LAYER metal1 ;
        RECT 203.800 126.200 204.200 129.900 ;
        RECT 203.900 125.100 204.200 126.200 ;
        RECT 203.800 121.100 204.200 125.100 ;
      LAYER via1 ;
        RECT 203.800 128.800 204.200 129.200 ;
      LAYER metal2 ;
        RECT 203.800 129.100 204.200 129.200 ;
        RECT 204.600 129.100 205.000 129.200 ;
        RECT 203.800 128.800 205.000 129.100 ;
      LAYER via2 ;
        RECT 204.600 128.800 205.000 129.200 ;
      LAYER metal3 ;
        RECT 264.600 130.100 265.000 130.200 ;
        RECT 267.800 130.100 268.200 130.200 ;
        RECT 264.600 129.800 268.200 130.100 ;
        RECT 204.600 129.100 205.000 129.200 ;
        RECT 207.800 129.100 208.200 129.200 ;
        RECT 203.800 128.800 208.200 129.100 ;
      LAYER via3 ;
        RECT 207.800 128.800 208.200 129.200 ;
      LAYER metal4 ;
        RECT 264.600 129.800 265.000 130.200 ;
        RECT 264.600 129.200 264.900 129.800 ;
        RECT 207.800 129.100 208.200 129.200 ;
        RECT 208.600 129.100 209.000 129.200 ;
        RECT 207.800 128.800 209.000 129.100 ;
        RECT 264.600 128.800 265.000 129.200 ;
      LAYER via4 ;
        RECT 208.600 128.800 209.000 129.200 ;
      LAYER metal5 ;
        RECT 208.600 129.100 209.000 129.200 ;
        RECT 264.600 129.100 265.000 129.200 ;
        RECT 208.600 128.800 265.000 129.100 ;
    END
  END dataout[3]
  PIN dataout[4]
    PORT
      LAYER metal1 ;
        RECT 256.600 95.900 257.000 99.900 ;
        RECT 256.700 94.800 257.000 95.900 ;
        RECT 256.600 91.100 257.000 94.800 ;
      LAYER via1 ;
        RECT 256.600 98.800 257.000 99.200 ;
      LAYER metal2 ;
        RECT 256.600 98.800 257.000 99.200 ;
        RECT 256.600 98.200 256.900 98.800 ;
        RECT 256.600 97.800 257.000 98.200 ;
      LAYER metal3 ;
        RECT 267.800 99.100 268.200 99.200 ;
        RECT 256.600 98.800 268.200 99.100 ;
        RECT 256.600 98.200 256.900 98.800 ;
        RECT 256.600 97.800 257.000 98.200 ;
    END
  END dataout[4]
  PIN dataout[5]
    PORT
      LAYER metal1 ;
        RECT 261.400 166.200 261.800 169.900 ;
        RECT 261.500 165.100 261.800 166.200 ;
        RECT 261.400 161.100 261.800 165.100 ;
      LAYER via1 ;
        RECT 261.400 166.800 261.800 167.200 ;
      LAYER metal2 ;
        RECT 261.400 167.800 261.800 168.200 ;
        RECT 261.400 167.200 261.700 167.800 ;
        RECT 261.400 166.800 261.800 167.200 ;
      LAYER metal3 ;
        RECT 261.400 167.800 261.800 168.200 ;
        RECT 261.400 167.100 261.700 167.800 ;
        RECT 267.800 167.100 268.200 167.200 ;
        RECT 261.400 166.800 268.200 167.100 ;
    END
  END dataout[5]
  PIN dataout[6]
    PORT
      LAYER metal1 ;
        RECT 263.000 139.100 263.400 139.900 ;
        RECT 263.800 139.100 264.200 139.200 ;
        RECT 263.000 138.800 264.200 139.100 ;
        RECT 263.000 135.900 263.400 138.800 ;
        RECT 263.100 134.800 263.400 135.900 ;
        RECT 263.000 131.100 263.400 134.800 ;
      LAYER via1 ;
        RECT 263.800 138.800 264.200 139.200 ;
      LAYER metal2 ;
        RECT 263.800 139.100 264.200 139.200 ;
        RECT 264.600 139.100 265.000 139.200 ;
        RECT 263.800 138.800 265.000 139.100 ;
      LAYER via2 ;
        RECT 264.600 138.800 265.000 139.200 ;
      LAYER metal3 ;
        RECT 264.600 139.100 265.000 139.200 ;
        RECT 267.800 139.100 268.200 139.200 ;
        RECT 264.600 138.800 268.200 139.100 ;
    END
  END dataout[6]
  PIN dataout[7]
    PORT
      LAYER metal1 ;
        RECT 153.400 195.900 153.800 199.900 ;
        RECT 153.500 194.800 153.800 195.900 ;
        RECT 153.400 191.100 153.800 194.800 ;
      LAYER via1 ;
        RECT 153.400 198.800 153.800 199.200 ;
      LAYER metal2 ;
        RECT 152.600 242.800 153.000 243.200 ;
        RECT 152.600 240.200 152.900 242.800 ;
        RECT 152.600 239.800 153.000 240.200 ;
        RECT 153.400 202.800 153.800 203.200 ;
        RECT 153.400 199.200 153.700 202.800 ;
        RECT 153.400 198.800 153.800 199.200 ;
      LAYER metal3 ;
        RECT 152.600 240.100 153.000 240.200 ;
        RECT 153.400 240.100 153.800 240.200 ;
        RECT 152.600 239.800 153.800 240.100 ;
        RECT 152.600 203.100 153.000 203.200 ;
        RECT 153.400 203.100 153.800 203.200 ;
        RECT 152.600 202.800 153.800 203.100 ;
      LAYER via3 ;
        RECT 153.400 239.800 153.800 240.200 ;
      LAYER metal4 ;
        RECT 153.400 240.100 153.800 240.200 ;
        RECT 152.600 239.800 153.800 240.100 ;
        RECT 152.600 203.200 152.900 239.800 ;
        RECT 152.600 202.800 153.000 203.200 ;
    END
  END dataout[7]
  OBS
      LAYER metal1 ;
        RECT 1.400 235.600 1.800 239.900 ;
        RECT 3.000 235.600 3.400 239.900 ;
        RECT 4.600 235.600 5.000 239.900 ;
        RECT 6.200 235.600 6.600 239.900 ;
        RECT 8.600 235.600 9.000 239.900 ;
        RECT 10.200 235.600 10.600 239.900 ;
        RECT 11.800 235.600 12.200 239.900 ;
        RECT 13.400 235.600 13.800 239.900 ;
        RECT 15.800 235.600 16.200 239.900 ;
        RECT 17.400 235.600 17.800 239.900 ;
        RECT 19.000 235.600 19.400 239.900 ;
        RECT 20.600 235.600 21.000 239.900 ;
        RECT 1.400 235.200 2.300 235.600 ;
        RECT 3.000 235.200 4.100 235.600 ;
        RECT 4.600 235.200 5.700 235.600 ;
        RECT 6.200 235.200 7.400 235.600 ;
        RECT 8.600 235.200 9.500 235.600 ;
        RECT 10.200 235.200 11.300 235.600 ;
        RECT 11.800 235.200 12.900 235.600 ;
        RECT 13.400 235.200 14.600 235.600 ;
        RECT 1.900 234.500 2.300 235.200 ;
        RECT 3.700 234.500 4.100 235.200 ;
        RECT 5.300 234.500 5.700 235.200 ;
        RECT 1.900 234.100 3.200 234.500 ;
        RECT 3.700 234.100 4.900 234.500 ;
        RECT 5.300 234.100 6.600 234.500 ;
        RECT 1.900 233.800 2.300 234.100 ;
        RECT 3.700 233.800 4.100 234.100 ;
        RECT 5.300 233.800 5.700 234.100 ;
        RECT 7.000 233.800 7.400 235.200 ;
        RECT 9.100 234.500 9.500 235.200 ;
        RECT 10.900 234.500 11.300 235.200 ;
        RECT 12.500 234.500 12.900 235.200 ;
        RECT 9.100 234.100 10.400 234.500 ;
        RECT 10.900 234.100 12.100 234.500 ;
        RECT 12.500 234.100 13.800 234.500 ;
        RECT 9.100 233.800 9.500 234.100 ;
        RECT 10.900 233.800 11.300 234.100 ;
        RECT 12.500 233.800 12.900 234.100 ;
        RECT 14.200 233.800 14.600 235.200 ;
        RECT 1.400 233.400 2.300 233.800 ;
        RECT 3.000 233.400 4.100 233.800 ;
        RECT 4.600 233.400 5.700 233.800 ;
        RECT 6.200 233.400 7.400 233.800 ;
        RECT 8.600 233.400 9.500 233.800 ;
        RECT 10.200 233.400 11.300 233.800 ;
        RECT 11.800 233.400 12.900 233.800 ;
        RECT 13.400 233.400 14.600 233.800 ;
        RECT 15.000 235.200 16.200 235.600 ;
        RECT 16.700 235.200 17.800 235.600 ;
        RECT 18.300 235.200 19.400 235.600 ;
        RECT 20.100 235.200 21.000 235.600 ;
        RECT 23.000 235.600 23.400 239.900 ;
        RECT 24.600 235.600 25.000 239.900 ;
        RECT 26.200 235.600 26.600 239.900 ;
        RECT 27.800 235.600 28.200 239.900 ;
        RECT 30.200 235.600 30.600 239.900 ;
        RECT 31.800 235.600 32.200 239.900 ;
        RECT 33.400 235.600 33.800 239.900 ;
        RECT 35.000 235.600 35.400 239.900 ;
        RECT 37.400 235.600 37.800 239.900 ;
        RECT 39.000 235.600 39.400 239.900 ;
        RECT 40.600 235.600 41.000 239.900 ;
        RECT 42.200 235.600 42.600 239.900 ;
        RECT 43.800 235.700 44.200 239.900 ;
        RECT 46.000 238.200 46.400 239.900 ;
        RECT 45.400 237.900 46.400 238.200 ;
        RECT 48.200 237.900 48.600 239.900 ;
        RECT 50.300 237.900 50.900 239.900 ;
        RECT 45.400 237.500 45.800 237.900 ;
        RECT 48.200 237.600 48.500 237.900 ;
        RECT 47.100 237.300 48.900 237.600 ;
        RECT 50.200 237.500 50.600 237.900 ;
        RECT 47.100 237.200 47.500 237.300 ;
        RECT 48.500 237.200 48.900 237.300 ;
        RECT 45.400 236.500 45.800 236.600 ;
        RECT 47.700 236.500 48.100 236.600 ;
        RECT 45.400 236.200 48.100 236.500 ;
        RECT 48.400 236.500 49.500 236.800 ;
        RECT 48.400 235.900 48.700 236.500 ;
        RECT 49.100 236.400 49.500 236.500 ;
        RECT 50.300 236.600 51.000 237.000 ;
        RECT 50.300 236.100 50.600 236.600 ;
        RECT 46.300 235.700 48.700 235.900 ;
        RECT 43.800 235.600 48.700 235.700 ;
        RECT 49.400 235.800 50.600 236.100 ;
        RECT 23.000 235.200 23.900 235.600 ;
        RECT 24.600 235.200 25.700 235.600 ;
        RECT 26.200 235.200 27.300 235.600 ;
        RECT 27.800 235.200 29.000 235.600 ;
        RECT 30.200 235.200 31.100 235.600 ;
        RECT 31.800 235.200 32.900 235.600 ;
        RECT 33.400 235.200 34.500 235.600 ;
        RECT 35.000 235.200 36.200 235.600 ;
        RECT 37.400 235.200 38.300 235.600 ;
        RECT 39.000 235.200 40.100 235.600 ;
        RECT 40.600 235.200 41.700 235.600 ;
        RECT 42.200 235.200 43.400 235.600 ;
        RECT 43.800 235.500 46.700 235.600 ;
        RECT 43.800 235.400 46.600 235.500 ;
        RECT 15.000 233.800 15.400 235.200 ;
        RECT 16.700 234.500 17.100 235.200 ;
        RECT 18.300 234.500 18.700 235.200 ;
        RECT 20.100 234.500 20.500 235.200 ;
        RECT 23.500 234.500 23.900 235.200 ;
        RECT 25.300 234.500 25.700 235.200 ;
        RECT 26.900 234.500 27.300 235.200 ;
        RECT 15.800 234.100 17.100 234.500 ;
        RECT 17.500 234.100 18.700 234.500 ;
        RECT 19.200 234.100 20.500 234.500 ;
        RECT 20.900 234.100 21.800 234.500 ;
        RECT 16.700 233.800 17.100 234.100 ;
        RECT 18.300 233.800 18.700 234.100 ;
        RECT 20.100 233.800 20.500 234.100 ;
        RECT 21.400 233.800 21.800 234.100 ;
        RECT 23.500 234.100 24.800 234.500 ;
        RECT 25.300 234.100 26.500 234.500 ;
        RECT 26.900 234.100 28.200 234.500 ;
        RECT 23.500 233.800 23.900 234.100 ;
        RECT 25.300 233.800 25.700 234.100 ;
        RECT 26.900 233.800 27.300 234.100 ;
        RECT 28.600 233.800 29.000 235.200 ;
        RECT 30.700 234.500 31.100 235.200 ;
        RECT 32.500 234.500 32.900 235.200 ;
        RECT 34.100 234.500 34.500 235.200 ;
        RECT 29.400 234.100 30.300 234.500 ;
        RECT 30.700 234.100 32.000 234.500 ;
        RECT 32.500 234.100 33.700 234.500 ;
        RECT 34.100 234.100 35.400 234.500 ;
        RECT 29.400 233.800 29.800 234.100 ;
        RECT 30.700 233.800 31.100 234.100 ;
        RECT 32.500 233.800 32.900 234.100 ;
        RECT 34.100 233.800 34.500 234.100 ;
        RECT 35.800 233.800 36.200 235.200 ;
        RECT 37.900 234.500 38.300 235.200 ;
        RECT 39.700 234.500 40.100 235.200 ;
        RECT 41.300 234.500 41.700 235.200 ;
        RECT 36.600 234.100 37.500 234.500 ;
        RECT 37.900 234.100 39.200 234.500 ;
        RECT 39.700 234.100 40.900 234.500 ;
        RECT 41.300 234.100 42.600 234.500 ;
        RECT 36.600 233.800 37.000 234.100 ;
        RECT 37.900 233.800 38.300 234.100 ;
        RECT 39.700 233.800 40.100 234.100 ;
        RECT 41.300 233.800 41.700 234.100 ;
        RECT 43.000 233.800 43.400 235.200 ;
        RECT 47.000 235.100 47.400 235.200 ;
        RECT 44.900 234.800 47.400 235.100 ;
        RECT 44.900 234.700 45.300 234.800 ;
        RECT 45.700 234.200 46.100 234.300 ;
        RECT 49.400 234.200 49.700 235.800 ;
        RECT 52.600 235.600 53.000 239.900 ;
        RECT 50.900 235.300 53.000 235.600 ;
        RECT 50.900 235.200 51.300 235.300 ;
        RECT 51.700 234.900 52.100 235.000 ;
        RECT 50.200 234.600 52.100 234.900 ;
        RECT 50.200 234.500 50.600 234.600 ;
        RECT 44.200 233.900 49.800 234.200 ;
        RECT 44.200 233.800 45.000 233.900 ;
        RECT 15.000 233.400 16.200 233.800 ;
        RECT 16.700 233.400 17.800 233.800 ;
        RECT 18.300 233.400 19.400 233.800 ;
        RECT 20.100 233.400 21.000 233.800 ;
        RECT 1.400 231.100 1.800 233.400 ;
        RECT 3.000 231.100 3.400 233.400 ;
        RECT 4.600 231.100 5.000 233.400 ;
        RECT 6.200 231.100 6.600 233.400 ;
        RECT 8.600 231.100 9.000 233.400 ;
        RECT 10.200 231.100 10.600 233.400 ;
        RECT 11.800 231.100 12.200 233.400 ;
        RECT 13.400 231.100 13.800 233.400 ;
        RECT 15.800 231.100 16.200 233.400 ;
        RECT 17.400 231.100 17.800 233.400 ;
        RECT 19.000 231.100 19.400 233.400 ;
        RECT 20.600 231.100 21.000 233.400 ;
        RECT 23.000 233.400 23.900 233.800 ;
        RECT 24.600 233.400 25.700 233.800 ;
        RECT 26.200 233.400 27.300 233.800 ;
        RECT 27.800 233.400 29.000 233.800 ;
        RECT 30.200 233.400 31.100 233.800 ;
        RECT 31.800 233.400 32.900 233.800 ;
        RECT 33.400 233.400 34.500 233.800 ;
        RECT 35.000 233.400 36.200 233.800 ;
        RECT 37.400 233.400 38.300 233.800 ;
        RECT 39.000 233.400 40.100 233.800 ;
        RECT 40.600 233.400 41.700 233.800 ;
        RECT 42.200 233.400 43.400 233.800 ;
        RECT 23.000 231.100 23.400 233.400 ;
        RECT 24.600 231.100 25.000 233.400 ;
        RECT 26.200 231.100 26.600 233.400 ;
        RECT 27.800 231.100 28.200 233.400 ;
        RECT 30.200 231.100 30.600 233.400 ;
        RECT 31.800 231.100 32.200 233.400 ;
        RECT 33.400 231.100 33.800 233.400 ;
        RECT 35.000 231.100 35.400 233.400 ;
        RECT 37.400 231.100 37.800 233.400 ;
        RECT 39.000 231.100 39.400 233.400 ;
        RECT 40.600 231.100 41.000 233.400 ;
        RECT 42.200 231.100 42.600 233.400 ;
        RECT 43.800 231.100 44.200 233.500 ;
        RECT 46.300 232.800 46.600 233.900 ;
        RECT 49.100 233.800 49.800 233.900 ;
        RECT 52.600 233.600 53.000 235.300 ;
        RECT 55.800 235.600 56.200 239.900 ;
        RECT 57.400 235.600 57.800 239.900 ;
        RECT 59.000 235.600 59.400 239.900 ;
        RECT 60.600 235.600 61.000 239.900 ;
        RECT 63.500 236.200 63.900 239.900 ;
        RECT 64.200 236.800 64.600 237.200 ;
        RECT 64.300 236.200 64.600 236.800 ;
        RECT 63.500 235.900 64.000 236.200 ;
        RECT 64.300 235.900 65.000 236.200 ;
        RECT 55.800 235.200 56.700 235.600 ;
        RECT 57.400 235.200 58.500 235.600 ;
        RECT 59.000 235.200 60.100 235.600 ;
        RECT 60.600 235.200 61.800 235.600 ;
        RECT 56.300 234.500 56.700 235.200 ;
        RECT 58.100 234.500 58.500 235.200 ;
        RECT 59.700 234.500 60.100 235.200 ;
        RECT 53.400 234.100 53.800 234.200 ;
        RECT 55.000 234.100 55.900 234.500 ;
        RECT 56.300 234.100 57.600 234.500 ;
        RECT 58.100 234.100 59.300 234.500 ;
        RECT 59.700 234.100 61.000 234.500 ;
        RECT 53.400 233.800 55.400 234.100 ;
        RECT 56.300 233.800 56.700 234.100 ;
        RECT 58.100 233.800 58.500 234.100 ;
        RECT 59.700 233.800 60.100 234.100 ;
        RECT 61.400 233.800 61.800 235.200 ;
        RECT 62.200 235.100 62.600 235.200 ;
        RECT 63.000 235.100 63.400 235.200 ;
        RECT 62.200 234.800 63.400 235.100 ;
        RECT 63.000 234.400 63.400 234.800 ;
        RECT 63.700 234.200 64.000 235.900 ;
        RECT 64.600 235.800 65.000 235.900 ;
        RECT 65.400 235.800 65.800 236.600 ;
        RECT 64.600 235.100 64.900 235.800 ;
        RECT 66.200 235.100 66.600 239.900 ;
        RECT 67.800 235.700 68.200 239.900 ;
        RECT 70.000 238.200 70.400 239.900 ;
        RECT 69.400 237.900 70.400 238.200 ;
        RECT 72.200 237.900 72.600 239.900 ;
        RECT 74.300 237.900 74.900 239.900 ;
        RECT 69.400 237.500 69.800 237.900 ;
        RECT 72.200 237.600 72.500 237.900 ;
        RECT 71.100 237.300 72.900 237.600 ;
        RECT 74.200 237.500 74.600 237.900 ;
        RECT 71.100 237.200 71.500 237.300 ;
        RECT 72.500 237.200 72.900 237.300 ;
        RECT 69.400 236.500 69.800 236.600 ;
        RECT 71.700 236.500 72.100 236.600 ;
        RECT 69.400 236.200 72.100 236.500 ;
        RECT 72.400 236.500 73.500 236.800 ;
        RECT 72.400 235.900 72.700 236.500 ;
        RECT 73.100 236.400 73.500 236.500 ;
        RECT 74.300 236.600 75.000 237.000 ;
        RECT 74.300 236.100 74.600 236.600 ;
        RECT 70.300 235.700 72.700 235.900 ;
        RECT 67.800 235.600 72.700 235.700 ;
        RECT 73.400 235.800 74.600 236.100 ;
        RECT 67.800 235.500 70.700 235.600 ;
        RECT 67.800 235.400 70.600 235.500 ;
        RECT 71.000 235.100 71.400 235.200 ;
        RECT 64.600 234.800 66.600 235.100 ;
        RECT 62.200 234.100 62.600 234.200 ;
        RECT 62.200 233.800 63.000 234.100 ;
        RECT 63.700 233.800 65.000 234.200 ;
        RECT 51.100 233.300 53.000 233.600 ;
        RECT 51.100 233.200 51.500 233.300 ;
        RECT 45.400 232.100 45.800 232.500 ;
        RECT 46.200 232.400 46.600 232.800 ;
        RECT 47.100 232.700 47.500 232.800 ;
        RECT 47.100 232.400 48.500 232.700 ;
        RECT 48.200 232.100 48.500 232.400 ;
        RECT 50.200 232.100 50.600 232.500 ;
        RECT 45.400 231.800 46.400 232.100 ;
        RECT 46.000 231.100 46.400 231.800 ;
        RECT 48.200 231.100 48.600 232.100 ;
        RECT 50.200 231.800 50.900 232.100 ;
        RECT 50.300 231.100 50.900 231.800 ;
        RECT 52.600 231.100 53.000 233.300 ;
        RECT 55.800 233.400 56.700 233.800 ;
        RECT 57.400 233.400 58.500 233.800 ;
        RECT 59.000 233.400 60.100 233.800 ;
        RECT 60.600 233.400 61.800 233.800 ;
        RECT 62.600 233.600 63.000 233.800 ;
        RECT 55.800 231.100 56.200 233.400 ;
        RECT 57.400 231.100 57.800 233.400 ;
        RECT 59.000 231.100 59.400 233.400 ;
        RECT 60.600 231.100 61.000 233.400 ;
        RECT 62.300 233.100 64.100 233.300 ;
        RECT 64.600 233.100 64.900 233.800 ;
        RECT 66.200 233.100 66.600 234.800 ;
        RECT 68.900 234.800 71.400 235.100 ;
        RECT 68.900 234.700 69.300 234.800 ;
        RECT 69.700 234.200 70.100 234.300 ;
        RECT 73.400 234.200 73.700 235.800 ;
        RECT 76.600 235.600 77.000 239.900 ;
        RECT 74.900 235.300 77.000 235.600 ;
        RECT 77.400 235.700 77.800 239.900 ;
        RECT 79.600 238.200 80.000 239.900 ;
        RECT 79.000 237.900 80.000 238.200 ;
        RECT 81.800 237.900 82.200 239.900 ;
        RECT 83.900 237.900 84.500 239.900 ;
        RECT 79.000 237.500 79.400 237.900 ;
        RECT 81.800 237.600 82.100 237.900 ;
        RECT 80.700 237.300 82.500 237.600 ;
        RECT 83.800 237.500 84.200 237.900 ;
        RECT 80.700 237.200 81.100 237.300 ;
        RECT 82.100 237.200 82.500 237.300 ;
        RECT 79.000 236.500 79.400 236.600 ;
        RECT 81.300 236.500 81.700 236.600 ;
        RECT 79.000 236.200 81.700 236.500 ;
        RECT 82.000 236.500 83.100 236.800 ;
        RECT 82.000 235.900 82.300 236.500 ;
        RECT 82.700 236.400 83.100 236.500 ;
        RECT 83.900 236.600 84.600 237.000 ;
        RECT 83.900 236.100 84.200 236.600 ;
        RECT 79.900 235.700 82.300 235.900 ;
        RECT 77.400 235.600 82.300 235.700 ;
        RECT 83.000 235.800 84.200 236.100 ;
        RECT 77.400 235.500 80.300 235.600 ;
        RECT 77.400 235.400 80.200 235.500 ;
        RECT 74.900 235.200 75.300 235.300 ;
        RECT 75.700 234.900 76.100 235.000 ;
        RECT 74.200 234.600 76.100 234.900 ;
        RECT 74.200 234.500 74.600 234.600 ;
        RECT 67.000 233.400 67.400 234.200 ;
        RECT 68.200 233.900 73.700 234.200 ;
        RECT 68.200 233.800 69.000 233.900 ;
        RECT 62.200 233.000 64.200 233.100 ;
        RECT 62.200 231.100 62.600 233.000 ;
        RECT 63.800 231.100 64.200 233.000 ;
        RECT 64.600 231.100 65.000 233.100 ;
        RECT 65.700 232.800 66.600 233.100 ;
        RECT 65.700 231.100 66.100 232.800 ;
        RECT 67.800 231.100 68.200 233.500 ;
        RECT 70.300 232.800 70.600 233.900 ;
        RECT 73.100 233.800 73.500 233.900 ;
        RECT 76.600 233.600 77.000 235.300 ;
        RECT 83.000 235.200 83.300 235.800 ;
        RECT 86.200 235.600 86.600 239.900 ;
        RECT 84.500 235.300 86.600 235.600 ;
        RECT 84.500 235.200 84.900 235.300 ;
        RECT 80.600 235.100 81.000 235.200 ;
        RECT 78.500 234.800 81.000 235.100 ;
        RECT 83.000 234.800 83.400 235.200 ;
        RECT 85.300 234.900 85.700 235.000 ;
        RECT 78.500 234.700 78.900 234.800 ;
        RECT 79.300 234.200 79.700 234.300 ;
        RECT 83.000 234.200 83.300 234.800 ;
        RECT 83.800 234.600 85.700 234.900 ;
        RECT 83.800 234.500 84.200 234.600 ;
        RECT 77.800 233.900 83.300 234.200 ;
        RECT 77.800 233.800 78.600 233.900 ;
        RECT 75.100 233.300 77.000 233.600 ;
        RECT 75.100 233.200 75.500 233.300 ;
        RECT 69.400 232.100 69.800 232.500 ;
        RECT 70.200 232.400 70.600 232.800 ;
        RECT 71.100 232.700 71.500 232.800 ;
        RECT 71.100 232.400 72.500 232.700 ;
        RECT 72.200 232.100 72.500 232.400 ;
        RECT 74.200 232.100 74.600 232.500 ;
        RECT 69.400 231.800 70.400 232.100 ;
        RECT 70.000 231.100 70.400 231.800 ;
        RECT 72.200 231.100 72.600 232.100 ;
        RECT 74.200 231.800 74.900 232.100 ;
        RECT 74.300 231.100 74.900 231.800 ;
        RECT 76.600 231.100 77.000 233.300 ;
        RECT 77.400 231.100 77.800 233.500 ;
        RECT 79.900 232.800 80.200 233.900 ;
        RECT 82.700 233.800 83.100 233.900 ;
        RECT 86.200 233.600 86.600 235.300 ;
        RECT 84.700 233.300 86.600 233.600 ;
        RECT 84.700 233.200 85.100 233.300 ;
        RECT 86.200 233.100 86.600 233.300 ;
        RECT 87.800 235.100 88.200 239.900 ;
        RECT 90.500 236.400 90.900 239.900 ;
        RECT 92.600 237.500 93.000 239.500 ;
        RECT 90.100 236.100 90.900 236.400 ;
        RECT 89.400 235.100 89.800 235.600 ;
        RECT 87.800 234.800 89.800 235.100 ;
        RECT 87.000 233.100 87.400 233.200 ;
        RECT 86.200 232.800 87.400 233.100 ;
        RECT 79.000 232.100 79.400 232.500 ;
        RECT 79.800 232.400 80.200 232.800 ;
        RECT 80.700 232.700 81.100 232.800 ;
        RECT 80.700 232.400 82.100 232.700 ;
        RECT 81.800 232.100 82.100 232.400 ;
        RECT 83.800 232.100 84.200 232.500 ;
        RECT 79.000 231.800 80.000 232.100 ;
        RECT 79.600 231.100 80.000 231.800 ;
        RECT 81.800 231.100 82.200 232.100 ;
        RECT 83.800 231.800 84.500 232.100 ;
        RECT 83.900 231.100 84.500 231.800 ;
        RECT 86.200 231.100 86.600 232.800 ;
        RECT 87.000 232.400 87.400 232.800 ;
        RECT 87.800 231.100 88.200 234.800 ;
        RECT 90.100 234.200 90.400 236.100 ;
        RECT 92.700 235.800 93.000 237.500 ;
        RECT 91.100 235.500 93.000 235.800 ;
        RECT 93.400 235.700 93.800 239.900 ;
        RECT 95.600 238.200 96.000 239.900 ;
        RECT 95.000 237.900 96.000 238.200 ;
        RECT 97.800 237.900 98.200 239.900 ;
        RECT 99.900 237.900 100.500 239.900 ;
        RECT 95.000 237.500 95.400 237.900 ;
        RECT 97.800 237.600 98.100 237.900 ;
        RECT 96.700 237.300 98.500 237.600 ;
        RECT 99.800 237.500 100.200 237.900 ;
        RECT 96.700 237.200 97.100 237.300 ;
        RECT 98.100 237.200 98.500 237.300 ;
        RECT 95.000 236.500 95.400 236.600 ;
        RECT 97.300 236.500 97.700 236.600 ;
        RECT 95.000 236.200 97.700 236.500 ;
        RECT 98.000 236.500 99.100 236.800 ;
        RECT 98.000 235.900 98.300 236.500 ;
        RECT 98.700 236.400 99.100 236.500 ;
        RECT 99.900 236.600 100.600 237.000 ;
        RECT 99.900 236.100 100.200 236.600 ;
        RECT 95.900 235.700 98.300 235.900 ;
        RECT 93.400 235.600 98.300 235.700 ;
        RECT 99.000 235.800 100.200 236.100 ;
        RECT 93.400 235.500 96.300 235.600 ;
        RECT 91.100 234.500 91.400 235.500 ;
        RECT 93.400 235.400 96.200 235.500 ;
        RECT 88.600 234.100 89.000 234.200 ;
        RECT 89.400 234.100 90.400 234.200 ;
        RECT 90.700 234.100 91.400 234.500 ;
        RECT 91.800 234.400 92.200 235.200 ;
        RECT 92.600 234.400 93.000 235.200 ;
        RECT 96.600 235.100 97.000 235.200 ;
        RECT 97.400 235.100 97.800 235.200 ;
        RECT 94.500 234.800 97.800 235.100 ;
        RECT 94.500 234.700 94.900 234.800 ;
        RECT 95.300 234.200 95.700 234.300 ;
        RECT 99.000 234.200 99.300 235.800 ;
        RECT 102.200 235.600 102.600 239.900 ;
        RECT 103.400 236.800 103.800 237.200 ;
        RECT 103.400 236.200 103.700 236.800 ;
        RECT 104.100 236.200 104.500 239.900 ;
        RECT 103.000 235.900 103.700 236.200 ;
        RECT 104.000 235.900 104.500 236.200 ;
        RECT 103.000 235.800 103.400 235.900 ;
        RECT 100.500 235.300 102.600 235.600 ;
        RECT 100.500 235.200 100.900 235.300 ;
        RECT 101.300 234.900 101.700 235.000 ;
        RECT 99.800 234.600 101.700 234.900 ;
        RECT 99.800 234.500 100.200 234.600 ;
        RECT 88.600 233.800 90.400 234.100 ;
        RECT 90.100 233.500 90.400 233.800 ;
        RECT 90.900 233.900 91.400 234.100 ;
        RECT 93.800 233.900 99.300 234.200 ;
        RECT 90.900 233.600 93.000 233.900 ;
        RECT 93.800 233.800 94.600 233.900 ;
        RECT 90.100 233.300 90.500 233.500 ;
        RECT 90.100 233.000 90.900 233.300 ;
        RECT 90.500 231.500 90.900 233.000 ;
        RECT 92.700 232.500 93.000 233.600 ;
        RECT 92.600 231.500 93.000 232.500 ;
        RECT 93.400 231.100 93.800 233.500 ;
        RECT 95.900 232.800 96.200 233.900 ;
        RECT 97.400 233.800 97.800 233.900 ;
        RECT 98.700 233.800 99.100 233.900 ;
        RECT 102.200 233.600 102.600 235.300 ;
        RECT 103.000 235.100 103.400 235.200 ;
        RECT 104.000 235.100 104.300 235.900 ;
        RECT 107.800 235.800 108.200 236.600 ;
        RECT 108.600 236.100 109.000 239.900 ;
        RECT 111.500 236.200 111.900 239.900 ;
        RECT 112.200 236.800 112.600 237.200 ;
        RECT 112.300 236.200 112.600 236.800 ;
        RECT 109.400 236.100 109.800 236.200 ;
        RECT 108.600 235.800 109.800 236.100 ;
        RECT 111.500 235.900 112.000 236.200 ;
        RECT 112.300 235.900 113.000 236.200 ;
        RECT 103.000 234.800 104.300 235.100 ;
        RECT 104.000 234.200 104.300 234.800 ;
        RECT 104.600 235.100 105.000 235.200 ;
        RECT 107.800 235.100 108.200 235.200 ;
        RECT 104.600 234.800 108.200 235.100 ;
        RECT 104.600 234.400 105.000 234.800 ;
        RECT 103.000 233.800 104.300 234.200 ;
        RECT 105.400 234.100 105.800 234.200 ;
        RECT 107.800 234.100 108.200 234.200 ;
        RECT 105.000 233.800 108.200 234.100 ;
        RECT 100.700 233.300 102.600 233.600 ;
        RECT 100.700 233.200 101.100 233.300 ;
        RECT 95.000 232.100 95.400 232.500 ;
        RECT 95.800 232.400 96.200 232.800 ;
        RECT 96.700 232.700 97.100 232.800 ;
        RECT 96.700 232.400 98.100 232.700 ;
        RECT 97.800 232.100 98.100 232.400 ;
        RECT 99.800 232.100 100.200 232.500 ;
        RECT 95.000 231.800 96.000 232.100 ;
        RECT 95.600 231.100 96.000 231.800 ;
        RECT 97.800 231.100 98.200 232.100 ;
        RECT 99.800 231.800 100.500 232.100 ;
        RECT 99.900 231.100 100.500 231.800 ;
        RECT 102.200 231.100 102.600 233.300 ;
        RECT 103.100 233.100 103.400 233.800 ;
        RECT 105.000 233.600 105.400 233.800 ;
        RECT 103.900 233.100 105.700 233.300 ;
        RECT 108.600 233.100 109.000 235.800 ;
        RECT 111.000 234.400 111.400 235.200 ;
        RECT 111.700 234.200 112.000 235.900 ;
        RECT 112.600 235.800 113.000 235.900 ;
        RECT 113.400 235.700 113.800 239.900 ;
        RECT 115.600 238.200 116.000 239.900 ;
        RECT 115.000 237.900 116.000 238.200 ;
        RECT 117.800 237.900 118.200 239.900 ;
        RECT 119.900 237.900 120.500 239.900 ;
        RECT 115.000 237.500 115.400 237.900 ;
        RECT 117.800 237.600 118.100 237.900 ;
        RECT 116.700 237.300 118.500 237.600 ;
        RECT 119.800 237.500 120.200 237.900 ;
        RECT 116.700 237.200 117.100 237.300 ;
        RECT 118.100 237.200 118.500 237.300 ;
        RECT 115.000 236.500 115.400 236.600 ;
        RECT 117.300 236.500 117.700 236.600 ;
        RECT 115.000 236.200 117.700 236.500 ;
        RECT 118.000 236.500 119.100 236.800 ;
        RECT 118.000 235.900 118.300 236.500 ;
        RECT 118.700 236.400 119.100 236.500 ;
        RECT 119.900 236.600 120.600 237.000 ;
        RECT 119.900 236.100 120.200 236.600 ;
        RECT 115.900 235.700 118.300 235.900 ;
        RECT 113.400 235.600 118.300 235.700 ;
        RECT 119.000 235.800 120.200 236.100 ;
        RECT 113.400 235.500 116.300 235.600 ;
        RECT 113.400 235.400 116.200 235.500 ;
        RECT 116.600 235.100 117.000 235.200 ;
        RECT 118.200 235.100 118.600 235.200 ;
        RECT 114.500 234.800 118.600 235.100 ;
        RECT 114.500 234.700 114.900 234.800 ;
        RECT 115.300 234.200 115.700 234.300 ;
        RECT 119.000 234.200 119.300 235.800 ;
        RECT 122.200 235.600 122.600 239.900 ;
        RECT 124.300 236.200 124.700 239.900 ;
        RECT 125.000 236.800 125.400 237.200 ;
        RECT 125.100 236.200 125.400 236.800 ;
        RECT 124.300 235.900 124.800 236.200 ;
        RECT 125.100 235.900 125.800 236.200 ;
        RECT 120.500 235.300 122.600 235.600 ;
        RECT 120.500 235.200 120.900 235.300 ;
        RECT 121.300 234.900 121.700 235.000 ;
        RECT 119.800 234.600 121.700 234.900 ;
        RECT 119.800 234.500 120.200 234.600 ;
        RECT 109.400 233.400 109.800 234.200 ;
        RECT 110.200 234.100 110.600 234.200 ;
        RECT 110.200 233.800 111.000 234.100 ;
        RECT 111.700 233.800 113.000 234.200 ;
        RECT 113.800 233.900 119.300 234.200 ;
        RECT 113.800 233.800 114.600 233.900 ;
        RECT 110.600 233.600 111.000 233.800 ;
        RECT 110.300 233.100 112.100 233.300 ;
        RECT 112.600 233.100 112.900 233.800 ;
        RECT 103.000 231.100 103.400 233.100 ;
        RECT 103.800 233.000 105.800 233.100 ;
        RECT 103.800 231.100 104.200 233.000 ;
        RECT 105.400 231.100 105.800 233.000 ;
        RECT 108.100 232.800 109.000 233.100 ;
        RECT 110.200 233.000 112.200 233.100 ;
        RECT 108.100 231.100 108.500 232.800 ;
        RECT 110.200 231.100 110.600 233.000 ;
        RECT 111.800 231.100 112.200 233.000 ;
        RECT 112.600 231.100 113.000 233.100 ;
        RECT 113.400 231.100 113.800 233.500 ;
        RECT 115.900 233.200 116.200 233.900 ;
        RECT 118.700 233.800 119.100 233.900 ;
        RECT 122.200 233.600 122.600 235.300 ;
        RECT 124.500 235.200 124.800 235.900 ;
        RECT 125.400 235.800 125.800 235.900 ;
        RECT 126.200 235.800 126.600 236.600 ;
        RECT 123.800 234.400 124.200 235.200 ;
        RECT 124.500 234.800 125.000 235.200 ;
        RECT 125.400 235.100 125.700 235.800 ;
        RECT 127.000 235.100 127.400 239.900 ;
        RECT 128.600 235.700 129.000 239.900 ;
        RECT 130.800 238.200 131.200 239.900 ;
        RECT 130.200 237.900 131.200 238.200 ;
        RECT 133.000 237.900 133.400 239.900 ;
        RECT 135.100 237.900 135.700 239.900 ;
        RECT 130.200 237.500 130.600 237.900 ;
        RECT 133.000 237.600 133.300 237.900 ;
        RECT 131.900 237.300 133.700 237.600 ;
        RECT 135.000 237.500 135.400 237.900 ;
        RECT 131.900 237.200 132.300 237.300 ;
        RECT 133.300 237.200 133.700 237.300 ;
        RECT 137.400 237.100 137.800 239.900 ;
        RECT 138.200 237.100 138.600 237.200 ;
        RECT 130.200 236.500 130.600 236.600 ;
        RECT 132.500 236.500 132.900 236.600 ;
        RECT 130.200 236.200 132.900 236.500 ;
        RECT 133.200 236.500 134.300 236.800 ;
        RECT 133.200 235.900 133.500 236.500 ;
        RECT 133.900 236.400 134.300 236.500 ;
        RECT 135.100 236.600 135.800 237.000 ;
        RECT 137.400 236.800 138.600 237.100 ;
        RECT 135.100 236.100 135.400 236.600 ;
        RECT 131.100 235.700 133.500 235.900 ;
        RECT 128.600 235.600 133.500 235.700 ;
        RECT 134.200 235.800 135.400 236.100 ;
        RECT 128.600 235.500 131.500 235.600 ;
        RECT 128.600 235.400 131.400 235.500 ;
        RECT 131.800 235.100 132.200 235.200 ;
        RECT 125.400 234.800 127.400 235.100 ;
        RECT 124.500 234.200 124.800 234.800 ;
        RECT 123.000 234.100 123.400 234.200 ;
        RECT 123.000 233.800 123.800 234.100 ;
        RECT 124.500 233.800 125.800 234.200 ;
        RECT 123.400 233.600 123.800 233.800 ;
        RECT 120.700 233.300 122.600 233.600 ;
        RECT 120.700 233.200 121.100 233.300 ;
        RECT 115.000 232.100 115.400 232.500 ;
        RECT 115.800 232.400 116.200 233.200 ;
        RECT 116.700 232.700 117.100 232.800 ;
        RECT 116.700 232.400 118.100 232.700 ;
        RECT 117.800 232.100 118.100 232.400 ;
        RECT 119.800 232.100 120.200 232.500 ;
        RECT 115.000 231.800 116.000 232.100 ;
        RECT 115.600 231.100 116.000 231.800 ;
        RECT 117.800 231.100 118.200 232.100 ;
        RECT 119.800 231.800 120.500 232.100 ;
        RECT 119.900 231.100 120.500 231.800 ;
        RECT 122.200 231.100 122.600 233.300 ;
        RECT 123.100 233.100 124.900 233.300 ;
        RECT 125.400 233.100 125.700 233.800 ;
        RECT 127.000 233.100 127.400 234.800 ;
        RECT 129.700 234.800 132.200 235.100 ;
        RECT 129.700 234.700 130.100 234.800 ;
        RECT 130.500 234.200 130.900 234.300 ;
        RECT 134.200 234.200 134.500 235.800 ;
        RECT 137.400 235.600 137.800 236.800 ;
        RECT 135.700 235.300 137.800 235.600 ;
        RECT 135.700 235.200 136.100 235.300 ;
        RECT 136.500 234.900 136.900 235.000 ;
        RECT 135.000 234.600 136.900 234.900 ;
        RECT 135.000 234.500 135.400 234.600 ;
        RECT 127.800 233.400 128.200 234.200 ;
        RECT 129.000 233.900 134.500 234.200 ;
        RECT 129.000 233.800 129.800 233.900 ;
        RECT 123.000 233.000 125.000 233.100 ;
        RECT 123.000 231.100 123.400 233.000 ;
        RECT 124.600 231.100 125.000 233.000 ;
        RECT 125.400 231.100 125.800 233.100 ;
        RECT 126.500 232.800 127.400 233.100 ;
        RECT 126.500 231.100 126.900 232.800 ;
        RECT 128.600 231.100 129.000 233.500 ;
        RECT 131.100 232.800 131.400 233.900 ;
        RECT 133.900 233.800 134.300 233.900 ;
        RECT 137.400 233.600 137.800 235.300 ;
        RECT 139.000 235.100 139.400 239.900 ;
        RECT 141.000 236.800 141.400 237.200 ;
        RECT 139.800 235.800 140.200 236.600 ;
        RECT 141.000 236.200 141.300 236.800 ;
        RECT 141.700 236.200 142.100 239.900 ;
        RECT 140.600 235.900 141.300 236.200 ;
        RECT 141.600 235.900 142.100 236.200 ;
        RECT 143.800 236.200 144.200 239.900 ;
        RECT 145.400 236.200 145.800 239.900 ;
        RECT 143.800 235.900 145.800 236.200 ;
        RECT 140.600 235.800 141.000 235.900 ;
        RECT 140.600 235.100 140.900 235.800 ;
        RECT 139.000 234.800 140.900 235.100 ;
        RECT 135.900 233.300 137.800 233.600 ;
        RECT 138.200 233.400 138.600 234.200 ;
        RECT 135.900 233.200 136.300 233.300 ;
        RECT 130.200 232.100 130.600 232.500 ;
        RECT 131.000 232.400 131.400 232.800 ;
        RECT 131.900 232.700 132.300 232.800 ;
        RECT 131.900 232.400 133.300 232.700 ;
        RECT 133.000 232.100 133.300 232.400 ;
        RECT 135.000 232.100 135.400 232.500 ;
        RECT 130.200 231.800 131.200 232.100 ;
        RECT 130.800 231.100 131.200 231.800 ;
        RECT 133.000 231.100 133.400 232.100 ;
        RECT 135.000 231.800 135.700 232.100 ;
        RECT 135.100 231.100 135.700 231.800 ;
        RECT 137.400 231.100 137.800 233.300 ;
        RECT 139.000 233.100 139.400 234.800 ;
        RECT 141.600 234.200 141.900 235.900 ;
        RECT 146.200 235.800 146.600 239.900 ;
        RECT 148.300 236.300 148.700 239.900 ;
        RECT 147.800 235.900 148.700 236.300 ;
        RECT 144.200 235.200 144.600 235.400 ;
        RECT 146.200 235.200 146.500 235.800 ;
        RECT 142.200 234.400 142.600 235.200 ;
        RECT 143.800 235.100 144.600 235.200 ;
        RECT 143.000 234.900 144.600 235.100 ;
        RECT 145.400 234.900 146.600 235.200 ;
        RECT 143.000 234.800 144.200 234.900 ;
        RECT 139.800 234.100 140.200 234.200 ;
        RECT 140.600 234.100 141.900 234.200 ;
        RECT 143.000 234.200 143.300 234.800 ;
        RECT 143.000 234.100 143.400 234.200 ;
        RECT 139.800 233.800 141.900 234.100 ;
        RECT 142.600 233.800 143.400 234.100 ;
        RECT 144.600 233.800 145.000 234.600 ;
        RECT 140.700 233.100 141.000 233.800 ;
        RECT 142.600 233.600 143.000 233.800 ;
        RECT 141.500 233.100 143.300 233.300 ;
        RECT 145.400 233.100 145.700 234.900 ;
        RECT 146.200 234.800 146.600 234.900 ;
        RECT 147.900 234.200 148.200 235.900 ;
        RECT 149.400 235.600 149.800 239.900 ;
        RECT 151.500 237.900 152.100 239.900 ;
        RECT 153.800 237.900 154.200 239.900 ;
        RECT 156.000 238.200 156.400 239.900 ;
        RECT 156.000 237.900 157.000 238.200 ;
        RECT 151.800 237.500 152.200 237.900 ;
        RECT 153.900 237.600 154.200 237.900 ;
        RECT 153.500 237.300 155.300 237.600 ;
        RECT 156.600 237.500 157.000 237.900 ;
        RECT 153.500 237.200 153.900 237.300 ;
        RECT 154.900 237.200 155.300 237.300 ;
        RECT 151.400 236.600 152.100 237.000 ;
        RECT 151.800 236.100 152.100 236.600 ;
        RECT 152.900 236.500 154.000 236.800 ;
        RECT 152.900 236.400 153.300 236.500 ;
        RECT 151.800 235.800 153.000 236.100 ;
        RECT 148.600 234.800 149.000 235.600 ;
        RECT 149.400 235.300 151.500 235.600 ;
        RECT 147.800 234.100 148.200 234.200 ;
        RECT 146.200 233.800 148.200 234.100 ;
        RECT 146.200 233.200 146.500 233.800 ;
        RECT 139.000 232.800 139.900 233.100 ;
        RECT 139.500 231.100 139.900 232.800 ;
        RECT 140.600 231.100 141.000 233.100 ;
        RECT 141.400 233.000 143.400 233.100 ;
        RECT 141.400 231.100 141.800 233.000 ;
        RECT 143.000 231.100 143.400 233.000 ;
        RECT 145.400 231.100 145.800 233.100 ;
        RECT 146.200 232.800 146.600 233.200 ;
        RECT 146.100 232.400 146.500 232.800 ;
        RECT 147.000 232.400 147.400 233.200 ;
        RECT 147.900 232.100 148.200 233.800 ;
        RECT 147.800 231.100 148.200 232.100 ;
        RECT 149.400 233.600 149.800 235.300 ;
        RECT 151.100 235.200 151.500 235.300 ;
        RECT 152.700 235.200 153.000 235.800 ;
        RECT 153.700 235.900 154.000 236.500 ;
        RECT 154.300 236.500 154.700 236.600 ;
        RECT 156.600 236.500 157.000 236.600 ;
        RECT 154.300 236.200 157.000 236.500 ;
        RECT 153.700 235.700 156.100 235.900 ;
        RECT 158.200 235.700 158.600 239.900 ;
        RECT 160.600 235.800 161.000 236.600 ;
        RECT 161.400 236.100 161.800 239.900 ;
        RECT 163.400 236.800 163.800 237.200 ;
        RECT 163.400 236.200 163.700 236.800 ;
        RECT 164.100 236.200 164.500 239.900 ;
        RECT 163.000 236.100 163.700 236.200 ;
        RECT 161.400 235.900 163.700 236.100 ;
        RECT 164.000 235.900 164.500 236.200 ;
        RECT 161.400 235.800 163.400 235.900 ;
        RECT 153.700 235.600 158.600 235.700 ;
        RECT 155.700 235.500 158.600 235.600 ;
        RECT 155.800 235.400 158.600 235.500 ;
        RECT 150.300 234.900 150.700 235.000 ;
        RECT 150.300 234.600 152.200 234.900 ;
        RECT 152.600 234.800 153.000 235.200 ;
        RECT 153.400 235.100 153.800 235.200 ;
        RECT 155.000 235.100 155.400 235.200 ;
        RECT 153.400 234.800 157.500 235.100 ;
        RECT 151.800 234.500 152.200 234.600 ;
        RECT 152.700 234.200 153.000 234.800 ;
        RECT 157.100 234.700 157.500 234.800 ;
        RECT 156.300 234.200 156.700 234.300 ;
        RECT 152.700 233.900 158.200 234.200 ;
        RECT 152.900 233.800 153.300 233.900 ;
        RECT 149.400 233.300 151.300 233.600 ;
        RECT 149.400 231.100 149.800 233.300 ;
        RECT 150.900 233.200 151.300 233.300 ;
        RECT 155.800 232.800 156.100 233.900 ;
        RECT 157.400 233.800 158.200 233.900 ;
        RECT 154.900 232.700 155.300 232.800 ;
        RECT 151.800 232.100 152.200 232.500 ;
        RECT 153.900 232.400 155.300 232.700 ;
        RECT 155.800 232.400 156.200 232.800 ;
        RECT 153.900 232.100 154.200 232.400 ;
        RECT 156.600 232.100 157.000 232.500 ;
        RECT 151.500 231.800 152.200 232.100 ;
        RECT 151.500 231.100 152.100 231.800 ;
        RECT 153.800 231.100 154.200 232.100 ;
        RECT 156.000 231.800 157.000 232.100 ;
        RECT 156.000 231.100 156.400 231.800 ;
        RECT 158.200 231.100 158.600 233.500 ;
        RECT 161.400 233.100 161.800 235.800 ;
        RECT 164.000 235.200 164.300 235.900 ;
        RECT 166.200 235.700 166.600 239.900 ;
        RECT 168.400 238.200 168.800 239.900 ;
        RECT 167.800 237.900 168.800 238.200 ;
        RECT 170.600 237.900 171.000 239.900 ;
        RECT 172.700 237.900 173.300 239.900 ;
        RECT 167.800 237.500 168.200 237.900 ;
        RECT 170.600 237.600 170.900 237.900 ;
        RECT 169.500 237.300 171.300 237.600 ;
        RECT 172.600 237.500 173.000 237.900 ;
        RECT 169.500 237.200 169.900 237.300 ;
        RECT 170.900 237.200 171.300 237.300 ;
        RECT 167.800 236.500 168.200 236.600 ;
        RECT 170.100 236.500 170.500 236.600 ;
        RECT 167.800 236.200 170.500 236.500 ;
        RECT 170.800 236.500 171.900 236.800 ;
        RECT 170.800 235.900 171.100 236.500 ;
        RECT 171.500 236.400 171.900 236.500 ;
        RECT 172.700 236.600 173.400 237.000 ;
        RECT 172.700 236.100 173.000 236.600 ;
        RECT 168.700 235.700 171.100 235.900 ;
        RECT 166.200 235.600 171.100 235.700 ;
        RECT 171.800 235.800 173.000 236.100 ;
        RECT 166.200 235.500 169.100 235.600 ;
        RECT 166.200 235.400 169.000 235.500 ;
        RECT 163.800 234.800 164.300 235.200 ;
        RECT 164.000 234.200 164.300 234.800 ;
        RECT 164.600 234.400 165.000 235.200 ;
        RECT 169.400 235.100 169.800 235.200 ;
        RECT 167.300 234.800 169.800 235.100 ;
        RECT 167.300 234.700 167.700 234.800 ;
        RECT 168.600 234.700 169.000 234.800 ;
        RECT 168.100 234.200 168.500 234.300 ;
        RECT 171.800 234.200 172.100 235.800 ;
        RECT 175.000 235.600 175.400 239.900 ;
        RECT 173.300 235.300 175.400 235.600 ;
        RECT 175.800 237.500 176.200 239.500 ;
        RECT 175.800 235.800 176.100 237.500 ;
        RECT 177.900 236.400 178.300 239.900 ;
        RECT 177.900 236.100 178.700 236.400 ;
        RECT 175.800 235.500 177.700 235.800 ;
        RECT 173.300 235.200 173.700 235.300 ;
        RECT 174.100 234.900 174.500 235.000 ;
        RECT 172.600 234.600 174.500 234.900 ;
        RECT 172.600 234.500 173.000 234.600 ;
        RECT 162.200 233.400 162.600 234.200 ;
        RECT 163.000 233.800 164.300 234.200 ;
        RECT 165.400 234.100 165.800 234.200 ;
        RECT 165.000 233.800 165.800 234.100 ;
        RECT 166.600 233.900 172.100 234.200 ;
        RECT 166.600 233.800 167.400 233.900 ;
        RECT 163.100 233.100 163.400 233.800 ;
        RECT 165.000 233.600 165.400 233.800 ;
        RECT 163.900 233.100 165.700 233.300 ;
        RECT 160.900 232.800 161.800 233.100 ;
        RECT 160.900 231.100 161.300 232.800 ;
        RECT 163.000 231.100 163.400 233.100 ;
        RECT 163.800 233.000 165.800 233.100 ;
        RECT 163.800 231.100 164.200 233.000 ;
        RECT 165.400 231.100 165.800 233.000 ;
        RECT 166.200 231.100 166.600 233.500 ;
        RECT 168.700 233.200 169.000 233.900 ;
        RECT 171.500 233.800 171.900 233.900 ;
        RECT 175.000 233.600 175.400 235.300 ;
        RECT 175.800 234.400 176.200 235.200 ;
        RECT 176.600 234.400 177.000 235.200 ;
        RECT 177.400 234.500 177.700 235.500 ;
        RECT 177.400 234.100 178.100 234.500 ;
        RECT 178.400 234.200 178.700 236.100 ;
        RECT 179.000 235.100 179.400 235.600 ;
        RECT 181.400 235.100 181.800 239.900 ;
        RECT 183.400 236.800 183.800 237.200 ;
        RECT 182.200 235.800 182.600 236.600 ;
        RECT 183.400 236.200 183.700 236.800 ;
        RECT 184.100 236.200 184.500 239.900 ;
        RECT 183.000 235.900 183.700 236.200 ;
        RECT 183.000 235.800 183.400 235.900 ;
        RECT 184.000 235.800 185.000 236.200 ;
        RECT 183.000 235.100 183.300 235.800 ;
        RECT 179.000 234.800 180.100 235.100 ;
        RECT 177.400 233.900 177.900 234.100 ;
        RECT 173.500 233.300 175.400 233.600 ;
        RECT 173.500 233.200 173.900 233.300 ;
        RECT 167.800 232.100 168.200 232.500 ;
        RECT 168.600 232.400 169.000 233.200 ;
        RECT 169.500 232.700 169.900 232.800 ;
        RECT 169.500 232.400 170.900 232.700 ;
        RECT 170.600 232.100 170.900 232.400 ;
        RECT 172.600 232.100 173.000 232.500 ;
        RECT 167.800 231.800 168.800 232.100 ;
        RECT 168.400 231.100 168.800 231.800 ;
        RECT 170.600 231.100 171.000 232.100 ;
        RECT 172.600 231.800 173.300 232.100 ;
        RECT 172.700 231.100 173.300 231.800 ;
        RECT 175.000 231.100 175.400 233.300 ;
        RECT 175.800 233.600 177.900 233.900 ;
        RECT 178.400 233.800 179.400 234.200 ;
        RECT 179.800 234.100 180.100 234.800 ;
        RECT 181.400 234.800 183.300 235.100 ;
        RECT 180.600 234.100 181.000 234.200 ;
        RECT 179.800 233.800 181.000 234.100 ;
        RECT 175.800 232.500 176.100 233.600 ;
        RECT 178.400 233.500 178.700 233.800 ;
        RECT 178.300 233.300 178.700 233.500 ;
        RECT 180.600 233.400 181.000 233.800 ;
        RECT 177.900 233.000 178.700 233.300 ;
        RECT 181.400 233.100 181.800 234.800 ;
        RECT 184.000 234.200 184.300 235.800 ;
        RECT 186.200 235.700 186.600 239.900 ;
        RECT 188.400 238.200 188.800 239.900 ;
        RECT 187.800 237.900 188.800 238.200 ;
        RECT 190.600 237.900 191.000 239.900 ;
        RECT 192.700 237.900 193.300 239.900 ;
        RECT 187.800 237.500 188.200 237.900 ;
        RECT 190.600 237.600 190.900 237.900 ;
        RECT 189.500 237.300 191.300 237.600 ;
        RECT 192.600 237.500 193.000 237.900 ;
        RECT 189.500 237.200 189.900 237.300 ;
        RECT 190.900 237.200 191.300 237.300 ;
        RECT 187.800 236.500 188.200 236.600 ;
        RECT 190.100 236.500 190.500 236.600 ;
        RECT 187.800 236.200 190.500 236.500 ;
        RECT 190.800 236.500 191.900 236.800 ;
        RECT 190.800 235.900 191.100 236.500 ;
        RECT 191.500 236.400 191.900 236.500 ;
        RECT 192.700 236.600 193.400 237.000 ;
        RECT 192.700 236.100 193.000 236.600 ;
        RECT 188.700 235.700 191.100 235.900 ;
        RECT 186.200 235.600 191.100 235.700 ;
        RECT 191.800 235.800 193.000 236.100 ;
        RECT 186.200 235.500 189.100 235.600 ;
        RECT 186.200 235.400 189.000 235.500 ;
        RECT 184.600 234.400 185.000 235.200 ;
        RECT 189.400 235.100 189.800 235.200 ;
        RECT 187.300 234.800 189.800 235.100 ;
        RECT 187.300 234.700 187.700 234.800 ;
        RECT 188.600 234.700 189.000 234.800 ;
        RECT 188.100 234.200 188.500 234.300 ;
        RECT 191.800 234.200 192.100 235.800 ;
        RECT 195.000 235.600 195.400 239.900 ;
        RECT 193.300 235.300 195.400 235.600 ;
        RECT 193.300 235.200 193.700 235.300 ;
        RECT 194.100 234.900 194.500 235.000 ;
        RECT 192.600 234.600 194.500 234.900 ;
        RECT 192.600 234.500 193.000 234.600 ;
        RECT 183.000 233.800 184.300 234.200 ;
        RECT 185.400 234.100 185.800 234.200 ;
        RECT 185.000 233.800 185.800 234.100 ;
        RECT 186.600 233.900 192.100 234.200 ;
        RECT 186.600 233.800 187.400 233.900 ;
        RECT 183.100 233.100 183.400 233.800 ;
        RECT 185.000 233.600 185.400 233.800 ;
        RECT 183.900 233.100 185.700 233.300 ;
        RECT 175.800 231.500 176.200 232.500 ;
        RECT 177.900 232.200 178.300 233.000 ;
        RECT 181.400 232.800 182.300 233.100 ;
        RECT 177.400 231.800 178.300 232.200 ;
        RECT 177.900 231.500 178.300 231.800 ;
        RECT 181.900 231.100 182.300 232.800 ;
        RECT 183.000 231.100 183.400 233.100 ;
        RECT 183.800 233.000 185.800 233.100 ;
        RECT 183.800 231.100 184.200 233.000 ;
        RECT 185.400 231.100 185.800 233.000 ;
        RECT 186.200 231.100 186.600 233.500 ;
        RECT 188.700 232.800 189.000 233.900 ;
        RECT 191.500 233.800 191.900 233.900 ;
        RECT 195.000 233.600 195.400 235.300 ;
        RECT 193.500 233.300 195.400 233.600 ;
        RECT 193.500 233.200 193.900 233.300 ;
        RECT 187.800 232.100 188.200 232.500 ;
        RECT 188.600 232.400 189.000 232.800 ;
        RECT 189.500 232.700 189.900 232.800 ;
        RECT 189.500 232.400 190.900 232.700 ;
        RECT 190.600 232.100 190.900 232.400 ;
        RECT 192.600 232.100 193.000 232.500 ;
        RECT 187.800 231.800 188.800 232.100 ;
        RECT 188.400 231.100 188.800 231.800 ;
        RECT 190.600 231.100 191.000 232.100 ;
        RECT 192.600 231.800 193.300 232.100 ;
        RECT 192.700 231.100 193.300 231.800 ;
        RECT 195.000 231.100 195.400 233.300 ;
        RECT 195.800 235.600 196.200 239.900 ;
        RECT 197.900 237.900 198.500 239.900 ;
        RECT 200.200 237.900 200.600 239.900 ;
        RECT 202.400 238.200 202.800 239.900 ;
        RECT 202.400 237.900 203.400 238.200 ;
        RECT 198.200 237.500 198.600 237.900 ;
        RECT 200.300 237.600 200.600 237.900 ;
        RECT 199.900 237.300 201.700 237.600 ;
        RECT 203.000 237.500 203.400 237.900 ;
        RECT 199.900 237.200 200.300 237.300 ;
        RECT 201.300 237.200 201.700 237.300 ;
        RECT 197.800 236.600 198.500 237.000 ;
        RECT 198.200 236.100 198.500 236.600 ;
        RECT 199.300 236.500 200.400 236.800 ;
        RECT 199.300 236.400 199.700 236.500 ;
        RECT 198.200 235.800 199.400 236.100 ;
        RECT 195.800 235.300 197.900 235.600 ;
        RECT 195.800 233.600 196.200 235.300 ;
        RECT 197.500 235.200 197.900 235.300 ;
        RECT 196.700 234.900 197.100 235.000 ;
        RECT 196.700 234.600 198.600 234.900 ;
        RECT 198.200 234.500 198.600 234.600 ;
        RECT 199.100 234.200 199.400 235.800 ;
        RECT 200.100 235.900 200.400 236.500 ;
        RECT 200.700 236.500 201.100 236.600 ;
        RECT 203.000 236.500 203.400 236.600 ;
        RECT 200.700 236.200 203.400 236.500 ;
        RECT 200.100 235.700 202.500 235.900 ;
        RECT 204.600 235.700 205.000 239.900 ;
        RECT 200.100 235.600 205.000 235.700 ;
        RECT 207.800 235.600 208.200 239.900 ;
        RECT 209.400 235.600 209.800 239.900 ;
        RECT 211.000 235.600 211.400 239.900 ;
        RECT 212.600 235.600 213.000 239.900 ;
        RECT 215.000 235.600 215.400 239.900 ;
        RECT 216.600 235.600 217.000 239.900 ;
        RECT 218.200 235.600 218.600 239.900 ;
        RECT 219.800 235.600 220.200 239.900 ;
        RECT 222.700 236.200 223.100 239.900 ;
        RECT 223.400 236.800 223.800 237.200 ;
        RECT 223.500 236.200 223.800 236.800 ;
        RECT 222.700 235.900 223.200 236.200 ;
        RECT 223.500 235.900 224.200 236.200 ;
        RECT 202.100 235.500 205.000 235.600 ;
        RECT 202.200 235.400 205.000 235.500 ;
        RECT 207.000 235.200 208.200 235.600 ;
        RECT 208.700 235.200 209.800 235.600 ;
        RECT 210.300 235.200 211.400 235.600 ;
        RECT 212.100 235.200 213.000 235.600 ;
        RECT 214.200 235.200 215.400 235.600 ;
        RECT 215.900 235.200 217.000 235.600 ;
        RECT 217.500 235.200 218.600 235.600 ;
        RECT 219.300 235.200 220.200 235.600 ;
        RECT 199.800 235.100 200.200 235.200 ;
        RECT 201.400 235.100 201.800 235.200 ;
        RECT 206.200 235.100 206.600 235.200 ;
        RECT 207.000 235.100 207.400 235.200 ;
        RECT 199.800 234.800 203.900 235.100 ;
        RECT 206.200 234.800 207.400 235.100 ;
        RECT 203.500 234.700 203.900 234.800 ;
        RECT 202.700 234.200 203.100 234.300 ;
        RECT 199.100 233.900 204.600 234.200 ;
        RECT 199.300 233.800 199.700 233.900 ;
        RECT 195.800 233.300 197.700 233.600 ;
        RECT 195.800 231.100 196.200 233.300 ;
        RECT 197.300 233.200 197.700 233.300 ;
        RECT 202.200 232.800 202.500 233.900 ;
        RECT 203.800 233.800 204.600 233.900 ;
        RECT 207.000 233.800 207.400 234.800 ;
        RECT 208.700 234.500 209.100 235.200 ;
        RECT 210.300 234.500 210.700 235.200 ;
        RECT 212.100 234.500 212.500 235.200 ;
        RECT 207.800 234.100 209.100 234.500 ;
        RECT 209.500 234.100 210.700 234.500 ;
        RECT 211.200 234.100 212.500 234.500 ;
        RECT 212.900 234.100 213.800 234.500 ;
        RECT 208.700 233.800 209.100 234.100 ;
        RECT 210.300 233.800 210.700 234.100 ;
        RECT 212.100 233.800 212.500 234.100 ;
        RECT 213.400 233.800 213.800 234.100 ;
        RECT 214.200 233.800 214.600 235.200 ;
        RECT 215.900 234.500 216.300 235.200 ;
        RECT 217.500 234.500 217.900 235.200 ;
        RECT 219.300 234.500 219.700 235.200 ;
        RECT 215.000 234.100 216.300 234.500 ;
        RECT 216.700 234.100 217.900 234.500 ;
        RECT 218.400 234.100 219.700 234.500 ;
        RECT 220.100 234.100 221.000 234.500 ;
        RECT 222.200 234.400 222.600 235.200 ;
        RECT 222.900 234.200 223.200 235.900 ;
        RECT 223.800 235.800 224.200 235.900 ;
        RECT 224.600 235.800 225.000 236.600 ;
        RECT 223.800 235.100 224.100 235.800 ;
        RECT 225.400 235.100 225.800 239.900 ;
        RECT 227.800 235.600 228.200 239.900 ;
        RECT 229.400 235.600 229.800 239.900 ;
        RECT 231.000 235.600 231.400 239.900 ;
        RECT 232.600 235.600 233.000 239.900 ;
        RECT 223.800 234.800 225.800 235.100 ;
        RECT 215.900 233.800 216.300 234.100 ;
        RECT 217.500 233.800 217.900 234.100 ;
        RECT 219.300 233.800 219.700 234.100 ;
        RECT 220.600 233.800 221.000 234.100 ;
        RECT 221.400 234.100 221.800 234.200 ;
        RECT 221.400 233.800 222.200 234.100 ;
        RECT 222.900 233.800 224.200 234.200 ;
        RECT 201.300 232.700 201.700 232.800 ;
        RECT 198.200 232.100 198.600 232.500 ;
        RECT 200.300 232.400 201.700 232.700 ;
        RECT 202.200 232.400 202.600 232.800 ;
        RECT 200.300 232.100 200.600 232.400 ;
        RECT 203.000 232.100 203.400 232.500 ;
        RECT 197.900 231.800 198.600 232.100 ;
        RECT 197.900 231.100 198.500 231.800 ;
        RECT 200.200 231.100 200.600 232.100 ;
        RECT 202.400 231.800 203.400 232.100 ;
        RECT 202.400 231.100 202.800 231.800 ;
        RECT 204.600 231.100 205.000 233.500 ;
        RECT 207.000 233.400 208.200 233.800 ;
        RECT 208.700 233.400 209.800 233.800 ;
        RECT 210.300 233.400 211.400 233.800 ;
        RECT 212.100 233.400 213.000 233.800 ;
        RECT 214.200 233.400 215.400 233.800 ;
        RECT 215.900 233.400 217.000 233.800 ;
        RECT 217.500 233.400 218.600 233.800 ;
        RECT 219.300 233.400 220.200 233.800 ;
        RECT 221.800 233.600 222.200 233.800 ;
        RECT 207.800 231.100 208.200 233.400 ;
        RECT 209.400 231.100 209.800 233.400 ;
        RECT 211.000 231.100 211.400 233.400 ;
        RECT 212.600 231.100 213.000 233.400 ;
        RECT 215.000 231.100 215.400 233.400 ;
        RECT 216.600 231.100 217.000 233.400 ;
        RECT 218.200 231.100 218.600 233.400 ;
        RECT 219.800 231.100 220.200 233.400 ;
        RECT 221.500 233.100 223.300 233.300 ;
        RECT 223.800 233.100 224.100 233.800 ;
        RECT 225.400 233.100 225.800 234.800 ;
        RECT 227.000 235.200 228.200 235.600 ;
        RECT 228.700 235.200 229.800 235.600 ;
        RECT 230.300 235.200 231.400 235.600 ;
        RECT 232.100 235.200 233.000 235.600 ;
        RECT 234.200 235.700 234.600 239.900 ;
        RECT 236.400 238.200 236.800 239.900 ;
        RECT 235.800 237.900 236.800 238.200 ;
        RECT 238.600 237.900 239.000 239.900 ;
        RECT 240.700 237.900 241.300 239.900 ;
        RECT 235.800 237.500 236.200 237.900 ;
        RECT 238.600 237.600 238.900 237.900 ;
        RECT 237.500 237.300 239.300 237.600 ;
        RECT 240.600 237.500 241.000 237.900 ;
        RECT 237.500 237.200 237.900 237.300 ;
        RECT 238.900 237.200 239.300 237.300 ;
        RECT 235.800 236.500 236.200 236.600 ;
        RECT 238.100 236.500 238.500 236.600 ;
        RECT 235.800 236.200 238.500 236.500 ;
        RECT 238.800 236.500 239.900 236.800 ;
        RECT 238.800 235.900 239.100 236.500 ;
        RECT 239.500 236.400 239.900 236.500 ;
        RECT 240.700 236.600 241.400 237.000 ;
        RECT 240.700 236.100 241.000 236.600 ;
        RECT 236.700 235.700 239.100 235.900 ;
        RECT 234.200 235.600 239.100 235.700 ;
        RECT 239.800 235.800 241.000 236.100 ;
        RECT 234.200 235.500 237.100 235.600 ;
        RECT 234.200 235.400 237.000 235.500 ;
        RECT 226.200 233.400 226.600 234.200 ;
        RECT 227.000 233.800 227.400 235.200 ;
        RECT 228.700 234.500 229.100 235.200 ;
        RECT 230.300 234.500 230.700 235.200 ;
        RECT 232.100 234.500 232.500 235.200 ;
        RECT 237.400 235.100 237.800 235.200 ;
        RECT 238.200 235.100 238.600 235.200 ;
        RECT 235.300 234.800 238.600 235.100 ;
        RECT 235.300 234.700 235.700 234.800 ;
        RECT 227.800 234.100 229.100 234.500 ;
        RECT 229.500 234.100 230.700 234.500 ;
        RECT 231.200 234.100 232.500 234.500 ;
        RECT 236.100 234.200 236.500 234.300 ;
        RECT 239.800 234.200 240.100 235.800 ;
        RECT 243.000 235.600 243.400 239.900 ;
        RECT 241.300 235.300 243.400 235.600 ;
        RECT 241.300 235.200 241.700 235.300 ;
        RECT 242.100 234.900 242.500 235.000 ;
        RECT 240.600 234.600 242.500 234.900 ;
        RECT 240.600 234.500 241.000 234.600 ;
        RECT 228.700 233.800 229.100 234.100 ;
        RECT 230.300 233.800 230.700 234.100 ;
        RECT 232.100 233.800 232.500 234.100 ;
        RECT 234.600 233.900 240.100 234.200 ;
        RECT 234.600 233.800 235.400 233.900 ;
        RECT 227.000 233.400 228.200 233.800 ;
        RECT 228.700 233.400 229.800 233.800 ;
        RECT 230.300 233.400 231.400 233.800 ;
        RECT 232.100 233.400 233.000 233.800 ;
        RECT 221.400 233.000 223.400 233.100 ;
        RECT 221.400 231.100 221.800 233.000 ;
        RECT 223.000 231.100 223.400 233.000 ;
        RECT 223.800 231.100 224.200 233.100 ;
        RECT 224.900 232.800 225.800 233.100 ;
        RECT 224.900 231.100 225.300 232.800 ;
        RECT 227.800 231.100 228.200 233.400 ;
        RECT 229.400 231.100 229.800 233.400 ;
        RECT 231.000 231.100 231.400 233.400 ;
        RECT 232.600 231.100 233.000 233.400 ;
        RECT 234.200 231.100 234.600 233.500 ;
        RECT 236.700 232.800 237.000 233.900 ;
        RECT 237.400 233.800 237.800 233.900 ;
        RECT 239.500 233.800 239.900 233.900 ;
        RECT 243.000 233.600 243.400 235.300 ;
        RECT 241.500 233.300 243.400 233.600 ;
        RECT 241.500 233.200 241.900 233.300 ;
        RECT 235.800 232.100 236.200 232.500 ;
        RECT 236.600 232.400 237.000 232.800 ;
        RECT 237.500 232.700 237.900 232.800 ;
        RECT 237.500 232.400 238.900 232.700 ;
        RECT 238.600 232.100 238.900 232.400 ;
        RECT 240.600 232.100 241.000 232.500 ;
        RECT 235.800 231.800 236.800 232.100 ;
        RECT 236.400 231.100 236.800 231.800 ;
        RECT 238.600 231.100 239.000 232.100 ;
        RECT 240.600 231.800 241.300 232.100 ;
        RECT 240.700 231.100 241.300 231.800 ;
        RECT 243.000 231.100 243.400 233.300 ;
        RECT 243.800 235.600 244.200 239.900 ;
        RECT 245.900 237.900 246.500 239.900 ;
        RECT 248.200 237.900 248.600 239.900 ;
        RECT 250.400 238.200 250.800 239.900 ;
        RECT 250.400 237.900 251.400 238.200 ;
        RECT 246.200 237.500 246.600 237.900 ;
        RECT 248.300 237.600 248.600 237.900 ;
        RECT 247.900 237.300 249.700 237.600 ;
        RECT 251.000 237.500 251.400 237.900 ;
        RECT 247.900 237.200 248.300 237.300 ;
        RECT 249.300 237.200 249.700 237.300 ;
        RECT 245.800 236.600 246.500 237.000 ;
        RECT 246.200 236.100 246.500 236.600 ;
        RECT 247.300 236.500 248.400 236.800 ;
        RECT 247.300 236.400 247.700 236.500 ;
        RECT 246.200 235.800 247.400 236.100 ;
        RECT 243.800 235.300 245.900 235.600 ;
        RECT 243.800 233.600 244.200 235.300 ;
        RECT 245.500 235.200 245.900 235.300 ;
        RECT 244.700 234.900 245.100 235.000 ;
        RECT 244.700 234.600 246.600 234.900 ;
        RECT 246.200 234.500 246.600 234.600 ;
        RECT 247.100 234.200 247.400 235.800 ;
        RECT 248.100 235.900 248.400 236.500 ;
        RECT 248.700 236.500 249.100 236.600 ;
        RECT 251.000 236.500 251.400 236.600 ;
        RECT 248.700 236.200 251.400 236.500 ;
        RECT 248.100 235.700 250.500 235.900 ;
        RECT 252.600 235.700 253.000 239.900 ;
        RECT 253.400 235.800 253.800 236.600 ;
        RECT 248.100 235.600 253.000 235.700 ;
        RECT 250.100 235.500 253.000 235.600 ;
        RECT 250.200 235.400 253.000 235.500 ;
        RECT 248.600 235.100 249.000 235.200 ;
        RECT 249.400 235.100 249.800 235.200 ;
        RECT 248.600 234.800 251.900 235.100 ;
        RECT 251.500 234.700 251.900 234.800 ;
        RECT 250.700 234.200 251.100 234.300 ;
        RECT 247.100 233.900 252.600 234.200 ;
        RECT 247.300 233.800 247.700 233.900 ;
        RECT 243.800 233.300 245.700 233.600 ;
        RECT 243.800 231.100 244.200 233.300 ;
        RECT 245.300 233.200 245.700 233.300 ;
        RECT 250.200 233.200 250.500 233.900 ;
        RECT 251.800 233.800 252.600 233.900 ;
        RECT 249.300 232.700 249.700 232.800 ;
        RECT 246.200 232.100 246.600 232.500 ;
        RECT 248.300 232.400 249.700 232.700 ;
        RECT 250.200 232.400 250.600 233.200 ;
        RECT 248.300 232.100 248.600 232.400 ;
        RECT 251.000 232.100 251.400 232.500 ;
        RECT 245.900 231.800 246.600 232.100 ;
        RECT 245.900 231.100 246.500 231.800 ;
        RECT 248.200 231.100 248.600 232.100 ;
        RECT 250.400 231.800 251.400 232.100 ;
        RECT 250.400 231.100 250.800 231.800 ;
        RECT 252.600 231.100 253.000 233.500 ;
        RECT 254.200 233.100 254.600 239.900 ;
        RECT 256.600 235.600 257.000 239.900 ;
        RECT 258.200 235.600 258.600 239.900 ;
        RECT 259.800 235.600 260.200 239.900 ;
        RECT 261.400 235.600 261.800 239.900 ;
        RECT 256.600 235.200 257.500 235.600 ;
        RECT 258.200 235.200 259.300 235.600 ;
        RECT 259.800 235.200 260.900 235.600 ;
        RECT 261.400 235.200 262.600 235.600 ;
        RECT 257.100 234.500 257.500 235.200 ;
        RECT 258.900 234.500 259.300 235.200 ;
        RECT 260.500 234.500 260.900 235.200 ;
        RECT 255.000 233.400 255.400 234.200 ;
        RECT 257.100 234.100 258.400 234.500 ;
        RECT 258.900 234.100 260.100 234.500 ;
        RECT 260.500 234.100 261.800 234.500 ;
        RECT 257.100 233.800 257.500 234.100 ;
        RECT 258.900 233.800 259.300 234.100 ;
        RECT 260.500 233.800 260.900 234.100 ;
        RECT 262.200 233.800 262.600 235.200 ;
        RECT 256.600 233.400 257.500 233.800 ;
        RECT 258.200 233.400 259.300 233.800 ;
        RECT 259.800 233.400 260.900 233.800 ;
        RECT 261.400 233.400 262.600 233.800 ;
        RECT 253.700 232.800 254.600 233.100 ;
        RECT 253.700 232.200 254.100 232.800 ;
        RECT 253.400 231.800 254.100 232.200 ;
        RECT 253.700 231.100 254.100 231.800 ;
        RECT 256.600 231.100 257.000 233.400 ;
        RECT 258.200 231.100 258.600 233.400 ;
        RECT 259.800 231.100 260.200 233.400 ;
        RECT 261.400 231.100 261.800 233.400 ;
        RECT 1.400 227.600 1.800 229.900 ;
        RECT 3.000 227.600 3.400 229.900 ;
        RECT 4.600 227.600 5.000 229.900 ;
        RECT 6.200 227.600 6.600 229.900 ;
        RECT 1.400 227.200 2.300 227.600 ;
        RECT 3.000 227.200 4.100 227.600 ;
        RECT 4.600 227.200 5.700 227.600 ;
        RECT 6.200 227.200 7.400 227.600 ;
        RECT 7.800 227.500 8.200 229.900 ;
        RECT 10.000 229.200 10.400 229.900 ;
        RECT 9.400 228.900 10.400 229.200 ;
        RECT 12.200 228.900 12.600 229.900 ;
        RECT 14.300 229.200 14.900 229.900 ;
        RECT 14.200 228.900 14.900 229.200 ;
        RECT 9.400 228.500 9.800 228.900 ;
        RECT 12.200 228.600 12.500 228.900 ;
        RECT 10.200 228.200 10.600 228.600 ;
        RECT 11.100 228.300 12.500 228.600 ;
        RECT 14.200 228.500 14.600 228.900 ;
        RECT 11.100 228.200 11.500 228.300 ;
        RECT 0.600 226.900 1.000 227.200 ;
        RECT 1.900 226.900 2.300 227.200 ;
        RECT 3.700 226.900 4.100 227.200 ;
        RECT 5.300 226.900 5.700 227.200 ;
        RECT 0.600 226.500 1.500 226.900 ;
        RECT 1.900 226.500 3.200 226.900 ;
        RECT 3.700 226.500 4.900 226.900 ;
        RECT 5.300 226.500 6.600 226.900 ;
        RECT 1.900 225.800 2.300 226.500 ;
        RECT 3.700 225.800 4.100 226.500 ;
        RECT 5.300 225.800 5.700 226.500 ;
        RECT 7.000 225.800 7.400 227.200 ;
        RECT 8.200 227.100 9.000 227.200 ;
        RECT 10.300 227.100 10.600 228.200 ;
        RECT 15.100 227.700 15.500 227.800 ;
        RECT 16.600 227.700 17.000 229.900 ;
        RECT 15.100 227.400 17.000 227.700 ;
        RECT 13.100 227.100 13.500 227.200 ;
        RECT 8.200 226.800 13.700 227.100 ;
        RECT 9.700 226.700 10.100 226.800 ;
        RECT 8.900 226.200 9.300 226.300 ;
        RECT 8.900 226.100 11.400 226.200 ;
        RECT 12.600 226.100 13.000 226.200 ;
        RECT 8.900 225.900 13.000 226.100 ;
        RECT 11.000 225.800 13.000 225.900 ;
        RECT 1.400 225.400 2.300 225.800 ;
        RECT 3.000 225.400 4.100 225.800 ;
        RECT 4.600 225.400 5.700 225.800 ;
        RECT 6.200 225.400 7.400 225.800 ;
        RECT 7.800 225.500 10.600 225.600 ;
        RECT 7.800 225.400 10.700 225.500 ;
        RECT 1.400 221.100 1.800 225.400 ;
        RECT 3.000 221.100 3.400 225.400 ;
        RECT 4.600 221.100 5.000 225.400 ;
        RECT 6.200 221.100 6.600 225.400 ;
        RECT 7.800 225.300 12.700 225.400 ;
        RECT 7.800 221.100 8.200 225.300 ;
        RECT 10.300 225.100 12.700 225.300 ;
        RECT 9.400 224.500 12.100 224.800 ;
        RECT 9.400 224.400 9.800 224.500 ;
        RECT 11.700 224.400 12.100 224.500 ;
        RECT 12.400 224.500 12.700 225.100 ;
        RECT 13.400 225.200 13.700 226.800 ;
        RECT 14.200 226.400 14.600 226.500 ;
        RECT 14.200 226.100 16.100 226.400 ;
        RECT 15.700 226.000 16.100 226.100 ;
        RECT 14.900 225.700 15.300 225.800 ;
        RECT 16.600 225.700 17.000 227.400 ;
        RECT 19.000 227.900 19.400 229.900 ;
        RECT 21.400 228.900 21.800 229.900 ;
        RECT 19.700 228.200 20.100 228.600 ;
        RECT 19.800 228.100 20.200 228.200 ;
        RECT 21.400 228.100 21.700 228.900 ;
        RECT 19.000 227.200 19.300 227.900 ;
        RECT 19.800 227.800 21.700 228.100 ;
        RECT 22.200 227.800 22.600 228.600 ;
        RECT 21.400 227.200 21.700 227.800 ;
        RECT 23.000 227.500 23.400 229.900 ;
        RECT 25.200 229.200 25.600 229.900 ;
        RECT 24.600 228.900 25.600 229.200 ;
        RECT 27.400 228.900 27.800 229.900 ;
        RECT 29.500 229.200 30.100 229.900 ;
        RECT 29.400 228.900 30.100 229.200 ;
        RECT 24.600 228.500 25.000 228.900 ;
        RECT 27.400 228.600 27.700 228.900 ;
        RECT 25.400 227.800 25.800 228.600 ;
        RECT 26.300 228.300 27.700 228.600 ;
        RECT 29.400 228.500 29.800 228.900 ;
        RECT 26.300 228.200 26.700 228.300 ;
        RECT 18.200 226.400 18.600 227.200 ;
        RECT 19.000 226.800 19.400 227.200 ;
        RECT 21.400 226.800 21.800 227.200 ;
        RECT 23.400 227.100 24.200 227.200 ;
        RECT 25.500 227.100 25.800 227.800 ;
        RECT 30.300 227.700 30.700 227.800 ;
        RECT 31.800 227.700 32.200 229.900 ;
        RECT 30.300 227.400 32.200 227.700 ;
        RECT 28.300 227.100 28.700 227.200 ;
        RECT 23.400 226.800 28.900 227.100 ;
        RECT 17.400 226.100 17.800 226.200 ;
        RECT 19.000 226.100 19.300 226.800 ;
        RECT 19.800 226.100 20.200 226.200 ;
        RECT 17.400 225.800 18.200 226.100 ;
        RECT 19.000 225.800 20.200 226.100 ;
        RECT 14.900 225.400 17.000 225.700 ;
        RECT 17.800 225.600 18.200 225.800 ;
        RECT 13.400 224.900 14.600 225.200 ;
        RECT 13.100 224.500 13.500 224.600 ;
        RECT 12.400 224.200 13.500 224.500 ;
        RECT 14.300 224.400 14.600 224.900 ;
        RECT 14.300 224.000 15.000 224.400 ;
        RECT 11.100 223.700 11.500 223.800 ;
        RECT 12.500 223.700 12.900 223.800 ;
        RECT 9.400 223.100 9.800 223.500 ;
        RECT 11.100 223.400 12.900 223.700 ;
        RECT 12.200 223.100 12.500 223.400 ;
        RECT 14.200 223.100 14.600 223.500 ;
        RECT 9.400 222.800 10.400 223.100 ;
        RECT 10.000 221.100 10.400 222.800 ;
        RECT 12.200 221.100 12.600 223.100 ;
        RECT 14.300 221.100 14.900 223.100 ;
        RECT 16.600 221.100 17.000 225.400 ;
        RECT 19.800 225.100 20.100 225.800 ;
        RECT 20.600 225.400 21.000 226.200 ;
        RECT 21.400 225.100 21.700 226.800 ;
        RECT 24.900 226.700 25.300 226.800 ;
        RECT 24.100 226.200 24.500 226.300 ;
        RECT 24.100 225.900 26.600 226.200 ;
        RECT 26.200 225.800 26.600 225.900 ;
        RECT 23.000 225.500 25.800 225.600 ;
        RECT 23.000 225.400 25.900 225.500 ;
        RECT 23.000 225.300 27.900 225.400 ;
        RECT 17.400 224.800 19.400 225.100 ;
        RECT 17.400 221.100 17.800 224.800 ;
        RECT 19.000 221.100 19.400 224.800 ;
        RECT 19.800 221.100 20.200 225.100 ;
        RECT 20.900 224.700 21.800 225.100 ;
        RECT 20.900 221.100 21.300 224.700 ;
        RECT 23.000 221.100 23.400 225.300 ;
        RECT 25.500 225.100 27.900 225.300 ;
        RECT 24.600 224.500 27.300 224.800 ;
        RECT 24.600 224.400 25.000 224.500 ;
        RECT 26.900 224.400 27.300 224.500 ;
        RECT 27.600 224.500 27.900 225.100 ;
        RECT 28.600 225.200 28.900 226.800 ;
        RECT 29.400 226.400 29.800 226.500 ;
        RECT 29.400 226.100 31.300 226.400 ;
        RECT 30.900 226.000 31.300 226.100 ;
        RECT 30.100 225.700 30.500 225.800 ;
        RECT 31.800 225.700 32.200 227.400 ;
        RECT 32.600 228.500 33.000 229.500 ;
        RECT 32.600 227.400 32.900 228.500 ;
        RECT 34.700 228.000 35.100 229.500 ;
        RECT 34.700 227.700 35.500 228.000 ;
        RECT 35.100 227.500 35.500 227.700 ;
        RECT 32.600 227.100 34.700 227.400 ;
        RECT 34.200 226.900 34.700 227.100 ;
        RECT 35.200 227.200 35.500 227.500 ;
        RECT 32.600 225.800 33.000 226.600 ;
        RECT 33.400 225.800 33.800 226.600 ;
        RECT 34.200 226.500 34.900 226.900 ;
        RECT 35.200 226.800 36.200 227.200 ;
        RECT 30.100 225.400 32.200 225.700 ;
        RECT 34.200 225.500 34.500 226.500 ;
        RECT 28.600 224.900 29.800 225.200 ;
        RECT 28.300 224.500 28.700 224.600 ;
        RECT 27.600 224.200 28.700 224.500 ;
        RECT 29.500 224.400 29.800 224.900 ;
        RECT 29.500 224.200 30.200 224.400 ;
        RECT 29.500 224.000 30.600 224.200 ;
        RECT 29.900 223.800 30.600 224.000 ;
        RECT 26.300 223.700 26.700 223.800 ;
        RECT 27.700 223.700 28.100 223.800 ;
        RECT 24.600 223.100 25.000 223.500 ;
        RECT 26.300 223.400 28.100 223.700 ;
        RECT 27.400 223.100 27.700 223.400 ;
        RECT 29.400 223.100 29.800 223.500 ;
        RECT 24.600 222.800 25.600 223.100 ;
        RECT 25.200 221.100 25.600 222.800 ;
        RECT 27.400 221.100 27.800 223.100 ;
        RECT 29.500 221.100 30.100 223.100 ;
        RECT 31.800 221.100 32.200 225.400 ;
        RECT 32.600 225.200 34.500 225.500 ;
        RECT 32.600 223.500 32.900 225.200 ;
        RECT 35.200 224.900 35.500 226.800 ;
        RECT 35.800 226.100 36.200 226.200 ;
        RECT 37.400 226.100 37.800 229.900 ;
        RECT 38.200 227.800 38.600 228.600 ;
        RECT 39.000 228.500 39.400 229.500 ;
        RECT 39.000 227.400 39.300 228.500 ;
        RECT 41.100 228.000 41.500 229.500 ;
        RECT 44.600 228.200 45.000 229.900 ;
        RECT 41.100 227.700 41.900 228.000 ;
        RECT 41.500 227.500 41.900 227.700 ;
        RECT 39.000 227.100 41.100 227.400 ;
        RECT 40.600 226.900 41.100 227.100 ;
        RECT 41.600 227.200 41.900 227.500 ;
        RECT 44.500 227.900 45.000 228.200 ;
        RECT 44.500 227.200 44.800 227.900 ;
        RECT 46.200 227.600 46.600 229.900 ;
        RECT 45.300 227.300 46.600 227.600 ;
        RECT 35.800 225.800 37.800 226.100 ;
        RECT 38.200 226.100 38.600 226.200 ;
        RECT 39.000 226.100 39.400 226.600 ;
        RECT 38.200 225.800 39.400 226.100 ;
        RECT 39.800 225.800 40.200 226.600 ;
        RECT 40.600 226.500 41.300 226.900 ;
        RECT 41.600 226.800 42.600 227.200 ;
        RECT 43.000 227.100 43.400 227.200 ;
        RECT 44.500 227.100 45.000 227.200 ;
        RECT 43.000 226.800 45.000 227.100 ;
        RECT 35.800 225.400 36.200 225.800 ;
        RECT 34.700 224.600 35.500 224.900 ;
        RECT 34.700 224.200 35.100 224.600 ;
        RECT 34.200 223.800 35.100 224.200 ;
        RECT 32.600 221.500 33.000 223.500 ;
        RECT 34.700 221.100 35.100 223.800 ;
        RECT 37.400 221.100 37.800 225.800 ;
        RECT 40.600 225.500 40.900 226.500 ;
        RECT 39.000 225.200 40.900 225.500 ;
        RECT 39.000 223.500 39.300 225.200 ;
        RECT 41.600 224.900 41.900 226.800 ;
        RECT 42.200 225.400 42.600 226.200 ;
        RECT 41.100 224.600 41.900 224.900 ;
        RECT 44.500 225.100 44.800 226.800 ;
        RECT 45.300 226.500 45.600 227.300 ;
        RECT 45.100 226.100 45.600 226.500 ;
        RECT 45.300 225.100 45.600 226.100 ;
        RECT 46.100 226.200 46.500 226.600 ;
        RECT 46.100 225.800 46.600 226.200 ;
        RECT 44.500 224.600 45.000 225.100 ;
        RECT 45.300 224.800 46.600 225.100 ;
        RECT 39.000 221.500 39.400 223.500 ;
        RECT 41.100 222.200 41.500 224.600 ;
        RECT 40.600 221.800 41.500 222.200 ;
        RECT 41.100 221.100 41.500 221.800 ;
        RECT 44.600 221.100 45.000 224.600 ;
        RECT 46.200 221.100 46.600 224.800 ;
        RECT 47.000 221.100 47.400 229.900 ;
        RECT 47.800 227.800 48.200 228.600 ;
        RECT 49.400 227.600 49.800 229.900 ;
        RECT 51.000 227.600 51.400 229.900 ;
        RECT 49.400 227.200 51.400 227.600 ;
        RECT 54.200 227.500 54.600 229.900 ;
        RECT 56.400 229.200 56.800 229.900 ;
        RECT 55.800 228.900 56.800 229.200 ;
        RECT 58.600 228.900 59.000 229.900 ;
        RECT 60.700 229.200 61.300 229.900 ;
        RECT 60.600 228.900 61.300 229.200 ;
        RECT 55.800 228.500 56.200 228.900 ;
        RECT 58.600 228.600 58.900 228.900 ;
        RECT 56.600 228.200 57.000 228.600 ;
        RECT 57.500 228.300 58.900 228.600 ;
        RECT 60.600 228.500 61.000 228.900 ;
        RECT 57.500 228.200 57.900 228.300 ;
        RECT 56.700 227.200 57.000 228.200 ;
        RECT 61.500 227.700 61.900 227.800 ;
        RECT 63.000 227.700 63.400 229.900 ;
        RECT 63.800 228.000 64.200 229.900 ;
        RECT 65.400 228.000 65.800 229.900 ;
        RECT 63.800 227.900 65.800 228.000 ;
        RECT 66.200 227.900 66.600 229.900 ;
        RECT 67.300 228.200 67.700 229.900 ;
        RECT 67.300 227.900 68.200 228.200 ;
        RECT 71.300 228.000 71.700 229.500 ;
        RECT 73.400 228.500 73.800 229.500 ;
        RECT 63.900 227.700 65.700 227.900 ;
        RECT 61.500 227.400 63.400 227.700 ;
        RECT 51.000 225.800 51.400 227.200 ;
        RECT 54.600 227.100 55.400 227.200 ;
        RECT 56.600 227.100 57.000 227.200 ;
        RECT 59.500 227.100 59.900 227.200 ;
        RECT 54.600 226.800 60.100 227.100 ;
        RECT 56.100 226.700 56.500 226.800 ;
        RECT 55.300 226.200 55.700 226.300 ;
        RECT 55.300 225.900 57.800 226.200 ;
        RECT 57.400 225.800 57.800 225.900 ;
        RECT 49.400 225.400 51.400 225.800 ;
        RECT 49.400 221.100 49.800 225.400 ;
        RECT 51.000 221.100 51.400 225.400 ;
        RECT 54.200 225.500 57.000 225.600 ;
        RECT 54.200 225.400 57.100 225.500 ;
        RECT 54.200 225.300 59.100 225.400 ;
        RECT 54.200 221.100 54.600 225.300 ;
        RECT 56.700 225.100 59.100 225.300 ;
        RECT 55.800 224.500 58.500 224.800 ;
        RECT 55.800 224.400 56.200 224.500 ;
        RECT 58.100 224.400 58.500 224.500 ;
        RECT 58.800 224.500 59.100 225.100 ;
        RECT 59.800 225.200 60.100 226.800 ;
        RECT 60.600 226.400 61.000 226.500 ;
        RECT 60.600 226.100 62.500 226.400 ;
        RECT 62.100 226.000 62.500 226.100 ;
        RECT 61.300 225.700 61.700 225.800 ;
        RECT 63.000 225.700 63.400 227.400 ;
        RECT 64.200 227.200 64.600 227.400 ;
        RECT 66.200 227.200 66.500 227.900 ;
        RECT 63.800 226.900 64.600 227.200 ;
        RECT 63.800 226.800 64.200 226.900 ;
        RECT 65.300 226.800 66.600 227.200 ;
        RECT 64.600 225.800 65.000 226.600 ;
        RECT 61.300 225.400 63.400 225.700 ;
        RECT 59.800 224.900 61.000 225.200 ;
        RECT 59.500 224.500 59.900 224.600 ;
        RECT 58.800 224.200 59.900 224.500 ;
        RECT 60.700 224.400 61.000 224.900 ;
        RECT 60.700 224.000 61.400 224.400 ;
        RECT 57.500 223.700 57.900 223.800 ;
        RECT 58.900 223.700 59.300 223.800 ;
        RECT 55.800 223.100 56.200 223.500 ;
        RECT 57.500 223.400 59.300 223.700 ;
        RECT 58.600 223.100 58.900 223.400 ;
        RECT 60.600 223.100 61.000 223.500 ;
        RECT 55.800 222.800 56.800 223.100 ;
        RECT 56.400 221.100 56.800 222.800 ;
        RECT 58.600 221.100 59.000 223.100 ;
        RECT 60.700 221.100 61.300 223.100 ;
        RECT 63.000 221.100 63.400 225.400 ;
        RECT 65.300 225.100 65.600 226.800 ;
        RECT 67.800 226.100 68.200 227.900 ;
        RECT 70.900 227.700 71.700 228.000 ;
        RECT 68.600 227.100 69.000 227.600 ;
        RECT 70.900 227.500 71.300 227.700 ;
        RECT 70.900 227.200 71.200 227.500 ;
        RECT 73.500 227.400 73.800 228.500 ;
        RECT 68.600 226.800 69.700 227.100 ;
        RECT 70.200 226.800 71.200 227.200 ;
        RECT 71.700 227.100 73.800 227.400 ;
        RECT 74.200 227.700 74.600 229.900 ;
        RECT 76.300 229.200 76.900 229.900 ;
        RECT 76.300 228.900 77.000 229.200 ;
        RECT 78.600 228.900 79.000 229.900 ;
        RECT 80.800 229.200 81.200 229.900 ;
        RECT 80.800 228.900 81.800 229.200 ;
        RECT 76.600 228.500 77.000 228.900 ;
        RECT 78.700 228.600 79.000 228.900 ;
        RECT 78.700 228.300 80.100 228.600 ;
        RECT 79.700 228.200 80.100 228.300 ;
        RECT 80.600 228.200 81.000 228.600 ;
        RECT 81.400 228.500 81.800 228.900 ;
        RECT 75.700 227.700 76.100 227.800 ;
        RECT 74.200 227.400 76.100 227.700 ;
        RECT 71.700 226.900 72.200 227.100 ;
        RECT 66.200 225.800 68.200 226.100 ;
        RECT 69.400 226.100 69.700 226.800 ;
        RECT 70.200 226.100 70.600 226.200 ;
        RECT 69.400 225.800 70.600 226.100 ;
        RECT 66.200 225.200 66.500 225.800 ;
        RECT 66.200 225.100 66.600 225.200 ;
        RECT 65.100 224.800 65.600 225.100 ;
        RECT 65.900 224.800 66.600 225.100 ;
        RECT 65.100 221.100 65.500 224.800 ;
        RECT 65.900 224.200 66.200 224.800 ;
        RECT 67.000 224.400 67.400 225.200 ;
        RECT 65.800 223.800 66.200 224.200 ;
        RECT 67.800 221.100 68.200 225.800 ;
        RECT 70.200 225.400 70.600 225.800 ;
        RECT 70.900 224.900 71.200 226.800 ;
        RECT 71.500 226.500 72.200 226.900 ;
        RECT 71.900 225.500 72.200 226.500 ;
        RECT 72.600 225.800 73.000 226.600 ;
        RECT 73.400 225.800 73.800 226.600 ;
        RECT 74.200 225.700 74.600 227.400 ;
        RECT 77.700 227.100 78.100 227.200 ;
        RECT 79.800 227.100 80.200 227.200 ;
        RECT 80.600 227.100 80.900 228.200 ;
        RECT 83.000 227.500 83.400 229.900 ;
        RECT 84.600 228.900 85.000 229.900 ;
        RECT 83.800 227.800 84.200 228.600 ;
        RECT 84.700 228.100 85.000 228.900 ;
        RECT 86.300 228.200 86.700 228.600 ;
        RECT 86.200 228.100 86.600 228.200 ;
        RECT 84.600 227.800 86.600 228.100 ;
        RECT 87.000 227.900 87.400 229.900 ;
        RECT 84.700 227.200 85.000 227.800 ;
        RECT 87.100 227.200 87.400 227.900 ;
        RECT 90.200 227.600 90.600 229.900 ;
        RECT 91.800 227.600 92.200 229.900 ;
        RECT 93.400 227.600 93.800 229.900 ;
        RECT 95.000 227.600 95.400 229.900 ;
        RECT 90.200 227.200 91.100 227.600 ;
        RECT 91.800 227.200 92.900 227.600 ;
        RECT 93.400 227.200 94.500 227.600 ;
        RECT 95.000 227.200 96.200 227.600 ;
        RECT 96.600 227.500 97.000 229.900 ;
        RECT 98.800 229.200 99.200 229.900 ;
        RECT 98.200 228.900 99.200 229.200 ;
        RECT 101.000 228.900 101.400 229.900 ;
        RECT 103.100 229.200 103.700 229.900 ;
        RECT 103.000 228.900 103.700 229.200 ;
        RECT 98.200 228.500 98.600 228.900 ;
        RECT 101.000 228.600 101.300 228.900 ;
        RECT 99.000 228.200 99.400 228.600 ;
        RECT 99.900 228.300 101.300 228.600 ;
        RECT 103.000 228.500 103.400 228.900 ;
        RECT 99.900 228.200 100.300 228.300 ;
        RECT 82.200 227.100 83.000 227.200 ;
        RECT 77.500 226.800 83.000 227.100 ;
        RECT 84.600 226.800 85.000 227.200 ;
        RECT 87.000 226.800 87.400 227.200 ;
        RECT 76.600 226.400 77.000 226.500 ;
        RECT 75.100 226.100 77.000 226.400 ;
        RECT 75.100 226.000 75.500 226.100 ;
        RECT 75.900 225.700 76.300 225.800 ;
        RECT 71.900 225.200 73.800 225.500 ;
        RECT 70.900 224.600 71.700 224.900 ;
        RECT 71.300 222.200 71.700 224.600 ;
        RECT 73.500 223.500 73.800 225.200 ;
        RECT 71.300 221.800 72.200 222.200 ;
        RECT 71.300 221.100 71.700 221.800 ;
        RECT 73.400 221.500 73.800 223.500 ;
        RECT 74.200 225.400 76.300 225.700 ;
        RECT 74.200 221.100 74.600 225.400 ;
        RECT 77.500 225.200 77.800 226.800 ;
        RECT 81.100 226.700 81.500 226.800 ;
        RECT 80.600 226.200 81.000 226.300 ;
        RECT 81.900 226.200 82.300 226.300 ;
        RECT 79.800 225.900 82.300 226.200 ;
        RECT 79.800 225.800 80.200 225.900 ;
        RECT 80.600 225.500 83.400 225.600 ;
        RECT 80.500 225.400 83.400 225.500 ;
        RECT 76.600 224.900 77.800 225.200 ;
        RECT 78.500 225.300 83.400 225.400 ;
        RECT 78.500 225.100 80.900 225.300 ;
        RECT 76.600 224.400 76.900 224.900 ;
        RECT 76.200 224.000 76.900 224.400 ;
        RECT 77.700 224.500 78.100 224.600 ;
        RECT 78.500 224.500 78.800 225.100 ;
        RECT 77.700 224.200 78.800 224.500 ;
        RECT 79.100 224.500 81.800 224.800 ;
        RECT 79.100 224.400 79.500 224.500 ;
        RECT 81.400 224.400 81.800 224.500 ;
        RECT 78.300 223.700 78.700 223.800 ;
        RECT 79.700 223.700 80.100 223.800 ;
        RECT 76.600 223.100 77.000 223.500 ;
        RECT 78.300 223.400 80.100 223.700 ;
        RECT 78.700 223.100 79.000 223.400 ;
        RECT 81.400 223.100 81.800 223.500 ;
        RECT 76.300 221.100 76.900 223.100 ;
        RECT 78.600 221.100 79.000 223.100 ;
        RECT 80.800 222.800 81.800 223.100 ;
        RECT 80.800 221.100 81.200 222.800 ;
        RECT 83.000 221.100 83.400 225.300 ;
        RECT 84.700 225.100 85.000 226.800 ;
        RECT 85.400 225.400 85.800 226.200 ;
        RECT 86.200 226.100 86.600 226.200 ;
        RECT 87.100 226.100 87.400 226.800 ;
        RECT 87.800 226.400 88.200 227.200 ;
        RECT 89.400 226.900 89.800 227.200 ;
        RECT 90.700 226.900 91.100 227.200 ;
        RECT 92.500 226.900 92.900 227.200 ;
        RECT 94.100 226.900 94.500 227.200 ;
        RECT 89.400 226.500 90.300 226.900 ;
        RECT 90.700 226.500 92.000 226.900 ;
        RECT 92.500 226.500 93.700 226.900 ;
        RECT 94.100 226.500 95.400 226.900 ;
        RECT 88.600 226.100 89.000 226.200 ;
        RECT 86.200 225.800 87.400 226.100 ;
        RECT 88.200 225.800 89.000 226.100 ;
        RECT 90.700 225.800 91.100 226.500 ;
        RECT 92.500 225.800 92.900 226.500 ;
        RECT 94.100 225.800 94.500 226.500 ;
        RECT 95.800 225.800 96.200 227.200 ;
        RECT 97.000 227.100 97.800 227.200 ;
        RECT 99.100 227.100 99.400 228.200 ;
        RECT 103.900 227.700 104.300 227.800 ;
        RECT 105.400 227.700 105.800 229.900 ;
        RECT 103.900 227.400 105.800 227.700 ;
        RECT 101.900 227.100 102.300 227.200 ;
        RECT 97.000 226.800 102.500 227.100 ;
        RECT 98.500 226.700 98.900 226.800 ;
        RECT 97.700 226.200 98.100 226.300 ;
        RECT 97.700 226.100 100.200 226.200 ;
        RECT 100.600 226.100 101.000 226.200 ;
        RECT 97.700 225.900 101.000 226.100 ;
        RECT 99.800 225.800 101.000 225.900 ;
        RECT 86.300 225.100 86.600 225.800 ;
        RECT 88.200 225.600 88.600 225.800 ;
        RECT 90.200 225.400 91.100 225.800 ;
        RECT 91.800 225.400 92.900 225.800 ;
        RECT 93.400 225.400 94.500 225.800 ;
        RECT 95.000 225.400 96.200 225.800 ;
        RECT 96.600 225.500 99.400 225.600 ;
        RECT 96.600 225.400 99.500 225.500 ;
        RECT 84.600 224.700 85.500 225.100 ;
        RECT 85.100 221.100 85.500 224.700 ;
        RECT 86.200 221.100 86.600 225.100 ;
        RECT 87.000 224.800 89.000 225.100 ;
        RECT 87.000 221.100 87.400 224.800 ;
        RECT 88.600 221.100 89.000 224.800 ;
        RECT 90.200 221.100 90.600 225.400 ;
        RECT 91.800 221.100 92.200 225.400 ;
        RECT 93.400 221.100 93.800 225.400 ;
        RECT 95.000 221.100 95.400 225.400 ;
        RECT 96.600 225.300 101.500 225.400 ;
        RECT 96.600 221.100 97.000 225.300 ;
        RECT 99.100 225.100 101.500 225.300 ;
        RECT 98.200 224.500 100.900 224.800 ;
        RECT 98.200 224.400 98.600 224.500 ;
        RECT 100.500 224.400 100.900 224.500 ;
        RECT 101.200 224.500 101.500 225.100 ;
        RECT 102.200 225.200 102.500 226.800 ;
        RECT 103.000 226.400 103.400 226.500 ;
        RECT 103.000 226.100 104.900 226.400 ;
        RECT 104.500 226.000 104.900 226.100 ;
        RECT 103.700 225.700 104.100 225.800 ;
        RECT 105.400 225.700 105.800 227.400 ;
        RECT 107.800 228.500 108.200 229.500 ;
        RECT 109.900 229.200 110.300 229.500 ;
        RECT 113.900 229.200 114.300 229.900 ;
        RECT 109.900 228.800 110.600 229.200 ;
        RECT 113.400 228.800 114.300 229.200 ;
        RECT 107.800 227.400 108.100 228.500 ;
        RECT 109.900 228.000 110.300 228.800 ;
        RECT 113.900 228.200 114.300 228.800 ;
        RECT 109.900 227.700 110.700 228.000 ;
        RECT 110.300 227.500 110.700 227.700 ;
        RECT 113.400 227.900 114.300 228.200 ;
        RECT 107.800 227.100 109.900 227.400 ;
        RECT 109.400 226.900 109.900 227.100 ;
        RECT 110.400 227.200 110.700 227.500 ;
        RECT 107.800 225.800 108.200 226.600 ;
        RECT 108.600 225.800 109.000 226.600 ;
        RECT 109.400 226.500 110.100 226.900 ;
        RECT 110.400 226.800 111.400 227.200 ;
        RECT 112.600 227.100 113.000 227.600 ;
        RECT 111.800 226.800 113.000 227.100 ;
        RECT 103.700 225.400 105.800 225.700 ;
        RECT 109.400 225.500 109.700 226.500 ;
        RECT 102.200 224.900 103.400 225.200 ;
        RECT 101.900 224.500 102.300 224.600 ;
        RECT 101.200 224.200 102.300 224.500 ;
        RECT 103.100 224.400 103.400 224.900 ;
        RECT 103.100 224.000 103.800 224.400 ;
        RECT 105.400 224.100 105.800 225.400 ;
        RECT 107.800 225.200 109.700 225.500 ;
        RECT 107.000 224.100 107.400 224.200 ;
        RECT 105.400 223.800 107.400 224.100 ;
        RECT 99.900 223.700 100.300 223.800 ;
        RECT 101.300 223.700 101.700 223.800 ;
        RECT 98.200 223.100 98.600 223.500 ;
        RECT 99.900 223.400 101.700 223.700 ;
        RECT 101.000 223.100 101.300 223.400 ;
        RECT 103.000 223.100 103.400 223.500 ;
        RECT 98.200 222.800 99.200 223.100 ;
        RECT 98.800 221.100 99.200 222.800 ;
        RECT 101.000 221.100 101.400 223.100 ;
        RECT 103.100 221.100 103.700 223.100 ;
        RECT 105.400 221.100 105.800 223.800 ;
        RECT 107.800 223.500 108.100 225.200 ;
        RECT 110.400 224.900 110.700 226.800 ;
        RECT 111.000 226.100 111.400 226.200 ;
        RECT 111.800 226.100 112.100 226.800 ;
        RECT 111.000 225.800 112.100 226.100 ;
        RECT 111.000 225.400 111.400 225.800 ;
        RECT 109.900 224.600 110.700 224.900 ;
        RECT 107.800 221.500 108.200 223.500 ;
        RECT 109.900 221.100 110.300 224.600 ;
        RECT 113.400 221.100 113.800 227.900 ;
        RECT 115.000 227.600 115.400 229.900 ;
        RECT 116.600 228.200 117.000 229.900 ;
        RECT 116.600 227.900 117.100 228.200 ;
        RECT 115.000 227.300 116.300 227.600 ;
        RECT 115.100 226.200 115.500 226.600 ;
        RECT 115.000 225.800 115.500 226.200 ;
        RECT 116.000 226.500 116.300 227.300 ;
        RECT 116.800 227.200 117.100 227.900 ;
        RECT 119.000 227.600 119.400 229.900 ;
        RECT 120.600 227.600 121.000 229.900 ;
        RECT 124.100 228.000 124.500 229.500 ;
        RECT 126.200 228.500 126.600 229.500 ;
        RECT 119.000 227.200 121.000 227.600 ;
        RECT 123.700 227.700 124.500 228.000 ;
        RECT 123.700 227.500 124.100 227.700 ;
        RECT 123.700 227.200 124.000 227.500 ;
        RECT 126.300 227.400 126.600 228.500 ;
        RECT 116.600 226.800 117.100 227.200 ;
        RECT 116.000 226.100 116.500 226.500 ;
        RECT 114.200 224.400 114.600 225.200 ;
        RECT 116.000 225.100 116.300 226.100 ;
        RECT 116.800 225.100 117.100 226.800 ;
        RECT 120.600 225.800 121.000 227.200 ;
        RECT 123.000 226.800 124.000 227.200 ;
        RECT 124.500 227.100 126.600 227.400 ;
        RECT 127.000 228.500 127.400 229.500 ;
        RECT 127.000 227.400 127.300 228.500 ;
        RECT 129.100 228.000 129.500 229.500 ;
        RECT 131.800 228.500 132.200 229.500 ;
        RECT 129.100 227.700 129.900 228.000 ;
        RECT 129.500 227.500 129.900 227.700 ;
        RECT 127.000 227.100 129.100 227.400 ;
        RECT 124.500 226.900 125.000 227.100 ;
        RECT 122.200 226.100 122.600 226.200 ;
        RECT 123.000 226.100 123.400 226.200 ;
        RECT 122.200 225.800 123.400 226.100 ;
        RECT 115.000 224.800 116.300 225.100 ;
        RECT 115.000 221.100 115.400 224.800 ;
        RECT 116.600 224.600 117.100 225.100 ;
        RECT 119.000 225.400 121.000 225.800 ;
        RECT 123.000 225.400 123.400 225.800 ;
        RECT 116.600 221.100 117.000 224.600 ;
        RECT 119.000 221.100 119.400 225.400 ;
        RECT 120.600 221.100 121.000 225.400 ;
        RECT 123.700 224.900 124.000 226.800 ;
        RECT 124.300 226.500 125.000 226.900 ;
        RECT 128.600 226.900 129.100 227.100 ;
        RECT 129.600 227.200 129.900 227.500 ;
        RECT 131.800 227.400 132.100 228.500 ;
        RECT 133.900 228.000 134.300 229.500 ;
        RECT 137.900 228.200 138.300 229.900 ;
        RECT 133.900 227.700 134.700 228.000 ;
        RECT 134.300 227.500 134.700 227.700 ;
        RECT 137.400 227.900 138.300 228.200 ;
        RECT 139.000 227.900 139.400 229.900 ;
        RECT 139.800 228.000 140.200 229.900 ;
        RECT 141.400 228.000 141.800 229.900 ;
        RECT 139.800 227.900 141.800 228.000 ;
        RECT 124.700 225.500 125.000 226.500 ;
        RECT 125.400 225.800 125.800 226.600 ;
        RECT 126.200 225.800 126.600 226.600 ;
        RECT 127.000 225.800 127.400 226.600 ;
        RECT 127.800 225.800 128.200 226.600 ;
        RECT 128.600 226.500 129.300 226.900 ;
        RECT 129.600 226.800 130.600 227.200 ;
        RECT 131.800 227.100 133.900 227.400 ;
        RECT 133.400 226.900 133.900 227.100 ;
        RECT 134.400 227.200 134.700 227.500 ;
        RECT 128.600 225.500 128.900 226.500 ;
        RECT 124.700 225.200 126.600 225.500 ;
        RECT 123.700 224.600 124.500 224.900 ;
        RECT 124.100 222.200 124.500 224.600 ;
        RECT 126.300 223.500 126.600 225.200 ;
        RECT 123.800 221.800 124.500 222.200 ;
        RECT 124.100 221.100 124.500 221.800 ;
        RECT 126.200 221.500 126.600 223.500 ;
        RECT 127.000 225.200 128.900 225.500 ;
        RECT 127.000 223.500 127.300 225.200 ;
        RECT 129.600 224.900 129.900 226.800 ;
        RECT 130.200 225.400 130.600 226.200 ;
        RECT 131.800 225.800 132.200 226.600 ;
        RECT 132.600 225.800 133.000 226.600 ;
        RECT 133.400 226.500 134.100 226.900 ;
        RECT 134.400 226.800 135.400 227.200 ;
        RECT 135.800 227.100 136.200 227.200 ;
        RECT 136.600 227.100 137.000 227.600 ;
        RECT 135.800 226.800 137.000 227.100 ;
        RECT 133.400 225.500 133.700 226.500 ;
        RECT 129.100 224.600 129.900 224.900 ;
        RECT 131.800 225.200 133.700 225.500 ;
        RECT 127.000 221.500 127.400 223.500 ;
        RECT 129.100 222.200 129.500 224.600 ;
        RECT 131.800 223.500 132.100 225.200 ;
        RECT 134.400 224.900 134.700 226.800 ;
        RECT 135.000 226.100 135.400 226.200 ;
        RECT 136.600 226.100 137.000 226.200 ;
        RECT 135.000 225.800 137.000 226.100 ;
        RECT 137.400 226.100 137.800 227.900 ;
        RECT 139.100 227.200 139.400 227.900 ;
        RECT 139.900 227.700 141.700 227.900 ;
        RECT 142.200 227.700 142.600 229.900 ;
        RECT 144.300 229.200 144.900 229.900 ;
        RECT 144.300 228.900 145.000 229.200 ;
        RECT 146.600 228.900 147.000 229.900 ;
        RECT 148.800 229.200 149.200 229.900 ;
        RECT 148.800 228.900 149.800 229.200 ;
        RECT 144.600 228.500 145.000 228.900 ;
        RECT 146.700 228.600 147.000 228.900 ;
        RECT 146.700 228.300 148.100 228.600 ;
        RECT 147.700 228.200 148.100 228.300 ;
        RECT 148.600 228.200 149.000 228.600 ;
        RECT 149.400 228.500 149.800 228.900 ;
        RECT 143.700 227.700 144.100 227.800 ;
        RECT 142.200 227.400 144.100 227.700 ;
        RECT 141.000 227.200 141.400 227.400 ;
        RECT 139.000 226.800 140.300 227.200 ;
        RECT 141.000 226.900 141.800 227.200 ;
        RECT 141.400 226.800 141.800 226.900 ;
        RECT 137.400 225.800 139.300 226.100 ;
        RECT 135.000 225.400 135.400 225.800 ;
        RECT 133.900 224.600 134.700 224.900 ;
        RECT 129.100 221.800 129.800 222.200 ;
        RECT 129.100 221.100 129.500 221.800 ;
        RECT 131.800 221.500 132.200 223.500 ;
        RECT 133.900 222.200 134.300 224.600 ;
        RECT 133.900 221.800 134.600 222.200 ;
        RECT 133.900 221.100 134.300 221.800 ;
        RECT 137.400 221.100 137.800 225.800 ;
        RECT 139.000 225.200 139.300 225.800 ;
        RECT 140.000 225.200 140.300 226.800 ;
        RECT 140.600 225.800 141.000 226.600 ;
        RECT 142.200 225.700 142.600 227.400 ;
        RECT 148.600 227.200 148.900 228.200 ;
        RECT 151.000 227.500 151.400 229.900 ;
        RECT 151.800 228.500 152.200 229.500 ;
        RECT 151.800 227.400 152.100 228.500 ;
        RECT 153.900 228.000 154.300 229.500 ;
        RECT 160.100 228.000 160.500 229.500 ;
        RECT 162.200 228.500 162.600 229.500 ;
        RECT 153.900 227.700 154.700 228.000 ;
        RECT 154.300 227.500 154.700 227.700 ;
        RECT 145.700 227.100 146.100 227.200 ;
        RECT 148.600 227.100 149.000 227.200 ;
        RECT 150.200 227.100 151.000 227.200 ;
        RECT 151.800 227.100 153.900 227.400 ;
        RECT 145.500 226.800 151.000 227.100 ;
        RECT 153.400 226.900 153.900 227.100 ;
        RECT 154.400 227.200 154.700 227.500 ;
        RECT 159.700 227.700 160.500 228.000 ;
        RECT 159.700 227.500 160.100 227.700 ;
        RECT 159.700 227.200 160.000 227.500 ;
        RECT 162.300 227.400 162.600 228.500 ;
        RECT 144.600 226.400 145.000 226.500 ;
        RECT 143.100 226.100 145.000 226.400 ;
        RECT 143.100 226.000 143.500 226.100 ;
        RECT 143.900 225.700 144.300 225.800 ;
        RECT 142.200 225.400 144.300 225.700 ;
        RECT 138.200 224.400 138.600 225.200 ;
        RECT 139.000 225.100 139.400 225.200 ;
        RECT 139.000 224.800 139.700 225.100 ;
        RECT 140.000 224.800 141.000 225.200 ;
        RECT 139.400 224.200 139.700 224.800 ;
        RECT 139.400 223.800 139.800 224.200 ;
        RECT 140.100 221.100 140.500 224.800 ;
        RECT 142.200 221.100 142.600 225.400 ;
        RECT 145.500 225.200 145.800 226.800 ;
        RECT 149.100 226.700 149.500 226.800 ;
        RECT 149.900 226.200 150.300 226.300 ;
        RECT 147.800 225.900 150.300 226.200 ;
        RECT 147.800 225.800 148.200 225.900 ;
        RECT 151.800 225.800 152.200 226.600 ;
        RECT 152.600 225.800 153.000 226.600 ;
        RECT 153.400 226.500 154.100 226.900 ;
        RECT 154.400 226.800 155.400 227.200 ;
        RECT 155.800 227.100 156.200 227.200 ;
        RECT 159.000 227.100 160.000 227.200 ;
        RECT 155.800 226.800 160.000 227.100 ;
        RECT 160.500 227.100 162.600 227.400 ;
        RECT 163.000 227.700 163.400 229.900 ;
        RECT 165.100 229.200 165.700 229.900 ;
        RECT 165.100 228.900 165.800 229.200 ;
        RECT 167.400 228.900 167.800 229.900 ;
        RECT 169.600 229.200 170.000 229.900 ;
        RECT 169.600 228.900 170.600 229.200 ;
        RECT 165.400 228.500 165.800 228.900 ;
        RECT 167.500 228.600 167.800 228.900 ;
        RECT 167.500 228.300 168.900 228.600 ;
        RECT 168.500 228.200 168.900 228.300 ;
        RECT 169.400 228.200 169.800 228.600 ;
        RECT 170.200 228.500 170.600 228.900 ;
        RECT 164.500 227.700 164.900 227.800 ;
        RECT 163.000 227.400 164.900 227.700 ;
        RECT 160.500 226.900 161.000 227.100 ;
        RECT 148.600 225.500 151.400 225.600 ;
        RECT 153.400 225.500 153.700 226.500 ;
        RECT 148.500 225.400 151.400 225.500 ;
        RECT 144.600 224.900 145.800 225.200 ;
        RECT 146.500 225.300 151.400 225.400 ;
        RECT 146.500 225.100 148.900 225.300 ;
        RECT 144.600 224.400 144.900 224.900 ;
        RECT 144.200 224.000 144.900 224.400 ;
        RECT 145.700 224.500 146.100 224.600 ;
        RECT 146.500 224.500 146.800 225.100 ;
        RECT 145.700 224.200 146.800 224.500 ;
        RECT 147.100 224.500 149.800 224.800 ;
        RECT 147.100 224.400 147.500 224.500 ;
        RECT 149.400 224.400 149.800 224.500 ;
        RECT 146.300 223.700 146.700 223.800 ;
        RECT 147.700 223.700 148.100 223.800 ;
        RECT 144.600 223.100 145.000 223.500 ;
        RECT 146.300 223.400 148.100 223.700 ;
        RECT 146.700 223.100 147.000 223.400 ;
        RECT 149.400 223.100 149.800 223.500 ;
        RECT 144.300 221.100 144.900 223.100 ;
        RECT 146.600 221.100 147.000 223.100 ;
        RECT 148.800 222.800 149.800 223.100 ;
        RECT 148.800 221.100 149.200 222.800 ;
        RECT 151.000 221.100 151.400 225.300 ;
        RECT 151.800 225.200 153.700 225.500 ;
        RECT 151.800 223.500 152.100 225.200 ;
        RECT 154.400 224.900 154.700 226.800 ;
        RECT 155.000 225.400 155.400 226.200 ;
        RECT 159.000 225.400 159.400 226.200 ;
        RECT 153.900 224.600 154.700 224.900 ;
        RECT 159.700 224.900 160.000 226.800 ;
        RECT 160.300 226.500 161.000 226.900 ;
        RECT 160.700 225.500 161.000 226.500 ;
        RECT 161.400 225.800 161.800 226.600 ;
        RECT 162.200 225.800 162.600 226.600 ;
        RECT 163.000 225.700 163.400 227.400 ;
        RECT 166.500 227.100 166.900 227.200 ;
        RECT 168.600 227.100 169.000 227.200 ;
        RECT 169.400 227.100 169.700 228.200 ;
        RECT 171.800 227.500 172.200 229.900 ;
        RECT 173.400 228.900 173.800 229.900 ;
        RECT 172.600 227.800 173.000 228.600 ;
        RECT 173.500 228.100 173.800 228.900 ;
        RECT 175.100 228.200 175.500 228.600 ;
        RECT 175.000 228.100 175.400 228.200 ;
        RECT 173.400 227.800 175.400 228.100 ;
        RECT 175.800 227.900 176.200 229.900 ;
        RECT 180.100 228.000 180.500 229.500 ;
        RECT 182.200 228.500 182.600 229.500 ;
        RECT 173.500 227.200 173.800 227.800 ;
        RECT 171.000 227.100 171.800 227.200 ;
        RECT 166.300 226.800 171.800 227.100 ;
        RECT 173.400 226.800 173.800 227.200 ;
        RECT 165.400 226.400 165.800 226.500 ;
        RECT 163.900 226.100 165.800 226.400 ;
        RECT 166.300 226.200 166.600 226.800 ;
        RECT 169.900 226.700 170.300 226.800 ;
        RECT 169.400 226.200 169.800 226.300 ;
        RECT 170.700 226.200 171.100 226.300 ;
        RECT 163.900 226.000 164.300 226.100 ;
        RECT 166.200 225.800 166.600 226.200 ;
        RECT 168.600 225.900 171.100 226.200 ;
        RECT 168.600 225.800 169.000 225.900 ;
        RECT 164.700 225.700 165.100 225.800 ;
        RECT 160.700 225.200 162.600 225.500 ;
        RECT 159.700 224.600 160.500 224.900 ;
        RECT 151.800 221.500 152.200 223.500 ;
        RECT 153.900 222.200 154.300 224.600 ;
        RECT 153.400 221.800 154.300 222.200 ;
        RECT 153.900 221.100 154.300 221.800 ;
        RECT 160.100 221.100 160.500 224.600 ;
        RECT 162.300 223.500 162.600 225.200 ;
        RECT 162.200 221.500 162.600 223.500 ;
        RECT 163.000 225.400 165.100 225.700 ;
        RECT 163.000 221.100 163.400 225.400 ;
        RECT 166.300 225.200 166.600 225.800 ;
        RECT 169.400 225.500 172.200 225.600 ;
        RECT 169.300 225.400 172.200 225.500 ;
        RECT 165.400 224.900 166.600 225.200 ;
        RECT 167.300 225.300 172.200 225.400 ;
        RECT 167.300 225.100 169.700 225.300 ;
        RECT 165.400 224.400 165.700 224.900 ;
        RECT 165.000 224.000 165.700 224.400 ;
        RECT 166.500 224.500 166.900 224.600 ;
        RECT 167.300 224.500 167.600 225.100 ;
        RECT 166.500 224.200 167.600 224.500 ;
        RECT 167.900 224.500 170.600 224.800 ;
        RECT 167.900 224.400 168.300 224.500 ;
        RECT 170.200 224.400 170.600 224.500 ;
        RECT 167.100 223.700 167.500 223.800 ;
        RECT 168.500 223.700 168.900 223.800 ;
        RECT 165.400 223.100 165.800 223.500 ;
        RECT 167.100 223.400 168.900 223.700 ;
        RECT 167.500 223.100 167.800 223.400 ;
        RECT 170.200 223.100 170.600 223.500 ;
        RECT 165.100 221.100 165.700 223.100 ;
        RECT 167.400 221.100 167.800 223.100 ;
        RECT 169.600 222.800 170.600 223.100 ;
        RECT 169.600 221.100 170.000 222.800 ;
        RECT 171.800 221.100 172.200 225.300 ;
        RECT 173.500 225.100 173.800 226.800 ;
        RECT 174.200 225.400 174.600 226.200 ;
        RECT 175.000 226.100 175.400 226.200 ;
        RECT 175.900 226.100 176.200 227.900 ;
        RECT 179.700 227.700 180.500 228.000 ;
        RECT 179.700 227.500 180.100 227.700 ;
        RECT 179.700 227.200 180.000 227.500 ;
        RECT 182.300 227.400 182.600 228.500 ;
        RECT 183.300 228.200 183.700 229.900 ;
        RECT 183.300 227.900 184.200 228.200 ;
        RECT 176.600 226.400 177.000 227.200 ;
        RECT 178.200 227.100 178.600 227.200 ;
        RECT 179.000 227.100 180.000 227.200 ;
        RECT 178.200 226.800 180.000 227.100 ;
        RECT 180.500 227.100 182.600 227.400 ;
        RECT 180.500 226.900 181.000 227.100 ;
        RECT 177.400 226.100 177.800 226.200 ;
        RECT 178.200 226.100 178.600 226.200 ;
        RECT 175.000 225.800 176.200 226.100 ;
        RECT 177.000 225.800 178.600 226.100 ;
        RECT 175.100 225.100 175.400 225.800 ;
        RECT 177.000 225.600 177.400 225.800 ;
        RECT 179.000 225.400 179.400 226.200 ;
        RECT 173.400 224.700 174.300 225.100 ;
        RECT 173.900 221.100 174.300 224.700 ;
        RECT 175.000 221.100 175.400 225.100 ;
        RECT 175.800 224.800 177.800 225.100 ;
        RECT 175.800 221.100 176.200 224.800 ;
        RECT 177.400 221.100 177.800 224.800 ;
        RECT 179.700 224.900 180.000 226.800 ;
        RECT 180.300 226.500 181.000 226.900 ;
        RECT 180.700 225.500 181.000 226.500 ;
        RECT 181.400 225.800 181.800 226.600 ;
        RECT 182.200 225.800 182.600 226.600 ;
        RECT 180.700 225.200 182.600 225.500 ;
        RECT 179.700 224.600 180.500 224.900 ;
        RECT 180.100 221.100 180.500 224.600 ;
        RECT 182.300 223.500 182.600 225.200 ;
        RECT 183.000 224.400 183.400 225.200 ;
        RECT 182.200 221.500 182.600 223.500 ;
        RECT 183.800 221.100 184.200 227.900 ;
        RECT 185.400 227.700 185.800 229.900 ;
        RECT 187.500 229.200 188.100 229.900 ;
        RECT 187.500 228.900 188.200 229.200 ;
        RECT 189.800 228.900 190.200 229.900 ;
        RECT 192.000 229.200 192.400 229.900 ;
        RECT 192.000 228.900 193.000 229.200 ;
        RECT 187.800 228.500 188.200 228.900 ;
        RECT 189.900 228.600 190.200 228.900 ;
        RECT 189.900 228.300 191.300 228.600 ;
        RECT 190.900 228.200 191.300 228.300 ;
        RECT 191.800 228.200 192.200 228.600 ;
        RECT 192.600 228.500 193.000 228.900 ;
        RECT 186.900 227.700 187.300 227.800 ;
        RECT 184.600 227.100 185.000 227.600 ;
        RECT 185.400 227.400 187.300 227.700 ;
        RECT 185.400 227.100 185.800 227.400 ;
        RECT 188.900 227.100 189.300 227.200 ;
        RECT 191.000 227.100 191.400 227.200 ;
        RECT 191.800 227.100 192.100 228.200 ;
        RECT 194.200 227.500 194.600 229.900 ;
        RECT 195.800 228.900 196.200 229.900 ;
        RECT 195.000 227.800 195.400 228.600 ;
        RECT 195.900 228.100 196.200 228.900 ;
        RECT 197.500 228.200 197.900 228.600 ;
        RECT 197.400 228.100 197.800 228.200 ;
        RECT 195.800 227.800 197.800 228.100 ;
        RECT 198.200 227.900 198.600 229.900 ;
        RECT 195.900 227.200 196.200 227.800 ;
        RECT 193.400 227.100 194.200 227.200 ;
        RECT 184.600 226.800 185.800 227.100 ;
        RECT 184.600 226.200 184.900 226.800 ;
        RECT 184.600 225.800 185.000 226.200 ;
        RECT 185.400 225.700 185.800 226.800 ;
        RECT 188.700 226.800 194.200 227.100 ;
        RECT 195.800 226.800 196.200 227.200 ;
        RECT 187.800 226.400 188.200 226.500 ;
        RECT 186.300 226.100 188.200 226.400 ;
        RECT 186.300 226.000 186.700 226.100 ;
        RECT 187.100 225.700 187.500 225.800 ;
        RECT 185.400 225.400 187.500 225.700 ;
        RECT 185.400 221.100 185.800 225.400 ;
        RECT 188.700 225.200 189.000 226.800 ;
        RECT 192.300 226.700 192.700 226.800 ;
        RECT 193.100 226.200 193.500 226.300 ;
        RECT 190.200 226.100 190.600 226.200 ;
        RECT 191.000 226.100 193.500 226.200 ;
        RECT 190.200 225.900 193.500 226.100 ;
        RECT 190.200 225.800 191.400 225.900 ;
        RECT 191.800 225.500 194.600 225.600 ;
        RECT 191.700 225.400 194.600 225.500 ;
        RECT 187.800 224.900 189.000 225.200 ;
        RECT 189.700 225.300 194.600 225.400 ;
        RECT 189.700 225.100 192.100 225.300 ;
        RECT 187.800 224.400 188.100 224.900 ;
        RECT 187.400 224.000 188.100 224.400 ;
        RECT 188.900 224.500 189.300 224.600 ;
        RECT 189.700 224.500 190.000 225.100 ;
        RECT 188.900 224.200 190.000 224.500 ;
        RECT 190.300 224.500 193.000 224.800 ;
        RECT 190.300 224.400 190.700 224.500 ;
        RECT 192.600 224.400 193.000 224.500 ;
        RECT 189.500 223.700 189.900 223.800 ;
        RECT 190.900 223.700 191.300 223.800 ;
        RECT 187.800 223.100 188.200 223.500 ;
        RECT 189.500 223.400 191.300 223.700 ;
        RECT 189.900 223.100 190.200 223.400 ;
        RECT 192.600 223.100 193.000 223.500 ;
        RECT 187.500 221.100 188.100 223.100 ;
        RECT 189.800 221.100 190.200 223.100 ;
        RECT 192.000 222.800 193.000 223.100 ;
        RECT 192.000 221.100 192.400 222.800 ;
        RECT 194.200 221.100 194.600 225.300 ;
        RECT 195.900 225.100 196.200 226.800 ;
        RECT 196.600 225.400 197.000 226.200 ;
        RECT 197.400 226.100 197.800 226.200 ;
        RECT 198.300 226.100 198.600 227.900 ;
        RECT 200.600 227.700 201.000 229.900 ;
        RECT 202.700 229.200 203.300 229.900 ;
        RECT 202.700 228.900 203.400 229.200 ;
        RECT 205.000 228.900 205.400 229.900 ;
        RECT 207.200 229.200 207.600 229.900 ;
        RECT 207.200 228.900 208.200 229.200 ;
        RECT 203.000 228.500 203.400 228.900 ;
        RECT 205.100 228.600 205.400 228.900 ;
        RECT 205.100 228.300 206.500 228.600 ;
        RECT 206.100 228.200 206.500 228.300 ;
        RECT 207.000 228.200 207.400 228.600 ;
        RECT 207.800 228.500 208.200 228.900 ;
        RECT 202.100 227.700 202.500 227.800 ;
        RECT 200.600 227.400 202.500 227.700 ;
        RECT 199.000 226.400 199.400 227.200 ;
        RECT 199.800 226.100 200.200 226.200 ;
        RECT 197.400 225.800 198.600 226.100 ;
        RECT 199.400 225.800 200.200 226.100 ;
        RECT 197.500 225.100 197.800 225.800 ;
        RECT 199.400 225.600 199.800 225.800 ;
        RECT 200.600 225.700 201.000 227.400 ;
        RECT 204.100 227.100 204.500 227.200 ;
        RECT 207.000 227.100 207.300 228.200 ;
        RECT 209.400 227.500 209.800 229.900 ;
        RECT 212.600 228.900 213.000 229.900 ;
        RECT 210.200 228.100 210.600 228.200 ;
        RECT 211.800 228.100 212.200 228.600 ;
        RECT 212.700 228.100 213.000 228.900 ;
        RECT 214.300 228.200 214.700 228.600 ;
        RECT 214.200 228.100 214.600 228.200 ;
        RECT 210.200 227.800 212.200 228.100 ;
        RECT 212.600 227.800 214.600 228.100 ;
        RECT 215.000 227.800 215.400 229.900 ;
        RECT 212.700 227.200 213.000 227.800 ;
        RECT 208.600 227.100 209.400 227.200 ;
        RECT 203.900 226.800 209.400 227.100 ;
        RECT 212.600 226.800 213.000 227.200 ;
        RECT 203.000 226.400 203.400 226.500 ;
        RECT 201.500 226.100 203.400 226.400 ;
        RECT 201.500 226.000 201.900 226.100 ;
        RECT 202.300 225.700 202.700 225.800 ;
        RECT 200.600 225.400 202.700 225.700 ;
        RECT 195.800 224.700 196.700 225.100 ;
        RECT 196.300 221.100 196.700 224.700 ;
        RECT 197.400 221.100 197.800 225.100 ;
        RECT 198.200 224.800 200.200 225.100 ;
        RECT 198.200 221.100 198.600 224.800 ;
        RECT 199.800 221.100 200.200 224.800 ;
        RECT 200.600 221.100 201.000 225.400 ;
        RECT 203.900 225.200 204.200 226.800 ;
        RECT 207.500 226.700 207.900 226.800 ;
        RECT 207.000 226.200 207.400 226.300 ;
        RECT 208.300 226.200 208.700 226.300 ;
        RECT 206.200 225.900 208.700 226.200 ;
        RECT 206.200 225.800 206.600 225.900 ;
        RECT 207.000 225.500 209.800 225.600 ;
        RECT 206.900 225.400 209.800 225.500 ;
        RECT 203.000 224.900 204.200 225.200 ;
        RECT 204.900 225.300 209.800 225.400 ;
        RECT 204.900 225.100 207.300 225.300 ;
        RECT 203.000 224.400 203.300 224.900 ;
        RECT 202.600 224.000 203.300 224.400 ;
        RECT 204.100 224.500 204.500 224.600 ;
        RECT 204.900 224.500 205.200 225.100 ;
        RECT 204.100 224.200 205.200 224.500 ;
        RECT 205.500 224.500 208.200 224.800 ;
        RECT 205.500 224.400 205.900 224.500 ;
        RECT 207.800 224.400 208.200 224.500 ;
        RECT 204.700 223.700 205.100 223.800 ;
        RECT 206.100 223.700 206.500 223.800 ;
        RECT 203.000 223.100 203.400 223.500 ;
        RECT 204.700 223.400 206.500 223.700 ;
        RECT 205.100 223.100 205.400 223.400 ;
        RECT 207.800 223.100 208.200 223.500 ;
        RECT 202.700 221.100 203.300 223.100 ;
        RECT 205.000 221.100 205.400 223.100 ;
        RECT 207.200 222.800 208.200 223.100 ;
        RECT 207.200 221.100 207.600 222.800 ;
        RECT 209.400 221.100 209.800 225.300 ;
        RECT 212.700 225.100 213.000 226.800 ;
        RECT 213.400 225.400 213.800 226.200 ;
        RECT 214.200 226.100 214.600 226.200 ;
        RECT 215.100 226.100 215.400 227.800 ;
        RECT 217.400 227.500 217.800 229.900 ;
        RECT 219.600 229.200 220.000 229.900 ;
        RECT 219.000 228.900 220.000 229.200 ;
        RECT 221.800 228.900 222.200 229.900 ;
        RECT 223.900 229.200 224.500 229.900 ;
        RECT 223.800 228.900 224.500 229.200 ;
        RECT 219.000 228.500 219.400 228.900 ;
        RECT 221.800 228.600 222.100 228.900 ;
        RECT 219.800 228.200 220.200 228.600 ;
        RECT 220.700 228.300 222.100 228.600 ;
        RECT 223.800 228.500 224.200 228.900 ;
        RECT 220.700 228.200 221.100 228.300 ;
        RECT 215.800 226.400 216.200 227.200 ;
        RECT 217.800 227.100 218.600 227.200 ;
        RECT 219.900 227.100 220.200 228.200 ;
        RECT 224.700 227.700 225.100 227.800 ;
        RECT 226.200 227.700 226.600 229.900 ;
        RECT 224.700 227.400 226.600 227.700 ;
        RECT 220.600 227.100 221.000 227.200 ;
        RECT 222.700 227.100 223.100 227.200 ;
        RECT 217.800 226.800 223.300 227.100 ;
        RECT 219.300 226.700 219.700 226.800 ;
        RECT 218.500 226.200 218.900 226.300 ;
        RECT 216.600 226.100 217.000 226.200 ;
        RECT 214.200 225.800 215.400 226.100 ;
        RECT 216.200 225.800 217.000 226.100 ;
        RECT 218.500 226.100 221.000 226.200 ;
        RECT 221.400 226.100 221.800 226.200 ;
        RECT 218.500 225.900 221.800 226.100 ;
        RECT 220.600 225.800 221.800 225.900 ;
        RECT 214.300 225.100 214.600 225.800 ;
        RECT 216.200 225.600 216.600 225.800 ;
        RECT 217.400 225.500 220.200 225.600 ;
        RECT 217.400 225.400 220.300 225.500 ;
        RECT 217.400 225.300 222.300 225.400 ;
        RECT 212.600 224.700 213.500 225.100 ;
        RECT 213.100 221.100 213.500 224.700 ;
        RECT 214.200 221.100 214.600 225.100 ;
        RECT 215.000 224.800 217.000 225.100 ;
        RECT 215.000 221.100 215.400 224.800 ;
        RECT 216.600 221.100 217.000 224.800 ;
        RECT 217.400 221.100 217.800 225.300 ;
        RECT 219.900 225.100 222.300 225.300 ;
        RECT 219.000 224.500 221.700 224.800 ;
        RECT 219.000 224.400 219.400 224.500 ;
        RECT 221.300 224.400 221.700 224.500 ;
        RECT 222.000 224.500 222.300 225.100 ;
        RECT 223.000 225.200 223.300 226.800 ;
        RECT 223.800 226.400 224.200 226.500 ;
        RECT 223.800 226.100 225.700 226.400 ;
        RECT 225.300 226.000 225.700 226.100 ;
        RECT 224.500 225.700 224.900 225.800 ;
        RECT 226.200 225.700 226.600 227.400 ;
        RECT 224.500 225.400 226.600 225.700 ;
        RECT 223.000 224.900 224.200 225.200 ;
        RECT 222.700 224.500 223.100 224.600 ;
        RECT 222.000 224.200 223.100 224.500 ;
        RECT 223.900 224.400 224.200 224.900 ;
        RECT 223.900 224.000 224.600 224.400 ;
        RECT 220.700 223.700 221.100 223.800 ;
        RECT 222.100 223.700 222.500 223.800 ;
        RECT 219.000 223.100 219.400 223.500 ;
        RECT 220.700 223.400 222.500 223.700 ;
        RECT 221.800 223.100 222.100 223.400 ;
        RECT 223.800 223.100 224.200 223.500 ;
        RECT 219.000 222.800 220.000 223.100 ;
        RECT 219.600 221.100 220.000 222.800 ;
        RECT 221.800 221.100 222.200 223.100 ;
        RECT 223.900 221.100 224.500 223.100 ;
        RECT 226.200 221.100 226.600 225.400 ;
        RECT 227.800 227.600 228.200 229.900 ;
        RECT 229.400 227.600 229.800 229.900 ;
        RECT 232.900 228.000 233.300 229.500 ;
        RECT 235.000 228.500 235.400 229.500 ;
        RECT 227.800 227.200 229.800 227.600 ;
        RECT 232.500 227.700 233.300 228.000 ;
        RECT 232.500 227.500 232.900 227.700 ;
        RECT 232.500 227.200 232.800 227.500 ;
        RECT 235.100 227.400 235.400 228.500 ;
        RECT 235.800 228.000 236.200 229.900 ;
        RECT 237.400 228.000 237.800 229.900 ;
        RECT 235.800 227.900 237.800 228.000 ;
        RECT 238.200 227.900 238.600 229.900 ;
        RECT 239.300 228.200 239.700 229.900 ;
        RECT 242.700 228.200 243.100 229.900 ;
        RECT 239.300 227.900 240.200 228.200 ;
        RECT 235.900 227.700 237.700 227.900 ;
        RECT 227.800 225.800 228.200 227.200 ;
        RECT 231.800 226.800 232.800 227.200 ;
        RECT 233.300 227.100 235.400 227.400 ;
        RECT 236.200 227.200 236.600 227.400 ;
        RECT 238.200 227.200 238.500 227.900 ;
        RECT 233.300 226.900 233.800 227.100 ;
        RECT 227.800 225.400 229.800 225.800 ;
        RECT 231.800 225.400 232.200 226.200 ;
        RECT 227.800 221.100 228.200 225.400 ;
        RECT 229.400 221.100 229.800 225.400 ;
        RECT 232.500 224.900 232.800 226.800 ;
        RECT 233.100 226.500 233.800 226.900 ;
        RECT 235.800 226.900 236.600 227.200 ;
        RECT 235.800 226.800 236.200 226.900 ;
        RECT 237.300 226.800 238.600 227.200 ;
        RECT 233.500 225.500 233.800 226.500 ;
        RECT 234.200 225.800 234.600 226.600 ;
        RECT 235.000 225.800 235.400 226.600 ;
        RECT 236.600 225.800 237.000 226.600 ;
        RECT 233.500 225.200 235.400 225.500 ;
        RECT 232.500 224.600 233.300 224.900 ;
        RECT 232.900 222.200 233.300 224.600 ;
        RECT 235.100 223.500 235.400 225.200 ;
        RECT 237.300 225.100 237.600 226.800 ;
        RECT 239.800 226.100 240.200 227.900 ;
        RECT 242.200 227.900 243.100 228.200 ;
        RECT 243.800 227.900 244.200 229.900 ;
        RECT 244.600 228.000 245.000 229.900 ;
        RECT 246.200 228.000 246.600 229.900 ;
        RECT 244.600 227.900 246.600 228.000 ;
        RECT 240.600 226.800 241.000 227.600 ;
        RECT 241.400 226.800 241.800 227.600 ;
        RECT 238.200 225.800 240.200 226.100 ;
        RECT 238.200 225.200 238.500 225.800 ;
        RECT 238.200 225.100 238.600 225.200 ;
        RECT 232.600 221.800 233.300 222.200 ;
        RECT 232.900 221.100 233.300 221.800 ;
        RECT 235.000 221.500 235.400 223.500 ;
        RECT 237.100 224.800 237.600 225.100 ;
        RECT 237.900 224.800 238.600 225.100 ;
        RECT 237.100 221.100 237.500 224.800 ;
        RECT 237.900 224.200 238.200 224.800 ;
        RECT 239.000 224.400 239.400 225.200 ;
        RECT 237.800 223.800 238.200 224.200 ;
        RECT 239.800 221.100 240.200 225.800 ;
        RECT 242.200 226.100 242.600 227.900 ;
        RECT 243.900 227.200 244.200 227.900 ;
        RECT 244.700 227.700 246.500 227.900 ;
        RECT 247.800 227.600 248.200 229.900 ;
        RECT 249.400 227.600 249.800 229.900 ;
        RECT 251.000 227.600 251.400 229.900 ;
        RECT 252.600 227.600 253.000 229.900 ;
        RECT 254.500 228.200 254.900 229.900 ;
        RECT 254.500 227.900 255.400 228.200 ;
        RECT 245.800 227.200 246.200 227.400 ;
        RECT 247.000 227.200 248.200 227.600 ;
        RECT 248.700 227.200 249.800 227.600 ;
        RECT 250.300 227.200 251.400 227.600 ;
        RECT 252.100 227.200 253.000 227.600 ;
        RECT 243.800 226.800 245.100 227.200 ;
        RECT 245.800 226.900 246.600 227.200 ;
        RECT 246.200 226.800 246.600 226.900 ;
        RECT 242.200 225.800 244.100 226.100 ;
        RECT 242.200 221.100 242.600 225.800 ;
        RECT 243.800 225.200 244.100 225.800 ;
        RECT 243.000 224.400 243.400 225.200 ;
        RECT 243.800 225.100 244.200 225.200 ;
        RECT 244.800 225.100 245.100 226.800 ;
        RECT 245.400 225.800 245.800 226.600 ;
        RECT 247.000 225.800 247.400 227.200 ;
        RECT 248.700 226.900 249.100 227.200 ;
        RECT 250.300 226.900 250.700 227.200 ;
        RECT 252.100 226.900 252.500 227.200 ;
        RECT 253.400 226.900 253.800 227.200 ;
        RECT 247.800 226.500 249.100 226.900 ;
        RECT 249.500 226.500 250.700 226.900 ;
        RECT 251.200 226.500 252.500 226.900 ;
        RECT 252.900 226.500 253.800 226.900 ;
        RECT 248.700 225.800 249.100 226.500 ;
        RECT 250.300 225.800 250.700 226.500 ;
        RECT 252.100 225.800 252.500 226.500 ;
        RECT 247.000 225.400 248.200 225.800 ;
        RECT 248.700 225.400 249.800 225.800 ;
        RECT 250.300 225.400 251.400 225.800 ;
        RECT 252.100 225.400 253.000 225.800 ;
        RECT 243.800 224.800 244.500 225.100 ;
        RECT 244.800 224.800 245.300 225.100 ;
        RECT 244.200 224.200 244.500 224.800 ;
        RECT 244.200 223.800 244.600 224.200 ;
        RECT 244.900 221.100 245.300 224.800 ;
        RECT 247.800 221.100 248.200 225.400 ;
        RECT 249.400 221.100 249.800 225.400 ;
        RECT 251.000 221.100 251.400 225.400 ;
        RECT 252.600 221.100 253.000 225.400 ;
        RECT 254.200 224.400 254.600 225.200 ;
        RECT 255.000 221.100 255.400 227.900 ;
        RECT 257.400 227.600 257.800 229.900 ;
        RECT 259.000 227.600 259.400 229.900 ;
        RECT 260.600 227.600 261.000 229.900 ;
        RECT 262.200 227.600 262.600 229.900 ;
        RECT 255.800 226.800 256.200 227.600 ;
        RECT 257.400 227.200 258.300 227.600 ;
        RECT 259.000 227.200 260.100 227.600 ;
        RECT 260.600 227.200 261.700 227.600 ;
        RECT 262.200 227.200 263.400 227.600 ;
        RECT 256.600 226.900 257.000 227.200 ;
        RECT 257.900 226.900 258.300 227.200 ;
        RECT 259.700 226.900 260.100 227.200 ;
        RECT 261.300 226.900 261.700 227.200 ;
        RECT 256.600 226.500 257.500 226.900 ;
        RECT 257.900 226.500 259.200 226.900 ;
        RECT 259.700 226.500 260.900 226.900 ;
        RECT 261.300 226.500 262.600 226.900 ;
        RECT 257.900 225.800 258.300 226.500 ;
        RECT 259.700 225.800 260.100 226.500 ;
        RECT 261.300 225.800 261.700 226.500 ;
        RECT 263.000 225.800 263.400 227.200 ;
        RECT 257.400 225.400 258.300 225.800 ;
        RECT 259.000 225.400 260.100 225.800 ;
        RECT 260.600 225.400 261.700 225.800 ;
        RECT 262.200 225.400 263.400 225.800 ;
        RECT 257.400 221.100 257.800 225.400 ;
        RECT 259.000 221.100 259.400 225.400 ;
        RECT 260.600 221.100 261.000 225.400 ;
        RECT 262.200 221.100 262.600 225.400 ;
        RECT 0.600 215.600 1.000 219.900 ;
        RECT 2.700 217.900 3.300 219.900 ;
        RECT 5.000 217.900 5.400 219.900 ;
        RECT 7.200 218.200 7.600 219.900 ;
        RECT 7.200 217.900 8.200 218.200 ;
        RECT 3.000 217.500 3.400 217.900 ;
        RECT 5.100 217.600 5.400 217.900 ;
        RECT 4.700 217.300 6.500 217.600 ;
        RECT 7.800 217.500 8.200 217.900 ;
        RECT 4.700 217.200 5.100 217.300 ;
        RECT 6.100 217.200 6.500 217.300 ;
        RECT 2.600 216.600 3.300 217.000 ;
        RECT 3.000 216.100 3.300 216.600 ;
        RECT 4.100 216.500 5.200 216.800 ;
        RECT 4.100 216.400 4.500 216.500 ;
        RECT 3.000 215.800 4.200 216.100 ;
        RECT 0.600 215.300 2.700 215.600 ;
        RECT 0.600 213.600 1.000 215.300 ;
        RECT 2.300 215.200 2.700 215.300 ;
        RECT 1.500 214.900 1.900 215.000 ;
        RECT 1.500 214.600 3.400 214.900 ;
        RECT 3.000 214.500 3.400 214.600 ;
        RECT 3.900 214.200 4.200 215.800 ;
        RECT 4.900 215.900 5.200 216.500 ;
        RECT 5.500 216.500 5.900 216.600 ;
        RECT 7.800 216.500 8.200 216.600 ;
        RECT 5.500 216.200 8.200 216.500 ;
        RECT 4.900 215.700 7.300 215.900 ;
        RECT 9.400 215.700 9.800 219.900 ;
        RECT 11.500 216.300 11.900 219.900 ;
        RECT 11.000 215.900 11.900 216.300 ;
        RECT 12.600 215.900 13.000 219.900 ;
        RECT 13.400 216.200 13.800 219.900 ;
        RECT 15.000 216.200 15.400 219.900 ;
        RECT 13.400 215.900 15.400 216.200 ;
        RECT 4.900 215.600 9.800 215.700 ;
        RECT 6.900 215.500 9.800 215.600 ;
        RECT 7.000 215.400 9.800 215.500 ;
        RECT 6.200 215.100 6.600 215.200 ;
        RECT 6.200 214.800 8.700 215.100 ;
        RECT 7.000 214.700 7.400 214.800 ;
        RECT 8.300 214.700 8.700 214.800 ;
        RECT 7.500 214.200 7.900 214.300 ;
        RECT 11.100 214.200 11.400 215.900 ;
        RECT 11.800 214.800 12.200 215.600 ;
        RECT 12.700 215.200 13.000 215.900 ;
        RECT 15.800 215.600 16.200 219.900 ;
        RECT 17.900 217.900 18.500 219.900 ;
        RECT 20.200 217.900 20.600 219.900 ;
        RECT 22.400 218.200 22.800 219.900 ;
        RECT 22.400 217.900 23.400 218.200 ;
        RECT 18.200 217.500 18.600 217.900 ;
        RECT 20.300 217.600 20.600 217.900 ;
        RECT 19.900 217.300 21.700 217.600 ;
        RECT 23.000 217.500 23.400 217.900 ;
        RECT 19.900 217.200 20.300 217.300 ;
        RECT 21.300 217.200 21.700 217.300 ;
        RECT 17.800 216.600 18.500 217.000 ;
        RECT 18.200 216.100 18.500 216.600 ;
        RECT 19.300 216.500 20.400 216.800 ;
        RECT 19.300 216.400 19.700 216.500 ;
        RECT 18.200 215.800 19.400 216.100 ;
        RECT 14.600 215.200 15.000 215.400 ;
        RECT 15.800 215.300 17.900 215.600 ;
        RECT 12.600 214.900 13.800 215.200 ;
        RECT 14.600 214.900 15.400 215.200 ;
        RECT 12.600 214.800 13.000 214.900 ;
        RECT 3.900 213.900 9.400 214.200 ;
        RECT 4.100 213.800 4.500 213.900 ;
        RECT 6.200 213.800 6.600 213.900 ;
        RECT 0.600 213.300 2.500 213.600 ;
        RECT 0.600 211.100 1.000 213.300 ;
        RECT 2.100 213.200 2.500 213.300 ;
        RECT 7.000 212.800 7.300 213.900 ;
        RECT 8.600 213.800 9.400 213.900 ;
        RECT 11.000 213.800 11.400 214.200 ;
        RECT 12.600 214.200 12.900 214.800 ;
        RECT 12.600 213.800 13.000 214.200 ;
        RECT 6.100 212.700 6.500 212.800 ;
        RECT 3.000 212.100 3.400 212.500 ;
        RECT 5.100 212.400 6.500 212.700 ;
        RECT 7.000 212.400 7.400 212.800 ;
        RECT 5.100 212.100 5.400 212.400 ;
        RECT 7.800 212.100 8.200 212.500 ;
        RECT 2.700 211.800 3.400 212.100 ;
        RECT 2.700 211.100 3.300 211.800 ;
        RECT 5.000 211.100 5.400 212.100 ;
        RECT 7.200 211.800 8.200 212.100 ;
        RECT 7.200 211.100 7.600 211.800 ;
        RECT 9.400 211.100 9.800 213.500 ;
        RECT 10.200 212.400 10.600 213.200 ;
        RECT 11.100 213.100 11.400 213.800 ;
        RECT 12.600 213.100 13.000 213.200 ;
        RECT 13.500 213.100 13.800 214.900 ;
        RECT 15.000 214.800 15.400 214.900 ;
        RECT 14.200 213.800 14.600 214.600 ;
        RECT 11.000 212.800 13.000 213.100 ;
        RECT 11.100 212.100 11.400 212.800 ;
        RECT 12.700 212.400 13.100 212.800 ;
        RECT 11.000 211.100 11.400 212.100 ;
        RECT 13.400 211.100 13.800 213.100 ;
        RECT 15.800 213.600 16.200 215.300 ;
        RECT 17.500 215.200 17.900 215.300 ;
        RECT 16.700 214.900 17.100 215.000 ;
        RECT 16.700 214.600 18.600 214.900 ;
        RECT 18.200 214.500 18.600 214.600 ;
        RECT 19.100 214.200 19.400 215.800 ;
        RECT 20.100 215.900 20.400 216.500 ;
        RECT 20.700 216.500 21.100 216.600 ;
        RECT 23.000 216.500 23.400 216.600 ;
        RECT 20.700 216.200 23.400 216.500 ;
        RECT 20.100 215.700 22.500 215.900 ;
        RECT 24.600 215.700 25.000 219.900 ;
        RECT 20.100 215.600 25.000 215.700 ;
        RECT 22.100 215.500 25.000 215.600 ;
        RECT 22.200 215.400 25.000 215.500 ;
        RECT 25.400 215.600 25.800 219.900 ;
        RECT 27.500 217.900 28.100 219.900 ;
        RECT 29.800 217.900 30.200 219.900 ;
        RECT 32.000 218.200 32.400 219.900 ;
        RECT 32.000 217.900 33.000 218.200 ;
        RECT 27.800 217.500 28.200 217.900 ;
        RECT 29.900 217.600 30.200 217.900 ;
        RECT 29.500 217.300 31.300 217.600 ;
        RECT 32.600 217.500 33.000 217.900 ;
        RECT 29.500 217.200 29.900 217.300 ;
        RECT 30.900 217.200 31.300 217.300 ;
        RECT 27.400 216.600 28.100 217.000 ;
        RECT 27.800 216.100 28.100 216.600 ;
        RECT 28.900 216.500 30.000 216.800 ;
        RECT 28.900 216.400 29.300 216.500 ;
        RECT 27.800 215.800 29.000 216.100 ;
        RECT 25.400 215.300 27.500 215.600 ;
        RECT 19.800 215.100 20.200 215.200 ;
        RECT 21.400 215.100 21.800 215.200 ;
        RECT 19.800 214.800 23.900 215.100 ;
        RECT 23.500 214.700 23.900 214.800 ;
        RECT 22.700 214.200 23.100 214.300 ;
        RECT 19.100 213.900 24.600 214.200 ;
        RECT 19.300 213.800 19.700 213.900 ;
        RECT 15.800 213.300 17.700 213.600 ;
        RECT 15.800 211.100 16.200 213.300 ;
        RECT 17.300 213.200 17.700 213.300 ;
        RECT 22.200 212.800 22.500 213.900 ;
        RECT 23.800 213.800 24.600 213.900 ;
        RECT 25.400 213.600 25.800 215.300 ;
        RECT 27.100 215.200 27.500 215.300 ;
        RECT 26.300 214.900 26.700 215.000 ;
        RECT 26.300 214.600 28.200 214.900 ;
        RECT 27.800 214.500 28.200 214.600 ;
        RECT 28.700 214.200 29.000 215.800 ;
        RECT 29.700 215.900 30.000 216.500 ;
        RECT 30.300 216.500 30.700 216.600 ;
        RECT 32.600 216.500 33.000 216.600 ;
        RECT 30.300 216.200 33.000 216.500 ;
        RECT 29.700 215.700 32.100 215.900 ;
        RECT 34.200 215.700 34.600 219.900 ;
        RECT 29.700 215.600 34.600 215.700 ;
        RECT 31.700 215.500 34.600 215.600 ;
        RECT 31.800 215.400 34.600 215.500 ;
        RECT 31.000 215.100 31.400 215.200 ;
        RECT 35.800 215.100 36.200 219.900 ;
        RECT 37.800 216.800 38.200 217.200 ;
        RECT 36.600 215.800 37.000 216.600 ;
        RECT 37.800 216.200 38.100 216.800 ;
        RECT 38.500 216.200 38.900 219.900 ;
        RECT 41.400 216.400 41.800 219.900 ;
        RECT 37.400 215.900 38.100 216.200 ;
        RECT 38.400 215.900 38.900 216.200 ;
        RECT 41.300 215.900 41.800 216.400 ;
        RECT 43.000 216.200 43.400 219.900 ;
        RECT 42.100 215.900 43.400 216.200 ;
        RECT 43.800 217.500 44.200 219.500 ;
        RECT 45.900 219.200 46.300 219.900 ;
        RECT 45.900 218.800 46.600 219.200 ;
        RECT 37.400 215.800 37.800 215.900 ;
        RECT 37.400 215.100 37.700 215.800 ;
        RECT 31.000 214.800 33.500 215.100 ;
        RECT 31.800 214.700 32.200 214.800 ;
        RECT 33.100 214.700 33.500 214.800 ;
        RECT 35.800 214.800 37.700 215.100 ;
        RECT 32.300 214.200 32.700 214.300 ;
        RECT 28.700 213.900 34.200 214.200 ;
        RECT 28.900 213.800 29.300 213.900 ;
        RECT 30.200 213.800 30.600 213.900 ;
        RECT 21.300 212.700 21.700 212.800 ;
        RECT 18.200 212.100 18.600 212.500 ;
        RECT 20.300 212.400 21.700 212.700 ;
        RECT 22.200 212.400 22.600 212.800 ;
        RECT 20.300 212.100 20.600 212.400 ;
        RECT 23.000 212.100 23.400 212.500 ;
        RECT 17.900 211.800 18.600 212.100 ;
        RECT 17.900 211.100 18.500 211.800 ;
        RECT 20.200 211.100 20.600 212.100 ;
        RECT 22.400 211.800 23.400 212.100 ;
        RECT 22.400 211.100 22.800 211.800 ;
        RECT 24.600 211.100 25.000 213.500 ;
        RECT 25.400 213.300 27.300 213.600 ;
        RECT 25.400 211.100 25.800 213.300 ;
        RECT 26.900 213.200 27.300 213.300 ;
        RECT 31.800 212.800 32.100 213.900 ;
        RECT 33.400 213.800 34.200 213.900 ;
        RECT 30.900 212.700 31.300 212.800 ;
        RECT 27.800 212.100 28.200 212.500 ;
        RECT 29.900 212.400 31.300 212.700 ;
        RECT 31.800 212.400 32.200 212.800 ;
        RECT 29.900 212.100 30.200 212.400 ;
        RECT 32.600 212.100 33.000 212.500 ;
        RECT 27.500 211.800 28.200 212.100 ;
        RECT 27.500 211.100 28.100 211.800 ;
        RECT 29.800 211.100 30.200 212.100 ;
        RECT 32.000 211.800 33.000 212.100 ;
        RECT 32.000 211.100 32.400 211.800 ;
        RECT 34.200 211.100 34.600 213.500 ;
        RECT 35.000 213.400 35.400 214.200 ;
        RECT 35.800 213.100 36.200 214.800 ;
        RECT 38.400 214.200 38.700 215.900 ;
        RECT 39.000 214.400 39.400 215.200 ;
        RECT 41.300 214.200 41.600 215.900 ;
        RECT 42.100 214.900 42.400 215.900 ;
        RECT 43.800 215.800 44.100 217.500 ;
        RECT 45.900 216.400 46.300 218.800 ;
        RECT 45.900 216.100 46.700 216.400 ;
        RECT 43.800 215.500 45.700 215.800 ;
        RECT 41.900 214.500 42.400 214.900 ;
        RECT 37.400 213.800 38.700 214.200 ;
        RECT 39.800 214.100 40.200 214.200 ;
        RECT 41.300 214.100 41.800 214.200 ;
        RECT 39.400 213.800 41.800 214.100 ;
        RECT 37.500 213.100 37.800 213.800 ;
        RECT 39.400 213.600 39.800 213.800 ;
        RECT 38.300 213.100 40.100 213.300 ;
        RECT 41.300 213.100 41.600 213.800 ;
        RECT 42.100 213.700 42.400 214.500 ;
        RECT 42.900 214.800 43.400 215.200 ;
        RECT 42.900 214.400 43.300 214.800 ;
        RECT 43.800 214.400 44.200 215.200 ;
        RECT 44.600 214.400 45.000 215.200 ;
        RECT 45.400 214.500 45.700 215.500 ;
        RECT 45.400 214.100 46.100 214.500 ;
        RECT 46.400 214.200 46.700 216.100 ;
        RECT 48.600 215.700 49.000 219.900 ;
        RECT 50.800 218.200 51.200 219.900 ;
        RECT 50.200 217.900 51.200 218.200 ;
        RECT 53.000 217.900 53.400 219.900 ;
        RECT 55.100 217.900 55.700 219.900 ;
        RECT 50.200 217.500 50.600 217.900 ;
        RECT 53.000 217.600 53.300 217.900 ;
        RECT 51.900 217.300 53.700 217.600 ;
        RECT 55.000 217.500 55.400 217.900 ;
        RECT 51.900 217.200 52.300 217.300 ;
        RECT 53.300 217.200 53.700 217.300 ;
        RECT 55.500 217.000 56.200 217.200 ;
        RECT 55.100 216.800 56.200 217.000 ;
        RECT 50.200 216.500 50.600 216.600 ;
        RECT 52.500 216.500 52.900 216.600 ;
        RECT 50.200 216.200 52.900 216.500 ;
        RECT 53.200 216.500 54.300 216.800 ;
        RECT 53.200 215.900 53.500 216.500 ;
        RECT 53.900 216.400 54.300 216.500 ;
        RECT 55.100 216.600 55.800 216.800 ;
        RECT 55.100 216.100 55.400 216.600 ;
        RECT 51.100 215.700 53.500 215.900 ;
        RECT 48.600 215.600 53.500 215.700 ;
        RECT 54.200 215.800 55.400 216.100 ;
        RECT 47.000 214.800 47.400 215.600 ;
        RECT 48.600 215.500 51.500 215.600 ;
        RECT 48.600 215.400 51.400 215.500 ;
        RECT 51.800 215.100 52.200 215.200 ;
        RECT 53.400 215.100 53.800 215.200 ;
        RECT 49.700 214.800 53.800 215.100 ;
        RECT 49.700 214.700 50.100 214.800 ;
        RECT 50.500 214.200 50.900 214.300 ;
        RECT 54.200 214.200 54.500 215.800 ;
        RECT 57.400 215.600 57.800 219.900 ;
        RECT 55.700 215.300 57.800 215.600 ;
        RECT 55.700 215.200 56.100 215.300 ;
        RECT 56.500 214.900 56.900 215.000 ;
        RECT 55.000 214.600 56.900 214.900 ;
        RECT 55.000 214.500 55.400 214.600 ;
        RECT 45.400 213.900 45.900 214.100 ;
        RECT 42.100 213.400 43.400 213.700 ;
        RECT 35.800 212.800 36.700 213.100 ;
        RECT 36.300 211.100 36.700 212.800 ;
        RECT 37.400 211.100 37.800 213.100 ;
        RECT 38.200 213.000 40.200 213.100 ;
        RECT 38.200 211.100 38.600 213.000 ;
        RECT 39.800 211.100 40.200 213.000 ;
        RECT 41.300 212.800 41.800 213.100 ;
        RECT 41.400 211.100 41.800 212.800 ;
        RECT 43.000 211.100 43.400 213.400 ;
        RECT 43.800 213.600 45.900 213.900 ;
        RECT 46.400 213.800 47.400 214.200 ;
        RECT 49.000 213.900 54.500 214.200 ;
        RECT 57.400 214.100 57.800 215.300 ;
        RECT 60.600 215.100 61.000 219.900 ;
        RECT 62.600 216.800 63.000 217.200 ;
        RECT 61.400 215.800 61.800 216.600 ;
        RECT 62.600 216.200 62.900 216.800 ;
        RECT 63.300 216.200 63.700 219.900 ;
        RECT 62.200 215.900 62.900 216.200 ;
        RECT 63.200 215.900 63.700 216.200 ;
        RECT 66.700 216.200 67.100 219.900 ;
        RECT 67.400 216.800 67.800 217.200 ;
        RECT 67.500 216.200 67.800 216.800 ;
        RECT 66.700 215.900 67.200 216.200 ;
        RECT 67.500 215.900 68.200 216.200 ;
        RECT 62.200 215.800 62.600 215.900 ;
        RECT 62.200 215.100 62.500 215.800 ;
        RECT 60.600 214.800 62.500 215.100 ;
        RECT 59.800 214.100 60.200 214.200 ;
        RECT 49.000 213.800 49.800 213.900 ;
        RECT 43.800 212.500 44.100 213.600 ;
        RECT 46.400 213.500 46.700 213.800 ;
        RECT 46.300 213.300 46.700 213.500 ;
        RECT 45.900 213.000 46.700 213.300 ;
        RECT 43.800 211.500 44.200 212.500 ;
        RECT 45.900 211.500 46.300 213.000 ;
        RECT 48.600 211.100 49.000 213.500 ;
        RECT 51.100 212.800 51.400 213.900 ;
        RECT 53.900 213.800 54.300 213.900 ;
        RECT 57.400 213.800 60.200 214.100 ;
        RECT 57.400 213.600 57.800 213.800 ;
        RECT 55.900 213.300 57.800 213.600 ;
        RECT 59.800 213.400 60.200 213.800 ;
        RECT 55.900 213.200 56.300 213.300 ;
        RECT 50.200 212.100 50.600 212.500 ;
        RECT 51.000 212.400 51.400 212.800 ;
        RECT 51.900 212.700 52.300 212.800 ;
        RECT 51.900 212.400 53.300 212.700 ;
        RECT 53.000 212.100 53.300 212.400 ;
        RECT 55.000 212.100 55.400 212.500 ;
        RECT 57.400 212.100 57.800 213.300 ;
        RECT 60.600 213.100 61.000 214.800 ;
        RECT 63.200 214.200 63.500 215.900 ;
        RECT 63.800 214.400 64.200 215.200 ;
        RECT 66.200 214.400 66.600 215.200 ;
        RECT 66.900 214.200 67.200 215.900 ;
        RECT 67.800 215.800 68.200 215.900 ;
        RECT 68.600 215.800 69.000 216.600 ;
        RECT 67.800 215.100 68.100 215.800 ;
        RECT 69.400 215.100 69.800 219.900 ;
        RECT 70.200 217.100 70.600 217.200 ;
        RECT 71.000 217.100 71.400 219.900 ;
        RECT 73.100 217.900 73.700 219.900 ;
        RECT 75.400 217.900 75.800 219.900 ;
        RECT 77.600 218.200 78.000 219.900 ;
        RECT 77.600 217.900 78.600 218.200 ;
        RECT 73.400 217.500 73.800 217.900 ;
        RECT 75.500 217.600 75.800 217.900 ;
        RECT 75.100 217.300 76.900 217.600 ;
        RECT 78.200 217.500 78.600 217.900 ;
        RECT 75.100 217.200 75.500 217.300 ;
        RECT 76.500 217.200 76.900 217.300 ;
        RECT 70.200 216.800 71.400 217.100 ;
        RECT 67.800 214.800 69.800 215.100 ;
        RECT 62.200 213.800 63.500 214.200 ;
        RECT 64.600 214.100 65.000 214.200 ;
        RECT 65.400 214.100 65.800 214.200 ;
        RECT 66.900 214.100 68.200 214.200 ;
        RECT 68.600 214.100 69.000 214.200 ;
        RECT 64.200 213.800 66.200 214.100 ;
        RECT 66.900 213.800 69.000 214.100 ;
        RECT 62.300 213.100 62.600 213.800 ;
        RECT 64.200 213.600 64.600 213.800 ;
        RECT 65.800 213.600 66.200 213.800 ;
        RECT 63.100 213.100 64.900 213.300 ;
        RECT 65.500 213.100 67.300 213.300 ;
        RECT 67.800 213.100 68.100 213.800 ;
        RECT 69.400 213.100 69.800 214.800 ;
        RECT 71.000 215.600 71.400 216.800 ;
        RECT 73.000 216.600 73.700 217.000 ;
        RECT 73.400 216.100 73.700 216.600 ;
        RECT 74.500 216.500 75.600 216.800 ;
        RECT 74.500 216.400 74.900 216.500 ;
        RECT 73.400 215.800 74.600 216.100 ;
        RECT 71.000 215.300 73.100 215.600 ;
        RECT 70.200 213.400 70.600 214.200 ;
        RECT 71.000 213.600 71.400 215.300 ;
        RECT 72.700 215.200 73.100 215.300 ;
        RECT 74.300 215.100 74.600 215.800 ;
        RECT 75.300 215.900 75.600 216.500 ;
        RECT 75.900 216.500 76.300 216.600 ;
        RECT 78.200 216.500 78.600 216.600 ;
        RECT 75.900 216.200 78.600 216.500 ;
        RECT 75.300 215.700 77.700 215.900 ;
        RECT 79.800 215.700 80.200 219.900 ;
        RECT 75.300 215.600 80.200 215.700 ;
        RECT 77.300 215.500 80.200 215.600 ;
        RECT 77.400 215.400 80.200 215.500 ;
        RECT 80.600 215.600 81.000 219.900 ;
        RECT 82.700 217.900 83.300 219.900 ;
        RECT 85.000 217.900 85.400 219.900 ;
        RECT 87.200 218.200 87.600 219.900 ;
        RECT 87.200 217.900 88.200 218.200 ;
        RECT 83.000 217.500 83.400 217.900 ;
        RECT 85.100 217.600 85.400 217.900 ;
        RECT 84.700 217.300 86.500 217.600 ;
        RECT 87.800 217.500 88.200 217.900 ;
        RECT 84.700 217.200 85.100 217.300 ;
        RECT 86.100 217.200 86.500 217.300 ;
        RECT 82.600 216.600 83.300 217.000 ;
        RECT 83.000 216.100 83.300 216.600 ;
        RECT 84.100 216.500 85.200 216.800 ;
        RECT 84.100 216.400 84.500 216.500 ;
        RECT 83.000 215.800 84.200 216.100 ;
        RECT 80.600 215.300 82.700 215.600 ;
        RECT 75.000 215.100 75.400 215.200 ;
        RECT 71.900 214.900 72.300 215.000 ;
        RECT 71.900 214.600 73.800 214.900 ;
        RECT 74.200 214.800 75.400 215.100 ;
        RECT 76.600 215.100 77.000 215.200 ;
        RECT 76.600 214.800 79.100 215.100 ;
        RECT 73.400 214.500 73.800 214.600 ;
        RECT 74.300 214.200 74.600 214.800 ;
        RECT 78.700 214.700 79.100 214.800 ;
        RECT 77.900 214.200 78.300 214.300 ;
        RECT 74.300 213.900 79.800 214.200 ;
        RECT 74.500 213.800 74.900 213.900 ;
        RECT 60.600 212.800 61.500 213.100 ;
        RECT 59.000 212.100 59.400 212.200 ;
        RECT 50.200 211.800 51.200 212.100 ;
        RECT 50.800 211.100 51.200 211.800 ;
        RECT 53.000 211.100 53.400 212.100 ;
        RECT 55.000 211.800 55.700 212.100 ;
        RECT 55.100 211.100 55.700 211.800 ;
        RECT 57.400 211.800 59.400 212.100 ;
        RECT 57.400 211.100 57.800 211.800 ;
        RECT 61.100 211.100 61.500 212.800 ;
        RECT 62.200 211.100 62.600 213.100 ;
        RECT 63.000 213.000 65.000 213.100 ;
        RECT 63.000 211.100 63.400 213.000 ;
        RECT 64.600 211.100 65.000 213.000 ;
        RECT 65.400 213.000 67.400 213.100 ;
        RECT 65.400 211.100 65.800 213.000 ;
        RECT 67.000 211.100 67.400 213.000 ;
        RECT 67.800 211.100 68.200 213.100 ;
        RECT 68.900 212.800 69.800 213.100 ;
        RECT 71.000 213.300 72.900 213.600 ;
        RECT 68.900 211.100 69.300 212.800 ;
        RECT 71.000 211.100 71.400 213.300 ;
        RECT 72.500 213.200 72.900 213.300 ;
        RECT 77.400 212.800 77.700 213.900 ;
        RECT 79.000 213.800 79.800 213.900 ;
        RECT 80.600 213.600 81.000 215.300 ;
        RECT 82.300 215.200 82.700 215.300 ;
        RECT 83.900 215.200 84.200 215.800 ;
        RECT 84.900 215.900 85.200 216.500 ;
        RECT 85.500 216.500 85.900 216.600 ;
        RECT 87.800 216.500 88.200 216.600 ;
        RECT 85.500 216.200 88.200 216.500 ;
        RECT 84.900 215.700 87.300 215.900 ;
        RECT 89.400 215.700 89.800 219.900 ;
        RECT 84.900 215.600 89.800 215.700 ;
        RECT 86.900 215.500 89.800 215.600 ;
        RECT 87.000 215.400 89.800 215.500 ;
        RECT 90.200 215.700 90.600 219.900 ;
        RECT 92.400 218.200 92.800 219.900 ;
        RECT 91.800 217.900 92.800 218.200 ;
        RECT 94.600 217.900 95.000 219.900 ;
        RECT 96.700 217.900 97.300 219.900 ;
        RECT 91.800 217.500 92.200 217.900 ;
        RECT 94.600 217.600 94.900 217.900 ;
        RECT 93.500 217.300 95.300 217.600 ;
        RECT 96.600 217.500 97.000 217.900 ;
        RECT 93.500 217.200 93.900 217.300 ;
        RECT 94.900 217.200 95.300 217.300 ;
        RECT 91.800 216.500 92.200 216.600 ;
        RECT 94.100 216.500 94.500 216.600 ;
        RECT 91.800 216.200 94.500 216.500 ;
        RECT 94.800 216.500 95.900 216.800 ;
        RECT 94.800 215.900 95.100 216.500 ;
        RECT 95.500 216.400 95.900 216.500 ;
        RECT 96.700 216.600 97.400 217.000 ;
        RECT 96.700 216.100 97.000 216.600 ;
        RECT 92.700 215.700 95.100 215.900 ;
        RECT 90.200 215.600 95.100 215.700 ;
        RECT 95.800 215.800 97.000 216.100 ;
        RECT 90.200 215.500 93.100 215.600 ;
        RECT 90.200 215.400 93.000 215.500 ;
        RECT 81.500 214.900 81.900 215.000 ;
        RECT 81.500 214.600 83.400 214.900 ;
        RECT 83.800 214.800 84.200 215.200 ;
        RECT 86.200 215.100 86.600 215.200 ;
        RECT 93.400 215.100 93.800 215.200 ;
        RECT 86.200 214.800 88.700 215.100 ;
        RECT 83.000 214.500 83.400 214.600 ;
        RECT 83.900 214.200 84.200 214.800 ;
        RECT 88.300 214.700 88.700 214.800 ;
        RECT 91.300 214.800 93.800 215.100 ;
        RECT 91.300 214.700 91.700 214.800 ;
        RECT 87.500 214.200 87.900 214.300 ;
        RECT 92.100 214.200 92.500 214.300 ;
        RECT 95.800 214.200 96.100 215.800 ;
        RECT 99.000 215.600 99.400 219.900 ;
        RECT 99.800 215.900 100.200 219.900 ;
        RECT 100.600 216.200 101.000 219.900 ;
        RECT 102.200 216.200 102.600 219.900 ;
        RECT 100.600 215.900 102.600 216.200 ;
        RECT 97.300 215.300 99.400 215.600 ;
        RECT 97.300 215.200 97.700 215.300 ;
        RECT 98.100 214.900 98.500 215.000 ;
        RECT 96.600 214.600 98.500 214.900 ;
        RECT 96.600 214.500 97.000 214.600 ;
        RECT 83.900 214.100 89.400 214.200 ;
        RECT 90.600 214.100 96.100 214.200 ;
        RECT 83.900 213.900 96.100 214.100 ;
        RECT 84.100 213.800 84.500 213.900 ;
        RECT 76.500 212.700 76.900 212.800 ;
        RECT 73.400 212.100 73.800 212.500 ;
        RECT 75.500 212.400 76.900 212.700 ;
        RECT 77.400 212.400 77.800 212.800 ;
        RECT 75.500 212.100 75.800 212.400 ;
        RECT 78.200 212.100 78.600 212.500 ;
        RECT 73.100 211.800 73.800 212.100 ;
        RECT 73.100 211.100 73.700 211.800 ;
        RECT 75.400 211.100 75.800 212.100 ;
        RECT 77.600 211.800 78.600 212.100 ;
        RECT 77.600 211.100 78.000 211.800 ;
        RECT 79.800 211.100 80.200 213.500 ;
        RECT 80.600 213.300 82.500 213.600 ;
        RECT 80.600 211.100 81.000 213.300 ;
        RECT 82.100 213.200 82.500 213.300 ;
        RECT 87.000 212.800 87.300 213.900 ;
        RECT 88.600 213.800 91.400 213.900 ;
        RECT 86.100 212.700 86.500 212.800 ;
        RECT 83.000 212.100 83.400 212.500 ;
        RECT 85.100 212.400 86.500 212.700 ;
        RECT 87.000 212.400 87.400 212.800 ;
        RECT 85.100 212.100 85.400 212.400 ;
        RECT 87.800 212.100 88.200 212.500 ;
        RECT 82.700 211.800 83.400 212.100 ;
        RECT 82.700 211.100 83.300 211.800 ;
        RECT 85.000 211.100 85.400 212.100 ;
        RECT 87.200 211.800 88.200 212.100 ;
        RECT 87.200 211.100 87.600 211.800 ;
        RECT 89.400 211.100 89.800 213.500 ;
        RECT 90.200 211.100 90.600 213.500 ;
        RECT 92.700 212.800 93.000 213.900 ;
        RECT 95.500 213.800 95.900 213.900 ;
        RECT 99.000 213.600 99.400 215.300 ;
        RECT 99.900 215.200 100.200 215.900 ;
        RECT 104.600 215.600 105.000 219.900 ;
        RECT 106.700 217.900 107.300 219.900 ;
        RECT 109.000 217.900 109.400 219.900 ;
        RECT 111.200 218.200 111.600 219.900 ;
        RECT 111.200 217.900 112.200 218.200 ;
        RECT 107.000 217.500 107.400 217.900 ;
        RECT 109.100 217.600 109.400 217.900 ;
        RECT 108.700 217.300 110.500 217.600 ;
        RECT 111.800 217.500 112.200 217.900 ;
        RECT 108.700 217.200 109.100 217.300 ;
        RECT 110.100 217.200 110.500 217.300 ;
        RECT 106.600 216.600 107.300 217.000 ;
        RECT 107.000 216.100 107.300 216.600 ;
        RECT 108.100 216.500 109.200 216.800 ;
        RECT 108.100 216.400 108.500 216.500 ;
        RECT 107.000 215.800 108.200 216.100 ;
        RECT 101.800 215.200 102.200 215.400 ;
        RECT 104.600 215.300 106.700 215.600 ;
        RECT 99.800 214.900 101.000 215.200 ;
        RECT 101.800 214.900 102.600 215.200 ;
        RECT 99.800 214.800 100.200 214.900 ;
        RECT 99.800 214.100 100.200 214.200 ;
        RECT 100.700 214.100 101.000 214.900 ;
        RECT 102.200 214.800 102.600 214.900 ;
        RECT 99.800 213.800 101.000 214.100 ;
        RECT 101.400 213.800 101.800 214.600 ;
        RECT 97.500 213.300 99.400 213.600 ;
        RECT 97.500 213.200 97.900 213.300 ;
        RECT 91.800 212.100 92.200 212.500 ;
        RECT 92.600 212.400 93.000 212.800 ;
        RECT 93.500 212.700 93.900 212.800 ;
        RECT 93.500 212.400 94.900 212.700 ;
        RECT 94.600 212.100 94.900 212.400 ;
        RECT 96.600 212.100 97.000 212.500 ;
        RECT 91.800 211.800 92.800 212.100 ;
        RECT 92.400 211.100 92.800 211.800 ;
        RECT 94.600 211.100 95.000 212.100 ;
        RECT 96.600 211.800 97.300 212.100 ;
        RECT 96.700 211.100 97.300 211.800 ;
        RECT 99.000 211.100 99.400 213.300 ;
        RECT 99.800 212.800 100.200 213.200 ;
        RECT 100.700 213.100 101.000 213.800 ;
        RECT 99.900 212.400 100.300 212.800 ;
        RECT 100.600 211.100 101.000 213.100 ;
        RECT 104.600 213.600 105.000 215.300 ;
        RECT 106.300 215.200 106.700 215.300 ;
        RECT 107.900 215.200 108.200 215.800 ;
        RECT 108.900 215.900 109.200 216.500 ;
        RECT 109.500 216.500 109.900 216.600 ;
        RECT 111.800 216.500 112.200 216.600 ;
        RECT 109.500 216.200 112.200 216.500 ;
        RECT 108.900 215.700 111.300 215.900 ;
        RECT 113.400 215.700 113.800 219.900 ;
        RECT 108.900 215.600 113.800 215.700 ;
        RECT 110.900 215.500 113.800 215.600 ;
        RECT 111.000 215.400 113.800 215.500 ;
        RECT 105.500 214.900 105.900 215.000 ;
        RECT 105.500 214.600 107.400 214.900 ;
        RECT 107.800 214.800 108.200 215.200 ;
        RECT 110.200 215.100 110.600 215.200 ;
        RECT 110.200 214.800 112.700 215.100 ;
        RECT 107.000 214.500 107.400 214.600 ;
        RECT 107.900 214.200 108.200 214.800 ;
        RECT 111.000 214.700 111.400 214.800 ;
        RECT 112.300 214.700 112.700 214.800 ;
        RECT 111.500 214.200 111.900 214.300 ;
        RECT 107.900 213.900 113.400 214.200 ;
        RECT 108.100 213.800 108.500 213.900 ;
        RECT 104.600 213.300 106.500 213.600 ;
        RECT 104.600 211.100 105.000 213.300 ;
        RECT 106.100 213.200 106.500 213.300 ;
        RECT 111.000 212.800 111.300 213.900 ;
        RECT 112.600 213.800 113.400 213.900 ;
        RECT 114.200 213.800 114.600 214.200 ;
        RECT 110.100 212.700 110.500 212.800 ;
        RECT 107.000 212.100 107.400 212.500 ;
        RECT 109.100 212.400 110.500 212.700 ;
        RECT 111.000 212.400 111.400 212.800 ;
        RECT 109.100 212.100 109.400 212.400 ;
        RECT 111.800 212.100 112.200 212.500 ;
        RECT 106.700 211.800 107.400 212.100 ;
        RECT 106.700 211.100 107.300 211.800 ;
        RECT 109.000 211.100 109.400 212.100 ;
        RECT 111.200 211.800 112.200 212.100 ;
        RECT 111.200 211.100 111.600 211.800 ;
        RECT 113.400 211.100 113.800 213.500 ;
        RECT 114.200 213.200 114.500 213.800 ;
        RECT 114.200 212.400 114.600 213.200 ;
        RECT 115.000 211.100 115.400 219.900 ;
        RECT 117.100 216.300 117.500 219.900 ;
        RECT 116.600 215.900 117.500 216.300 ;
        RECT 118.200 215.900 118.600 219.900 ;
        RECT 119.000 216.200 119.400 219.900 ;
        RECT 120.600 216.200 121.000 219.900 ;
        RECT 119.000 215.900 121.000 216.200 ;
        RECT 116.700 214.200 117.000 215.900 ;
        RECT 117.400 214.800 117.800 215.600 ;
        RECT 118.300 215.200 118.600 215.900 ;
        RECT 121.400 215.600 121.800 219.900 ;
        RECT 123.500 217.900 124.100 219.900 ;
        RECT 125.800 217.900 126.200 219.900 ;
        RECT 128.000 218.200 128.400 219.900 ;
        RECT 128.000 217.900 129.000 218.200 ;
        RECT 123.800 217.500 124.200 217.900 ;
        RECT 125.900 217.600 126.200 217.900 ;
        RECT 125.500 217.300 127.300 217.600 ;
        RECT 128.600 217.500 129.000 217.900 ;
        RECT 125.500 217.200 125.900 217.300 ;
        RECT 126.900 217.200 127.300 217.300 ;
        RECT 123.400 216.600 124.100 217.000 ;
        RECT 123.800 216.100 124.100 216.600 ;
        RECT 124.900 216.500 126.000 216.800 ;
        RECT 124.900 216.400 125.300 216.500 ;
        RECT 123.800 215.800 125.000 216.100 ;
        RECT 120.200 215.200 120.600 215.400 ;
        RECT 121.400 215.300 123.500 215.600 ;
        RECT 118.200 214.900 119.400 215.200 ;
        RECT 120.200 214.900 121.000 215.200 ;
        RECT 118.200 214.800 118.600 214.900 ;
        RECT 116.600 213.800 117.000 214.200 ;
        RECT 118.200 214.100 118.600 214.200 ;
        RECT 119.100 214.100 119.400 214.900 ;
        RECT 120.600 214.800 121.000 214.900 ;
        RECT 118.200 213.800 119.400 214.100 ;
        RECT 119.800 213.800 120.200 214.600 ;
        RECT 115.800 212.400 116.200 213.200 ;
        RECT 116.700 213.100 117.000 213.800 ;
        RECT 118.200 213.100 118.600 213.200 ;
        RECT 119.100 213.100 119.400 213.800 ;
        RECT 116.600 212.800 118.600 213.100 ;
        RECT 116.700 212.100 117.000 212.800 ;
        RECT 118.300 212.400 118.700 212.800 ;
        RECT 116.600 211.100 117.000 212.100 ;
        RECT 119.000 211.100 119.400 213.100 ;
        RECT 121.400 213.600 121.800 215.300 ;
        RECT 123.100 215.200 123.500 215.300 ;
        RECT 122.300 214.900 122.700 215.000 ;
        RECT 122.300 214.600 124.200 214.900 ;
        RECT 123.800 214.500 124.200 214.600 ;
        RECT 124.700 214.200 125.000 215.800 ;
        RECT 125.700 215.900 126.000 216.500 ;
        RECT 126.300 216.500 126.700 216.600 ;
        RECT 128.600 216.500 129.000 216.600 ;
        RECT 126.300 216.200 129.000 216.500 ;
        RECT 125.700 215.700 128.100 215.900 ;
        RECT 130.200 215.700 130.600 219.900 ;
        RECT 132.900 216.400 133.300 219.900 ;
        RECT 135.000 217.500 135.400 219.500 ;
        RECT 125.700 215.600 130.600 215.700 ;
        RECT 132.500 216.100 133.300 216.400 ;
        RECT 127.700 215.500 130.600 215.600 ;
        RECT 127.800 215.400 130.600 215.500 ;
        RECT 127.000 215.100 127.400 215.200 ;
        RECT 127.000 214.800 129.500 215.100 ;
        RECT 131.800 214.800 132.200 215.600 ;
        RECT 129.100 214.700 129.500 214.800 ;
        RECT 128.300 214.200 128.700 214.300 ;
        RECT 132.500 214.200 132.800 216.100 ;
        RECT 135.100 215.800 135.400 217.500 ;
        RECT 136.600 216.400 137.000 219.900 ;
        RECT 133.500 215.500 135.400 215.800 ;
        RECT 136.500 215.900 137.000 216.400 ;
        RECT 138.200 216.200 138.600 219.900 ;
        RECT 137.300 215.900 138.600 216.200 ;
        RECT 139.000 216.200 139.400 219.900 ;
        RECT 140.600 216.400 141.000 219.900 ;
        RECT 139.000 215.900 140.300 216.200 ;
        RECT 140.600 215.900 141.100 216.400 ;
        RECT 133.500 214.500 133.800 215.500 ;
        RECT 124.700 213.900 130.200 214.200 ;
        RECT 124.900 213.800 125.300 213.900 ;
        RECT 121.400 213.300 123.300 213.600 ;
        RECT 121.400 211.100 121.800 213.300 ;
        RECT 122.900 213.200 123.300 213.300 ;
        RECT 127.800 212.800 128.100 213.900 ;
        RECT 129.400 213.800 130.200 213.900 ;
        RECT 131.800 213.800 132.800 214.200 ;
        RECT 133.100 214.100 133.800 214.500 ;
        RECT 134.200 214.400 134.600 215.200 ;
        RECT 135.000 214.400 135.400 215.200 ;
        RECT 132.500 213.500 132.800 213.800 ;
        RECT 133.300 213.900 133.800 214.100 ;
        RECT 136.500 214.200 136.800 215.900 ;
        RECT 137.300 214.900 137.600 215.900 ;
        RECT 137.100 214.500 137.600 214.900 ;
        RECT 133.300 213.600 135.400 213.900 ;
        RECT 126.900 212.700 127.300 212.800 ;
        RECT 123.800 212.100 124.200 212.500 ;
        RECT 125.900 212.400 127.300 212.700 ;
        RECT 127.800 212.400 128.200 212.800 ;
        RECT 125.900 212.100 126.200 212.400 ;
        RECT 128.600 212.100 129.000 212.500 ;
        RECT 123.500 211.800 124.200 212.100 ;
        RECT 123.500 211.100 124.100 211.800 ;
        RECT 125.800 211.100 126.200 212.100 ;
        RECT 128.000 211.800 129.000 212.100 ;
        RECT 128.000 211.100 128.400 211.800 ;
        RECT 130.200 211.100 130.600 213.500 ;
        RECT 132.500 213.300 132.900 213.500 ;
        RECT 132.500 213.000 133.300 213.300 ;
        RECT 132.900 212.200 133.300 213.000 ;
        RECT 135.100 212.500 135.400 213.600 ;
        RECT 136.500 213.800 137.000 214.200 ;
        RECT 136.500 213.100 136.800 213.800 ;
        RECT 137.300 213.700 137.600 214.500 ;
        RECT 138.100 215.100 138.600 215.200 ;
        RECT 139.000 215.100 139.500 215.200 ;
        RECT 138.100 214.800 139.500 215.100 ;
        RECT 138.100 214.400 138.500 214.800 ;
        RECT 139.100 214.400 139.500 214.800 ;
        RECT 140.000 214.900 140.300 215.900 ;
        RECT 140.000 214.500 140.500 214.900 ;
        RECT 140.000 213.700 140.300 214.500 ;
        RECT 140.800 214.200 141.100 215.900 ;
        RECT 143.000 215.600 143.400 219.900 ;
        RECT 144.600 215.600 145.000 219.900 ;
        RECT 146.200 215.600 146.600 219.900 ;
        RECT 147.800 215.600 148.200 219.900 ;
        RECT 140.600 213.800 141.100 214.200 ;
        RECT 137.300 213.400 138.600 213.700 ;
        RECT 136.500 212.800 137.000 213.100 ;
        RECT 132.600 211.800 133.300 212.200 ;
        RECT 132.900 211.500 133.300 211.800 ;
        RECT 135.000 211.500 135.400 212.500 ;
        RECT 136.600 211.100 137.000 212.800 ;
        RECT 138.200 211.100 138.600 213.400 ;
        RECT 139.000 213.400 140.300 213.700 ;
        RECT 139.000 211.100 139.400 213.400 ;
        RECT 140.800 213.100 141.100 213.800 ;
        RECT 142.200 215.200 143.400 215.600 ;
        RECT 143.900 215.200 145.000 215.600 ;
        RECT 145.500 215.200 146.600 215.600 ;
        RECT 147.300 215.200 148.200 215.600 ;
        RECT 149.400 215.600 149.800 219.900 ;
        RECT 151.500 217.900 152.100 219.900 ;
        RECT 153.800 217.900 154.200 219.900 ;
        RECT 156.000 218.200 156.400 219.900 ;
        RECT 156.000 217.900 157.000 218.200 ;
        RECT 151.800 217.500 152.200 217.900 ;
        RECT 153.900 217.600 154.200 217.900 ;
        RECT 153.500 217.300 155.300 217.600 ;
        RECT 156.600 217.500 157.000 217.900 ;
        RECT 153.500 217.200 153.900 217.300 ;
        RECT 154.900 217.200 155.300 217.300 ;
        RECT 151.400 216.600 152.100 217.000 ;
        RECT 151.800 216.100 152.100 216.600 ;
        RECT 152.900 216.500 154.000 216.800 ;
        RECT 152.900 216.400 153.300 216.500 ;
        RECT 151.800 215.800 153.000 216.100 ;
        RECT 149.400 215.300 151.500 215.600 ;
        RECT 142.200 213.800 142.600 215.200 ;
        RECT 143.900 214.500 144.300 215.200 ;
        RECT 145.500 214.500 145.900 215.200 ;
        RECT 147.300 214.500 147.700 215.200 ;
        RECT 143.000 214.100 144.300 214.500 ;
        RECT 144.700 214.100 145.900 214.500 ;
        RECT 146.400 214.100 147.700 214.500 ;
        RECT 148.100 214.100 149.000 214.500 ;
        RECT 143.900 213.800 144.300 214.100 ;
        RECT 145.500 213.800 145.900 214.100 ;
        RECT 147.300 213.800 147.700 214.100 ;
        RECT 148.600 213.800 149.000 214.100 ;
        RECT 142.200 213.400 143.400 213.800 ;
        RECT 143.900 213.400 145.000 213.800 ;
        RECT 145.500 213.400 146.600 213.800 ;
        RECT 147.300 213.400 148.200 213.800 ;
        RECT 140.600 212.800 141.100 213.100 ;
        RECT 140.600 211.100 141.000 212.800 ;
        RECT 143.000 211.100 143.400 213.400 ;
        RECT 144.600 211.100 145.000 213.400 ;
        RECT 146.200 211.100 146.600 213.400 ;
        RECT 147.800 211.100 148.200 213.400 ;
        RECT 149.400 213.600 149.800 215.300 ;
        RECT 151.100 215.200 151.500 215.300 ;
        RECT 152.700 215.200 153.000 215.800 ;
        RECT 153.700 215.900 154.000 216.500 ;
        RECT 154.300 216.500 154.700 216.600 ;
        RECT 156.600 216.500 157.000 216.600 ;
        RECT 154.300 216.200 157.000 216.500 ;
        RECT 153.700 215.700 156.100 215.900 ;
        RECT 158.200 215.700 158.600 219.900 ;
        RECT 153.700 215.600 158.600 215.700 ;
        RECT 161.400 215.600 161.800 219.900 ;
        RECT 163.000 215.600 163.400 219.900 ;
        RECT 164.600 215.600 165.000 219.900 ;
        RECT 166.200 215.600 166.600 219.900 ;
        RECT 155.700 215.500 158.600 215.600 ;
        RECT 155.800 215.400 158.600 215.500 ;
        RECT 160.600 215.200 161.800 215.600 ;
        RECT 162.300 215.200 163.400 215.600 ;
        RECT 163.900 215.200 165.000 215.600 ;
        RECT 165.700 215.200 166.600 215.600 ;
        RECT 167.800 215.600 168.200 219.900 ;
        RECT 169.900 217.900 170.500 219.900 ;
        RECT 172.200 217.900 172.600 219.900 ;
        RECT 174.400 218.200 174.800 219.900 ;
        RECT 174.400 217.900 175.400 218.200 ;
        RECT 170.200 217.500 170.600 217.900 ;
        RECT 172.300 217.600 172.600 217.900 ;
        RECT 171.900 217.300 173.700 217.600 ;
        RECT 175.000 217.500 175.400 217.900 ;
        RECT 171.900 217.200 172.300 217.300 ;
        RECT 173.300 217.200 173.700 217.300 ;
        RECT 169.800 216.600 170.500 217.000 ;
        RECT 170.200 216.100 170.500 216.600 ;
        RECT 171.300 216.500 172.400 216.800 ;
        RECT 171.300 216.400 171.700 216.500 ;
        RECT 170.200 215.800 171.400 216.100 ;
        RECT 167.800 215.300 169.900 215.600 ;
        RECT 150.300 214.900 150.700 215.000 ;
        RECT 150.300 214.600 152.200 214.900 ;
        RECT 152.600 214.800 153.000 215.200 ;
        RECT 155.000 215.100 155.400 215.200 ;
        RECT 155.000 214.800 157.500 215.100 ;
        RECT 151.800 214.500 152.200 214.600 ;
        RECT 152.700 214.200 153.000 214.800 ;
        RECT 157.100 214.700 157.500 214.800 ;
        RECT 156.300 214.200 156.700 214.300 ;
        RECT 152.700 213.900 158.200 214.200 ;
        RECT 152.900 213.800 153.300 213.900 ;
        RECT 149.400 213.300 151.300 213.600 ;
        RECT 149.400 211.100 149.800 213.300 ;
        RECT 150.900 213.200 151.300 213.300 ;
        RECT 155.800 212.800 156.100 213.900 ;
        RECT 157.400 213.800 158.200 213.900 ;
        RECT 160.600 213.800 161.000 215.200 ;
        RECT 162.300 214.500 162.700 215.200 ;
        RECT 163.900 214.500 164.300 215.200 ;
        RECT 165.700 214.500 166.100 215.200 ;
        RECT 161.400 214.100 162.700 214.500 ;
        RECT 163.100 214.100 164.300 214.500 ;
        RECT 164.800 214.100 166.100 214.500 ;
        RECT 162.300 213.800 162.700 214.100 ;
        RECT 163.900 213.800 164.300 214.100 ;
        RECT 165.700 213.800 166.100 214.100 ;
        RECT 154.900 212.700 155.300 212.800 ;
        RECT 151.800 212.100 152.200 212.500 ;
        RECT 153.900 212.400 155.300 212.700 ;
        RECT 155.800 212.400 156.200 212.800 ;
        RECT 153.900 212.100 154.200 212.400 ;
        RECT 156.600 212.100 157.000 212.500 ;
        RECT 151.500 211.800 152.200 212.100 ;
        RECT 151.500 211.100 152.100 211.800 ;
        RECT 153.800 211.100 154.200 212.100 ;
        RECT 156.000 211.800 157.000 212.100 ;
        RECT 156.000 211.100 156.400 211.800 ;
        RECT 158.200 211.100 158.600 213.500 ;
        RECT 160.600 213.400 161.800 213.800 ;
        RECT 162.300 213.400 163.400 213.800 ;
        RECT 163.900 213.400 165.000 213.800 ;
        RECT 165.700 213.400 166.600 213.800 ;
        RECT 161.400 211.100 161.800 213.400 ;
        RECT 163.000 211.100 163.400 213.400 ;
        RECT 164.600 211.100 165.000 213.400 ;
        RECT 166.200 211.100 166.600 213.400 ;
        RECT 167.800 213.600 168.200 215.300 ;
        RECT 169.500 215.200 169.900 215.300 ;
        RECT 168.700 214.900 169.100 215.000 ;
        RECT 168.700 214.600 170.600 214.900 ;
        RECT 170.200 214.500 170.600 214.600 ;
        RECT 171.100 214.200 171.400 215.800 ;
        RECT 172.100 215.900 172.400 216.500 ;
        RECT 172.700 216.500 173.100 216.600 ;
        RECT 175.000 216.500 175.400 216.600 ;
        RECT 172.700 216.200 175.400 216.500 ;
        RECT 172.100 215.700 174.500 215.900 ;
        RECT 176.600 215.700 177.000 219.900 ;
        RECT 172.100 215.600 177.000 215.700 ;
        RECT 174.100 215.500 177.000 215.600 ;
        RECT 174.200 215.400 177.000 215.500 ;
        RECT 173.400 215.100 173.800 215.200 ;
        RECT 178.200 215.100 178.600 219.900 ;
        RECT 180.200 216.800 180.600 217.200 ;
        RECT 179.000 215.800 179.400 216.600 ;
        RECT 180.200 216.200 180.500 216.800 ;
        RECT 180.900 216.200 181.300 219.900 ;
        RECT 184.100 219.200 184.500 219.900 ;
        RECT 184.100 218.800 185.000 219.200 ;
        RECT 183.400 216.800 183.800 217.200 ;
        RECT 183.400 216.200 183.700 216.800 ;
        RECT 184.100 216.200 184.500 218.800 ;
        RECT 179.800 215.900 180.500 216.200 ;
        RECT 180.800 215.900 181.300 216.200 ;
        RECT 183.000 215.900 183.700 216.200 ;
        RECT 184.000 215.900 184.500 216.200 ;
        RECT 179.800 215.800 180.200 215.900 ;
        RECT 179.800 215.100 180.100 215.800 ;
        RECT 173.400 214.800 175.900 215.100 ;
        RECT 174.200 214.700 174.600 214.800 ;
        RECT 175.500 214.700 175.900 214.800 ;
        RECT 178.200 214.800 180.100 215.100 ;
        RECT 174.700 214.200 175.100 214.300 ;
        RECT 171.100 213.900 176.600 214.200 ;
        RECT 171.300 213.800 172.200 213.900 ;
        RECT 167.800 213.300 169.700 213.600 ;
        RECT 167.800 211.100 168.200 213.300 ;
        RECT 169.300 213.200 169.700 213.300 ;
        RECT 174.200 212.800 174.500 213.900 ;
        RECT 175.800 213.800 176.600 213.900 ;
        RECT 173.300 212.700 173.700 212.800 ;
        RECT 170.200 212.100 170.600 212.500 ;
        RECT 172.300 212.400 173.700 212.700 ;
        RECT 174.200 212.400 174.600 212.800 ;
        RECT 172.300 212.100 172.600 212.400 ;
        RECT 175.000 212.100 175.400 212.500 ;
        RECT 169.900 211.800 170.600 212.100 ;
        RECT 169.900 211.100 170.500 211.800 ;
        RECT 172.200 211.100 172.600 212.100 ;
        RECT 174.400 211.800 175.400 212.100 ;
        RECT 174.400 211.100 174.800 211.800 ;
        RECT 176.600 211.100 177.000 213.500 ;
        RECT 177.400 213.400 177.800 214.200 ;
        RECT 178.200 213.100 178.600 214.800 ;
        RECT 180.800 214.200 181.100 215.900 ;
        RECT 183.000 215.800 183.400 215.900 ;
        RECT 181.400 214.400 181.800 215.200 ;
        RECT 184.000 214.200 184.300 215.900 ;
        RECT 187.000 215.600 187.400 219.900 ;
        RECT 188.600 215.600 189.000 219.900 ;
        RECT 190.200 215.600 190.600 219.900 ;
        RECT 191.800 215.600 192.200 219.900 ;
        RECT 194.700 216.200 195.100 219.900 ;
        RECT 195.400 216.800 195.800 217.200 ;
        RECT 195.500 216.200 195.800 216.800 ;
        RECT 194.700 215.900 195.200 216.200 ;
        RECT 195.500 215.900 196.200 216.200 ;
        RECT 186.200 215.200 187.400 215.600 ;
        RECT 187.900 215.200 189.000 215.600 ;
        RECT 189.500 215.200 190.600 215.600 ;
        RECT 191.300 215.200 192.200 215.600 ;
        RECT 184.600 214.400 185.000 215.200 ;
        RECT 179.000 214.100 179.400 214.200 ;
        RECT 179.800 214.100 181.100 214.200 ;
        RECT 182.200 214.100 182.600 214.200 ;
        RECT 179.000 213.800 181.100 214.100 ;
        RECT 181.800 213.800 182.600 214.100 ;
        RECT 183.000 213.800 184.300 214.200 ;
        RECT 185.400 214.100 185.800 214.200 ;
        RECT 185.000 213.800 185.800 214.100 ;
        RECT 186.200 213.800 186.600 215.200 ;
        RECT 187.900 214.500 188.300 215.200 ;
        RECT 189.500 214.500 189.900 215.200 ;
        RECT 191.300 214.500 191.700 215.200 ;
        RECT 187.000 214.100 188.300 214.500 ;
        RECT 188.700 214.100 189.900 214.500 ;
        RECT 190.400 214.100 191.700 214.500 ;
        RECT 192.100 214.100 193.000 214.500 ;
        RECT 194.200 214.400 194.600 215.200 ;
        RECT 194.900 214.200 195.200 215.900 ;
        RECT 195.800 215.800 196.200 215.900 ;
        RECT 196.600 215.800 197.000 216.600 ;
        RECT 195.800 215.100 196.100 215.800 ;
        RECT 197.400 215.100 197.800 219.900 ;
        RECT 195.800 214.800 197.800 215.100 ;
        RECT 187.900 213.800 188.300 214.100 ;
        RECT 189.500 213.800 189.900 214.100 ;
        RECT 191.300 213.800 191.700 214.100 ;
        RECT 192.600 213.800 193.000 214.100 ;
        RECT 193.400 214.100 193.800 214.200 ;
        RECT 193.400 213.800 194.200 214.100 ;
        RECT 194.900 213.800 196.200 214.200 ;
        RECT 179.900 213.100 180.200 213.800 ;
        RECT 181.800 213.600 182.200 213.800 ;
        RECT 180.700 213.100 182.500 213.300 ;
        RECT 183.100 213.100 183.400 213.800 ;
        RECT 185.000 213.600 185.400 213.800 ;
        RECT 186.200 213.400 187.400 213.800 ;
        RECT 187.900 213.400 189.000 213.800 ;
        RECT 189.500 213.400 190.600 213.800 ;
        RECT 191.300 213.400 192.200 213.800 ;
        RECT 193.800 213.600 194.200 213.800 ;
        RECT 183.900 213.100 185.700 213.300 ;
        RECT 178.200 212.800 179.100 213.100 ;
        RECT 178.700 211.100 179.100 212.800 ;
        RECT 179.800 211.100 180.200 213.100 ;
        RECT 180.600 213.000 182.600 213.100 ;
        RECT 180.600 211.100 181.000 213.000 ;
        RECT 182.200 211.100 182.600 213.000 ;
        RECT 183.000 211.100 183.400 213.100 ;
        RECT 183.800 213.000 185.800 213.100 ;
        RECT 183.800 211.100 184.200 213.000 ;
        RECT 185.400 211.100 185.800 213.000 ;
        RECT 187.000 211.100 187.400 213.400 ;
        RECT 188.600 211.100 189.000 213.400 ;
        RECT 190.200 211.100 190.600 213.400 ;
        RECT 191.800 211.100 192.200 213.400 ;
        RECT 193.500 213.100 195.300 213.300 ;
        RECT 195.800 213.100 196.100 213.800 ;
        RECT 197.400 213.100 197.800 214.800 ;
        RECT 199.000 215.600 199.400 219.900 ;
        RECT 201.100 217.900 201.700 219.900 ;
        RECT 203.400 217.900 203.800 219.900 ;
        RECT 205.600 218.200 206.000 219.900 ;
        RECT 205.600 217.900 206.600 218.200 ;
        RECT 201.400 217.500 201.800 217.900 ;
        RECT 203.500 217.600 203.800 217.900 ;
        RECT 203.100 217.300 204.900 217.600 ;
        RECT 206.200 217.500 206.600 217.900 ;
        RECT 203.100 217.200 203.500 217.300 ;
        RECT 204.500 217.200 204.900 217.300 ;
        RECT 201.000 216.600 201.700 217.000 ;
        RECT 201.400 216.100 201.700 216.600 ;
        RECT 202.500 216.500 203.600 216.800 ;
        RECT 202.500 216.400 202.900 216.500 ;
        RECT 201.400 215.800 202.600 216.100 ;
        RECT 199.000 215.300 201.100 215.600 ;
        RECT 198.200 213.400 198.600 214.200 ;
        RECT 199.000 213.600 199.400 215.300 ;
        RECT 200.700 215.200 201.100 215.300 ;
        RECT 199.900 214.900 200.300 215.000 ;
        RECT 199.900 214.600 201.800 214.900 ;
        RECT 201.400 214.500 201.800 214.600 ;
        RECT 202.300 214.200 202.600 215.800 ;
        RECT 203.300 215.900 203.600 216.500 ;
        RECT 203.900 216.500 204.300 216.600 ;
        RECT 206.200 216.500 206.600 216.600 ;
        RECT 203.900 216.200 206.600 216.500 ;
        RECT 203.300 215.700 205.700 215.900 ;
        RECT 207.800 215.700 208.200 219.900 ;
        RECT 203.300 215.600 208.200 215.700 ;
        RECT 205.300 215.500 208.200 215.600 ;
        RECT 205.400 215.400 208.200 215.500 ;
        RECT 210.200 215.700 210.600 219.900 ;
        RECT 212.400 218.200 212.800 219.900 ;
        RECT 211.800 217.900 212.800 218.200 ;
        RECT 214.600 217.900 215.000 219.900 ;
        RECT 216.700 217.900 217.300 219.900 ;
        RECT 211.800 217.500 212.200 217.900 ;
        RECT 214.600 217.600 214.900 217.900 ;
        RECT 213.500 217.300 215.300 217.600 ;
        RECT 216.600 217.500 217.000 217.900 ;
        RECT 213.500 217.200 213.900 217.300 ;
        RECT 214.900 217.200 215.300 217.300 ;
        RECT 211.800 216.500 212.200 216.600 ;
        RECT 214.100 216.500 214.500 216.600 ;
        RECT 211.800 216.200 214.500 216.500 ;
        RECT 214.800 216.500 215.900 216.800 ;
        RECT 214.800 215.900 215.100 216.500 ;
        RECT 215.500 216.400 215.900 216.500 ;
        RECT 216.700 216.600 217.400 217.000 ;
        RECT 216.700 216.100 217.000 216.600 ;
        RECT 212.700 215.700 215.100 215.900 ;
        RECT 210.200 215.600 215.100 215.700 ;
        RECT 215.800 215.800 217.000 216.100 ;
        RECT 210.200 215.500 213.100 215.600 ;
        RECT 210.200 215.400 213.000 215.500 ;
        RECT 203.000 215.100 203.400 215.200 ;
        RECT 204.600 215.100 205.000 215.200 ;
        RECT 213.400 215.100 213.800 215.200 ;
        RECT 203.000 214.800 207.100 215.100 ;
        RECT 206.700 214.700 207.100 214.800 ;
        RECT 211.300 214.800 213.800 215.100 ;
        RECT 215.000 215.100 215.400 215.200 ;
        RECT 215.800 215.100 216.100 215.800 ;
        RECT 219.000 215.600 219.400 219.900 ;
        RECT 219.800 216.200 220.200 219.900 ;
        RECT 221.400 216.400 221.800 219.900 ;
        RECT 223.800 216.400 224.200 219.900 ;
        RECT 219.800 215.900 221.100 216.200 ;
        RECT 221.400 215.900 221.900 216.400 ;
        RECT 217.300 215.300 219.400 215.600 ;
        RECT 217.300 215.200 217.700 215.300 ;
        RECT 215.000 214.800 216.100 215.100 ;
        RECT 218.100 214.900 218.500 215.000 ;
        RECT 211.300 214.700 211.700 214.800 ;
        RECT 212.600 214.700 213.000 214.800 ;
        RECT 205.900 214.200 206.300 214.300 ;
        RECT 212.100 214.200 212.500 214.300 ;
        RECT 215.800 214.200 216.100 214.800 ;
        RECT 216.600 214.600 218.500 214.900 ;
        RECT 216.600 214.500 217.000 214.600 ;
        RECT 202.300 213.900 207.800 214.200 ;
        RECT 202.500 213.800 202.900 213.900 ;
        RECT 203.800 213.800 204.200 213.900 ;
        RECT 193.400 213.000 195.400 213.100 ;
        RECT 193.400 211.100 193.800 213.000 ;
        RECT 195.000 211.100 195.400 213.000 ;
        RECT 195.800 211.100 196.200 213.100 ;
        RECT 196.900 212.800 197.800 213.100 ;
        RECT 199.000 213.300 200.900 213.600 ;
        RECT 196.900 211.100 197.300 212.800 ;
        RECT 199.000 211.100 199.400 213.300 ;
        RECT 200.500 213.200 200.900 213.300 ;
        RECT 205.400 212.800 205.700 213.900 ;
        RECT 207.000 213.800 207.800 213.900 ;
        RECT 208.600 214.100 209.000 214.200 ;
        RECT 210.600 214.100 216.100 214.200 ;
        RECT 208.600 213.900 216.100 214.100 ;
        RECT 208.600 213.800 211.400 213.900 ;
        RECT 204.500 212.700 204.900 212.800 ;
        RECT 201.400 212.100 201.800 212.500 ;
        RECT 203.500 212.400 204.900 212.700 ;
        RECT 205.400 212.400 205.800 212.800 ;
        RECT 203.500 212.100 203.800 212.400 ;
        RECT 206.200 212.100 206.600 212.500 ;
        RECT 201.100 211.800 201.800 212.100 ;
        RECT 201.100 211.100 201.700 211.800 ;
        RECT 203.400 211.100 203.800 212.100 ;
        RECT 205.600 211.800 206.600 212.100 ;
        RECT 205.600 211.100 206.000 211.800 ;
        RECT 207.800 211.100 208.200 213.500 ;
        RECT 210.200 211.100 210.600 213.500 ;
        RECT 212.700 212.800 213.000 213.900 ;
        RECT 215.500 213.800 215.900 213.900 ;
        RECT 219.000 213.600 219.400 215.300 ;
        RECT 219.800 214.800 220.300 215.200 ;
        RECT 219.900 214.400 220.300 214.800 ;
        RECT 220.800 214.900 221.100 215.900 ;
        RECT 220.800 214.500 221.300 214.900 ;
        RECT 220.800 213.700 221.100 214.500 ;
        RECT 221.600 214.200 221.900 215.900 ;
        RECT 221.400 213.800 221.900 214.200 ;
        RECT 217.500 213.300 219.400 213.600 ;
        RECT 217.500 213.200 217.900 213.300 ;
        RECT 211.800 212.100 212.200 212.500 ;
        RECT 212.600 212.400 213.000 212.800 ;
        RECT 213.500 212.700 213.900 212.800 ;
        RECT 213.500 212.400 214.900 212.700 ;
        RECT 214.600 212.100 214.900 212.400 ;
        RECT 216.600 212.100 217.000 212.500 ;
        RECT 211.800 211.800 212.800 212.100 ;
        RECT 212.400 211.100 212.800 211.800 ;
        RECT 214.600 211.100 215.000 212.100 ;
        RECT 216.600 211.800 217.300 212.100 ;
        RECT 216.700 211.100 217.300 211.800 ;
        RECT 219.000 211.100 219.400 213.300 ;
        RECT 219.800 213.400 221.100 213.700 ;
        RECT 219.800 211.100 220.200 213.400 ;
        RECT 221.600 213.100 221.900 213.800 ;
        RECT 221.400 212.800 221.900 213.100 ;
        RECT 223.700 215.900 224.200 216.400 ;
        RECT 225.400 216.200 225.800 219.900 ;
        RECT 224.500 215.900 225.800 216.200 ;
        RECT 223.700 214.200 224.000 215.900 ;
        RECT 224.500 214.900 224.800 215.900 ;
        RECT 226.200 215.600 226.600 219.900 ;
        RECT 228.300 217.900 228.900 219.900 ;
        RECT 230.600 217.900 231.000 219.900 ;
        RECT 232.800 218.200 233.200 219.900 ;
        RECT 232.800 217.900 233.800 218.200 ;
        RECT 228.600 217.500 229.000 217.900 ;
        RECT 230.700 217.600 231.000 217.900 ;
        RECT 230.300 217.300 232.100 217.600 ;
        RECT 233.400 217.500 233.800 217.900 ;
        RECT 230.300 217.200 230.700 217.300 ;
        RECT 231.700 217.200 232.100 217.300 ;
        RECT 228.200 216.600 228.900 217.000 ;
        RECT 228.600 216.100 228.900 216.600 ;
        RECT 229.700 216.500 230.800 216.800 ;
        RECT 229.700 216.400 230.100 216.500 ;
        RECT 228.600 215.800 229.800 216.100 ;
        RECT 226.200 215.300 228.300 215.600 ;
        RECT 224.300 214.500 224.800 214.900 ;
        RECT 223.700 213.800 224.200 214.200 ;
        RECT 223.700 213.100 224.000 213.800 ;
        RECT 224.500 213.700 224.800 214.500 ;
        RECT 225.300 214.800 225.800 215.200 ;
        RECT 225.300 214.400 225.700 214.800 ;
        RECT 224.500 213.400 225.800 213.700 ;
        RECT 223.700 212.800 224.200 213.100 ;
        RECT 221.400 211.100 221.800 212.800 ;
        RECT 223.800 211.100 224.200 212.800 ;
        RECT 225.400 211.100 225.800 213.400 ;
        RECT 226.200 213.600 226.600 215.300 ;
        RECT 227.900 215.200 228.300 215.300 ;
        RECT 227.100 214.900 227.500 215.000 ;
        RECT 227.100 214.600 229.000 214.900 ;
        RECT 228.600 214.500 229.000 214.600 ;
        RECT 229.500 214.200 229.800 215.800 ;
        RECT 230.500 215.900 230.800 216.500 ;
        RECT 231.100 216.500 231.500 216.600 ;
        RECT 233.400 216.500 233.800 216.600 ;
        RECT 231.100 216.200 233.800 216.500 ;
        RECT 230.500 215.700 232.900 215.900 ;
        RECT 235.000 215.700 235.400 219.900 ;
        RECT 230.500 215.600 235.400 215.700 ;
        RECT 232.500 215.500 235.400 215.600 ;
        RECT 232.600 215.400 235.400 215.500 ;
        RECT 235.800 215.600 236.200 219.900 ;
        RECT 237.900 217.900 238.500 219.900 ;
        RECT 240.200 217.900 240.600 219.900 ;
        RECT 242.400 218.200 242.800 219.900 ;
        RECT 242.400 217.900 243.400 218.200 ;
        RECT 238.200 217.500 238.600 217.900 ;
        RECT 240.300 217.600 240.600 217.900 ;
        RECT 239.900 217.300 241.700 217.600 ;
        RECT 243.000 217.500 243.400 217.900 ;
        RECT 239.900 217.200 240.300 217.300 ;
        RECT 241.300 217.200 241.700 217.300 ;
        RECT 237.400 217.000 238.100 217.200 ;
        RECT 237.400 216.800 238.500 217.000 ;
        RECT 237.800 216.600 238.500 216.800 ;
        RECT 238.200 216.100 238.500 216.600 ;
        RECT 239.300 216.500 240.400 216.800 ;
        RECT 239.300 216.400 239.700 216.500 ;
        RECT 238.200 215.800 239.400 216.100 ;
        RECT 235.800 215.300 237.900 215.600 ;
        RECT 231.800 215.100 232.200 215.200 ;
        RECT 231.800 214.800 234.300 215.100 ;
        RECT 233.900 214.700 234.300 214.800 ;
        RECT 233.100 214.200 233.500 214.300 ;
        RECT 229.500 213.900 235.000 214.200 ;
        RECT 229.700 213.800 230.100 213.900 ;
        RECT 226.200 213.300 228.100 213.600 ;
        RECT 226.200 211.100 226.600 213.300 ;
        RECT 227.700 213.200 228.100 213.300 ;
        RECT 232.600 212.800 232.900 213.900 ;
        RECT 234.200 213.800 235.000 213.900 ;
        RECT 235.800 213.600 236.200 215.300 ;
        RECT 237.500 215.200 237.900 215.300 ;
        RECT 236.700 214.900 237.100 215.000 ;
        RECT 236.700 214.600 238.600 214.900 ;
        RECT 238.200 214.500 238.600 214.600 ;
        RECT 239.100 214.200 239.400 215.800 ;
        RECT 240.100 215.900 240.400 216.500 ;
        RECT 240.700 216.500 241.100 216.600 ;
        RECT 243.000 216.500 243.400 216.600 ;
        RECT 240.700 216.200 243.400 216.500 ;
        RECT 240.100 215.700 242.500 215.900 ;
        RECT 244.600 215.700 245.000 219.900 ;
        RECT 240.100 215.600 245.000 215.700 ;
        RECT 242.100 215.500 245.000 215.600 ;
        RECT 242.200 215.400 245.000 215.500 ;
        RECT 245.400 215.700 245.800 219.900 ;
        RECT 247.600 218.200 248.000 219.900 ;
        RECT 247.000 217.900 248.000 218.200 ;
        RECT 249.800 217.900 250.200 219.900 ;
        RECT 251.900 217.900 252.500 219.900 ;
        RECT 247.000 217.500 247.400 217.900 ;
        RECT 249.800 217.600 250.100 217.900 ;
        RECT 248.700 217.300 250.500 217.600 ;
        RECT 251.800 217.500 252.200 217.900 ;
        RECT 248.700 217.200 249.100 217.300 ;
        RECT 250.100 217.200 250.500 217.300 ;
        RECT 247.000 216.500 247.400 216.600 ;
        RECT 249.300 216.500 249.700 216.600 ;
        RECT 247.000 216.200 249.700 216.500 ;
        RECT 250.000 216.500 251.100 216.800 ;
        RECT 250.000 215.900 250.300 216.500 ;
        RECT 250.700 216.400 251.100 216.500 ;
        RECT 251.900 216.600 252.600 217.000 ;
        RECT 251.900 216.100 252.200 216.600 ;
        RECT 247.900 215.700 250.300 215.900 ;
        RECT 245.400 215.600 250.300 215.700 ;
        RECT 251.000 215.800 252.200 216.100 ;
        RECT 245.400 215.500 248.300 215.600 ;
        RECT 245.400 215.400 248.200 215.500 ;
        RECT 241.400 215.100 241.800 215.200 ;
        RECT 248.600 215.100 249.000 215.200 ;
        RECT 241.400 214.800 243.900 215.100 ;
        RECT 243.500 214.700 243.900 214.800 ;
        RECT 246.500 214.800 249.000 215.100 ;
        RECT 246.500 214.700 246.900 214.800 ;
        RECT 247.800 214.700 248.200 214.800 ;
        RECT 242.700 214.200 243.100 214.300 ;
        RECT 247.300 214.200 247.700 214.300 ;
        RECT 251.000 214.200 251.300 215.800 ;
        RECT 254.200 215.600 254.600 219.900 ;
        RECT 252.500 215.300 254.600 215.600 ;
        RECT 255.000 215.700 255.400 219.900 ;
        RECT 257.200 218.200 257.600 219.900 ;
        RECT 256.600 217.900 257.600 218.200 ;
        RECT 259.400 217.900 259.800 219.900 ;
        RECT 261.500 217.900 262.100 219.900 ;
        RECT 256.600 217.500 257.000 217.900 ;
        RECT 259.400 217.600 259.700 217.900 ;
        RECT 258.300 217.300 260.100 217.600 ;
        RECT 261.400 217.500 261.800 217.900 ;
        RECT 258.300 217.200 258.700 217.300 ;
        RECT 259.700 217.200 260.100 217.300 ;
        RECT 256.600 216.500 257.000 216.600 ;
        RECT 258.900 216.500 259.300 216.600 ;
        RECT 256.600 216.200 259.300 216.500 ;
        RECT 259.600 216.500 260.700 216.800 ;
        RECT 259.600 215.900 259.900 216.500 ;
        RECT 260.300 216.400 260.700 216.500 ;
        RECT 261.500 216.600 262.200 217.000 ;
        RECT 261.500 216.100 261.800 216.600 ;
        RECT 257.500 215.700 259.900 215.900 ;
        RECT 255.000 215.600 259.900 215.700 ;
        RECT 260.600 215.800 261.800 216.100 ;
        RECT 255.000 215.500 257.900 215.600 ;
        RECT 255.000 215.400 257.800 215.500 ;
        RECT 252.500 215.200 252.900 215.300 ;
        RECT 253.300 214.900 253.700 215.000 ;
        RECT 251.800 214.600 253.700 214.900 ;
        RECT 251.800 214.500 252.200 214.600 ;
        RECT 239.000 214.100 244.600 214.200 ;
        RECT 245.800 214.100 251.300 214.200 ;
        RECT 239.000 213.900 251.300 214.100 ;
        RECT 239.000 213.800 239.700 213.900 ;
        RECT 231.700 212.700 232.100 212.800 ;
        RECT 228.600 212.100 229.000 212.500 ;
        RECT 230.700 212.400 232.100 212.700 ;
        RECT 232.600 212.400 233.000 212.800 ;
        RECT 230.700 212.100 231.000 212.400 ;
        RECT 233.400 212.100 233.800 212.500 ;
        RECT 228.300 211.800 229.000 212.100 ;
        RECT 228.300 211.100 228.900 211.800 ;
        RECT 230.600 211.100 231.000 212.100 ;
        RECT 232.800 211.800 233.800 212.100 ;
        RECT 232.800 211.100 233.200 211.800 ;
        RECT 235.000 211.100 235.400 213.500 ;
        RECT 235.800 213.300 237.700 213.600 ;
        RECT 235.800 211.100 236.200 213.300 ;
        RECT 237.300 213.200 237.700 213.300 ;
        RECT 239.000 213.200 239.300 213.800 ;
        RECT 239.000 212.800 239.400 213.200 ;
        RECT 242.200 212.800 242.500 213.900 ;
        RECT 243.800 213.800 246.600 213.900 ;
        RECT 241.300 212.700 241.700 212.800 ;
        RECT 238.200 212.100 238.600 212.500 ;
        RECT 240.300 212.400 241.700 212.700 ;
        RECT 242.200 212.400 242.600 212.800 ;
        RECT 240.300 212.100 240.600 212.400 ;
        RECT 243.000 212.100 243.400 212.500 ;
        RECT 237.900 211.800 238.600 212.100 ;
        RECT 237.900 211.100 238.500 211.800 ;
        RECT 240.200 211.100 240.600 212.100 ;
        RECT 242.400 211.800 243.400 212.100 ;
        RECT 242.400 211.100 242.800 211.800 ;
        RECT 244.600 211.100 245.000 213.500 ;
        RECT 245.400 211.100 245.800 213.500 ;
        RECT 247.900 212.800 248.200 213.900 ;
        RECT 250.700 213.800 251.100 213.900 ;
        RECT 254.200 213.600 254.600 215.300 ;
        RECT 258.200 215.100 258.600 215.200 ;
        RECT 256.100 214.800 258.600 215.100 ;
        RECT 256.100 214.700 256.500 214.800 ;
        RECT 256.900 214.200 257.300 214.300 ;
        RECT 260.600 214.200 260.900 215.800 ;
        RECT 263.800 215.600 264.200 219.900 ;
        RECT 262.100 215.300 264.200 215.600 ;
        RECT 262.100 215.200 262.500 215.300 ;
        RECT 262.900 214.900 263.300 215.000 ;
        RECT 261.400 214.600 263.300 214.900 ;
        RECT 261.400 214.500 261.800 214.600 ;
        RECT 255.400 213.900 260.900 214.200 ;
        RECT 255.400 213.800 256.200 213.900 ;
        RECT 252.600 213.300 254.600 213.600 ;
        RECT 252.600 213.200 253.100 213.300 ;
        RECT 252.600 212.800 253.000 213.200 ;
        RECT 247.000 212.100 247.400 212.500 ;
        RECT 247.800 212.400 248.200 212.800 ;
        RECT 248.700 212.700 249.100 212.800 ;
        RECT 248.700 212.400 250.100 212.700 ;
        RECT 249.800 212.100 250.100 212.400 ;
        RECT 251.800 212.100 252.200 212.500 ;
        RECT 247.000 211.800 248.000 212.100 ;
        RECT 247.600 211.100 248.000 211.800 ;
        RECT 249.800 211.100 250.200 212.100 ;
        RECT 251.800 211.800 252.500 212.100 ;
        RECT 251.900 211.100 252.500 211.800 ;
        RECT 254.200 211.100 254.600 213.300 ;
        RECT 255.000 211.100 255.400 213.500 ;
        RECT 257.500 212.800 257.800 213.900 ;
        RECT 259.000 213.800 259.400 213.900 ;
        RECT 260.300 213.800 260.700 213.900 ;
        RECT 263.800 213.600 264.200 215.300 ;
        RECT 262.300 213.300 264.200 213.600 ;
        RECT 262.300 213.200 262.700 213.300 ;
        RECT 256.600 212.100 257.000 212.500 ;
        RECT 257.400 212.400 257.800 212.800 ;
        RECT 258.300 212.700 258.700 212.800 ;
        RECT 258.300 212.400 259.700 212.700 ;
        RECT 259.400 212.100 259.700 212.400 ;
        RECT 261.400 212.100 261.800 212.500 ;
        RECT 256.600 211.800 257.600 212.100 ;
        RECT 257.200 211.100 257.600 211.800 ;
        RECT 259.400 211.100 259.800 212.100 ;
        RECT 261.400 211.800 262.100 212.100 ;
        RECT 261.500 211.100 262.100 211.800 ;
        RECT 263.800 211.100 264.200 213.300 ;
        RECT 0.600 207.500 1.000 209.900 ;
        RECT 2.800 209.200 3.200 209.900 ;
        RECT 2.200 208.900 3.200 209.200 ;
        RECT 5.000 208.900 5.400 209.900 ;
        RECT 7.100 209.200 7.700 209.900 ;
        RECT 7.000 208.900 7.700 209.200 ;
        RECT 2.200 208.500 2.600 208.900 ;
        RECT 5.000 208.600 5.300 208.900 ;
        RECT 3.000 208.200 3.400 208.600 ;
        RECT 3.900 208.300 5.300 208.600 ;
        RECT 7.000 208.500 7.400 208.900 ;
        RECT 3.900 208.200 4.300 208.300 ;
        RECT 1.000 207.100 1.800 207.200 ;
        RECT 3.100 207.100 3.400 208.200 ;
        RECT 7.900 207.700 8.300 207.800 ;
        RECT 9.400 207.700 9.800 209.900 ;
        RECT 10.200 207.900 10.600 209.900 ;
        RECT 11.000 208.000 11.400 209.900 ;
        RECT 12.600 208.000 13.000 209.900 ;
        RECT 11.000 207.900 13.000 208.000 ;
        RECT 13.700 208.200 14.100 209.900 ;
        RECT 13.700 207.900 14.600 208.200 ;
        RECT 7.900 207.400 9.800 207.700 ;
        RECT 5.900 207.100 6.300 207.200 ;
        RECT 1.000 206.800 6.500 207.100 ;
        RECT 2.500 206.700 2.900 206.800 ;
        RECT 1.700 206.200 2.100 206.300 ;
        RECT 6.200 206.200 6.500 206.800 ;
        RECT 7.000 206.400 7.400 206.500 ;
        RECT 1.700 206.100 4.200 206.200 ;
        RECT 4.600 206.100 5.000 206.200 ;
        RECT 1.700 205.900 5.000 206.100 ;
        RECT 3.800 205.800 5.000 205.900 ;
        RECT 6.200 205.800 6.600 206.200 ;
        RECT 7.000 206.100 8.900 206.400 ;
        RECT 8.500 206.000 8.900 206.100 ;
        RECT 0.600 205.500 3.400 205.600 ;
        RECT 0.600 205.400 3.500 205.500 ;
        RECT 0.600 205.300 5.500 205.400 ;
        RECT 0.600 201.100 1.000 205.300 ;
        RECT 3.100 205.100 5.500 205.300 ;
        RECT 2.200 204.500 4.900 204.800 ;
        RECT 2.200 204.400 2.600 204.500 ;
        RECT 4.500 204.400 4.900 204.500 ;
        RECT 5.200 204.500 5.500 205.100 ;
        RECT 6.200 205.200 6.500 205.800 ;
        RECT 7.700 205.700 8.100 205.800 ;
        RECT 9.400 205.700 9.800 207.400 ;
        RECT 10.300 207.200 10.600 207.900 ;
        RECT 11.100 207.700 12.900 207.900 ;
        RECT 12.200 207.200 12.600 207.400 ;
        RECT 10.200 206.800 11.500 207.200 ;
        RECT 12.200 206.900 13.000 207.200 ;
        RECT 12.600 206.800 13.000 206.900 ;
        RECT 13.400 207.100 13.800 207.200 ;
        RECT 14.200 207.100 14.600 207.900 ;
        RECT 13.400 206.800 14.600 207.100 ;
        RECT 15.000 206.800 15.400 207.600 ;
        RECT 11.200 206.200 11.500 206.800 ;
        RECT 11.000 205.800 11.500 206.200 ;
        RECT 11.800 206.100 12.200 206.600 ;
        RECT 11.800 205.800 13.700 206.100 ;
        RECT 7.700 205.400 9.800 205.700 ;
        RECT 6.200 204.900 7.400 205.200 ;
        RECT 5.900 204.500 6.300 204.600 ;
        RECT 5.200 204.200 6.300 204.500 ;
        RECT 7.100 204.400 7.400 204.900 ;
        RECT 7.100 204.000 7.800 204.400 ;
        RECT 3.900 203.700 4.300 203.800 ;
        RECT 5.300 203.700 5.700 203.800 ;
        RECT 2.200 203.100 2.600 203.500 ;
        RECT 3.900 203.400 5.700 203.700 ;
        RECT 5.000 203.100 5.300 203.400 ;
        RECT 7.000 203.100 7.400 203.500 ;
        RECT 2.200 202.800 3.200 203.100 ;
        RECT 2.800 201.100 3.200 202.800 ;
        RECT 5.000 201.100 5.400 203.100 ;
        RECT 7.100 201.100 7.700 203.100 ;
        RECT 9.400 201.100 9.800 205.400 ;
        RECT 10.200 205.100 10.600 205.200 ;
        RECT 11.200 205.100 11.500 205.800 ;
        RECT 13.400 205.200 13.700 205.800 ;
        RECT 10.200 204.800 10.900 205.100 ;
        RECT 11.200 204.800 11.700 205.100 ;
        RECT 10.600 204.200 10.900 204.800 ;
        RECT 10.600 203.800 11.000 204.200 ;
        RECT 11.300 201.100 11.700 204.800 ;
        RECT 13.400 204.400 13.800 205.200 ;
        RECT 14.200 201.100 14.600 206.800 ;
        RECT 15.800 206.100 16.200 209.900 ;
        RECT 19.300 209.200 19.700 209.500 ;
        RECT 19.300 208.800 20.200 209.200 ;
        RECT 16.600 207.800 17.000 208.600 ;
        RECT 19.300 208.000 19.700 208.800 ;
        RECT 21.400 208.500 21.800 209.500 ;
        RECT 18.900 207.700 19.700 208.000 ;
        RECT 18.900 207.500 19.300 207.700 ;
        RECT 18.900 207.200 19.200 207.500 ;
        RECT 21.500 207.400 21.800 208.500 ;
        RECT 24.100 208.000 24.500 209.500 ;
        RECT 26.200 208.500 26.600 209.500 ;
        RECT 18.200 206.800 19.200 207.200 ;
        RECT 19.700 207.100 21.800 207.400 ;
        RECT 23.700 207.700 24.500 208.000 ;
        RECT 23.700 207.500 24.100 207.700 ;
        RECT 23.700 207.200 24.000 207.500 ;
        RECT 26.300 207.400 26.600 208.500 ;
        RECT 28.900 208.000 29.300 209.500 ;
        RECT 31.000 208.500 31.400 209.500 ;
        RECT 19.700 206.900 20.200 207.100 ;
        RECT 18.200 206.100 18.600 206.200 ;
        RECT 15.800 205.800 18.600 206.100 ;
        RECT 15.800 201.100 16.200 205.800 ;
        RECT 18.200 205.400 18.600 205.800 ;
        RECT 18.900 204.900 19.200 206.800 ;
        RECT 19.500 206.500 20.200 206.900 ;
        RECT 23.000 206.800 24.000 207.200 ;
        RECT 24.500 207.100 26.600 207.400 ;
        RECT 28.500 207.700 29.300 208.000 ;
        RECT 28.500 207.500 28.900 207.700 ;
        RECT 28.500 207.200 28.800 207.500 ;
        RECT 31.100 207.400 31.400 208.500 ;
        RECT 31.800 207.500 32.200 209.900 ;
        RECT 34.000 209.200 34.400 209.900 ;
        RECT 33.400 208.900 34.400 209.200 ;
        RECT 36.200 208.900 36.600 209.900 ;
        RECT 38.300 209.200 38.900 209.900 ;
        RECT 38.200 208.900 38.900 209.200 ;
        RECT 33.400 208.500 33.800 208.900 ;
        RECT 36.200 208.600 36.500 208.900 ;
        RECT 34.200 208.200 34.600 208.600 ;
        RECT 35.100 208.300 36.500 208.600 ;
        RECT 38.200 208.500 38.600 208.900 ;
        RECT 35.100 208.200 35.500 208.300 ;
        RECT 24.500 206.900 25.000 207.100 ;
        RECT 19.900 205.500 20.200 206.500 ;
        RECT 20.600 205.800 21.000 206.600 ;
        RECT 21.400 205.800 21.800 206.600 ;
        RECT 22.200 206.100 22.600 206.200 ;
        RECT 23.000 206.100 23.400 206.200 ;
        RECT 22.200 205.800 23.400 206.100 ;
        RECT 19.900 205.200 21.800 205.500 ;
        RECT 23.000 205.400 23.400 205.800 ;
        RECT 18.900 204.600 19.700 204.900 ;
        RECT 19.300 201.100 19.700 204.600 ;
        RECT 21.500 203.500 21.800 205.200 ;
        RECT 23.700 204.900 24.000 206.800 ;
        RECT 24.300 206.500 25.000 206.900 ;
        RECT 27.800 206.800 28.800 207.200 ;
        RECT 29.300 207.100 31.400 207.400 ;
        RECT 32.200 207.100 33.000 207.200 ;
        RECT 34.300 207.100 34.600 208.200 ;
        RECT 39.100 207.700 39.500 207.800 ;
        RECT 40.600 207.700 41.000 209.900 ;
        RECT 39.100 207.400 41.000 207.700 ;
        RECT 37.100 207.100 37.800 207.200 ;
        RECT 29.300 206.900 29.800 207.100 ;
        RECT 24.700 205.500 25.000 206.500 ;
        RECT 25.400 205.800 25.800 206.600 ;
        RECT 26.200 205.800 26.600 206.600 ;
        RECT 24.700 205.200 26.600 205.500 ;
        RECT 27.800 205.400 28.200 206.200 ;
        RECT 23.700 204.600 24.500 204.900 ;
        RECT 21.400 201.500 21.800 203.500 ;
        RECT 24.100 202.200 24.500 204.600 ;
        RECT 26.300 203.500 26.600 205.200 ;
        RECT 28.500 204.900 28.800 206.800 ;
        RECT 29.100 206.500 29.800 206.900 ;
        RECT 32.200 206.800 37.800 207.100 ;
        RECT 33.700 206.700 34.100 206.800 ;
        RECT 29.500 205.500 29.800 206.500 ;
        RECT 30.200 205.800 30.600 206.600 ;
        RECT 31.000 205.800 31.400 206.600 ;
        RECT 32.900 206.200 33.300 206.300 ;
        RECT 32.900 205.900 35.400 206.200 ;
        RECT 35.000 205.800 35.400 205.900 ;
        RECT 31.800 205.500 34.600 205.600 ;
        RECT 29.500 205.200 31.400 205.500 ;
        RECT 28.500 204.600 29.300 204.900 ;
        RECT 23.800 201.800 24.500 202.200 ;
        RECT 24.100 201.100 24.500 201.800 ;
        RECT 26.200 201.500 26.600 203.500 ;
        RECT 28.900 202.200 29.300 204.600 ;
        RECT 31.100 203.500 31.400 205.200 ;
        RECT 28.900 201.800 29.800 202.200 ;
        RECT 28.900 201.100 29.300 201.800 ;
        RECT 31.000 201.500 31.400 203.500 ;
        RECT 31.800 205.400 34.700 205.500 ;
        RECT 31.800 205.300 36.700 205.400 ;
        RECT 31.800 201.100 32.200 205.300 ;
        RECT 34.300 205.100 36.700 205.300 ;
        RECT 33.400 204.500 36.100 204.800 ;
        RECT 33.400 204.400 33.800 204.500 ;
        RECT 35.700 204.400 36.100 204.500 ;
        RECT 36.400 204.500 36.700 205.100 ;
        RECT 37.400 205.200 37.700 206.800 ;
        RECT 38.200 206.400 38.600 206.500 ;
        RECT 38.200 206.100 40.100 206.400 ;
        RECT 39.700 206.000 40.100 206.100 ;
        RECT 38.900 205.700 39.300 205.800 ;
        RECT 40.600 205.700 41.000 207.400 ;
        RECT 41.400 208.500 41.800 209.500 ;
        RECT 41.400 207.400 41.700 208.500 ;
        RECT 43.500 208.200 43.900 209.500 ;
        RECT 43.000 208.000 43.900 208.200 ;
        RECT 43.000 207.800 44.300 208.000 ;
        RECT 43.500 207.700 44.300 207.800 ;
        RECT 43.900 207.500 44.300 207.700 ;
        RECT 41.400 207.100 43.500 207.400 ;
        RECT 43.000 206.900 43.500 207.100 ;
        RECT 44.000 207.200 44.300 207.500 ;
        RECT 41.400 205.800 41.800 206.600 ;
        RECT 42.200 205.800 42.600 206.600 ;
        RECT 43.000 206.500 43.700 206.900 ;
        RECT 44.000 206.800 45.000 207.200 ;
        RECT 38.900 205.400 41.000 205.700 ;
        RECT 43.000 205.500 43.300 206.500 ;
        RECT 37.400 204.900 38.600 205.200 ;
        RECT 37.100 204.500 37.500 204.600 ;
        RECT 36.400 204.200 37.500 204.500 ;
        RECT 38.300 204.400 38.600 204.900 ;
        RECT 38.300 204.000 39.000 204.400 ;
        RECT 35.100 203.700 35.500 203.800 ;
        RECT 36.500 203.700 36.900 203.800 ;
        RECT 33.400 203.100 33.800 203.500 ;
        RECT 35.100 203.400 36.900 203.700 ;
        RECT 36.200 203.100 36.500 203.400 ;
        RECT 38.200 203.100 38.600 203.500 ;
        RECT 33.400 202.800 34.400 203.100 ;
        RECT 34.000 201.100 34.400 202.800 ;
        RECT 36.200 201.100 36.600 203.100 ;
        RECT 38.300 201.100 38.900 203.100 ;
        RECT 40.600 201.100 41.000 205.400 ;
        RECT 41.400 205.200 43.300 205.500 ;
        RECT 41.400 203.500 41.700 205.200 ;
        RECT 44.000 204.900 44.300 206.800 ;
        RECT 44.600 206.100 45.000 206.200 ;
        RECT 46.200 206.100 46.600 209.900 ;
        RECT 47.000 207.800 47.400 208.600 ;
        RECT 47.800 208.500 48.200 209.500 ;
        RECT 47.800 207.400 48.100 208.500 ;
        RECT 49.900 208.000 50.300 209.500 ;
        RECT 49.900 207.700 50.700 208.000 ;
        RECT 50.300 207.500 50.700 207.700 ;
        RECT 54.200 207.500 54.600 209.900 ;
        RECT 56.400 209.200 56.800 209.900 ;
        RECT 55.800 208.900 56.800 209.200 ;
        RECT 58.600 208.900 59.000 209.900 ;
        RECT 60.700 209.200 61.300 209.900 ;
        RECT 60.600 208.900 61.300 209.200 ;
        RECT 55.800 208.500 56.200 208.900 ;
        RECT 58.600 208.600 58.900 208.900 ;
        RECT 56.600 208.200 57.000 208.600 ;
        RECT 57.500 208.300 58.900 208.600 ;
        RECT 60.600 208.500 61.000 208.900 ;
        RECT 57.500 208.200 57.900 208.300 ;
        RECT 47.800 207.100 49.900 207.400 ;
        RECT 49.400 206.900 49.900 207.100 ;
        RECT 50.400 207.200 50.700 207.500 ;
        RECT 44.600 205.800 46.600 206.100 ;
        RECT 47.800 205.800 48.200 206.600 ;
        RECT 48.600 205.800 49.000 206.600 ;
        RECT 49.400 206.500 50.100 206.900 ;
        RECT 50.400 206.800 51.400 207.200 ;
        RECT 52.600 207.100 53.000 207.200 ;
        RECT 54.600 207.100 55.400 207.200 ;
        RECT 56.700 207.100 57.000 208.200 ;
        RECT 63.000 208.100 63.400 209.900 ;
        RECT 63.800 208.100 64.200 208.600 ;
        RECT 63.000 207.800 64.200 208.100 ;
        RECT 61.500 207.700 61.900 207.800 ;
        RECT 63.000 207.700 63.400 207.800 ;
        RECT 61.500 207.400 63.400 207.700 ;
        RECT 59.500 207.100 59.900 207.200 ;
        RECT 52.600 206.800 60.100 207.100 ;
        RECT 44.600 205.400 45.000 205.800 ;
        RECT 43.500 204.600 44.300 204.900 ;
        RECT 41.400 201.500 41.800 203.500 ;
        RECT 43.500 201.100 43.900 204.600 ;
        RECT 46.200 201.100 46.600 205.800 ;
        RECT 49.400 205.500 49.700 206.500 ;
        RECT 47.800 205.200 49.700 205.500 ;
        RECT 47.800 203.500 48.100 205.200 ;
        RECT 50.400 204.900 50.700 206.800 ;
        RECT 56.100 206.700 56.500 206.800 ;
        RECT 55.300 206.200 55.700 206.300 ;
        RECT 59.800 206.200 60.100 206.800 ;
        RECT 60.600 206.400 61.000 206.500 ;
        RECT 51.000 206.100 51.400 206.200 ;
        RECT 51.800 206.100 52.200 206.200 ;
        RECT 51.000 205.800 52.200 206.100 ;
        RECT 55.300 205.900 57.800 206.200 ;
        RECT 57.400 205.800 57.800 205.900 ;
        RECT 59.800 205.800 60.200 206.200 ;
        RECT 60.600 206.100 62.500 206.400 ;
        RECT 62.100 206.000 62.500 206.100 ;
        RECT 51.000 205.400 51.400 205.800 ;
        RECT 54.200 205.500 57.000 205.600 ;
        RECT 54.200 205.400 57.100 205.500 ;
        RECT 49.900 204.600 50.700 204.900 ;
        RECT 54.200 205.300 59.100 205.400 ;
        RECT 47.800 201.500 48.200 203.500 ;
        RECT 49.900 202.200 50.300 204.600 ;
        RECT 49.400 201.800 50.300 202.200 ;
        RECT 49.900 201.100 50.300 201.800 ;
        RECT 54.200 201.100 54.600 205.300 ;
        RECT 56.700 205.100 59.100 205.300 ;
        RECT 55.800 204.500 58.500 204.800 ;
        RECT 55.800 204.400 56.200 204.500 ;
        RECT 58.100 204.400 58.500 204.500 ;
        RECT 58.800 204.500 59.100 205.100 ;
        RECT 59.800 205.200 60.100 205.800 ;
        RECT 61.300 205.700 61.700 205.800 ;
        RECT 63.000 205.700 63.400 207.400 ;
        RECT 63.800 207.200 64.100 207.800 ;
        RECT 63.800 206.800 64.200 207.200 ;
        RECT 61.300 205.400 63.400 205.700 ;
        RECT 59.800 204.900 61.000 205.200 ;
        RECT 59.500 204.500 59.900 204.600 ;
        RECT 58.800 204.200 59.900 204.500 ;
        RECT 60.700 204.400 61.000 204.900 ;
        RECT 60.700 204.000 61.400 204.400 ;
        RECT 57.500 203.700 57.900 203.800 ;
        RECT 58.900 203.700 59.300 203.800 ;
        RECT 55.800 203.100 56.200 203.500 ;
        RECT 57.500 203.400 59.300 203.700 ;
        RECT 58.600 203.100 58.900 203.400 ;
        RECT 60.600 203.100 61.000 203.500 ;
        RECT 55.800 202.800 56.800 203.100 ;
        RECT 56.400 201.100 56.800 202.800 ;
        RECT 58.600 201.100 59.000 203.100 ;
        RECT 60.700 201.100 61.300 203.100 ;
        RECT 63.000 201.100 63.400 205.400 ;
        RECT 64.600 206.100 65.000 209.900 ;
        RECT 67.300 208.000 67.700 209.500 ;
        RECT 69.400 208.500 69.800 209.500 ;
        RECT 66.900 207.700 67.700 208.000 ;
        RECT 66.900 207.500 67.300 207.700 ;
        RECT 66.900 207.200 67.200 207.500 ;
        RECT 69.500 207.400 69.800 208.500 ;
        RECT 72.100 208.000 72.500 209.500 ;
        RECT 74.200 208.500 74.600 209.500 ;
        RECT 75.800 208.900 76.200 209.900 ;
        RECT 65.400 207.100 65.800 207.200 ;
        RECT 66.200 207.100 67.200 207.200 ;
        RECT 65.400 206.800 67.200 207.100 ;
        RECT 67.700 207.100 69.800 207.400 ;
        RECT 71.700 207.700 72.500 208.000 ;
        RECT 71.700 207.500 72.100 207.700 ;
        RECT 71.700 207.200 72.000 207.500 ;
        RECT 74.300 207.400 74.600 208.500 ;
        RECT 67.700 206.900 68.200 207.100 ;
        RECT 66.200 206.100 66.600 206.200 ;
        RECT 64.600 205.800 66.600 206.100 ;
        RECT 64.600 201.100 65.000 205.800 ;
        RECT 66.200 205.400 66.600 205.800 ;
        RECT 66.900 204.900 67.200 206.800 ;
        RECT 67.500 206.500 68.200 206.900 ;
        RECT 71.000 206.800 72.000 207.200 ;
        RECT 72.500 207.100 74.600 207.400 ;
        RECT 75.000 207.800 75.400 208.600 ;
        RECT 75.900 208.100 76.200 208.900 ;
        RECT 77.500 208.200 77.900 208.600 ;
        RECT 77.400 208.100 77.800 208.200 ;
        RECT 75.800 207.800 77.800 208.100 ;
        RECT 78.200 207.900 78.600 209.900 ;
        RECT 75.000 207.200 75.300 207.800 ;
        RECT 75.900 207.200 76.200 207.800 ;
        RECT 72.500 206.900 73.000 207.100 ;
        RECT 67.900 205.500 68.200 206.500 ;
        RECT 68.600 205.800 69.000 206.600 ;
        RECT 69.400 205.800 69.800 206.600 ;
        RECT 67.900 205.200 69.800 205.500 ;
        RECT 71.000 205.400 71.400 206.200 ;
        RECT 66.900 204.600 67.700 204.900 ;
        RECT 67.300 201.100 67.700 204.600 ;
        RECT 69.500 203.500 69.800 205.200 ;
        RECT 71.700 204.900 72.000 206.800 ;
        RECT 72.300 206.500 73.000 206.900 ;
        RECT 75.000 206.800 75.400 207.200 ;
        RECT 75.800 206.800 76.200 207.200 ;
        RECT 72.700 205.500 73.000 206.500 ;
        RECT 73.400 205.800 73.800 206.600 ;
        RECT 74.200 205.800 74.600 206.600 ;
        RECT 72.700 205.200 74.600 205.500 ;
        RECT 71.700 204.600 72.500 204.900 ;
        RECT 69.400 201.500 69.800 203.500 ;
        RECT 72.100 202.200 72.500 204.600 ;
        RECT 74.300 203.500 74.600 205.200 ;
        RECT 75.900 205.100 76.200 206.800 ;
        RECT 76.600 205.400 77.000 206.200 ;
        RECT 77.400 206.100 77.800 206.200 ;
        RECT 78.300 206.100 78.600 207.900 ;
        RECT 80.600 207.500 81.000 209.900 ;
        RECT 82.800 209.200 83.200 209.900 ;
        RECT 82.200 208.900 83.200 209.200 ;
        RECT 85.000 208.900 85.400 209.900 ;
        RECT 87.100 209.200 87.700 209.900 ;
        RECT 87.000 208.900 87.700 209.200 ;
        RECT 82.200 208.500 82.600 208.900 ;
        RECT 85.000 208.600 85.300 208.900 ;
        RECT 83.000 208.200 83.400 208.600 ;
        RECT 83.900 208.300 85.300 208.600 ;
        RECT 87.000 208.500 87.400 208.900 ;
        RECT 83.900 208.200 84.300 208.300 ;
        RECT 79.000 206.400 79.400 207.200 ;
        RECT 81.000 207.100 81.800 207.200 ;
        RECT 83.100 207.100 83.400 208.200 ;
        RECT 87.900 207.700 88.300 207.800 ;
        RECT 89.400 207.700 89.800 209.900 ;
        RECT 90.200 207.900 90.600 209.900 ;
        RECT 91.000 208.000 91.400 209.900 ;
        RECT 92.600 208.000 93.000 209.900 ;
        RECT 91.000 207.900 93.000 208.000 ;
        RECT 93.400 208.500 93.800 209.500 ;
        RECT 87.900 207.400 89.800 207.700 ;
        RECT 85.900 207.100 86.300 207.200 ;
        RECT 81.000 206.800 86.500 207.100 ;
        RECT 82.500 206.700 82.900 206.800 ;
        RECT 81.700 206.200 82.100 206.300 ;
        RECT 79.800 206.100 80.200 206.200 ;
        RECT 77.400 205.800 78.600 206.100 ;
        RECT 79.400 205.800 80.200 206.100 ;
        RECT 81.700 206.100 84.200 206.200 ;
        RECT 84.600 206.100 85.000 206.200 ;
        RECT 81.700 205.900 85.000 206.100 ;
        RECT 83.800 205.800 85.000 205.900 ;
        RECT 77.500 205.100 77.800 205.800 ;
        RECT 79.400 205.600 79.800 205.800 ;
        RECT 80.600 205.500 83.400 205.600 ;
        RECT 80.600 205.400 83.500 205.500 ;
        RECT 80.600 205.300 85.500 205.400 ;
        RECT 75.800 204.700 76.700 205.100 ;
        RECT 72.100 201.800 73.000 202.200 ;
        RECT 72.100 201.100 72.500 201.800 ;
        RECT 74.200 201.500 74.600 203.500 ;
        RECT 76.300 201.100 76.700 204.700 ;
        RECT 77.400 201.100 77.800 205.100 ;
        RECT 78.200 204.800 80.200 205.100 ;
        RECT 78.200 201.100 78.600 204.800 ;
        RECT 79.800 201.100 80.200 204.800 ;
        RECT 80.600 201.100 81.000 205.300 ;
        RECT 83.100 205.100 85.500 205.300 ;
        RECT 82.200 204.500 84.900 204.800 ;
        RECT 82.200 204.400 82.600 204.500 ;
        RECT 84.500 204.400 84.900 204.500 ;
        RECT 85.200 204.500 85.500 205.100 ;
        RECT 86.200 205.200 86.500 206.800 ;
        RECT 87.000 206.400 87.400 206.500 ;
        RECT 87.000 206.100 88.900 206.400 ;
        RECT 88.500 206.000 88.900 206.100 ;
        RECT 87.700 205.700 88.100 205.800 ;
        RECT 89.400 205.700 89.800 207.400 ;
        RECT 90.300 207.200 90.600 207.900 ;
        RECT 91.100 207.700 92.900 207.900 ;
        RECT 93.400 207.400 93.700 208.500 ;
        RECT 95.500 208.000 95.900 209.500 ;
        RECT 99.000 208.800 99.400 209.900 ;
        RECT 95.500 207.700 96.300 208.000 ;
        RECT 98.200 207.800 98.600 208.600 ;
        RECT 95.900 207.500 96.300 207.700 ;
        RECT 92.200 207.200 92.600 207.400 ;
        RECT 90.200 206.800 91.500 207.200 ;
        RECT 92.200 206.900 93.000 207.200 ;
        RECT 93.400 207.100 95.500 207.400 ;
        RECT 92.600 206.800 93.000 206.900 ;
        RECT 95.000 206.900 95.500 207.100 ;
        RECT 96.000 207.200 96.300 207.500 ;
        RECT 99.100 207.200 99.400 208.800 ;
        RECT 102.500 208.000 102.900 209.500 ;
        RECT 104.600 208.500 105.000 209.500 ;
        RECT 102.100 207.700 102.900 208.000 ;
        RECT 102.100 207.500 102.500 207.700 ;
        RECT 102.100 207.200 102.400 207.500 ;
        RECT 104.700 207.400 105.000 208.500 ;
        RECT 87.700 205.400 89.800 205.700 ;
        RECT 86.200 204.900 87.400 205.200 ;
        RECT 85.900 204.500 86.300 204.600 ;
        RECT 85.200 204.200 86.300 204.500 ;
        RECT 87.100 204.400 87.400 204.900 ;
        RECT 87.100 204.000 87.800 204.400 ;
        RECT 83.900 203.700 84.300 203.800 ;
        RECT 85.300 203.700 85.700 203.800 ;
        RECT 82.200 203.100 82.600 203.500 ;
        RECT 83.900 203.400 85.700 203.700 ;
        RECT 85.000 203.100 85.300 203.400 ;
        RECT 87.000 203.100 87.400 203.500 ;
        RECT 82.200 202.800 83.200 203.100 ;
        RECT 82.800 201.100 83.200 202.800 ;
        RECT 85.000 201.100 85.400 203.100 ;
        RECT 87.100 201.100 87.700 203.100 ;
        RECT 89.400 201.100 89.800 205.400 ;
        RECT 90.200 205.100 90.600 205.200 ;
        RECT 91.200 205.100 91.500 206.800 ;
        RECT 91.800 205.800 92.200 206.600 ;
        RECT 93.400 205.800 93.800 206.600 ;
        RECT 94.200 205.800 94.600 206.600 ;
        RECT 95.000 206.500 95.700 206.900 ;
        RECT 96.000 206.800 97.000 207.200 ;
        RECT 99.000 206.800 99.400 207.200 ;
        RECT 101.400 206.800 102.400 207.200 ;
        RECT 102.900 207.100 105.000 207.400 ;
        RECT 107.000 208.500 107.400 209.500 ;
        RECT 107.000 207.400 107.300 208.500 ;
        RECT 109.100 208.000 109.500 209.500 ;
        RECT 111.800 208.500 112.200 209.500 ;
        RECT 113.900 209.200 114.300 209.500 ;
        RECT 113.900 208.800 114.600 209.200 ;
        RECT 109.100 207.700 109.900 208.000 ;
        RECT 109.500 207.500 109.900 207.700 ;
        RECT 107.000 207.100 109.100 207.400 ;
        RECT 102.900 206.900 103.400 207.100 ;
        RECT 95.000 205.500 95.300 206.500 ;
        RECT 93.400 205.200 95.300 205.500 ;
        RECT 90.200 204.800 90.900 205.100 ;
        RECT 91.200 204.800 91.700 205.100 ;
        RECT 90.600 204.200 90.900 204.800 ;
        RECT 90.600 203.800 91.000 204.200 ;
        RECT 91.300 201.100 91.700 204.800 ;
        RECT 93.400 203.500 93.700 205.200 ;
        RECT 96.000 204.900 96.300 206.800 ;
        RECT 96.600 205.400 97.000 206.200 ;
        RECT 99.100 205.100 99.400 206.800 ;
        RECT 99.800 205.400 100.200 206.200 ;
        RECT 101.400 205.400 101.800 206.200 ;
        RECT 95.500 204.600 96.300 204.900 ;
        RECT 99.000 204.700 99.900 205.100 ;
        RECT 93.400 201.500 93.800 203.500 ;
        RECT 95.500 202.200 95.900 204.600 ;
        RECT 95.000 201.800 95.900 202.200 ;
        RECT 95.500 201.100 95.900 201.800 ;
        RECT 99.500 201.100 99.900 204.700 ;
        RECT 102.100 204.900 102.400 206.800 ;
        RECT 102.700 206.500 103.400 206.900 ;
        RECT 108.600 206.900 109.100 207.100 ;
        RECT 109.600 207.200 109.900 207.500 ;
        RECT 111.800 207.400 112.100 208.500 ;
        RECT 113.900 208.000 114.300 208.800 ;
        RECT 116.600 208.000 117.000 209.900 ;
        RECT 118.200 208.000 118.600 209.900 ;
        RECT 113.900 207.700 114.700 208.000 ;
        RECT 116.600 207.900 118.600 208.000 ;
        RECT 116.700 207.700 118.500 207.900 ;
        RECT 119.000 207.800 119.400 209.900 ;
        RECT 120.100 208.200 120.500 209.900 ;
        RECT 120.100 207.900 121.000 208.200 ;
        RECT 114.300 207.500 114.700 207.700 ;
        RECT 103.100 205.500 103.400 206.500 ;
        RECT 103.800 205.800 104.200 206.600 ;
        RECT 104.600 205.800 105.000 206.600 ;
        RECT 107.000 205.800 107.400 206.600 ;
        RECT 107.800 205.800 108.200 206.600 ;
        RECT 108.600 206.500 109.300 206.900 ;
        RECT 109.600 206.800 110.600 207.200 ;
        RECT 111.800 207.100 113.900 207.400 ;
        RECT 113.400 206.900 113.900 207.100 ;
        RECT 114.400 207.200 114.700 207.500 ;
        RECT 117.000 207.200 117.400 207.400 ;
        RECT 119.000 207.200 119.300 207.800 ;
        RECT 108.600 205.500 108.900 206.500 ;
        RECT 103.100 205.200 105.000 205.500 ;
        RECT 102.100 204.600 102.900 204.900 ;
        RECT 102.500 202.200 102.900 204.600 ;
        RECT 104.700 203.500 105.000 205.200 ;
        RECT 102.200 201.800 102.900 202.200 ;
        RECT 102.500 201.100 102.900 201.800 ;
        RECT 104.600 201.500 105.000 203.500 ;
        RECT 107.000 205.200 108.900 205.500 ;
        RECT 107.000 203.500 107.300 205.200 ;
        RECT 109.600 204.900 109.900 206.800 ;
        RECT 110.200 206.100 110.600 206.200 ;
        RECT 111.000 206.100 111.400 206.200 ;
        RECT 110.200 205.800 111.400 206.100 ;
        RECT 111.800 205.800 112.200 206.600 ;
        RECT 112.600 205.800 113.000 206.600 ;
        RECT 113.400 206.500 114.100 206.900 ;
        RECT 114.400 206.800 115.400 207.200 ;
        RECT 116.600 206.900 117.400 207.200 ;
        RECT 116.600 206.800 117.000 206.900 ;
        RECT 118.100 206.800 119.400 207.200 ;
        RECT 110.200 205.400 110.600 205.800 ;
        RECT 113.400 205.500 113.700 206.500 ;
        RECT 109.100 204.600 109.900 204.900 ;
        RECT 111.800 205.200 113.700 205.500 ;
        RECT 107.000 201.500 107.400 203.500 ;
        RECT 109.100 202.200 109.500 204.600 ;
        RECT 108.600 201.800 109.500 202.200 ;
        RECT 109.100 201.100 109.500 201.800 ;
        RECT 111.800 203.500 112.100 205.200 ;
        RECT 114.400 204.900 114.700 206.800 ;
        RECT 115.000 205.400 115.400 206.200 ;
        RECT 117.400 205.800 117.800 206.600 ;
        RECT 118.100 205.100 118.400 206.800 ;
        RECT 120.600 206.100 121.000 207.900 ;
        RECT 122.200 207.700 122.600 209.900 ;
        RECT 124.300 209.200 124.900 209.900 ;
        RECT 124.300 208.900 125.000 209.200 ;
        RECT 126.600 208.900 127.000 209.900 ;
        RECT 128.800 209.200 129.200 209.900 ;
        RECT 128.800 208.900 129.800 209.200 ;
        RECT 124.600 208.500 125.000 208.900 ;
        RECT 126.700 208.600 127.000 208.900 ;
        RECT 126.700 208.300 128.100 208.600 ;
        RECT 127.700 208.200 128.100 208.300 ;
        RECT 128.600 208.200 129.000 208.600 ;
        RECT 129.400 208.500 129.800 208.900 ;
        RECT 123.700 207.700 124.100 207.800 ;
        RECT 121.400 207.100 121.800 207.600 ;
        RECT 122.200 207.400 124.100 207.700 ;
        RECT 122.200 207.100 122.600 207.400 ;
        RECT 125.700 207.100 126.100 207.200 ;
        RECT 128.600 207.100 128.900 208.200 ;
        RECT 131.000 207.500 131.400 209.900 ;
        RECT 131.800 207.500 132.200 209.900 ;
        RECT 134.000 209.200 134.400 209.900 ;
        RECT 133.400 208.900 134.400 209.200 ;
        RECT 136.200 208.900 136.600 209.900 ;
        RECT 138.300 209.200 138.900 209.900 ;
        RECT 138.200 208.900 138.900 209.200 ;
        RECT 133.400 208.500 133.800 208.900 ;
        RECT 136.200 208.600 136.500 208.900 ;
        RECT 134.200 208.200 134.600 208.600 ;
        RECT 135.100 208.300 136.500 208.600 ;
        RECT 138.200 208.500 138.600 208.900 ;
        RECT 135.100 208.200 135.500 208.300 ;
        RECT 130.200 207.100 131.000 207.200 ;
        RECT 121.400 206.800 122.600 207.100 ;
        RECT 119.000 205.800 121.000 206.100 ;
        RECT 119.000 205.200 119.300 205.800 ;
        RECT 119.000 205.100 119.400 205.200 ;
        RECT 113.900 204.600 114.700 204.900 ;
        RECT 117.900 204.800 118.400 205.100 ;
        RECT 118.700 204.800 119.400 205.100 ;
        RECT 111.800 201.500 112.200 203.500 ;
        RECT 113.900 201.100 114.300 204.600 ;
        RECT 117.900 201.100 118.300 204.800 ;
        RECT 118.700 204.200 119.000 204.800 ;
        RECT 119.800 204.400 120.200 205.200 ;
        RECT 118.600 203.800 119.000 204.200 ;
        RECT 120.600 201.100 121.000 205.800 ;
        RECT 122.200 205.700 122.600 206.800 ;
        RECT 125.500 206.800 131.000 207.100 ;
        RECT 132.200 207.100 133.000 207.200 ;
        RECT 134.300 207.100 134.600 208.200 ;
        RECT 139.100 207.700 139.500 207.800 ;
        RECT 140.600 207.700 141.000 209.900 ;
        RECT 141.400 208.000 141.800 209.900 ;
        RECT 143.000 208.000 143.400 209.900 ;
        RECT 141.400 207.900 143.400 208.000 ;
        RECT 143.800 207.900 144.200 209.900 ;
        RECT 144.900 208.200 145.300 209.900 ;
        RECT 147.000 208.500 147.400 209.500 ;
        RECT 144.900 207.900 145.800 208.200 ;
        RECT 141.500 207.700 143.300 207.900 ;
        RECT 139.100 207.400 141.000 207.700 ;
        RECT 135.800 207.100 136.200 207.200 ;
        RECT 137.100 207.100 137.500 207.200 ;
        RECT 132.200 206.800 137.700 207.100 ;
        RECT 124.600 206.400 125.000 206.500 ;
        RECT 123.100 206.100 125.000 206.400 ;
        RECT 123.100 206.000 123.500 206.100 ;
        RECT 123.900 205.700 124.300 205.800 ;
        RECT 122.200 205.400 124.300 205.700 ;
        RECT 122.200 201.100 122.600 205.400 ;
        RECT 125.500 205.200 125.800 206.800 ;
        RECT 129.100 206.700 129.500 206.800 ;
        RECT 133.700 206.700 134.100 206.800 ;
        RECT 129.900 206.200 130.300 206.300 ;
        RECT 127.800 205.900 130.300 206.200 ;
        RECT 132.900 206.200 133.300 206.300 ;
        RECT 132.900 205.900 135.400 206.200 ;
        RECT 127.800 205.800 128.200 205.900 ;
        RECT 135.000 205.800 135.400 205.900 ;
        RECT 128.600 205.500 131.400 205.600 ;
        RECT 128.500 205.400 131.400 205.500 ;
        RECT 124.600 204.900 125.800 205.200 ;
        RECT 126.500 205.300 131.400 205.400 ;
        RECT 126.500 205.100 128.900 205.300 ;
        RECT 124.600 204.400 124.900 204.900 ;
        RECT 124.200 204.000 124.900 204.400 ;
        RECT 125.700 204.500 126.100 204.600 ;
        RECT 126.500 204.500 126.800 205.100 ;
        RECT 125.700 204.200 126.800 204.500 ;
        RECT 127.100 204.500 129.800 204.800 ;
        RECT 127.100 204.400 127.500 204.500 ;
        RECT 129.400 204.400 129.800 204.500 ;
        RECT 126.300 203.700 126.700 203.800 ;
        RECT 127.700 203.700 128.100 203.800 ;
        RECT 124.600 203.100 125.000 203.500 ;
        RECT 126.300 203.400 128.100 203.700 ;
        RECT 126.700 203.100 127.000 203.400 ;
        RECT 129.400 203.100 129.800 203.500 ;
        RECT 124.300 201.100 124.900 203.100 ;
        RECT 126.600 201.100 127.000 203.100 ;
        RECT 128.800 202.800 129.800 203.100 ;
        RECT 128.800 201.100 129.200 202.800 ;
        RECT 131.000 201.100 131.400 205.300 ;
        RECT 131.800 205.500 134.600 205.600 ;
        RECT 131.800 205.400 134.700 205.500 ;
        RECT 131.800 205.300 136.700 205.400 ;
        RECT 131.800 201.100 132.200 205.300 ;
        RECT 134.300 205.100 136.700 205.300 ;
        RECT 133.400 204.500 136.100 204.800 ;
        RECT 133.400 204.400 133.800 204.500 ;
        RECT 135.700 204.400 136.100 204.500 ;
        RECT 136.400 204.500 136.700 205.100 ;
        RECT 137.400 205.200 137.700 206.800 ;
        RECT 138.200 206.400 138.600 206.500 ;
        RECT 138.200 206.100 140.100 206.400 ;
        RECT 139.700 206.000 140.100 206.100 ;
        RECT 138.900 205.700 139.300 205.800 ;
        RECT 140.600 205.700 141.000 207.400 ;
        RECT 141.800 207.200 142.200 207.400 ;
        RECT 143.800 207.200 144.100 207.900 ;
        RECT 141.400 206.900 142.200 207.200 ;
        RECT 141.400 206.800 141.800 206.900 ;
        RECT 142.900 206.800 144.200 207.200 ;
        RECT 142.200 205.800 142.600 206.600 ;
        RECT 138.900 205.400 141.000 205.700 ;
        RECT 137.400 204.900 138.600 205.200 ;
        RECT 137.100 204.500 137.500 204.600 ;
        RECT 136.400 204.200 137.500 204.500 ;
        RECT 138.300 204.400 138.600 204.900 ;
        RECT 138.300 204.000 139.000 204.400 ;
        RECT 135.100 203.700 135.500 203.800 ;
        RECT 136.500 203.700 136.900 203.800 ;
        RECT 133.400 203.100 133.800 203.500 ;
        RECT 135.100 203.400 136.900 203.700 ;
        RECT 136.200 203.100 136.500 203.400 ;
        RECT 138.200 203.100 138.600 203.500 ;
        RECT 133.400 202.800 134.400 203.100 ;
        RECT 134.000 201.100 134.400 202.800 ;
        RECT 136.200 201.100 136.600 203.100 ;
        RECT 138.300 201.100 138.900 203.100 ;
        RECT 140.600 201.100 141.000 205.400 ;
        RECT 142.900 205.100 143.200 206.800 ;
        RECT 145.400 206.100 145.800 207.900 ;
        RECT 146.200 206.800 146.600 207.600 ;
        RECT 147.000 207.400 147.300 208.500 ;
        RECT 149.100 208.000 149.500 209.500 ;
        RECT 149.100 207.700 149.900 208.000 ;
        RECT 151.800 207.900 152.200 209.900 ;
        RECT 152.600 208.000 153.000 209.900 ;
        RECT 154.200 208.000 154.600 209.900 ;
        RECT 152.600 207.900 154.600 208.000 ;
        RECT 155.000 207.900 155.400 209.900 ;
        RECT 155.800 208.000 156.200 209.900 ;
        RECT 157.400 208.000 157.800 209.900 ;
        RECT 155.800 207.900 157.800 208.000 ;
        RECT 159.800 208.000 160.200 209.900 ;
        RECT 161.400 208.000 161.800 209.900 ;
        RECT 159.800 207.900 161.800 208.000 ;
        RECT 162.200 207.900 162.600 209.900 ;
        RECT 163.300 208.200 163.700 209.900 ;
        RECT 163.300 207.900 164.200 208.200 ;
        RECT 149.500 207.500 149.900 207.700 ;
        RECT 147.000 207.100 149.100 207.400 ;
        RECT 148.600 206.900 149.100 207.100 ;
        RECT 149.600 207.200 149.900 207.500 ;
        RECT 151.900 207.200 152.200 207.900 ;
        RECT 152.700 207.700 154.500 207.900 ;
        RECT 153.800 207.200 154.200 207.400 ;
        RECT 155.100 207.200 155.400 207.900 ;
        RECT 155.900 207.700 157.700 207.900 ;
        RECT 159.900 207.700 161.700 207.900 ;
        RECT 157.000 207.200 157.400 207.400 ;
        RECT 160.200 207.200 160.600 207.400 ;
        RECT 162.200 207.200 162.500 207.900 ;
        RECT 143.800 205.800 145.800 206.100 ;
        RECT 147.000 205.800 147.400 206.600 ;
        RECT 147.800 205.800 148.200 206.600 ;
        RECT 148.600 206.500 149.300 206.900 ;
        RECT 149.600 206.800 150.600 207.200 ;
        RECT 151.800 206.800 153.100 207.200 ;
        RECT 153.800 206.900 154.600 207.200 ;
        RECT 154.200 206.800 154.600 206.900 ;
        RECT 155.000 206.800 156.300 207.200 ;
        RECT 157.000 206.900 157.800 207.200 ;
        RECT 157.400 206.800 157.800 206.900 ;
        RECT 159.800 206.900 160.600 207.200 ;
        RECT 161.300 207.100 162.600 207.200 ;
        RECT 163.000 207.100 163.400 207.200 ;
        RECT 159.800 206.800 160.200 206.900 ;
        RECT 161.300 206.800 163.400 207.100 ;
        RECT 143.800 205.200 144.100 205.800 ;
        RECT 143.800 205.100 144.200 205.200 ;
        RECT 142.700 204.800 143.200 205.100 ;
        RECT 143.500 204.800 144.200 205.100 ;
        RECT 142.700 204.200 143.100 204.800 ;
        RECT 143.500 204.200 143.800 204.800 ;
        RECT 144.600 204.400 145.000 205.200 ;
        RECT 142.200 203.800 143.100 204.200 ;
        RECT 143.400 203.800 143.800 204.200 ;
        RECT 142.700 201.100 143.100 203.800 ;
        RECT 145.400 201.100 145.800 205.800 ;
        RECT 148.600 205.500 148.900 206.500 ;
        RECT 147.000 205.200 148.900 205.500 ;
        RECT 147.000 203.500 147.300 205.200 ;
        RECT 149.600 204.900 149.900 206.800 ;
        RECT 150.200 206.100 150.600 206.200 ;
        RECT 151.000 206.100 151.400 206.200 ;
        RECT 150.200 205.800 152.100 206.100 ;
        RECT 150.200 205.400 150.600 205.800 ;
        RECT 149.100 204.600 149.900 204.900 ;
        RECT 151.800 205.200 152.100 205.800 ;
        RECT 152.800 205.200 153.100 206.800 ;
        RECT 153.400 206.100 153.800 206.600 ;
        RECT 154.200 206.100 154.600 206.200 ;
        RECT 153.400 205.800 154.600 206.100 ;
        RECT 151.800 205.100 152.200 205.200 ;
        RECT 151.800 204.800 152.500 205.100 ;
        RECT 152.800 204.800 153.800 205.200 ;
        RECT 155.000 205.100 155.400 205.200 ;
        RECT 156.000 205.100 156.300 206.800 ;
        RECT 156.600 206.100 157.000 206.600 ;
        RECT 159.800 206.100 160.200 206.200 ;
        RECT 156.600 205.800 160.200 206.100 ;
        RECT 160.600 205.800 161.000 206.600 ;
        RECT 161.300 205.100 161.600 206.800 ;
        RECT 163.800 206.100 164.200 207.900 ;
        RECT 165.400 207.700 165.800 209.900 ;
        RECT 167.500 209.200 168.100 209.900 ;
        RECT 167.500 208.900 168.200 209.200 ;
        RECT 169.800 208.900 170.200 209.900 ;
        RECT 172.000 209.200 172.400 209.900 ;
        RECT 172.000 208.900 173.000 209.200 ;
        RECT 167.800 208.500 168.200 208.900 ;
        RECT 169.900 208.600 170.200 208.900 ;
        RECT 169.900 208.300 171.300 208.600 ;
        RECT 170.900 208.200 171.300 208.300 ;
        RECT 171.800 207.800 172.200 208.600 ;
        RECT 172.600 208.500 173.000 208.900 ;
        RECT 166.900 207.700 167.300 207.800 ;
        RECT 164.600 206.800 165.000 207.600 ;
        RECT 165.400 207.400 167.300 207.700 ;
        RECT 162.200 205.800 164.200 206.100 ;
        RECT 162.200 205.200 162.500 205.800 ;
        RECT 162.200 205.100 162.600 205.200 ;
        RECT 155.000 204.800 155.700 205.100 ;
        RECT 156.000 204.800 156.500 205.100 ;
        RECT 147.000 201.500 147.400 203.500 ;
        RECT 149.100 201.100 149.500 204.600 ;
        RECT 152.200 204.200 152.500 204.800 ;
        RECT 152.200 203.800 152.600 204.200 ;
        RECT 152.900 201.100 153.300 204.800 ;
        RECT 155.400 204.200 155.700 204.800 ;
        RECT 155.400 203.800 155.800 204.200 ;
        RECT 156.100 201.100 156.500 204.800 ;
        RECT 161.100 204.800 161.600 205.100 ;
        RECT 161.900 204.800 162.600 205.100 ;
        RECT 161.100 201.100 161.500 204.800 ;
        RECT 161.900 204.200 162.200 204.800 ;
        RECT 163.000 204.400 163.400 205.200 ;
        RECT 161.800 203.800 162.200 204.200 ;
        RECT 163.800 201.100 164.200 205.800 ;
        RECT 165.400 205.700 165.800 207.400 ;
        RECT 168.900 207.100 169.300 207.200 ;
        RECT 171.800 207.100 172.100 207.800 ;
        RECT 174.200 207.500 174.600 209.900 ;
        RECT 175.000 207.700 175.400 209.900 ;
        RECT 177.100 209.200 177.700 209.900 ;
        RECT 177.100 208.900 177.800 209.200 ;
        RECT 179.400 208.900 179.800 209.900 ;
        RECT 181.600 209.200 182.000 209.900 ;
        RECT 181.600 208.900 182.600 209.200 ;
        RECT 177.400 208.500 177.800 208.900 ;
        RECT 179.500 208.600 179.800 208.900 ;
        RECT 179.500 208.300 180.900 208.600 ;
        RECT 180.500 208.200 180.900 208.300 ;
        RECT 181.400 208.200 181.800 208.600 ;
        RECT 182.200 208.500 182.600 208.900 ;
        RECT 176.500 207.700 176.900 207.800 ;
        RECT 175.000 207.400 176.900 207.700 ;
        RECT 173.400 207.100 174.200 207.200 ;
        RECT 168.700 206.800 174.200 207.100 ;
        RECT 167.800 206.400 168.200 206.500 ;
        RECT 166.300 206.100 168.200 206.400 ;
        RECT 168.700 206.100 169.000 206.800 ;
        RECT 172.300 206.700 172.700 206.800 ;
        RECT 173.100 206.200 173.500 206.300 ;
        RECT 169.400 206.100 169.800 206.200 ;
        RECT 166.300 206.000 166.700 206.100 ;
        RECT 168.600 205.800 169.800 206.100 ;
        RECT 171.000 205.900 173.500 206.200 ;
        RECT 171.000 205.800 171.400 205.900 ;
        RECT 167.100 205.700 167.500 205.800 ;
        RECT 165.400 205.400 167.500 205.700 ;
        RECT 164.600 204.100 165.000 204.200 ;
        RECT 165.400 204.100 165.800 205.400 ;
        RECT 168.700 205.200 169.000 205.800 ;
        RECT 175.000 205.700 175.400 207.400 ;
        RECT 178.500 207.100 178.900 207.200 ;
        RECT 181.400 207.100 181.700 208.200 ;
        RECT 183.800 207.500 184.200 209.900 ;
        RECT 184.600 207.700 185.000 209.900 ;
        RECT 186.700 209.200 187.300 209.900 ;
        RECT 186.700 208.900 187.400 209.200 ;
        RECT 189.000 208.900 189.400 209.900 ;
        RECT 191.200 209.200 191.600 209.900 ;
        RECT 191.200 208.900 192.200 209.200 ;
        RECT 187.000 208.500 187.400 208.900 ;
        RECT 189.100 208.600 189.400 208.900 ;
        RECT 189.100 208.300 190.500 208.600 ;
        RECT 190.100 208.200 190.500 208.300 ;
        RECT 191.000 207.800 191.400 208.600 ;
        RECT 191.800 208.500 192.200 208.900 ;
        RECT 186.100 207.700 186.500 207.800 ;
        RECT 184.600 207.400 186.500 207.700 ;
        RECT 183.000 207.100 183.800 207.200 ;
        RECT 178.300 206.800 183.800 207.100 ;
        RECT 177.400 206.400 177.800 206.500 ;
        RECT 175.900 206.100 177.800 206.400 ;
        RECT 175.900 206.000 176.300 206.100 ;
        RECT 176.700 205.700 177.100 205.800 ;
        RECT 171.800 205.500 174.600 205.600 ;
        RECT 171.700 205.400 174.600 205.500 ;
        RECT 167.800 204.900 169.000 205.200 ;
        RECT 169.700 205.300 174.600 205.400 ;
        RECT 169.700 205.100 172.100 205.300 ;
        RECT 167.800 204.400 168.100 204.900 ;
        RECT 164.600 203.800 165.800 204.100 ;
        RECT 167.400 204.000 168.100 204.400 ;
        RECT 168.900 204.500 169.300 204.600 ;
        RECT 169.700 204.500 170.000 205.100 ;
        RECT 168.900 204.200 170.000 204.500 ;
        RECT 170.300 204.500 173.000 204.800 ;
        RECT 170.300 204.400 170.700 204.500 ;
        RECT 172.600 204.400 173.000 204.500 ;
        RECT 165.400 201.100 165.800 203.800 ;
        RECT 169.500 203.700 169.900 203.800 ;
        RECT 170.900 203.700 171.300 203.800 ;
        RECT 167.800 203.100 168.200 203.500 ;
        RECT 169.500 203.400 171.300 203.700 ;
        RECT 169.900 203.100 170.200 203.400 ;
        RECT 172.600 203.100 173.000 203.500 ;
        RECT 167.500 201.100 168.100 203.100 ;
        RECT 169.800 201.100 170.200 203.100 ;
        RECT 172.000 202.800 173.000 203.100 ;
        RECT 172.000 201.100 172.400 202.800 ;
        RECT 174.200 201.100 174.600 205.300 ;
        RECT 175.000 205.400 177.100 205.700 ;
        RECT 175.000 201.100 175.400 205.400 ;
        RECT 178.300 205.200 178.600 206.800 ;
        RECT 181.900 206.700 182.300 206.800 ;
        RECT 182.700 206.200 183.100 206.300 ;
        RECT 179.000 206.100 179.400 206.200 ;
        RECT 180.600 206.100 183.100 206.200 ;
        RECT 179.000 205.900 183.100 206.100 ;
        RECT 179.000 205.800 181.000 205.900 ;
        RECT 184.600 205.700 185.000 207.400 ;
        RECT 188.100 207.100 188.500 207.200 ;
        RECT 191.000 207.100 191.300 207.800 ;
        RECT 193.400 207.500 193.800 209.900 ;
        RECT 194.200 208.000 194.600 209.900 ;
        RECT 195.800 208.000 196.200 209.900 ;
        RECT 194.200 207.900 196.200 208.000 ;
        RECT 196.600 207.900 197.000 209.900 ;
        RECT 197.400 207.900 197.800 209.900 ;
        RECT 198.200 208.000 198.600 209.900 ;
        RECT 199.800 208.000 200.200 209.900 ;
        RECT 198.200 207.900 200.200 208.000 ;
        RECT 200.600 208.500 201.000 209.500 ;
        RECT 194.300 207.700 196.100 207.900 ;
        RECT 194.600 207.200 195.000 207.400 ;
        RECT 196.600 207.200 196.900 207.900 ;
        RECT 197.500 207.200 197.800 207.900 ;
        RECT 198.300 207.700 200.100 207.900 ;
        RECT 200.600 207.400 200.900 208.500 ;
        RECT 202.700 208.000 203.100 209.500 ;
        RECT 202.700 207.700 203.500 208.000 ;
        RECT 205.400 207.800 205.800 208.600 ;
        RECT 203.100 207.500 203.500 207.700 ;
        RECT 199.400 207.200 199.800 207.400 ;
        RECT 192.600 207.100 193.400 207.200 ;
        RECT 187.900 206.800 193.400 207.100 ;
        RECT 194.200 206.900 195.000 207.200 ;
        RECT 194.200 206.800 194.600 206.900 ;
        RECT 195.700 206.800 197.000 207.200 ;
        RECT 197.400 206.800 198.700 207.200 ;
        RECT 199.400 206.900 200.200 207.200 ;
        RECT 200.600 207.100 202.700 207.400 ;
        RECT 199.800 206.800 200.200 206.900 ;
        RECT 202.200 206.900 202.700 207.100 ;
        RECT 203.200 207.200 203.500 207.500 ;
        RECT 187.000 206.400 187.400 206.500 ;
        RECT 185.500 206.100 187.400 206.400 ;
        RECT 185.500 206.000 185.900 206.100 ;
        RECT 186.300 205.700 186.700 205.800 ;
        RECT 181.400 205.500 184.200 205.600 ;
        RECT 181.300 205.400 184.200 205.500 ;
        RECT 177.400 204.900 178.600 205.200 ;
        RECT 179.300 205.300 184.200 205.400 ;
        RECT 179.300 205.100 181.700 205.300 ;
        RECT 177.400 204.400 177.700 204.900 ;
        RECT 177.000 204.000 177.700 204.400 ;
        RECT 178.500 204.500 178.900 204.600 ;
        RECT 179.300 204.500 179.600 205.100 ;
        RECT 178.500 204.200 179.600 204.500 ;
        RECT 179.900 204.500 182.600 204.800 ;
        RECT 179.900 204.400 180.300 204.500 ;
        RECT 182.200 204.400 182.600 204.500 ;
        RECT 179.100 203.700 179.500 203.800 ;
        RECT 180.500 203.700 180.900 203.800 ;
        RECT 177.400 203.100 177.800 203.500 ;
        RECT 179.100 203.400 180.900 203.700 ;
        RECT 179.500 203.100 179.800 203.400 ;
        RECT 182.200 203.100 182.600 203.500 ;
        RECT 177.100 201.100 177.700 203.100 ;
        RECT 179.400 201.100 179.800 203.100 ;
        RECT 181.600 202.800 182.600 203.100 ;
        RECT 181.600 201.100 182.000 202.800 ;
        RECT 183.800 201.100 184.200 205.300 ;
        RECT 184.600 205.400 186.700 205.700 ;
        RECT 184.600 201.100 185.000 205.400 ;
        RECT 187.900 205.200 188.200 206.800 ;
        RECT 191.500 206.700 191.900 206.800 ;
        RECT 192.300 206.200 192.700 206.300 ;
        RECT 190.200 205.900 192.700 206.200 ;
        RECT 190.200 205.800 190.600 205.900 ;
        RECT 195.000 205.800 195.400 206.600 ;
        RECT 191.000 205.500 193.800 205.600 ;
        RECT 190.900 205.400 193.800 205.500 ;
        RECT 187.000 204.900 188.200 205.200 ;
        RECT 188.900 205.300 193.800 205.400 ;
        RECT 188.900 205.100 191.300 205.300 ;
        RECT 187.000 204.400 187.300 204.900 ;
        RECT 186.600 204.000 187.300 204.400 ;
        RECT 188.100 204.500 188.500 204.600 ;
        RECT 188.900 204.500 189.200 205.100 ;
        RECT 188.100 204.200 189.200 204.500 ;
        RECT 189.500 204.500 192.200 204.800 ;
        RECT 189.500 204.400 189.900 204.500 ;
        RECT 191.800 204.400 192.200 204.500 ;
        RECT 188.700 203.700 189.100 203.800 ;
        RECT 190.100 203.700 190.500 203.800 ;
        RECT 187.000 203.100 187.400 203.500 ;
        RECT 188.700 203.400 190.500 203.700 ;
        RECT 189.100 203.100 189.400 203.400 ;
        RECT 191.800 203.100 192.200 203.500 ;
        RECT 186.700 201.100 187.300 203.100 ;
        RECT 189.000 201.100 189.400 203.100 ;
        RECT 191.200 202.800 192.200 203.100 ;
        RECT 191.200 201.100 191.600 202.800 ;
        RECT 193.400 201.100 193.800 205.300 ;
        RECT 195.700 205.100 196.000 206.800 ;
        RECT 198.400 206.100 198.700 206.800 ;
        RECT 196.600 205.800 198.700 206.100 ;
        RECT 199.000 205.800 199.400 206.600 ;
        RECT 200.600 205.800 201.000 206.600 ;
        RECT 201.400 205.800 201.800 206.600 ;
        RECT 202.200 206.500 202.900 206.900 ;
        RECT 203.200 206.800 204.200 207.200 ;
        RECT 196.600 205.200 196.900 205.800 ;
        RECT 196.600 205.100 197.000 205.200 ;
        RECT 195.500 204.800 196.000 205.100 ;
        RECT 196.300 204.800 197.000 205.100 ;
        RECT 197.400 205.100 197.800 205.200 ;
        RECT 198.400 205.100 198.700 205.800 ;
        RECT 202.200 205.500 202.500 206.500 ;
        RECT 200.600 205.200 202.500 205.500 ;
        RECT 197.400 204.800 198.100 205.100 ;
        RECT 198.400 204.800 198.900 205.100 ;
        RECT 195.500 201.100 195.900 204.800 ;
        RECT 196.300 204.200 196.600 204.800 ;
        RECT 196.200 203.800 196.600 204.200 ;
        RECT 197.800 204.200 198.100 204.800 ;
        RECT 197.800 203.800 198.200 204.200 ;
        RECT 198.500 201.100 198.900 204.800 ;
        RECT 200.600 203.500 200.900 205.200 ;
        RECT 203.200 204.900 203.500 206.800 ;
        RECT 203.800 206.100 204.200 206.200 ;
        RECT 204.600 206.100 205.000 206.200 ;
        RECT 203.800 205.800 205.000 206.100 ;
        RECT 206.200 206.100 206.600 209.900 ;
        RECT 210.500 209.200 210.900 209.500 ;
        RECT 210.500 208.800 211.400 209.200 ;
        RECT 210.500 208.000 210.900 208.800 ;
        RECT 212.600 208.500 213.000 209.500 ;
        RECT 214.200 208.900 214.600 209.900 ;
        RECT 210.100 207.700 210.900 208.000 ;
        RECT 210.100 207.500 210.500 207.700 ;
        RECT 210.100 207.200 210.400 207.500 ;
        RECT 212.700 207.400 213.000 208.500 ;
        RECT 213.400 207.800 213.800 208.600 ;
        RECT 214.300 208.100 214.600 208.900 ;
        RECT 215.900 208.200 216.300 208.600 ;
        RECT 215.800 208.100 216.200 208.200 ;
        RECT 214.200 207.800 216.200 208.100 ;
        RECT 216.600 207.900 217.000 209.900 ;
        RECT 209.400 206.800 210.400 207.200 ;
        RECT 210.900 207.100 213.000 207.400 ;
        RECT 214.300 207.200 214.600 207.800 ;
        RECT 210.900 206.900 211.400 207.100 ;
        RECT 209.400 206.100 209.800 206.200 ;
        RECT 206.200 205.800 209.800 206.100 ;
        RECT 203.800 205.400 204.200 205.800 ;
        RECT 202.700 204.600 203.500 204.900 ;
        RECT 200.600 201.500 201.000 203.500 ;
        RECT 202.700 202.200 203.100 204.600 ;
        RECT 202.200 201.800 203.100 202.200 ;
        RECT 202.700 201.100 203.100 201.800 ;
        RECT 206.200 201.100 206.600 205.800 ;
        RECT 209.400 205.400 209.800 205.800 ;
        RECT 210.100 204.900 210.400 206.800 ;
        RECT 210.700 206.500 211.400 206.900 ;
        RECT 214.200 206.800 214.600 207.200 ;
        RECT 211.100 205.500 211.400 206.500 ;
        RECT 211.800 205.800 212.200 206.600 ;
        RECT 212.600 205.800 213.000 206.600 ;
        RECT 211.100 205.200 213.000 205.500 ;
        RECT 210.100 204.600 210.900 204.900 ;
        RECT 210.500 201.100 210.900 204.600 ;
        RECT 212.700 203.500 213.000 205.200 ;
        RECT 214.300 205.100 214.600 206.800 ;
        RECT 215.000 205.400 215.400 206.200 ;
        RECT 215.800 206.100 216.200 206.200 ;
        RECT 216.700 206.100 217.000 207.900 ;
        RECT 219.000 208.500 219.400 209.500 ;
        RECT 219.000 207.400 219.300 208.500 ;
        RECT 221.100 208.000 221.500 209.500 ;
        RECT 223.800 208.000 224.200 209.900 ;
        RECT 225.400 208.000 225.800 209.900 ;
        RECT 221.100 207.700 221.900 208.000 ;
        RECT 223.800 207.900 225.800 208.000 ;
        RECT 226.200 207.900 226.600 209.900 ;
        RECT 227.000 207.900 227.400 209.900 ;
        RECT 227.800 208.000 228.200 209.900 ;
        RECT 229.400 208.000 229.800 209.900 ;
        RECT 227.800 207.900 229.800 208.000 ;
        RECT 223.900 207.700 225.700 207.900 ;
        RECT 221.500 207.500 221.900 207.700 ;
        RECT 217.400 206.400 217.800 207.200 ;
        RECT 218.200 206.800 218.600 207.200 ;
        RECT 219.000 207.100 221.100 207.400 ;
        RECT 220.600 206.900 221.100 207.100 ;
        RECT 221.600 207.200 221.900 207.500 ;
        RECT 224.200 207.200 224.600 207.400 ;
        RECT 226.200 207.200 226.500 207.900 ;
        RECT 227.100 207.200 227.400 207.900 ;
        RECT 227.900 207.700 229.700 207.900 ;
        RECT 230.200 207.700 230.600 209.900 ;
        RECT 232.300 209.200 232.900 209.900 ;
        RECT 232.300 208.900 233.000 209.200 ;
        RECT 234.600 208.900 235.000 209.900 ;
        RECT 236.800 209.200 237.200 209.900 ;
        RECT 236.800 208.900 237.800 209.200 ;
        RECT 232.600 208.500 233.000 208.900 ;
        RECT 234.700 208.600 235.000 208.900 ;
        RECT 234.700 208.300 236.100 208.600 ;
        RECT 235.700 208.200 236.100 208.300 ;
        RECT 236.600 208.200 237.000 208.600 ;
        RECT 237.400 208.500 237.800 208.900 ;
        RECT 231.700 207.700 232.100 207.800 ;
        RECT 230.200 207.400 232.100 207.700 ;
        RECT 229.000 207.200 229.400 207.400 ;
        RECT 218.200 206.200 218.500 206.800 ;
        RECT 218.200 206.100 218.600 206.200 ;
        RECT 215.800 205.800 217.000 206.100 ;
        RECT 217.800 205.800 218.600 206.100 ;
        RECT 219.000 205.800 219.400 206.600 ;
        RECT 219.800 205.800 220.200 206.600 ;
        RECT 220.600 206.500 221.300 206.900 ;
        RECT 221.600 206.800 222.600 207.200 ;
        RECT 223.800 206.900 224.600 207.200 ;
        RECT 223.800 206.800 224.200 206.900 ;
        RECT 225.300 206.800 226.600 207.200 ;
        RECT 227.000 206.800 228.300 207.200 ;
        RECT 229.000 206.900 229.800 207.200 ;
        RECT 229.400 206.800 229.800 206.900 ;
        RECT 215.900 205.100 216.200 205.800 ;
        RECT 217.800 205.600 218.200 205.800 ;
        RECT 220.600 205.500 220.900 206.500 ;
        RECT 219.000 205.200 220.900 205.500 ;
        RECT 214.200 204.700 215.100 205.100 ;
        RECT 212.600 201.500 213.000 203.500 ;
        RECT 214.700 201.100 215.100 204.700 ;
        RECT 215.800 201.100 216.200 205.100 ;
        RECT 216.600 204.800 218.600 205.100 ;
        RECT 216.600 201.100 217.000 204.800 ;
        RECT 218.200 201.100 218.600 204.800 ;
        RECT 219.000 203.500 219.300 205.200 ;
        RECT 221.600 204.900 221.900 206.800 ;
        RECT 222.200 206.100 222.600 206.200 ;
        RECT 223.000 206.100 223.400 206.200 ;
        RECT 222.200 205.800 223.400 206.100 ;
        RECT 224.600 205.800 225.000 206.600 ;
        RECT 225.300 206.100 225.600 206.800 ;
        RECT 228.000 206.200 228.300 206.800 ;
        RECT 225.300 205.800 227.300 206.100 ;
        RECT 227.800 205.800 228.300 206.200 ;
        RECT 228.600 205.800 229.000 206.600 ;
        RECT 222.200 205.400 222.600 205.800 ;
        RECT 225.300 205.100 225.600 205.800 ;
        RECT 227.000 205.200 227.300 205.800 ;
        RECT 226.200 205.100 226.600 205.200 ;
        RECT 221.100 204.600 221.900 204.900 ;
        RECT 225.100 204.800 225.600 205.100 ;
        RECT 225.900 204.800 226.600 205.100 ;
        RECT 227.000 205.100 227.400 205.200 ;
        RECT 228.000 205.100 228.300 205.800 ;
        RECT 230.200 205.700 230.600 207.400 ;
        RECT 233.700 207.100 234.100 207.200 ;
        RECT 236.600 207.100 236.900 208.200 ;
        RECT 239.000 207.500 239.400 209.900 ;
        RECT 239.800 208.500 240.200 209.500 ;
        RECT 239.800 207.400 240.100 208.500 ;
        RECT 241.900 208.000 242.300 209.500 ;
        RECT 241.900 207.700 242.700 208.000 ;
        RECT 242.300 207.500 242.700 207.700 ;
        RECT 238.200 207.100 239.000 207.200 ;
        RECT 239.800 207.100 241.900 207.400 ;
        RECT 233.500 206.800 239.000 207.100 ;
        RECT 241.400 206.900 241.900 207.100 ;
        RECT 242.400 207.200 242.700 207.500 ;
        RECT 242.400 207.100 243.400 207.200 ;
        RECT 243.800 207.100 244.200 207.200 ;
        RECT 232.600 206.400 233.000 206.500 ;
        RECT 231.100 206.100 233.000 206.400 ;
        RECT 231.100 206.000 231.500 206.100 ;
        RECT 231.900 205.700 232.300 205.800 ;
        RECT 230.200 205.400 232.300 205.700 ;
        RECT 227.000 204.800 227.700 205.100 ;
        RECT 228.000 204.800 228.500 205.100 ;
        RECT 219.000 201.500 219.400 203.500 ;
        RECT 221.100 202.200 221.500 204.600 ;
        RECT 220.600 201.800 221.500 202.200 ;
        RECT 221.100 201.100 221.500 201.800 ;
        RECT 225.100 201.100 225.500 204.800 ;
        RECT 225.900 204.200 226.200 204.800 ;
        RECT 225.800 203.800 226.200 204.200 ;
        RECT 227.400 204.200 227.700 204.800 ;
        RECT 227.400 203.800 227.800 204.200 ;
        RECT 228.100 201.100 228.500 204.800 ;
        RECT 230.200 201.100 230.600 205.400 ;
        RECT 233.500 205.200 233.800 206.800 ;
        RECT 237.100 206.700 237.500 206.800 ;
        RECT 237.900 206.200 238.300 206.300 ;
        RECT 235.000 206.100 235.400 206.200 ;
        RECT 235.800 206.100 238.300 206.200 ;
        RECT 235.000 205.900 238.300 206.100 ;
        RECT 235.000 205.800 236.200 205.900 ;
        RECT 239.800 205.800 240.200 206.600 ;
        RECT 240.600 205.800 241.000 206.600 ;
        RECT 241.400 206.500 242.100 206.900 ;
        RECT 242.400 206.800 244.200 207.100 ;
        RECT 236.600 205.500 239.400 205.600 ;
        RECT 241.400 205.500 241.700 206.500 ;
        RECT 236.500 205.400 239.400 205.500 ;
        RECT 232.600 204.900 233.800 205.200 ;
        RECT 234.500 205.300 239.400 205.400 ;
        RECT 234.500 205.100 236.900 205.300 ;
        RECT 232.600 204.400 232.900 204.900 ;
        RECT 232.200 204.000 232.900 204.400 ;
        RECT 233.700 204.500 234.100 204.600 ;
        RECT 234.500 204.500 234.800 205.100 ;
        RECT 233.700 204.200 234.800 204.500 ;
        RECT 235.100 204.500 237.800 204.800 ;
        RECT 235.100 204.400 235.500 204.500 ;
        RECT 237.400 204.400 237.800 204.500 ;
        RECT 234.300 203.700 234.700 203.800 ;
        RECT 235.700 203.700 236.100 203.800 ;
        RECT 232.600 203.100 233.000 203.500 ;
        RECT 234.300 203.400 236.100 203.700 ;
        RECT 234.700 203.100 235.000 203.400 ;
        RECT 237.400 203.100 237.800 203.500 ;
        RECT 232.300 201.100 232.900 203.100 ;
        RECT 234.600 201.100 235.000 203.100 ;
        RECT 236.800 202.800 237.800 203.100 ;
        RECT 236.800 201.100 237.200 202.800 ;
        RECT 239.000 201.100 239.400 205.300 ;
        RECT 239.800 205.200 241.700 205.500 ;
        RECT 239.800 203.500 240.100 205.200 ;
        RECT 242.400 204.900 242.700 206.800 ;
        RECT 243.000 206.100 243.400 206.200 ;
        RECT 244.600 206.100 245.000 209.900 ;
        RECT 245.400 208.100 245.800 208.600 ;
        RECT 246.200 208.100 246.600 209.900 ;
        RECT 248.300 209.200 248.900 209.900 ;
        RECT 248.300 208.900 249.000 209.200 ;
        RECT 250.600 208.900 251.000 209.900 ;
        RECT 252.800 209.200 253.200 209.900 ;
        RECT 252.800 208.900 253.800 209.200 ;
        RECT 248.600 208.500 249.000 208.900 ;
        RECT 250.700 208.600 251.000 208.900 ;
        RECT 250.700 208.300 252.100 208.600 ;
        RECT 251.700 208.200 252.100 208.300 ;
        RECT 252.600 208.200 253.000 208.600 ;
        RECT 253.400 208.500 253.800 208.900 ;
        RECT 245.400 207.800 246.600 208.100 ;
        RECT 243.000 205.800 245.000 206.100 ;
        RECT 243.000 205.400 243.400 205.800 ;
        RECT 241.900 204.600 242.700 204.900 ;
        RECT 239.800 201.500 240.200 203.500 ;
        RECT 241.900 201.100 242.300 204.600 ;
        RECT 244.600 201.100 245.000 205.800 ;
        RECT 246.200 207.700 246.600 207.800 ;
        RECT 247.700 207.700 248.100 207.800 ;
        RECT 246.200 207.400 248.100 207.700 ;
        RECT 246.200 205.700 246.600 207.400 ;
        RECT 249.700 207.100 250.100 207.200 ;
        RECT 252.600 207.100 252.900 208.200 ;
        RECT 255.000 207.500 255.400 209.900 ;
        RECT 256.600 207.600 257.000 209.900 ;
        RECT 258.200 207.600 258.600 209.900 ;
        RECT 259.800 207.600 260.200 209.900 ;
        RECT 261.400 207.600 261.800 209.900 ;
        RECT 256.600 207.200 257.500 207.600 ;
        RECT 258.200 207.200 259.300 207.600 ;
        RECT 259.800 207.200 260.900 207.600 ;
        RECT 261.400 207.200 262.600 207.600 ;
        RECT 254.200 207.100 255.000 207.200 ;
        RECT 249.500 206.800 255.000 207.100 ;
        RECT 255.800 206.900 256.200 207.200 ;
        RECT 257.100 206.900 257.500 207.200 ;
        RECT 258.900 206.900 259.300 207.200 ;
        RECT 260.500 206.900 260.900 207.200 ;
        RECT 248.600 206.400 249.000 206.500 ;
        RECT 247.100 206.100 249.000 206.400 ;
        RECT 247.100 206.000 247.500 206.100 ;
        RECT 247.900 205.700 248.300 205.800 ;
        RECT 246.200 205.400 248.300 205.700 ;
        RECT 246.200 201.100 246.600 205.400 ;
        RECT 249.500 205.200 249.800 206.800 ;
        RECT 253.100 206.700 253.500 206.800 ;
        RECT 255.800 206.500 256.700 206.900 ;
        RECT 257.100 206.500 258.400 206.900 ;
        RECT 258.900 206.500 260.100 206.900 ;
        RECT 260.500 206.500 261.800 206.900 ;
        RECT 253.900 206.200 254.300 206.300 ;
        RECT 251.800 205.900 254.300 206.200 ;
        RECT 251.800 205.800 252.200 205.900 ;
        RECT 257.100 205.800 257.500 206.500 ;
        RECT 258.900 205.800 259.300 206.500 ;
        RECT 260.500 205.800 260.900 206.500 ;
        RECT 262.200 205.800 262.600 207.200 ;
        RECT 252.600 205.500 255.400 205.600 ;
        RECT 252.500 205.400 255.400 205.500 ;
        RECT 248.600 204.900 249.800 205.200 ;
        RECT 250.500 205.300 255.400 205.400 ;
        RECT 250.500 205.100 252.900 205.300 ;
        RECT 248.600 204.400 248.900 204.900 ;
        RECT 248.200 204.000 248.900 204.400 ;
        RECT 249.700 204.500 250.100 204.600 ;
        RECT 250.500 204.500 250.800 205.100 ;
        RECT 249.700 204.200 250.800 204.500 ;
        RECT 251.100 204.500 253.800 204.800 ;
        RECT 251.100 204.400 251.500 204.500 ;
        RECT 253.400 204.400 253.800 204.500 ;
        RECT 250.300 203.700 250.700 203.800 ;
        RECT 251.700 203.700 252.100 203.800 ;
        RECT 248.600 203.100 249.000 203.500 ;
        RECT 250.300 203.400 252.100 203.700 ;
        RECT 250.700 203.100 251.000 203.400 ;
        RECT 253.400 203.100 253.800 203.500 ;
        RECT 248.300 201.100 248.900 203.100 ;
        RECT 250.600 201.100 251.000 203.100 ;
        RECT 252.800 202.800 253.800 203.100 ;
        RECT 252.800 201.100 253.200 202.800 ;
        RECT 255.000 201.100 255.400 205.300 ;
        RECT 256.600 205.400 257.500 205.800 ;
        RECT 258.200 205.400 259.300 205.800 ;
        RECT 259.800 205.400 260.900 205.800 ;
        RECT 261.400 205.400 262.600 205.800 ;
        RECT 256.600 201.100 257.000 205.400 ;
        RECT 258.200 201.100 258.600 205.400 ;
        RECT 259.800 201.100 260.200 205.400 ;
        RECT 261.400 201.100 261.800 205.400 ;
        RECT 1.400 195.600 1.800 199.900 ;
        RECT 3.000 195.600 3.400 199.900 ;
        RECT 4.600 195.600 5.000 199.900 ;
        RECT 6.200 195.600 6.600 199.900 ;
        RECT 7.800 195.700 8.200 199.900 ;
        RECT 10.000 198.200 10.400 199.900 ;
        RECT 9.400 197.900 10.400 198.200 ;
        RECT 12.200 197.900 12.600 199.900 ;
        RECT 14.300 197.900 14.900 199.900 ;
        RECT 9.400 197.500 9.800 197.900 ;
        RECT 12.200 197.600 12.500 197.900 ;
        RECT 11.100 197.300 12.900 197.600 ;
        RECT 14.200 197.500 14.600 197.900 ;
        RECT 11.100 197.200 11.500 197.300 ;
        RECT 12.500 197.200 12.900 197.300 ;
        RECT 9.400 196.500 9.800 196.600 ;
        RECT 11.700 196.500 12.100 196.600 ;
        RECT 9.400 196.200 12.100 196.500 ;
        RECT 12.400 196.500 13.500 196.800 ;
        RECT 12.400 195.900 12.700 196.500 ;
        RECT 13.100 196.400 13.500 196.500 ;
        RECT 14.300 196.600 15.000 197.000 ;
        RECT 14.300 196.100 14.600 196.600 ;
        RECT 10.300 195.700 12.700 195.900 ;
        RECT 7.800 195.600 12.700 195.700 ;
        RECT 13.400 195.800 14.600 196.100 ;
        RECT 1.400 195.200 2.300 195.600 ;
        RECT 3.000 195.200 4.100 195.600 ;
        RECT 4.600 195.200 5.700 195.600 ;
        RECT 6.200 195.200 7.400 195.600 ;
        RECT 7.800 195.500 10.700 195.600 ;
        RECT 7.800 195.400 10.600 195.500 ;
        RECT 0.600 194.800 1.000 195.200 ;
        RECT 0.600 194.500 0.900 194.800 ;
        RECT 1.900 194.500 2.300 195.200 ;
        RECT 3.700 194.500 4.100 195.200 ;
        RECT 5.300 194.500 5.700 195.200 ;
        RECT 0.600 194.100 1.500 194.500 ;
        RECT 1.900 194.100 3.200 194.500 ;
        RECT 3.700 194.100 4.900 194.500 ;
        RECT 5.300 194.100 6.600 194.500 ;
        RECT 0.600 193.800 1.000 194.100 ;
        RECT 1.900 193.800 2.300 194.100 ;
        RECT 3.700 193.800 4.100 194.100 ;
        RECT 5.300 193.800 5.700 194.100 ;
        RECT 7.000 193.800 7.400 195.200 ;
        RECT 11.000 195.100 11.400 195.200 ;
        RECT 8.900 194.800 11.400 195.100 ;
        RECT 8.900 194.700 9.300 194.800 ;
        RECT 9.700 194.200 10.100 194.300 ;
        RECT 13.400 194.200 13.700 195.800 ;
        RECT 16.600 195.600 17.000 199.900 ;
        RECT 18.700 196.300 19.100 199.900 ;
        RECT 18.200 195.900 19.100 196.300 ;
        RECT 19.800 195.900 20.200 199.900 ;
        RECT 20.600 196.200 21.000 199.900 ;
        RECT 22.200 196.200 22.600 199.900 ;
        RECT 20.600 195.900 22.600 196.200 ;
        RECT 14.900 195.300 17.000 195.600 ;
        RECT 14.900 195.200 15.300 195.300 ;
        RECT 15.700 194.900 16.100 195.000 ;
        RECT 14.200 194.600 16.100 194.900 ;
        RECT 14.200 194.500 14.600 194.600 ;
        RECT 8.200 193.900 13.700 194.200 ;
        RECT 8.200 193.800 9.000 193.900 ;
        RECT 1.400 193.400 2.300 193.800 ;
        RECT 3.000 193.400 4.100 193.800 ;
        RECT 4.600 193.400 5.700 193.800 ;
        RECT 6.200 193.400 7.400 193.800 ;
        RECT 1.400 191.100 1.800 193.400 ;
        RECT 3.000 191.100 3.400 193.400 ;
        RECT 4.600 191.100 5.000 193.400 ;
        RECT 6.200 191.100 6.600 193.400 ;
        RECT 7.800 191.100 8.200 193.500 ;
        RECT 10.300 192.800 10.600 193.900 ;
        RECT 13.100 193.800 13.500 193.900 ;
        RECT 16.600 193.600 17.000 195.300 ;
        RECT 18.300 194.200 18.600 195.900 ;
        RECT 19.000 194.800 19.400 195.600 ;
        RECT 19.900 195.200 20.200 195.900 ;
        RECT 21.800 195.200 22.200 195.400 ;
        RECT 19.800 194.900 21.000 195.200 ;
        RECT 21.800 194.900 22.600 195.200 ;
        RECT 19.800 194.800 20.200 194.900 ;
        RECT 18.200 193.800 18.600 194.200 ;
        RECT 19.800 194.200 20.100 194.800 ;
        RECT 19.800 193.800 20.200 194.200 ;
        RECT 15.000 193.300 17.000 193.600 ;
        RECT 15.000 193.200 15.500 193.300 ;
        RECT 15.000 192.800 15.400 193.200 ;
        RECT 16.600 193.100 17.000 193.300 ;
        RECT 17.400 193.100 17.800 193.200 ;
        RECT 18.300 193.100 18.600 193.800 ;
        RECT 19.800 193.100 20.200 193.200 ;
        RECT 20.700 193.100 21.000 194.900 ;
        RECT 22.200 194.800 22.600 194.900 ;
        RECT 23.800 195.100 24.200 199.900 ;
        RECT 25.800 196.800 26.200 197.200 ;
        RECT 24.600 195.800 25.000 196.600 ;
        RECT 25.800 196.200 26.100 196.800 ;
        RECT 26.500 196.200 26.900 199.900 ;
        RECT 25.400 195.900 26.100 196.200 ;
        RECT 25.400 195.800 25.800 195.900 ;
        RECT 26.400 195.800 27.400 196.200 ;
        RECT 25.400 195.100 25.700 195.800 ;
        RECT 23.800 194.800 25.700 195.100 ;
        RECT 21.400 193.800 21.800 194.600 ;
        RECT 23.000 193.400 23.400 194.200 ;
        RECT 16.600 192.800 17.800 193.100 ;
        RECT 18.200 192.800 20.200 193.100 ;
        RECT 9.400 192.100 9.800 192.500 ;
        RECT 10.200 192.400 10.600 192.800 ;
        RECT 11.100 192.700 11.500 192.800 ;
        RECT 11.100 192.400 12.500 192.700 ;
        RECT 12.200 192.100 12.500 192.400 ;
        RECT 14.200 192.100 14.600 192.500 ;
        RECT 9.400 191.800 10.400 192.100 ;
        RECT 10.000 191.100 10.400 191.800 ;
        RECT 12.200 191.100 12.600 192.100 ;
        RECT 14.200 191.800 14.900 192.100 ;
        RECT 14.300 191.100 14.900 191.800 ;
        RECT 16.600 191.100 17.000 192.800 ;
        RECT 17.400 192.400 17.800 192.800 ;
        RECT 18.300 192.100 18.600 192.800 ;
        RECT 19.900 192.400 20.300 192.800 ;
        RECT 18.200 191.100 18.600 192.100 ;
        RECT 20.600 191.100 21.000 193.100 ;
        RECT 23.800 193.100 24.200 194.800 ;
        RECT 26.400 194.200 26.700 195.800 ;
        RECT 28.600 195.600 29.000 199.900 ;
        RECT 30.700 197.900 31.300 199.900 ;
        RECT 33.000 197.900 33.400 199.900 ;
        RECT 35.200 198.200 35.600 199.900 ;
        RECT 35.200 197.900 36.200 198.200 ;
        RECT 31.000 197.500 31.400 197.900 ;
        RECT 33.100 197.600 33.400 197.900 ;
        RECT 32.700 197.300 34.500 197.600 ;
        RECT 35.800 197.500 36.200 197.900 ;
        RECT 32.700 197.200 33.100 197.300 ;
        RECT 34.100 197.200 34.500 197.300 ;
        RECT 30.600 196.600 31.300 197.000 ;
        RECT 31.000 196.100 31.300 196.600 ;
        RECT 32.100 196.500 33.200 196.800 ;
        RECT 32.100 196.400 32.500 196.500 ;
        RECT 31.000 195.800 32.200 196.100 ;
        RECT 28.600 195.300 30.700 195.600 ;
        RECT 27.000 194.400 27.400 195.200 ;
        RECT 25.400 193.800 26.700 194.200 ;
        RECT 27.800 194.100 28.200 194.200 ;
        RECT 27.400 193.800 28.200 194.100 ;
        RECT 25.500 193.100 25.800 193.800 ;
        RECT 27.400 193.600 27.800 193.800 ;
        RECT 28.600 193.600 29.000 195.300 ;
        RECT 30.300 195.200 30.700 195.300 ;
        RECT 29.500 194.900 29.900 195.000 ;
        RECT 29.500 194.600 31.400 194.900 ;
        RECT 31.000 194.500 31.400 194.600 ;
        RECT 31.900 194.200 32.200 195.800 ;
        RECT 32.900 195.900 33.200 196.500 ;
        RECT 33.500 196.500 33.900 196.600 ;
        RECT 35.800 196.500 36.200 196.600 ;
        RECT 33.500 196.200 36.200 196.500 ;
        RECT 32.900 195.700 35.300 195.900 ;
        RECT 37.400 195.700 37.800 199.900 ;
        RECT 32.900 195.600 37.800 195.700 ;
        RECT 34.900 195.500 37.800 195.600 ;
        RECT 35.000 195.400 37.800 195.500 ;
        RECT 38.200 195.700 38.600 199.900 ;
        RECT 40.400 198.200 40.800 199.900 ;
        RECT 39.800 197.900 40.800 198.200 ;
        RECT 42.600 197.900 43.000 199.900 ;
        RECT 44.700 197.900 45.300 199.900 ;
        RECT 39.800 197.500 40.200 197.900 ;
        RECT 42.600 197.600 42.900 197.900 ;
        RECT 41.500 197.300 43.300 197.600 ;
        RECT 44.600 197.500 45.000 197.900 ;
        RECT 41.500 197.200 41.900 197.300 ;
        RECT 42.900 197.200 43.300 197.300 ;
        RECT 39.800 196.500 40.200 196.600 ;
        RECT 42.100 196.500 42.500 196.600 ;
        RECT 39.800 196.200 42.500 196.500 ;
        RECT 42.800 196.500 43.900 196.800 ;
        RECT 42.800 195.900 43.100 196.500 ;
        RECT 43.500 196.400 43.900 196.500 ;
        RECT 44.700 196.600 45.400 197.000 ;
        RECT 44.700 196.100 45.000 196.600 ;
        RECT 40.700 195.700 43.100 195.900 ;
        RECT 38.200 195.600 43.100 195.700 ;
        RECT 43.800 195.800 45.000 196.100 ;
        RECT 38.200 195.500 41.100 195.600 ;
        RECT 38.200 195.400 41.000 195.500 ;
        RECT 34.200 195.100 34.600 195.200 ;
        RECT 41.400 195.100 41.800 195.200 ;
        RECT 34.200 194.800 36.700 195.100 ;
        RECT 36.300 194.700 36.700 194.800 ;
        RECT 39.300 194.800 41.800 195.100 ;
        RECT 39.300 194.700 39.700 194.800 ;
        RECT 35.500 194.200 35.900 194.300 ;
        RECT 40.100 194.200 40.500 194.300 ;
        RECT 43.800 194.200 44.100 195.800 ;
        RECT 47.000 195.600 47.400 199.900 ;
        RECT 48.200 196.800 48.600 197.200 ;
        RECT 48.200 196.200 48.500 196.800 ;
        RECT 48.900 196.200 49.300 199.900 ;
        RECT 47.800 195.900 48.500 196.200 ;
        RECT 48.800 195.900 49.300 196.200 ;
        RECT 47.800 195.800 48.200 195.900 ;
        RECT 45.300 195.300 47.400 195.600 ;
        RECT 45.300 195.200 45.700 195.300 ;
        RECT 46.100 194.900 46.500 195.000 ;
        RECT 44.600 194.600 46.500 194.900 ;
        RECT 44.600 194.500 45.000 194.600 ;
        RECT 31.900 193.900 37.400 194.200 ;
        RECT 32.100 193.800 32.500 193.900 ;
        RECT 28.600 193.300 30.500 193.600 ;
        RECT 26.300 193.100 28.100 193.300 ;
        RECT 23.800 192.800 24.700 193.100 ;
        RECT 24.300 191.100 24.700 192.800 ;
        RECT 25.400 191.100 25.800 193.100 ;
        RECT 26.200 193.000 28.200 193.100 ;
        RECT 26.200 191.100 26.600 193.000 ;
        RECT 27.800 191.100 28.200 193.000 ;
        RECT 28.600 191.100 29.000 193.300 ;
        RECT 30.100 193.200 30.500 193.300 ;
        RECT 35.000 192.800 35.300 193.900 ;
        RECT 36.600 193.800 37.400 193.900 ;
        RECT 38.600 193.900 44.100 194.200 ;
        RECT 38.600 193.800 39.400 193.900 ;
        RECT 34.100 192.700 34.500 192.800 ;
        RECT 31.000 192.100 31.400 192.500 ;
        RECT 33.100 192.400 34.500 192.700 ;
        RECT 35.000 192.400 35.400 192.800 ;
        RECT 33.100 192.100 33.400 192.400 ;
        RECT 35.800 192.100 36.200 192.500 ;
        RECT 30.700 191.800 31.400 192.100 ;
        RECT 30.700 191.100 31.300 191.800 ;
        RECT 33.000 191.100 33.400 192.100 ;
        RECT 35.200 191.800 36.200 192.100 ;
        RECT 35.200 191.100 35.600 191.800 ;
        RECT 37.400 191.100 37.800 193.500 ;
        RECT 38.200 191.100 38.600 193.500 ;
        RECT 40.700 192.800 41.000 193.900 ;
        RECT 43.500 193.800 43.900 193.900 ;
        RECT 47.000 193.600 47.400 195.300 ;
        RECT 48.800 194.200 49.100 195.900 ;
        RECT 52.600 195.600 53.000 199.900 ;
        RECT 54.700 197.900 55.300 199.900 ;
        RECT 57.000 197.900 57.400 199.900 ;
        RECT 59.200 198.200 59.600 199.900 ;
        RECT 59.200 197.900 60.200 198.200 ;
        RECT 55.000 197.500 55.400 197.900 ;
        RECT 57.100 197.600 57.400 197.900 ;
        RECT 56.700 197.300 58.500 197.600 ;
        RECT 59.800 197.500 60.200 197.900 ;
        RECT 56.700 197.200 57.100 197.300 ;
        RECT 58.100 197.200 58.500 197.300 ;
        RECT 54.600 196.600 55.300 197.000 ;
        RECT 55.000 196.100 55.300 196.600 ;
        RECT 56.100 196.500 57.200 196.800 ;
        RECT 56.100 196.400 56.500 196.500 ;
        RECT 55.000 195.800 56.200 196.100 ;
        RECT 52.600 195.300 54.700 195.600 ;
        RECT 49.400 195.100 49.800 195.200 ;
        RECT 51.800 195.100 52.200 195.200 ;
        RECT 49.400 194.800 52.200 195.100 ;
        RECT 49.400 194.400 49.800 194.800 ;
        RECT 47.800 193.800 49.100 194.200 ;
        RECT 50.200 194.100 50.600 194.200 ;
        RECT 51.000 194.100 51.400 194.200 ;
        RECT 49.800 193.800 51.400 194.100 ;
        RECT 45.500 193.300 47.400 193.600 ;
        RECT 45.500 193.200 45.900 193.300 ;
        RECT 39.800 192.100 40.200 192.500 ;
        RECT 40.600 192.400 41.000 192.800 ;
        RECT 41.500 192.700 41.900 192.800 ;
        RECT 41.500 192.400 42.900 192.700 ;
        RECT 42.600 192.100 42.900 192.400 ;
        RECT 44.600 192.100 45.000 192.500 ;
        RECT 39.800 191.800 40.800 192.100 ;
        RECT 40.400 191.100 40.800 191.800 ;
        RECT 42.600 191.100 43.000 192.100 ;
        RECT 44.600 191.800 45.300 192.100 ;
        RECT 44.700 191.100 45.300 191.800 ;
        RECT 47.000 191.100 47.400 193.300 ;
        RECT 47.900 193.100 48.200 193.800 ;
        RECT 49.800 193.600 50.200 193.800 ;
        RECT 52.600 193.600 53.000 195.300 ;
        RECT 54.300 195.200 54.700 195.300 ;
        RECT 53.500 194.900 53.900 195.000 ;
        RECT 53.500 194.600 55.400 194.900 ;
        RECT 55.000 194.500 55.400 194.600 ;
        RECT 55.900 194.200 56.200 195.800 ;
        RECT 56.900 195.900 57.200 196.500 ;
        RECT 57.500 196.500 57.900 196.600 ;
        RECT 59.800 196.500 60.200 196.600 ;
        RECT 57.500 196.200 60.200 196.500 ;
        RECT 56.900 195.700 59.300 195.900 ;
        RECT 61.400 195.700 61.800 199.900 ;
        RECT 62.200 196.200 62.600 199.900 ;
        RECT 63.800 196.200 64.200 199.900 ;
        RECT 62.200 195.900 64.200 196.200 ;
        RECT 64.600 195.900 65.000 199.900 ;
        RECT 66.700 196.300 67.100 199.900 ;
        RECT 66.200 195.900 67.100 196.300 ;
        RECT 68.200 196.800 68.600 197.200 ;
        RECT 68.200 196.200 68.500 196.800 ;
        RECT 68.900 196.200 69.300 199.900 ;
        RECT 67.800 195.900 68.500 196.200 ;
        RECT 68.800 195.900 69.300 196.200 ;
        RECT 56.900 195.600 61.800 195.700 ;
        RECT 58.900 195.500 61.800 195.600 ;
        RECT 59.000 195.400 61.800 195.500 ;
        RECT 62.600 195.200 63.000 195.400 ;
        RECT 64.600 195.200 64.900 195.900 ;
        RECT 57.400 195.100 57.800 195.200 ;
        RECT 58.200 195.100 58.600 195.200 ;
        RECT 57.400 194.800 60.700 195.100 ;
        RECT 62.200 194.900 63.000 195.200 ;
        RECT 63.800 194.900 65.000 195.200 ;
        RECT 62.200 194.800 62.600 194.900 ;
        RECT 63.800 194.800 64.200 194.900 ;
        RECT 64.600 194.800 65.000 194.900 ;
        RECT 60.300 194.700 60.700 194.800 ;
        RECT 59.500 194.200 59.900 194.300 ;
        RECT 55.900 193.900 61.400 194.200 ;
        RECT 56.100 193.800 56.500 193.900 ;
        RECT 58.200 193.800 58.600 193.900 ;
        RECT 52.600 193.300 54.500 193.600 ;
        RECT 48.700 193.100 50.500 193.300 ;
        RECT 47.800 191.100 48.200 193.100 ;
        RECT 48.600 193.000 50.600 193.100 ;
        RECT 48.600 191.100 49.000 193.000 ;
        RECT 50.200 191.100 50.600 193.000 ;
        RECT 52.600 191.100 53.000 193.300 ;
        RECT 54.100 193.200 54.500 193.300 ;
        RECT 59.000 192.800 59.300 193.900 ;
        RECT 60.600 193.800 61.400 193.900 ;
        RECT 63.000 193.800 63.400 194.600 ;
        RECT 58.100 192.700 58.500 192.800 ;
        RECT 55.000 192.100 55.400 192.500 ;
        RECT 57.100 192.400 58.500 192.700 ;
        RECT 59.000 192.400 59.400 192.800 ;
        RECT 57.100 192.100 57.400 192.400 ;
        RECT 59.800 192.100 60.200 192.500 ;
        RECT 54.700 191.800 55.400 192.100 ;
        RECT 54.700 191.100 55.300 191.800 ;
        RECT 57.000 191.100 57.400 192.100 ;
        RECT 59.200 191.800 60.200 192.100 ;
        RECT 59.200 191.100 59.600 191.800 ;
        RECT 61.400 191.100 61.800 193.500 ;
        RECT 63.800 193.100 64.100 194.800 ;
        RECT 66.300 194.200 66.600 195.900 ;
        RECT 67.800 195.800 68.200 195.900 ;
        RECT 67.000 194.800 67.400 195.600 ;
        RECT 68.800 195.200 69.100 195.900 ;
        RECT 71.000 195.600 71.400 199.900 ;
        RECT 73.100 197.900 73.700 199.900 ;
        RECT 75.400 197.900 75.800 199.900 ;
        RECT 77.600 198.200 78.000 199.900 ;
        RECT 77.600 197.900 78.600 198.200 ;
        RECT 73.400 197.500 73.800 197.900 ;
        RECT 75.500 197.600 75.800 197.900 ;
        RECT 75.100 197.300 76.900 197.600 ;
        RECT 78.200 197.500 78.600 197.900 ;
        RECT 75.100 197.200 75.500 197.300 ;
        RECT 76.500 197.200 76.900 197.300 ;
        RECT 73.000 196.600 73.700 197.000 ;
        RECT 73.400 196.100 73.700 196.600 ;
        RECT 74.500 196.500 75.600 196.800 ;
        RECT 74.500 196.400 74.900 196.500 ;
        RECT 73.400 195.800 74.600 196.100 ;
        RECT 71.000 195.300 73.100 195.600 ;
        RECT 68.600 194.800 69.100 195.200 ;
        RECT 68.800 194.200 69.100 194.800 ;
        RECT 69.400 194.400 69.800 195.200 ;
        RECT 66.200 194.100 66.600 194.200 ;
        RECT 64.600 193.800 66.600 194.100 ;
        RECT 67.800 193.800 69.100 194.200 ;
        RECT 70.200 194.100 70.600 194.200 ;
        RECT 69.800 193.800 70.600 194.100 ;
        RECT 64.600 193.200 64.900 193.800 ;
        RECT 63.800 191.100 64.200 193.100 ;
        RECT 64.600 192.800 65.000 193.200 ;
        RECT 64.500 192.400 64.900 192.800 ;
        RECT 65.400 192.400 65.800 193.200 ;
        RECT 66.300 192.100 66.600 193.800 ;
        RECT 67.900 193.100 68.200 193.800 ;
        RECT 69.800 193.600 70.200 193.800 ;
        RECT 71.000 193.600 71.400 195.300 ;
        RECT 72.700 195.200 73.100 195.300 ;
        RECT 71.900 194.900 72.300 195.000 ;
        RECT 71.900 194.600 73.800 194.900 ;
        RECT 73.400 194.500 73.800 194.600 ;
        RECT 74.300 194.200 74.600 195.800 ;
        RECT 75.300 195.900 75.600 196.500 ;
        RECT 75.900 196.500 76.300 196.600 ;
        RECT 78.200 196.500 78.600 196.600 ;
        RECT 75.900 196.200 78.600 196.500 ;
        RECT 75.300 195.700 77.700 195.900 ;
        RECT 79.800 195.700 80.200 199.900 ;
        RECT 75.300 195.600 80.200 195.700 ;
        RECT 77.300 195.500 80.200 195.600 ;
        RECT 80.600 197.500 81.000 199.500 ;
        RECT 80.600 195.800 80.900 197.500 ;
        RECT 82.700 196.400 83.100 199.900 ;
        RECT 82.700 196.100 83.500 196.400 ;
        RECT 80.600 195.500 82.500 195.800 ;
        RECT 77.400 195.400 80.200 195.500 ;
        RECT 76.600 195.100 77.000 195.200 ;
        RECT 76.600 194.800 79.100 195.100 ;
        RECT 78.700 194.700 79.100 194.800 ;
        RECT 80.600 194.400 81.000 195.200 ;
        RECT 81.400 194.400 81.800 195.200 ;
        RECT 82.200 194.500 82.500 195.500 ;
        RECT 77.900 194.200 78.300 194.300 ;
        RECT 74.300 193.900 79.800 194.200 ;
        RECT 82.200 194.100 82.900 194.500 ;
        RECT 83.200 194.200 83.500 196.100 ;
        RECT 85.400 195.800 85.800 196.600 ;
        RECT 83.800 194.800 84.200 195.600 ;
        RECT 82.200 193.900 82.700 194.100 ;
        RECT 74.500 193.800 74.900 193.900 ;
        RECT 77.400 193.800 77.800 193.900 ;
        RECT 79.000 193.800 79.800 193.900 ;
        RECT 71.000 193.300 72.900 193.600 ;
        RECT 68.700 193.100 70.500 193.300 ;
        RECT 66.200 191.100 66.600 192.100 ;
        RECT 67.800 191.100 68.200 193.100 ;
        RECT 68.600 193.000 70.600 193.100 ;
        RECT 68.600 191.100 69.000 193.000 ;
        RECT 70.200 191.100 70.600 193.000 ;
        RECT 71.000 191.100 71.400 193.300 ;
        RECT 72.500 193.200 72.900 193.300 ;
        RECT 77.400 192.800 77.700 193.800 ;
        RECT 80.600 193.600 82.700 193.900 ;
        RECT 83.200 193.800 84.200 194.200 ;
        RECT 76.500 192.700 76.900 192.800 ;
        RECT 73.400 192.100 73.800 192.500 ;
        RECT 75.500 192.400 76.900 192.700 ;
        RECT 77.400 192.400 77.800 192.800 ;
        RECT 75.500 192.100 75.800 192.400 ;
        RECT 78.200 192.100 78.600 192.500 ;
        RECT 73.100 191.800 73.800 192.100 ;
        RECT 73.100 191.100 73.700 191.800 ;
        RECT 75.400 191.100 75.800 192.100 ;
        RECT 77.600 191.800 78.600 192.100 ;
        RECT 77.600 191.100 78.000 191.800 ;
        RECT 79.800 191.100 80.200 193.500 ;
        RECT 80.600 192.500 80.900 193.600 ;
        RECT 83.200 193.500 83.500 193.800 ;
        RECT 83.100 193.300 83.500 193.500 ;
        RECT 82.700 193.000 83.500 193.300 ;
        RECT 86.200 193.100 86.600 199.900 ;
        RECT 87.800 197.500 88.200 199.500 ;
        RECT 87.800 195.800 88.100 197.500 ;
        RECT 89.900 196.400 90.300 199.900 ;
        RECT 89.900 196.100 90.700 196.400 ;
        RECT 87.800 195.500 89.700 195.800 ;
        RECT 87.800 194.400 88.200 195.200 ;
        RECT 88.600 194.400 89.000 195.200 ;
        RECT 89.400 194.500 89.700 195.500 ;
        RECT 87.000 193.400 87.400 194.200 ;
        RECT 89.400 194.100 90.100 194.500 ;
        RECT 90.400 194.200 90.700 196.100 ;
        RECT 91.000 195.100 91.400 195.600 ;
        RECT 92.600 195.100 93.000 199.900 ;
        RECT 91.000 194.800 93.000 195.100 ;
        RECT 90.400 194.100 91.400 194.200 ;
        RECT 91.800 194.100 92.200 194.200 ;
        RECT 89.400 193.900 89.900 194.100 ;
        RECT 87.800 193.600 89.900 193.900 ;
        RECT 90.400 193.800 92.200 194.100 ;
        RECT 80.600 191.500 81.000 192.500 ;
        RECT 82.700 192.200 83.100 193.000 ;
        RECT 85.700 192.800 86.600 193.100 ;
        RECT 82.700 191.800 83.400 192.200 ;
        RECT 82.700 191.500 83.100 191.800 ;
        RECT 85.700 191.100 86.100 192.800 ;
        RECT 87.800 192.500 88.100 193.600 ;
        RECT 90.400 193.500 90.700 193.800 ;
        RECT 90.300 193.300 90.700 193.500 ;
        RECT 89.900 193.000 90.700 193.300 ;
        RECT 87.800 191.500 88.200 192.500 ;
        RECT 89.900 191.500 90.300 193.000 ;
        RECT 92.600 191.100 93.000 194.800 ;
        RECT 94.200 195.600 94.600 199.900 ;
        RECT 96.300 197.900 96.900 199.900 ;
        RECT 98.600 197.900 99.000 199.900 ;
        RECT 100.800 198.200 101.200 199.900 ;
        RECT 100.800 197.900 101.800 198.200 ;
        RECT 96.600 197.500 97.000 197.900 ;
        RECT 98.700 197.600 99.000 197.900 ;
        RECT 98.300 197.300 100.100 197.600 ;
        RECT 101.400 197.500 101.800 197.900 ;
        RECT 98.300 197.200 98.700 197.300 ;
        RECT 99.700 197.200 100.100 197.300 ;
        RECT 96.200 196.600 96.900 197.000 ;
        RECT 95.800 195.600 96.200 196.200 ;
        RECT 96.600 196.100 96.900 196.600 ;
        RECT 97.700 196.500 98.800 196.800 ;
        RECT 97.700 196.400 98.100 196.500 ;
        RECT 96.600 195.800 97.800 196.100 ;
        RECT 94.200 195.300 96.300 195.600 ;
        RECT 94.200 193.600 94.600 195.300 ;
        RECT 95.900 195.200 96.300 195.300 ;
        RECT 95.100 194.900 95.500 195.000 ;
        RECT 95.100 194.600 97.000 194.900 ;
        RECT 96.600 194.500 97.000 194.600 ;
        RECT 97.500 194.200 97.800 195.800 ;
        RECT 98.500 195.900 98.800 196.500 ;
        RECT 99.100 196.500 99.500 196.600 ;
        RECT 101.400 196.500 101.800 196.600 ;
        RECT 99.100 196.200 101.800 196.500 ;
        RECT 98.500 195.700 100.900 195.900 ;
        RECT 103.000 195.700 103.400 199.900 ;
        RECT 104.600 196.400 105.000 199.900 ;
        RECT 98.500 195.600 103.400 195.700 ;
        RECT 100.500 195.500 103.400 195.600 ;
        RECT 100.600 195.400 103.400 195.500 ;
        RECT 104.500 195.900 105.000 196.400 ;
        RECT 106.200 196.200 106.600 199.900 ;
        RECT 105.300 195.900 106.600 196.200 ;
        RECT 99.800 195.100 100.200 195.200 ;
        RECT 99.800 194.800 102.300 195.100 ;
        RECT 101.900 194.700 102.300 194.800 ;
        RECT 101.100 194.200 101.500 194.300 ;
        RECT 104.500 194.200 104.800 195.900 ;
        RECT 105.300 194.900 105.600 195.900 ;
        RECT 108.600 195.600 109.000 199.900 ;
        RECT 110.700 197.900 111.300 199.900 ;
        RECT 113.000 197.900 113.400 199.900 ;
        RECT 115.200 198.200 115.600 199.900 ;
        RECT 115.200 197.900 116.200 198.200 ;
        RECT 111.000 197.500 111.400 197.900 ;
        RECT 113.100 197.600 113.400 197.900 ;
        RECT 112.700 197.300 114.500 197.600 ;
        RECT 115.800 197.500 116.200 197.900 ;
        RECT 112.700 197.200 113.100 197.300 ;
        RECT 114.100 197.200 114.500 197.300 ;
        RECT 110.200 197.000 110.900 197.200 ;
        RECT 110.200 196.800 111.300 197.000 ;
        RECT 110.600 196.600 111.300 196.800 ;
        RECT 111.000 196.100 111.300 196.600 ;
        RECT 112.100 196.500 113.200 196.800 ;
        RECT 112.100 196.400 112.500 196.500 ;
        RECT 111.000 195.800 112.200 196.100 ;
        RECT 108.600 195.300 110.700 195.600 ;
        RECT 105.100 194.500 105.600 194.900 ;
        RECT 97.500 193.900 103.000 194.200 ;
        RECT 97.700 193.800 98.100 193.900 ;
        RECT 100.600 193.800 101.000 193.900 ;
        RECT 102.200 193.800 103.000 193.900 ;
        RECT 104.500 193.800 105.000 194.200 ;
        RECT 94.200 193.300 96.100 193.600 ;
        RECT 93.400 193.100 93.800 193.200 ;
        RECT 94.200 193.100 94.600 193.300 ;
        RECT 95.700 193.200 96.100 193.300 ;
        RECT 93.400 192.800 94.600 193.100 ;
        RECT 100.600 192.800 100.900 193.800 ;
        RECT 93.400 192.400 93.800 192.800 ;
        RECT 94.200 191.100 94.600 192.800 ;
        RECT 99.700 192.700 100.100 192.800 ;
        RECT 96.600 192.100 97.000 192.500 ;
        RECT 98.700 192.400 100.100 192.700 ;
        RECT 100.600 192.400 101.000 192.800 ;
        RECT 98.700 192.100 99.000 192.400 ;
        RECT 101.400 192.100 101.800 192.500 ;
        RECT 96.300 191.800 97.000 192.100 ;
        RECT 96.300 191.100 96.900 191.800 ;
        RECT 98.600 191.100 99.000 192.100 ;
        RECT 100.800 191.800 101.800 192.100 ;
        RECT 100.800 191.100 101.200 191.800 ;
        RECT 103.000 191.100 103.400 193.500 ;
        RECT 104.500 193.100 104.800 193.800 ;
        RECT 105.300 193.700 105.600 194.500 ;
        RECT 106.100 195.100 106.600 195.200 ;
        RECT 107.800 195.100 108.200 195.200 ;
        RECT 106.100 194.800 108.200 195.100 ;
        RECT 106.100 194.400 106.500 194.800 ;
        RECT 105.300 193.400 106.600 193.700 ;
        RECT 104.500 192.800 105.000 193.100 ;
        RECT 104.600 191.100 105.000 192.800 ;
        RECT 106.200 191.100 106.600 193.400 ;
        RECT 108.600 193.600 109.000 195.300 ;
        RECT 110.300 195.200 110.700 195.300 ;
        RECT 109.500 194.900 109.900 195.000 ;
        RECT 109.500 194.600 111.400 194.900 ;
        RECT 111.000 194.500 111.400 194.600 ;
        RECT 111.900 194.200 112.200 195.800 ;
        RECT 112.900 195.900 113.200 196.500 ;
        RECT 113.500 196.500 113.900 196.600 ;
        RECT 115.800 196.500 116.200 196.600 ;
        RECT 113.500 196.200 116.200 196.500 ;
        RECT 112.900 195.700 115.300 195.900 ;
        RECT 117.400 195.700 117.800 199.900 ;
        RECT 112.900 195.600 117.800 195.700 ;
        RECT 114.900 195.500 117.800 195.600 ;
        RECT 115.000 195.400 117.800 195.500 ;
        RECT 114.200 195.100 114.600 195.200 ;
        RECT 119.000 195.100 119.400 199.900 ;
        RECT 121.000 196.800 121.400 197.200 ;
        RECT 119.800 195.800 120.200 196.600 ;
        RECT 121.000 196.200 121.300 196.800 ;
        RECT 121.700 196.200 122.100 199.900 ;
        RECT 124.600 196.400 125.000 199.900 ;
        RECT 120.600 195.900 121.300 196.200 ;
        RECT 121.600 195.900 122.100 196.200 ;
        RECT 124.500 195.900 125.000 196.400 ;
        RECT 126.200 196.200 126.600 199.900 ;
        RECT 125.300 195.900 126.600 196.200 ;
        RECT 120.600 195.800 121.000 195.900 ;
        RECT 120.600 195.100 120.900 195.800 ;
        RECT 121.600 195.200 121.900 195.900 ;
        RECT 114.200 194.800 116.700 195.100 ;
        RECT 115.000 194.700 115.400 194.800 ;
        RECT 116.300 194.700 116.700 194.800 ;
        RECT 119.000 194.800 120.900 195.100 ;
        RECT 121.400 194.800 121.900 195.200 ;
        RECT 115.500 194.200 115.900 194.300 ;
        RECT 111.900 193.900 117.400 194.200 ;
        RECT 112.100 193.800 112.500 193.900 ;
        RECT 114.200 193.800 114.600 193.900 ;
        RECT 108.600 193.300 110.500 193.600 ;
        RECT 108.600 191.100 109.000 193.300 ;
        RECT 110.100 193.200 110.500 193.300 ;
        RECT 115.000 192.800 115.300 193.900 ;
        RECT 116.600 193.800 117.400 193.900 ;
        RECT 114.100 192.700 114.500 192.800 ;
        RECT 111.000 192.100 111.400 192.500 ;
        RECT 113.100 192.400 114.500 192.700 ;
        RECT 115.000 192.400 115.400 192.800 ;
        RECT 113.100 192.100 113.400 192.400 ;
        RECT 115.800 192.100 116.200 192.500 ;
        RECT 110.700 191.800 111.400 192.100 ;
        RECT 110.700 191.100 111.300 191.800 ;
        RECT 113.000 191.100 113.400 192.100 ;
        RECT 115.200 191.800 116.200 192.100 ;
        RECT 115.200 191.100 115.600 191.800 ;
        RECT 117.400 191.100 117.800 193.500 ;
        RECT 118.200 193.400 118.600 194.200 ;
        RECT 119.000 193.100 119.400 194.800 ;
        RECT 121.600 194.200 121.900 194.800 ;
        RECT 122.200 194.400 122.600 195.200 ;
        RECT 124.500 194.200 124.800 195.900 ;
        RECT 125.300 194.900 125.600 195.900 ;
        RECT 127.000 195.800 127.400 196.600 ;
        RECT 127.800 196.100 128.200 199.900 ;
        RECT 129.800 196.800 130.200 197.200 ;
        RECT 129.800 196.200 130.100 196.800 ;
        RECT 130.500 196.200 130.900 199.900 ;
        RECT 129.400 196.100 130.100 196.200 ;
        RECT 127.800 195.900 130.100 196.100 ;
        RECT 127.800 195.800 129.800 195.900 ;
        RECT 130.400 195.800 131.400 196.200 ;
        RECT 125.100 194.500 125.600 194.900 ;
        RECT 120.600 193.800 121.900 194.200 ;
        RECT 123.000 194.100 123.400 194.200 ;
        RECT 124.500 194.100 125.000 194.200 ;
        RECT 122.600 193.800 125.000 194.100 ;
        RECT 120.700 193.100 121.000 193.800 ;
        RECT 122.600 193.600 123.000 193.800 ;
        RECT 121.500 193.100 123.300 193.300 ;
        RECT 124.500 193.100 124.800 193.800 ;
        RECT 125.300 193.700 125.600 194.500 ;
        RECT 126.100 194.800 126.600 195.200 ;
        RECT 126.100 194.400 126.500 194.800 ;
        RECT 125.300 193.400 126.600 193.700 ;
        RECT 119.000 192.800 119.900 193.100 ;
        RECT 119.500 191.100 119.900 192.800 ;
        RECT 120.600 191.100 121.000 193.100 ;
        RECT 121.400 193.000 123.400 193.100 ;
        RECT 121.400 191.100 121.800 193.000 ;
        RECT 123.000 191.100 123.400 193.000 ;
        RECT 124.500 192.800 125.000 193.100 ;
        RECT 124.600 191.100 125.000 192.800 ;
        RECT 126.200 191.100 126.600 193.400 ;
        RECT 127.800 193.100 128.200 195.800 ;
        RECT 130.400 194.200 130.700 195.800 ;
        RECT 132.600 195.700 133.000 199.900 ;
        RECT 134.800 198.200 135.200 199.900 ;
        RECT 134.200 197.900 135.200 198.200 ;
        RECT 137.000 197.900 137.400 199.900 ;
        RECT 139.100 197.900 139.700 199.900 ;
        RECT 134.200 197.500 134.600 197.900 ;
        RECT 137.000 197.600 137.300 197.900 ;
        RECT 135.900 197.300 137.700 197.600 ;
        RECT 139.000 197.500 139.400 197.900 ;
        RECT 135.900 197.200 136.300 197.300 ;
        RECT 137.300 197.200 137.700 197.300 ;
        RECT 134.200 196.500 134.600 196.600 ;
        RECT 136.500 196.500 136.900 196.600 ;
        RECT 134.200 196.200 136.900 196.500 ;
        RECT 137.200 196.500 138.300 196.800 ;
        RECT 137.200 195.900 137.500 196.500 ;
        RECT 137.900 196.400 138.300 196.500 ;
        RECT 139.100 196.600 139.800 197.000 ;
        RECT 139.100 196.100 139.400 196.600 ;
        RECT 135.100 195.700 137.500 195.900 ;
        RECT 132.600 195.600 137.500 195.700 ;
        RECT 138.200 195.800 139.400 196.100 ;
        RECT 132.600 195.500 135.500 195.600 ;
        RECT 132.600 195.400 135.400 195.500 ;
        RECT 131.000 194.400 131.400 195.200 ;
        RECT 135.800 195.100 136.200 195.200 ;
        RECT 133.700 194.800 136.200 195.100 ;
        RECT 133.700 194.700 134.100 194.800 ;
        RECT 135.000 194.700 135.400 194.800 ;
        RECT 134.500 194.200 134.900 194.300 ;
        RECT 138.200 194.200 138.500 195.800 ;
        RECT 141.400 195.600 141.800 199.900 ;
        RECT 139.700 195.300 141.800 195.600 ;
        RECT 142.200 197.500 142.600 199.500 ;
        RECT 142.200 195.800 142.500 197.500 ;
        RECT 144.300 196.400 144.700 199.900 ;
        RECT 148.900 196.400 149.300 199.900 ;
        RECT 151.000 197.500 151.400 199.500 ;
        RECT 144.300 196.100 145.100 196.400 ;
        RECT 142.200 195.500 144.100 195.800 ;
        RECT 139.700 195.200 140.100 195.300 ;
        RECT 140.500 194.900 140.900 195.000 ;
        RECT 139.000 194.600 140.900 194.900 ;
        RECT 139.000 194.500 139.400 194.600 ;
        RECT 128.600 193.400 129.000 194.200 ;
        RECT 129.400 193.800 130.700 194.200 ;
        RECT 131.800 194.100 132.200 194.200 ;
        RECT 131.400 193.800 132.200 194.100 ;
        RECT 133.000 193.900 138.500 194.200 ;
        RECT 133.000 193.800 133.800 193.900 ;
        RECT 129.500 193.100 129.800 193.800 ;
        RECT 131.400 193.600 131.800 193.800 ;
        RECT 130.300 193.100 132.100 193.300 ;
        RECT 127.300 192.800 128.200 193.100 ;
        RECT 127.300 191.100 127.700 192.800 ;
        RECT 129.400 191.100 129.800 193.100 ;
        RECT 130.200 193.000 132.200 193.100 ;
        RECT 130.200 191.100 130.600 193.000 ;
        RECT 131.800 191.100 132.200 193.000 ;
        RECT 132.600 191.100 133.000 193.500 ;
        RECT 135.100 192.800 135.400 193.900 ;
        RECT 135.800 193.800 136.200 193.900 ;
        RECT 137.900 193.800 138.300 193.900 ;
        RECT 141.400 193.600 141.800 195.300 ;
        RECT 142.200 194.400 142.600 195.200 ;
        RECT 143.000 194.400 143.400 195.200 ;
        RECT 143.800 194.500 144.100 195.500 ;
        RECT 143.800 194.100 144.500 194.500 ;
        RECT 144.800 194.200 145.100 196.100 ;
        RECT 148.500 196.100 149.300 196.400 ;
        RECT 145.400 194.800 145.800 195.600 ;
        RECT 147.800 195.100 148.200 195.600 ;
        RECT 147.000 194.800 148.200 195.100 ;
        RECT 144.800 194.100 145.800 194.200 ;
        RECT 147.000 194.100 147.300 194.800 ;
        RECT 148.500 194.200 148.800 196.100 ;
        RECT 151.100 195.800 151.400 197.500 ;
        RECT 151.800 196.200 152.200 199.900 ;
        RECT 155.500 196.200 155.900 199.900 ;
        RECT 156.200 196.800 156.600 197.200 ;
        RECT 156.300 196.200 156.600 196.800 ;
        RECT 151.800 195.900 152.900 196.200 ;
        RECT 155.500 195.900 156.000 196.200 ;
        RECT 156.300 196.100 157.000 196.200 ;
        RECT 157.400 196.100 157.800 196.200 ;
        RECT 156.300 195.900 157.800 196.100 ;
        RECT 149.500 195.500 151.400 195.800 ;
        RECT 152.600 195.600 152.900 195.900 ;
        RECT 149.500 194.500 149.800 195.500 ;
        RECT 152.600 195.200 153.200 195.600 ;
        RECT 143.800 193.900 144.300 194.100 ;
        RECT 139.900 193.300 141.800 193.600 ;
        RECT 139.900 193.200 140.300 193.300 ;
        RECT 134.200 192.100 134.600 192.500 ;
        RECT 135.000 192.400 135.400 192.800 ;
        RECT 135.900 192.700 136.300 192.800 ;
        RECT 135.900 192.400 137.300 192.700 ;
        RECT 137.000 192.100 137.300 192.400 ;
        RECT 139.000 192.100 139.400 192.500 ;
        RECT 134.200 191.800 135.200 192.100 ;
        RECT 134.800 191.100 135.200 191.800 ;
        RECT 137.000 191.100 137.400 192.100 ;
        RECT 139.000 191.800 139.700 192.100 ;
        RECT 139.100 191.100 139.700 191.800 ;
        RECT 141.400 191.100 141.800 193.300 ;
        RECT 142.200 193.600 144.300 193.900 ;
        RECT 144.800 193.800 147.300 194.100 ;
        RECT 147.800 193.800 148.800 194.200 ;
        RECT 149.100 194.100 149.800 194.500 ;
        RECT 150.200 194.400 150.600 195.200 ;
        RECT 151.000 194.400 151.400 195.200 ;
        RECT 151.800 194.400 152.200 195.200 ;
        RECT 142.200 192.500 142.500 193.600 ;
        RECT 144.800 193.500 145.100 193.800 ;
        RECT 144.700 193.300 145.100 193.500 ;
        RECT 144.300 193.000 145.100 193.300 ;
        RECT 148.500 193.500 148.800 193.800 ;
        RECT 149.300 193.900 149.800 194.100 ;
        RECT 149.300 193.600 151.400 193.900 ;
        RECT 152.600 193.700 152.900 195.200 ;
        RECT 155.000 194.400 155.400 195.200 ;
        RECT 155.700 195.100 156.000 195.900 ;
        RECT 156.600 195.800 157.800 195.900 ;
        RECT 159.000 195.800 159.400 196.600 ;
        RECT 158.200 195.100 158.600 195.200 ;
        RECT 155.700 194.800 158.600 195.100 ;
        RECT 155.700 194.200 156.000 194.800 ;
        RECT 154.200 194.100 154.600 194.200 ;
        RECT 154.200 193.800 155.000 194.100 ;
        RECT 155.700 193.800 157.000 194.200 ;
        RECT 157.400 194.100 157.800 194.200 ;
        RECT 159.800 194.100 160.200 199.900 ;
        RECT 160.600 197.100 161.000 197.200 ;
        RECT 161.400 197.100 161.800 199.900 ;
        RECT 163.500 197.900 164.100 199.900 ;
        RECT 165.800 197.900 166.200 199.900 ;
        RECT 168.000 198.200 168.400 199.900 ;
        RECT 168.000 197.900 169.000 198.200 ;
        RECT 163.800 197.500 164.200 197.900 ;
        RECT 165.900 197.600 166.200 197.900 ;
        RECT 165.500 197.300 167.300 197.600 ;
        RECT 168.600 197.500 169.000 197.900 ;
        RECT 165.500 197.200 165.900 197.300 ;
        RECT 166.900 197.200 167.300 197.300 ;
        RECT 160.600 196.800 161.800 197.100 ;
        RECT 161.400 195.600 161.800 196.800 ;
        RECT 163.400 196.600 164.100 197.000 ;
        RECT 163.800 196.100 164.100 196.600 ;
        RECT 164.900 196.500 166.000 196.800 ;
        RECT 164.900 196.400 165.300 196.500 ;
        RECT 163.800 195.800 165.000 196.100 ;
        RECT 161.400 195.300 163.500 195.600 ;
        RECT 157.400 193.800 160.200 194.100 ;
        RECT 148.500 193.300 148.900 193.500 ;
        RECT 148.500 193.000 149.300 193.300 ;
        RECT 142.200 191.500 142.600 192.500 ;
        RECT 144.300 191.500 144.700 193.000 ;
        RECT 148.900 192.200 149.300 193.000 ;
        RECT 151.100 192.500 151.400 193.600 ;
        RECT 148.600 191.800 149.300 192.200 ;
        RECT 148.900 191.500 149.300 191.800 ;
        RECT 151.000 191.500 151.400 192.500 ;
        RECT 151.800 193.400 152.900 193.700 ;
        RECT 154.600 193.600 155.000 193.800 ;
        RECT 151.800 191.100 152.200 193.400 ;
        RECT 154.300 193.100 156.100 193.300 ;
        RECT 156.600 193.100 156.900 193.800 ;
        RECT 159.800 193.100 160.200 193.800 ;
        RECT 160.600 193.400 161.000 194.200 ;
        RECT 161.400 193.600 161.800 195.300 ;
        RECT 163.100 195.200 163.500 195.300 ;
        RECT 162.300 194.900 162.700 195.000 ;
        RECT 162.300 194.600 164.200 194.900 ;
        RECT 163.800 194.500 164.200 194.600 ;
        RECT 164.700 194.200 165.000 195.800 ;
        RECT 165.700 195.900 166.000 196.500 ;
        RECT 166.300 196.500 166.700 196.600 ;
        RECT 168.600 196.500 169.000 196.600 ;
        RECT 166.300 196.200 169.000 196.500 ;
        RECT 165.700 195.700 168.100 195.900 ;
        RECT 170.200 195.700 170.600 199.900 ;
        RECT 171.800 196.400 172.200 199.900 ;
        RECT 165.700 195.600 170.600 195.700 ;
        RECT 167.700 195.500 170.600 195.600 ;
        RECT 167.800 195.400 170.600 195.500 ;
        RECT 171.700 195.900 172.200 196.400 ;
        RECT 173.400 196.200 173.800 199.900 ;
        RECT 172.500 195.900 173.800 196.200 ;
        RECT 167.000 195.100 167.400 195.200 ;
        RECT 167.000 194.800 169.500 195.100 ;
        RECT 169.100 194.700 169.500 194.800 ;
        RECT 168.300 194.200 168.700 194.300 ;
        RECT 171.700 194.200 172.000 195.900 ;
        RECT 172.500 194.900 172.800 195.900 ;
        RECT 172.300 194.500 172.800 194.900 ;
        RECT 164.700 193.900 170.200 194.200 ;
        RECT 164.900 193.800 165.300 193.900 ;
        RECT 154.200 193.000 156.200 193.100 ;
        RECT 154.200 191.100 154.600 193.000 ;
        RECT 155.800 191.100 156.200 193.000 ;
        RECT 156.600 191.100 157.000 193.100 ;
        RECT 159.300 192.800 160.200 193.100 ;
        RECT 161.400 193.300 163.300 193.600 ;
        RECT 159.300 191.100 159.700 192.800 ;
        RECT 161.400 191.100 161.800 193.300 ;
        RECT 162.900 193.200 163.300 193.300 ;
        RECT 167.800 192.800 168.100 193.900 ;
        RECT 169.400 193.800 170.200 193.900 ;
        RECT 171.700 193.800 172.200 194.200 ;
        RECT 166.900 192.700 167.300 192.800 ;
        RECT 163.800 192.100 164.200 192.500 ;
        RECT 165.900 192.400 167.300 192.700 ;
        RECT 167.800 192.400 168.200 192.800 ;
        RECT 165.900 192.100 166.200 192.400 ;
        RECT 168.600 192.100 169.000 192.500 ;
        RECT 163.500 191.800 164.200 192.100 ;
        RECT 163.500 191.100 164.100 191.800 ;
        RECT 165.800 191.100 166.200 192.100 ;
        RECT 168.000 191.800 169.000 192.100 ;
        RECT 168.000 191.100 168.400 191.800 ;
        RECT 170.200 191.100 170.600 193.500 ;
        RECT 171.700 193.100 172.000 193.800 ;
        RECT 172.500 193.700 172.800 194.500 ;
        RECT 173.300 194.800 173.800 195.200 ;
        RECT 175.000 195.100 175.400 199.900 ;
        RECT 177.700 199.200 178.100 199.900 ;
        RECT 177.700 198.800 178.600 199.200 ;
        RECT 177.700 196.400 178.100 198.800 ;
        RECT 179.800 197.500 180.200 199.500 ;
        RECT 177.300 196.100 178.100 196.400 ;
        RECT 176.600 195.100 177.000 195.600 ;
        RECT 175.000 194.800 177.000 195.100 ;
        RECT 173.300 194.400 173.700 194.800 ;
        RECT 172.500 193.400 173.800 193.700 ;
        RECT 171.700 192.800 172.200 193.100 ;
        RECT 171.800 191.100 172.200 192.800 ;
        RECT 173.400 191.100 173.800 193.400 ;
        RECT 174.200 192.400 174.600 193.200 ;
        RECT 175.000 191.100 175.400 194.800 ;
        RECT 177.300 194.200 177.600 196.100 ;
        RECT 179.900 195.800 180.200 197.500 ;
        RECT 178.300 195.500 180.200 195.800 ;
        RECT 178.300 194.500 178.600 195.500 ;
        RECT 176.600 193.800 177.600 194.200 ;
        RECT 177.900 194.100 178.600 194.500 ;
        RECT 179.000 194.400 179.400 195.200 ;
        RECT 179.800 194.400 180.200 195.200 ;
        RECT 181.400 195.100 181.800 199.900 ;
        RECT 184.100 199.200 184.500 199.900 ;
        RECT 184.100 198.800 185.000 199.200 ;
        RECT 183.400 196.800 183.800 197.200 ;
        RECT 182.200 195.800 182.600 196.600 ;
        RECT 183.400 196.200 183.700 196.800 ;
        RECT 184.100 196.200 184.500 198.800 ;
        RECT 183.000 195.900 183.700 196.200 ;
        RECT 184.000 195.900 184.500 196.200 ;
        RECT 186.200 197.500 186.600 199.500 ;
        RECT 183.000 195.800 183.400 195.900 ;
        RECT 183.000 195.100 183.300 195.800 ;
        RECT 181.400 194.800 183.300 195.100 ;
        RECT 177.300 193.500 177.600 193.800 ;
        RECT 178.100 193.900 178.600 194.100 ;
        RECT 178.100 193.600 180.200 193.900 ;
        RECT 177.300 193.300 177.700 193.500 ;
        RECT 177.300 193.000 178.100 193.300 ;
        RECT 177.700 191.500 178.100 193.000 ;
        RECT 179.900 192.500 180.200 193.600 ;
        RECT 180.600 193.400 181.000 194.200 ;
        RECT 181.400 193.100 181.800 194.800 ;
        RECT 184.000 194.200 184.300 195.900 ;
        RECT 186.200 195.800 186.500 197.500 ;
        RECT 188.300 196.400 188.700 199.900 ;
        RECT 188.300 196.100 189.100 196.400 ;
        RECT 186.200 195.500 188.100 195.800 ;
        RECT 184.600 194.400 185.000 195.200 ;
        RECT 186.200 194.400 186.600 195.200 ;
        RECT 187.000 194.400 187.400 195.200 ;
        RECT 187.800 194.500 188.100 195.500 ;
        RECT 183.000 193.800 184.300 194.200 ;
        RECT 185.400 194.100 185.800 194.200 ;
        RECT 185.000 193.800 185.800 194.100 ;
        RECT 187.800 194.100 188.500 194.500 ;
        RECT 188.800 194.200 189.100 196.100 ;
        RECT 189.400 195.100 189.800 195.600 ;
        RECT 191.000 195.100 191.400 199.900 ;
        RECT 189.400 194.800 191.400 195.100 ;
        RECT 188.800 194.100 189.800 194.200 ;
        RECT 190.200 194.100 190.600 194.200 ;
        RECT 187.800 193.900 188.300 194.100 ;
        RECT 183.100 193.100 183.400 193.800 ;
        RECT 185.000 193.600 185.400 193.800 ;
        RECT 186.200 193.600 188.300 193.900 ;
        RECT 188.800 193.800 190.600 194.100 ;
        RECT 183.900 193.100 185.700 193.300 ;
        RECT 181.400 192.800 182.300 193.100 ;
        RECT 179.800 191.500 180.200 192.500 ;
        RECT 181.900 191.100 182.300 192.800 ;
        RECT 183.000 191.100 183.400 193.100 ;
        RECT 183.800 193.000 185.800 193.100 ;
        RECT 183.800 191.100 184.200 193.000 ;
        RECT 185.400 191.100 185.800 193.000 ;
        RECT 186.200 192.500 186.500 193.600 ;
        RECT 188.800 193.500 189.100 193.800 ;
        RECT 188.700 193.300 189.100 193.500 ;
        RECT 188.300 193.000 189.100 193.300 ;
        RECT 186.200 191.500 186.600 192.500 ;
        RECT 188.300 191.500 188.700 193.000 ;
        RECT 191.000 191.100 191.400 194.800 ;
        RECT 192.600 195.600 193.000 199.900 ;
        RECT 194.700 197.900 195.300 199.900 ;
        RECT 197.000 197.900 197.400 199.900 ;
        RECT 199.200 198.200 199.600 199.900 ;
        RECT 199.200 197.900 200.200 198.200 ;
        RECT 195.000 197.500 195.400 197.900 ;
        RECT 197.100 197.600 197.400 197.900 ;
        RECT 196.700 197.300 198.500 197.600 ;
        RECT 199.800 197.500 200.200 197.900 ;
        RECT 196.700 197.200 197.100 197.300 ;
        RECT 198.100 197.200 198.500 197.300 ;
        RECT 194.600 196.600 195.300 197.000 ;
        RECT 195.000 196.100 195.300 196.600 ;
        RECT 196.100 196.500 197.200 196.800 ;
        RECT 196.100 196.400 196.500 196.500 ;
        RECT 195.000 195.800 196.200 196.100 ;
        RECT 192.600 195.300 194.700 195.600 ;
        RECT 192.600 193.600 193.000 195.300 ;
        RECT 194.300 195.200 194.700 195.300 ;
        RECT 193.500 194.900 193.900 195.000 ;
        RECT 193.500 194.600 195.400 194.900 ;
        RECT 195.000 194.500 195.400 194.600 ;
        RECT 195.900 194.200 196.200 195.800 ;
        RECT 196.900 195.900 197.200 196.500 ;
        RECT 197.500 196.500 197.900 196.600 ;
        RECT 199.800 196.500 200.200 196.600 ;
        RECT 197.500 196.200 200.200 196.500 ;
        RECT 196.900 195.700 199.300 195.900 ;
        RECT 201.400 195.700 201.800 199.900 ;
        RECT 196.900 195.600 201.800 195.700 ;
        RECT 198.900 195.500 201.800 195.600 ;
        RECT 199.000 195.400 201.800 195.500 ;
        RECT 202.200 195.600 202.600 199.900 ;
        RECT 204.300 197.900 204.900 199.900 ;
        RECT 206.600 197.900 207.000 199.900 ;
        RECT 208.800 198.200 209.200 199.900 ;
        RECT 208.800 197.900 209.800 198.200 ;
        RECT 204.600 197.500 205.000 197.900 ;
        RECT 206.700 197.600 207.000 197.900 ;
        RECT 206.300 197.300 208.100 197.600 ;
        RECT 209.400 197.500 209.800 197.900 ;
        RECT 206.300 197.200 206.700 197.300 ;
        RECT 207.700 197.200 208.100 197.300 ;
        RECT 204.200 196.600 204.900 197.000 ;
        RECT 204.600 196.100 204.900 196.600 ;
        RECT 205.700 196.500 206.800 196.800 ;
        RECT 205.700 196.400 206.100 196.500 ;
        RECT 204.600 195.800 205.800 196.100 ;
        RECT 202.200 195.300 204.300 195.600 ;
        RECT 198.200 195.100 198.600 195.200 ;
        RECT 198.200 194.800 200.700 195.100 ;
        RECT 200.300 194.700 200.700 194.800 ;
        RECT 199.500 194.200 199.900 194.300 ;
        RECT 195.900 193.900 201.400 194.200 ;
        RECT 196.100 193.800 196.500 193.900 ;
        RECT 192.600 193.300 194.500 193.600 ;
        RECT 191.800 193.100 192.200 193.200 ;
        RECT 192.600 193.100 193.000 193.300 ;
        RECT 194.100 193.200 194.500 193.300 ;
        RECT 191.800 192.800 193.000 193.100 ;
        RECT 199.000 192.800 199.300 193.900 ;
        RECT 200.600 193.800 201.400 193.900 ;
        RECT 202.200 193.600 202.600 195.300 ;
        RECT 203.900 195.200 204.300 195.300 ;
        RECT 203.100 194.900 203.500 195.000 ;
        RECT 203.100 194.600 205.000 194.900 ;
        RECT 204.600 194.500 205.000 194.600 ;
        RECT 205.500 194.200 205.800 195.800 ;
        RECT 206.500 195.900 206.800 196.500 ;
        RECT 207.100 196.500 207.500 196.600 ;
        RECT 209.400 196.500 209.800 196.600 ;
        RECT 207.100 196.200 209.800 196.500 ;
        RECT 206.500 195.700 208.900 195.900 ;
        RECT 211.000 195.700 211.400 199.900 ;
        RECT 206.500 195.600 211.400 195.700 ;
        RECT 208.500 195.500 211.400 195.600 ;
        RECT 208.600 195.400 211.400 195.500 ;
        RECT 207.800 195.100 208.200 195.200 ;
        RECT 214.200 195.100 214.600 199.900 ;
        RECT 216.200 196.800 216.600 197.200 ;
        RECT 215.000 195.800 215.400 196.600 ;
        RECT 216.200 196.200 216.500 196.800 ;
        RECT 216.900 196.200 217.300 199.900 ;
        RECT 215.800 195.900 216.500 196.200 ;
        RECT 216.800 195.900 217.300 196.200 ;
        RECT 219.000 197.500 219.400 199.500 ;
        RECT 215.800 195.800 216.200 195.900 ;
        RECT 215.800 195.100 216.100 195.800 ;
        RECT 207.800 194.800 210.300 195.100 ;
        RECT 208.600 194.700 209.000 194.800 ;
        RECT 209.900 194.700 210.300 194.800 ;
        RECT 214.200 194.800 216.100 195.100 ;
        RECT 209.100 194.200 209.500 194.300 ;
        RECT 205.500 193.900 211.000 194.200 ;
        RECT 205.700 193.800 206.100 193.900 ;
        RECT 207.000 193.800 207.400 193.900 ;
        RECT 191.800 192.400 192.200 192.800 ;
        RECT 192.600 191.100 193.000 192.800 ;
        RECT 198.100 192.700 198.500 192.800 ;
        RECT 195.000 192.100 195.400 192.500 ;
        RECT 197.100 192.400 198.500 192.700 ;
        RECT 199.000 192.400 199.400 192.800 ;
        RECT 197.100 192.100 197.400 192.400 ;
        RECT 199.800 192.100 200.200 192.500 ;
        RECT 194.700 191.800 195.400 192.100 ;
        RECT 194.700 191.100 195.300 191.800 ;
        RECT 197.000 191.100 197.400 192.100 ;
        RECT 199.200 191.800 200.200 192.100 ;
        RECT 199.200 191.100 199.600 191.800 ;
        RECT 201.400 191.100 201.800 193.500 ;
        RECT 202.200 193.300 204.100 193.600 ;
        RECT 202.200 191.100 202.600 193.300 ;
        RECT 203.700 193.200 204.100 193.300 ;
        RECT 208.600 192.800 208.900 193.900 ;
        RECT 210.200 193.800 211.000 193.900 ;
        RECT 211.800 194.100 212.200 194.200 ;
        RECT 213.400 194.100 213.800 194.200 ;
        RECT 211.800 193.800 213.800 194.100 ;
        RECT 207.700 192.700 208.100 192.800 ;
        RECT 204.600 192.100 205.000 192.500 ;
        RECT 206.700 192.400 208.100 192.700 ;
        RECT 208.600 192.400 209.000 192.800 ;
        RECT 206.700 192.100 207.000 192.400 ;
        RECT 209.400 192.100 209.800 192.500 ;
        RECT 204.300 191.800 205.000 192.100 ;
        RECT 204.300 191.100 204.900 191.800 ;
        RECT 206.600 191.100 207.000 192.100 ;
        RECT 208.800 191.800 209.800 192.100 ;
        RECT 208.800 191.100 209.200 191.800 ;
        RECT 211.000 191.100 211.400 193.500 ;
        RECT 213.400 193.400 213.800 193.800 ;
        RECT 214.200 193.100 214.600 194.800 ;
        RECT 216.800 194.200 217.100 195.900 ;
        RECT 219.000 195.800 219.300 197.500 ;
        RECT 221.100 196.400 221.500 199.900 ;
        RECT 221.100 196.100 221.900 196.400 ;
        RECT 219.000 195.500 220.900 195.800 ;
        RECT 217.400 194.400 217.800 195.200 ;
        RECT 219.000 194.400 219.400 195.200 ;
        RECT 219.800 194.400 220.200 195.200 ;
        RECT 220.600 194.500 220.900 195.500 ;
        RECT 215.000 194.100 215.400 194.200 ;
        RECT 215.800 194.100 217.100 194.200 ;
        RECT 218.200 194.100 218.600 194.200 ;
        RECT 215.000 193.800 217.100 194.100 ;
        RECT 217.800 193.800 218.600 194.100 ;
        RECT 220.600 194.100 221.300 194.500 ;
        RECT 221.600 194.200 221.900 196.100 ;
        RECT 223.800 196.200 224.200 199.900 ;
        RECT 225.400 196.400 225.800 199.900 ;
        RECT 223.800 195.900 225.100 196.200 ;
        RECT 225.400 195.900 225.900 196.400 ;
        RECT 228.300 196.200 228.700 199.900 ;
        RECT 229.000 196.800 229.400 197.200 ;
        RECT 229.100 196.200 229.400 196.800 ;
        RECT 228.300 195.900 228.800 196.200 ;
        RECT 229.100 195.900 229.800 196.200 ;
        RECT 222.200 194.800 222.600 195.600 ;
        RECT 223.800 194.800 224.300 195.200 ;
        RECT 223.900 194.400 224.300 194.800 ;
        RECT 224.800 194.900 225.100 195.900 ;
        RECT 224.800 194.500 225.300 194.900 ;
        RECT 220.600 193.900 221.100 194.100 ;
        RECT 215.900 193.100 216.200 193.800 ;
        RECT 217.800 193.600 218.200 193.800 ;
        RECT 219.000 193.600 221.100 193.900 ;
        RECT 221.600 193.800 222.600 194.200 ;
        RECT 216.700 193.100 218.500 193.300 ;
        RECT 214.200 192.800 215.100 193.100 ;
        RECT 214.700 191.100 215.100 192.800 ;
        RECT 215.800 191.100 216.200 193.100 ;
        RECT 216.600 193.000 218.600 193.100 ;
        RECT 216.600 191.100 217.000 193.000 ;
        RECT 218.200 191.100 218.600 193.000 ;
        RECT 219.000 192.500 219.300 193.600 ;
        RECT 221.600 193.500 221.900 193.800 ;
        RECT 224.800 193.700 225.100 194.500 ;
        RECT 225.600 194.200 225.900 195.900 ;
        RECT 227.000 195.100 227.400 195.200 ;
        RECT 227.800 195.100 228.200 195.200 ;
        RECT 227.000 194.800 228.200 195.100 ;
        RECT 227.800 194.400 228.200 194.800 ;
        RECT 228.500 194.200 228.800 195.900 ;
        RECT 229.400 195.800 229.800 195.900 ;
        RECT 230.200 195.800 230.600 196.600 ;
        RECT 229.400 195.100 229.700 195.800 ;
        RECT 231.000 195.100 231.400 199.900 ;
        RECT 231.800 197.100 232.200 197.200 ;
        RECT 232.600 197.100 233.000 199.900 ;
        RECT 234.700 197.900 235.300 199.900 ;
        RECT 237.000 197.900 237.400 199.900 ;
        RECT 239.200 198.200 239.600 199.900 ;
        RECT 239.200 197.900 240.200 198.200 ;
        RECT 235.000 197.500 235.400 197.900 ;
        RECT 237.100 197.600 237.400 197.900 ;
        RECT 236.700 197.300 238.500 197.600 ;
        RECT 239.800 197.500 240.200 197.900 ;
        RECT 236.700 197.200 237.100 197.300 ;
        RECT 238.100 197.200 238.500 197.300 ;
        RECT 231.800 196.800 233.000 197.100 ;
        RECT 229.400 194.800 231.400 195.100 ;
        RECT 225.400 193.800 225.900 194.200 ;
        RECT 227.000 194.100 227.400 194.200 ;
        RECT 228.500 194.100 229.800 194.200 ;
        RECT 230.200 194.100 230.600 194.200 ;
        RECT 227.000 193.800 227.800 194.100 ;
        RECT 228.500 193.800 230.600 194.100 ;
        RECT 221.500 193.300 221.900 193.500 ;
        RECT 221.100 193.000 221.900 193.300 ;
        RECT 223.800 193.400 225.100 193.700 ;
        RECT 219.000 191.500 219.400 192.500 ;
        RECT 221.100 192.200 221.500 193.000 ;
        RECT 220.600 191.800 221.500 192.200 ;
        RECT 221.100 191.500 221.500 191.800 ;
        RECT 223.800 191.100 224.200 193.400 ;
        RECT 225.600 193.100 225.900 193.800 ;
        RECT 227.400 193.600 227.800 193.800 ;
        RECT 227.100 193.100 228.900 193.300 ;
        RECT 229.400 193.100 229.700 193.800 ;
        RECT 231.000 193.100 231.400 194.800 ;
        RECT 232.600 195.600 233.000 196.800 ;
        RECT 234.600 196.600 235.300 197.000 ;
        RECT 235.000 196.100 235.300 196.600 ;
        RECT 236.100 196.500 237.200 196.800 ;
        RECT 236.100 196.400 236.500 196.500 ;
        RECT 235.000 195.800 236.200 196.100 ;
        RECT 232.600 195.300 234.700 195.600 ;
        RECT 231.800 193.400 232.200 194.200 ;
        RECT 232.600 193.600 233.000 195.300 ;
        RECT 234.300 195.200 234.700 195.300 ;
        RECT 233.500 194.900 233.900 195.000 ;
        RECT 233.500 194.600 235.400 194.900 ;
        RECT 235.000 194.500 235.400 194.600 ;
        RECT 235.900 194.200 236.200 195.800 ;
        RECT 236.900 195.900 237.200 196.500 ;
        RECT 237.500 196.500 237.900 196.600 ;
        RECT 239.800 196.500 240.200 196.600 ;
        RECT 237.500 196.200 240.200 196.500 ;
        RECT 236.900 195.700 239.300 195.900 ;
        RECT 241.400 195.700 241.800 199.900 ;
        RECT 236.900 195.600 241.800 195.700 ;
        RECT 238.900 195.500 241.800 195.600 ;
        RECT 242.200 197.500 242.600 199.500 ;
        RECT 242.200 195.800 242.500 197.500 ;
        RECT 244.300 196.400 244.700 199.900 ;
        RECT 248.300 199.200 248.700 199.900 ;
        RECT 247.800 198.800 248.700 199.200 ;
        RECT 244.300 196.100 245.100 196.400 ;
        RECT 242.200 195.500 244.100 195.800 ;
        RECT 239.000 195.400 241.800 195.500 ;
        RECT 238.200 195.100 238.600 195.200 ;
        RECT 238.200 194.800 240.700 195.100 ;
        RECT 240.300 194.700 240.700 194.800 ;
        RECT 242.200 194.400 242.600 195.200 ;
        RECT 243.000 194.400 243.400 195.200 ;
        RECT 243.800 194.500 244.100 195.500 ;
        RECT 239.500 194.200 239.900 194.300 ;
        RECT 235.900 193.900 241.400 194.200 ;
        RECT 243.800 194.100 244.500 194.500 ;
        RECT 244.800 194.200 245.100 196.100 ;
        RECT 248.300 196.200 248.700 198.800 ;
        RECT 249.000 196.800 249.400 197.200 ;
        RECT 249.100 196.200 249.400 196.800 ;
        RECT 248.300 195.900 248.800 196.200 ;
        RECT 249.100 195.900 249.800 196.200 ;
        RECT 245.400 194.800 245.800 195.600 ;
        RECT 247.800 194.400 248.200 195.200 ;
        RECT 248.500 194.200 248.800 195.900 ;
        RECT 249.400 195.800 249.800 195.900 ;
        RECT 249.400 195.100 249.800 195.200 ;
        RECT 250.200 195.100 250.600 199.900 ;
        RECT 249.400 194.800 250.600 195.100 ;
        RECT 244.800 194.100 245.800 194.200 ;
        RECT 246.200 194.100 246.600 194.200 ;
        RECT 243.800 193.900 244.300 194.100 ;
        RECT 236.100 193.800 236.500 193.900 ;
        RECT 225.400 192.800 225.900 193.100 ;
        RECT 227.000 193.000 229.000 193.100 ;
        RECT 225.400 191.100 225.800 192.800 ;
        RECT 227.000 191.100 227.400 193.000 ;
        RECT 228.600 191.100 229.000 193.000 ;
        RECT 229.400 191.100 229.800 193.100 ;
        RECT 230.500 192.800 231.400 193.100 ;
        RECT 232.600 193.300 234.500 193.600 ;
        RECT 230.500 191.100 230.900 192.800 ;
        RECT 232.600 191.100 233.000 193.300 ;
        RECT 234.100 193.200 234.500 193.300 ;
        RECT 239.000 192.800 239.300 193.900 ;
        RECT 240.600 193.800 241.400 193.900 ;
        RECT 242.200 193.600 244.300 193.900 ;
        RECT 244.800 193.800 246.600 194.100 ;
        RECT 247.000 194.100 247.400 194.200 ;
        RECT 247.000 193.800 247.800 194.100 ;
        RECT 248.500 193.800 249.800 194.200 ;
        RECT 238.100 192.700 238.500 192.800 ;
        RECT 235.000 192.100 235.400 192.500 ;
        RECT 237.100 192.400 238.500 192.700 ;
        RECT 239.000 192.400 239.400 192.800 ;
        RECT 237.100 192.100 237.400 192.400 ;
        RECT 239.800 192.100 240.200 192.500 ;
        RECT 234.700 191.800 235.400 192.100 ;
        RECT 234.700 191.100 235.300 191.800 ;
        RECT 237.000 191.100 237.400 192.100 ;
        RECT 239.200 191.800 240.200 192.100 ;
        RECT 239.200 191.100 239.600 191.800 ;
        RECT 241.400 191.100 241.800 193.500 ;
        RECT 242.200 192.500 242.500 193.600 ;
        RECT 244.800 193.500 245.100 193.800 ;
        RECT 247.400 193.600 247.800 193.800 ;
        RECT 244.700 193.300 245.100 193.500 ;
        RECT 244.300 193.000 245.100 193.300 ;
        RECT 247.100 193.100 248.900 193.300 ;
        RECT 249.400 193.100 249.700 193.800 ;
        RECT 247.000 193.000 249.000 193.100 ;
        RECT 242.200 191.500 242.600 192.500 ;
        RECT 244.300 191.500 244.700 193.000 ;
        RECT 247.000 191.100 247.400 193.000 ;
        RECT 248.600 191.100 249.000 193.000 ;
        RECT 249.400 191.100 249.800 193.100 ;
        RECT 250.200 191.100 250.600 194.800 ;
        RECT 251.800 195.600 252.200 199.900 ;
        RECT 253.900 197.900 254.500 199.900 ;
        RECT 256.200 197.900 256.600 199.900 ;
        RECT 258.400 198.200 258.800 199.900 ;
        RECT 258.400 197.900 259.400 198.200 ;
        RECT 254.200 197.500 254.600 197.900 ;
        RECT 256.300 197.600 256.600 197.900 ;
        RECT 255.900 197.300 257.700 197.600 ;
        RECT 259.000 197.500 259.400 197.900 ;
        RECT 255.900 197.200 256.300 197.300 ;
        RECT 257.300 197.200 257.700 197.300 ;
        RECT 253.400 197.000 254.100 197.200 ;
        RECT 253.400 196.800 254.500 197.000 ;
        RECT 253.800 196.600 254.500 196.800 ;
        RECT 254.200 196.100 254.500 196.600 ;
        RECT 255.300 196.500 256.400 196.800 ;
        RECT 255.300 196.400 255.700 196.500 ;
        RECT 254.200 195.800 255.400 196.100 ;
        RECT 251.800 195.300 253.900 195.600 ;
        RECT 251.800 193.600 252.200 195.300 ;
        RECT 253.500 195.200 253.900 195.300 ;
        RECT 252.700 194.900 253.100 195.000 ;
        RECT 252.700 194.600 254.600 194.900 ;
        RECT 254.200 194.500 254.600 194.600 ;
        RECT 255.100 194.200 255.400 195.800 ;
        RECT 256.100 195.900 256.400 196.500 ;
        RECT 256.700 196.500 257.100 196.600 ;
        RECT 259.000 196.500 259.400 196.600 ;
        RECT 256.700 196.200 259.400 196.500 ;
        RECT 256.100 195.700 258.500 195.900 ;
        RECT 260.600 195.700 261.000 199.900 ;
        RECT 262.700 199.200 263.100 199.900 ;
        RECT 262.200 198.800 263.100 199.200 ;
        RECT 262.700 196.200 263.100 198.800 ;
        RECT 263.400 196.800 263.800 197.200 ;
        RECT 263.500 196.200 263.800 196.800 ;
        RECT 262.700 195.900 263.200 196.200 ;
        RECT 263.500 196.100 264.200 196.200 ;
        RECT 264.600 196.100 265.000 196.200 ;
        RECT 263.500 195.900 265.000 196.100 ;
        RECT 256.100 195.600 261.000 195.700 ;
        RECT 258.100 195.500 261.000 195.600 ;
        RECT 258.200 195.400 261.000 195.500 ;
        RECT 257.400 195.100 257.800 195.200 ;
        RECT 257.400 194.800 259.900 195.100 ;
        RECT 259.500 194.700 259.900 194.800 ;
        RECT 262.200 194.400 262.600 195.200 ;
        RECT 258.700 194.200 259.100 194.300 ;
        RECT 262.900 194.200 263.200 195.900 ;
        RECT 263.800 195.800 265.000 195.900 ;
        RECT 255.100 193.900 260.600 194.200 ;
        RECT 255.300 193.800 255.700 193.900 ;
        RECT 251.800 193.300 253.700 193.600 ;
        RECT 251.000 193.100 251.400 193.200 ;
        RECT 251.800 193.100 252.200 193.300 ;
        RECT 253.300 193.200 253.700 193.300 ;
        RECT 251.000 192.800 252.200 193.100 ;
        RECT 258.200 192.800 258.500 193.900 ;
        RECT 259.800 193.800 260.600 193.900 ;
        RECT 261.400 194.100 261.800 194.200 ;
        RECT 261.400 193.800 262.200 194.100 ;
        RECT 262.900 193.800 264.200 194.200 ;
        RECT 261.800 193.600 262.200 193.800 ;
        RECT 251.000 192.400 251.400 192.800 ;
        RECT 251.800 191.100 252.200 192.800 ;
        RECT 257.300 192.700 257.700 192.800 ;
        RECT 254.200 192.100 254.600 192.500 ;
        RECT 256.300 192.400 257.700 192.700 ;
        RECT 258.200 192.400 258.600 192.800 ;
        RECT 256.300 192.100 256.600 192.400 ;
        RECT 259.000 192.100 259.400 192.500 ;
        RECT 253.900 191.800 254.600 192.100 ;
        RECT 253.900 191.100 254.500 191.800 ;
        RECT 256.200 191.100 256.600 192.100 ;
        RECT 258.400 191.800 259.400 192.100 ;
        RECT 258.400 191.100 258.800 191.800 ;
        RECT 260.600 191.100 261.000 193.500 ;
        RECT 261.500 193.100 263.300 193.300 ;
        RECT 263.800 193.100 264.100 193.800 ;
        RECT 261.400 193.000 263.400 193.100 ;
        RECT 261.400 191.100 261.800 193.000 ;
        RECT 263.000 191.100 263.400 193.000 ;
        RECT 263.800 191.100 264.200 193.100 ;
        RECT 0.600 187.500 1.000 189.900 ;
        RECT 2.800 189.200 3.200 189.900 ;
        RECT 2.200 188.900 3.200 189.200 ;
        RECT 5.000 188.900 5.400 189.900 ;
        RECT 7.100 189.200 7.700 189.900 ;
        RECT 7.000 188.900 7.700 189.200 ;
        RECT 2.200 188.500 2.600 188.900 ;
        RECT 5.000 188.600 5.300 188.900 ;
        RECT 3.000 188.200 3.400 188.600 ;
        RECT 3.900 188.300 5.300 188.600 ;
        RECT 7.000 188.500 7.400 188.900 ;
        RECT 3.900 188.200 4.300 188.300 ;
        RECT 1.000 187.100 1.800 187.200 ;
        RECT 3.100 187.100 3.400 188.200 ;
        RECT 9.400 188.100 9.800 189.900 ;
        RECT 10.200 188.100 10.600 188.600 ;
        RECT 9.400 187.800 10.600 188.100 ;
        RECT 7.900 187.700 8.300 187.800 ;
        RECT 9.400 187.700 9.800 187.800 ;
        RECT 7.900 187.400 9.800 187.700 ;
        RECT 5.900 187.100 6.300 187.200 ;
        RECT 1.000 186.800 6.500 187.100 ;
        RECT 2.500 186.700 2.900 186.800 ;
        RECT 1.700 186.200 2.100 186.300 ;
        RECT 6.200 186.200 6.500 186.800 ;
        RECT 7.000 186.400 7.400 186.500 ;
        RECT 1.700 185.900 4.200 186.200 ;
        RECT 3.800 185.800 4.200 185.900 ;
        RECT 6.200 185.800 6.600 186.200 ;
        RECT 7.000 186.100 8.900 186.400 ;
        RECT 8.500 186.000 8.900 186.100 ;
        RECT 9.400 186.100 9.800 187.400 ;
        RECT 10.200 186.800 10.600 187.200 ;
        RECT 10.200 186.100 10.500 186.800 ;
        RECT 9.400 185.800 10.500 186.100 ;
        RECT 0.600 185.500 3.400 185.600 ;
        RECT 0.600 185.400 3.500 185.500 ;
        RECT 0.600 185.300 5.500 185.400 ;
        RECT 0.600 181.100 1.000 185.300 ;
        RECT 3.100 185.100 5.500 185.300 ;
        RECT 2.200 184.500 4.900 184.800 ;
        RECT 2.200 184.400 2.600 184.500 ;
        RECT 4.500 184.400 4.900 184.500 ;
        RECT 5.200 184.500 5.500 185.100 ;
        RECT 6.200 185.200 6.500 185.800 ;
        RECT 7.700 185.700 8.100 185.800 ;
        RECT 9.400 185.700 9.800 185.800 ;
        RECT 7.700 185.400 9.800 185.700 ;
        RECT 6.200 184.900 7.400 185.200 ;
        RECT 5.900 184.500 6.300 184.600 ;
        RECT 5.200 184.200 6.300 184.500 ;
        RECT 7.100 184.400 7.400 184.900 ;
        RECT 7.100 184.000 7.800 184.400 ;
        RECT 3.900 183.700 4.300 183.800 ;
        RECT 5.300 183.700 5.700 183.800 ;
        RECT 2.200 183.100 2.600 183.500 ;
        RECT 3.900 183.400 5.700 183.700 ;
        RECT 5.000 183.100 5.300 183.400 ;
        RECT 7.000 183.100 7.400 183.500 ;
        RECT 2.200 182.800 3.200 183.100 ;
        RECT 2.800 181.100 3.200 182.800 ;
        RECT 5.000 181.100 5.400 183.100 ;
        RECT 7.100 181.100 7.700 183.100 ;
        RECT 9.400 181.100 9.800 185.400 ;
        RECT 11.000 181.100 11.400 189.900 ;
        RECT 13.700 188.200 14.100 189.500 ;
        RECT 15.800 188.500 16.200 189.500 ;
        RECT 13.700 188.000 14.600 188.200 ;
        RECT 13.300 187.800 14.600 188.000 ;
        RECT 13.300 187.700 14.100 187.800 ;
        RECT 13.300 187.500 13.700 187.700 ;
        RECT 13.300 187.200 13.600 187.500 ;
        RECT 15.900 187.400 16.200 188.500 ;
        RECT 16.600 187.500 17.000 189.900 ;
        RECT 18.800 189.200 19.200 189.900 ;
        RECT 18.200 188.900 19.200 189.200 ;
        RECT 21.000 188.900 21.400 189.900 ;
        RECT 23.100 189.200 23.700 189.900 ;
        RECT 23.000 188.900 23.700 189.200 ;
        RECT 18.200 188.500 18.600 188.900 ;
        RECT 21.000 188.600 21.300 188.900 ;
        RECT 19.000 188.200 19.400 188.600 ;
        RECT 19.900 188.300 21.300 188.600 ;
        RECT 23.000 188.500 23.400 188.900 ;
        RECT 19.900 188.200 20.300 188.300 ;
        RECT 12.600 186.800 13.600 187.200 ;
        RECT 14.100 187.100 16.200 187.400 ;
        RECT 17.000 187.100 17.800 187.200 ;
        RECT 19.100 187.100 19.400 188.200 ;
        RECT 23.900 187.700 24.300 187.800 ;
        RECT 25.400 187.700 25.800 189.900 ;
        RECT 23.900 187.400 25.800 187.700 ;
        RECT 21.900 187.100 22.300 187.200 ;
        RECT 14.100 186.900 14.600 187.100 ;
        RECT 12.600 185.400 13.000 186.200 ;
        RECT 13.300 184.900 13.600 186.800 ;
        RECT 13.900 186.500 14.600 186.900 ;
        RECT 17.000 186.800 22.500 187.100 ;
        RECT 18.500 186.700 18.900 186.800 ;
        RECT 14.300 185.500 14.600 186.500 ;
        RECT 15.000 185.800 15.400 186.600 ;
        RECT 15.800 185.800 16.200 186.600 ;
        RECT 17.700 186.200 18.100 186.300 ;
        RECT 17.700 185.900 20.200 186.200 ;
        RECT 19.800 185.800 20.200 185.900 ;
        RECT 16.600 185.500 19.400 185.600 ;
        RECT 14.300 185.200 16.200 185.500 ;
        RECT 13.300 184.600 14.100 184.900 ;
        RECT 13.700 181.100 14.100 184.600 ;
        RECT 15.900 183.500 16.200 185.200 ;
        RECT 15.800 181.500 16.200 183.500 ;
        RECT 16.600 185.400 19.500 185.500 ;
        RECT 16.600 185.300 21.500 185.400 ;
        RECT 16.600 181.100 17.000 185.300 ;
        RECT 19.100 185.100 21.500 185.300 ;
        RECT 18.200 184.500 20.900 184.800 ;
        RECT 18.200 184.400 18.600 184.500 ;
        RECT 20.500 184.400 20.900 184.500 ;
        RECT 21.200 184.500 21.500 185.100 ;
        RECT 22.200 185.200 22.500 186.800 ;
        RECT 23.000 186.400 23.400 186.500 ;
        RECT 23.000 186.100 24.900 186.400 ;
        RECT 24.500 186.000 24.900 186.100 ;
        RECT 23.700 185.700 24.100 185.800 ;
        RECT 25.400 185.700 25.800 187.400 ;
        RECT 26.200 188.500 26.600 189.500 ;
        RECT 26.200 187.400 26.500 188.500 ;
        RECT 28.300 188.200 28.700 189.500 ;
        RECT 27.800 188.000 28.700 188.200 ;
        RECT 27.800 187.800 29.100 188.000 ;
        RECT 28.300 187.700 29.100 187.800 ;
        RECT 28.700 187.500 29.100 187.700 ;
        RECT 26.200 187.100 28.300 187.400 ;
        RECT 27.800 186.900 28.300 187.100 ;
        RECT 28.800 187.200 29.100 187.500 ;
        RECT 26.200 185.800 26.600 186.600 ;
        RECT 27.000 185.800 27.400 186.600 ;
        RECT 27.800 186.500 28.500 186.900 ;
        RECT 28.800 186.800 29.800 187.200 ;
        RECT 23.700 185.400 25.800 185.700 ;
        RECT 27.800 185.500 28.100 186.500 ;
        RECT 22.200 184.900 23.400 185.200 ;
        RECT 21.900 184.500 22.300 184.600 ;
        RECT 21.200 184.200 22.300 184.500 ;
        RECT 23.100 184.400 23.400 184.900 ;
        RECT 23.100 184.000 23.800 184.400 ;
        RECT 19.900 183.700 20.300 183.800 ;
        RECT 21.300 183.700 21.700 183.800 ;
        RECT 18.200 183.100 18.600 183.500 ;
        RECT 19.900 183.400 21.700 183.700 ;
        RECT 21.000 183.100 21.300 183.400 ;
        RECT 23.000 183.100 23.400 183.500 ;
        RECT 18.200 182.800 19.200 183.100 ;
        RECT 18.800 181.100 19.200 182.800 ;
        RECT 21.000 181.100 21.400 183.100 ;
        RECT 23.100 181.100 23.700 183.100 ;
        RECT 25.400 181.100 25.800 185.400 ;
        RECT 26.200 185.200 28.100 185.500 ;
        RECT 26.200 183.500 26.500 185.200 ;
        RECT 28.800 184.900 29.100 186.800 ;
        RECT 29.400 186.100 29.800 186.200 ;
        RECT 31.000 186.100 31.400 189.900 ;
        RECT 31.800 187.800 32.200 188.600 ;
        RECT 34.500 188.000 34.900 189.500 ;
        RECT 36.600 188.500 37.000 189.500 ;
        RECT 34.100 187.700 34.900 188.000 ;
        RECT 34.100 187.500 34.500 187.700 ;
        RECT 34.100 187.200 34.400 187.500 ;
        RECT 36.700 187.400 37.000 188.500 ;
        RECT 39.300 188.000 39.700 189.500 ;
        RECT 41.400 188.500 41.800 189.500 ;
        RECT 33.400 186.800 34.400 187.200 ;
        RECT 34.900 187.100 37.000 187.400 ;
        RECT 38.900 187.700 39.700 188.000 ;
        RECT 38.900 187.500 39.300 187.700 ;
        RECT 38.900 187.200 39.200 187.500 ;
        RECT 41.500 187.400 41.800 188.500 ;
        RECT 34.900 186.900 35.400 187.100 ;
        RECT 29.400 185.800 31.400 186.100 ;
        RECT 29.400 185.400 29.800 185.800 ;
        RECT 28.300 184.600 29.100 184.900 ;
        RECT 26.200 181.500 26.600 183.500 ;
        RECT 28.300 181.100 28.700 184.600 ;
        RECT 31.000 181.100 31.400 185.800 ;
        RECT 33.400 185.400 33.800 186.200 ;
        RECT 34.100 184.900 34.400 186.800 ;
        RECT 34.700 186.500 35.400 186.900 ;
        RECT 38.200 186.800 39.200 187.200 ;
        RECT 39.700 187.100 41.800 187.400 ;
        RECT 42.200 188.500 42.600 189.500 ;
        RECT 42.200 187.400 42.500 188.500 ;
        RECT 44.300 188.200 44.700 189.500 ;
        RECT 48.300 189.200 48.700 189.900 ;
        RECT 47.800 188.800 48.700 189.200 ;
        RECT 48.300 188.200 48.700 188.800 ;
        RECT 43.800 188.000 44.700 188.200 ;
        RECT 43.800 187.800 45.100 188.000 ;
        RECT 44.300 187.700 45.100 187.800 ;
        RECT 44.700 187.500 45.100 187.700 ;
        RECT 47.800 187.900 48.700 188.200 ;
        RECT 49.400 188.500 49.800 189.500 ;
        RECT 42.200 187.100 44.300 187.400 ;
        RECT 39.700 186.900 40.200 187.100 ;
        RECT 35.100 185.500 35.400 186.500 ;
        RECT 35.800 185.800 36.200 186.600 ;
        RECT 36.600 185.800 37.000 186.600 ;
        RECT 35.100 185.200 37.000 185.500 ;
        RECT 38.200 185.400 38.600 186.200 ;
        RECT 34.100 184.600 34.900 184.900 ;
        RECT 34.500 182.200 34.900 184.600 ;
        RECT 36.700 183.500 37.000 185.200 ;
        RECT 38.900 184.900 39.200 186.800 ;
        RECT 39.500 186.500 40.200 186.900 ;
        RECT 43.800 186.900 44.300 187.100 ;
        RECT 44.800 187.200 45.100 187.500 ;
        RECT 39.900 185.500 40.200 186.500 ;
        RECT 40.600 185.800 41.000 186.600 ;
        RECT 41.400 185.800 41.800 186.600 ;
        RECT 42.200 185.800 42.600 186.600 ;
        RECT 43.000 185.800 43.400 186.600 ;
        RECT 43.800 186.500 44.500 186.900 ;
        RECT 44.800 186.800 45.800 187.200 ;
        RECT 47.000 186.800 47.400 187.600 ;
        RECT 43.800 185.500 44.100 186.500 ;
        RECT 39.900 185.200 41.800 185.500 ;
        RECT 38.900 184.600 39.700 184.900 ;
        RECT 34.500 181.800 35.400 182.200 ;
        RECT 34.500 181.100 34.900 181.800 ;
        RECT 36.600 181.500 37.000 183.500 ;
        RECT 39.300 182.200 39.700 184.600 ;
        RECT 41.500 183.500 41.800 185.200 ;
        RECT 39.300 181.800 40.200 182.200 ;
        RECT 39.300 181.100 39.700 181.800 ;
        RECT 41.400 181.500 41.800 183.500 ;
        RECT 42.200 185.200 44.100 185.500 ;
        RECT 42.200 183.500 42.500 185.200 ;
        RECT 44.800 184.900 45.100 186.800 ;
        RECT 45.400 185.400 45.800 186.200 ;
        RECT 44.300 184.600 45.100 184.900 ;
        RECT 42.200 181.500 42.600 183.500 ;
        RECT 44.300 181.100 44.700 184.600 ;
        RECT 47.800 181.100 48.200 187.900 ;
        RECT 49.400 187.400 49.700 188.500 ;
        RECT 51.500 188.000 51.900 189.500 ;
        RECT 55.800 188.500 56.200 189.500 ;
        RECT 51.500 187.700 52.300 188.000 ;
        RECT 51.900 187.500 52.300 187.700 ;
        RECT 49.400 187.100 51.500 187.400 ;
        RECT 51.000 186.900 51.500 187.100 ;
        RECT 52.000 187.200 52.300 187.500 ;
        RECT 55.800 187.400 56.100 188.500 ;
        RECT 57.900 188.000 58.300 189.500 ;
        RECT 60.600 188.500 61.000 189.500 ;
        RECT 57.900 187.700 58.700 188.000 ;
        RECT 58.300 187.500 58.700 187.700 ;
        RECT 52.000 187.100 53.000 187.200 ;
        RECT 55.000 187.100 55.400 187.200 ;
        RECT 55.800 187.100 57.900 187.400 ;
        RECT 49.400 185.800 49.800 186.600 ;
        RECT 50.200 185.800 50.600 186.600 ;
        RECT 51.000 186.500 51.700 186.900 ;
        RECT 52.000 186.800 55.400 187.100 ;
        RECT 57.400 186.900 57.900 187.100 ;
        RECT 58.400 187.200 58.700 187.500 ;
        RECT 60.600 187.400 60.900 188.500 ;
        RECT 62.700 188.000 63.100 189.500 ;
        RECT 66.700 189.200 67.100 189.900 ;
        RECT 66.700 188.800 67.400 189.200 ;
        RECT 66.700 188.200 67.100 188.800 ;
        RECT 62.700 187.700 63.500 188.000 ;
        RECT 63.100 187.500 63.500 187.700 ;
        RECT 66.200 187.900 67.100 188.200 ;
        RECT 67.800 188.500 68.200 189.500 ;
        RECT 51.000 185.500 51.300 186.500 ;
        RECT 49.400 185.200 51.300 185.500 ;
        RECT 48.600 184.400 49.000 185.200 ;
        RECT 49.400 183.500 49.700 185.200 ;
        RECT 52.000 184.900 52.300 186.800 ;
        RECT 52.600 185.400 53.000 186.200 ;
        RECT 55.800 185.800 56.200 186.600 ;
        RECT 56.600 185.800 57.000 186.600 ;
        RECT 57.400 186.500 58.100 186.900 ;
        RECT 58.400 186.800 59.400 187.200 ;
        RECT 60.600 187.100 62.700 187.400 ;
        RECT 62.200 186.900 62.700 187.100 ;
        RECT 63.200 187.200 63.500 187.500 ;
        RECT 57.400 185.500 57.700 186.500 ;
        RECT 51.500 184.600 52.300 184.900 ;
        RECT 55.800 185.200 57.700 185.500 ;
        RECT 49.400 181.500 49.800 183.500 ;
        RECT 51.500 181.100 51.900 184.600 ;
        RECT 55.800 183.500 56.100 185.200 ;
        RECT 58.400 184.900 58.700 186.800 ;
        RECT 59.000 185.400 59.400 186.200 ;
        RECT 60.600 185.800 61.000 186.600 ;
        RECT 61.400 185.800 61.800 186.600 ;
        RECT 62.200 186.500 62.900 186.900 ;
        RECT 63.200 186.800 64.200 187.200 ;
        RECT 65.400 186.800 65.800 187.600 ;
        RECT 62.200 185.500 62.500 186.500 ;
        RECT 63.200 186.200 63.500 186.800 ;
        RECT 63.000 185.800 63.500 186.200 ;
        RECT 57.900 184.600 58.700 184.900 ;
        RECT 60.600 185.200 62.500 185.500 ;
        RECT 55.800 181.500 56.200 183.500 ;
        RECT 57.900 182.200 58.300 184.600 ;
        RECT 60.600 183.500 60.900 185.200 ;
        RECT 63.200 184.900 63.500 185.800 ;
        RECT 63.800 186.100 64.200 186.200 ;
        RECT 64.600 186.100 65.000 186.200 ;
        RECT 63.800 185.800 65.000 186.100 ;
        RECT 63.800 185.400 64.200 185.800 ;
        RECT 62.700 184.600 63.500 184.900 ;
        RECT 57.900 181.800 58.600 182.200 ;
        RECT 57.900 181.100 58.300 181.800 ;
        RECT 60.600 181.500 61.000 183.500 ;
        RECT 62.700 181.100 63.100 184.600 ;
        RECT 66.200 181.100 66.600 187.900 ;
        RECT 67.800 187.400 68.100 188.500 ;
        RECT 69.900 188.000 70.300 189.500 ;
        RECT 69.900 187.700 70.700 188.000 ;
        RECT 70.300 187.500 70.700 187.700 ;
        RECT 67.800 187.100 69.900 187.400 ;
        RECT 69.400 186.900 69.900 187.100 ;
        RECT 70.400 187.200 70.700 187.500 ;
        RECT 70.400 187.100 71.400 187.200 ;
        RECT 71.800 187.100 72.200 187.200 ;
        RECT 67.800 185.800 68.200 186.600 ;
        RECT 68.600 185.800 69.000 186.600 ;
        RECT 69.400 186.500 70.100 186.900 ;
        RECT 70.400 186.800 72.200 187.100 ;
        RECT 69.400 185.500 69.700 186.500 ;
        RECT 67.800 185.200 69.700 185.500 ;
        RECT 67.000 184.400 67.400 185.200 ;
        RECT 67.800 183.500 68.100 185.200 ;
        RECT 70.400 184.900 70.700 186.800 ;
        RECT 71.000 186.100 71.400 186.200 ;
        RECT 72.600 186.100 73.000 189.900 ;
        RECT 73.400 187.800 73.800 188.600 ;
        RECT 74.200 187.500 74.600 189.900 ;
        RECT 76.400 189.200 76.800 189.900 ;
        RECT 75.800 188.900 76.800 189.200 ;
        RECT 78.600 188.900 79.000 189.900 ;
        RECT 80.700 189.200 81.300 189.900 ;
        RECT 80.600 188.900 81.300 189.200 ;
        RECT 75.800 188.500 76.200 188.900 ;
        RECT 78.600 188.600 78.900 188.900 ;
        RECT 76.600 188.200 77.000 188.600 ;
        RECT 77.500 188.300 78.900 188.600 ;
        RECT 80.600 188.500 81.000 188.900 ;
        RECT 77.500 188.200 77.900 188.300 ;
        RECT 74.600 187.100 75.400 187.200 ;
        RECT 76.700 187.100 77.000 188.200 ;
        RECT 81.500 187.700 81.900 187.800 ;
        RECT 83.000 187.700 83.400 189.900 ;
        RECT 81.500 187.400 83.400 187.700 ;
        RECT 79.500 187.100 79.900 187.200 ;
        RECT 74.600 186.800 80.100 187.100 ;
        RECT 76.100 186.700 76.500 186.800 ;
        RECT 71.000 185.800 73.000 186.100 ;
        RECT 75.300 186.200 75.700 186.300 ;
        RECT 76.600 186.200 77.000 186.300 ;
        RECT 79.800 186.200 80.100 186.800 ;
        RECT 80.600 186.400 81.000 186.500 ;
        RECT 75.300 185.900 77.800 186.200 ;
        RECT 77.400 185.800 77.800 185.900 ;
        RECT 79.800 185.800 80.200 186.200 ;
        RECT 80.600 186.100 82.500 186.400 ;
        RECT 82.100 186.000 82.500 186.100 ;
        RECT 71.000 185.400 71.400 185.800 ;
        RECT 69.900 184.600 70.700 184.900 ;
        RECT 67.800 181.500 68.200 183.500 ;
        RECT 69.900 181.100 70.300 184.600 ;
        RECT 72.600 181.100 73.000 185.800 ;
        RECT 74.200 185.500 77.000 185.600 ;
        RECT 74.200 185.400 77.100 185.500 ;
        RECT 74.200 185.300 79.100 185.400 ;
        RECT 74.200 181.100 74.600 185.300 ;
        RECT 76.700 185.100 79.100 185.300 ;
        RECT 75.800 184.500 78.500 184.800 ;
        RECT 75.800 184.400 76.200 184.500 ;
        RECT 78.100 184.400 78.500 184.500 ;
        RECT 78.800 184.500 79.100 185.100 ;
        RECT 79.800 185.200 80.100 185.800 ;
        RECT 81.300 185.700 81.700 185.800 ;
        RECT 83.000 185.700 83.400 187.400 ;
        RECT 83.800 188.500 84.200 189.500 ;
        RECT 83.800 187.400 84.100 188.500 ;
        RECT 85.900 188.000 86.300 189.500 ;
        RECT 85.900 187.700 86.700 188.000 ;
        RECT 88.600 187.800 89.000 188.600 ;
        RECT 86.300 187.500 86.700 187.700 ;
        RECT 83.800 187.100 85.900 187.400 ;
        RECT 85.400 186.900 85.900 187.100 ;
        RECT 86.400 187.200 86.700 187.500 ;
        RECT 83.800 185.800 84.200 186.600 ;
        RECT 84.600 185.800 85.000 186.600 ;
        RECT 85.400 186.500 86.100 186.900 ;
        RECT 86.400 186.800 87.400 187.200 ;
        RECT 81.300 185.400 83.400 185.700 ;
        RECT 85.400 185.500 85.700 186.500 ;
        RECT 79.800 184.900 81.000 185.200 ;
        RECT 79.500 184.500 79.900 184.600 ;
        RECT 78.800 184.200 79.900 184.500 ;
        RECT 80.700 184.400 81.000 184.900 ;
        RECT 80.700 184.000 81.400 184.400 ;
        RECT 77.500 183.700 77.900 183.800 ;
        RECT 78.900 183.700 79.300 183.800 ;
        RECT 75.800 183.100 76.200 183.500 ;
        RECT 77.500 183.400 79.300 183.700 ;
        RECT 78.600 183.100 78.900 183.400 ;
        RECT 80.600 183.100 81.000 183.500 ;
        RECT 75.800 182.800 76.800 183.100 ;
        RECT 76.400 181.100 76.800 182.800 ;
        RECT 78.600 181.100 79.000 183.100 ;
        RECT 80.700 181.100 81.300 183.100 ;
        RECT 83.000 181.100 83.400 185.400 ;
        RECT 83.800 185.200 85.700 185.500 ;
        RECT 83.800 183.500 84.100 185.200 ;
        RECT 86.400 184.900 86.700 186.800 ;
        RECT 87.000 185.400 87.400 186.200 ;
        RECT 89.400 186.100 89.800 189.900 ;
        RECT 92.100 188.000 92.500 189.500 ;
        RECT 94.200 188.500 94.600 189.500 ;
        RECT 91.700 187.700 92.500 188.000 ;
        RECT 91.700 187.500 92.100 187.700 ;
        RECT 91.700 187.200 92.000 187.500 ;
        RECT 94.300 187.400 94.600 188.500 ;
        RECT 96.900 188.000 97.300 189.500 ;
        RECT 99.000 188.500 99.400 189.500 ;
        RECT 91.000 186.800 92.000 187.200 ;
        RECT 92.500 187.100 94.600 187.400 ;
        RECT 96.500 187.700 97.300 188.000 ;
        RECT 96.500 187.500 96.900 187.700 ;
        RECT 96.500 187.200 96.800 187.500 ;
        RECT 99.100 187.400 99.400 188.500 ;
        RECT 101.700 188.000 102.100 189.500 ;
        RECT 103.800 188.500 104.200 189.500 ;
        RECT 92.500 186.900 93.000 187.100 ;
        RECT 91.000 186.100 91.400 186.200 ;
        RECT 89.400 185.800 91.400 186.100 ;
        RECT 85.900 184.600 86.700 184.900 ;
        RECT 83.800 181.500 84.200 183.500 ;
        RECT 85.900 182.200 86.300 184.600 ;
        RECT 85.900 181.800 86.600 182.200 ;
        RECT 85.900 181.100 86.300 181.800 ;
        RECT 89.400 181.100 89.800 185.800 ;
        RECT 91.000 185.400 91.400 185.800 ;
        RECT 91.700 184.900 92.000 186.800 ;
        RECT 92.300 186.500 93.000 186.900 ;
        RECT 95.800 186.800 96.800 187.200 ;
        RECT 97.300 187.100 99.400 187.400 ;
        RECT 101.300 187.700 102.100 188.000 ;
        RECT 101.300 187.500 101.700 187.700 ;
        RECT 101.300 187.200 101.600 187.500 ;
        RECT 103.900 187.400 104.200 188.500 ;
        RECT 97.300 186.900 97.800 187.100 ;
        RECT 92.700 185.500 93.000 186.500 ;
        RECT 93.400 185.800 93.800 186.600 ;
        RECT 94.200 185.800 94.600 186.600 ;
        RECT 95.000 186.100 95.400 186.200 ;
        RECT 95.800 186.100 96.200 186.200 ;
        RECT 95.000 185.800 96.200 186.100 ;
        RECT 92.700 185.200 94.600 185.500 ;
        RECT 95.800 185.400 96.200 185.800 ;
        RECT 91.700 184.600 92.500 184.900 ;
        RECT 92.100 182.200 92.500 184.600 ;
        RECT 94.300 183.500 94.600 185.200 ;
        RECT 96.500 184.900 96.800 186.800 ;
        RECT 97.100 186.500 97.800 186.900 ;
        RECT 100.600 186.800 101.600 187.200 ;
        RECT 102.100 187.100 104.200 187.400 ;
        RECT 106.200 187.700 106.600 189.900 ;
        RECT 108.300 189.200 108.900 189.900 ;
        RECT 108.300 188.900 109.000 189.200 ;
        RECT 110.600 188.900 111.000 189.900 ;
        RECT 112.800 189.200 113.200 189.900 ;
        RECT 112.800 188.900 113.800 189.200 ;
        RECT 108.600 188.500 109.000 188.900 ;
        RECT 110.700 188.600 111.000 188.900 ;
        RECT 110.700 188.300 112.100 188.600 ;
        RECT 111.700 188.200 112.100 188.300 ;
        RECT 112.600 188.200 113.000 188.600 ;
        RECT 113.400 188.500 113.800 188.900 ;
        RECT 107.700 187.700 108.100 187.800 ;
        RECT 106.200 187.400 108.100 187.700 ;
        RECT 102.100 186.900 102.600 187.100 ;
        RECT 97.500 185.500 97.800 186.500 ;
        RECT 98.200 185.800 98.600 186.600 ;
        RECT 99.000 185.800 99.400 186.600 ;
        RECT 97.500 185.200 99.400 185.500 ;
        RECT 100.600 185.400 101.000 186.200 ;
        RECT 96.500 184.600 97.300 184.900 ;
        RECT 91.800 181.800 92.500 182.200 ;
        RECT 92.100 181.100 92.500 181.800 ;
        RECT 94.200 181.500 94.600 183.500 ;
        RECT 96.900 182.200 97.300 184.600 ;
        RECT 99.100 183.500 99.400 185.200 ;
        RECT 101.300 184.900 101.600 186.800 ;
        RECT 101.900 186.500 102.600 186.900 ;
        RECT 102.300 185.500 102.600 186.500 ;
        RECT 103.000 185.800 103.400 186.600 ;
        RECT 103.800 186.100 104.200 186.600 ;
        RECT 104.600 186.100 105.000 186.200 ;
        RECT 103.800 185.800 105.000 186.100 ;
        RECT 106.200 185.700 106.600 187.400 ;
        RECT 109.700 187.100 110.100 187.200 ;
        RECT 112.600 187.100 112.900 188.200 ;
        RECT 115.000 187.500 115.400 189.900 ;
        RECT 117.100 188.200 117.500 189.900 ;
        RECT 116.600 187.900 117.500 188.200 ;
        RECT 118.200 187.900 118.600 189.900 ;
        RECT 119.000 188.000 119.400 189.900 ;
        RECT 120.600 188.000 121.000 189.900 ;
        RECT 119.000 187.900 121.000 188.000 ;
        RECT 114.200 187.100 115.000 187.200 ;
        RECT 109.500 186.800 115.000 187.100 ;
        RECT 115.800 186.800 116.200 187.600 ;
        RECT 108.600 186.400 109.000 186.500 ;
        RECT 107.100 186.100 109.000 186.400 ;
        RECT 109.500 186.200 109.800 186.800 ;
        RECT 113.100 186.700 113.500 186.800 ;
        RECT 112.600 186.200 113.000 186.300 ;
        RECT 113.900 186.200 114.300 186.300 ;
        RECT 107.100 186.000 107.500 186.100 ;
        RECT 109.400 185.800 109.800 186.200 ;
        RECT 111.800 185.900 114.300 186.200 ;
        RECT 116.600 186.100 117.000 187.900 ;
        RECT 118.300 187.200 118.600 187.900 ;
        RECT 119.100 187.700 120.900 187.900 ;
        RECT 122.200 187.600 122.600 189.900 ;
        RECT 123.800 187.600 124.200 189.900 ;
        RECT 125.400 187.600 125.800 189.900 ;
        RECT 127.000 187.600 127.400 189.900 ;
        RECT 120.200 187.200 120.600 187.400 ;
        RECT 122.200 187.200 123.100 187.600 ;
        RECT 123.800 187.200 124.900 187.600 ;
        RECT 125.400 187.200 126.500 187.600 ;
        RECT 127.000 187.200 128.200 187.600 ;
        RECT 128.600 187.500 129.000 189.900 ;
        RECT 130.800 189.200 131.200 189.900 ;
        RECT 130.200 188.900 131.200 189.200 ;
        RECT 133.000 188.900 133.400 189.900 ;
        RECT 135.100 189.200 135.700 189.900 ;
        RECT 135.000 188.900 135.700 189.200 ;
        RECT 130.200 188.500 130.600 188.900 ;
        RECT 133.000 188.600 133.300 188.900 ;
        RECT 131.000 187.800 131.400 188.600 ;
        RECT 131.900 188.300 133.300 188.600 ;
        RECT 135.000 188.500 135.400 188.900 ;
        RECT 131.900 188.200 132.300 188.300 ;
        RECT 117.400 187.100 117.800 187.200 ;
        RECT 118.200 187.100 119.500 187.200 ;
        RECT 117.400 186.800 119.500 187.100 ;
        RECT 120.200 186.900 121.000 187.200 ;
        RECT 120.600 186.800 121.000 186.900 ;
        RECT 121.400 186.900 121.800 187.200 ;
        RECT 122.700 186.900 123.100 187.200 ;
        RECT 124.500 186.900 124.900 187.200 ;
        RECT 126.100 186.900 126.500 187.200 ;
        RECT 111.800 185.800 112.200 185.900 ;
        RECT 116.600 185.800 118.500 186.100 ;
        RECT 107.900 185.700 108.300 185.800 ;
        RECT 102.300 185.200 104.200 185.500 ;
        RECT 101.300 184.600 102.100 184.900 ;
        RECT 96.900 181.800 97.800 182.200 ;
        RECT 96.900 181.100 97.300 181.800 ;
        RECT 99.000 181.500 99.400 183.500 ;
        RECT 101.700 182.200 102.100 184.600 ;
        RECT 103.900 183.500 104.200 185.200 ;
        RECT 101.400 181.800 102.100 182.200 ;
        RECT 101.700 181.100 102.100 181.800 ;
        RECT 103.800 181.500 104.200 183.500 ;
        RECT 106.200 185.400 108.300 185.700 ;
        RECT 106.200 181.100 106.600 185.400 ;
        RECT 109.500 185.200 109.800 185.800 ;
        RECT 112.600 185.500 115.400 185.600 ;
        RECT 112.500 185.400 115.400 185.500 ;
        RECT 108.600 184.900 109.800 185.200 ;
        RECT 110.500 185.300 115.400 185.400 ;
        RECT 110.500 185.100 112.900 185.300 ;
        RECT 108.600 184.400 108.900 184.900 ;
        RECT 108.200 184.000 108.900 184.400 ;
        RECT 109.700 184.500 110.100 184.600 ;
        RECT 110.500 184.500 110.800 185.100 ;
        RECT 109.700 184.200 110.800 184.500 ;
        RECT 111.100 184.500 113.800 184.800 ;
        RECT 111.100 184.400 111.500 184.500 ;
        RECT 113.400 184.400 113.800 184.500 ;
        RECT 110.300 183.700 110.700 183.800 ;
        RECT 111.700 183.700 112.100 183.800 ;
        RECT 108.600 183.100 109.000 183.500 ;
        RECT 110.300 183.400 112.100 183.700 ;
        RECT 110.700 183.100 111.000 183.400 ;
        RECT 113.400 183.100 113.800 183.500 ;
        RECT 108.300 181.100 108.900 183.100 ;
        RECT 110.600 181.100 111.000 183.100 ;
        RECT 112.800 182.800 113.800 183.100 ;
        RECT 112.800 181.100 113.200 182.800 ;
        RECT 115.000 181.100 115.400 185.300 ;
        RECT 116.600 181.100 117.000 185.800 ;
        RECT 118.200 185.200 118.500 185.800 ;
        RECT 117.400 184.400 117.800 185.200 ;
        RECT 118.200 185.100 118.600 185.200 ;
        RECT 119.200 185.100 119.500 186.800 ;
        RECT 119.800 185.800 120.200 186.600 ;
        RECT 121.400 186.500 122.300 186.900 ;
        RECT 122.700 186.500 124.000 186.900 ;
        RECT 124.500 186.500 125.700 186.900 ;
        RECT 126.100 186.500 127.400 186.900 ;
        RECT 122.700 185.800 123.100 186.500 ;
        RECT 124.500 185.800 124.900 186.500 ;
        RECT 126.100 185.800 126.500 186.500 ;
        RECT 127.800 185.800 128.200 187.200 ;
        RECT 129.000 187.100 129.800 187.200 ;
        RECT 131.100 187.100 131.400 187.800 ;
        RECT 135.900 187.700 136.300 187.800 ;
        RECT 137.400 187.700 137.800 189.900 ;
        RECT 138.200 188.000 138.600 189.900 ;
        RECT 139.800 188.000 140.200 189.900 ;
        RECT 138.200 187.900 140.200 188.000 ;
        RECT 140.600 187.900 141.000 189.900 ;
        RECT 141.700 188.200 142.100 189.900 ;
        RECT 141.700 187.900 142.600 188.200 ;
        RECT 138.300 187.700 140.100 187.900 ;
        RECT 135.900 187.400 137.800 187.700 ;
        RECT 133.900 187.100 134.300 187.200 ;
        RECT 129.000 186.800 134.500 187.100 ;
        RECT 130.500 186.700 130.900 186.800 ;
        RECT 129.700 186.200 130.100 186.300 ;
        RECT 129.700 185.900 132.200 186.200 ;
        RECT 131.800 185.800 132.200 185.900 ;
        RECT 122.200 185.400 123.100 185.800 ;
        RECT 123.800 185.400 124.900 185.800 ;
        RECT 125.400 185.400 126.500 185.800 ;
        RECT 127.000 185.400 128.200 185.800 ;
        RECT 128.600 185.500 131.400 185.600 ;
        RECT 128.600 185.400 131.500 185.500 ;
        RECT 118.200 184.800 118.900 185.100 ;
        RECT 119.200 184.800 119.700 185.100 ;
        RECT 118.600 184.200 118.900 184.800 ;
        RECT 118.600 183.800 119.000 184.200 ;
        RECT 119.300 181.100 119.700 184.800 ;
        RECT 122.200 181.100 122.600 185.400 ;
        RECT 123.800 181.100 124.200 185.400 ;
        RECT 125.400 181.100 125.800 185.400 ;
        RECT 127.000 181.100 127.400 185.400 ;
        RECT 128.600 185.300 133.500 185.400 ;
        RECT 128.600 181.100 129.000 185.300 ;
        RECT 131.100 185.100 133.500 185.300 ;
        RECT 130.200 184.500 132.900 184.800 ;
        RECT 130.200 184.400 130.600 184.500 ;
        RECT 132.500 184.400 132.900 184.500 ;
        RECT 133.200 184.500 133.500 185.100 ;
        RECT 134.200 185.200 134.500 186.800 ;
        RECT 135.000 186.400 135.400 186.500 ;
        RECT 135.000 186.100 136.900 186.400 ;
        RECT 136.500 186.000 136.900 186.100 ;
        RECT 135.700 185.700 136.100 185.800 ;
        RECT 137.400 185.700 137.800 187.400 ;
        RECT 138.600 187.200 139.000 187.400 ;
        RECT 140.600 187.200 140.900 187.900 ;
        RECT 138.200 186.900 139.000 187.200 ;
        RECT 138.200 186.800 138.600 186.900 ;
        RECT 139.700 186.800 141.000 187.200 ;
        RECT 139.000 185.800 139.400 186.600 ;
        RECT 139.700 186.200 140.000 186.800 ;
        RECT 139.700 185.800 140.200 186.200 ;
        RECT 142.200 186.100 142.600 187.900 ;
        RECT 143.000 186.800 143.400 187.600 ;
        RECT 143.800 187.500 144.200 189.900 ;
        RECT 146.000 189.200 146.400 189.900 ;
        RECT 145.400 188.900 146.400 189.200 ;
        RECT 148.200 188.900 148.600 189.900 ;
        RECT 150.300 189.200 150.900 189.900 ;
        RECT 150.200 188.900 150.900 189.200 ;
        RECT 145.400 188.500 145.800 188.900 ;
        RECT 148.200 188.600 148.500 188.900 ;
        RECT 146.200 187.800 146.600 188.600 ;
        RECT 147.100 188.300 148.500 188.600 ;
        RECT 150.200 188.500 150.600 188.900 ;
        RECT 147.100 188.200 147.500 188.300 ;
        RECT 144.200 187.100 145.000 187.200 ;
        RECT 146.300 187.100 146.600 187.800 ;
        RECT 151.100 187.700 151.500 187.800 ;
        RECT 152.600 187.700 153.000 189.900 ;
        RECT 151.100 187.400 153.000 187.700 ;
        RECT 155.000 187.500 155.400 189.900 ;
        RECT 157.200 189.200 157.600 189.900 ;
        RECT 156.600 188.900 157.600 189.200 ;
        RECT 159.400 188.900 159.800 189.900 ;
        RECT 161.500 189.200 162.100 189.900 ;
        RECT 161.400 188.900 162.100 189.200 ;
        RECT 156.600 188.500 157.000 188.900 ;
        RECT 159.400 188.600 159.700 188.900 ;
        RECT 157.400 188.200 157.800 188.600 ;
        RECT 158.300 188.300 159.700 188.600 ;
        RECT 161.400 188.500 161.800 188.900 ;
        RECT 158.300 188.200 158.700 188.300 ;
        RECT 149.100 187.100 149.500 187.200 ;
        RECT 144.200 186.800 149.700 187.100 ;
        RECT 151.800 186.800 152.200 187.400 ;
        RECT 145.700 186.700 146.100 186.800 ;
        RECT 140.600 185.800 142.600 186.100 ;
        RECT 144.900 186.200 145.300 186.300 ;
        RECT 144.900 185.900 147.400 186.200 ;
        RECT 147.000 185.800 147.400 185.900 ;
        RECT 135.700 185.400 137.800 185.700 ;
        RECT 134.200 184.900 135.400 185.200 ;
        RECT 133.900 184.500 134.300 184.600 ;
        RECT 133.200 184.200 134.300 184.500 ;
        RECT 135.100 184.400 135.400 184.900 ;
        RECT 135.100 184.000 135.800 184.400 ;
        RECT 131.900 183.700 132.300 183.800 ;
        RECT 133.300 183.700 133.700 183.800 ;
        RECT 130.200 183.100 130.600 183.500 ;
        RECT 131.900 183.400 133.700 183.700 ;
        RECT 133.000 183.100 133.300 183.400 ;
        RECT 135.000 183.100 135.400 183.500 ;
        RECT 130.200 182.800 131.200 183.100 ;
        RECT 130.800 181.100 131.200 182.800 ;
        RECT 133.000 181.100 133.400 183.100 ;
        RECT 135.100 181.100 135.700 183.100 ;
        RECT 137.400 181.100 137.800 185.400 ;
        RECT 139.700 185.100 140.000 185.800 ;
        RECT 140.600 185.200 140.900 185.800 ;
        RECT 140.600 185.100 141.000 185.200 ;
        RECT 139.500 184.800 140.000 185.100 ;
        RECT 140.300 184.800 141.000 185.100 ;
        RECT 139.500 181.100 139.900 184.800 ;
        RECT 140.300 184.200 140.600 184.800 ;
        RECT 141.400 184.400 141.800 185.200 ;
        RECT 140.200 183.800 140.600 184.200 ;
        RECT 142.200 181.100 142.600 185.800 ;
        RECT 143.800 185.500 146.600 185.600 ;
        RECT 143.800 185.400 146.700 185.500 ;
        RECT 143.800 185.300 148.700 185.400 ;
        RECT 143.800 181.100 144.200 185.300 ;
        RECT 146.300 185.100 148.700 185.300 ;
        RECT 145.400 184.500 148.100 184.800 ;
        RECT 145.400 184.400 145.800 184.500 ;
        RECT 147.700 184.400 148.100 184.500 ;
        RECT 148.400 184.500 148.700 185.100 ;
        RECT 149.400 185.200 149.700 186.800 ;
        RECT 150.200 186.400 150.600 186.500 ;
        RECT 150.200 186.100 152.100 186.400 ;
        RECT 151.700 186.000 152.100 186.100 ;
        RECT 150.900 185.700 151.300 185.800 ;
        RECT 152.600 185.700 153.000 187.400 ;
        RECT 155.400 187.100 156.200 187.200 ;
        RECT 157.500 187.100 157.800 188.200 ;
        RECT 162.300 187.700 162.700 187.800 ;
        RECT 163.800 187.700 164.200 189.900 ;
        RECT 164.600 187.800 165.000 188.600 ;
        RECT 162.300 187.400 164.200 187.700 ;
        RECT 160.300 187.100 160.700 187.200 ;
        RECT 155.400 186.800 160.900 187.100 ;
        RECT 156.900 186.700 157.300 186.800 ;
        RECT 156.100 186.200 156.500 186.300 ;
        RECT 156.100 186.100 158.600 186.200 ;
        RECT 159.800 186.100 160.200 186.200 ;
        RECT 156.100 185.900 160.200 186.100 ;
        RECT 158.200 185.800 160.200 185.900 ;
        RECT 150.900 185.400 153.000 185.700 ;
        RECT 149.400 184.900 150.600 185.200 ;
        RECT 149.100 184.500 149.500 184.600 ;
        RECT 148.400 184.200 149.500 184.500 ;
        RECT 150.300 184.400 150.600 184.900 ;
        RECT 150.300 184.000 151.000 184.400 ;
        RECT 147.100 183.700 147.500 183.800 ;
        RECT 148.500 183.700 148.900 183.800 ;
        RECT 145.400 183.100 145.800 183.500 ;
        RECT 147.100 183.400 148.900 183.700 ;
        RECT 148.200 183.100 148.500 183.400 ;
        RECT 150.200 183.100 150.600 183.500 ;
        RECT 145.400 182.800 146.400 183.100 ;
        RECT 146.000 181.100 146.400 182.800 ;
        RECT 148.200 181.100 148.600 183.100 ;
        RECT 150.300 181.100 150.900 183.100 ;
        RECT 152.600 181.100 153.000 185.400 ;
        RECT 155.000 185.500 157.800 185.600 ;
        RECT 155.000 185.400 157.900 185.500 ;
        RECT 155.000 185.300 159.900 185.400 ;
        RECT 155.000 181.100 155.400 185.300 ;
        RECT 157.500 185.100 159.900 185.300 ;
        RECT 156.600 184.500 159.300 184.800 ;
        RECT 156.600 184.400 157.000 184.500 ;
        RECT 158.900 184.400 159.300 184.500 ;
        RECT 159.600 184.500 159.900 185.100 ;
        RECT 160.600 185.200 160.900 186.800 ;
        RECT 161.400 186.400 161.800 186.500 ;
        RECT 161.400 186.100 163.300 186.400 ;
        RECT 162.900 186.000 163.300 186.100 ;
        RECT 162.100 185.700 162.500 185.800 ;
        RECT 163.800 185.700 164.200 187.400 ;
        RECT 162.100 185.400 164.200 185.700 ;
        RECT 160.600 184.900 161.800 185.200 ;
        RECT 160.300 184.500 160.700 184.600 ;
        RECT 159.600 184.200 160.700 184.500 ;
        RECT 161.500 184.400 161.800 184.900 ;
        RECT 161.500 184.200 162.200 184.400 ;
        RECT 161.500 184.000 162.600 184.200 ;
        RECT 161.900 183.800 162.600 184.000 ;
        RECT 158.300 183.700 158.700 183.800 ;
        RECT 159.700 183.700 160.100 183.800 ;
        RECT 156.600 183.100 157.000 183.500 ;
        RECT 158.300 183.400 160.100 183.700 ;
        RECT 159.400 183.100 159.700 183.400 ;
        RECT 161.400 183.100 161.800 183.500 ;
        RECT 156.600 182.800 157.600 183.100 ;
        RECT 157.200 181.100 157.600 182.800 ;
        RECT 159.400 181.100 159.800 183.100 ;
        RECT 161.500 181.100 162.100 183.100 ;
        RECT 163.800 181.100 164.200 185.400 ;
        RECT 165.400 186.100 165.800 189.900 ;
        RECT 168.100 188.000 168.500 189.500 ;
        RECT 170.200 188.500 170.600 189.500 ;
        RECT 167.700 187.700 168.500 188.000 ;
        RECT 167.700 187.500 168.100 187.700 ;
        RECT 167.700 187.200 168.000 187.500 ;
        RECT 170.300 187.400 170.600 188.500 ;
        RECT 172.900 188.000 173.300 189.500 ;
        RECT 175.000 188.500 175.400 189.500 ;
        RECT 166.200 187.100 166.600 187.200 ;
        RECT 167.000 187.100 168.000 187.200 ;
        RECT 166.200 186.800 168.000 187.100 ;
        RECT 168.500 187.100 170.600 187.400 ;
        RECT 172.500 187.700 173.300 188.000 ;
        RECT 172.500 187.500 172.900 187.700 ;
        RECT 172.500 187.200 172.800 187.500 ;
        RECT 175.100 187.400 175.400 188.500 ;
        RECT 168.500 186.900 169.000 187.100 ;
        RECT 167.000 186.100 167.400 186.200 ;
        RECT 165.400 185.800 167.400 186.100 ;
        RECT 165.400 181.100 165.800 185.800 ;
        RECT 167.000 185.400 167.400 185.800 ;
        RECT 167.700 184.900 168.000 186.800 ;
        RECT 168.300 186.500 169.000 186.900 ;
        RECT 171.800 186.800 172.800 187.200 ;
        RECT 173.300 187.100 175.400 187.400 ;
        RECT 175.800 188.500 176.200 189.500 ;
        RECT 175.800 187.400 176.100 188.500 ;
        RECT 177.900 188.000 178.300 189.500 ;
        RECT 180.600 188.500 181.000 189.500 ;
        RECT 177.900 187.700 178.700 188.000 ;
        RECT 178.300 187.500 178.700 187.700 ;
        RECT 175.800 187.100 177.900 187.400 ;
        RECT 173.300 186.900 173.800 187.100 ;
        RECT 168.700 185.500 169.000 186.500 ;
        RECT 169.400 185.800 169.800 186.600 ;
        RECT 170.200 185.800 170.600 186.600 ;
        RECT 171.000 186.100 171.400 186.200 ;
        RECT 171.800 186.100 172.200 186.200 ;
        RECT 171.000 185.800 172.200 186.100 ;
        RECT 168.700 185.200 170.600 185.500 ;
        RECT 171.800 185.400 172.200 185.800 ;
        RECT 167.700 184.600 168.500 184.900 ;
        RECT 168.100 181.100 168.500 184.600 ;
        RECT 170.300 183.500 170.600 185.200 ;
        RECT 172.500 184.900 172.800 186.800 ;
        RECT 173.100 186.500 173.800 186.900 ;
        RECT 177.400 186.900 177.900 187.100 ;
        RECT 178.400 187.200 178.700 187.500 ;
        RECT 180.600 187.400 180.900 188.500 ;
        RECT 182.700 188.000 183.100 189.500 ;
        RECT 182.700 187.700 183.500 188.000 ;
        RECT 183.100 187.500 183.500 187.700 ;
        RECT 173.500 185.500 173.800 186.500 ;
        RECT 174.200 185.800 174.600 186.600 ;
        RECT 175.000 185.800 175.400 186.600 ;
        RECT 175.800 185.800 176.200 186.600 ;
        RECT 176.600 185.800 177.000 186.600 ;
        RECT 177.400 186.500 178.100 186.900 ;
        RECT 178.400 186.800 179.400 187.200 ;
        RECT 180.600 187.100 182.700 187.400 ;
        RECT 182.200 186.900 182.700 187.100 ;
        RECT 183.200 187.200 183.500 187.500 ;
        RECT 185.400 187.600 185.800 189.900 ;
        RECT 187.000 188.200 187.400 189.900 ;
        RECT 188.600 188.500 189.000 189.500 ;
        RECT 187.000 187.900 187.500 188.200 ;
        RECT 185.400 187.300 186.700 187.600 ;
        RECT 177.400 185.500 177.700 186.500 ;
        RECT 173.500 185.200 175.400 185.500 ;
        RECT 172.500 184.600 173.300 184.900 ;
        RECT 170.200 181.500 170.600 183.500 ;
        RECT 172.900 182.200 173.300 184.600 ;
        RECT 175.100 183.500 175.400 185.200 ;
        RECT 172.900 181.800 173.800 182.200 ;
        RECT 172.900 181.100 173.300 181.800 ;
        RECT 175.000 181.500 175.400 183.500 ;
        RECT 175.800 185.200 177.700 185.500 ;
        RECT 175.800 183.500 176.100 185.200 ;
        RECT 178.400 184.900 178.700 186.800 ;
        RECT 179.000 185.400 179.400 186.200 ;
        RECT 179.800 186.100 180.200 186.200 ;
        RECT 180.600 186.100 181.000 186.600 ;
        RECT 179.800 185.800 181.000 186.100 ;
        RECT 181.400 185.800 181.800 186.600 ;
        RECT 182.200 186.500 182.900 186.900 ;
        RECT 183.200 186.800 184.200 187.200 ;
        RECT 182.200 185.500 182.500 186.500 ;
        RECT 177.900 184.600 178.700 184.900 ;
        RECT 180.600 185.200 182.500 185.500 ;
        RECT 175.800 181.500 176.200 183.500 ;
        RECT 177.900 182.200 178.300 184.600 ;
        RECT 180.600 183.500 180.900 185.200 ;
        RECT 183.200 184.900 183.500 186.800 ;
        RECT 185.500 186.200 185.900 186.600 ;
        RECT 183.800 185.400 184.200 186.200 ;
        RECT 185.400 185.800 185.900 186.200 ;
        RECT 186.400 186.500 186.700 187.300 ;
        RECT 187.200 187.200 187.500 187.900 ;
        RECT 187.000 186.800 187.500 187.200 ;
        RECT 188.600 187.400 188.900 188.500 ;
        RECT 190.700 188.000 191.100 189.500 ;
        RECT 195.300 188.000 195.700 189.500 ;
        RECT 197.400 188.500 197.800 189.500 ;
        RECT 190.700 187.700 191.500 188.000 ;
        RECT 191.100 187.500 191.500 187.700 ;
        RECT 188.600 187.100 190.700 187.400 ;
        RECT 186.400 186.100 186.900 186.500 ;
        RECT 186.400 185.100 186.700 186.100 ;
        RECT 187.200 185.100 187.500 186.800 ;
        RECT 190.200 186.900 190.700 187.100 ;
        RECT 191.200 187.200 191.500 187.500 ;
        RECT 194.900 187.700 195.700 188.000 ;
        RECT 194.900 187.500 195.300 187.700 ;
        RECT 194.900 187.200 195.200 187.500 ;
        RECT 197.500 187.400 197.800 188.500 ;
        RECT 200.100 188.200 200.500 189.500 ;
        RECT 202.200 188.500 202.600 189.500 ;
        RECT 200.100 188.000 201.000 188.200 ;
        RECT 191.200 187.100 192.200 187.200 ;
        RECT 188.600 185.800 189.000 186.600 ;
        RECT 189.400 185.800 189.800 186.600 ;
        RECT 190.200 186.500 190.900 186.900 ;
        RECT 191.200 186.800 193.700 187.100 ;
        RECT 194.200 186.800 195.200 187.200 ;
        RECT 195.700 187.100 197.800 187.400 ;
        RECT 199.700 187.800 201.000 188.000 ;
        RECT 199.700 187.700 200.500 187.800 ;
        RECT 199.700 187.500 200.100 187.700 ;
        RECT 199.700 187.200 200.000 187.500 ;
        RECT 202.300 187.400 202.600 188.500 ;
        RECT 195.700 186.900 196.200 187.100 ;
        RECT 190.200 185.500 190.500 186.500 ;
        RECT 182.700 184.600 183.500 184.900 ;
        RECT 185.400 184.800 186.700 185.100 ;
        RECT 177.900 181.800 178.600 182.200 ;
        RECT 177.900 181.100 178.300 181.800 ;
        RECT 180.600 181.500 181.000 183.500 ;
        RECT 182.700 182.200 183.100 184.600 ;
        RECT 182.200 181.800 183.100 182.200 ;
        RECT 182.700 181.100 183.100 181.800 ;
        RECT 185.400 181.100 185.800 184.800 ;
        RECT 187.000 184.600 187.500 185.100 ;
        RECT 188.600 185.200 190.500 185.500 ;
        RECT 187.000 181.100 187.400 184.600 ;
        RECT 188.600 183.500 188.900 185.200 ;
        RECT 191.200 184.900 191.500 186.800 ;
        RECT 191.800 185.400 192.200 186.200 ;
        RECT 193.400 186.100 193.700 186.800 ;
        RECT 194.200 186.100 194.600 186.200 ;
        RECT 193.400 185.800 194.600 186.100 ;
        RECT 194.200 185.400 194.600 185.800 ;
        RECT 190.700 184.600 191.500 184.900 ;
        RECT 194.900 184.900 195.200 186.800 ;
        RECT 195.500 186.500 196.200 186.900 ;
        RECT 199.000 186.800 200.000 187.200 ;
        RECT 200.500 187.100 202.600 187.400 ;
        RECT 203.000 188.500 203.400 189.500 ;
        RECT 203.000 187.400 203.300 188.500 ;
        RECT 205.100 188.000 205.500 189.500 ;
        RECT 209.400 188.500 209.800 189.500 ;
        RECT 205.100 187.700 205.900 188.000 ;
        RECT 205.500 187.500 205.900 187.700 ;
        RECT 203.000 187.100 205.100 187.400 ;
        RECT 200.500 186.900 201.000 187.100 ;
        RECT 195.900 185.500 196.200 186.500 ;
        RECT 196.600 185.800 197.000 186.600 ;
        RECT 197.400 185.800 197.800 186.600 ;
        RECT 195.900 185.200 197.800 185.500 ;
        RECT 199.000 185.400 199.400 186.200 ;
        RECT 194.900 184.600 195.700 184.900 ;
        RECT 188.600 181.500 189.000 183.500 ;
        RECT 190.700 181.100 191.100 184.600 ;
        RECT 195.300 182.200 195.700 184.600 ;
        RECT 197.500 183.500 197.800 185.200 ;
        RECT 199.700 184.900 200.000 186.800 ;
        RECT 200.300 186.500 201.000 186.900 ;
        RECT 204.600 186.900 205.100 187.100 ;
        RECT 205.600 187.200 205.900 187.500 ;
        RECT 209.400 187.400 209.700 188.500 ;
        RECT 211.500 188.000 211.900 189.500 ;
        RECT 214.200 188.500 214.600 189.500 ;
        RECT 211.500 187.700 212.300 188.000 ;
        RECT 211.900 187.500 212.300 187.700 ;
        RECT 200.700 185.500 201.000 186.500 ;
        RECT 201.400 185.800 201.800 186.600 ;
        RECT 202.200 185.800 202.600 186.600 ;
        RECT 203.000 185.800 203.400 186.600 ;
        RECT 203.800 185.800 204.200 186.600 ;
        RECT 204.600 186.500 205.300 186.900 ;
        RECT 205.600 186.800 206.600 187.200 ;
        RECT 209.400 187.100 211.500 187.400 ;
        RECT 211.000 186.900 211.500 187.100 ;
        RECT 212.000 187.200 212.300 187.500 ;
        RECT 214.200 187.400 214.500 188.500 ;
        RECT 216.300 188.000 216.700 189.500 ;
        RECT 216.300 187.700 217.100 188.000 ;
        RECT 216.700 187.500 217.100 187.700 ;
        RECT 219.000 187.500 219.400 189.900 ;
        RECT 221.200 189.200 221.600 189.900 ;
        RECT 220.600 188.900 221.600 189.200 ;
        RECT 223.400 188.900 223.800 189.900 ;
        RECT 225.500 189.200 226.100 189.900 ;
        RECT 225.400 188.900 226.100 189.200 ;
        RECT 220.600 188.500 221.000 188.900 ;
        RECT 223.400 188.600 223.700 188.900 ;
        RECT 221.400 188.200 221.800 188.600 ;
        RECT 222.300 188.300 223.700 188.600 ;
        RECT 225.400 188.500 225.800 188.900 ;
        RECT 222.300 188.200 222.700 188.300 ;
        RECT 212.000 187.100 213.000 187.200 ;
        RECT 213.400 187.100 213.800 187.200 ;
        RECT 214.200 187.100 216.300 187.400 ;
        RECT 204.600 185.500 204.900 186.500 ;
        RECT 200.700 185.200 202.600 185.500 ;
        RECT 199.700 184.600 200.500 184.900 ;
        RECT 195.300 181.800 196.200 182.200 ;
        RECT 195.300 181.100 195.700 181.800 ;
        RECT 197.400 181.500 197.800 183.500 ;
        RECT 200.100 181.100 200.500 184.600 ;
        RECT 202.300 183.500 202.600 185.200 ;
        RECT 202.200 181.500 202.600 183.500 ;
        RECT 203.000 185.200 204.900 185.500 ;
        RECT 203.000 183.500 203.300 185.200 ;
        RECT 205.600 184.900 205.900 186.800 ;
        RECT 206.200 185.400 206.600 186.200 ;
        RECT 209.400 185.800 209.800 186.600 ;
        RECT 210.200 185.800 210.600 186.600 ;
        RECT 211.000 186.500 211.700 186.900 ;
        RECT 212.000 186.800 213.800 187.100 ;
        RECT 215.800 186.900 216.300 187.100 ;
        RECT 216.800 187.200 217.100 187.500 ;
        RECT 211.000 185.500 211.300 186.500 ;
        RECT 205.100 184.600 205.900 184.900 ;
        RECT 209.400 185.200 211.300 185.500 ;
        RECT 203.000 181.500 203.400 183.500 ;
        RECT 205.100 182.200 205.500 184.600 ;
        RECT 209.400 183.500 209.700 185.200 ;
        RECT 212.000 184.900 212.300 186.800 ;
        RECT 212.600 185.400 213.000 186.200 ;
        RECT 214.200 185.800 214.600 186.600 ;
        RECT 215.000 185.800 215.400 186.600 ;
        RECT 215.800 186.500 216.500 186.900 ;
        RECT 216.800 186.800 217.800 187.200 ;
        RECT 219.400 187.100 220.200 187.200 ;
        RECT 221.500 187.100 221.800 188.200 ;
        RECT 226.300 187.700 226.700 187.800 ;
        RECT 227.800 187.700 228.200 189.900 ;
        RECT 230.500 188.000 230.900 189.500 ;
        RECT 232.600 188.500 233.000 189.500 ;
        RECT 226.300 187.400 228.200 187.700 ;
        RECT 222.200 187.100 222.600 187.200 ;
        RECT 224.300 187.100 224.700 187.200 ;
        RECT 219.400 186.800 224.900 187.100 ;
        RECT 215.800 185.500 216.100 186.500 ;
        RECT 211.500 184.600 212.300 184.900 ;
        RECT 214.200 185.200 216.100 185.500 ;
        RECT 205.100 181.800 205.800 182.200 ;
        RECT 205.100 181.100 205.500 181.800 ;
        RECT 209.400 181.500 209.800 183.500 ;
        RECT 211.500 181.100 211.900 184.600 ;
        RECT 214.200 183.500 214.500 185.200 ;
        RECT 216.800 184.900 217.100 186.800 ;
        RECT 220.900 186.700 221.300 186.800 ;
        RECT 220.100 186.200 220.500 186.300 ;
        RECT 224.600 186.200 224.900 186.800 ;
        RECT 225.400 186.400 225.800 186.500 ;
        RECT 217.400 185.400 217.800 186.200 ;
        RECT 220.100 186.100 222.600 186.200 ;
        RECT 223.800 186.100 224.200 186.200 ;
        RECT 220.100 185.900 224.200 186.100 ;
        RECT 222.200 185.800 224.200 185.900 ;
        RECT 224.600 185.800 225.000 186.200 ;
        RECT 225.400 186.100 227.300 186.400 ;
        RECT 226.900 186.000 227.300 186.100 ;
        RECT 219.000 185.500 221.800 185.600 ;
        RECT 219.000 185.400 221.900 185.500 ;
        RECT 216.300 184.600 217.100 184.900 ;
        RECT 219.000 185.300 223.900 185.400 ;
        RECT 214.200 181.500 214.600 183.500 ;
        RECT 216.300 182.200 216.700 184.600 ;
        RECT 216.300 181.800 217.000 182.200 ;
        RECT 216.300 181.100 216.700 181.800 ;
        RECT 219.000 181.100 219.400 185.300 ;
        RECT 221.500 185.100 223.900 185.300 ;
        RECT 220.600 184.500 223.300 184.800 ;
        RECT 220.600 184.400 221.000 184.500 ;
        RECT 222.900 184.400 223.300 184.500 ;
        RECT 223.600 184.500 223.900 185.100 ;
        RECT 224.600 185.200 224.900 185.800 ;
        RECT 226.100 185.700 226.500 185.800 ;
        RECT 227.800 185.700 228.200 187.400 ;
        RECT 230.100 187.700 230.900 188.000 ;
        RECT 230.100 187.500 230.500 187.700 ;
        RECT 230.100 187.200 230.400 187.500 ;
        RECT 232.700 187.400 233.000 188.500 ;
        RECT 235.300 188.000 235.700 189.500 ;
        RECT 237.400 188.500 237.800 189.500 ;
        RECT 229.400 186.800 230.400 187.200 ;
        RECT 230.900 187.100 233.000 187.400 ;
        RECT 234.900 187.700 235.700 188.000 ;
        RECT 234.900 187.500 235.300 187.700 ;
        RECT 234.900 187.200 235.200 187.500 ;
        RECT 237.500 187.400 237.800 188.500 ;
        RECT 239.500 188.200 239.900 189.900 ;
        RECT 239.000 187.900 239.900 188.200 ;
        RECT 240.600 187.900 241.000 189.900 ;
        RECT 241.400 188.000 241.800 189.900 ;
        RECT 243.000 188.000 243.400 189.900 ;
        RECT 241.400 187.900 243.400 188.000 ;
        RECT 233.400 187.100 233.800 187.200 ;
        RECT 234.200 187.100 235.200 187.200 ;
        RECT 230.900 186.900 231.400 187.100 ;
        RECT 226.100 185.400 228.200 185.700 ;
        RECT 229.400 185.400 229.800 186.200 ;
        RECT 224.600 184.900 225.800 185.200 ;
        RECT 224.300 184.500 224.700 184.600 ;
        RECT 223.600 184.200 224.700 184.500 ;
        RECT 225.500 184.400 225.800 184.900 ;
        RECT 225.500 184.000 226.200 184.400 ;
        RECT 222.300 183.700 222.700 183.800 ;
        RECT 223.700 183.700 224.100 183.800 ;
        RECT 220.600 183.100 221.000 183.500 ;
        RECT 222.300 183.400 224.100 183.700 ;
        RECT 223.400 183.100 223.700 183.400 ;
        RECT 225.400 183.100 225.800 183.500 ;
        RECT 220.600 182.800 221.600 183.100 ;
        RECT 221.200 181.100 221.600 182.800 ;
        RECT 223.400 181.100 223.800 183.100 ;
        RECT 225.500 181.100 226.100 183.100 ;
        RECT 227.800 181.100 228.200 185.400 ;
        RECT 230.100 184.900 230.400 186.800 ;
        RECT 230.700 186.500 231.400 186.900 ;
        RECT 233.400 186.800 235.200 187.100 ;
        RECT 235.700 187.100 237.800 187.400 ;
        RECT 235.700 186.900 236.200 187.100 ;
        RECT 231.100 185.500 231.400 186.500 ;
        RECT 231.800 185.800 232.200 186.600 ;
        RECT 232.600 186.100 233.000 186.600 ;
        RECT 233.400 186.100 233.800 186.200 ;
        RECT 232.600 185.800 233.800 186.100 ;
        RECT 231.100 185.200 233.000 185.500 ;
        RECT 234.200 185.400 234.600 186.200 ;
        RECT 230.100 184.600 230.900 184.900 ;
        RECT 230.500 182.200 230.900 184.600 ;
        RECT 232.700 183.500 233.000 185.200 ;
        RECT 234.900 184.900 235.200 186.800 ;
        RECT 235.500 186.500 236.200 186.900 ;
        RECT 238.200 186.800 238.600 187.600 ;
        RECT 235.900 185.500 236.200 186.500 ;
        RECT 236.600 185.800 237.000 186.600 ;
        RECT 237.400 185.800 237.800 186.600 ;
        RECT 238.200 186.200 238.500 186.800 ;
        RECT 238.200 185.800 238.600 186.200 ;
        RECT 239.000 186.100 239.400 187.900 ;
        RECT 240.700 187.200 241.000 187.900 ;
        RECT 241.500 187.700 243.300 187.900 ;
        RECT 243.800 187.700 244.200 189.900 ;
        RECT 245.900 189.200 246.500 189.900 ;
        RECT 245.900 188.900 246.600 189.200 ;
        RECT 248.200 188.900 248.600 189.900 ;
        RECT 250.400 189.200 250.800 189.900 ;
        RECT 250.400 188.900 251.400 189.200 ;
        RECT 246.200 188.500 246.600 188.900 ;
        RECT 248.300 188.600 248.600 188.900 ;
        RECT 248.300 188.300 249.700 188.600 ;
        RECT 249.300 188.200 249.700 188.300 ;
        RECT 250.200 188.200 250.600 188.600 ;
        RECT 251.000 188.500 251.400 188.900 ;
        RECT 245.300 187.700 245.700 187.800 ;
        RECT 243.800 187.400 245.700 187.700 ;
        RECT 242.600 187.200 243.000 187.400 ;
        RECT 240.600 186.800 241.900 187.200 ;
        RECT 242.600 186.900 243.400 187.200 ;
        RECT 243.000 186.800 243.400 186.900 ;
        RECT 239.000 185.800 240.900 186.100 ;
        RECT 235.900 185.200 237.800 185.500 ;
        RECT 234.900 184.600 235.700 184.900 ;
        RECT 230.200 181.800 230.900 182.200 ;
        RECT 230.500 181.100 230.900 181.800 ;
        RECT 232.600 181.500 233.000 183.500 ;
        RECT 235.300 181.100 235.700 184.600 ;
        RECT 237.500 183.500 237.800 185.200 ;
        RECT 237.400 181.500 237.800 183.500 ;
        RECT 239.000 181.100 239.400 185.800 ;
        RECT 240.600 185.200 240.900 185.800 ;
        RECT 241.600 185.200 241.900 186.800 ;
        RECT 242.200 186.100 242.600 186.600 ;
        RECT 243.000 186.100 243.400 186.200 ;
        RECT 242.200 185.800 243.400 186.100 ;
        RECT 243.800 185.700 244.200 187.400 ;
        RECT 247.300 187.100 247.700 187.200 ;
        RECT 250.200 187.100 250.500 188.200 ;
        RECT 252.600 187.500 253.000 189.900 ;
        RECT 254.200 187.600 254.600 189.900 ;
        RECT 255.800 187.600 256.200 189.900 ;
        RECT 257.400 187.600 257.800 189.900 ;
        RECT 259.000 187.600 259.400 189.900 ;
        RECT 260.900 189.200 261.300 189.900 ;
        RECT 260.900 188.800 261.800 189.200 ;
        RECT 260.900 188.200 261.300 188.800 ;
        RECT 260.900 187.900 261.800 188.200 ;
        RECT 254.200 187.200 255.100 187.600 ;
        RECT 255.800 187.200 256.900 187.600 ;
        RECT 257.400 187.200 258.500 187.600 ;
        RECT 259.000 187.200 260.200 187.600 ;
        RECT 251.800 187.100 252.600 187.200 ;
        RECT 247.100 186.800 252.600 187.100 ;
        RECT 253.400 186.900 253.800 187.200 ;
        RECT 254.700 186.900 255.100 187.200 ;
        RECT 256.500 186.900 256.900 187.200 ;
        RECT 258.100 186.900 258.500 187.200 ;
        RECT 246.200 186.400 246.600 186.500 ;
        RECT 244.700 186.100 246.600 186.400 ;
        RECT 244.700 186.000 245.100 186.100 ;
        RECT 245.500 185.700 245.900 185.800 ;
        RECT 243.800 185.400 245.900 185.700 ;
        RECT 239.800 184.400 240.200 185.200 ;
        RECT 240.600 185.100 241.000 185.200 ;
        RECT 240.600 184.800 241.300 185.100 ;
        RECT 241.600 184.800 242.600 185.200 ;
        RECT 241.000 184.200 241.300 184.800 ;
        RECT 241.000 183.800 241.400 184.200 ;
        RECT 241.700 181.100 242.100 184.800 ;
        RECT 243.800 181.100 244.200 185.400 ;
        RECT 247.100 185.200 247.400 186.800 ;
        RECT 250.700 186.700 251.100 186.800 ;
        RECT 253.400 186.500 254.300 186.900 ;
        RECT 254.700 186.500 256.000 186.900 ;
        RECT 256.500 186.500 257.700 186.900 ;
        RECT 258.100 186.500 259.400 186.900 ;
        RECT 251.500 186.200 251.900 186.300 ;
        RECT 249.400 185.900 251.900 186.200 ;
        RECT 249.400 185.800 249.800 185.900 ;
        RECT 254.700 185.800 255.100 186.500 ;
        RECT 256.500 185.800 256.900 186.500 ;
        RECT 258.100 185.800 258.500 186.500 ;
        RECT 259.800 185.800 260.200 187.200 ;
        RECT 250.200 185.500 253.000 185.600 ;
        RECT 250.100 185.400 253.000 185.500 ;
        RECT 246.200 184.900 247.400 185.200 ;
        RECT 248.100 185.300 253.000 185.400 ;
        RECT 248.100 185.100 250.500 185.300 ;
        RECT 246.200 184.400 246.500 184.900 ;
        RECT 245.800 184.000 246.500 184.400 ;
        RECT 247.300 184.500 247.700 184.600 ;
        RECT 248.100 184.500 248.400 185.100 ;
        RECT 247.300 184.200 248.400 184.500 ;
        RECT 248.700 184.500 251.400 184.800 ;
        RECT 248.700 184.400 249.100 184.500 ;
        RECT 251.000 184.400 251.400 184.500 ;
        RECT 247.900 183.700 248.300 183.800 ;
        RECT 249.300 183.700 249.700 183.800 ;
        RECT 246.200 183.100 246.600 183.500 ;
        RECT 247.900 183.400 249.700 183.700 ;
        RECT 248.300 183.100 248.600 183.400 ;
        RECT 251.000 183.100 251.400 183.500 ;
        RECT 245.900 181.100 246.500 183.100 ;
        RECT 248.200 181.100 248.600 183.100 ;
        RECT 250.400 182.800 251.400 183.100 ;
        RECT 250.400 181.100 250.800 182.800 ;
        RECT 252.600 181.100 253.000 185.300 ;
        RECT 254.200 185.400 255.100 185.800 ;
        RECT 255.800 185.400 256.900 185.800 ;
        RECT 257.400 185.400 258.500 185.800 ;
        RECT 259.000 185.400 260.200 185.800 ;
        RECT 254.200 181.100 254.600 185.400 ;
        RECT 255.800 181.100 256.200 185.400 ;
        RECT 257.400 181.100 257.800 185.400 ;
        RECT 259.000 181.100 259.400 185.400 ;
        RECT 260.600 184.400 261.000 185.200 ;
        RECT 261.400 181.100 261.800 187.900 ;
        RECT 262.200 187.100 262.600 187.600 ;
        RECT 263.800 187.100 264.200 187.200 ;
        RECT 262.200 186.800 264.200 187.100 ;
        RECT 0.600 175.600 1.000 179.900 ;
        RECT 2.700 177.900 3.300 179.900 ;
        RECT 5.000 177.900 5.400 179.900 ;
        RECT 7.200 178.200 7.600 179.900 ;
        RECT 7.200 177.900 8.200 178.200 ;
        RECT 3.000 177.500 3.400 177.900 ;
        RECT 5.100 177.600 5.400 177.900 ;
        RECT 4.700 177.300 6.500 177.600 ;
        RECT 7.800 177.500 8.200 177.900 ;
        RECT 4.700 177.200 5.100 177.300 ;
        RECT 6.100 177.200 6.500 177.300 ;
        RECT 2.600 176.600 3.300 177.000 ;
        RECT 3.000 176.100 3.300 176.600 ;
        RECT 4.100 176.500 5.200 176.800 ;
        RECT 4.100 176.400 4.500 176.500 ;
        RECT 3.000 175.800 4.200 176.100 ;
        RECT 0.600 175.300 2.700 175.600 ;
        RECT 0.600 173.600 1.000 175.300 ;
        RECT 2.300 175.200 2.700 175.300 ;
        RECT 1.500 174.900 1.900 175.000 ;
        RECT 1.500 174.600 3.400 174.900 ;
        RECT 3.000 174.500 3.400 174.600 ;
        RECT 3.900 174.200 4.200 175.800 ;
        RECT 4.900 175.900 5.200 176.500 ;
        RECT 5.500 176.500 5.900 176.600 ;
        RECT 7.800 176.500 8.200 176.600 ;
        RECT 5.500 176.200 8.200 176.500 ;
        RECT 4.900 175.700 7.300 175.900 ;
        RECT 9.400 175.700 9.800 179.900 ;
        RECT 12.100 179.200 12.500 179.900 ;
        RECT 11.800 178.800 12.500 179.200 ;
        RECT 12.100 176.400 12.500 178.800 ;
        RECT 14.200 177.500 14.600 179.500 ;
        RECT 4.900 175.600 9.800 175.700 ;
        RECT 11.700 176.100 12.500 176.400 ;
        RECT 6.900 175.500 9.800 175.600 ;
        RECT 7.000 175.400 9.800 175.500 ;
        RECT 6.200 175.100 6.600 175.200 ;
        RECT 6.200 174.800 8.700 175.100 ;
        RECT 11.000 174.800 11.400 175.600 ;
        RECT 7.000 174.700 7.400 174.800 ;
        RECT 8.300 174.700 8.700 174.800 ;
        RECT 7.500 174.200 7.900 174.300 ;
        RECT 11.700 174.200 12.000 176.100 ;
        RECT 14.300 175.800 14.600 177.500 ;
        RECT 12.700 175.500 14.600 175.800 ;
        RECT 15.000 177.500 15.400 179.500 ;
        RECT 15.000 175.800 15.300 177.500 ;
        RECT 17.100 176.400 17.500 179.900 ;
        RECT 21.700 176.400 22.100 179.900 ;
        RECT 23.800 177.500 24.200 179.500 ;
        RECT 17.100 176.100 17.900 176.400 ;
        RECT 15.000 175.500 16.900 175.800 ;
        RECT 12.700 174.500 13.000 175.500 ;
        RECT 3.900 173.900 9.400 174.200 ;
        RECT 4.100 173.800 4.500 173.900 ;
        RECT 0.600 173.300 2.500 173.600 ;
        RECT 0.600 171.100 1.000 173.300 ;
        RECT 2.100 173.200 2.500 173.300 ;
        RECT 7.000 172.800 7.300 173.900 ;
        RECT 8.600 173.800 9.400 173.900 ;
        RECT 11.000 173.800 12.000 174.200 ;
        RECT 12.300 174.100 13.000 174.500 ;
        RECT 13.400 174.400 13.800 175.200 ;
        RECT 14.200 174.400 14.600 175.200 ;
        RECT 15.000 174.400 15.400 175.200 ;
        RECT 15.800 174.400 16.200 175.200 ;
        RECT 16.600 174.500 16.900 175.500 ;
        RECT 11.700 173.500 12.000 173.800 ;
        RECT 12.500 173.900 13.000 174.100 ;
        RECT 16.600 174.100 17.300 174.500 ;
        RECT 17.600 174.200 17.900 176.100 ;
        RECT 21.300 176.100 22.100 176.400 ;
        RECT 18.200 175.100 18.600 175.600 ;
        RECT 19.000 175.100 19.400 175.200 ;
        RECT 20.600 175.100 21.000 175.600 ;
        RECT 18.200 174.800 19.400 175.100 ;
        RECT 19.800 174.800 21.000 175.100 ;
        RECT 17.600 174.100 18.600 174.200 ;
        RECT 19.800 174.100 20.100 174.800 ;
        RECT 21.300 174.200 21.600 176.100 ;
        RECT 23.900 175.800 24.200 177.500 ;
        RECT 26.500 176.400 26.900 179.900 ;
        RECT 28.600 177.500 29.000 179.500 ;
        RECT 22.300 175.500 24.200 175.800 ;
        RECT 26.100 176.100 26.900 176.400 ;
        RECT 26.100 175.800 26.600 176.100 ;
        RECT 28.700 175.800 29.000 177.500 ;
        RECT 31.300 178.200 31.700 179.900 ;
        RECT 31.300 177.800 32.200 178.200 ;
        RECT 31.300 176.400 31.700 177.800 ;
        RECT 33.400 177.500 33.800 179.500 ;
        RECT 22.300 174.500 22.600 175.500 ;
        RECT 16.600 173.900 17.100 174.100 ;
        RECT 12.500 173.600 14.600 173.900 ;
        RECT 6.100 172.700 6.500 172.800 ;
        RECT 3.000 172.100 3.400 172.500 ;
        RECT 5.100 172.400 6.500 172.700 ;
        RECT 7.000 172.400 7.400 172.800 ;
        RECT 5.100 172.100 5.400 172.400 ;
        RECT 7.800 172.100 8.200 172.500 ;
        RECT 2.700 171.800 3.400 172.100 ;
        RECT 2.700 171.100 3.300 171.800 ;
        RECT 5.000 171.100 5.400 172.100 ;
        RECT 7.200 171.800 8.200 172.100 ;
        RECT 7.200 171.100 7.600 171.800 ;
        RECT 9.400 171.100 9.800 173.500 ;
        RECT 11.700 173.300 12.100 173.500 ;
        RECT 11.700 173.000 12.500 173.300 ;
        RECT 12.100 171.500 12.500 173.000 ;
        RECT 14.300 172.500 14.600 173.600 ;
        RECT 14.200 171.500 14.600 172.500 ;
        RECT 15.000 173.600 17.100 173.900 ;
        RECT 17.600 173.800 20.100 174.100 ;
        RECT 20.600 173.800 21.600 174.200 ;
        RECT 21.900 174.100 22.600 174.500 ;
        RECT 23.000 174.400 23.400 175.200 ;
        RECT 23.800 174.400 24.200 175.200 ;
        RECT 25.400 174.800 25.800 175.600 ;
        RECT 26.100 174.200 26.400 175.800 ;
        RECT 27.100 175.500 29.000 175.800 ;
        RECT 30.900 176.100 31.700 176.400 ;
        RECT 27.100 174.500 27.400 175.500 ;
        RECT 15.000 172.500 15.300 173.600 ;
        RECT 17.600 173.500 17.900 173.800 ;
        RECT 17.500 173.300 17.900 173.500 ;
        RECT 17.100 173.000 17.900 173.300 ;
        RECT 21.300 173.500 21.600 173.800 ;
        RECT 22.100 173.900 22.600 174.100 ;
        RECT 22.100 173.600 24.200 173.900 ;
        RECT 25.400 173.800 26.400 174.200 ;
        RECT 26.700 174.100 27.400 174.500 ;
        RECT 27.800 174.400 28.200 175.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 29.400 175.100 29.800 175.200 ;
        RECT 28.600 174.800 29.800 175.100 ;
        RECT 30.200 174.800 30.600 175.600 ;
        RECT 28.600 174.400 29.000 174.800 ;
        RECT 30.900 174.200 31.200 176.100 ;
        RECT 33.500 175.800 33.800 177.500 ;
        RECT 34.200 175.800 34.600 176.600 ;
        RECT 31.900 175.500 33.800 175.800 ;
        RECT 31.900 174.500 32.200 175.500 ;
        RECT 21.300 173.300 21.700 173.500 ;
        RECT 21.300 173.200 22.100 173.300 ;
        RECT 21.300 173.000 22.600 173.200 ;
        RECT 15.000 171.500 15.400 172.500 ;
        RECT 17.100 171.500 17.500 173.000 ;
        RECT 21.700 172.800 22.600 173.000 ;
        RECT 21.700 171.500 22.100 172.800 ;
        RECT 23.900 172.500 24.200 173.600 ;
        RECT 26.100 173.500 26.400 173.800 ;
        RECT 26.900 173.900 27.400 174.100 ;
        RECT 26.900 173.600 29.000 173.900 ;
        RECT 30.200 173.800 31.200 174.200 ;
        RECT 31.500 174.100 32.200 174.500 ;
        RECT 32.600 174.400 33.000 175.200 ;
        RECT 33.400 174.400 33.800 175.200 ;
        RECT 26.100 173.300 26.500 173.500 ;
        RECT 26.100 173.000 26.900 173.300 ;
        RECT 23.800 171.500 24.200 172.500 ;
        RECT 26.500 171.500 26.900 173.000 ;
        RECT 28.700 172.500 29.000 173.600 ;
        RECT 30.900 173.500 31.200 173.800 ;
        RECT 31.700 173.900 32.200 174.100 ;
        RECT 31.700 173.600 33.800 173.900 ;
        RECT 30.900 173.300 31.300 173.500 ;
        RECT 30.900 173.000 31.700 173.300 ;
        RECT 28.600 171.500 29.000 172.500 ;
        RECT 31.300 171.500 31.700 173.000 ;
        RECT 33.500 172.500 33.800 173.600 ;
        RECT 35.000 173.100 35.400 179.900 ;
        RECT 36.600 176.200 37.000 179.900 ;
        RECT 38.200 179.600 40.200 179.900 ;
        RECT 38.200 176.200 38.600 179.600 ;
        RECT 36.600 175.900 38.600 176.200 ;
        RECT 39.000 175.900 39.400 179.300 ;
        RECT 39.800 175.900 40.200 179.600 ;
        RECT 40.600 176.200 41.000 179.900 ;
        RECT 42.200 179.600 44.200 179.900 ;
        RECT 42.200 176.200 42.600 179.600 ;
        RECT 40.600 175.900 42.600 176.200 ;
        RECT 43.000 175.900 43.400 179.300 ;
        RECT 43.800 175.900 44.200 179.600 ;
        RECT 45.400 176.400 45.800 179.900 ;
        RECT 45.300 175.900 45.800 176.400 ;
        RECT 47.000 176.200 47.400 179.900 ;
        RECT 46.100 175.900 47.400 176.200 ;
        RECT 48.100 176.300 48.500 179.900 ;
        RECT 52.100 177.200 52.500 179.900 ;
        RECT 54.200 177.500 54.600 179.500 ;
        RECT 52.100 176.800 53.000 177.200 ;
        RECT 52.100 176.400 52.500 176.800 ;
        RECT 48.100 175.900 49.000 176.300 ;
        RECT 51.700 176.100 52.500 176.400 ;
        RECT 39.000 175.600 39.300 175.900 ;
        RECT 43.000 175.600 43.300 175.900 ;
        RECT 37.000 175.200 37.400 175.400 ;
        RECT 38.300 175.300 39.300 175.600 ;
        RECT 38.300 175.200 38.600 175.300 ;
        RECT 35.800 175.100 36.200 175.200 ;
        RECT 36.600 175.100 37.400 175.200 ;
        RECT 35.800 174.900 37.400 175.100 ;
        RECT 35.800 174.800 37.000 174.900 ;
        RECT 38.200 174.800 38.600 175.200 ;
        RECT 39.800 174.800 40.200 175.600 ;
        RECT 41.000 175.200 41.400 175.400 ;
        RECT 42.300 175.300 43.300 175.600 ;
        RECT 42.300 175.200 42.600 175.300 ;
        RECT 40.600 174.900 41.400 175.200 ;
        RECT 40.600 174.800 41.000 174.900 ;
        RECT 42.200 174.800 42.600 175.200 ;
        RECT 43.800 174.800 44.200 175.600 ;
        RECT 35.800 174.100 36.200 174.200 ;
        RECT 36.600 174.100 37.000 174.200 ;
        RECT 35.800 173.800 37.000 174.100 ;
        RECT 37.400 173.800 37.800 174.600 ;
        RECT 35.800 173.400 36.200 173.800 ;
        RECT 38.300 173.100 38.600 174.800 ;
        RECT 38.900 174.400 39.300 174.800 ;
        RECT 39.000 174.200 39.300 174.400 ;
        RECT 39.000 174.100 39.400 174.200 ;
        RECT 39.800 174.100 40.200 174.200 ;
        RECT 39.000 173.800 40.200 174.100 ;
        RECT 41.400 173.800 41.800 174.600 ;
        RECT 42.300 173.100 42.600 174.800 ;
        RECT 42.900 174.400 43.300 174.800 ;
        RECT 43.000 174.200 43.300 174.400 ;
        RECT 45.300 174.200 45.600 175.900 ;
        RECT 46.100 174.900 46.400 175.900 ;
        RECT 45.900 174.500 46.400 174.900 ;
        RECT 43.000 173.800 43.400 174.200 ;
        RECT 45.300 173.800 45.800 174.200 ;
        RECT 45.300 173.100 45.600 173.800 ;
        RECT 46.100 173.700 46.400 174.500 ;
        RECT 46.900 174.800 47.400 175.200 ;
        RECT 47.800 174.800 48.200 175.600 ;
        RECT 46.900 174.400 47.300 174.800 ;
        RECT 48.600 174.200 48.900 175.900 ;
        RECT 49.400 175.100 49.800 175.200 ;
        RECT 51.000 175.100 51.400 175.600 ;
        RECT 49.400 174.800 51.400 175.100 ;
        RECT 51.700 174.200 52.000 176.100 ;
        RECT 54.300 175.800 54.600 177.500 ;
        RECT 52.700 175.500 54.600 175.800 ;
        RECT 56.600 177.500 57.000 179.500 ;
        RECT 56.600 175.800 56.900 177.500 ;
        RECT 58.700 176.400 59.100 179.900 ;
        RECT 63.300 176.400 63.700 179.900 ;
        RECT 65.400 177.500 65.800 179.500 ;
        RECT 58.700 176.100 59.500 176.400 ;
        RECT 56.600 175.500 58.500 175.800 ;
        RECT 52.700 174.500 53.000 175.500 ;
        RECT 48.600 173.800 49.000 174.200 ;
        RECT 51.000 173.800 52.000 174.200 ;
        RECT 52.300 174.100 53.000 174.500 ;
        RECT 53.400 174.400 53.800 175.200 ;
        RECT 54.200 174.400 54.600 175.200 ;
        RECT 55.800 175.100 56.200 175.200 ;
        RECT 56.600 175.100 57.000 175.200 ;
        RECT 55.800 174.800 57.000 175.100 ;
        RECT 56.600 174.400 57.000 174.800 ;
        RECT 57.400 174.400 57.800 175.200 ;
        RECT 58.200 174.500 58.500 175.500 ;
        RECT 46.100 173.400 47.400 173.700 ;
        RECT 33.400 171.500 33.800 172.500 ;
        RECT 34.500 172.800 35.400 173.100 ;
        RECT 34.500 172.200 34.900 172.800 ;
        RECT 38.100 172.200 38.900 173.100 ;
        RECT 42.100 172.200 42.900 173.100 ;
        RECT 45.300 172.800 45.800 173.100 ;
        RECT 34.500 171.800 35.400 172.200 ;
        RECT 38.100 171.800 39.400 172.200 ;
        RECT 42.100 171.800 43.400 172.200 ;
        RECT 34.500 171.100 34.900 171.800 ;
        RECT 38.100 171.100 38.900 171.800 ;
        RECT 42.100 171.100 42.900 171.800 ;
        RECT 45.400 171.100 45.800 172.800 ;
        RECT 47.000 171.100 47.400 173.400 ;
        RECT 48.600 172.200 48.900 173.800 ;
        RECT 51.700 173.500 52.000 173.800 ;
        RECT 52.500 173.900 53.000 174.100 ;
        RECT 58.200 174.100 58.900 174.500 ;
        RECT 59.200 174.200 59.500 176.100 ;
        RECT 62.900 176.100 63.700 176.400 ;
        RECT 59.800 175.100 60.200 175.600 ;
        RECT 59.800 174.800 60.900 175.100 ;
        RECT 62.200 174.800 62.600 175.600 ;
        RECT 58.200 173.900 58.700 174.100 ;
        RECT 52.500 173.600 54.600 173.900 ;
        RECT 51.700 173.300 52.100 173.500 ;
        RECT 49.400 172.400 49.800 173.200 ;
        RECT 51.700 173.000 52.500 173.300 ;
        RECT 48.600 171.100 49.000 172.200 ;
        RECT 52.100 171.500 52.500 173.000 ;
        RECT 54.300 172.500 54.600 173.600 ;
        RECT 54.200 171.500 54.600 172.500 ;
        RECT 56.600 173.600 58.700 173.900 ;
        RECT 59.200 173.800 60.200 174.200 ;
        RECT 60.600 174.100 60.900 174.800 ;
        RECT 62.900 174.200 63.200 176.100 ;
        RECT 65.500 175.800 65.800 177.500 ;
        RECT 63.900 175.500 65.800 175.800 ;
        RECT 63.900 174.500 64.200 175.500 ;
        RECT 62.200 174.100 63.200 174.200 ;
        RECT 63.500 174.100 64.200 174.500 ;
        RECT 64.600 174.400 65.000 175.200 ;
        RECT 65.400 174.400 65.800 175.200 ;
        RECT 67.000 175.100 67.400 179.900 ;
        RECT 69.000 176.800 69.400 177.200 ;
        RECT 67.800 175.800 68.200 176.600 ;
        RECT 69.000 176.200 69.300 176.800 ;
        RECT 69.700 176.200 70.100 179.900 ;
        RECT 68.600 175.900 69.300 176.200 ;
        RECT 69.600 175.900 70.100 176.200 ;
        RECT 68.600 175.800 69.000 175.900 ;
        RECT 68.600 175.100 68.900 175.800 ;
        RECT 67.000 174.800 68.900 175.100 ;
        RECT 60.600 173.800 63.200 174.100 ;
        RECT 56.600 172.500 56.900 173.600 ;
        RECT 59.200 173.500 59.500 173.800 ;
        RECT 59.100 173.300 59.500 173.500 ;
        RECT 58.700 173.000 59.500 173.300 ;
        RECT 62.900 173.500 63.200 173.800 ;
        RECT 63.700 173.900 64.200 174.100 ;
        RECT 63.700 173.600 65.800 173.900 ;
        RECT 62.900 173.300 63.300 173.500 ;
        RECT 62.900 173.000 63.700 173.300 ;
        RECT 56.600 171.500 57.000 172.500 ;
        RECT 58.700 172.200 59.100 173.000 ;
        RECT 58.700 171.800 59.400 172.200 ;
        RECT 58.700 171.500 59.100 171.800 ;
        RECT 63.300 171.500 63.700 173.000 ;
        RECT 65.500 172.500 65.800 173.600 ;
        RECT 66.200 173.400 66.600 174.200 ;
        RECT 67.000 173.100 67.400 174.800 ;
        RECT 69.600 174.200 69.900 175.900 ;
        RECT 71.800 175.600 72.200 179.900 ;
        RECT 73.900 177.900 74.500 179.900 ;
        RECT 76.200 177.900 76.600 179.900 ;
        RECT 78.400 178.200 78.800 179.900 ;
        RECT 78.400 177.900 79.400 178.200 ;
        RECT 74.200 177.500 74.600 177.900 ;
        RECT 76.300 177.600 76.600 177.900 ;
        RECT 75.900 177.300 77.700 177.600 ;
        RECT 79.000 177.500 79.400 177.900 ;
        RECT 75.900 177.200 76.300 177.300 ;
        RECT 77.300 177.200 77.700 177.300 ;
        RECT 73.800 176.600 74.500 177.000 ;
        RECT 74.200 176.100 74.500 176.600 ;
        RECT 75.300 176.500 76.400 176.800 ;
        RECT 75.300 176.400 75.700 176.500 ;
        RECT 74.200 175.800 75.400 176.100 ;
        RECT 71.800 175.300 73.900 175.600 ;
        RECT 70.200 174.400 70.600 175.200 ;
        RECT 68.600 173.800 69.900 174.200 ;
        RECT 71.000 174.100 71.400 174.200 ;
        RECT 70.600 173.800 71.400 174.100 ;
        RECT 68.700 173.100 69.000 173.800 ;
        RECT 70.600 173.600 71.000 173.800 ;
        RECT 71.800 173.600 72.200 175.300 ;
        RECT 73.500 175.200 73.900 175.300 ;
        RECT 72.700 174.900 73.100 175.000 ;
        RECT 72.700 174.600 74.600 174.900 ;
        RECT 74.200 174.500 74.600 174.600 ;
        RECT 75.100 174.200 75.400 175.800 ;
        RECT 76.100 175.900 76.400 176.500 ;
        RECT 76.700 176.500 77.100 176.600 ;
        RECT 79.000 176.500 79.400 176.600 ;
        RECT 76.700 176.200 79.400 176.500 ;
        RECT 76.100 175.700 78.500 175.900 ;
        RECT 80.600 175.700 81.000 179.900 ;
        RECT 81.400 179.600 83.400 179.900 ;
        RECT 81.400 175.900 81.800 179.600 ;
        RECT 82.200 175.900 82.600 179.300 ;
        RECT 83.000 176.200 83.400 179.600 ;
        RECT 84.600 176.200 85.000 179.900 ;
        RECT 83.000 175.900 85.000 176.200 ;
        RECT 76.100 175.600 81.000 175.700 ;
        RECT 82.300 175.600 82.600 175.900 ;
        RECT 85.400 175.600 85.800 179.900 ;
        RECT 87.500 177.900 88.100 179.900 ;
        RECT 89.800 177.900 90.200 179.900 ;
        RECT 92.000 178.200 92.400 179.900 ;
        RECT 92.000 177.900 93.000 178.200 ;
        RECT 87.800 177.500 88.200 177.900 ;
        RECT 89.900 177.600 90.200 177.900 ;
        RECT 89.500 177.300 91.300 177.600 ;
        RECT 92.600 177.500 93.000 177.900 ;
        RECT 89.500 177.200 89.900 177.300 ;
        RECT 90.900 177.200 91.300 177.300 ;
        RECT 87.400 176.600 88.100 177.000 ;
        RECT 87.800 176.100 88.100 176.600 ;
        RECT 88.900 176.500 90.000 176.800 ;
        RECT 88.900 176.400 89.300 176.500 ;
        RECT 87.800 175.800 89.000 176.100 ;
        RECT 78.100 175.500 81.000 175.600 ;
        RECT 78.200 175.400 81.000 175.500 ;
        RECT 76.600 175.100 77.000 175.200 ;
        RECT 77.400 175.100 77.800 175.200 ;
        RECT 76.600 174.800 79.900 175.100 ;
        RECT 81.400 174.800 81.800 175.600 ;
        RECT 82.300 175.300 83.300 175.600 ;
        RECT 83.000 175.200 83.300 175.300 ;
        RECT 84.200 175.200 84.600 175.400 ;
        RECT 85.400 175.300 87.500 175.600 ;
        RECT 83.000 174.800 83.400 175.200 ;
        RECT 84.200 174.900 85.000 175.200 ;
        RECT 84.600 174.800 85.000 174.900 ;
        RECT 79.500 174.700 79.900 174.800 ;
        RECT 82.300 174.400 82.700 174.800 ;
        RECT 78.700 174.200 79.100 174.300 ;
        RECT 82.300 174.200 82.600 174.400 ;
        RECT 75.100 173.900 80.600 174.200 ;
        RECT 75.300 173.800 75.700 173.900 ;
        RECT 71.800 173.300 73.700 173.600 ;
        RECT 69.500 173.100 71.300 173.300 ;
        RECT 67.000 172.800 67.900 173.100 ;
        RECT 65.400 171.500 65.800 172.500 ;
        RECT 67.500 171.100 67.900 172.800 ;
        RECT 68.600 171.100 69.000 173.100 ;
        RECT 69.400 173.000 71.400 173.100 ;
        RECT 69.400 171.100 69.800 173.000 ;
        RECT 71.000 171.100 71.400 173.000 ;
        RECT 71.800 171.100 72.200 173.300 ;
        RECT 73.300 173.200 73.700 173.300 ;
        RECT 78.200 172.800 78.500 173.900 ;
        RECT 79.800 173.800 80.600 173.900 ;
        RECT 82.200 173.800 82.600 174.200 ;
        RECT 77.300 172.700 77.700 172.800 ;
        RECT 74.200 172.100 74.600 172.500 ;
        RECT 76.300 172.400 77.700 172.700 ;
        RECT 78.200 172.400 78.600 172.800 ;
        RECT 76.300 172.100 76.600 172.400 ;
        RECT 79.000 172.100 79.400 172.500 ;
        RECT 73.900 171.800 74.600 172.100 ;
        RECT 73.900 171.100 74.500 171.800 ;
        RECT 76.200 171.100 76.600 172.100 ;
        RECT 78.400 171.800 79.400 172.100 ;
        RECT 78.400 171.100 78.800 171.800 ;
        RECT 80.600 171.100 81.000 173.500 ;
        RECT 83.000 173.100 83.300 174.800 ;
        RECT 83.800 174.100 84.200 174.600 ;
        RECT 84.600 174.100 85.000 174.200 ;
        RECT 83.800 173.800 85.000 174.100 ;
        RECT 85.400 173.600 85.800 175.300 ;
        RECT 87.100 175.200 87.500 175.300 ;
        RECT 88.700 175.200 89.000 175.800 ;
        RECT 89.700 175.900 90.000 176.500 ;
        RECT 90.300 176.500 90.700 176.600 ;
        RECT 92.600 176.500 93.000 176.600 ;
        RECT 90.300 176.200 93.000 176.500 ;
        RECT 89.700 175.700 92.100 175.900 ;
        RECT 94.200 175.700 94.600 179.900 ;
        RECT 95.000 179.600 97.000 179.900 ;
        RECT 95.000 175.900 95.400 179.600 ;
        RECT 95.800 175.900 96.200 179.300 ;
        RECT 96.600 176.200 97.000 179.600 ;
        RECT 98.200 176.200 98.600 179.900 ;
        RECT 100.900 176.400 101.300 179.900 ;
        RECT 103.000 177.500 103.400 179.500 ;
        RECT 96.600 175.900 98.600 176.200 ;
        RECT 100.500 176.100 101.300 176.400 ;
        RECT 89.700 175.600 94.600 175.700 ;
        RECT 95.900 175.600 96.200 175.900 ;
        RECT 91.700 175.500 94.600 175.600 ;
        RECT 91.800 175.400 94.600 175.500 ;
        RECT 86.300 174.900 86.700 175.000 ;
        RECT 86.300 174.600 88.200 174.900 ;
        RECT 88.600 174.800 89.000 175.200 ;
        RECT 91.000 175.100 91.400 175.200 ;
        RECT 91.000 174.800 93.500 175.100 ;
        RECT 95.000 174.800 95.400 175.600 ;
        RECT 95.900 175.300 96.900 175.600 ;
        RECT 96.600 175.200 96.900 175.300 ;
        RECT 97.800 175.200 98.200 175.400 ;
        RECT 96.600 174.800 97.000 175.200 ;
        RECT 97.800 174.900 98.600 175.200 ;
        RECT 98.200 174.800 98.600 174.900 ;
        RECT 99.800 174.800 100.200 175.600 ;
        RECT 87.800 174.500 88.200 174.600 ;
        RECT 88.700 174.200 89.000 174.800 ;
        RECT 91.800 174.700 92.200 174.800 ;
        RECT 93.100 174.700 93.500 174.800 ;
        RECT 95.900 174.400 96.300 174.800 ;
        RECT 92.300 174.200 92.700 174.300 ;
        RECT 95.900 174.200 96.200 174.400 ;
        RECT 88.700 173.900 94.200 174.200 ;
        RECT 88.900 173.800 89.300 173.900 ;
        RECT 85.400 173.300 87.300 173.600 ;
        RECT 82.700 171.100 83.500 173.100 ;
        RECT 85.400 171.100 85.800 173.300 ;
        RECT 86.900 173.200 87.300 173.300 ;
        RECT 91.800 172.800 92.100 173.900 ;
        RECT 93.400 173.800 94.200 173.900 ;
        RECT 95.800 173.800 96.200 174.200 ;
        RECT 90.900 172.700 91.300 172.800 ;
        RECT 87.800 172.100 88.200 172.500 ;
        RECT 89.900 172.400 91.300 172.700 ;
        RECT 91.800 172.400 92.200 172.800 ;
        RECT 89.900 172.100 90.200 172.400 ;
        RECT 92.600 172.100 93.000 172.500 ;
        RECT 87.500 171.800 88.200 172.100 ;
        RECT 87.500 171.100 88.100 171.800 ;
        RECT 89.800 171.100 90.200 172.100 ;
        RECT 92.000 171.800 93.000 172.100 ;
        RECT 92.000 171.100 92.400 171.800 ;
        RECT 94.200 171.100 94.600 173.500 ;
        RECT 96.600 173.100 96.900 174.800 ;
        RECT 97.400 173.800 97.800 174.600 ;
        RECT 98.200 174.100 98.500 174.800 ;
        RECT 100.500 174.200 100.800 176.100 ;
        RECT 103.100 175.800 103.400 177.500 ;
        RECT 101.500 175.500 103.400 175.800 ;
        RECT 101.500 174.500 101.800 175.500 ;
        RECT 99.800 174.100 100.800 174.200 ;
        RECT 101.100 174.100 101.800 174.500 ;
        RECT 102.200 174.400 102.600 175.200 ;
        RECT 103.000 174.400 103.400 175.200 ;
        RECT 98.200 173.800 100.800 174.100 ;
        RECT 100.500 173.500 100.800 173.800 ;
        RECT 101.300 173.900 101.800 174.100 ;
        RECT 101.300 173.600 103.400 173.900 ;
        RECT 100.500 173.300 100.900 173.500 ;
        RECT 96.300 171.100 97.100 173.100 ;
        RECT 100.500 173.000 101.300 173.300 ;
        RECT 100.900 171.500 101.300 173.000 ;
        RECT 103.100 172.500 103.400 173.600 ;
        RECT 103.800 173.400 104.200 174.200 ;
        RECT 104.600 173.100 105.000 179.900 ;
        RECT 107.800 179.600 109.800 179.900 ;
        RECT 105.400 176.100 105.800 176.600 ;
        RECT 106.200 176.100 106.600 176.200 ;
        RECT 105.400 175.800 106.600 176.100 ;
        RECT 107.800 175.900 108.200 179.600 ;
        RECT 108.600 175.800 109.000 179.300 ;
        RECT 109.400 176.200 109.800 179.600 ;
        RECT 111.000 176.200 111.400 179.900 ;
        RECT 109.400 175.900 111.400 176.200 ;
        RECT 108.700 175.600 109.000 175.800 ;
        RECT 107.800 174.800 108.200 175.600 ;
        RECT 108.700 175.300 109.700 175.600 ;
        RECT 109.400 175.200 109.700 175.300 ;
        RECT 110.600 175.200 111.000 175.400 ;
        RECT 109.400 174.800 109.800 175.200 ;
        RECT 110.600 174.900 111.400 175.200 ;
        RECT 111.000 174.800 111.400 174.900 ;
        RECT 108.700 174.400 109.100 174.800 ;
        RECT 108.700 174.200 109.000 174.400 ;
        RECT 105.400 174.100 105.800 174.200 ;
        RECT 108.600 174.100 109.000 174.200 ;
        RECT 105.400 173.800 109.000 174.100 ;
        RECT 109.400 173.100 109.700 174.800 ;
        RECT 110.200 173.800 110.600 174.600 ;
        RECT 111.800 173.400 112.200 174.200 ;
        RECT 112.600 173.100 113.000 179.900 ;
        RECT 114.200 179.600 116.200 179.900 ;
        RECT 113.400 175.800 113.800 176.600 ;
        RECT 114.200 175.900 114.600 179.600 ;
        RECT 115.000 175.800 115.400 179.300 ;
        RECT 115.800 176.200 116.200 179.600 ;
        RECT 117.400 176.200 117.800 179.900 ;
        RECT 115.800 175.900 117.800 176.200 ;
        RECT 115.100 175.600 115.400 175.800 ;
        RECT 118.200 175.600 118.600 179.900 ;
        RECT 120.300 177.900 120.900 179.900 ;
        RECT 122.600 177.900 123.000 179.900 ;
        RECT 124.800 178.200 125.200 179.900 ;
        RECT 124.800 177.900 125.800 178.200 ;
        RECT 120.600 177.500 121.000 177.900 ;
        RECT 122.700 177.600 123.000 177.900 ;
        RECT 122.300 177.300 124.100 177.600 ;
        RECT 125.400 177.500 125.800 177.900 ;
        RECT 122.300 177.200 122.700 177.300 ;
        RECT 123.700 177.200 124.100 177.300 ;
        RECT 120.200 176.600 120.900 177.000 ;
        RECT 120.600 176.100 120.900 176.600 ;
        RECT 121.700 176.500 122.800 176.800 ;
        RECT 121.700 176.400 122.100 176.500 ;
        RECT 120.600 175.800 121.800 176.100 ;
        RECT 113.400 175.100 113.800 175.200 ;
        RECT 114.200 175.100 114.600 175.600 ;
        RECT 115.100 175.300 116.100 175.600 ;
        RECT 113.400 174.800 114.600 175.100 ;
        RECT 115.800 175.200 116.100 175.300 ;
        RECT 117.000 175.200 117.400 175.400 ;
        RECT 118.200 175.300 120.300 175.600 ;
        RECT 115.800 174.800 116.200 175.200 ;
        RECT 117.000 174.900 117.800 175.200 ;
        RECT 117.400 174.800 117.800 174.900 ;
        RECT 115.100 174.400 115.500 174.800 ;
        RECT 115.100 174.200 115.400 174.400 ;
        RECT 114.200 174.100 114.600 174.200 ;
        RECT 115.000 174.100 115.400 174.200 ;
        RECT 114.200 173.800 115.400 174.100 ;
        RECT 115.800 173.100 116.100 174.800 ;
        RECT 116.600 173.800 117.000 174.600 ;
        RECT 118.200 173.600 118.600 175.300 ;
        RECT 119.900 175.200 120.300 175.300 ;
        RECT 119.100 174.900 119.500 175.000 ;
        RECT 119.100 174.600 121.000 174.900 ;
        RECT 120.600 174.500 121.000 174.600 ;
        RECT 121.500 174.200 121.800 175.800 ;
        RECT 122.500 175.900 122.800 176.500 ;
        RECT 123.100 176.500 123.500 176.600 ;
        RECT 125.400 176.500 125.800 176.600 ;
        RECT 123.100 176.200 125.800 176.500 ;
        RECT 122.500 175.700 124.900 175.900 ;
        RECT 127.000 175.700 127.400 179.900 ;
        RECT 129.100 176.300 129.500 179.900 ;
        RECT 128.600 175.900 129.500 176.300 ;
        RECT 130.200 175.900 130.600 179.900 ;
        RECT 131.000 176.200 131.400 179.900 ;
        RECT 132.600 176.200 133.000 179.900 ;
        RECT 131.000 175.900 133.000 176.200 ;
        RECT 122.500 175.600 127.400 175.700 ;
        RECT 124.500 175.500 127.400 175.600 ;
        RECT 124.600 175.400 127.400 175.500 ;
        RECT 123.800 175.100 124.200 175.200 ;
        RECT 123.800 174.800 126.300 175.100 ;
        RECT 124.600 174.700 125.000 174.800 ;
        RECT 125.900 174.700 126.300 174.800 ;
        RECT 125.100 174.200 125.500 174.300 ;
        RECT 128.700 174.200 129.000 175.900 ;
        RECT 129.400 174.800 129.800 175.600 ;
        RECT 130.300 175.200 130.600 175.900 ;
        RECT 133.400 175.700 133.800 179.900 ;
        RECT 135.600 178.200 136.000 179.900 ;
        RECT 135.000 177.900 136.000 178.200 ;
        RECT 137.800 177.900 138.200 179.900 ;
        RECT 139.900 177.900 140.500 179.900 ;
        RECT 135.000 177.500 135.400 177.900 ;
        RECT 137.800 177.600 138.100 177.900 ;
        RECT 136.700 177.300 138.500 177.600 ;
        RECT 139.800 177.500 140.200 177.900 ;
        RECT 136.700 177.200 137.100 177.300 ;
        RECT 138.100 177.200 138.500 177.300 ;
        RECT 135.000 176.500 135.400 176.600 ;
        RECT 137.300 176.500 137.700 176.600 ;
        RECT 135.000 176.200 137.700 176.500 ;
        RECT 138.000 176.500 139.100 176.800 ;
        RECT 138.000 175.900 138.300 176.500 ;
        RECT 138.700 176.400 139.100 176.500 ;
        RECT 139.900 176.600 140.600 177.000 ;
        RECT 139.900 176.100 140.200 176.600 ;
        RECT 135.900 175.700 138.300 175.900 ;
        RECT 133.400 175.600 138.300 175.700 ;
        RECT 139.000 175.800 140.200 176.100 ;
        RECT 133.400 175.500 136.300 175.600 ;
        RECT 133.400 175.400 136.200 175.500 ;
        RECT 132.200 175.200 132.600 175.400 ;
        RECT 130.200 174.900 131.400 175.200 ;
        RECT 132.200 174.900 133.000 175.200 ;
        RECT 136.600 175.100 137.000 175.200 ;
        RECT 130.200 174.800 130.600 174.900 ;
        RECT 121.500 173.900 127.000 174.200 ;
        RECT 121.700 173.800 122.100 173.900 ;
        RECT 118.200 173.300 120.100 173.600 ;
        RECT 104.600 172.800 105.500 173.100 ;
        RECT 103.000 171.500 103.400 172.500 ;
        RECT 105.100 172.200 105.500 172.800 ;
        RECT 104.600 171.800 105.500 172.200 ;
        RECT 105.100 171.100 105.500 171.800 ;
        RECT 109.100 171.100 109.900 173.100 ;
        RECT 112.600 172.800 113.500 173.100 ;
        RECT 113.100 172.200 113.500 172.800 ;
        RECT 113.100 171.800 113.800 172.200 ;
        RECT 113.100 171.100 113.500 171.800 ;
        RECT 115.500 171.100 116.300 173.100 ;
        RECT 118.200 171.100 118.600 173.300 ;
        RECT 119.700 173.200 120.100 173.300 ;
        RECT 124.600 172.800 124.900 173.900 ;
        RECT 126.200 173.800 127.000 173.900 ;
        RECT 128.600 173.800 129.000 174.200 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 131.100 174.100 131.400 174.900 ;
        RECT 132.600 174.800 133.000 174.900 ;
        RECT 134.500 174.800 137.000 175.100 ;
        RECT 134.500 174.700 134.900 174.800 ;
        RECT 130.200 173.800 131.400 174.100 ;
        RECT 131.800 174.100 132.200 174.600 ;
        RECT 135.300 174.200 135.700 174.300 ;
        RECT 139.000 174.200 139.300 175.800 ;
        RECT 142.200 175.600 142.600 179.900 ;
        RECT 140.500 175.300 142.600 175.600 ;
        RECT 140.500 175.200 140.900 175.300 ;
        RECT 141.300 174.900 141.700 175.000 ;
        RECT 139.800 174.600 141.700 174.900 ;
        RECT 139.800 174.500 140.200 174.600 ;
        RECT 132.600 174.100 133.000 174.200 ;
        RECT 131.800 173.800 133.000 174.100 ;
        RECT 133.800 173.900 139.300 174.200 ;
        RECT 133.800 173.800 134.600 173.900 ;
        RECT 123.700 172.700 124.100 172.800 ;
        RECT 120.600 172.100 121.000 172.500 ;
        RECT 122.700 172.400 124.100 172.700 ;
        RECT 124.600 172.400 125.000 172.800 ;
        RECT 122.700 172.100 123.000 172.400 ;
        RECT 125.400 172.100 125.800 172.500 ;
        RECT 120.300 171.800 121.000 172.100 ;
        RECT 120.300 171.100 120.900 171.800 ;
        RECT 122.600 171.100 123.000 172.100 ;
        RECT 124.800 171.800 125.800 172.100 ;
        RECT 124.800 171.100 125.200 171.800 ;
        RECT 127.000 171.100 127.400 173.500 ;
        RECT 127.800 172.400 128.200 173.200 ;
        RECT 128.700 173.100 129.000 173.800 ;
        RECT 130.200 173.100 130.600 173.200 ;
        RECT 131.100 173.100 131.400 173.800 ;
        RECT 128.600 172.800 130.600 173.100 ;
        RECT 128.700 172.100 129.000 172.800 ;
        RECT 130.300 172.400 130.700 172.800 ;
        RECT 128.600 171.100 129.000 172.100 ;
        RECT 131.000 171.100 131.400 173.100 ;
        RECT 133.400 171.100 133.800 173.500 ;
        RECT 135.900 172.800 136.200 173.900 ;
        RECT 138.700 173.800 139.100 173.900 ;
        RECT 142.200 173.600 142.600 175.300 ;
        RECT 140.600 173.300 142.600 173.600 ;
        RECT 140.600 173.200 141.100 173.300 ;
        RECT 139.000 173.100 139.400 173.200 ;
        RECT 140.600 173.100 141.000 173.200 ;
        RECT 139.000 172.800 141.000 173.100 ;
        RECT 142.200 173.100 142.600 173.300 ;
        RECT 143.800 175.100 144.200 179.900 ;
        RECT 146.500 176.400 146.900 179.900 ;
        RECT 148.600 177.500 149.000 179.500 ;
        RECT 146.100 176.100 146.900 176.400 ;
        RECT 145.400 175.100 145.800 175.600 ;
        RECT 143.800 174.800 145.800 175.100 ;
        RECT 143.000 173.100 143.400 173.200 ;
        RECT 142.200 172.800 143.400 173.100 ;
        RECT 135.000 172.100 135.400 172.500 ;
        RECT 135.800 172.400 136.200 172.800 ;
        RECT 136.700 172.700 137.100 172.800 ;
        RECT 136.700 172.400 138.100 172.700 ;
        RECT 137.800 172.100 138.100 172.400 ;
        RECT 139.800 172.100 140.200 172.500 ;
        RECT 135.000 171.800 136.000 172.100 ;
        RECT 135.600 171.100 136.000 171.800 ;
        RECT 137.800 171.100 138.200 172.100 ;
        RECT 139.800 171.800 140.500 172.100 ;
        RECT 139.900 171.100 140.500 171.800 ;
        RECT 142.200 171.100 142.600 172.800 ;
        RECT 143.000 172.400 143.400 172.800 ;
        RECT 143.800 171.100 144.200 174.800 ;
        RECT 146.100 174.200 146.400 176.100 ;
        RECT 148.700 175.800 149.000 177.500 ;
        RECT 149.400 176.200 149.800 179.900 ;
        RECT 151.000 176.200 151.400 179.900 ;
        RECT 149.400 175.900 151.400 176.200 ;
        RECT 151.800 175.900 152.200 179.900 ;
        RECT 147.100 175.500 149.000 175.800 ;
        RECT 147.100 174.500 147.400 175.500 ;
        RECT 149.800 175.200 150.200 175.400 ;
        RECT 151.800 175.200 152.100 175.900 ;
        RECT 152.600 175.800 153.000 177.200 ;
        RECT 144.600 174.100 145.000 174.200 ;
        RECT 145.400 174.100 146.400 174.200 ;
        RECT 146.700 174.100 147.400 174.500 ;
        RECT 147.800 174.400 148.200 175.200 ;
        RECT 148.600 174.400 149.000 175.200 ;
        RECT 149.400 174.900 150.200 175.200 ;
        RECT 151.000 174.900 152.200 175.200 ;
        RECT 153.400 175.100 153.800 179.900 ;
        RECT 156.600 175.700 157.000 179.900 ;
        RECT 158.800 178.200 159.200 179.900 ;
        RECT 158.200 177.900 159.200 178.200 ;
        RECT 161.000 177.900 161.400 179.900 ;
        RECT 163.100 177.900 163.700 179.900 ;
        RECT 158.200 177.500 158.600 177.900 ;
        RECT 161.000 177.600 161.300 177.900 ;
        RECT 159.900 177.300 161.700 177.600 ;
        RECT 163.000 177.500 163.400 177.900 ;
        RECT 159.900 177.200 160.300 177.300 ;
        RECT 161.300 177.200 161.700 177.300 ;
        RECT 158.200 176.500 158.600 176.600 ;
        RECT 160.500 176.500 160.900 176.600 ;
        RECT 158.200 176.200 160.900 176.500 ;
        RECT 161.200 176.500 162.300 176.800 ;
        RECT 161.200 175.900 161.500 176.500 ;
        RECT 161.900 176.400 162.300 176.500 ;
        RECT 163.100 176.600 163.800 177.000 ;
        RECT 163.100 176.100 163.400 176.600 ;
        RECT 159.100 175.700 161.500 175.900 ;
        RECT 156.600 175.600 161.500 175.700 ;
        RECT 162.200 175.800 163.400 176.100 ;
        RECT 156.600 175.500 159.500 175.600 ;
        RECT 156.600 175.400 159.400 175.500 ;
        RECT 159.800 175.100 160.200 175.200 ;
        RECT 149.400 174.800 149.800 174.900 ;
        RECT 144.600 173.800 146.400 174.100 ;
        RECT 146.100 173.500 146.400 173.800 ;
        RECT 146.900 173.900 147.400 174.100 ;
        RECT 146.900 173.600 149.000 173.900 ;
        RECT 150.200 173.800 150.600 174.600 ;
        RECT 146.100 173.300 146.500 173.500 ;
        RECT 146.100 173.000 146.900 173.300 ;
        RECT 146.500 171.500 146.900 173.000 ;
        RECT 148.700 172.500 149.000 173.600 ;
        RECT 148.600 171.500 149.000 172.500 ;
        RECT 151.000 173.100 151.300 174.900 ;
        RECT 151.800 174.800 152.200 174.900 ;
        RECT 152.600 174.800 153.800 175.100 ;
        RECT 152.600 174.200 152.900 174.800 ;
        RECT 152.600 173.800 153.000 174.200 ;
        RECT 151.000 171.100 151.400 173.100 ;
        RECT 151.800 172.800 152.200 173.200 ;
        RECT 153.400 173.100 153.800 174.800 ;
        RECT 157.700 174.800 160.200 175.100 ;
        RECT 157.700 174.700 158.100 174.800 ;
        RECT 158.500 174.200 158.900 174.300 ;
        RECT 162.200 174.200 162.500 175.800 ;
        RECT 165.400 175.600 165.800 179.900 ;
        RECT 163.700 175.300 165.800 175.600 ;
        RECT 163.700 175.200 164.100 175.300 ;
        RECT 164.500 174.900 164.900 175.000 ;
        RECT 163.000 174.600 164.900 174.900 ;
        RECT 163.000 174.500 163.400 174.600 ;
        RECT 157.000 173.900 162.500 174.200 ;
        RECT 157.000 173.800 157.800 173.900 ;
        RECT 152.900 172.800 153.800 173.100 ;
        RECT 151.700 172.400 152.100 172.800 ;
        RECT 152.900 171.100 153.300 172.800 ;
        RECT 156.600 171.100 157.000 173.500 ;
        RECT 159.100 173.200 159.400 173.900 ;
        RECT 161.900 173.800 162.300 173.900 ;
        RECT 165.400 173.600 165.800 175.300 ;
        RECT 163.900 173.300 165.800 173.600 ;
        RECT 163.900 173.200 164.300 173.300 ;
        RECT 158.200 172.100 158.600 172.500 ;
        RECT 159.000 172.400 159.400 173.200 ;
        RECT 165.400 173.100 165.800 173.300 ;
        RECT 167.000 175.100 167.400 179.900 ;
        RECT 169.700 176.400 170.100 179.900 ;
        RECT 171.800 177.500 172.200 179.500 ;
        RECT 169.300 176.100 170.100 176.400 ;
        RECT 168.600 175.100 169.000 175.600 ;
        RECT 167.000 174.800 169.000 175.100 ;
        RECT 166.200 173.100 166.600 173.200 ;
        RECT 165.400 172.800 166.600 173.100 ;
        RECT 159.900 172.700 160.300 172.800 ;
        RECT 159.900 172.400 161.300 172.700 ;
        RECT 161.000 172.100 161.300 172.400 ;
        RECT 163.000 172.100 163.400 172.500 ;
        RECT 158.200 171.800 159.200 172.100 ;
        RECT 158.800 171.100 159.200 171.800 ;
        RECT 161.000 171.100 161.400 172.100 ;
        RECT 163.000 171.800 163.700 172.100 ;
        RECT 163.100 171.100 163.700 171.800 ;
        RECT 165.400 171.100 165.800 172.800 ;
        RECT 166.200 172.400 166.600 172.800 ;
        RECT 167.000 171.100 167.400 174.800 ;
        RECT 169.300 174.200 169.600 176.100 ;
        RECT 171.900 175.800 172.200 177.500 ;
        RECT 170.300 175.500 172.200 175.800 ;
        RECT 172.600 175.700 173.000 179.900 ;
        RECT 174.800 178.200 175.200 179.900 ;
        RECT 174.200 177.900 175.200 178.200 ;
        RECT 177.000 177.900 177.400 179.900 ;
        RECT 179.100 177.900 179.700 179.900 ;
        RECT 174.200 177.500 174.600 177.900 ;
        RECT 177.000 177.600 177.300 177.900 ;
        RECT 175.900 177.300 177.700 177.600 ;
        RECT 179.000 177.500 179.400 177.900 ;
        RECT 175.900 177.200 176.300 177.300 ;
        RECT 177.300 177.200 177.700 177.300 ;
        RECT 174.200 176.500 174.600 176.600 ;
        RECT 176.500 176.500 176.900 176.600 ;
        RECT 174.200 176.200 176.900 176.500 ;
        RECT 177.200 176.500 178.300 176.800 ;
        RECT 177.200 175.900 177.500 176.500 ;
        RECT 177.900 176.400 178.300 176.500 ;
        RECT 179.100 176.600 179.800 177.000 ;
        RECT 179.100 176.100 179.400 176.600 ;
        RECT 175.100 175.700 177.500 175.900 ;
        RECT 172.600 175.600 177.500 175.700 ;
        RECT 178.200 175.800 179.400 176.100 ;
        RECT 172.600 175.500 175.500 175.600 ;
        RECT 170.300 174.500 170.600 175.500 ;
        RECT 172.600 175.400 175.400 175.500 ;
        RECT 167.800 174.100 168.200 174.200 ;
        RECT 168.600 174.100 169.600 174.200 ;
        RECT 169.900 174.100 170.600 174.500 ;
        RECT 171.000 174.400 171.400 175.200 ;
        RECT 171.800 174.400 172.200 175.200 ;
        RECT 175.800 175.100 176.200 175.200 ;
        RECT 173.700 174.800 176.200 175.100 ;
        RECT 173.700 174.700 174.100 174.800 ;
        RECT 174.500 174.200 174.900 174.300 ;
        RECT 178.200 174.200 178.500 175.800 ;
        RECT 181.400 175.600 181.800 179.900 ;
        RECT 179.700 175.300 181.800 175.600 ;
        RECT 179.700 175.200 180.100 175.300 ;
        RECT 180.500 174.900 180.900 175.000 ;
        RECT 179.000 174.600 180.900 174.900 ;
        RECT 179.000 174.500 179.400 174.600 ;
        RECT 167.800 173.800 169.600 174.100 ;
        RECT 169.300 173.500 169.600 173.800 ;
        RECT 170.100 173.900 170.600 174.100 ;
        RECT 173.000 173.900 178.500 174.200 ;
        RECT 170.100 173.600 172.200 173.900 ;
        RECT 173.000 173.800 173.800 173.900 ;
        RECT 169.300 173.300 169.700 173.500 ;
        RECT 169.300 173.000 170.100 173.300 ;
        RECT 169.700 171.500 170.100 173.000 ;
        RECT 171.900 172.500 172.200 173.600 ;
        RECT 171.800 171.500 172.200 172.500 ;
        RECT 172.600 171.100 173.000 173.500 ;
        RECT 175.100 173.200 175.400 173.900 ;
        RECT 177.900 173.800 178.300 173.900 ;
        RECT 181.400 173.600 181.800 175.300 ;
        RECT 179.900 173.300 181.800 173.600 ;
        RECT 179.900 173.200 180.300 173.300 ;
        RECT 174.200 172.100 174.600 172.500 ;
        RECT 175.000 172.400 175.400 173.200 ;
        RECT 175.900 172.700 176.300 172.800 ;
        RECT 175.900 172.400 177.300 172.700 ;
        RECT 177.000 172.100 177.300 172.400 ;
        RECT 179.000 172.100 179.400 172.500 ;
        RECT 174.200 171.800 175.200 172.100 ;
        RECT 174.800 171.100 175.200 171.800 ;
        RECT 177.000 171.100 177.400 172.100 ;
        RECT 179.000 171.800 179.700 172.100 ;
        RECT 179.100 171.100 179.700 171.800 ;
        RECT 181.400 171.100 181.800 173.300 ;
        RECT 182.200 175.600 182.600 179.900 ;
        RECT 184.300 177.900 184.900 179.900 ;
        RECT 186.600 177.900 187.000 179.900 ;
        RECT 188.800 178.200 189.200 179.900 ;
        RECT 188.800 177.900 189.800 178.200 ;
        RECT 184.600 177.500 185.000 177.900 ;
        RECT 186.700 177.600 187.000 177.900 ;
        RECT 186.300 177.300 188.100 177.600 ;
        RECT 189.400 177.500 189.800 177.900 ;
        RECT 186.300 177.200 186.700 177.300 ;
        RECT 187.700 177.200 188.100 177.300 ;
        RECT 184.200 176.600 184.900 177.000 ;
        RECT 183.800 175.600 184.200 176.200 ;
        RECT 184.600 176.100 184.900 176.600 ;
        RECT 185.700 176.500 186.800 176.800 ;
        RECT 185.700 176.400 186.100 176.500 ;
        RECT 184.600 175.800 185.800 176.100 ;
        RECT 182.200 175.300 184.300 175.600 ;
        RECT 182.200 173.600 182.600 175.300 ;
        RECT 183.900 175.200 184.300 175.300 ;
        RECT 185.500 175.200 185.800 175.800 ;
        RECT 186.500 175.900 186.800 176.500 ;
        RECT 187.100 176.500 187.500 176.600 ;
        RECT 189.400 176.500 189.800 176.600 ;
        RECT 187.100 176.200 189.800 176.500 ;
        RECT 186.500 175.700 188.900 175.900 ;
        RECT 191.000 175.700 191.400 179.900 ;
        RECT 186.500 175.600 191.400 175.700 ;
        RECT 188.500 175.500 191.400 175.600 ;
        RECT 191.800 177.500 192.200 179.500 ;
        RECT 191.800 175.800 192.100 177.500 ;
        RECT 193.900 176.400 194.300 179.900 ;
        RECT 193.900 176.100 194.700 176.400 ;
        RECT 194.200 175.800 194.700 176.100 ;
        RECT 191.800 175.500 193.700 175.800 ;
        RECT 188.600 175.400 191.400 175.500 ;
        RECT 183.100 174.900 183.500 175.000 ;
        RECT 183.100 174.600 185.000 174.900 ;
        RECT 185.400 174.800 185.800 175.200 ;
        RECT 187.800 175.100 188.200 175.200 ;
        RECT 187.800 174.800 190.300 175.100 ;
        RECT 184.600 174.500 185.000 174.600 ;
        RECT 185.500 174.200 185.800 174.800 ;
        RECT 189.900 174.700 190.300 174.800 ;
        RECT 191.800 174.400 192.200 175.200 ;
        RECT 192.600 174.400 193.000 175.200 ;
        RECT 193.400 174.500 193.700 175.500 ;
        RECT 189.100 174.200 189.500 174.300 ;
        RECT 185.500 173.900 191.000 174.200 ;
        RECT 193.400 174.100 194.100 174.500 ;
        RECT 194.400 174.200 194.700 175.800 ;
        RECT 196.600 175.700 197.000 179.900 ;
        RECT 198.800 178.200 199.200 179.900 ;
        RECT 198.200 177.900 199.200 178.200 ;
        RECT 201.000 177.900 201.400 179.900 ;
        RECT 203.100 177.900 203.700 179.900 ;
        RECT 198.200 177.500 198.600 177.900 ;
        RECT 201.000 177.600 201.300 177.900 ;
        RECT 199.900 177.300 201.700 177.600 ;
        RECT 203.000 177.500 203.400 177.900 ;
        RECT 199.900 177.200 200.300 177.300 ;
        RECT 201.300 177.200 201.700 177.300 ;
        RECT 198.200 176.500 198.600 176.600 ;
        RECT 200.500 176.500 200.900 176.600 ;
        RECT 198.200 176.200 200.900 176.500 ;
        RECT 201.200 176.500 202.300 176.800 ;
        RECT 201.200 175.900 201.500 176.500 ;
        RECT 201.900 176.400 202.300 176.500 ;
        RECT 203.100 176.600 203.800 177.000 ;
        RECT 203.100 176.100 203.400 176.600 ;
        RECT 199.100 175.700 201.500 175.900 ;
        RECT 196.600 175.600 201.500 175.700 ;
        RECT 202.200 175.800 203.400 176.100 ;
        RECT 195.000 174.800 195.400 175.600 ;
        RECT 196.600 175.500 199.500 175.600 ;
        RECT 196.600 175.400 199.400 175.500 ;
        RECT 199.800 175.100 200.200 175.200 ;
        RECT 197.700 174.800 200.200 175.100 ;
        RECT 197.700 174.700 198.100 174.800 ;
        RECT 199.000 174.700 199.400 174.800 ;
        RECT 198.500 174.200 198.900 174.300 ;
        RECT 202.200 174.200 202.500 175.800 ;
        RECT 205.400 175.600 205.800 179.900 ;
        RECT 203.700 175.300 205.800 175.600 ;
        RECT 203.700 175.200 204.100 175.300 ;
        RECT 204.500 174.900 204.900 175.000 ;
        RECT 203.000 174.600 204.900 174.900 ;
        RECT 203.000 174.500 203.400 174.600 ;
        RECT 193.400 173.900 193.900 174.100 ;
        RECT 185.700 173.800 186.100 173.900 ;
        RECT 182.200 173.300 184.100 173.600 ;
        RECT 182.200 171.100 182.600 173.300 ;
        RECT 183.700 173.200 184.100 173.300 ;
        RECT 188.600 172.800 188.900 173.900 ;
        RECT 190.200 173.800 191.000 173.900 ;
        RECT 191.800 173.600 193.900 173.900 ;
        RECT 194.400 173.800 195.400 174.200 ;
        RECT 197.000 173.900 202.500 174.200 ;
        RECT 197.000 173.800 197.800 173.900 ;
        RECT 187.700 172.700 188.100 172.800 ;
        RECT 184.600 172.100 185.000 172.500 ;
        RECT 186.700 172.400 188.100 172.700 ;
        RECT 188.600 172.400 189.000 172.800 ;
        RECT 186.700 172.100 187.000 172.400 ;
        RECT 189.400 172.100 189.800 172.500 ;
        RECT 184.300 171.800 185.000 172.100 ;
        RECT 184.300 171.100 184.900 171.800 ;
        RECT 186.600 171.100 187.000 172.100 ;
        RECT 188.800 171.800 189.800 172.100 ;
        RECT 188.800 171.100 189.200 171.800 ;
        RECT 191.000 171.100 191.400 173.500 ;
        RECT 191.800 172.500 192.100 173.600 ;
        RECT 194.400 173.500 194.700 173.800 ;
        RECT 194.300 173.300 194.700 173.500 ;
        RECT 193.900 173.000 194.700 173.300 ;
        RECT 191.800 171.500 192.200 172.500 ;
        RECT 193.900 171.500 194.300 173.000 ;
        RECT 196.600 171.100 197.000 173.500 ;
        RECT 199.100 172.800 199.400 173.900 ;
        RECT 201.900 173.800 202.300 173.900 ;
        RECT 205.400 173.600 205.800 175.300 ;
        RECT 203.900 173.300 205.800 173.600 ;
        RECT 203.900 173.200 204.300 173.300 ;
        RECT 198.200 172.100 198.600 172.500 ;
        RECT 199.000 172.400 199.400 172.800 ;
        RECT 199.900 172.700 200.300 172.800 ;
        RECT 199.900 172.400 201.300 172.700 ;
        RECT 201.000 172.100 201.300 172.400 ;
        RECT 203.000 172.100 203.400 172.500 ;
        RECT 198.200 171.800 199.200 172.100 ;
        RECT 198.800 171.100 199.200 171.800 ;
        RECT 201.000 171.100 201.400 172.100 ;
        RECT 203.000 171.800 203.700 172.100 ;
        RECT 203.100 171.100 203.700 171.800 ;
        RECT 205.400 171.100 205.800 173.300 ;
        RECT 206.200 177.100 206.600 179.900 ;
        RECT 207.000 177.100 207.400 177.200 ;
        RECT 206.200 176.800 207.400 177.100 ;
        RECT 206.200 171.100 206.600 176.800 ;
        RECT 209.400 175.800 209.800 176.600 ;
        RECT 207.000 172.400 207.400 173.200 ;
        RECT 210.200 173.100 210.600 179.900 ;
        RECT 211.800 176.200 212.200 179.900 ;
        RECT 213.400 179.600 215.400 179.900 ;
        RECT 213.400 176.200 213.800 179.600 ;
        RECT 211.800 175.900 213.800 176.200 ;
        RECT 214.200 175.900 214.600 179.300 ;
        RECT 215.000 175.900 215.400 179.600 ;
        RECT 215.800 179.600 217.800 179.900 ;
        RECT 215.800 175.900 216.200 179.600 ;
        RECT 216.600 175.900 217.000 179.300 ;
        RECT 217.400 176.200 217.800 179.600 ;
        RECT 219.000 176.200 219.400 179.900 ;
        RECT 221.700 179.200 222.100 179.900 ;
        RECT 221.400 178.800 222.100 179.200 ;
        RECT 221.700 176.400 222.100 178.800 ;
        RECT 223.800 177.500 224.200 179.500 ;
        RECT 217.400 175.900 219.400 176.200 ;
        RECT 221.300 176.100 222.100 176.400 ;
        RECT 214.200 175.600 214.500 175.900 ;
        RECT 216.700 175.600 217.000 175.900 ;
        RECT 212.200 175.200 212.600 175.400 ;
        RECT 213.500 175.300 214.500 175.600 ;
        RECT 213.500 175.200 213.800 175.300 ;
        RECT 211.000 175.100 211.400 175.200 ;
        RECT 211.800 175.100 212.600 175.200 ;
        RECT 211.000 174.900 212.600 175.100 ;
        RECT 211.000 174.800 212.200 174.900 ;
        RECT 213.400 174.800 213.800 175.200 ;
        RECT 215.000 175.100 215.400 175.600 ;
        RECT 215.800 175.100 216.200 175.600 ;
        RECT 216.700 175.300 217.700 175.600 ;
        RECT 215.000 174.800 216.200 175.100 ;
        RECT 217.400 175.200 217.700 175.300 ;
        RECT 218.600 175.200 219.000 175.400 ;
        RECT 217.400 174.800 217.800 175.200 ;
        RECT 218.600 175.100 219.400 175.200 ;
        RECT 219.800 175.100 220.200 175.200 ;
        RECT 218.600 174.900 220.200 175.100 ;
        RECT 219.000 174.800 220.200 174.900 ;
        RECT 220.600 174.800 221.000 175.600 ;
        RECT 211.000 173.400 211.400 174.200 ;
        RECT 212.600 173.800 213.000 174.600 ;
        RECT 213.500 173.200 213.800 174.800 ;
        RECT 214.100 174.400 214.500 174.800 ;
        RECT 214.200 174.200 214.500 174.400 ;
        RECT 216.700 174.400 217.100 174.800 ;
        RECT 216.700 174.200 217.000 174.400 ;
        RECT 214.200 173.800 214.600 174.200 ;
        RECT 216.600 173.800 217.000 174.200 ;
        RECT 213.400 173.100 213.800 173.200 ;
        RECT 217.400 173.100 217.700 174.800 ;
        RECT 218.200 173.800 218.600 174.600 ;
        RECT 221.300 174.200 221.600 176.100 ;
        RECT 223.900 175.800 224.200 177.500 ;
        RECT 222.300 175.500 224.200 175.800 ;
        RECT 224.600 177.500 225.000 179.500 ;
        RECT 224.600 175.800 224.900 177.500 ;
        RECT 226.700 176.400 227.100 179.900 ;
        RECT 229.800 176.800 230.200 177.200 ;
        RECT 226.700 176.100 227.500 176.400 ;
        RECT 229.800 176.200 230.100 176.800 ;
        RECT 230.500 176.200 230.900 179.900 ;
        RECT 233.000 176.800 233.400 177.200 ;
        RECT 233.000 176.200 233.300 176.800 ;
        RECT 233.700 176.200 234.100 179.900 ;
        RECT 224.600 175.500 226.500 175.800 ;
        RECT 222.300 174.500 222.600 175.500 ;
        RECT 220.600 173.800 221.600 174.200 ;
        RECT 221.900 174.100 222.600 174.500 ;
        RECT 223.000 174.400 223.400 175.200 ;
        RECT 223.800 174.400 224.200 175.200 ;
        RECT 224.600 174.400 225.000 175.200 ;
        RECT 225.400 174.400 225.800 175.200 ;
        RECT 226.200 174.500 226.500 175.500 ;
        RECT 221.300 173.500 221.600 173.800 ;
        RECT 222.100 173.900 222.600 174.100 ;
        RECT 226.200 174.100 226.900 174.500 ;
        RECT 227.200 174.200 227.500 176.100 ;
        RECT 229.400 175.900 230.100 176.200 ;
        RECT 229.400 175.800 229.800 175.900 ;
        RECT 230.400 175.800 231.400 176.200 ;
        RECT 232.600 175.900 233.300 176.200 ;
        RECT 233.600 175.900 234.100 176.200 ;
        RECT 232.600 175.800 233.000 175.900 ;
        RECT 227.800 175.100 228.200 175.600 ;
        RECT 229.400 175.100 229.700 175.800 ;
        RECT 227.800 174.800 229.700 175.100 ;
        RECT 230.400 174.200 230.700 175.800 ;
        RECT 233.600 175.200 233.900 175.900 ;
        RECT 235.800 175.800 236.200 176.600 ;
        RECT 231.000 174.400 231.400 175.200 ;
        RECT 233.400 174.800 233.900 175.200 ;
        RECT 233.600 174.200 233.900 174.800 ;
        RECT 234.200 174.400 234.600 175.200 ;
        RECT 226.200 173.900 226.700 174.100 ;
        RECT 222.100 173.600 224.200 173.900 ;
        RECT 221.300 173.300 221.700 173.500 ;
        RECT 209.700 172.800 210.600 173.100 ;
        RECT 209.700 172.200 210.100 172.800 ;
        RECT 209.700 171.800 210.600 172.200 ;
        RECT 209.700 171.100 210.100 171.800 ;
        RECT 213.300 171.100 214.100 173.100 ;
        RECT 217.100 172.200 217.900 173.100 ;
        RECT 221.300 173.000 222.100 173.300 ;
        RECT 216.600 171.800 217.900 172.200 ;
        RECT 217.100 171.100 217.900 171.800 ;
        RECT 221.700 171.500 222.100 173.000 ;
        RECT 223.900 172.500 224.200 173.600 ;
        RECT 223.800 171.500 224.200 172.500 ;
        RECT 224.600 173.600 226.700 173.900 ;
        RECT 227.200 173.800 228.200 174.200 ;
        RECT 229.400 173.800 230.700 174.200 ;
        RECT 231.800 174.100 232.200 174.200 ;
        RECT 231.400 173.800 232.200 174.100 ;
        RECT 232.600 173.800 233.900 174.200 ;
        RECT 235.000 174.100 235.400 174.200 ;
        RECT 234.600 173.800 235.400 174.100 ;
        RECT 224.600 172.500 224.900 173.600 ;
        RECT 227.200 173.500 227.500 173.800 ;
        RECT 227.100 173.300 227.500 173.500 ;
        RECT 226.700 173.000 227.500 173.300 ;
        RECT 229.500 173.100 229.800 173.800 ;
        RECT 231.400 173.600 231.800 173.800 ;
        RECT 230.300 173.100 232.100 173.300 ;
        RECT 232.700 173.100 233.000 173.800 ;
        RECT 234.600 173.600 235.000 173.800 ;
        RECT 233.500 173.100 235.300 173.300 ;
        RECT 236.600 173.100 237.000 179.900 ;
        RECT 237.400 177.100 237.800 177.200 ;
        RECT 238.200 177.100 238.600 179.900 ;
        RECT 240.300 177.900 240.900 179.900 ;
        RECT 242.600 177.900 243.000 179.900 ;
        RECT 244.800 178.200 245.200 179.900 ;
        RECT 244.800 177.900 245.800 178.200 ;
        RECT 240.600 177.500 241.000 177.900 ;
        RECT 242.700 177.600 243.000 177.900 ;
        RECT 242.300 177.300 244.100 177.600 ;
        RECT 245.400 177.500 245.800 177.900 ;
        RECT 242.300 177.200 242.700 177.300 ;
        RECT 243.700 177.200 244.100 177.300 ;
        RECT 237.400 176.800 238.600 177.100 ;
        RECT 238.200 175.600 238.600 176.800 ;
        RECT 240.200 176.600 240.900 177.000 ;
        RECT 240.600 176.100 240.900 176.600 ;
        RECT 241.700 176.500 242.800 176.800 ;
        RECT 241.700 176.400 242.100 176.500 ;
        RECT 240.600 175.800 241.800 176.100 ;
        RECT 238.200 175.300 240.300 175.600 ;
        RECT 237.400 173.400 237.800 174.200 ;
        RECT 238.200 173.600 238.600 175.300 ;
        RECT 239.900 175.200 240.300 175.300 ;
        RECT 239.100 174.900 239.500 175.000 ;
        RECT 239.100 174.600 241.000 174.900 ;
        RECT 240.600 174.500 241.000 174.600 ;
        RECT 241.500 174.200 241.800 175.800 ;
        RECT 242.500 175.900 242.800 176.500 ;
        RECT 243.100 176.500 243.500 176.600 ;
        RECT 245.400 176.500 245.800 176.600 ;
        RECT 243.100 176.200 245.800 176.500 ;
        RECT 242.500 175.700 244.900 175.900 ;
        RECT 247.000 175.700 247.400 179.900 ;
        RECT 248.200 176.800 248.600 177.200 ;
        RECT 248.200 176.200 248.500 176.800 ;
        RECT 248.900 176.200 249.300 179.900 ;
        RECT 247.800 175.900 248.500 176.200 ;
        RECT 248.800 175.900 249.300 176.200 ;
        RECT 247.800 175.800 248.200 175.900 ;
        RECT 242.500 175.600 247.400 175.700 ;
        RECT 244.500 175.500 247.400 175.600 ;
        RECT 244.600 175.400 247.400 175.500 ;
        RECT 248.800 175.200 249.100 175.900 ;
        RECT 251.000 175.600 251.400 179.900 ;
        RECT 253.100 177.900 253.700 179.900 ;
        RECT 255.400 177.900 255.800 179.900 ;
        RECT 257.600 178.200 258.000 179.900 ;
        RECT 257.600 177.900 258.600 178.200 ;
        RECT 253.400 177.500 253.800 177.900 ;
        RECT 255.500 177.600 255.800 177.900 ;
        RECT 255.100 177.300 256.900 177.600 ;
        RECT 258.200 177.500 258.600 177.900 ;
        RECT 255.100 177.200 255.500 177.300 ;
        RECT 256.500 177.200 256.900 177.300 ;
        RECT 253.000 176.600 253.700 177.000 ;
        RECT 253.400 176.100 253.700 176.600 ;
        RECT 254.500 176.500 255.600 176.800 ;
        RECT 254.500 176.400 254.900 176.500 ;
        RECT 253.400 175.800 254.600 176.100 ;
        RECT 251.000 175.300 253.100 175.600 ;
        RECT 243.800 175.100 244.200 175.200 ;
        RECT 243.800 174.800 246.300 175.100 ;
        RECT 248.600 174.800 249.100 175.200 ;
        RECT 245.900 174.700 246.300 174.800 ;
        RECT 245.100 174.200 245.500 174.300 ;
        RECT 248.800 174.200 249.100 174.800 ;
        RECT 249.400 174.400 249.800 175.200 ;
        RECT 241.500 173.900 247.000 174.200 ;
        RECT 241.700 173.800 242.100 173.900 ;
        RECT 224.600 171.500 225.000 172.500 ;
        RECT 226.700 172.200 227.100 173.000 ;
        RECT 226.200 171.800 227.100 172.200 ;
        RECT 226.700 171.500 227.100 171.800 ;
        RECT 229.400 171.100 229.800 173.100 ;
        RECT 230.200 173.000 232.200 173.100 ;
        RECT 230.200 171.100 230.600 173.000 ;
        RECT 231.800 171.100 232.200 173.000 ;
        RECT 232.600 171.100 233.000 173.100 ;
        RECT 233.400 173.000 235.400 173.100 ;
        RECT 233.400 171.100 233.800 173.000 ;
        RECT 235.000 171.100 235.400 173.000 ;
        RECT 236.100 172.800 237.000 173.100 ;
        RECT 238.200 173.300 240.100 173.600 ;
        RECT 236.100 172.200 236.500 172.800 ;
        RECT 235.800 171.800 236.500 172.200 ;
        RECT 236.100 171.100 236.500 171.800 ;
        RECT 238.200 171.100 238.600 173.300 ;
        RECT 239.700 173.200 240.100 173.300 ;
        RECT 244.600 173.200 244.900 173.900 ;
        RECT 246.200 173.800 247.000 173.900 ;
        RECT 247.800 173.800 249.100 174.200 ;
        RECT 250.200 174.100 250.600 174.200 ;
        RECT 249.800 173.800 250.600 174.100 ;
        RECT 243.700 172.700 244.100 172.800 ;
        RECT 240.600 172.100 241.000 172.500 ;
        RECT 242.700 172.400 244.100 172.700 ;
        RECT 244.600 172.400 245.000 173.200 ;
        RECT 242.700 172.100 243.000 172.400 ;
        RECT 245.400 172.100 245.800 172.500 ;
        RECT 240.300 171.800 241.000 172.100 ;
        RECT 240.300 171.100 240.900 171.800 ;
        RECT 242.600 171.100 243.000 172.100 ;
        RECT 244.800 171.800 245.800 172.100 ;
        RECT 244.800 171.100 245.200 171.800 ;
        RECT 247.000 171.100 247.400 173.500 ;
        RECT 247.900 173.100 248.200 173.800 ;
        RECT 249.800 173.600 250.200 173.800 ;
        RECT 251.000 173.600 251.400 175.300 ;
        RECT 252.700 175.200 253.100 175.300 ;
        RECT 251.900 174.900 252.300 175.000 ;
        RECT 251.900 174.600 253.800 174.900 ;
        RECT 253.400 174.500 253.800 174.600 ;
        RECT 254.300 174.200 254.600 175.800 ;
        RECT 255.300 175.900 255.600 176.500 ;
        RECT 255.900 176.500 256.300 176.600 ;
        RECT 258.200 176.500 258.600 176.600 ;
        RECT 255.900 176.200 258.600 176.500 ;
        RECT 255.300 175.700 257.700 175.900 ;
        RECT 259.800 175.700 260.200 179.900 ;
        RECT 260.600 175.800 261.000 176.600 ;
        RECT 255.300 175.600 260.200 175.700 ;
        RECT 257.300 175.500 260.200 175.600 ;
        RECT 257.400 175.400 260.200 175.500 ;
        RECT 256.600 175.100 257.000 175.200 ;
        RECT 256.600 174.800 259.100 175.100 ;
        RECT 258.700 174.700 259.100 174.800 ;
        RECT 257.900 174.200 258.300 174.300 ;
        RECT 254.300 173.900 259.800 174.200 ;
        RECT 254.500 173.800 254.900 173.900 ;
        RECT 251.000 173.300 252.900 173.600 ;
        RECT 248.700 173.100 250.500 173.300 ;
        RECT 247.800 171.100 248.200 173.100 ;
        RECT 248.600 173.000 250.600 173.100 ;
        RECT 248.600 171.100 249.000 173.000 ;
        RECT 250.200 171.100 250.600 173.000 ;
        RECT 251.000 171.100 251.400 173.300 ;
        RECT 252.500 173.200 252.900 173.300 ;
        RECT 257.400 172.800 257.700 173.900 ;
        RECT 259.000 173.800 259.800 173.900 ;
        RECT 256.500 172.700 256.900 172.800 ;
        RECT 253.400 172.100 253.800 172.500 ;
        RECT 255.500 172.400 256.900 172.700 ;
        RECT 257.400 172.400 257.800 172.800 ;
        RECT 255.500 172.100 255.800 172.400 ;
        RECT 258.200 172.100 258.600 172.500 ;
        RECT 253.100 171.800 253.800 172.100 ;
        RECT 253.100 171.100 253.700 171.800 ;
        RECT 255.400 171.100 255.800 172.100 ;
        RECT 257.600 171.800 258.600 172.100 ;
        RECT 257.600 171.100 258.000 171.800 ;
        RECT 259.800 171.100 260.200 173.500 ;
        RECT 261.400 173.100 261.800 179.900 ;
        RECT 260.900 172.800 261.800 173.100 ;
        RECT 260.900 172.200 261.300 172.800 ;
        RECT 260.900 171.800 261.800 172.200 ;
        RECT 260.900 171.100 261.300 171.800 ;
        RECT 0.600 167.500 1.000 169.900 ;
        RECT 2.800 169.200 3.200 169.900 ;
        RECT 2.200 168.900 3.200 169.200 ;
        RECT 5.000 168.900 5.400 169.900 ;
        RECT 7.100 169.200 7.700 169.900 ;
        RECT 7.000 168.900 7.700 169.200 ;
        RECT 2.200 168.500 2.600 168.900 ;
        RECT 5.000 168.600 5.300 168.900 ;
        RECT 3.000 168.200 3.400 168.600 ;
        RECT 3.900 168.300 5.300 168.600 ;
        RECT 7.000 168.500 7.400 168.900 ;
        RECT 3.900 168.200 4.300 168.300 ;
        RECT 1.000 167.100 1.800 167.200 ;
        RECT 3.100 167.100 3.400 168.200 ;
        RECT 7.900 167.700 8.300 167.800 ;
        RECT 9.400 167.700 9.800 169.900 ;
        RECT 11.500 168.200 11.900 169.900 ;
        RECT 7.900 167.400 9.800 167.700 ;
        RECT 11.000 167.900 11.900 168.200 ;
        RECT 12.600 167.900 13.000 169.900 ;
        RECT 13.400 168.000 13.800 169.900 ;
        RECT 15.000 168.000 15.400 169.900 ;
        RECT 13.400 167.900 15.400 168.000 ;
        RECT 5.900 167.100 6.300 167.200 ;
        RECT 9.400 167.100 9.800 167.400 ;
        RECT 10.200 167.100 10.600 167.600 ;
        RECT 1.000 166.800 6.500 167.100 ;
        RECT 2.500 166.700 2.900 166.800 ;
        RECT 1.700 166.200 2.100 166.300 ;
        RECT 1.700 165.900 4.200 166.200 ;
        RECT 3.800 165.800 4.200 165.900 ;
        RECT 0.600 165.500 3.400 165.600 ;
        RECT 0.600 165.400 3.500 165.500 ;
        RECT 0.600 165.300 5.500 165.400 ;
        RECT 0.600 161.100 1.000 165.300 ;
        RECT 3.100 165.100 5.500 165.300 ;
        RECT 2.200 164.500 4.900 164.800 ;
        RECT 2.200 164.400 2.600 164.500 ;
        RECT 4.500 164.400 4.900 164.500 ;
        RECT 5.200 164.500 5.500 165.100 ;
        RECT 6.200 165.200 6.500 166.800 ;
        RECT 9.400 166.800 10.600 167.100 ;
        RECT 7.000 166.400 7.400 166.500 ;
        RECT 7.000 166.100 8.900 166.400 ;
        RECT 8.500 166.000 8.900 166.100 ;
        RECT 7.700 165.700 8.100 165.800 ;
        RECT 9.400 165.700 9.800 166.800 ;
        RECT 7.700 165.400 9.800 165.700 ;
        RECT 6.200 164.900 7.400 165.200 ;
        RECT 5.900 164.500 6.300 164.600 ;
        RECT 5.200 164.200 6.300 164.500 ;
        RECT 7.100 164.400 7.400 164.900 ;
        RECT 7.100 164.000 7.800 164.400 ;
        RECT 3.900 163.700 4.300 163.800 ;
        RECT 5.300 163.700 5.700 163.800 ;
        RECT 2.200 163.100 2.600 163.500 ;
        RECT 3.900 163.400 5.700 163.700 ;
        RECT 5.000 163.100 5.300 163.400 ;
        RECT 7.000 163.100 7.400 163.500 ;
        RECT 2.200 162.800 3.200 163.100 ;
        RECT 2.800 161.100 3.200 162.800 ;
        RECT 5.000 161.100 5.400 163.100 ;
        RECT 7.100 161.100 7.700 163.100 ;
        RECT 9.400 161.100 9.800 165.400 ;
        RECT 11.000 166.100 11.400 167.900 ;
        RECT 12.700 167.200 13.000 167.900 ;
        RECT 13.500 167.700 15.300 167.900 ;
        RECT 15.800 167.500 16.200 169.900 ;
        RECT 18.000 169.200 18.400 169.900 ;
        RECT 17.400 168.900 18.400 169.200 ;
        RECT 20.200 168.900 20.600 169.900 ;
        RECT 22.300 169.200 22.900 169.900 ;
        RECT 22.200 168.900 22.900 169.200 ;
        RECT 17.400 168.500 17.800 168.900 ;
        RECT 20.200 168.600 20.500 168.900 ;
        RECT 18.200 168.200 18.600 168.600 ;
        RECT 19.100 168.300 20.500 168.600 ;
        RECT 22.200 168.500 22.600 168.900 ;
        RECT 19.100 168.200 19.500 168.300 ;
        RECT 14.600 167.200 15.000 167.400 ;
        RECT 11.800 167.100 12.200 167.200 ;
        RECT 12.600 167.100 13.900 167.200 ;
        RECT 11.800 166.800 13.900 167.100 ;
        RECT 14.600 166.900 15.400 167.200 ;
        RECT 15.000 166.800 15.400 166.900 ;
        RECT 16.200 167.100 17.000 167.200 ;
        RECT 18.300 167.100 18.600 168.200 ;
        RECT 24.600 168.100 25.000 169.900 ;
        RECT 25.400 168.100 25.800 168.600 ;
        RECT 24.600 167.800 25.800 168.100 ;
        RECT 23.100 167.700 23.500 167.800 ;
        RECT 24.600 167.700 25.000 167.800 ;
        RECT 23.100 167.400 25.000 167.700 ;
        RECT 21.100 167.100 21.500 167.200 ;
        RECT 16.200 166.800 21.700 167.100 ;
        RECT 11.000 165.800 12.900 166.100 ;
        RECT 11.000 161.100 11.400 165.800 ;
        RECT 12.600 165.200 12.900 165.800 ;
        RECT 11.800 164.400 12.200 165.200 ;
        RECT 12.600 165.100 13.000 165.200 ;
        RECT 13.600 165.100 13.900 166.800 ;
        RECT 17.700 166.700 18.100 166.800 ;
        RECT 14.200 165.800 14.600 166.600 ;
        RECT 16.900 166.200 17.300 166.300 ;
        RECT 16.900 166.100 19.400 166.200 ;
        RECT 20.600 166.100 21.000 166.200 ;
        RECT 16.900 165.900 21.000 166.100 ;
        RECT 19.000 165.800 21.000 165.900 ;
        RECT 15.800 165.500 18.600 165.600 ;
        RECT 15.800 165.400 18.700 165.500 ;
        RECT 15.800 165.300 20.700 165.400 ;
        RECT 12.600 164.800 13.300 165.100 ;
        RECT 13.600 164.800 14.100 165.100 ;
        RECT 13.000 164.200 13.300 164.800 ;
        RECT 13.000 163.800 13.400 164.200 ;
        RECT 13.700 161.100 14.100 164.800 ;
        RECT 15.800 161.100 16.200 165.300 ;
        RECT 18.300 165.100 20.700 165.300 ;
        RECT 17.400 164.500 20.100 164.800 ;
        RECT 17.400 164.400 17.800 164.500 ;
        RECT 19.700 164.400 20.100 164.500 ;
        RECT 20.400 164.500 20.700 165.100 ;
        RECT 21.400 165.200 21.700 166.800 ;
        RECT 22.200 166.400 22.600 166.500 ;
        RECT 22.200 166.100 24.100 166.400 ;
        RECT 23.700 166.000 24.100 166.100 ;
        RECT 22.900 165.700 23.300 165.800 ;
        RECT 24.600 165.700 25.000 167.400 ;
        RECT 22.900 165.400 25.000 165.700 ;
        RECT 21.400 164.900 22.600 165.200 ;
        RECT 21.100 164.500 21.500 164.600 ;
        RECT 20.400 164.200 21.500 164.500 ;
        RECT 22.300 164.400 22.600 164.900 ;
        RECT 22.300 164.000 23.000 164.400 ;
        RECT 19.100 163.700 19.500 163.800 ;
        RECT 20.500 163.700 20.900 163.800 ;
        RECT 17.400 163.100 17.800 163.500 ;
        RECT 19.100 163.400 20.900 163.700 ;
        RECT 20.200 163.100 20.500 163.400 ;
        RECT 22.200 163.100 22.600 163.500 ;
        RECT 17.400 162.800 18.400 163.100 ;
        RECT 18.000 161.100 18.400 162.800 ;
        RECT 20.200 161.100 20.600 163.100 ;
        RECT 22.300 161.100 22.900 163.100 ;
        RECT 24.600 161.100 25.000 165.400 ;
        RECT 26.200 166.100 26.600 169.900 ;
        RECT 28.900 168.000 29.300 169.500 ;
        RECT 31.000 168.500 31.400 169.500 ;
        RECT 28.500 167.700 29.300 168.000 ;
        RECT 28.500 167.500 28.900 167.700 ;
        RECT 28.500 167.200 28.800 167.500 ;
        RECT 31.100 167.400 31.400 168.500 ;
        RECT 33.100 168.200 33.500 169.900 ;
        RECT 32.600 167.900 33.500 168.200 ;
        RECT 27.800 166.800 28.800 167.200 ;
        RECT 29.300 167.100 31.400 167.400 ;
        RECT 29.300 166.900 29.800 167.100 ;
        RECT 27.800 166.100 28.200 166.200 ;
        RECT 26.200 165.800 28.200 166.100 ;
        RECT 26.200 161.100 26.600 165.800 ;
        RECT 27.800 165.400 28.200 165.800 ;
        RECT 28.500 165.200 28.800 166.800 ;
        RECT 29.100 166.500 29.800 166.900 ;
        RECT 31.800 166.800 32.200 167.600 ;
        RECT 29.500 165.500 29.800 166.500 ;
        RECT 30.200 165.800 30.600 166.600 ;
        RECT 31.000 166.100 31.400 166.600 ;
        RECT 31.800 166.100 32.200 166.200 ;
        RECT 31.000 165.800 32.200 166.100 ;
        RECT 32.600 166.100 33.000 167.900 ;
        RECT 34.200 167.800 34.600 169.900 ;
        RECT 35.000 168.000 35.400 169.900 ;
        RECT 36.600 168.000 37.000 169.900 ;
        RECT 35.000 167.900 37.000 168.000 ;
        RECT 37.400 167.900 37.800 169.900 ;
        RECT 38.200 168.000 38.600 169.900 ;
        RECT 39.800 168.000 40.200 169.900 ;
        RECT 38.200 167.900 40.200 168.000 ;
        RECT 34.300 167.200 34.600 167.800 ;
        RECT 35.100 167.700 36.900 167.900 ;
        RECT 36.200 167.200 36.600 167.400 ;
        RECT 37.500 167.200 37.800 167.900 ;
        RECT 38.300 167.700 40.100 167.900 ;
        RECT 40.600 167.700 41.000 169.900 ;
        RECT 42.700 169.200 43.300 169.900 ;
        RECT 42.700 168.900 43.400 169.200 ;
        RECT 45.000 168.900 45.400 169.900 ;
        RECT 47.200 169.200 47.600 169.900 ;
        RECT 47.200 168.900 48.200 169.200 ;
        RECT 43.000 168.500 43.400 168.900 ;
        RECT 45.100 168.600 45.400 168.900 ;
        RECT 45.100 168.300 46.500 168.600 ;
        RECT 46.100 168.200 46.500 168.300 ;
        RECT 47.000 168.200 47.400 168.600 ;
        RECT 47.800 168.500 48.200 168.900 ;
        RECT 42.100 167.700 42.500 167.800 ;
        RECT 40.600 167.400 42.500 167.700 ;
        RECT 39.400 167.200 39.800 167.400 ;
        RECT 34.200 166.800 35.500 167.200 ;
        RECT 36.200 166.900 37.000 167.200 ;
        RECT 36.600 166.800 37.000 166.900 ;
        RECT 37.400 166.800 38.700 167.200 ;
        RECT 39.400 166.900 40.200 167.200 ;
        RECT 39.800 166.800 40.200 166.900 ;
        RECT 32.600 165.800 34.500 166.100 ;
        RECT 29.500 165.200 31.400 165.500 ;
        RECT 28.500 164.900 29.000 165.200 ;
        RECT 28.500 164.600 29.300 164.900 ;
        RECT 28.900 161.100 29.300 164.600 ;
        RECT 31.100 163.500 31.400 165.200 ;
        RECT 31.000 161.500 31.400 163.500 ;
        RECT 32.600 161.100 33.000 165.800 ;
        RECT 34.200 165.200 34.500 165.800 ;
        RECT 33.400 164.400 33.800 165.200 ;
        RECT 34.200 165.100 34.600 165.200 ;
        RECT 35.200 165.100 35.500 166.800 ;
        RECT 35.800 165.800 36.200 166.600 ;
        RECT 38.400 165.200 38.700 166.800 ;
        RECT 39.000 165.800 39.400 166.600 ;
        RECT 40.600 165.700 41.000 167.400 ;
        RECT 44.100 167.100 44.500 167.200 ;
        RECT 47.000 167.100 47.300 168.200 ;
        RECT 49.400 167.500 49.800 169.900 ;
        RECT 50.300 168.200 50.700 168.600 ;
        RECT 50.200 167.800 50.600 168.200 ;
        RECT 51.000 167.900 51.400 169.900 ;
        RECT 48.600 167.100 49.400 167.200 ;
        RECT 43.900 166.800 49.400 167.100 ;
        RECT 43.000 166.400 43.400 166.500 ;
        RECT 41.500 166.100 43.400 166.400 ;
        RECT 41.500 166.000 41.900 166.100 ;
        RECT 42.300 165.700 42.700 165.800 ;
        RECT 40.600 165.400 42.700 165.700 ;
        RECT 37.400 165.100 37.800 165.200 ;
        RECT 34.200 164.800 34.900 165.100 ;
        RECT 35.200 164.800 35.700 165.100 ;
        RECT 37.400 164.800 38.100 165.100 ;
        RECT 38.400 164.800 39.400 165.200 ;
        RECT 34.600 164.200 34.900 164.800 ;
        RECT 34.600 163.800 35.000 164.200 ;
        RECT 35.300 161.100 35.700 164.800 ;
        RECT 37.800 164.200 38.100 164.800 ;
        RECT 37.800 163.800 38.200 164.200 ;
        RECT 38.500 161.100 38.900 164.800 ;
        RECT 40.600 161.100 41.000 165.400 ;
        RECT 43.900 165.200 44.200 166.800 ;
        RECT 47.500 166.700 47.900 166.800 ;
        RECT 48.300 166.200 48.700 166.300 ;
        RECT 51.100 166.200 51.400 167.900 ;
        RECT 55.000 167.700 55.400 169.900 ;
        RECT 57.100 169.200 57.700 169.900 ;
        RECT 57.100 168.900 57.800 169.200 ;
        RECT 59.400 168.900 59.800 169.900 ;
        RECT 61.600 169.200 62.000 169.900 ;
        RECT 61.600 168.900 62.600 169.200 ;
        RECT 57.400 168.500 57.800 168.900 ;
        RECT 59.500 168.600 59.800 168.900 ;
        RECT 59.500 168.300 60.900 168.600 ;
        RECT 60.500 168.200 60.900 168.300 ;
        RECT 61.400 168.200 61.800 168.600 ;
        RECT 62.200 168.500 62.600 168.900 ;
        RECT 56.500 167.700 56.900 167.800 ;
        RECT 55.000 167.400 56.900 167.700 ;
        RECT 51.800 166.400 52.200 167.200 ;
        RECT 46.200 165.900 48.700 166.200 ;
        RECT 50.200 166.100 50.600 166.200 ;
        RECT 51.000 166.100 51.400 166.200 ;
        RECT 52.600 166.100 53.000 166.200 ;
        RECT 53.400 166.100 53.800 166.200 ;
        RECT 46.200 165.800 46.600 165.900 ;
        RECT 50.200 165.800 51.400 166.100 ;
        RECT 52.200 165.800 53.800 166.100 ;
        RECT 47.000 165.500 49.800 165.600 ;
        RECT 46.900 165.400 49.800 165.500 ;
        RECT 43.000 164.900 44.200 165.200 ;
        RECT 44.900 165.300 49.800 165.400 ;
        RECT 44.900 165.100 47.300 165.300 ;
        RECT 43.000 164.400 43.300 164.900 ;
        RECT 42.600 164.000 43.300 164.400 ;
        RECT 44.100 164.500 44.500 164.600 ;
        RECT 44.900 164.500 45.200 165.100 ;
        RECT 44.100 164.200 45.200 164.500 ;
        RECT 45.500 164.500 48.200 164.800 ;
        RECT 45.500 164.400 45.900 164.500 ;
        RECT 47.800 164.400 48.200 164.500 ;
        RECT 44.700 163.700 45.100 163.800 ;
        RECT 46.100 163.700 46.500 163.800 ;
        RECT 43.000 163.100 43.400 163.500 ;
        RECT 44.700 163.400 46.500 163.700 ;
        RECT 45.100 163.100 45.400 163.400 ;
        RECT 47.800 163.100 48.200 163.500 ;
        RECT 42.700 161.100 43.300 163.100 ;
        RECT 45.000 161.100 45.400 163.100 ;
        RECT 47.200 162.800 48.200 163.100 ;
        RECT 47.200 161.100 47.600 162.800 ;
        RECT 49.400 161.100 49.800 165.300 ;
        RECT 50.300 165.100 50.600 165.800 ;
        RECT 52.200 165.600 52.600 165.800 ;
        RECT 55.000 165.700 55.400 167.400 ;
        RECT 58.500 167.100 58.900 167.200 ;
        RECT 61.400 167.100 61.700 168.200 ;
        RECT 63.800 167.500 64.200 169.900 ;
        RECT 65.900 168.200 66.300 169.900 ;
        RECT 65.400 167.900 66.300 168.200 ;
        RECT 67.000 167.900 67.400 169.900 ;
        RECT 67.800 168.000 68.200 169.900 ;
        RECT 69.400 168.000 69.800 169.900 ;
        RECT 67.800 167.900 69.800 168.000 ;
        RECT 63.000 167.100 63.800 167.200 ;
        RECT 58.300 166.800 63.800 167.100 ;
        RECT 64.600 166.800 65.000 167.600 ;
        RECT 57.400 166.400 57.800 166.500 ;
        RECT 55.900 166.100 57.800 166.400 ;
        RECT 58.300 166.200 58.600 166.800 ;
        RECT 61.900 166.700 62.300 166.800 ;
        RECT 62.700 166.200 63.100 166.300 ;
        RECT 55.900 166.000 56.300 166.100 ;
        RECT 58.200 165.800 58.600 166.200 ;
        RECT 59.800 166.100 60.200 166.200 ;
        RECT 60.600 166.100 63.100 166.200 ;
        RECT 59.800 165.900 63.100 166.100 ;
        RECT 65.400 166.100 65.800 167.900 ;
        RECT 67.100 167.200 67.400 167.900 ;
        RECT 67.900 167.700 69.700 167.900 ;
        RECT 70.200 167.700 70.600 169.900 ;
        RECT 72.300 169.200 72.900 169.900 ;
        RECT 72.300 168.900 73.000 169.200 ;
        RECT 74.600 168.900 75.000 169.900 ;
        RECT 76.800 169.200 77.200 169.900 ;
        RECT 76.800 168.900 77.800 169.200 ;
        RECT 72.600 168.500 73.000 168.900 ;
        RECT 74.700 168.600 75.000 168.900 ;
        RECT 74.700 168.300 76.100 168.600 ;
        RECT 75.700 168.200 76.100 168.300 ;
        RECT 76.600 167.800 77.000 168.600 ;
        RECT 77.400 168.500 77.800 168.900 ;
        RECT 71.700 167.700 72.100 167.800 ;
        RECT 70.200 167.400 72.100 167.700 ;
        RECT 69.000 167.200 69.400 167.400 ;
        RECT 67.000 166.800 68.300 167.200 ;
        RECT 69.000 166.900 69.800 167.200 ;
        RECT 69.400 166.800 69.800 166.900 ;
        RECT 68.000 166.200 68.300 166.800 ;
        RECT 59.800 165.800 61.000 165.900 ;
        RECT 65.400 165.800 67.300 166.100 ;
        RECT 67.800 165.800 68.300 166.200 ;
        RECT 68.600 166.100 69.000 166.600 ;
        RECT 69.400 166.100 69.800 166.200 ;
        RECT 68.600 165.800 69.800 166.100 ;
        RECT 56.700 165.700 57.100 165.800 ;
        RECT 55.000 165.400 57.100 165.700 ;
        RECT 50.200 161.100 50.600 165.100 ;
        RECT 51.000 164.800 53.000 165.100 ;
        RECT 51.000 161.100 51.400 164.800 ;
        RECT 52.600 161.100 53.000 164.800 ;
        RECT 55.000 161.100 55.400 165.400 ;
        RECT 58.300 165.200 58.600 165.800 ;
        RECT 61.400 165.500 64.200 165.600 ;
        RECT 61.300 165.400 64.200 165.500 ;
        RECT 57.400 164.900 58.600 165.200 ;
        RECT 59.300 165.300 64.200 165.400 ;
        RECT 59.300 165.100 61.700 165.300 ;
        RECT 57.400 164.400 57.700 164.900 ;
        RECT 57.000 164.000 57.700 164.400 ;
        RECT 58.500 164.500 58.900 164.600 ;
        RECT 59.300 164.500 59.600 165.100 ;
        RECT 58.500 164.200 59.600 164.500 ;
        RECT 59.900 164.500 62.600 164.800 ;
        RECT 59.900 164.400 60.300 164.500 ;
        RECT 62.200 164.400 62.600 164.500 ;
        RECT 59.100 163.700 59.500 163.800 ;
        RECT 60.500 163.700 60.900 163.800 ;
        RECT 57.400 163.100 57.800 163.500 ;
        RECT 59.100 163.400 60.900 163.700 ;
        RECT 59.500 163.100 59.800 163.400 ;
        RECT 62.200 163.100 62.600 163.500 ;
        RECT 57.100 161.100 57.700 163.100 ;
        RECT 59.400 161.100 59.800 163.100 ;
        RECT 61.600 162.800 62.600 163.100 ;
        RECT 61.600 161.100 62.000 162.800 ;
        RECT 63.800 161.100 64.200 165.300 ;
        RECT 65.400 161.100 65.800 165.800 ;
        RECT 67.000 165.200 67.300 165.800 ;
        RECT 66.200 164.400 66.600 165.200 ;
        RECT 67.000 165.100 67.400 165.200 ;
        RECT 68.000 165.100 68.300 165.800 ;
        RECT 70.200 165.700 70.600 167.400 ;
        RECT 73.700 167.100 74.100 167.200 ;
        RECT 76.600 167.100 76.900 167.800 ;
        RECT 79.000 167.500 79.400 169.900 ;
        RECT 80.600 167.600 81.000 169.900 ;
        RECT 82.200 167.600 82.600 169.900 ;
        RECT 83.800 167.600 84.200 169.900 ;
        RECT 85.400 167.600 85.800 169.900 ;
        RECT 88.900 168.000 89.300 169.500 ;
        RECT 91.000 168.500 91.400 169.500 ;
        RECT 88.500 167.700 89.300 168.000 ;
        RECT 80.600 167.200 81.500 167.600 ;
        RECT 82.200 167.200 83.300 167.600 ;
        RECT 83.800 167.200 84.900 167.600 ;
        RECT 85.400 167.200 86.600 167.600 ;
        RECT 88.500 167.500 88.900 167.700 ;
        RECT 88.500 167.200 88.800 167.500 ;
        RECT 91.100 167.400 91.400 168.500 ;
        RECT 93.700 168.000 94.100 169.500 ;
        RECT 95.800 168.500 96.200 169.500 ;
        RECT 78.200 167.100 79.000 167.200 ;
        RECT 73.500 166.800 79.000 167.100 ;
        RECT 79.800 166.900 80.200 167.200 ;
        RECT 81.100 166.900 81.500 167.200 ;
        RECT 82.900 166.900 83.300 167.200 ;
        RECT 84.500 166.900 84.900 167.200 ;
        RECT 72.600 166.400 73.000 166.500 ;
        RECT 71.100 166.100 73.000 166.400 ;
        RECT 71.100 166.000 71.500 166.100 ;
        RECT 71.900 165.700 72.300 165.800 ;
        RECT 70.200 165.400 72.300 165.700 ;
        RECT 67.000 164.800 67.700 165.100 ;
        RECT 68.000 164.800 68.500 165.100 ;
        RECT 67.400 164.200 67.700 164.800 ;
        RECT 67.400 163.800 67.800 164.200 ;
        RECT 68.100 161.100 68.500 164.800 ;
        RECT 70.200 161.100 70.600 165.400 ;
        RECT 73.500 165.200 73.800 166.800 ;
        RECT 77.100 166.700 77.500 166.800 ;
        RECT 79.800 166.500 80.700 166.900 ;
        RECT 81.100 166.500 82.400 166.900 ;
        RECT 82.900 166.500 84.100 166.900 ;
        RECT 84.500 166.500 85.800 166.900 ;
        RECT 77.900 166.200 78.300 166.300 ;
        RECT 75.800 165.900 78.300 166.200 ;
        RECT 75.800 165.800 76.200 165.900 ;
        RECT 81.100 165.800 81.500 166.500 ;
        RECT 82.900 165.800 83.300 166.500 ;
        RECT 84.500 165.800 84.900 166.500 ;
        RECT 86.200 165.800 86.600 167.200 ;
        RECT 87.000 166.800 87.400 167.200 ;
        RECT 87.800 166.800 88.800 167.200 ;
        RECT 89.300 167.100 91.400 167.400 ;
        RECT 93.300 167.700 94.100 168.000 ;
        RECT 93.300 167.500 93.700 167.700 ;
        RECT 93.300 167.200 93.600 167.500 ;
        RECT 95.900 167.400 96.200 168.500 ;
        RECT 97.900 168.200 98.300 169.900 ;
        RECT 97.400 167.900 98.300 168.200 ;
        RECT 99.000 168.500 99.400 169.500 ;
        RECT 89.300 166.900 89.800 167.100 ;
        RECT 87.000 166.100 87.300 166.800 ;
        RECT 87.800 166.100 88.200 166.200 ;
        RECT 87.000 165.800 88.200 166.100 ;
        RECT 76.600 165.500 79.400 165.600 ;
        RECT 76.500 165.400 79.400 165.500 ;
        RECT 72.600 164.900 73.800 165.200 ;
        RECT 74.500 165.300 79.400 165.400 ;
        RECT 74.500 165.100 76.900 165.300 ;
        RECT 72.600 164.400 72.900 164.900 ;
        RECT 72.200 164.000 72.900 164.400 ;
        RECT 73.700 164.500 74.100 164.600 ;
        RECT 74.500 164.500 74.800 165.100 ;
        RECT 73.700 164.200 74.800 164.500 ;
        RECT 75.100 164.500 77.800 164.800 ;
        RECT 75.100 164.400 75.500 164.500 ;
        RECT 77.400 164.400 77.800 164.500 ;
        RECT 74.300 163.700 74.700 163.800 ;
        RECT 75.700 163.700 76.100 163.800 ;
        RECT 72.600 163.100 73.000 163.500 ;
        RECT 74.300 163.400 76.100 163.700 ;
        RECT 74.700 163.100 75.000 163.400 ;
        RECT 77.400 163.100 77.800 163.500 ;
        RECT 72.300 161.100 72.900 163.100 ;
        RECT 74.600 161.100 75.000 163.100 ;
        RECT 76.800 162.800 77.800 163.100 ;
        RECT 76.800 161.100 77.200 162.800 ;
        RECT 79.000 161.100 79.400 165.300 ;
        RECT 80.600 165.400 81.500 165.800 ;
        RECT 82.200 165.400 83.300 165.800 ;
        RECT 83.800 165.400 84.900 165.800 ;
        RECT 85.400 165.400 86.600 165.800 ;
        RECT 87.800 165.400 88.200 165.800 ;
        RECT 80.600 161.100 81.000 165.400 ;
        RECT 82.200 161.100 82.600 165.400 ;
        RECT 83.800 161.100 84.200 165.400 ;
        RECT 85.400 161.100 85.800 165.400 ;
        RECT 88.500 165.200 88.800 166.800 ;
        RECT 89.100 166.500 89.800 166.900 ;
        RECT 92.600 166.800 93.600 167.200 ;
        RECT 94.100 167.100 96.200 167.400 ;
        RECT 94.100 166.900 94.600 167.100 ;
        RECT 89.500 165.500 89.800 166.500 ;
        RECT 90.200 165.800 90.600 166.600 ;
        RECT 91.000 165.800 91.400 166.600 ;
        RECT 93.300 166.200 93.600 166.800 ;
        RECT 93.900 166.500 94.600 166.900 ;
        RECT 96.600 166.800 97.000 167.600 ;
        RECT 89.500 165.200 91.400 165.500 ;
        RECT 92.600 165.400 93.000 166.200 ;
        RECT 93.300 165.800 93.800 166.200 ;
        RECT 88.500 164.900 89.000 165.200 ;
        RECT 88.500 164.600 89.300 164.900 ;
        RECT 88.900 161.100 89.300 164.600 ;
        RECT 91.100 163.500 91.400 165.200 ;
        RECT 93.300 164.900 93.600 165.800 ;
        RECT 94.300 165.500 94.600 166.500 ;
        RECT 95.000 165.800 95.400 166.600 ;
        RECT 95.800 165.800 96.200 166.600 ;
        RECT 94.300 165.200 96.200 165.500 ;
        RECT 93.300 164.600 94.100 164.900 ;
        RECT 91.000 161.500 91.400 163.500 ;
        RECT 93.700 161.100 94.100 164.600 ;
        RECT 95.900 163.500 96.200 165.200 ;
        RECT 95.800 161.500 96.200 163.500 ;
        RECT 97.400 161.100 97.800 167.900 ;
        RECT 99.000 167.400 99.300 168.500 ;
        RECT 101.100 168.000 101.500 169.500 ;
        RECT 101.100 167.700 101.900 168.000 ;
        RECT 101.500 167.500 101.900 167.700 ;
        RECT 105.400 167.500 105.800 169.900 ;
        RECT 107.600 169.200 108.000 169.900 ;
        RECT 107.000 168.900 108.000 169.200 ;
        RECT 109.800 168.900 110.200 169.900 ;
        RECT 111.900 169.200 112.500 169.900 ;
        RECT 111.800 168.900 112.500 169.200 ;
        RECT 107.000 168.500 107.400 168.900 ;
        RECT 109.800 168.600 110.100 168.900 ;
        RECT 107.800 168.200 108.200 168.600 ;
        RECT 108.700 168.300 110.100 168.600 ;
        RECT 111.800 168.500 112.200 168.900 ;
        RECT 108.700 168.200 109.100 168.300 ;
        RECT 99.000 167.100 101.100 167.400 ;
        RECT 100.600 166.900 101.100 167.100 ;
        RECT 101.600 167.200 101.900 167.500 ;
        RECT 101.600 167.100 102.600 167.200 ;
        RECT 104.600 167.100 105.000 167.200 ;
        RECT 99.000 165.800 99.400 166.600 ;
        RECT 99.800 165.800 100.200 166.600 ;
        RECT 100.600 166.500 101.300 166.900 ;
        RECT 101.600 166.800 105.000 167.100 ;
        RECT 105.800 167.100 106.600 167.200 ;
        RECT 107.900 167.100 108.200 168.200 ;
        RECT 114.200 168.100 114.600 169.900 ;
        RECT 115.000 168.100 115.400 168.600 ;
        RECT 114.200 167.800 115.400 168.100 ;
        RECT 112.700 167.700 113.100 167.800 ;
        RECT 114.200 167.700 114.600 167.800 ;
        RECT 112.700 167.400 114.600 167.700 ;
        RECT 110.700 167.100 111.100 167.200 ;
        RECT 105.800 166.800 111.300 167.100 ;
        RECT 100.600 165.500 100.900 166.500 ;
        RECT 99.000 165.200 100.900 165.500 ;
        RECT 98.200 164.400 98.600 165.200 ;
        RECT 99.000 163.500 99.300 165.200 ;
        RECT 101.600 164.900 101.900 166.800 ;
        RECT 107.300 166.700 107.700 166.800 ;
        RECT 106.500 166.200 106.900 166.300 ;
        RECT 102.200 165.400 102.600 166.200 ;
        RECT 106.500 165.900 109.000 166.200 ;
        RECT 108.600 165.800 109.000 165.900 ;
        RECT 105.400 165.500 108.200 165.600 ;
        RECT 105.400 165.400 108.300 165.500 ;
        RECT 101.100 164.600 101.900 164.900 ;
        RECT 105.400 165.300 110.300 165.400 ;
        RECT 99.000 161.500 99.400 163.500 ;
        RECT 101.100 161.100 101.500 164.600 ;
        RECT 105.400 161.100 105.800 165.300 ;
        RECT 107.900 165.100 110.300 165.300 ;
        RECT 107.000 164.500 109.700 164.800 ;
        RECT 107.000 164.400 107.400 164.500 ;
        RECT 109.300 164.400 109.700 164.500 ;
        RECT 110.000 164.500 110.300 165.100 ;
        RECT 111.000 165.200 111.300 166.800 ;
        RECT 111.800 166.400 112.200 166.500 ;
        RECT 111.800 166.100 113.700 166.400 ;
        RECT 113.300 166.000 113.700 166.100 ;
        RECT 114.200 166.100 114.600 167.400 ;
        RECT 115.000 166.800 115.400 167.200 ;
        RECT 115.000 166.100 115.300 166.800 ;
        RECT 114.200 165.800 115.300 166.100 ;
        RECT 115.800 166.100 116.200 169.900 ;
        RECT 118.500 168.000 118.900 169.500 ;
        RECT 120.600 168.500 121.000 169.500 ;
        RECT 118.100 167.700 118.900 168.000 ;
        RECT 118.100 167.500 118.500 167.700 ;
        RECT 118.100 167.200 118.400 167.500 ;
        RECT 120.700 167.400 121.000 168.500 ;
        RECT 116.600 167.100 117.000 167.200 ;
        RECT 117.400 167.100 118.400 167.200 ;
        RECT 116.600 166.800 118.400 167.100 ;
        RECT 118.900 167.100 121.000 167.400 ;
        RECT 121.400 167.600 121.800 169.900 ;
        RECT 123.000 168.200 123.400 169.900 ;
        RECT 124.600 168.500 125.000 169.500 ;
        RECT 123.000 167.900 123.500 168.200 ;
        RECT 121.400 167.300 122.700 167.600 ;
        RECT 118.900 166.900 119.400 167.100 ;
        RECT 117.400 166.100 117.800 166.200 ;
        RECT 115.800 165.800 117.800 166.100 ;
        RECT 112.500 165.700 112.900 165.800 ;
        RECT 114.200 165.700 114.600 165.800 ;
        RECT 112.500 165.400 114.600 165.700 ;
        RECT 111.000 164.900 112.200 165.200 ;
        RECT 110.700 164.500 111.100 164.600 ;
        RECT 110.000 164.200 111.100 164.500 ;
        RECT 111.900 164.400 112.200 164.900 ;
        RECT 111.900 164.000 112.600 164.400 ;
        RECT 108.700 163.700 109.100 163.800 ;
        RECT 110.100 163.700 110.500 163.800 ;
        RECT 107.000 163.100 107.400 163.500 ;
        RECT 108.700 163.400 110.500 163.700 ;
        RECT 109.800 163.100 110.100 163.400 ;
        RECT 111.800 163.100 112.200 163.500 ;
        RECT 107.000 162.800 108.000 163.100 ;
        RECT 107.600 161.100 108.000 162.800 ;
        RECT 109.800 161.100 110.200 163.100 ;
        RECT 111.900 161.100 112.500 163.100 ;
        RECT 114.200 161.100 114.600 165.400 ;
        RECT 115.800 161.100 116.200 165.800 ;
        RECT 117.400 165.400 117.800 165.800 ;
        RECT 118.100 164.900 118.400 166.800 ;
        RECT 118.700 166.500 119.400 166.900 ;
        RECT 119.100 165.500 119.400 166.500 ;
        RECT 119.800 165.800 120.200 166.600 ;
        RECT 120.600 165.800 121.000 166.600 ;
        RECT 121.500 166.200 121.900 166.600 ;
        RECT 121.400 165.800 121.900 166.200 ;
        RECT 122.400 166.500 122.700 167.300 ;
        RECT 123.200 167.200 123.500 167.900 ;
        RECT 123.000 166.800 123.500 167.200 ;
        RECT 124.600 167.400 124.900 168.500 ;
        RECT 126.700 168.000 127.100 169.500 ;
        RECT 129.400 168.500 129.800 169.500 ;
        RECT 126.700 167.700 127.500 168.000 ;
        RECT 127.100 167.500 127.500 167.700 ;
        RECT 124.600 167.100 126.700 167.400 ;
        RECT 122.400 166.100 122.900 166.500 ;
        RECT 119.100 165.200 121.000 165.500 ;
        RECT 118.100 164.600 118.900 164.900 ;
        RECT 118.500 161.100 118.900 164.600 ;
        RECT 120.700 163.500 121.000 165.200 ;
        RECT 122.400 165.100 122.700 166.100 ;
        RECT 123.200 165.100 123.500 166.800 ;
        RECT 126.200 166.900 126.700 167.100 ;
        RECT 127.200 167.200 127.500 167.500 ;
        RECT 129.400 167.400 129.700 168.500 ;
        RECT 131.500 168.000 131.900 169.500 ;
        RECT 136.100 168.200 136.500 169.500 ;
        RECT 138.200 168.500 138.600 169.500 ;
        RECT 136.100 168.000 137.000 168.200 ;
        RECT 131.500 167.700 132.300 168.000 ;
        RECT 131.900 167.500 132.300 167.700 ;
        RECT 127.200 167.100 128.200 167.200 ;
        RECT 128.600 167.100 129.000 167.200 ;
        RECT 129.400 167.100 131.500 167.400 ;
        RECT 124.600 165.800 125.000 166.600 ;
        RECT 125.400 165.800 125.800 166.600 ;
        RECT 126.200 166.500 126.900 166.900 ;
        RECT 127.200 166.800 129.000 167.100 ;
        RECT 131.000 166.900 131.500 167.100 ;
        RECT 132.000 167.200 132.300 167.500 ;
        RECT 135.700 167.800 137.000 168.000 ;
        RECT 135.700 167.700 136.500 167.800 ;
        RECT 135.700 167.500 136.100 167.700 ;
        RECT 135.700 167.200 136.000 167.500 ;
        RECT 138.300 167.400 138.600 168.500 ;
        RECT 140.300 167.900 141.100 169.900 ;
        RECT 144.300 168.200 144.700 169.900 ;
        RECT 143.800 167.900 144.700 168.200 ;
        RECT 145.400 168.000 145.800 169.900 ;
        RECT 147.000 168.000 147.400 169.900 ;
        RECT 145.400 167.900 147.400 168.000 ;
        RECT 147.800 167.900 148.200 169.900 ;
        RECT 150.100 167.900 150.900 169.900 ;
        RECT 154.500 168.000 154.900 169.500 ;
        RECT 156.600 168.500 157.000 169.500 ;
        RECT 160.900 169.200 161.300 169.500 ;
        RECT 160.600 168.800 161.300 169.200 ;
        RECT 132.000 167.100 133.000 167.200 ;
        RECT 126.200 165.500 126.500 166.500 ;
        RECT 120.600 161.500 121.000 163.500 ;
        RECT 121.400 164.800 122.700 165.100 ;
        RECT 121.400 161.100 121.800 164.800 ;
        RECT 123.000 164.600 123.500 165.100 ;
        RECT 124.600 165.200 126.500 165.500 ;
        RECT 123.000 161.100 123.400 164.600 ;
        RECT 124.600 163.500 124.900 165.200 ;
        RECT 127.200 164.900 127.500 166.800 ;
        RECT 127.800 165.400 128.200 166.200 ;
        RECT 129.400 165.800 129.800 166.600 ;
        RECT 130.200 165.800 130.600 166.600 ;
        RECT 131.000 166.500 131.700 166.900 ;
        RECT 132.000 166.800 134.500 167.100 ;
        RECT 135.000 166.800 136.000 167.200 ;
        RECT 136.500 167.100 138.600 167.400 ;
        RECT 140.600 167.200 140.900 167.900 ;
        RECT 136.500 166.900 137.000 167.100 ;
        RECT 131.000 165.500 131.300 166.500 ;
        RECT 126.700 164.600 127.500 164.900 ;
        RECT 129.400 165.200 131.300 165.500 ;
        RECT 124.600 161.500 125.000 163.500 ;
        RECT 126.700 161.100 127.100 164.600 ;
        RECT 129.400 163.500 129.700 165.200 ;
        RECT 132.000 164.900 132.300 166.800 ;
        RECT 132.600 165.400 133.000 166.200 ;
        RECT 134.200 166.100 134.500 166.800 ;
        RECT 135.000 166.100 135.400 166.200 ;
        RECT 134.200 165.800 135.400 166.100 ;
        RECT 135.000 165.400 135.400 165.800 ;
        RECT 131.500 164.600 132.300 164.900 ;
        RECT 135.700 164.900 136.000 166.800 ;
        RECT 136.300 166.500 137.000 166.900 ;
        RECT 139.800 166.800 140.200 167.200 ;
        RECT 139.900 166.600 140.200 166.800 ;
        RECT 140.600 166.800 141.000 167.200 ;
        RECT 136.700 165.500 137.000 166.500 ;
        RECT 137.400 165.800 137.800 166.600 ;
        RECT 138.200 165.800 138.600 166.600 ;
        RECT 139.900 166.200 140.300 166.600 ;
        RECT 140.600 166.200 140.900 166.800 ;
        RECT 141.400 166.400 141.800 167.200 ;
        RECT 143.000 166.800 143.400 167.600 ;
        RECT 143.800 167.100 144.200 167.900 ;
        RECT 145.500 167.700 147.300 167.900 ;
        RECT 145.800 167.200 146.200 167.400 ;
        RECT 147.800 167.200 148.100 167.900 ;
        RECT 150.300 167.200 150.600 167.900 ;
        RECT 154.100 167.700 154.900 168.000 ;
        RECT 154.100 167.500 154.500 167.700 ;
        RECT 154.100 167.200 154.400 167.500 ;
        RECT 156.700 167.400 157.000 168.500 ;
        RECT 160.900 168.000 161.300 168.800 ;
        RECT 163.000 168.500 163.400 169.500 ;
        RECT 145.400 167.100 146.200 167.200 ;
        RECT 143.800 166.900 146.200 167.100 ;
        RECT 143.800 166.800 145.800 166.900 ;
        RECT 146.900 166.800 148.200 167.200 ;
        RECT 136.700 165.200 138.600 165.500 ;
        RECT 139.000 165.400 139.400 166.200 ;
        RECT 140.600 165.800 141.000 166.200 ;
        RECT 142.200 166.100 142.600 166.200 ;
        RECT 141.800 165.800 142.600 166.100 ;
        RECT 140.600 165.700 140.900 165.800 ;
        RECT 139.900 165.400 140.900 165.700 ;
        RECT 141.800 165.600 142.200 165.800 ;
        RECT 135.700 164.600 136.500 164.900 ;
        RECT 129.400 161.500 129.800 163.500 ;
        RECT 131.500 161.100 131.900 164.600 ;
        RECT 136.100 161.100 136.500 164.600 ;
        RECT 138.300 163.500 138.600 165.200 ;
        RECT 139.900 165.100 140.200 165.400 ;
        RECT 138.200 161.500 138.600 163.500 ;
        RECT 139.000 161.400 139.400 165.100 ;
        RECT 139.800 161.700 140.200 165.100 ;
        RECT 140.600 164.800 142.600 165.100 ;
        RECT 140.600 161.400 141.000 164.800 ;
        RECT 139.000 161.100 141.000 161.400 ;
        RECT 142.200 161.100 142.600 164.800 ;
        RECT 143.800 161.100 144.200 166.800 ;
        RECT 146.200 165.800 146.600 166.600 ;
        RECT 144.600 164.400 145.000 165.200 ;
        RECT 146.900 165.100 147.200 166.800 ;
        RECT 149.400 166.400 149.800 167.200 ;
        RECT 150.200 166.800 150.600 167.200 ;
        RECT 150.300 166.200 150.600 166.800 ;
        RECT 151.000 167.100 151.400 167.200 ;
        RECT 152.600 167.100 153.000 167.200 ;
        RECT 151.000 166.800 153.000 167.100 ;
        RECT 153.400 166.800 154.400 167.200 ;
        RECT 154.900 167.100 157.000 167.400 ;
        RECT 160.500 167.700 161.300 168.000 ;
        RECT 160.500 167.500 160.900 167.700 ;
        RECT 160.500 167.200 160.800 167.500 ;
        RECT 163.100 167.400 163.400 168.500 ;
        RECT 154.900 166.900 155.400 167.100 ;
        RECT 151.000 166.600 151.300 166.800 ;
        RECT 150.900 166.200 151.300 166.600 ;
        RECT 148.600 166.100 149.000 166.200 ;
        RECT 148.600 165.800 149.400 166.100 ;
        RECT 150.200 165.800 150.600 166.200 ;
        RECT 149.000 165.600 149.400 165.800 ;
        RECT 150.300 165.700 150.600 165.800 ;
        RECT 150.300 165.400 151.300 165.700 ;
        RECT 151.800 165.400 152.200 166.200 ;
        RECT 153.400 165.400 153.800 166.200 ;
        RECT 147.800 165.100 148.200 165.200 ;
        RECT 151.000 165.100 151.300 165.400 ;
        RECT 154.100 165.200 154.400 166.800 ;
        RECT 154.700 166.500 155.400 166.900 ;
        RECT 159.800 166.800 160.800 167.200 ;
        RECT 161.300 167.100 163.400 167.400 ;
        RECT 163.800 168.500 164.200 169.500 ;
        RECT 163.800 167.400 164.100 168.500 ;
        RECT 165.900 168.000 166.300 169.500 ;
        RECT 168.600 168.000 169.000 169.900 ;
        RECT 170.200 168.000 170.600 169.900 ;
        RECT 165.900 167.700 166.700 168.000 ;
        RECT 168.600 167.900 170.600 168.000 ;
        RECT 171.000 167.900 171.400 169.900 ;
        RECT 171.800 168.500 172.200 169.500 ;
        RECT 168.700 167.700 170.500 167.900 ;
        RECT 166.300 167.500 166.700 167.700 ;
        RECT 163.800 167.100 165.900 167.400 ;
        RECT 161.300 166.900 161.800 167.100 ;
        RECT 155.100 165.500 155.400 166.500 ;
        RECT 155.800 165.800 156.200 166.600 ;
        RECT 156.600 166.100 157.000 166.600 ;
        RECT 158.200 166.100 158.600 166.200 ;
        RECT 156.600 165.800 158.600 166.100 ;
        RECT 155.100 165.200 157.000 165.500 ;
        RECT 159.800 165.400 160.200 166.200 ;
        RECT 146.700 164.800 147.200 165.100 ;
        RECT 147.500 164.800 148.200 165.100 ;
        RECT 148.600 164.800 150.600 165.100 ;
        RECT 146.700 161.100 147.100 164.800 ;
        RECT 147.500 164.200 147.800 164.800 ;
        RECT 147.400 163.800 147.800 164.200 ;
        RECT 148.600 161.100 149.000 164.800 ;
        RECT 150.200 161.400 150.600 164.800 ;
        RECT 151.000 161.700 151.400 165.100 ;
        RECT 151.800 161.400 152.200 165.100 ;
        RECT 154.100 164.900 154.600 165.200 ;
        RECT 154.100 164.600 154.900 164.900 ;
        RECT 150.200 161.100 152.200 161.400 ;
        RECT 154.500 161.100 154.900 164.600 ;
        RECT 156.700 163.500 157.000 165.200 ;
        RECT 160.500 164.900 160.800 166.800 ;
        RECT 161.100 166.500 161.800 166.900 ;
        RECT 165.400 166.900 165.900 167.100 ;
        RECT 166.400 167.200 166.700 167.500 ;
        RECT 169.000 167.200 169.400 167.400 ;
        RECT 171.000 167.200 171.300 167.900 ;
        RECT 171.800 167.400 172.100 168.500 ;
        RECT 173.900 168.000 174.300 169.500 ;
        RECT 176.600 168.500 177.000 169.500 ;
        RECT 178.700 169.200 179.100 169.500 ;
        RECT 178.700 168.800 179.400 169.200 ;
        RECT 173.900 167.700 174.700 168.000 ;
        RECT 174.300 167.500 174.700 167.700 ;
        RECT 161.500 165.500 161.800 166.500 ;
        RECT 162.200 165.800 162.600 166.600 ;
        RECT 163.000 165.800 163.400 166.600 ;
        RECT 163.800 165.800 164.200 166.600 ;
        RECT 164.600 165.800 165.000 166.600 ;
        RECT 165.400 166.500 166.100 166.900 ;
        RECT 166.400 166.800 167.400 167.200 ;
        RECT 168.600 166.900 169.400 167.200 ;
        RECT 168.600 166.800 169.000 166.900 ;
        RECT 170.100 166.800 171.400 167.200 ;
        RECT 171.800 167.100 173.900 167.400 ;
        RECT 173.400 166.900 173.900 167.100 ;
        RECT 174.400 167.200 174.700 167.500 ;
        RECT 176.600 167.400 176.900 168.500 ;
        RECT 178.700 168.000 179.100 168.800 ;
        RECT 178.700 167.700 179.500 168.000 ;
        RECT 179.100 167.500 179.500 167.700 ;
        RECT 165.400 165.500 165.700 166.500 ;
        RECT 161.500 165.200 163.400 165.500 ;
        RECT 160.500 164.600 161.300 164.900 ;
        RECT 156.600 161.500 157.000 163.500 ;
        RECT 160.900 161.100 161.300 164.600 ;
        RECT 163.100 163.500 163.400 165.200 ;
        RECT 163.000 161.500 163.400 163.500 ;
        RECT 163.800 165.200 165.700 165.500 ;
        RECT 163.800 163.500 164.100 165.200 ;
        RECT 166.400 164.900 166.700 166.800 ;
        RECT 167.000 166.100 167.400 166.200 ;
        RECT 167.800 166.100 168.200 166.200 ;
        RECT 167.000 165.800 168.200 166.100 ;
        RECT 169.400 165.800 169.800 166.600 ;
        RECT 167.000 165.400 167.400 165.800 ;
        RECT 170.100 165.100 170.400 166.800 ;
        RECT 171.800 165.800 172.200 166.600 ;
        RECT 172.600 165.800 173.000 166.600 ;
        RECT 173.400 166.500 174.100 166.900 ;
        RECT 174.400 166.800 175.400 167.200 ;
        RECT 176.600 167.100 178.700 167.400 ;
        RECT 178.200 166.900 178.700 167.100 ;
        RECT 179.200 167.200 179.500 167.500 ;
        RECT 183.000 167.900 183.400 169.900 ;
        RECT 185.400 168.900 185.800 169.900 ;
        RECT 183.700 168.200 184.100 168.600 ;
        RECT 173.400 165.500 173.700 166.500 ;
        RECT 171.800 165.200 173.700 165.500 ;
        RECT 174.400 165.200 174.700 166.800 ;
        RECT 175.000 165.400 175.400 166.200 ;
        RECT 176.600 165.800 177.000 166.600 ;
        RECT 177.400 165.800 177.800 166.600 ;
        RECT 178.200 166.500 178.900 166.900 ;
        RECT 179.200 166.800 180.200 167.200 ;
        RECT 178.200 165.500 178.500 166.500 ;
        RECT 171.000 165.100 171.400 165.200 ;
        RECT 165.900 164.600 166.700 164.900 ;
        RECT 169.900 164.800 170.400 165.100 ;
        RECT 170.700 164.800 171.400 165.100 ;
        RECT 163.800 161.500 164.200 163.500 ;
        RECT 165.900 163.200 166.300 164.600 ;
        RECT 165.400 162.800 166.300 163.200 ;
        RECT 165.900 161.100 166.300 162.800 ;
        RECT 169.900 161.100 170.300 164.800 ;
        RECT 170.700 164.200 171.000 164.800 ;
        RECT 170.600 163.800 171.000 164.200 ;
        RECT 171.800 163.500 172.100 165.200 ;
        RECT 174.200 164.900 174.700 165.200 ;
        RECT 173.900 164.600 174.700 164.900 ;
        RECT 176.600 165.200 178.500 165.500 ;
        RECT 171.800 161.500 172.200 163.500 ;
        RECT 173.900 161.100 174.300 164.600 ;
        RECT 176.600 163.500 176.900 165.200 ;
        RECT 179.200 164.900 179.500 166.800 ;
        RECT 182.200 166.400 182.600 167.200 ;
        RECT 179.800 165.400 180.200 166.200 ;
        RECT 181.400 166.100 181.800 166.200 ;
        RECT 183.000 166.100 183.300 167.900 ;
        RECT 183.800 167.800 184.200 168.200 ;
        RECT 184.600 167.800 185.000 168.600 ;
        RECT 183.800 167.100 184.100 167.800 ;
        RECT 185.500 167.200 185.800 168.900 ;
        RECT 188.500 167.900 189.300 169.900 ;
        RECT 191.300 168.200 191.700 169.900 ;
        RECT 191.300 167.900 192.200 168.200 ;
        RECT 193.400 168.000 193.800 169.900 ;
        RECT 195.000 168.000 195.400 169.900 ;
        RECT 193.400 167.900 195.400 168.000 ;
        RECT 195.800 167.900 196.200 169.900 ;
        RECT 198.100 169.200 198.900 169.900 ;
        RECT 198.100 168.800 199.400 169.200 ;
        RECT 198.100 167.900 198.900 168.800 ;
        RECT 200.600 167.900 201.000 169.900 ;
        RECT 201.400 168.000 201.800 169.900 ;
        RECT 203.000 168.000 203.400 169.900 ;
        RECT 201.400 167.900 203.400 168.000 ;
        RECT 185.400 167.100 185.800 167.200 ;
        RECT 183.800 166.800 185.800 167.100 ;
        RECT 183.800 166.100 184.200 166.200 ;
        RECT 181.400 165.800 182.200 166.100 ;
        RECT 183.000 165.800 184.200 166.100 ;
        RECT 181.800 165.600 182.200 165.800 ;
        RECT 183.800 165.100 184.100 165.800 ;
        RECT 185.500 165.100 185.800 166.800 ;
        RECT 187.800 166.400 188.200 167.200 ;
        RECT 188.700 166.200 189.000 167.900 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 189.400 166.600 189.700 166.800 ;
        RECT 189.300 166.200 189.700 166.600 ;
        RECT 186.200 165.400 186.600 166.200 ;
        RECT 187.000 166.100 187.400 166.200 ;
        RECT 187.000 165.800 187.800 166.100 ;
        RECT 188.600 165.800 189.000 166.200 ;
        RECT 187.400 165.600 187.800 165.800 ;
        RECT 188.700 165.700 189.000 165.800 ;
        RECT 188.700 165.400 189.700 165.700 ;
        RECT 190.200 165.400 190.600 166.200 ;
        RECT 191.800 166.100 192.200 167.900 ;
        RECT 193.500 167.700 195.300 167.900 ;
        RECT 192.600 166.800 193.000 167.600 ;
        RECT 193.800 167.200 194.200 167.400 ;
        RECT 195.800 167.200 196.100 167.900 ;
        RECT 193.400 166.900 194.200 167.200 ;
        RECT 193.400 166.800 193.800 166.900 ;
        RECT 194.900 166.800 196.200 167.200 ;
        RECT 196.600 167.100 197.000 167.200 ;
        RECT 197.400 167.100 197.800 167.200 ;
        RECT 196.600 166.800 197.800 167.100 ;
        RECT 193.400 166.100 193.700 166.800 ;
        RECT 191.800 165.800 193.700 166.100 ;
        RECT 194.200 165.800 194.600 166.600 ;
        RECT 189.400 165.200 189.700 165.400 ;
        RECT 178.700 164.600 179.500 164.900 ;
        RECT 181.400 164.800 183.400 165.100 ;
        RECT 176.600 161.500 177.000 163.500 ;
        RECT 178.700 161.100 179.100 164.600 ;
        RECT 181.400 161.100 181.800 164.800 ;
        RECT 183.000 161.100 183.400 164.800 ;
        RECT 183.800 161.100 184.200 165.100 ;
        RECT 185.400 164.700 186.300 165.100 ;
        RECT 185.900 161.100 186.300 164.700 ;
        RECT 187.000 164.800 189.000 165.100 ;
        RECT 187.000 161.100 187.400 164.800 ;
        RECT 188.600 161.400 189.000 164.800 ;
        RECT 189.400 161.700 189.800 165.200 ;
        RECT 190.200 161.400 190.600 165.100 ;
        RECT 191.000 164.400 191.400 165.200 ;
        RECT 188.600 161.100 190.600 161.400 ;
        RECT 191.800 161.100 192.200 165.800 ;
        RECT 194.900 165.100 195.200 166.800 ;
        RECT 197.400 166.400 197.800 166.800 ;
        RECT 198.300 166.200 198.600 167.900 ;
        RECT 200.700 167.200 201.000 167.900 ;
        RECT 201.500 167.700 203.300 167.900 ;
        RECT 205.400 167.700 205.800 169.900 ;
        RECT 207.500 169.200 208.100 169.900 ;
        RECT 207.500 168.900 208.200 169.200 ;
        RECT 209.800 168.900 210.200 169.900 ;
        RECT 212.000 169.200 212.400 169.900 ;
        RECT 212.000 168.900 213.000 169.200 ;
        RECT 207.800 168.500 208.200 168.900 ;
        RECT 209.900 168.600 210.200 168.900 ;
        RECT 209.900 168.300 211.300 168.600 ;
        RECT 210.900 168.200 211.300 168.300 ;
        RECT 211.800 168.200 212.200 168.600 ;
        RECT 212.600 168.500 213.000 168.900 ;
        RECT 206.900 167.700 207.300 167.800 ;
        RECT 205.400 167.400 207.300 167.700 ;
        RECT 202.600 167.200 203.000 167.400 ;
        RECT 199.000 166.800 199.400 167.200 ;
        RECT 200.600 166.800 201.900 167.200 ;
        RECT 202.600 166.900 203.400 167.200 ;
        RECT 203.000 166.800 203.400 166.900 ;
        RECT 199.000 166.600 199.300 166.800 ;
        RECT 198.900 166.200 199.300 166.600 ;
        RECT 195.800 166.100 196.200 166.200 ;
        RECT 196.600 166.100 197.000 166.200 ;
        RECT 195.800 165.800 197.400 166.100 ;
        RECT 198.200 165.800 198.600 166.200 ;
        RECT 197.000 165.600 197.400 165.800 ;
        RECT 198.300 165.700 198.600 165.800 ;
        RECT 198.300 165.400 199.300 165.700 ;
        RECT 199.800 165.400 200.200 166.200 ;
        RECT 200.600 165.800 201.000 166.200 ;
        RECT 195.800 165.100 196.200 165.200 ;
        RECT 199.000 165.100 199.300 165.400 ;
        RECT 200.600 165.200 200.900 165.800 ;
        RECT 200.600 165.100 201.000 165.200 ;
        RECT 201.600 165.100 201.900 166.800 ;
        RECT 202.200 165.800 202.600 166.600 ;
        RECT 205.400 165.700 205.800 167.400 ;
        RECT 208.900 167.100 209.300 167.200 ;
        RECT 211.800 167.100 212.100 168.200 ;
        RECT 214.200 167.500 214.600 169.900 ;
        RECT 215.000 167.800 215.400 168.600 ;
        RECT 215.000 167.200 215.300 167.800 ;
        RECT 213.400 167.100 214.200 167.200 ;
        RECT 208.700 166.800 214.200 167.100 ;
        RECT 215.000 166.800 215.400 167.200 ;
        RECT 207.800 166.400 208.200 166.500 ;
        RECT 206.300 166.100 208.200 166.400 ;
        RECT 206.300 166.000 206.700 166.100 ;
        RECT 207.100 165.700 207.500 165.800 ;
        RECT 205.400 165.400 207.500 165.700 ;
        RECT 194.700 164.800 195.200 165.100 ;
        RECT 195.500 164.800 196.200 165.100 ;
        RECT 196.600 164.800 198.600 165.100 ;
        RECT 194.700 161.100 195.100 164.800 ;
        RECT 195.500 164.200 195.800 164.800 ;
        RECT 195.400 163.800 195.800 164.200 ;
        RECT 196.600 161.100 197.000 164.800 ;
        RECT 198.200 161.400 198.600 164.800 ;
        RECT 199.000 161.700 199.400 165.100 ;
        RECT 199.800 161.400 200.200 165.100 ;
        RECT 200.600 164.800 201.300 165.100 ;
        RECT 201.600 164.800 202.100 165.100 ;
        RECT 201.000 164.200 201.300 164.800 ;
        RECT 201.000 163.800 201.400 164.200 ;
        RECT 198.200 161.100 200.200 161.400 ;
        RECT 201.700 162.200 202.100 164.800 ;
        RECT 201.700 161.800 202.600 162.200 ;
        RECT 201.700 161.100 202.100 161.800 ;
        RECT 205.400 161.100 205.800 165.400 ;
        RECT 208.700 165.200 209.000 166.800 ;
        RECT 212.300 166.700 212.700 166.800 ;
        RECT 211.800 166.200 212.200 166.300 ;
        RECT 213.100 166.200 213.500 166.300 ;
        RECT 211.000 165.900 213.500 166.200 ;
        RECT 215.800 166.100 216.200 169.900 ;
        RECT 218.500 168.000 218.900 169.500 ;
        RECT 220.600 168.500 221.000 169.500 ;
        RECT 218.100 167.700 218.900 168.000 ;
        RECT 218.100 167.500 218.500 167.700 ;
        RECT 218.100 167.200 218.400 167.500 ;
        RECT 220.700 167.400 221.000 168.500 ;
        RECT 223.300 168.000 223.700 169.500 ;
        RECT 225.400 168.500 225.800 169.500 ;
        RECT 216.600 167.100 217.000 167.200 ;
        RECT 217.400 167.100 218.400 167.200 ;
        RECT 216.600 166.800 218.400 167.100 ;
        RECT 218.900 167.100 221.000 167.400 ;
        RECT 222.900 167.700 223.700 168.000 ;
        RECT 222.900 167.500 223.300 167.700 ;
        RECT 222.900 167.200 223.200 167.500 ;
        RECT 225.500 167.400 225.800 168.500 ;
        RECT 228.100 168.000 228.500 169.500 ;
        RECT 230.200 168.500 230.600 169.500 ;
        RECT 218.900 166.900 219.400 167.100 ;
        RECT 217.400 166.100 217.800 166.200 ;
        RECT 211.000 165.800 211.400 165.900 ;
        RECT 215.800 165.800 217.800 166.100 ;
        RECT 211.800 165.500 214.600 165.600 ;
        RECT 211.700 165.400 214.600 165.500 ;
        RECT 207.800 164.900 209.000 165.200 ;
        RECT 209.700 165.300 214.600 165.400 ;
        RECT 209.700 165.100 212.100 165.300 ;
        RECT 207.800 164.400 208.100 164.900 ;
        RECT 207.400 164.000 208.100 164.400 ;
        RECT 208.900 164.500 209.300 164.600 ;
        RECT 209.700 164.500 210.000 165.100 ;
        RECT 208.900 164.200 210.000 164.500 ;
        RECT 210.300 164.500 213.000 164.800 ;
        RECT 210.300 164.400 210.700 164.500 ;
        RECT 212.600 164.400 213.000 164.500 ;
        RECT 209.500 163.700 209.900 163.800 ;
        RECT 210.900 163.700 211.300 163.800 ;
        RECT 207.800 163.100 208.200 163.500 ;
        RECT 209.500 163.400 211.300 163.700 ;
        RECT 209.900 163.100 210.200 163.400 ;
        RECT 212.600 163.100 213.000 163.500 ;
        RECT 207.500 161.100 208.100 163.100 ;
        RECT 209.800 161.100 210.200 163.100 ;
        RECT 212.000 162.800 213.000 163.100 ;
        RECT 212.000 161.100 212.400 162.800 ;
        RECT 214.200 161.100 214.600 165.300 ;
        RECT 215.800 161.100 216.200 165.800 ;
        RECT 217.400 165.400 217.800 165.800 ;
        RECT 218.100 164.900 218.400 166.800 ;
        RECT 218.700 166.500 219.400 166.900 ;
        RECT 222.200 166.800 223.200 167.200 ;
        RECT 223.700 167.100 225.800 167.400 ;
        RECT 227.700 167.700 228.500 168.000 ;
        RECT 227.700 167.500 228.100 167.700 ;
        RECT 227.700 167.200 228.000 167.500 ;
        RECT 230.300 167.400 230.600 168.500 ;
        RECT 232.900 168.000 233.300 169.500 ;
        RECT 235.000 168.500 235.400 169.500 ;
        RECT 223.700 166.900 224.200 167.100 ;
        RECT 219.100 165.500 219.400 166.500 ;
        RECT 219.800 165.800 220.200 166.600 ;
        RECT 220.600 165.800 221.000 166.600 ;
        RECT 219.100 165.200 221.000 165.500 ;
        RECT 222.200 165.400 222.600 166.200 ;
        RECT 218.100 164.600 218.900 164.900 ;
        RECT 218.500 161.100 218.900 164.600 ;
        RECT 220.700 163.500 221.000 165.200 ;
        RECT 222.900 164.900 223.200 166.800 ;
        RECT 223.500 166.500 224.200 166.900 ;
        RECT 227.000 166.800 228.000 167.200 ;
        RECT 228.500 167.100 230.600 167.400 ;
        RECT 232.500 167.700 233.300 168.000 ;
        RECT 232.500 167.500 232.900 167.700 ;
        RECT 232.500 167.200 232.800 167.500 ;
        RECT 235.100 167.400 235.400 168.500 ;
        RECT 235.800 167.900 236.200 169.900 ;
        RECT 236.600 168.000 237.000 169.900 ;
        RECT 238.200 168.000 238.600 169.900 ;
        RECT 236.600 167.900 238.600 168.000 ;
        RECT 239.800 168.900 240.200 169.900 ;
        RECT 228.500 166.900 229.000 167.100 ;
        RECT 223.900 165.500 224.200 166.500 ;
        RECT 224.600 165.800 225.000 166.600 ;
        RECT 225.400 165.800 225.800 166.600 ;
        RECT 223.900 165.200 225.800 165.500 ;
        RECT 227.000 165.400 227.400 166.200 ;
        RECT 222.900 164.600 223.700 164.900 ;
        RECT 223.300 164.200 223.700 164.600 ;
        RECT 223.000 163.800 223.700 164.200 ;
        RECT 220.600 161.500 221.000 163.500 ;
        RECT 223.300 161.100 223.700 163.800 ;
        RECT 225.500 163.500 225.800 165.200 ;
        RECT 227.700 164.900 228.000 166.800 ;
        RECT 228.300 166.500 229.000 166.900 ;
        RECT 231.800 166.800 232.800 167.200 ;
        RECT 233.300 167.100 235.400 167.400 ;
        RECT 235.900 167.200 236.200 167.900 ;
        RECT 236.700 167.700 238.500 167.900 ;
        RECT 237.800 167.200 238.200 167.400 ;
        RECT 239.800 167.200 240.100 168.900 ;
        RECT 240.600 167.800 241.000 168.600 ;
        RECT 241.500 168.200 241.900 168.600 ;
        RECT 241.400 167.800 241.800 168.200 ;
        RECT 242.200 167.900 242.600 169.900 ;
        RECT 245.900 169.200 246.300 169.900 ;
        RECT 245.900 168.800 246.600 169.200 ;
        RECT 245.900 168.200 246.300 168.800 ;
        RECT 233.300 166.900 233.800 167.100 ;
        RECT 228.700 165.500 229.000 166.500 ;
        RECT 229.400 165.800 229.800 166.600 ;
        RECT 230.200 165.800 230.600 166.600 ;
        RECT 231.000 166.100 231.400 166.200 ;
        RECT 231.800 166.100 232.200 166.200 ;
        RECT 231.000 165.800 232.200 166.100 ;
        RECT 228.700 165.200 230.600 165.500 ;
        RECT 231.800 165.400 232.200 165.800 ;
        RECT 227.700 164.600 228.500 164.900 ;
        RECT 225.400 161.500 225.800 163.500 ;
        RECT 228.100 162.200 228.500 164.600 ;
        RECT 230.300 163.500 230.600 165.200 ;
        RECT 232.500 164.900 232.800 166.800 ;
        RECT 233.100 166.500 233.800 166.900 ;
        RECT 235.800 166.800 237.100 167.200 ;
        RECT 237.800 166.900 238.600 167.200 ;
        RECT 238.200 166.800 238.600 166.900 ;
        RECT 239.800 167.100 240.200 167.200 ;
        RECT 241.400 167.100 241.700 167.800 ;
        RECT 239.800 166.800 241.700 167.100 ;
        RECT 233.500 165.500 233.800 166.500 ;
        RECT 234.200 165.800 234.600 166.600 ;
        RECT 235.000 165.800 235.400 166.600 ;
        RECT 233.500 165.200 235.400 165.500 ;
        RECT 232.500 164.600 233.300 164.900 ;
        RECT 227.800 161.800 228.500 162.200 ;
        RECT 228.100 161.100 228.500 161.800 ;
        RECT 230.200 161.500 230.600 163.500 ;
        RECT 232.900 161.100 233.300 164.600 ;
        RECT 235.100 163.500 235.400 165.200 ;
        RECT 235.800 165.100 236.200 165.200 ;
        RECT 236.800 165.100 237.100 166.800 ;
        RECT 237.400 165.800 237.800 166.600 ;
        RECT 239.000 165.400 239.400 166.200 ;
        RECT 239.800 165.100 240.100 166.800 ;
        RECT 242.300 166.200 242.600 167.900 ;
        RECT 245.400 167.900 246.300 168.200 ;
        RECT 243.000 166.400 243.400 167.200 ;
        RECT 244.600 166.800 245.000 167.600 ;
        RECT 241.400 166.100 241.800 166.200 ;
        RECT 242.200 166.100 242.600 166.200 ;
        RECT 243.800 166.100 244.200 166.200 ;
        RECT 241.400 165.800 242.600 166.100 ;
        RECT 243.400 165.800 244.200 166.100 ;
        RECT 241.500 165.100 241.800 165.800 ;
        RECT 243.400 165.600 243.800 165.800 ;
        RECT 235.800 164.800 236.500 165.100 ;
        RECT 236.800 164.800 237.300 165.100 ;
        RECT 236.200 164.200 236.500 164.800 ;
        RECT 236.200 163.800 236.600 164.200 ;
        RECT 235.000 161.500 235.400 163.500 ;
        RECT 236.900 161.100 237.300 164.800 ;
        RECT 239.300 164.700 240.200 165.100 ;
        RECT 239.300 161.100 239.700 164.700 ;
        RECT 241.400 161.100 241.800 165.100 ;
        RECT 242.200 164.800 244.200 165.100 ;
        RECT 242.200 161.100 242.600 164.800 ;
        RECT 243.800 161.100 244.200 164.800 ;
        RECT 245.400 161.100 245.800 167.900 ;
        RECT 247.000 167.700 247.400 169.900 ;
        RECT 249.100 169.200 249.700 169.900 ;
        RECT 249.100 168.900 249.800 169.200 ;
        RECT 251.400 168.900 251.800 169.900 ;
        RECT 253.600 169.200 254.000 169.900 ;
        RECT 253.600 168.900 254.600 169.200 ;
        RECT 249.400 168.500 249.800 168.900 ;
        RECT 251.500 168.600 251.800 168.900 ;
        RECT 251.500 168.300 252.900 168.600 ;
        RECT 252.500 168.200 252.900 168.300 ;
        RECT 253.400 168.200 253.800 168.600 ;
        RECT 254.200 168.500 254.600 168.900 ;
        RECT 248.500 167.700 248.900 167.800 ;
        RECT 247.000 167.400 248.900 167.700 ;
        RECT 247.000 165.700 247.400 167.400 ;
        RECT 250.500 167.100 250.900 167.200 ;
        RECT 252.600 167.100 253.000 167.200 ;
        RECT 253.400 167.100 253.700 168.200 ;
        RECT 255.800 167.500 256.200 169.900 ;
        RECT 256.700 168.200 257.100 168.600 ;
        RECT 256.600 167.800 257.000 168.200 ;
        RECT 257.400 167.900 257.800 169.900 ;
        RECT 255.000 167.100 255.800 167.200 ;
        RECT 250.300 166.800 255.800 167.100 ;
        RECT 249.400 166.400 249.800 166.500 ;
        RECT 247.900 166.100 249.800 166.400 ;
        RECT 250.300 166.100 250.600 166.800 ;
        RECT 253.900 166.700 254.300 166.800 ;
        RECT 254.700 166.200 255.100 166.300 ;
        RECT 251.000 166.100 251.400 166.200 ;
        RECT 247.900 166.000 248.300 166.100 ;
        RECT 250.200 165.800 251.400 166.100 ;
        RECT 252.600 165.900 255.100 166.200 ;
        RECT 256.600 166.100 257.000 166.200 ;
        RECT 257.500 166.100 257.800 167.900 ;
        RECT 259.800 167.600 260.200 169.900 ;
        RECT 262.200 167.600 262.600 169.900 ;
        RECT 259.800 167.300 260.900 167.600 ;
        RECT 262.200 167.300 263.300 167.600 ;
        RECT 258.200 166.400 258.600 167.200 ;
        RECT 259.000 166.100 259.400 166.200 ;
        RECT 252.600 165.800 253.000 165.900 ;
        RECT 256.600 165.800 257.800 166.100 ;
        RECT 258.600 165.800 259.400 166.100 ;
        RECT 259.800 165.800 260.200 166.600 ;
        RECT 260.600 165.800 260.900 167.300 ;
        RECT 262.200 165.800 262.600 166.600 ;
        RECT 263.000 165.800 263.300 167.300 ;
        RECT 248.700 165.700 249.100 165.800 ;
        RECT 247.000 165.400 249.100 165.700 ;
        RECT 246.200 164.400 246.600 165.200 ;
        RECT 247.000 161.100 247.400 165.400 ;
        RECT 250.300 165.200 250.600 165.800 ;
        RECT 253.400 165.500 256.200 165.600 ;
        RECT 253.300 165.400 256.200 165.500 ;
        RECT 249.400 164.900 250.600 165.200 ;
        RECT 251.300 165.300 256.200 165.400 ;
        RECT 251.300 165.100 253.700 165.300 ;
        RECT 249.400 164.400 249.700 164.900 ;
        RECT 249.000 164.000 249.700 164.400 ;
        RECT 250.500 164.500 250.900 164.600 ;
        RECT 251.300 164.500 251.600 165.100 ;
        RECT 250.500 164.200 251.600 164.500 ;
        RECT 251.900 164.500 254.600 164.800 ;
        RECT 251.900 164.400 252.300 164.500 ;
        RECT 254.200 164.400 254.600 164.500 ;
        RECT 251.100 163.700 251.500 163.800 ;
        RECT 252.500 163.700 252.900 163.800 ;
        RECT 249.400 163.100 249.800 163.500 ;
        RECT 251.100 163.400 252.900 163.700 ;
        RECT 251.500 163.100 251.800 163.400 ;
        RECT 254.200 163.100 254.600 163.500 ;
        RECT 249.100 161.100 249.700 163.100 ;
        RECT 251.400 161.100 251.800 163.100 ;
        RECT 253.600 162.800 254.600 163.100 ;
        RECT 253.600 161.100 254.000 162.800 ;
        RECT 255.800 161.100 256.200 165.300 ;
        RECT 256.700 165.100 257.000 165.800 ;
        RECT 258.600 165.600 259.000 165.800 ;
        RECT 260.600 165.400 261.200 165.800 ;
        RECT 263.000 165.400 263.600 165.800 ;
        RECT 260.600 165.100 260.900 165.400 ;
        RECT 263.000 165.100 263.300 165.400 ;
        RECT 256.600 161.100 257.000 165.100 ;
        RECT 257.400 164.800 259.400 165.100 ;
        RECT 257.400 161.100 257.800 164.800 ;
        RECT 259.000 161.100 259.400 164.800 ;
        RECT 259.800 164.800 260.900 165.100 ;
        RECT 262.200 164.800 263.300 165.100 ;
        RECT 259.800 161.100 260.200 164.800 ;
        RECT 262.200 161.100 262.600 164.800 ;
        RECT 0.600 155.700 1.000 159.900 ;
        RECT 2.800 158.200 3.200 159.900 ;
        RECT 2.200 157.900 3.200 158.200 ;
        RECT 5.000 157.900 5.400 159.900 ;
        RECT 7.100 157.900 7.700 159.900 ;
        RECT 2.200 157.500 2.600 157.900 ;
        RECT 5.000 157.600 5.300 157.900 ;
        RECT 3.900 157.300 5.700 157.600 ;
        RECT 7.000 157.500 7.400 157.900 ;
        RECT 3.900 157.200 4.300 157.300 ;
        RECT 5.300 157.200 5.700 157.300 ;
        RECT 9.400 157.100 9.800 159.900 ;
        RECT 10.200 157.100 10.600 157.200 ;
        RECT 2.200 156.500 2.600 156.600 ;
        RECT 4.500 156.500 4.900 156.600 ;
        RECT 2.200 156.200 4.900 156.500 ;
        RECT 5.200 156.500 6.300 156.800 ;
        RECT 5.200 155.900 5.500 156.500 ;
        RECT 5.900 156.400 6.300 156.500 ;
        RECT 7.100 156.600 7.800 157.000 ;
        RECT 9.400 156.800 10.600 157.100 ;
        RECT 7.100 156.100 7.400 156.600 ;
        RECT 3.100 155.700 5.500 155.900 ;
        RECT 0.600 155.600 5.500 155.700 ;
        RECT 6.200 155.800 7.400 156.100 ;
        RECT 0.600 155.500 3.500 155.600 ;
        RECT 0.600 155.400 3.400 155.500 ;
        RECT 6.200 155.200 6.500 155.800 ;
        RECT 9.400 155.600 9.800 156.800 ;
        RECT 7.700 155.300 9.800 155.600 ;
        RECT 7.700 155.200 8.100 155.300 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 1.700 154.800 4.200 155.100 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 8.500 154.900 8.900 155.000 ;
        RECT 1.700 154.700 2.100 154.800 ;
        RECT 2.500 154.200 2.900 154.300 ;
        RECT 6.200 154.200 6.500 154.800 ;
        RECT 7.000 154.600 8.900 154.900 ;
        RECT 7.000 154.500 7.400 154.600 ;
        RECT 1.000 153.900 6.500 154.200 ;
        RECT 1.000 153.800 1.800 153.900 ;
        RECT 0.600 151.100 1.000 153.500 ;
        RECT 3.100 152.800 3.400 153.900 ;
        RECT 5.900 153.800 6.300 153.900 ;
        RECT 9.400 153.600 9.800 155.300 ;
        RECT 7.900 153.300 9.800 153.600 ;
        RECT 10.200 153.400 10.600 154.200 ;
        RECT 7.900 153.200 8.300 153.300 ;
        RECT 2.200 152.100 2.600 152.500 ;
        RECT 3.000 152.400 3.400 152.800 ;
        RECT 3.900 152.700 4.300 152.800 ;
        RECT 3.900 152.400 5.300 152.700 ;
        RECT 5.000 152.100 5.300 152.400 ;
        RECT 7.000 152.100 7.400 152.500 ;
        RECT 2.200 151.800 3.200 152.100 ;
        RECT 2.800 151.100 3.200 151.800 ;
        RECT 5.000 151.100 5.400 152.100 ;
        RECT 7.000 151.800 7.700 152.100 ;
        RECT 7.100 151.100 7.700 151.800 ;
        RECT 9.400 151.100 9.800 153.300 ;
        RECT 11.000 153.100 11.400 159.900 ;
        RECT 11.800 155.800 12.200 156.600 ;
        RECT 13.400 155.600 13.800 159.900 ;
        RECT 15.000 155.600 15.400 159.900 ;
        RECT 16.600 155.600 17.000 159.900 ;
        RECT 18.200 155.600 18.600 159.900 ;
        RECT 19.800 155.700 20.200 159.900 ;
        RECT 22.000 158.200 22.400 159.900 ;
        RECT 21.400 157.900 22.400 158.200 ;
        RECT 24.200 157.900 24.600 159.900 ;
        RECT 26.300 157.900 26.900 159.900 ;
        RECT 21.400 157.500 21.800 157.900 ;
        RECT 24.200 157.600 24.500 157.900 ;
        RECT 23.100 157.300 24.900 157.600 ;
        RECT 26.200 157.500 26.600 157.900 ;
        RECT 23.100 157.200 23.500 157.300 ;
        RECT 24.500 157.200 24.900 157.300 ;
        RECT 21.400 156.500 21.800 156.600 ;
        RECT 23.700 156.500 24.100 156.600 ;
        RECT 21.400 156.200 24.100 156.500 ;
        RECT 24.400 156.500 25.500 156.800 ;
        RECT 24.400 155.900 24.700 156.500 ;
        RECT 25.100 156.400 25.500 156.500 ;
        RECT 26.300 156.600 27.000 157.000 ;
        RECT 26.300 156.100 26.600 156.600 ;
        RECT 22.300 155.700 24.700 155.900 ;
        RECT 19.800 155.600 24.700 155.700 ;
        RECT 25.400 155.800 26.600 156.100 ;
        RECT 13.400 155.200 14.300 155.600 ;
        RECT 15.000 155.200 16.100 155.600 ;
        RECT 16.600 155.200 17.700 155.600 ;
        RECT 18.200 155.200 19.400 155.600 ;
        RECT 19.800 155.500 22.700 155.600 ;
        RECT 19.800 155.400 22.600 155.500 ;
        RECT 25.400 155.200 25.700 155.800 ;
        RECT 28.600 155.600 29.000 159.900 ;
        RECT 26.900 155.300 29.000 155.600 ;
        RECT 29.400 155.700 29.800 159.900 ;
        RECT 31.600 158.200 32.000 159.900 ;
        RECT 31.000 157.900 32.000 158.200 ;
        RECT 33.800 157.900 34.200 159.900 ;
        RECT 35.900 157.900 36.500 159.900 ;
        RECT 31.000 157.500 31.400 157.900 ;
        RECT 33.800 157.600 34.100 157.900 ;
        RECT 32.700 157.300 34.500 157.600 ;
        RECT 35.800 157.500 36.200 157.900 ;
        RECT 32.700 157.200 33.100 157.300 ;
        RECT 34.100 157.200 34.500 157.300 ;
        RECT 31.000 156.500 31.400 156.600 ;
        RECT 33.300 156.500 33.700 156.600 ;
        RECT 31.000 156.200 33.700 156.500 ;
        RECT 34.000 156.500 35.100 156.800 ;
        RECT 34.000 155.900 34.300 156.500 ;
        RECT 34.700 156.400 35.100 156.500 ;
        RECT 35.900 156.600 36.600 157.000 ;
        RECT 35.900 156.100 36.200 156.600 ;
        RECT 31.900 155.700 34.300 155.900 ;
        RECT 29.400 155.600 34.300 155.700 ;
        RECT 35.000 155.800 36.200 156.100 ;
        RECT 29.400 155.500 32.300 155.600 ;
        RECT 29.400 155.400 32.200 155.500 ;
        RECT 26.900 155.200 27.300 155.300 ;
        RECT 13.900 154.500 14.300 155.200 ;
        RECT 15.700 154.500 16.100 155.200 ;
        RECT 17.300 154.500 17.700 155.200 ;
        RECT 12.600 154.100 13.500 154.500 ;
        RECT 13.900 154.100 15.200 154.500 ;
        RECT 15.700 154.100 16.900 154.500 ;
        RECT 17.300 154.100 18.600 154.500 ;
        RECT 12.600 153.800 13.000 154.100 ;
        RECT 13.900 153.800 14.300 154.100 ;
        RECT 15.700 153.800 16.100 154.100 ;
        RECT 17.300 153.800 17.700 154.100 ;
        RECT 19.000 153.800 19.400 155.200 ;
        RECT 23.000 155.100 23.400 155.200 ;
        RECT 20.900 154.800 23.400 155.100 ;
        RECT 25.400 154.800 25.800 155.200 ;
        RECT 27.700 154.900 28.100 155.000 ;
        RECT 20.900 154.700 21.300 154.800 ;
        RECT 21.700 154.200 22.100 154.300 ;
        RECT 25.400 154.200 25.700 154.800 ;
        RECT 26.200 154.600 28.100 154.900 ;
        RECT 26.200 154.500 26.600 154.600 ;
        RECT 20.200 153.900 25.700 154.200 ;
        RECT 20.200 153.800 21.000 153.900 ;
        RECT 13.400 153.400 14.300 153.800 ;
        RECT 15.000 153.400 16.100 153.800 ;
        RECT 16.600 153.400 17.700 153.800 ;
        RECT 18.200 153.400 19.400 153.800 ;
        RECT 11.000 152.800 11.900 153.100 ;
        RECT 11.500 152.200 11.900 152.800 ;
        RECT 11.000 151.800 11.900 152.200 ;
        RECT 11.500 151.100 11.900 151.800 ;
        RECT 13.400 151.100 13.800 153.400 ;
        RECT 15.000 151.100 15.400 153.400 ;
        RECT 16.600 151.100 17.000 153.400 ;
        RECT 18.200 151.100 18.600 153.400 ;
        RECT 19.800 151.100 20.200 153.500 ;
        RECT 22.300 152.800 22.600 153.900 ;
        RECT 25.100 153.800 25.500 153.900 ;
        RECT 28.600 153.600 29.000 155.300 ;
        RECT 32.600 155.100 33.000 155.200 ;
        RECT 30.500 154.800 33.000 155.100 ;
        RECT 30.500 154.700 30.900 154.800 ;
        RECT 31.300 154.200 31.700 154.300 ;
        RECT 35.000 154.200 35.300 155.800 ;
        RECT 38.200 155.600 38.600 159.900 ;
        RECT 40.300 156.300 40.700 159.900 ;
        RECT 39.800 155.900 40.700 156.300 ;
        RECT 41.400 155.900 41.800 159.900 ;
        RECT 42.200 156.200 42.600 159.900 ;
        RECT 43.800 156.200 44.200 159.900 ;
        RECT 45.400 156.400 45.800 159.900 ;
        RECT 42.200 155.900 44.200 156.200 ;
        RECT 36.500 155.300 38.600 155.600 ;
        RECT 36.500 155.200 36.900 155.300 ;
        RECT 37.300 154.900 37.700 155.000 ;
        RECT 35.800 154.600 37.700 154.900 ;
        RECT 35.800 154.500 36.200 154.600 ;
        RECT 29.800 153.900 35.300 154.200 ;
        RECT 29.800 153.800 30.600 153.900 ;
        RECT 27.100 153.300 29.000 153.600 ;
        RECT 27.100 153.200 27.500 153.300 ;
        RECT 21.400 152.100 21.800 152.500 ;
        RECT 22.200 152.400 22.600 152.800 ;
        RECT 23.100 152.700 23.500 152.800 ;
        RECT 23.100 152.400 24.500 152.700 ;
        RECT 24.200 152.100 24.500 152.400 ;
        RECT 26.200 152.100 26.600 152.500 ;
        RECT 21.400 151.800 22.400 152.100 ;
        RECT 22.000 151.100 22.400 151.800 ;
        RECT 24.200 151.100 24.600 152.100 ;
        RECT 26.200 151.800 26.900 152.100 ;
        RECT 26.300 151.100 26.900 151.800 ;
        RECT 28.600 151.100 29.000 153.300 ;
        RECT 29.400 151.100 29.800 153.500 ;
        RECT 31.900 152.800 32.200 153.900 ;
        RECT 34.700 153.800 35.100 153.900 ;
        RECT 38.200 153.600 38.600 155.300 ;
        RECT 39.900 154.200 40.200 155.900 ;
        RECT 40.600 154.800 41.000 155.600 ;
        RECT 41.500 155.200 41.800 155.900 ;
        RECT 45.300 155.800 45.800 156.400 ;
        RECT 47.000 156.200 47.400 159.900 ;
        RECT 46.100 155.900 47.400 156.200 ;
        RECT 47.800 157.500 48.200 159.500 ;
        RECT 43.400 155.200 43.800 155.400 ;
        RECT 41.400 154.900 42.600 155.200 ;
        RECT 43.400 154.900 44.200 155.200 ;
        RECT 41.400 154.800 41.800 154.900 ;
        RECT 39.800 153.800 40.200 154.200 ;
        RECT 36.700 153.300 38.600 153.600 ;
        RECT 36.700 153.200 37.100 153.300 ;
        RECT 31.000 152.100 31.400 152.500 ;
        RECT 31.800 152.400 32.200 152.800 ;
        RECT 32.700 152.700 33.100 152.800 ;
        RECT 32.700 152.400 34.100 152.700 ;
        RECT 33.800 152.100 34.100 152.400 ;
        RECT 35.800 152.100 36.200 152.500 ;
        RECT 31.000 151.800 32.000 152.100 ;
        RECT 31.600 151.100 32.000 151.800 ;
        RECT 33.800 151.100 34.200 152.100 ;
        RECT 35.800 151.800 36.500 152.100 ;
        RECT 35.900 151.100 36.500 151.800 ;
        RECT 38.200 151.100 38.600 153.300 ;
        RECT 39.000 152.400 39.400 153.200 ;
        RECT 39.900 153.100 40.200 153.800 ;
        RECT 42.300 153.200 42.600 154.900 ;
        RECT 43.800 154.800 44.200 154.900 ;
        RECT 43.000 153.800 43.400 154.600 ;
        RECT 43.800 154.100 44.100 154.800 ;
        RECT 45.300 154.200 45.600 155.800 ;
        RECT 46.100 154.900 46.400 155.900 ;
        RECT 47.800 155.800 48.100 157.500 ;
        RECT 49.900 156.400 50.300 159.900 ;
        RECT 49.900 156.100 50.700 156.400 ;
        RECT 47.800 155.500 49.700 155.800 ;
        RECT 45.900 154.500 46.400 154.900 ;
        RECT 45.300 154.100 45.800 154.200 ;
        RECT 43.800 153.800 45.800 154.100 ;
        RECT 41.400 153.100 41.800 153.200 ;
        RECT 39.800 152.800 41.800 153.100 ;
        RECT 39.900 152.100 40.200 152.800 ;
        RECT 41.500 152.400 41.900 152.800 ;
        RECT 39.800 151.100 40.200 152.100 ;
        RECT 42.200 151.100 42.600 153.200 ;
        RECT 45.300 153.100 45.600 153.800 ;
        RECT 46.100 153.700 46.400 154.500 ;
        RECT 46.900 154.800 47.400 155.200 ;
        RECT 46.900 154.400 47.300 154.800 ;
        RECT 47.800 154.400 48.200 155.200 ;
        RECT 48.600 154.400 49.000 155.200 ;
        RECT 49.400 154.500 49.700 155.500 ;
        RECT 49.400 154.100 50.100 154.500 ;
        RECT 50.400 154.200 50.700 156.100 ;
        RECT 51.000 155.100 51.400 155.600 ;
        RECT 52.600 155.100 53.000 159.900 ;
        RECT 55.800 155.700 56.200 159.900 ;
        RECT 58.000 158.200 58.400 159.900 ;
        RECT 57.400 157.900 58.400 158.200 ;
        RECT 60.200 157.900 60.600 159.900 ;
        RECT 62.300 157.900 62.900 159.900 ;
        RECT 57.400 157.500 57.800 157.900 ;
        RECT 60.200 157.600 60.500 157.900 ;
        RECT 59.100 157.300 60.900 157.600 ;
        RECT 62.200 157.500 62.600 157.900 ;
        RECT 59.100 157.200 59.500 157.300 ;
        RECT 60.500 157.200 60.900 157.300 ;
        RECT 57.400 156.500 57.800 156.600 ;
        RECT 59.700 156.500 60.100 156.600 ;
        RECT 57.400 156.200 60.100 156.500 ;
        RECT 60.400 156.500 61.500 156.800 ;
        RECT 60.400 155.900 60.700 156.500 ;
        RECT 61.100 156.400 61.500 156.500 ;
        RECT 62.300 156.600 63.000 157.000 ;
        RECT 62.300 156.100 62.600 156.600 ;
        RECT 58.300 155.700 60.700 155.900 ;
        RECT 55.800 155.600 60.700 155.700 ;
        RECT 61.400 155.800 62.600 156.100 ;
        RECT 55.800 155.500 58.700 155.600 ;
        RECT 55.800 155.400 58.600 155.500 ;
        RECT 59.000 155.100 59.400 155.200 ;
        RECT 51.000 154.800 53.000 155.100 ;
        RECT 49.400 153.900 49.900 154.100 ;
        RECT 46.100 153.400 47.400 153.700 ;
        RECT 45.300 152.800 45.800 153.100 ;
        RECT 45.400 151.100 45.800 152.800 ;
        RECT 47.000 151.100 47.400 153.400 ;
        RECT 47.800 153.600 49.900 153.900 ;
        RECT 50.400 153.800 51.400 154.200 ;
        RECT 47.800 152.500 48.100 153.600 ;
        RECT 50.400 153.500 50.700 153.800 ;
        RECT 50.300 153.300 50.700 153.500 ;
        RECT 49.900 153.000 50.700 153.300 ;
        RECT 47.800 151.500 48.200 152.500 ;
        RECT 49.900 151.500 50.300 153.000 ;
        RECT 52.600 151.100 53.000 154.800 ;
        RECT 56.900 154.800 59.400 155.100 ;
        RECT 56.900 154.700 57.300 154.800 ;
        RECT 58.200 154.700 58.600 154.800 ;
        RECT 57.700 154.200 58.100 154.300 ;
        RECT 61.400 154.200 61.700 155.800 ;
        RECT 64.600 155.600 65.000 159.900 ;
        RECT 62.900 155.300 65.000 155.600 ;
        RECT 65.400 155.700 65.800 159.900 ;
        RECT 67.600 158.200 68.000 159.900 ;
        RECT 67.000 157.900 68.000 158.200 ;
        RECT 69.800 157.900 70.200 159.900 ;
        RECT 71.900 157.900 72.500 159.900 ;
        RECT 67.000 157.500 67.400 157.900 ;
        RECT 69.800 157.600 70.100 157.900 ;
        RECT 68.700 157.300 70.500 157.600 ;
        RECT 71.800 157.500 72.200 157.900 ;
        RECT 68.700 157.200 69.100 157.300 ;
        RECT 70.100 157.200 70.500 157.300 ;
        RECT 67.000 156.500 67.400 156.600 ;
        RECT 69.300 156.500 69.700 156.600 ;
        RECT 67.000 156.200 69.700 156.500 ;
        RECT 70.000 156.500 71.100 156.800 ;
        RECT 70.000 155.900 70.300 156.500 ;
        RECT 70.700 156.400 71.100 156.500 ;
        RECT 71.900 156.600 72.600 157.000 ;
        RECT 71.900 156.100 72.200 156.600 ;
        RECT 67.900 155.700 70.300 155.900 ;
        RECT 65.400 155.600 70.300 155.700 ;
        RECT 71.000 155.800 72.200 156.100 ;
        RECT 65.400 155.500 68.300 155.600 ;
        RECT 65.400 155.400 68.200 155.500 ;
        RECT 62.900 155.200 63.300 155.300 ;
        RECT 63.700 154.900 64.100 155.000 ;
        RECT 62.200 154.600 64.100 154.900 ;
        RECT 62.200 154.500 62.600 154.600 ;
        RECT 56.200 153.900 61.700 154.200 ;
        RECT 56.200 153.800 57.000 153.900 ;
        RECT 53.400 152.400 53.800 153.200 ;
        RECT 55.800 151.100 56.200 153.500 ;
        RECT 58.300 152.800 58.600 153.900 ;
        RECT 61.100 153.800 61.500 153.900 ;
        RECT 64.600 153.600 65.000 155.300 ;
        RECT 68.600 155.100 69.000 155.200 ;
        RECT 66.500 154.800 69.000 155.100 ;
        RECT 66.500 154.700 66.900 154.800 ;
        RECT 67.300 154.200 67.700 154.300 ;
        RECT 71.000 154.200 71.300 155.800 ;
        RECT 74.200 155.600 74.600 159.900 ;
        RECT 76.900 159.200 77.300 159.900 ;
        RECT 76.600 158.800 77.300 159.200 ;
        RECT 76.900 156.400 77.300 158.800 ;
        RECT 79.000 157.500 79.400 159.500 ;
        RECT 76.500 156.100 77.300 156.400 ;
        RECT 72.500 155.300 74.600 155.600 ;
        RECT 72.500 155.200 72.900 155.300 ;
        RECT 73.300 154.900 73.700 155.000 ;
        RECT 71.800 154.600 73.700 154.900 ;
        RECT 71.800 154.500 72.200 154.600 ;
        RECT 65.800 153.900 71.300 154.200 ;
        RECT 65.800 153.800 66.600 153.900 ;
        RECT 63.100 153.300 65.000 153.600 ;
        RECT 63.100 153.200 63.500 153.300 ;
        RECT 57.400 152.100 57.800 152.500 ;
        RECT 58.200 152.400 58.600 152.800 ;
        RECT 59.100 152.700 59.500 152.800 ;
        RECT 59.100 152.400 60.500 152.700 ;
        RECT 60.200 152.100 60.500 152.400 ;
        RECT 62.200 152.100 62.600 152.500 ;
        RECT 57.400 151.800 58.400 152.100 ;
        RECT 58.000 151.100 58.400 151.800 ;
        RECT 60.200 151.100 60.600 152.100 ;
        RECT 62.200 151.800 62.900 152.100 ;
        RECT 62.300 151.100 62.900 151.800 ;
        RECT 64.600 151.100 65.000 153.300 ;
        RECT 65.400 151.100 65.800 153.500 ;
        RECT 67.900 152.800 68.200 153.900 ;
        RECT 70.700 153.800 71.100 153.900 ;
        RECT 74.200 153.600 74.600 155.300 ;
        RECT 75.800 155.100 76.200 155.600 ;
        RECT 75.000 154.800 76.200 155.100 ;
        RECT 75.000 154.200 75.300 154.800 ;
        RECT 76.500 154.200 76.800 156.100 ;
        RECT 79.100 155.800 79.400 157.500 ;
        RECT 77.500 155.500 79.400 155.800 ;
        RECT 77.500 154.500 77.800 155.500 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 75.800 153.800 76.800 154.200 ;
        RECT 77.100 154.100 77.800 154.500 ;
        RECT 78.200 154.400 78.600 155.200 ;
        RECT 79.000 154.400 79.400 155.200 ;
        RECT 79.800 154.800 80.200 155.200 ;
        RECT 80.600 155.100 81.000 159.900 ;
        RECT 82.600 156.800 83.000 157.200 ;
        RECT 81.400 155.800 81.800 156.600 ;
        RECT 82.600 156.200 82.900 156.800 ;
        RECT 83.300 156.200 83.700 159.900 ;
        RECT 87.300 157.200 87.700 159.900 ;
        RECT 89.400 157.500 89.800 159.500 ;
        RECT 87.300 156.800 88.200 157.200 ;
        RECT 87.300 156.400 87.700 156.800 ;
        RECT 82.200 155.900 82.900 156.200 ;
        RECT 83.200 155.900 83.700 156.200 ;
        RECT 86.900 156.100 87.700 156.400 ;
        RECT 82.200 155.800 82.600 155.900 ;
        RECT 82.200 155.100 82.500 155.800 ;
        RECT 80.600 154.800 82.500 155.100 ;
        RECT 72.700 153.300 74.600 153.600 ;
        RECT 72.700 153.200 73.100 153.300 ;
        RECT 67.000 152.100 67.400 152.500 ;
        RECT 67.800 152.400 68.200 152.800 ;
        RECT 68.700 152.700 69.100 152.800 ;
        RECT 68.700 152.400 70.100 152.700 ;
        RECT 69.800 152.100 70.100 152.400 ;
        RECT 71.800 152.100 72.200 152.500 ;
        RECT 67.000 151.800 68.000 152.100 ;
        RECT 67.600 151.100 68.000 151.800 ;
        RECT 69.800 151.100 70.200 152.100 ;
        RECT 71.800 151.800 72.500 152.100 ;
        RECT 71.900 151.100 72.500 151.800 ;
        RECT 74.200 151.100 74.600 153.300 ;
        RECT 76.500 153.500 76.800 153.800 ;
        RECT 77.300 153.900 77.800 154.100 ;
        RECT 79.800 154.200 80.100 154.800 ;
        RECT 77.300 153.600 79.400 153.900 ;
        RECT 76.500 153.300 76.900 153.500 ;
        RECT 76.500 153.000 77.300 153.300 ;
        RECT 76.900 151.500 77.300 153.000 ;
        RECT 79.100 152.500 79.400 153.600 ;
        RECT 79.800 153.400 80.200 154.200 ;
        RECT 80.600 153.100 81.000 154.800 ;
        RECT 83.200 154.200 83.500 155.900 ;
        RECT 83.800 154.400 84.200 155.200 ;
        RECT 86.200 154.800 86.600 155.600 ;
        RECT 86.900 154.200 87.200 156.100 ;
        RECT 89.500 155.800 89.800 157.500 ;
        RECT 87.900 155.500 89.800 155.800 ;
        RECT 90.200 155.700 90.600 159.900 ;
        RECT 92.400 158.200 92.800 159.900 ;
        RECT 91.800 157.900 92.800 158.200 ;
        RECT 94.600 157.900 95.000 159.900 ;
        RECT 96.700 157.900 97.300 159.900 ;
        RECT 91.800 157.500 92.200 157.900 ;
        RECT 94.600 157.600 94.900 157.900 ;
        RECT 93.500 157.300 95.300 157.600 ;
        RECT 96.600 157.500 97.000 157.900 ;
        RECT 93.500 157.200 93.900 157.300 ;
        RECT 94.900 157.200 95.300 157.300 ;
        RECT 91.800 156.500 92.200 156.600 ;
        RECT 94.100 156.500 94.500 156.600 ;
        RECT 91.800 156.200 94.500 156.500 ;
        RECT 94.800 156.500 95.900 156.800 ;
        RECT 94.800 155.900 95.100 156.500 ;
        RECT 95.500 156.400 95.900 156.500 ;
        RECT 96.700 156.600 97.400 157.000 ;
        RECT 96.700 156.100 97.000 156.600 ;
        RECT 92.700 155.700 95.100 155.900 ;
        RECT 90.200 155.600 95.100 155.700 ;
        RECT 95.800 155.800 97.000 156.100 ;
        RECT 90.200 155.500 93.100 155.600 ;
        RECT 87.900 154.500 88.200 155.500 ;
        RECT 90.200 155.400 93.000 155.500 ;
        RECT 82.200 153.800 83.500 154.200 ;
        RECT 84.600 154.100 85.000 154.200 ;
        RECT 84.200 153.800 85.000 154.100 ;
        RECT 86.200 153.800 87.200 154.200 ;
        RECT 87.500 154.100 88.200 154.500 ;
        RECT 88.600 154.400 89.000 155.200 ;
        RECT 89.400 154.400 89.800 155.200 ;
        RECT 93.400 155.100 93.800 155.200 ;
        RECT 91.300 154.800 93.800 155.100 ;
        RECT 91.300 154.700 91.700 154.800 ;
        RECT 92.100 154.200 92.500 154.300 ;
        RECT 95.800 154.200 96.100 155.800 ;
        RECT 99.000 155.600 99.400 159.900 ;
        RECT 97.300 155.300 99.400 155.600 ;
        RECT 99.800 157.500 100.200 159.500 ;
        RECT 101.900 159.200 102.300 159.900 ;
        RECT 101.400 158.800 102.300 159.200 ;
        RECT 99.800 155.800 100.100 157.500 ;
        RECT 101.900 156.400 102.300 158.800 ;
        RECT 101.900 156.100 102.700 156.400 ;
        RECT 99.800 155.500 101.700 155.800 ;
        RECT 97.300 155.200 97.700 155.300 ;
        RECT 98.100 154.900 98.500 155.000 ;
        RECT 96.600 154.600 98.500 154.900 ;
        RECT 96.600 154.500 97.000 154.600 ;
        RECT 82.300 153.100 82.600 153.800 ;
        RECT 84.200 153.600 84.600 153.800 ;
        RECT 86.900 153.500 87.200 153.800 ;
        RECT 87.700 153.900 88.200 154.100 ;
        RECT 90.600 153.900 96.100 154.200 ;
        RECT 87.700 153.600 89.800 153.900 ;
        RECT 90.600 153.800 91.400 153.900 ;
        RECT 86.900 153.300 87.300 153.500 ;
        RECT 83.100 153.100 84.900 153.300 ;
        RECT 80.600 152.800 81.500 153.100 ;
        RECT 79.000 151.500 79.400 152.500 ;
        RECT 81.100 151.100 81.500 152.800 ;
        RECT 82.200 151.100 82.600 153.100 ;
        RECT 83.000 153.000 85.000 153.100 ;
        RECT 86.900 153.000 87.700 153.300 ;
        RECT 83.000 151.100 83.400 153.000 ;
        RECT 84.600 151.100 85.000 153.000 ;
        RECT 87.300 151.500 87.700 153.000 ;
        RECT 89.500 152.500 89.800 153.600 ;
        RECT 89.400 151.500 89.800 152.500 ;
        RECT 90.200 151.100 90.600 153.500 ;
        RECT 92.700 152.800 93.000 153.900 ;
        RECT 95.500 153.800 95.900 153.900 ;
        RECT 99.000 153.600 99.400 155.300 ;
        RECT 99.800 154.400 100.200 155.200 ;
        RECT 100.600 154.400 101.000 155.200 ;
        RECT 101.400 154.500 101.700 155.500 ;
        RECT 101.400 154.100 102.100 154.500 ;
        RECT 102.400 154.200 102.700 156.100 ;
        RECT 103.000 155.100 103.400 155.600 ;
        RECT 104.600 155.100 105.000 155.200 ;
        RECT 103.000 154.800 105.000 155.100 ;
        RECT 105.400 155.100 105.800 159.900 ;
        RECT 109.000 156.800 109.400 157.200 ;
        RECT 106.200 155.800 106.600 156.600 ;
        RECT 109.000 156.200 109.300 156.800 ;
        RECT 109.700 156.200 110.100 159.900 ;
        RECT 108.600 155.900 109.300 156.200 ;
        RECT 109.600 155.900 110.100 156.200 ;
        RECT 108.600 155.800 109.000 155.900 ;
        RECT 108.600 155.100 108.900 155.800 ;
        RECT 105.400 154.800 108.900 155.100 ;
        RECT 101.400 153.900 101.900 154.100 ;
        RECT 97.500 153.300 99.400 153.600 ;
        RECT 97.500 153.200 97.900 153.300 ;
        RECT 91.800 152.100 92.200 152.500 ;
        RECT 92.600 152.400 93.000 152.800 ;
        RECT 93.500 152.700 93.900 152.800 ;
        RECT 93.500 152.400 94.900 152.700 ;
        RECT 94.600 152.100 94.900 152.400 ;
        RECT 96.600 152.100 97.000 152.500 ;
        RECT 91.800 151.800 92.800 152.100 ;
        RECT 92.400 151.100 92.800 151.800 ;
        RECT 94.600 151.100 95.000 152.100 ;
        RECT 96.600 151.800 97.300 152.100 ;
        RECT 96.700 151.100 97.300 151.800 ;
        RECT 99.000 151.100 99.400 153.300 ;
        RECT 99.800 153.600 101.900 153.900 ;
        RECT 102.400 153.800 103.400 154.200 ;
        RECT 103.800 154.100 104.200 154.200 ;
        RECT 104.600 154.100 105.000 154.200 ;
        RECT 103.800 153.800 105.000 154.100 ;
        RECT 99.800 152.500 100.100 153.600 ;
        RECT 102.400 153.500 102.700 153.800 ;
        RECT 102.300 153.300 102.700 153.500 ;
        RECT 104.600 153.400 105.000 153.800 ;
        RECT 101.900 153.000 102.700 153.300 ;
        RECT 105.400 153.100 105.800 154.800 ;
        RECT 109.600 154.200 109.900 155.900 ;
        RECT 110.200 154.400 110.600 155.200 ;
        RECT 107.000 154.100 107.400 154.200 ;
        RECT 108.600 154.100 109.900 154.200 ;
        RECT 111.000 154.100 111.400 154.200 ;
        RECT 107.000 153.800 109.900 154.100 ;
        RECT 110.600 153.800 111.400 154.100 ;
        RECT 108.700 153.100 109.000 153.800 ;
        RECT 110.600 153.600 111.000 153.800 ;
        RECT 111.800 153.400 112.200 154.200 ;
        RECT 109.500 153.100 111.300 153.300 ;
        RECT 112.600 153.100 113.000 159.900 ;
        RECT 113.400 155.800 113.800 156.600 ;
        RECT 115.500 156.300 115.900 159.900 ;
        RECT 115.000 155.900 115.900 156.300 ;
        RECT 115.100 154.200 115.400 155.900 ;
        RECT 116.600 155.700 117.000 159.900 ;
        RECT 118.800 158.200 119.200 159.900 ;
        RECT 118.200 157.900 119.200 158.200 ;
        RECT 121.000 157.900 121.400 159.900 ;
        RECT 123.100 157.900 123.700 159.900 ;
        RECT 118.200 157.500 118.600 157.900 ;
        RECT 121.000 157.600 121.300 157.900 ;
        RECT 119.900 157.300 121.700 157.600 ;
        RECT 123.000 157.500 123.400 157.900 ;
        RECT 119.900 157.200 120.300 157.300 ;
        RECT 121.300 157.200 121.700 157.300 ;
        RECT 118.200 156.500 118.600 156.600 ;
        RECT 120.500 156.500 120.900 156.600 ;
        RECT 118.200 156.200 120.900 156.500 ;
        RECT 121.200 156.500 122.300 156.800 ;
        RECT 121.200 155.900 121.500 156.500 ;
        RECT 121.900 156.400 122.300 156.500 ;
        RECT 123.100 156.600 123.800 157.000 ;
        RECT 123.100 156.100 123.400 156.600 ;
        RECT 119.100 155.700 121.500 155.900 ;
        RECT 116.600 155.600 121.500 155.700 ;
        RECT 122.200 155.800 123.400 156.100 ;
        RECT 115.800 154.800 116.200 155.600 ;
        RECT 116.600 155.500 119.500 155.600 ;
        RECT 116.600 155.400 119.400 155.500 ;
        RECT 119.800 155.100 120.200 155.200 ;
        RECT 120.600 155.100 121.000 155.200 ;
        RECT 117.700 154.800 121.000 155.100 ;
        RECT 117.700 154.700 118.100 154.800 ;
        RECT 118.500 154.200 118.900 154.300 ;
        RECT 122.200 154.200 122.500 155.800 ;
        RECT 125.400 155.600 125.800 159.900 ;
        RECT 127.500 157.200 127.900 159.900 ;
        RECT 127.000 156.800 127.900 157.200 ;
        RECT 128.200 156.800 128.600 157.200 ;
        RECT 129.400 156.800 130.200 157.200 ;
        RECT 127.500 156.200 127.900 156.800 ;
        RECT 128.300 156.200 128.600 156.800 ;
        RECT 129.800 156.200 130.100 156.800 ;
        RECT 130.500 156.200 130.900 159.900 ;
        RECT 127.500 155.900 128.000 156.200 ;
        RECT 128.300 155.900 129.000 156.200 ;
        RECT 123.700 155.300 125.800 155.600 ;
        RECT 123.700 155.200 124.100 155.300 ;
        RECT 124.500 154.900 124.900 155.000 ;
        RECT 123.000 154.600 124.900 154.900 ;
        RECT 123.000 154.500 123.400 154.600 ;
        RECT 115.000 153.800 115.400 154.200 ;
        RECT 117.000 153.900 122.600 154.200 ;
        RECT 117.000 153.800 117.800 153.900 ;
        RECT 99.800 151.500 100.200 152.500 ;
        RECT 101.900 151.500 102.300 153.000 ;
        RECT 105.400 152.800 106.300 153.100 ;
        RECT 105.900 151.100 106.300 152.800 ;
        RECT 108.600 151.100 109.000 153.100 ;
        RECT 109.400 153.000 111.400 153.100 ;
        RECT 109.400 151.100 109.800 153.000 ;
        RECT 111.000 151.100 111.400 153.000 ;
        RECT 112.600 152.800 113.500 153.100 ;
        RECT 113.100 152.200 113.500 152.800 ;
        RECT 114.200 152.400 114.600 153.200 ;
        RECT 115.100 152.200 115.400 153.800 ;
        RECT 112.600 151.800 113.500 152.200 ;
        RECT 113.100 151.100 113.500 151.800 ;
        RECT 115.000 151.100 115.400 152.200 ;
        RECT 116.600 151.100 117.000 153.500 ;
        RECT 119.100 152.800 119.400 153.900 ;
        RECT 121.900 153.800 122.600 153.900 ;
        RECT 125.400 153.600 125.800 155.300 ;
        RECT 127.000 154.400 127.400 155.200 ;
        RECT 127.700 154.200 128.000 155.900 ;
        RECT 128.600 155.800 129.000 155.900 ;
        RECT 129.400 155.900 130.100 156.200 ;
        RECT 130.400 155.900 130.900 156.200 ;
        RECT 129.400 155.800 129.800 155.900 ;
        RECT 128.600 155.100 128.900 155.800 ;
        RECT 130.400 155.100 130.700 155.900 ;
        RECT 132.600 155.700 133.000 159.900 ;
        RECT 134.800 158.200 135.200 159.900 ;
        RECT 134.200 157.900 135.200 158.200 ;
        RECT 137.000 157.900 137.400 159.900 ;
        RECT 139.100 157.900 139.700 159.900 ;
        RECT 134.200 157.500 134.600 157.900 ;
        RECT 137.000 157.600 137.300 157.900 ;
        RECT 135.900 157.300 137.700 157.600 ;
        RECT 139.000 157.500 139.400 157.900 ;
        RECT 135.900 157.200 136.300 157.300 ;
        RECT 137.300 157.200 137.700 157.300 ;
        RECT 134.200 156.500 134.600 156.600 ;
        RECT 136.500 156.500 136.900 156.600 ;
        RECT 134.200 156.200 136.900 156.500 ;
        RECT 137.200 156.500 138.300 156.800 ;
        RECT 137.200 155.900 137.500 156.500 ;
        RECT 137.900 156.400 138.300 156.500 ;
        RECT 139.100 156.600 139.800 157.000 ;
        RECT 139.100 156.100 139.400 156.600 ;
        RECT 135.100 155.700 137.500 155.900 ;
        RECT 132.600 155.600 137.500 155.700 ;
        RECT 138.200 155.800 139.400 156.100 ;
        RECT 132.600 155.500 135.500 155.600 ;
        RECT 132.600 155.400 135.400 155.500 ;
        RECT 128.600 154.800 130.700 155.100 ;
        RECT 130.400 154.200 130.700 154.800 ;
        RECT 131.000 154.400 131.400 155.200 ;
        RECT 135.800 155.100 136.200 155.200 ;
        RECT 133.700 154.800 136.200 155.100 ;
        RECT 133.700 154.700 134.100 154.800 ;
        RECT 134.500 154.200 134.900 154.300 ;
        RECT 138.200 154.200 138.500 155.800 ;
        RECT 141.400 155.600 141.800 159.900 ;
        RECT 142.200 155.800 142.600 156.600 ;
        RECT 139.700 155.300 141.800 155.600 ;
        RECT 139.700 155.200 140.100 155.300 ;
        RECT 140.500 154.900 140.900 155.000 ;
        RECT 139.000 154.600 140.900 154.900 ;
        RECT 139.000 154.500 139.400 154.600 ;
        RECT 126.200 154.100 126.600 154.200 ;
        RECT 126.200 153.800 127.000 154.100 ;
        RECT 127.700 153.800 129.000 154.200 ;
        RECT 129.400 153.800 130.700 154.200 ;
        RECT 131.800 154.100 132.200 154.200 ;
        RECT 131.400 153.800 132.200 154.100 ;
        RECT 133.000 153.900 138.500 154.200 ;
        RECT 133.000 153.800 133.800 153.900 ;
        RECT 126.600 153.600 127.000 153.800 ;
        RECT 123.900 153.300 125.800 153.600 ;
        RECT 123.900 153.200 124.300 153.300 ;
        RECT 118.200 152.100 118.600 152.500 ;
        RECT 119.000 152.400 119.400 152.800 ;
        RECT 119.900 152.700 120.300 152.800 ;
        RECT 119.900 152.400 121.300 152.700 ;
        RECT 121.000 152.100 121.300 152.400 ;
        RECT 123.000 152.100 123.400 152.500 ;
        RECT 118.200 151.800 119.200 152.100 ;
        RECT 118.800 151.100 119.200 151.800 ;
        RECT 121.000 151.100 121.400 152.100 ;
        RECT 123.000 151.800 123.700 152.100 ;
        RECT 123.100 151.100 123.700 151.800 ;
        RECT 125.400 151.100 125.800 153.300 ;
        RECT 126.300 153.100 128.100 153.300 ;
        RECT 128.600 153.100 128.900 153.800 ;
        RECT 129.500 153.100 129.800 153.800 ;
        RECT 131.400 153.600 131.800 153.800 ;
        RECT 130.300 153.100 132.100 153.300 ;
        RECT 126.200 153.000 128.200 153.100 ;
        RECT 126.200 151.100 126.600 153.000 ;
        RECT 127.800 151.100 128.200 153.000 ;
        RECT 128.600 151.100 129.000 153.100 ;
        RECT 129.400 151.100 129.800 153.100 ;
        RECT 130.200 153.000 132.200 153.100 ;
        RECT 130.200 151.100 130.600 153.000 ;
        RECT 131.800 151.100 132.200 153.000 ;
        RECT 132.600 151.100 133.000 153.500 ;
        RECT 135.100 152.800 135.400 153.900 ;
        RECT 137.900 153.800 138.300 153.900 ;
        RECT 141.400 153.600 141.800 155.300 ;
        RECT 139.900 153.300 141.800 153.600 ;
        RECT 139.900 153.200 140.300 153.300 ;
        RECT 134.200 152.100 134.600 152.500 ;
        RECT 135.000 152.400 135.400 152.800 ;
        RECT 135.900 152.700 136.300 152.800 ;
        RECT 135.900 152.400 137.300 152.700 ;
        RECT 137.000 152.100 137.300 152.400 ;
        RECT 139.000 152.100 139.400 152.500 ;
        RECT 134.200 151.800 135.200 152.100 ;
        RECT 134.800 151.100 135.200 151.800 ;
        RECT 137.000 151.100 137.400 152.100 ;
        RECT 139.000 151.800 139.700 152.100 ;
        RECT 139.100 151.100 139.700 151.800 ;
        RECT 141.400 151.100 141.800 153.300 ;
        RECT 143.000 153.100 143.400 159.900 ;
        RECT 145.400 155.100 145.800 159.900 ;
        RECT 147.400 156.800 147.800 157.200 ;
        RECT 146.200 155.800 146.600 156.600 ;
        RECT 147.400 156.200 147.700 156.800 ;
        RECT 148.100 156.200 148.500 159.900 ;
        RECT 147.000 155.900 147.700 156.200 ;
        RECT 148.000 155.900 148.500 156.200 ;
        RECT 147.000 155.800 147.400 155.900 ;
        RECT 147.000 155.100 147.300 155.800 ;
        RECT 145.400 154.800 147.300 155.100 ;
        RECT 143.800 153.400 144.200 154.200 ;
        RECT 144.600 153.400 145.000 154.200 ;
        RECT 142.500 152.800 143.400 153.100 ;
        RECT 145.400 153.100 145.800 154.800 ;
        RECT 148.000 154.200 148.300 155.900 ;
        RECT 150.200 155.800 150.600 156.600 ;
        RECT 148.600 155.100 149.000 155.200 ;
        RECT 149.400 155.100 149.800 155.200 ;
        RECT 151.000 155.100 151.400 159.900 ;
        RECT 148.600 154.800 151.400 155.100 ;
        RECT 148.600 154.400 149.000 154.800 ;
        RECT 146.200 154.100 146.600 154.200 ;
        RECT 147.000 154.100 148.300 154.200 ;
        RECT 149.400 154.100 149.800 154.200 ;
        RECT 146.200 153.800 148.300 154.100 ;
        RECT 149.000 153.800 149.800 154.100 ;
        RECT 147.100 153.100 147.400 153.800 ;
        RECT 149.000 153.600 149.400 153.800 ;
        RECT 147.900 153.100 149.700 153.300 ;
        RECT 151.000 153.100 151.400 154.800 ;
        RECT 154.200 155.600 154.600 159.900 ;
        RECT 156.300 157.900 156.900 159.900 ;
        RECT 158.600 157.900 159.000 159.900 ;
        RECT 160.800 158.200 161.200 159.900 ;
        RECT 160.800 157.900 161.800 158.200 ;
        RECT 156.600 157.500 157.000 157.900 ;
        RECT 158.700 157.600 159.000 157.900 ;
        RECT 158.300 157.300 160.100 157.600 ;
        RECT 161.400 157.500 161.800 157.900 ;
        RECT 158.300 157.200 158.700 157.300 ;
        RECT 159.700 157.200 160.100 157.300 ;
        RECT 156.200 156.600 156.900 157.000 ;
        RECT 156.600 156.100 156.900 156.600 ;
        RECT 157.700 156.500 158.800 156.800 ;
        RECT 157.700 156.400 158.100 156.500 ;
        RECT 156.600 155.800 157.800 156.100 ;
        RECT 154.200 155.300 156.300 155.600 ;
        RECT 151.800 153.400 152.200 154.200 ;
        RECT 154.200 153.600 154.600 155.300 ;
        RECT 155.900 155.200 156.300 155.300 ;
        RECT 155.100 154.900 155.500 155.000 ;
        RECT 155.100 154.600 157.000 154.900 ;
        RECT 156.600 154.500 157.000 154.600 ;
        RECT 157.500 154.200 157.800 155.800 ;
        RECT 158.500 155.900 158.800 156.500 ;
        RECT 159.100 156.500 159.500 156.600 ;
        RECT 161.400 156.500 161.800 156.600 ;
        RECT 159.100 156.200 161.800 156.500 ;
        RECT 158.500 155.700 160.900 155.900 ;
        RECT 163.000 155.700 163.400 159.900 ;
        RECT 163.800 155.800 164.200 156.600 ;
        RECT 164.600 156.100 165.000 159.900 ;
        RECT 166.600 156.800 167.000 157.200 ;
        RECT 166.600 156.200 166.900 156.800 ;
        RECT 167.300 156.200 167.700 159.900 ;
        RECT 170.700 156.300 171.100 159.900 ;
        RECT 166.200 156.100 166.900 156.200 ;
        RECT 164.600 155.900 166.900 156.100 ;
        RECT 167.200 155.900 167.700 156.200 ;
        RECT 170.200 155.900 171.100 156.300 ;
        RECT 171.800 156.200 172.200 159.900 ;
        RECT 173.400 156.200 173.800 159.900 ;
        RECT 171.800 155.900 173.800 156.200 ;
        RECT 174.200 155.900 174.600 159.900 ;
        RECT 176.300 159.200 176.700 159.900 ;
        RECT 180.100 159.200 180.500 159.900 ;
        RECT 175.800 158.800 176.700 159.200 ;
        RECT 179.800 158.800 180.500 159.200 ;
        RECT 176.300 156.200 176.700 158.800 ;
        RECT 177.000 156.800 177.800 157.200 ;
        RECT 177.100 156.200 177.400 156.800 ;
        RECT 180.100 156.400 180.500 158.800 ;
        RECT 182.200 157.500 182.600 159.500 ;
        RECT 176.300 155.900 176.800 156.200 ;
        RECT 177.100 155.900 177.800 156.200 ;
        RECT 164.600 155.800 166.600 155.900 ;
        RECT 158.500 155.600 163.400 155.700 ;
        RECT 160.500 155.500 163.400 155.600 ;
        RECT 160.600 155.400 163.400 155.500 ;
        RECT 159.800 155.100 160.200 155.200 ;
        RECT 159.800 154.800 162.300 155.100 ;
        RECT 160.600 154.700 161.000 154.800 ;
        RECT 161.900 154.700 162.300 154.800 ;
        RECT 161.100 154.200 161.500 154.300 ;
        RECT 157.500 153.900 163.000 154.200 ;
        RECT 157.700 153.800 158.100 153.900 ;
        RECT 145.400 152.800 146.300 153.100 ;
        RECT 142.500 151.100 142.900 152.800 ;
        RECT 145.900 151.100 146.300 152.800 ;
        RECT 147.000 151.100 147.400 153.100 ;
        RECT 147.800 153.000 149.800 153.100 ;
        RECT 147.800 151.100 148.200 153.000 ;
        RECT 149.400 151.100 149.800 153.000 ;
        RECT 150.500 152.800 151.400 153.100 ;
        RECT 154.200 153.300 156.100 153.600 ;
        RECT 150.500 151.100 150.900 152.800 ;
        RECT 154.200 151.100 154.600 153.300 ;
        RECT 155.700 153.200 156.100 153.300 ;
        RECT 160.600 152.800 160.900 153.900 ;
        RECT 162.200 153.800 163.000 153.900 ;
        RECT 159.700 152.700 160.100 152.800 ;
        RECT 156.600 152.100 157.000 152.500 ;
        RECT 158.700 152.400 160.100 152.700 ;
        RECT 160.600 152.400 161.000 152.800 ;
        RECT 158.700 152.100 159.000 152.400 ;
        RECT 161.400 152.100 161.800 152.500 ;
        RECT 156.300 151.800 157.000 152.100 ;
        RECT 156.300 151.100 156.900 151.800 ;
        RECT 158.600 151.100 159.000 152.100 ;
        RECT 160.800 151.800 161.800 152.100 ;
        RECT 160.800 151.100 161.200 151.800 ;
        RECT 163.000 151.100 163.400 153.500 ;
        RECT 164.600 153.100 165.000 155.800 ;
        RECT 166.200 155.100 166.600 155.200 ;
        RECT 167.200 155.100 167.500 155.900 ;
        RECT 166.200 154.800 167.500 155.100 ;
        RECT 167.200 154.200 167.500 154.800 ;
        RECT 167.800 155.100 168.200 155.200 ;
        RECT 168.600 155.100 169.000 155.200 ;
        RECT 167.800 154.800 169.000 155.100 ;
        RECT 167.800 154.400 168.200 154.800 ;
        RECT 170.300 154.200 170.600 155.900 ;
        RECT 165.400 153.400 165.800 154.200 ;
        RECT 166.200 153.800 167.500 154.200 ;
        RECT 168.600 154.100 169.000 154.200 ;
        RECT 169.400 154.100 169.800 154.200 ;
        RECT 168.200 153.800 169.800 154.100 ;
        RECT 170.200 153.800 170.600 154.200 ;
        RECT 171.000 154.800 171.400 155.600 ;
        RECT 172.200 155.200 172.600 155.400 ;
        RECT 174.200 155.200 174.500 155.900 ;
        RECT 171.800 154.900 172.600 155.200 ;
        RECT 173.400 154.900 174.600 155.200 ;
        RECT 171.800 154.800 172.200 154.900 ;
        RECT 171.000 154.100 171.300 154.800 ;
        RECT 172.600 154.100 173.000 154.600 ;
        RECT 171.000 153.800 173.000 154.100 ;
        RECT 166.300 153.100 166.600 153.800 ;
        RECT 168.200 153.600 168.600 153.800 ;
        RECT 167.100 153.100 168.900 153.300 ;
        RECT 170.300 153.200 170.600 153.800 ;
        RECT 164.100 152.800 165.000 153.100 ;
        RECT 164.100 151.100 164.500 152.800 ;
        RECT 166.200 151.100 166.600 153.100 ;
        RECT 167.000 153.000 169.000 153.100 ;
        RECT 167.000 151.100 167.400 153.000 ;
        RECT 168.600 151.100 169.000 153.000 ;
        RECT 169.400 152.400 169.800 153.200 ;
        RECT 170.200 152.800 170.600 153.200 ;
        RECT 170.300 152.100 170.600 152.800 ;
        RECT 170.200 151.100 170.600 152.100 ;
        RECT 173.400 153.100 173.700 154.900 ;
        RECT 174.200 154.800 174.600 154.900 ;
        RECT 175.800 154.400 176.200 155.200 ;
        RECT 176.500 154.200 176.800 155.900 ;
        RECT 177.400 155.800 177.800 155.900 ;
        RECT 179.700 156.100 180.500 156.400 ;
        RECT 179.000 154.800 179.400 155.600 ;
        RECT 179.700 154.200 180.000 156.100 ;
        RECT 182.300 155.800 182.600 157.500 ;
        RECT 180.700 155.500 182.600 155.800 ;
        RECT 183.000 155.700 183.400 159.900 ;
        RECT 185.200 158.200 185.600 159.900 ;
        RECT 184.600 157.900 185.600 158.200 ;
        RECT 187.400 157.900 187.800 159.900 ;
        RECT 189.500 157.900 190.100 159.900 ;
        RECT 184.600 157.500 185.000 157.900 ;
        RECT 187.400 157.600 187.700 157.900 ;
        RECT 186.300 157.300 188.100 157.600 ;
        RECT 189.400 157.500 189.800 157.900 ;
        RECT 186.300 157.200 186.700 157.300 ;
        RECT 187.700 157.200 188.100 157.300 ;
        RECT 184.600 156.500 185.000 156.600 ;
        RECT 186.900 156.500 187.300 156.600 ;
        RECT 184.600 156.200 187.300 156.500 ;
        RECT 187.600 156.500 188.700 156.800 ;
        RECT 187.600 155.900 187.900 156.500 ;
        RECT 188.300 156.400 188.700 156.500 ;
        RECT 189.500 156.600 190.200 157.000 ;
        RECT 189.500 156.100 189.800 156.600 ;
        RECT 185.500 155.700 187.900 155.900 ;
        RECT 183.000 155.600 187.900 155.700 ;
        RECT 188.600 155.800 189.800 156.100 ;
        RECT 183.000 155.500 185.900 155.600 ;
        RECT 180.700 154.500 181.000 155.500 ;
        RECT 183.000 155.400 185.800 155.500 ;
        RECT 175.000 154.100 175.400 154.200 ;
        RECT 175.000 153.800 175.800 154.100 ;
        RECT 176.500 153.800 177.800 154.200 ;
        RECT 179.000 153.800 180.000 154.200 ;
        RECT 180.300 154.100 181.000 154.500 ;
        RECT 181.400 154.400 181.800 155.200 ;
        RECT 182.200 154.400 182.600 155.200 ;
        RECT 186.200 155.100 186.600 155.200 ;
        RECT 184.100 154.800 186.600 155.100 ;
        RECT 184.100 154.700 184.500 154.800 ;
        RECT 184.900 154.200 185.300 154.300 ;
        RECT 188.600 154.200 188.900 155.800 ;
        RECT 191.800 155.600 192.200 159.900 ;
        RECT 193.900 156.200 194.300 159.900 ;
        RECT 194.600 156.800 195.000 157.200 ;
        RECT 194.700 156.200 195.000 156.800 ;
        RECT 197.100 156.200 197.500 159.900 ;
        RECT 197.800 156.800 198.200 157.200 ;
        RECT 197.900 156.200 198.200 156.800 ;
        RECT 193.900 155.900 194.400 156.200 ;
        RECT 194.700 155.900 195.400 156.200 ;
        RECT 197.100 155.900 197.600 156.200 ;
        RECT 197.900 156.100 198.600 156.200 ;
        RECT 199.800 156.100 200.200 159.900 ;
        RECT 201.400 156.800 202.200 157.200 ;
        RECT 197.900 155.900 200.200 156.100 ;
        RECT 190.100 155.300 192.200 155.600 ;
        RECT 190.100 155.200 190.500 155.300 ;
        RECT 190.900 154.900 191.300 155.000 ;
        RECT 189.400 154.600 191.300 154.900 ;
        RECT 189.400 154.500 189.800 154.600 ;
        RECT 175.400 153.600 175.800 153.800 ;
        RECT 173.400 151.100 173.800 153.100 ;
        RECT 174.200 152.800 174.600 153.200 ;
        RECT 175.100 153.100 176.900 153.300 ;
        RECT 177.400 153.100 177.700 153.800 ;
        RECT 179.700 153.500 180.000 153.800 ;
        RECT 180.500 153.900 181.000 154.100 ;
        RECT 183.400 153.900 188.900 154.200 ;
        RECT 180.500 153.600 182.600 153.900 ;
        RECT 183.400 153.800 184.200 153.900 ;
        RECT 179.700 153.300 180.100 153.500 ;
        RECT 175.000 153.000 177.000 153.100 ;
        RECT 174.100 152.400 174.500 152.800 ;
        RECT 175.000 151.100 175.400 153.000 ;
        RECT 176.600 151.100 177.000 153.000 ;
        RECT 177.400 151.100 177.800 153.100 ;
        RECT 179.700 153.000 180.500 153.300 ;
        RECT 180.100 151.500 180.500 153.000 ;
        RECT 182.300 152.500 182.600 153.600 ;
        RECT 182.200 151.500 182.600 152.500 ;
        RECT 183.000 151.100 183.400 153.500 ;
        RECT 185.500 152.800 185.800 153.900 ;
        RECT 187.000 153.800 187.400 153.900 ;
        RECT 188.300 153.800 188.700 153.900 ;
        RECT 191.800 153.600 192.200 155.300 ;
        RECT 193.400 154.400 193.800 155.200 ;
        RECT 194.100 155.100 194.400 155.900 ;
        RECT 195.000 155.800 195.400 155.900 ;
        RECT 195.000 155.100 195.400 155.200 ;
        RECT 194.100 154.800 195.400 155.100 ;
        RECT 194.100 154.200 194.400 154.800 ;
        RECT 196.600 154.400 197.000 155.200 ;
        RECT 197.300 154.200 197.600 155.900 ;
        RECT 198.200 155.800 200.200 155.900 ;
        RECT 200.600 155.800 201.000 156.600 ;
        RECT 201.800 156.200 202.100 156.800 ;
        RECT 202.500 156.200 202.900 159.900 ;
        RECT 206.500 156.400 206.900 159.900 ;
        RECT 211.000 159.600 213.000 159.900 ;
        RECT 208.600 157.500 209.000 159.500 ;
        RECT 201.400 155.900 202.100 156.200 ;
        RECT 202.400 155.900 202.900 156.200 ;
        RECT 206.100 156.100 206.900 156.400 ;
        RECT 201.400 155.800 201.800 155.900 ;
        RECT 192.600 154.100 193.000 154.200 ;
        RECT 192.600 153.800 193.400 154.100 ;
        RECT 194.100 153.800 195.400 154.200 ;
        RECT 195.800 154.100 196.200 154.200 ;
        RECT 195.800 153.800 196.600 154.100 ;
        RECT 197.300 153.800 198.600 154.200 ;
        RECT 193.000 153.600 193.400 153.800 ;
        RECT 190.300 153.300 192.200 153.600 ;
        RECT 190.300 153.200 190.700 153.300 ;
        RECT 184.600 152.100 185.000 152.500 ;
        RECT 185.400 152.400 185.800 152.800 ;
        RECT 186.300 152.700 186.700 152.800 ;
        RECT 186.300 152.400 187.700 152.700 ;
        RECT 187.400 152.100 187.700 152.400 ;
        RECT 189.400 152.100 189.800 152.500 ;
        RECT 184.600 151.800 185.600 152.100 ;
        RECT 185.200 151.100 185.600 151.800 ;
        RECT 187.400 151.100 187.800 152.100 ;
        RECT 189.400 151.800 190.100 152.100 ;
        RECT 189.500 151.100 190.100 151.800 ;
        RECT 191.800 151.100 192.200 153.300 ;
        RECT 192.700 153.100 194.500 153.300 ;
        RECT 195.000 153.100 195.300 153.800 ;
        RECT 196.200 153.600 196.600 153.800 ;
        RECT 195.900 153.100 197.700 153.300 ;
        RECT 198.200 153.100 198.500 153.800 ;
        RECT 199.000 153.400 199.400 154.200 ;
        RECT 199.800 153.100 200.200 155.800 ;
        RECT 201.400 155.100 201.800 155.200 ;
        RECT 202.400 155.100 202.700 155.900 ;
        RECT 201.400 154.800 202.700 155.100 ;
        RECT 202.400 154.200 202.700 154.800 ;
        RECT 203.000 154.400 203.400 155.200 ;
        RECT 204.600 155.100 205.000 155.200 ;
        RECT 205.400 155.100 205.800 155.600 ;
        RECT 204.600 154.800 205.800 155.100 ;
        RECT 206.100 155.200 206.400 156.100 ;
        RECT 208.700 155.800 209.000 157.500 ;
        RECT 211.000 155.900 211.400 159.600 ;
        RECT 211.800 155.900 212.200 159.300 ;
        RECT 212.600 156.200 213.000 159.600 ;
        RECT 214.200 156.200 214.600 159.900 ;
        RECT 212.600 155.900 214.600 156.200 ;
        RECT 215.000 157.500 215.400 159.500 ;
        RECT 207.100 155.500 209.000 155.800 ;
        RECT 211.900 155.600 212.200 155.900 ;
        RECT 215.000 155.800 215.300 157.500 ;
        RECT 217.100 156.400 217.500 159.900 ;
        RECT 221.700 159.200 222.100 159.900 ;
        RECT 221.400 158.800 222.100 159.200 ;
        RECT 221.700 156.400 222.100 158.800 ;
        RECT 223.800 157.500 224.200 159.500 ;
        RECT 217.100 156.100 217.900 156.400 ;
        RECT 206.100 154.800 206.600 155.200 ;
        RECT 206.100 154.200 206.400 154.800 ;
        RECT 207.100 154.500 207.400 155.500 ;
        RECT 201.400 153.800 202.700 154.200 ;
        RECT 203.800 154.100 204.200 154.200 ;
        RECT 203.400 153.800 204.200 154.100 ;
        RECT 205.400 153.800 206.400 154.200 ;
        RECT 206.700 154.100 207.400 154.500 ;
        RECT 207.800 154.400 208.200 155.200 ;
        RECT 208.600 154.400 209.000 155.200 ;
        RECT 211.000 154.800 211.400 155.600 ;
        RECT 211.900 155.300 212.900 155.600 ;
        RECT 215.000 155.500 216.900 155.800 ;
        RECT 212.600 155.200 212.900 155.300 ;
        RECT 213.800 155.200 214.200 155.400 ;
        RECT 212.600 154.800 213.000 155.200 ;
        RECT 213.800 154.900 214.600 155.200 ;
        RECT 214.200 154.800 214.600 154.900 ;
        RECT 211.900 154.400 212.300 154.800 ;
        RECT 211.900 154.200 212.200 154.400 ;
        RECT 201.500 153.100 201.800 153.800 ;
        RECT 203.400 153.600 203.800 153.800 ;
        RECT 206.100 153.500 206.400 153.800 ;
        RECT 206.900 153.900 207.400 154.100 ;
        RECT 206.900 153.600 209.000 153.900 ;
        RECT 211.800 153.800 212.200 154.200 ;
        RECT 206.100 153.300 206.500 153.500 ;
        RECT 202.300 153.100 204.100 153.300 ;
        RECT 192.600 153.000 194.600 153.100 ;
        RECT 192.600 151.100 193.000 153.000 ;
        RECT 194.200 151.100 194.600 153.000 ;
        RECT 195.000 151.100 195.400 153.100 ;
        RECT 195.800 153.000 197.800 153.100 ;
        RECT 195.800 151.100 196.200 153.000 ;
        RECT 197.400 151.100 197.800 153.000 ;
        RECT 198.200 151.100 198.600 153.100 ;
        RECT 199.800 152.800 200.700 153.100 ;
        RECT 200.300 151.100 200.700 152.800 ;
        RECT 201.400 151.100 201.800 153.100 ;
        RECT 202.200 153.000 204.200 153.100 ;
        RECT 206.100 153.000 206.900 153.300 ;
        RECT 202.200 151.100 202.600 153.000 ;
        RECT 203.800 151.100 204.200 153.000 ;
        RECT 206.500 151.500 206.900 153.000 ;
        RECT 208.700 152.500 209.000 153.600 ;
        RECT 212.600 153.100 212.900 154.800 ;
        RECT 213.400 153.800 213.800 154.600 ;
        RECT 215.000 154.400 215.400 155.200 ;
        RECT 215.800 154.400 216.200 155.200 ;
        RECT 216.600 154.500 216.900 155.500 ;
        RECT 216.600 154.100 217.300 154.500 ;
        RECT 217.600 154.200 217.900 156.100 ;
        RECT 221.300 156.100 222.100 156.400 ;
        RECT 218.200 155.100 218.600 155.600 ;
        RECT 219.000 155.100 219.400 155.200 ;
        RECT 218.200 154.800 219.400 155.100 ;
        RECT 220.600 154.800 221.000 155.600 ;
        RECT 221.300 154.200 221.600 156.100 ;
        RECT 223.900 155.800 224.200 157.500 ;
        RECT 222.300 155.500 224.200 155.800 ;
        RECT 224.600 157.500 225.000 159.500 ;
        RECT 226.700 159.200 227.100 159.900 ;
        RECT 226.200 158.800 227.100 159.200 ;
        RECT 224.600 155.800 224.900 157.500 ;
        RECT 226.700 156.400 227.100 158.800 ;
        RECT 226.700 156.100 227.500 156.400 ;
        RECT 224.600 155.500 226.500 155.800 ;
        RECT 222.300 154.500 222.600 155.500 ;
        RECT 216.600 153.900 217.100 154.100 ;
        RECT 215.000 153.600 217.100 153.900 ;
        RECT 217.600 153.800 218.600 154.200 ;
        RECT 220.600 153.800 221.600 154.200 ;
        RECT 221.900 154.100 222.600 154.500 ;
        RECT 223.000 154.400 223.400 155.200 ;
        RECT 223.800 154.400 224.200 155.200 ;
        RECT 224.600 154.400 225.000 155.200 ;
        RECT 225.400 154.400 225.800 155.200 ;
        RECT 226.200 154.500 226.500 155.500 ;
        RECT 208.600 151.500 209.000 152.500 ;
        RECT 212.300 151.100 213.100 153.100 ;
        RECT 215.000 152.500 215.300 153.600 ;
        RECT 217.600 153.500 217.900 153.800 ;
        RECT 217.500 153.300 217.900 153.500 ;
        RECT 217.100 153.200 217.900 153.300 ;
        RECT 216.600 153.000 217.900 153.200 ;
        RECT 221.300 153.500 221.600 153.800 ;
        RECT 222.100 153.900 222.600 154.100 ;
        RECT 226.200 154.100 226.900 154.500 ;
        RECT 227.200 154.200 227.500 156.100 ;
        RECT 229.400 155.900 229.800 159.900 ;
        RECT 230.200 156.200 230.600 159.900 ;
        RECT 231.800 156.200 232.200 159.900 ;
        RECT 230.200 155.900 232.200 156.200 ;
        RECT 227.800 154.800 228.200 155.600 ;
        RECT 229.500 155.200 229.800 155.900 ;
        RECT 232.600 155.700 233.000 159.900 ;
        RECT 234.800 158.200 235.200 159.900 ;
        RECT 234.200 157.900 235.200 158.200 ;
        RECT 237.000 157.900 237.400 159.900 ;
        RECT 239.100 157.900 239.700 159.900 ;
        RECT 234.200 157.500 234.600 157.900 ;
        RECT 237.000 157.600 237.300 157.900 ;
        RECT 235.900 157.300 237.700 157.600 ;
        RECT 239.000 157.500 239.400 157.900 ;
        RECT 235.900 157.200 236.300 157.300 ;
        RECT 237.300 157.200 237.700 157.300 ;
        RECT 241.400 157.100 241.800 159.900 ;
        RECT 234.200 156.500 234.600 156.600 ;
        RECT 236.500 156.500 236.900 156.600 ;
        RECT 234.200 156.200 236.900 156.500 ;
        RECT 237.200 156.500 238.300 156.800 ;
        RECT 237.200 155.900 237.500 156.500 ;
        RECT 237.900 156.400 238.300 156.500 ;
        RECT 239.100 156.600 239.800 157.000 ;
        RECT 241.400 156.800 242.600 157.100 ;
        RECT 239.100 156.100 239.400 156.600 ;
        RECT 235.100 155.700 237.500 155.900 ;
        RECT 232.600 155.600 237.500 155.700 ;
        RECT 238.200 155.800 239.400 156.100 ;
        RECT 232.600 155.500 235.500 155.600 ;
        RECT 232.600 155.400 235.400 155.500 ;
        RECT 231.400 155.200 231.800 155.400 ;
        RECT 229.400 154.900 230.600 155.200 ;
        RECT 231.400 154.900 232.200 155.200 ;
        RECT 235.800 155.100 236.200 155.200 ;
        RECT 229.400 154.800 229.800 154.900 ;
        RECT 230.200 154.800 230.600 154.900 ;
        RECT 231.800 154.800 232.200 154.900 ;
        RECT 233.700 154.800 236.200 155.100 ;
        RECT 226.200 153.900 226.700 154.100 ;
        RECT 222.100 153.600 224.200 153.900 ;
        RECT 221.300 153.300 221.700 153.500 ;
        RECT 221.300 153.000 222.100 153.300 ;
        RECT 216.600 152.800 217.500 153.000 ;
        RECT 215.000 151.500 215.400 152.500 ;
        RECT 217.100 151.500 217.500 152.800 ;
        RECT 221.700 151.500 222.100 153.000 ;
        RECT 223.900 152.500 224.200 153.600 ;
        RECT 223.800 151.500 224.200 152.500 ;
        RECT 224.600 153.600 226.700 153.900 ;
        RECT 227.200 153.800 228.200 154.200 ;
        RECT 224.600 152.500 224.900 153.600 ;
        RECT 227.200 153.500 227.500 153.800 ;
        RECT 227.100 153.300 227.500 153.500 ;
        RECT 226.700 153.000 227.500 153.300 ;
        RECT 224.600 151.500 225.000 152.500 ;
        RECT 226.700 151.500 227.100 153.000 ;
        RECT 229.400 152.800 229.800 153.200 ;
        RECT 230.300 153.100 230.600 154.800 ;
        RECT 233.700 154.700 234.100 154.800 ;
        RECT 235.000 154.700 235.400 154.800 ;
        RECT 231.000 153.800 231.400 154.600 ;
        RECT 234.500 154.200 234.900 154.300 ;
        RECT 238.200 154.200 238.500 155.800 ;
        RECT 241.400 155.600 241.800 156.800 ;
        RECT 242.200 155.800 242.600 156.800 ;
        RECT 239.700 155.300 241.800 155.600 ;
        RECT 239.700 155.200 240.100 155.300 ;
        RECT 240.500 154.900 240.900 155.000 ;
        RECT 239.000 154.600 240.900 154.900 ;
        RECT 239.000 154.500 239.400 154.600 ;
        RECT 233.000 153.900 238.500 154.200 ;
        RECT 233.000 153.800 233.800 153.900 ;
        RECT 229.500 152.400 229.900 152.800 ;
        RECT 230.200 151.100 230.600 153.100 ;
        RECT 232.600 151.100 233.000 153.500 ;
        RECT 235.100 152.800 235.400 153.900 ;
        RECT 237.900 153.800 238.300 153.900 ;
        RECT 241.400 153.600 241.800 155.300 ;
        RECT 243.000 155.100 243.400 159.900 ;
        RECT 242.200 154.800 243.400 155.100 ;
        RECT 242.200 154.200 242.500 154.800 ;
        RECT 242.200 153.800 242.600 154.200 ;
        RECT 239.900 153.300 241.800 153.600 ;
        RECT 239.900 153.200 240.300 153.300 ;
        RECT 234.200 152.100 234.600 152.500 ;
        RECT 235.000 152.400 235.400 152.800 ;
        RECT 235.900 152.700 236.300 152.800 ;
        RECT 235.900 152.400 237.300 152.700 ;
        RECT 237.000 152.100 237.300 152.400 ;
        RECT 239.000 152.100 239.400 152.500 ;
        RECT 234.200 151.800 235.200 152.100 ;
        RECT 234.800 151.100 235.200 151.800 ;
        RECT 237.000 151.100 237.400 152.100 ;
        RECT 239.000 151.800 239.700 152.100 ;
        RECT 239.100 151.100 239.700 151.800 ;
        RECT 241.400 151.100 241.800 153.300 ;
        RECT 243.000 153.100 243.400 154.800 ;
        RECT 245.400 155.100 245.800 159.900 ;
        RECT 247.400 156.800 247.800 157.200 ;
        RECT 246.200 155.800 246.600 156.600 ;
        RECT 247.400 156.200 247.700 156.800 ;
        RECT 248.100 156.200 248.500 159.900 ;
        RECT 247.000 155.900 247.700 156.200 ;
        RECT 248.000 155.900 248.500 156.200 ;
        RECT 247.000 155.800 247.400 155.900 ;
        RECT 247.000 155.100 247.300 155.800 ;
        RECT 245.400 154.800 247.300 155.100 ;
        RECT 244.600 153.400 245.000 154.200 ;
        RECT 242.500 152.800 243.400 153.100 ;
        RECT 245.400 153.100 245.800 154.800 ;
        RECT 248.000 154.200 248.300 155.900 ;
        RECT 248.600 154.400 249.000 155.200 ;
        RECT 251.000 155.100 251.400 159.900 ;
        RECT 253.000 156.800 253.400 157.200 ;
        RECT 251.800 155.800 252.200 156.600 ;
        RECT 253.000 156.200 253.300 156.800 ;
        RECT 253.700 156.200 254.100 159.900 ;
        RECT 252.600 155.900 253.300 156.200 ;
        RECT 253.600 155.900 254.100 156.200 ;
        RECT 252.600 155.800 253.000 155.900 ;
        RECT 252.600 155.100 252.900 155.800 ;
        RECT 251.000 154.800 252.900 155.100 ;
        RECT 247.000 153.800 248.300 154.200 ;
        RECT 249.400 154.100 249.800 154.200 ;
        RECT 249.000 153.800 249.800 154.100 ;
        RECT 247.100 153.100 247.400 153.800 ;
        RECT 249.000 153.600 249.400 153.800 ;
        RECT 250.200 153.400 250.600 154.200 ;
        RECT 247.900 153.100 249.700 153.300 ;
        RECT 251.000 153.100 251.400 154.800 ;
        RECT 253.600 154.200 253.900 155.900 ;
        RECT 255.800 155.600 256.200 159.900 ;
        RECT 257.900 157.900 258.500 159.900 ;
        RECT 260.200 157.900 260.600 159.900 ;
        RECT 262.400 158.200 262.800 159.900 ;
        RECT 262.400 157.900 263.400 158.200 ;
        RECT 258.200 157.500 258.600 157.900 ;
        RECT 260.300 157.600 260.600 157.900 ;
        RECT 259.900 157.300 261.700 157.600 ;
        RECT 263.000 157.500 263.400 157.900 ;
        RECT 259.900 157.200 260.300 157.300 ;
        RECT 261.300 157.200 261.700 157.300 ;
        RECT 257.800 156.600 258.500 157.000 ;
        RECT 258.200 156.100 258.500 156.600 ;
        RECT 259.300 156.500 260.400 156.800 ;
        RECT 259.300 156.400 259.700 156.500 ;
        RECT 258.200 155.800 259.400 156.100 ;
        RECT 255.800 155.300 257.900 155.600 ;
        RECT 254.200 154.400 254.600 155.200 ;
        RECT 252.600 153.800 253.900 154.200 ;
        RECT 255.000 154.100 255.400 154.200 ;
        RECT 254.600 153.800 255.400 154.100 ;
        RECT 252.700 153.100 253.000 153.800 ;
        RECT 254.600 153.600 255.000 153.800 ;
        RECT 255.800 153.600 256.200 155.300 ;
        RECT 257.500 155.200 257.900 155.300 ;
        RECT 259.100 155.200 259.400 155.800 ;
        RECT 260.100 155.900 260.400 156.500 ;
        RECT 260.700 156.500 261.100 156.600 ;
        RECT 263.000 156.500 263.400 156.600 ;
        RECT 260.700 156.200 263.400 156.500 ;
        RECT 260.100 155.700 262.500 155.900 ;
        RECT 264.600 155.700 265.000 159.900 ;
        RECT 260.100 155.600 265.000 155.700 ;
        RECT 262.100 155.500 265.000 155.600 ;
        RECT 262.200 155.400 265.000 155.500 ;
        RECT 256.700 154.900 257.100 155.000 ;
        RECT 256.700 154.600 258.600 154.900 ;
        RECT 259.000 154.800 259.400 155.200 ;
        RECT 259.800 155.100 260.200 155.200 ;
        RECT 261.400 155.100 261.800 155.200 ;
        RECT 259.800 154.800 263.900 155.100 ;
        RECT 258.200 154.500 258.600 154.600 ;
        RECT 259.100 154.200 259.400 154.800 ;
        RECT 263.500 154.700 263.900 154.800 ;
        RECT 262.700 154.200 263.100 154.300 ;
        RECT 259.100 153.900 264.600 154.200 ;
        RECT 259.300 153.800 259.700 153.900 ;
        RECT 255.800 153.300 257.700 153.600 ;
        RECT 253.500 153.100 255.300 153.300 ;
        RECT 245.400 152.800 246.300 153.100 ;
        RECT 242.500 151.100 242.900 152.800 ;
        RECT 245.900 151.100 246.300 152.800 ;
        RECT 247.000 151.100 247.400 153.100 ;
        RECT 247.800 153.000 249.800 153.100 ;
        RECT 247.800 151.100 248.200 153.000 ;
        RECT 249.400 151.100 249.800 153.000 ;
        RECT 251.000 152.800 251.900 153.100 ;
        RECT 251.500 151.100 251.900 152.800 ;
        RECT 252.600 151.100 253.000 153.100 ;
        RECT 253.400 153.000 255.400 153.100 ;
        RECT 253.400 151.100 253.800 153.000 ;
        RECT 255.000 151.100 255.400 153.000 ;
        RECT 255.800 151.100 256.200 153.300 ;
        RECT 257.300 153.200 257.700 153.300 ;
        RECT 262.200 152.800 262.500 153.900 ;
        RECT 263.800 153.800 264.600 153.900 ;
        RECT 261.300 152.700 261.700 152.800 ;
        RECT 258.200 152.100 258.600 152.500 ;
        RECT 260.300 152.400 261.700 152.700 ;
        RECT 262.200 152.400 262.600 152.800 ;
        RECT 260.300 152.100 260.600 152.400 ;
        RECT 263.000 152.100 263.400 152.500 ;
        RECT 257.900 151.800 258.600 152.100 ;
        RECT 257.900 151.100 258.500 151.800 ;
        RECT 260.200 151.100 260.600 152.100 ;
        RECT 262.400 151.800 263.400 152.100 ;
        RECT 262.400 151.100 262.800 151.800 ;
        RECT 264.600 151.100 265.000 153.500 ;
        RECT 0.600 147.500 1.000 149.900 ;
        RECT 2.800 149.200 3.200 149.900 ;
        RECT 2.200 148.900 3.200 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.100 149.200 7.700 149.900 ;
        RECT 7.000 148.900 7.700 149.200 ;
        RECT 2.200 148.500 2.600 148.900 ;
        RECT 5.000 148.600 5.300 148.900 ;
        RECT 3.000 148.200 3.400 148.600 ;
        RECT 3.900 148.300 5.300 148.600 ;
        RECT 7.000 148.500 7.400 148.900 ;
        RECT 3.900 148.200 4.300 148.300 ;
        RECT 1.000 147.100 1.800 147.200 ;
        RECT 3.100 147.100 3.400 148.200 ;
        RECT 7.900 147.700 8.300 147.800 ;
        RECT 9.400 147.700 9.800 149.900 ;
        RECT 10.200 147.800 10.600 149.900 ;
        RECT 11.000 148.000 11.400 149.900 ;
        RECT 12.600 148.000 13.000 149.900 ;
        RECT 11.000 147.900 13.000 148.000 ;
        RECT 13.400 148.000 13.800 149.900 ;
        RECT 15.000 148.000 15.400 149.900 ;
        RECT 13.400 147.900 15.400 148.000 ;
        RECT 15.800 147.900 16.200 149.900 ;
        RECT 16.900 148.200 17.300 149.900 ;
        RECT 19.000 148.500 19.400 149.500 ;
        RECT 16.900 147.900 17.800 148.200 ;
        RECT 7.900 147.400 9.800 147.700 ;
        RECT 5.900 147.100 6.300 147.200 ;
        RECT 1.000 146.800 6.500 147.100 ;
        RECT 2.500 146.700 2.900 146.800 ;
        RECT 1.700 146.200 2.100 146.300 ;
        RECT 1.700 145.900 4.200 146.200 ;
        RECT 3.800 145.800 4.200 145.900 ;
        RECT 0.600 145.500 3.400 145.600 ;
        RECT 0.600 145.400 3.500 145.500 ;
        RECT 0.600 145.300 5.500 145.400 ;
        RECT 0.600 141.100 1.000 145.300 ;
        RECT 3.100 145.100 5.500 145.300 ;
        RECT 2.200 144.500 4.900 144.800 ;
        RECT 2.200 144.400 2.600 144.500 ;
        RECT 4.500 144.400 4.900 144.500 ;
        RECT 5.200 144.500 5.500 145.100 ;
        RECT 6.200 145.200 6.500 146.800 ;
        RECT 7.000 146.400 7.400 146.500 ;
        RECT 7.000 146.100 8.900 146.400 ;
        RECT 8.500 146.000 8.900 146.100 ;
        RECT 7.700 145.700 8.100 145.800 ;
        RECT 9.400 145.700 9.800 147.400 ;
        RECT 10.300 147.200 10.600 147.800 ;
        RECT 11.100 147.700 12.900 147.900 ;
        RECT 13.500 147.700 15.300 147.900 ;
        RECT 12.200 147.200 12.600 147.400 ;
        RECT 13.800 147.200 14.200 147.400 ;
        RECT 15.800 147.200 16.100 147.900 ;
        RECT 10.200 146.800 11.500 147.200 ;
        RECT 12.200 147.100 13.000 147.200 ;
        RECT 13.400 147.100 14.200 147.200 ;
        RECT 12.200 146.900 14.200 147.100 ;
        RECT 12.600 146.800 13.800 146.900 ;
        RECT 14.900 146.800 16.200 147.200 ;
        RECT 7.700 145.400 9.800 145.700 ;
        RECT 6.200 144.900 7.400 145.200 ;
        RECT 5.900 144.500 6.300 144.600 ;
        RECT 5.200 144.200 6.300 144.500 ;
        RECT 7.100 144.400 7.400 144.900 ;
        RECT 7.100 144.000 7.800 144.400 ;
        RECT 3.900 143.700 4.300 143.800 ;
        RECT 5.300 143.700 5.700 143.800 ;
        RECT 2.200 143.100 2.600 143.500 ;
        RECT 3.900 143.400 5.700 143.700 ;
        RECT 5.000 143.100 5.300 143.400 ;
        RECT 7.000 143.100 7.400 143.500 ;
        RECT 2.200 142.800 3.200 143.100 ;
        RECT 2.800 141.100 3.200 142.800 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.100 141.100 7.700 143.100 ;
        RECT 9.400 141.100 9.800 145.400 ;
        RECT 10.200 145.100 10.600 145.200 ;
        RECT 11.200 145.100 11.500 146.800 ;
        RECT 11.800 145.800 12.200 146.600 ;
        RECT 14.200 145.800 14.600 146.600 ;
        RECT 14.900 145.200 15.200 146.800 ;
        RECT 17.400 146.100 17.800 147.900 ;
        RECT 18.200 146.800 18.600 147.600 ;
        RECT 19.000 147.400 19.300 148.500 ;
        RECT 21.100 148.000 21.500 149.500 ;
        RECT 21.100 147.700 21.900 148.000 ;
        RECT 21.500 147.500 21.900 147.700 ;
        RECT 19.000 147.100 21.100 147.400 ;
        RECT 20.600 146.900 21.100 147.100 ;
        RECT 21.600 147.200 21.900 147.500 ;
        RECT 24.600 147.600 25.000 149.900 ;
        RECT 26.200 147.600 26.600 149.900 ;
        RECT 27.800 147.600 28.200 149.900 ;
        RECT 29.400 147.600 29.800 149.900 ;
        RECT 31.000 148.500 31.400 149.500 ;
        RECT 33.100 149.200 33.500 149.500 ;
        RECT 32.600 148.800 33.500 149.200 ;
        RECT 24.600 147.200 25.500 147.600 ;
        RECT 26.200 147.200 27.300 147.600 ;
        RECT 27.800 147.200 28.900 147.600 ;
        RECT 29.400 147.200 30.600 147.600 ;
        RECT 10.200 144.800 10.900 145.100 ;
        RECT 11.200 144.800 11.700 145.100 ;
        RECT 14.200 144.800 15.200 145.200 ;
        RECT 15.800 145.800 17.800 146.100 ;
        RECT 19.000 145.800 19.400 146.600 ;
        RECT 19.800 145.800 20.200 146.600 ;
        RECT 20.600 146.500 21.300 146.900 ;
        RECT 21.600 146.800 22.600 147.200 ;
        RECT 23.800 146.900 24.200 147.200 ;
        RECT 25.100 146.900 25.500 147.200 ;
        RECT 26.900 146.900 27.300 147.200 ;
        RECT 28.500 146.900 28.900 147.200 ;
        RECT 15.800 145.200 16.100 145.800 ;
        RECT 15.800 145.100 16.200 145.200 ;
        RECT 15.500 144.800 16.200 145.100 ;
        RECT 10.600 144.200 10.900 144.800 ;
        RECT 10.600 143.800 11.000 144.200 ;
        RECT 11.300 141.100 11.700 144.800 ;
        RECT 14.700 141.100 15.100 144.800 ;
        RECT 15.500 144.200 15.800 144.800 ;
        RECT 16.600 144.400 17.000 145.200 ;
        RECT 15.400 143.800 15.800 144.200 ;
        RECT 17.400 141.100 17.800 145.800 ;
        RECT 20.600 145.500 20.900 146.500 ;
        RECT 19.000 145.200 20.900 145.500 ;
        RECT 19.000 143.500 19.300 145.200 ;
        RECT 21.600 144.900 21.900 146.800 ;
        RECT 23.800 146.500 24.700 146.900 ;
        RECT 25.100 146.500 26.400 146.900 ;
        RECT 26.900 146.500 28.100 146.900 ;
        RECT 28.500 146.500 29.800 146.900 ;
        RECT 22.200 145.400 22.600 146.200 ;
        RECT 25.100 145.800 25.500 146.500 ;
        RECT 26.900 145.800 27.300 146.500 ;
        RECT 28.500 145.800 28.900 146.500 ;
        RECT 30.200 145.800 30.600 147.200 ;
        RECT 31.000 147.400 31.300 148.500 ;
        RECT 33.100 148.000 33.500 148.800 ;
        RECT 33.100 147.700 33.900 148.000 ;
        RECT 33.500 147.500 33.900 147.700 ;
        RECT 31.000 147.100 33.100 147.400 ;
        RECT 32.600 146.900 33.100 147.100 ;
        RECT 33.600 147.200 33.900 147.500 ;
        RECT 31.000 145.800 31.400 146.600 ;
        RECT 31.800 145.800 32.200 146.600 ;
        RECT 32.600 146.500 33.300 146.900 ;
        RECT 33.600 146.800 34.600 147.200 ;
        RECT 24.600 145.400 25.500 145.800 ;
        RECT 26.200 145.400 27.300 145.800 ;
        RECT 27.800 145.400 28.900 145.800 ;
        RECT 29.400 145.400 30.600 145.800 ;
        RECT 32.600 145.500 32.900 146.500 ;
        RECT 21.100 144.600 21.900 144.900 ;
        RECT 19.000 141.500 19.400 143.500 ;
        RECT 21.100 142.200 21.500 144.600 ;
        RECT 21.100 141.800 21.800 142.200 ;
        RECT 21.100 141.100 21.500 141.800 ;
        RECT 24.600 141.100 25.000 145.400 ;
        RECT 26.200 141.100 26.600 145.400 ;
        RECT 27.800 141.100 28.200 145.400 ;
        RECT 29.400 141.100 29.800 145.400 ;
        RECT 31.000 145.200 32.900 145.500 ;
        RECT 31.000 143.500 31.300 145.200 ;
        RECT 33.600 144.900 33.900 146.800 ;
        RECT 34.200 146.100 34.600 146.200 ;
        RECT 35.800 146.100 36.200 149.900 ;
        RECT 36.600 147.800 37.000 148.600 ;
        RECT 37.400 148.500 37.800 149.500 ;
        RECT 39.500 149.200 39.900 149.500 ;
        RECT 39.500 148.800 40.200 149.200 ;
        RECT 37.400 147.400 37.700 148.500 ;
        RECT 39.500 148.000 39.900 148.800 ;
        RECT 39.500 147.700 40.300 148.000 ;
        RECT 39.900 147.500 40.300 147.700 ;
        RECT 37.400 147.100 39.500 147.400 ;
        RECT 39.000 146.900 39.500 147.100 ;
        RECT 40.000 147.200 40.300 147.500 ;
        RECT 43.000 147.600 43.400 149.900 ;
        RECT 44.600 147.600 45.000 149.900 ;
        RECT 46.200 147.600 46.600 149.900 ;
        RECT 47.800 147.600 48.200 149.900 ;
        RECT 43.000 147.200 43.900 147.600 ;
        RECT 44.600 147.200 45.700 147.600 ;
        RECT 46.200 147.200 47.300 147.600 ;
        RECT 47.800 147.200 49.000 147.600 ;
        RECT 49.400 147.500 49.800 149.900 ;
        RECT 51.600 149.200 52.000 149.900 ;
        RECT 51.000 148.900 52.000 149.200 ;
        RECT 53.800 148.900 54.200 149.900 ;
        RECT 55.900 149.200 56.500 149.900 ;
        RECT 55.800 148.900 56.500 149.200 ;
        RECT 51.000 148.500 51.400 148.900 ;
        RECT 53.800 148.600 54.100 148.900 ;
        RECT 51.800 148.200 52.200 148.600 ;
        RECT 52.700 148.300 54.100 148.600 ;
        RECT 55.800 148.500 56.200 148.900 ;
        RECT 52.700 148.200 53.100 148.300 ;
        RECT 34.200 145.800 36.200 146.100 ;
        RECT 37.400 145.800 37.800 146.600 ;
        RECT 38.200 145.800 38.600 146.600 ;
        RECT 39.000 146.500 39.700 146.900 ;
        RECT 40.000 146.800 41.000 147.200 ;
        RECT 42.200 146.900 42.600 147.200 ;
        RECT 43.500 146.900 43.900 147.200 ;
        RECT 45.300 146.900 45.700 147.200 ;
        RECT 46.900 146.900 47.300 147.200 ;
        RECT 34.200 145.400 34.600 145.800 ;
        RECT 33.100 144.600 33.900 144.900 ;
        RECT 31.000 141.500 31.400 143.500 ;
        RECT 33.100 141.100 33.500 144.600 ;
        RECT 35.800 141.100 36.200 145.800 ;
        RECT 39.000 145.500 39.300 146.500 ;
        RECT 37.400 145.200 39.300 145.500 ;
        RECT 37.400 143.500 37.700 145.200 ;
        RECT 40.000 144.900 40.300 146.800 ;
        RECT 42.200 146.500 43.100 146.900 ;
        RECT 43.500 146.500 44.800 146.900 ;
        RECT 45.300 146.500 46.500 146.900 ;
        RECT 46.900 146.500 48.200 146.900 ;
        RECT 40.600 145.400 41.000 146.200 ;
        RECT 43.500 145.800 43.900 146.500 ;
        RECT 45.300 145.800 45.700 146.500 ;
        RECT 46.900 145.800 47.300 146.500 ;
        RECT 48.600 145.800 49.000 147.200 ;
        RECT 49.800 147.100 50.600 147.200 ;
        RECT 51.900 147.100 52.200 148.200 ;
        RECT 56.700 147.700 57.100 147.800 ;
        RECT 58.200 147.700 58.600 149.900 ;
        RECT 60.600 148.000 61.000 149.900 ;
        RECT 62.200 148.000 62.600 149.900 ;
        RECT 60.600 147.900 62.600 148.000 ;
        RECT 63.000 147.900 63.400 149.900 ;
        RECT 64.100 148.200 64.500 149.900 ;
        RECT 66.200 148.500 66.600 149.500 ;
        RECT 64.100 147.900 65.000 148.200 ;
        RECT 60.700 147.700 62.500 147.900 ;
        RECT 56.700 147.400 58.600 147.700 ;
        RECT 54.700 147.100 55.100 147.200 ;
        RECT 49.800 146.800 55.300 147.100 ;
        RECT 51.300 146.700 51.700 146.800 ;
        RECT 50.500 146.200 50.900 146.300 ;
        RECT 50.500 145.900 53.000 146.200 ;
        RECT 52.600 145.800 53.000 145.900 ;
        RECT 43.000 145.400 43.900 145.800 ;
        RECT 44.600 145.400 45.700 145.800 ;
        RECT 46.200 145.400 47.300 145.800 ;
        RECT 47.800 145.400 49.000 145.800 ;
        RECT 49.400 145.500 52.200 145.600 ;
        RECT 49.400 145.400 52.300 145.500 ;
        RECT 39.500 144.600 40.300 144.900 ;
        RECT 37.400 141.500 37.800 143.500 ;
        RECT 39.500 141.100 39.900 144.600 ;
        RECT 43.000 141.100 43.400 145.400 ;
        RECT 44.600 141.100 45.000 145.400 ;
        RECT 46.200 141.100 46.600 145.400 ;
        RECT 47.800 141.100 48.200 145.400 ;
        RECT 49.400 145.300 54.300 145.400 ;
        RECT 49.400 141.100 49.800 145.300 ;
        RECT 51.900 145.100 54.300 145.300 ;
        RECT 51.000 144.500 53.700 144.800 ;
        RECT 51.000 144.400 51.400 144.500 ;
        RECT 53.300 144.400 53.700 144.500 ;
        RECT 54.000 144.500 54.300 145.100 ;
        RECT 55.000 145.200 55.300 146.800 ;
        RECT 55.800 146.400 56.200 146.500 ;
        RECT 55.800 146.100 57.700 146.400 ;
        RECT 57.300 146.000 57.700 146.100 ;
        RECT 56.500 145.700 56.900 145.800 ;
        RECT 58.200 145.700 58.600 147.400 ;
        RECT 61.000 147.200 61.400 147.400 ;
        RECT 63.000 147.200 63.300 147.900 ;
        RECT 59.800 147.100 60.200 147.200 ;
        RECT 60.600 147.100 61.400 147.200 ;
        RECT 59.800 146.900 61.400 147.100 ;
        RECT 59.800 146.800 61.000 146.900 ;
        RECT 62.100 146.800 63.400 147.200 ;
        RECT 61.400 145.800 61.800 146.600 ;
        RECT 62.100 146.200 62.400 146.800 ;
        RECT 62.100 145.800 62.600 146.200 ;
        RECT 64.600 146.100 65.000 147.900 ;
        RECT 63.000 145.800 65.000 146.100 ;
        RECT 65.400 146.800 65.800 147.600 ;
        RECT 66.200 147.400 66.500 148.500 ;
        RECT 68.300 148.000 68.700 149.500 ;
        RECT 71.000 148.500 71.400 149.500 ;
        RECT 68.300 147.700 69.100 148.000 ;
        RECT 68.700 147.500 69.100 147.700 ;
        RECT 66.200 147.100 68.300 147.400 ;
        RECT 67.800 146.900 68.300 147.100 ;
        RECT 68.800 147.200 69.100 147.500 ;
        RECT 71.000 147.400 71.300 148.500 ;
        RECT 73.100 148.000 73.500 149.500 ;
        RECT 73.100 147.700 73.900 148.000 ;
        RECT 73.500 147.500 73.900 147.700 ;
        RECT 65.400 146.200 65.700 146.800 ;
        RECT 65.400 145.800 65.800 146.200 ;
        RECT 66.200 145.800 66.600 146.600 ;
        RECT 67.000 145.800 67.400 146.600 ;
        RECT 67.800 146.500 68.500 146.900 ;
        RECT 68.800 146.800 69.800 147.200 ;
        RECT 71.000 147.100 73.100 147.400 ;
        RECT 72.600 146.900 73.100 147.100 ;
        RECT 73.600 147.200 73.900 147.500 ;
        RECT 75.800 147.700 76.200 149.900 ;
        RECT 77.900 149.200 78.500 149.900 ;
        RECT 77.900 148.900 78.600 149.200 ;
        RECT 80.200 148.900 80.600 149.900 ;
        RECT 82.400 149.200 82.800 149.900 ;
        RECT 82.400 148.900 83.400 149.200 ;
        RECT 78.200 148.500 78.600 148.900 ;
        RECT 80.300 148.600 80.600 148.900 ;
        RECT 80.300 148.300 81.700 148.600 ;
        RECT 81.300 148.200 81.700 148.300 ;
        RECT 82.200 148.200 82.600 148.600 ;
        RECT 83.000 148.500 83.400 148.900 ;
        RECT 77.300 147.700 77.700 147.800 ;
        RECT 75.800 147.400 77.700 147.700 ;
        RECT 56.500 145.400 58.600 145.700 ;
        RECT 55.000 144.900 56.200 145.200 ;
        RECT 54.700 144.500 55.100 144.600 ;
        RECT 54.000 144.200 55.100 144.500 ;
        RECT 55.900 144.400 56.200 144.900 ;
        RECT 55.900 144.000 56.600 144.400 ;
        RECT 52.700 143.700 53.100 143.800 ;
        RECT 54.100 143.700 54.500 143.800 ;
        RECT 51.000 143.100 51.400 143.500 ;
        RECT 52.700 143.400 54.500 143.700 ;
        RECT 53.800 143.100 54.100 143.400 ;
        RECT 55.800 143.100 56.200 143.500 ;
        RECT 51.000 142.800 52.000 143.100 ;
        RECT 51.600 141.100 52.000 142.800 ;
        RECT 53.800 141.100 54.200 143.100 ;
        RECT 55.900 141.100 56.500 143.100 ;
        RECT 58.200 141.100 58.600 145.400 ;
        RECT 62.100 145.100 62.400 145.800 ;
        RECT 63.000 145.200 63.300 145.800 ;
        RECT 63.000 145.100 63.400 145.200 ;
        RECT 61.900 144.800 62.400 145.100 ;
        RECT 62.700 144.800 63.400 145.100 ;
        RECT 61.900 141.100 62.300 144.800 ;
        RECT 62.700 144.200 63.000 144.800 ;
        RECT 63.800 144.400 64.200 145.200 ;
        RECT 62.600 143.800 63.000 144.200 ;
        RECT 64.600 141.100 65.000 145.800 ;
        RECT 67.800 145.500 68.100 146.500 ;
        RECT 66.200 145.200 68.100 145.500 ;
        RECT 66.200 143.500 66.500 145.200 ;
        RECT 68.800 144.900 69.100 146.800 ;
        RECT 69.400 146.100 69.800 146.200 ;
        RECT 70.200 146.100 70.600 146.200 ;
        RECT 69.400 145.800 70.600 146.100 ;
        RECT 71.000 145.800 71.400 146.600 ;
        RECT 71.800 145.800 72.200 146.600 ;
        RECT 72.600 146.500 73.300 146.900 ;
        RECT 73.600 146.800 74.600 147.200 ;
        RECT 69.400 145.400 69.800 145.800 ;
        RECT 72.600 145.500 72.900 146.500 ;
        RECT 68.300 144.600 69.100 144.900 ;
        RECT 71.000 145.200 72.900 145.500 ;
        RECT 66.200 141.500 66.600 143.500 ;
        RECT 68.300 142.200 68.700 144.600 ;
        RECT 67.800 141.800 68.700 142.200 ;
        RECT 68.300 141.100 68.700 141.800 ;
        RECT 71.000 143.500 71.300 145.200 ;
        RECT 73.600 144.900 73.900 146.800 ;
        RECT 74.200 145.400 74.600 146.200 ;
        RECT 75.800 145.700 76.200 147.400 ;
        RECT 79.300 147.100 79.700 147.200 ;
        RECT 80.600 147.100 81.000 147.200 ;
        RECT 82.200 147.100 82.500 148.200 ;
        RECT 84.600 147.500 85.000 149.900 ;
        RECT 85.400 147.800 85.800 148.600 ;
        RECT 83.800 147.100 84.600 147.200 ;
        RECT 79.100 146.800 84.600 147.100 ;
        RECT 78.200 146.400 78.600 146.500 ;
        RECT 76.700 146.100 78.600 146.400 ;
        RECT 76.700 146.000 77.100 146.100 ;
        RECT 77.500 145.700 77.900 145.800 ;
        RECT 75.800 145.400 77.900 145.700 ;
        RECT 73.100 144.600 73.900 144.900 ;
        RECT 71.000 141.500 71.400 143.500 ;
        RECT 73.100 142.200 73.500 144.600 ;
        RECT 73.100 141.800 73.800 142.200 ;
        RECT 73.100 141.100 73.500 141.800 ;
        RECT 75.800 141.100 76.200 145.400 ;
        RECT 79.100 145.200 79.400 146.800 ;
        RECT 82.700 146.700 83.100 146.800 ;
        RECT 82.200 146.200 82.600 146.300 ;
        RECT 83.500 146.200 83.900 146.300 ;
        RECT 81.400 145.900 83.900 146.200 ;
        RECT 86.200 146.100 86.600 149.900 ;
        RECT 88.900 148.000 89.300 149.500 ;
        RECT 91.000 148.500 91.400 149.500 ;
        RECT 88.500 147.700 89.300 148.000 ;
        RECT 88.500 147.500 88.900 147.700 ;
        RECT 88.500 147.200 88.800 147.500 ;
        RECT 91.100 147.400 91.400 148.500 ;
        RECT 91.800 147.800 92.200 148.600 ;
        RECT 87.000 147.100 87.400 147.200 ;
        RECT 87.800 147.100 88.800 147.200 ;
        RECT 87.000 146.800 88.800 147.100 ;
        RECT 89.300 147.100 91.400 147.400 ;
        RECT 89.300 146.900 89.800 147.100 ;
        RECT 87.800 146.100 88.200 146.200 ;
        RECT 81.400 145.800 81.800 145.900 ;
        RECT 86.200 145.800 88.200 146.100 ;
        RECT 82.200 145.500 85.000 145.600 ;
        RECT 82.100 145.400 85.000 145.500 ;
        RECT 78.200 144.900 79.400 145.200 ;
        RECT 80.100 145.300 85.000 145.400 ;
        RECT 80.100 145.100 82.500 145.300 ;
        RECT 78.200 144.400 78.500 144.900 ;
        RECT 77.800 144.000 78.500 144.400 ;
        RECT 79.300 144.500 79.700 144.600 ;
        RECT 80.100 144.500 80.400 145.100 ;
        RECT 79.300 144.200 80.400 144.500 ;
        RECT 80.700 144.500 83.400 144.800 ;
        RECT 80.700 144.400 81.100 144.500 ;
        RECT 83.000 144.400 83.400 144.500 ;
        RECT 79.900 143.700 80.300 143.800 ;
        RECT 81.300 143.700 81.700 143.800 ;
        RECT 78.200 143.100 78.600 143.500 ;
        RECT 79.900 143.400 81.700 143.700 ;
        RECT 80.300 143.100 80.600 143.400 ;
        RECT 83.000 143.100 83.400 143.500 ;
        RECT 77.900 141.100 78.500 143.100 ;
        RECT 80.200 141.100 80.600 143.100 ;
        RECT 82.400 142.800 83.400 143.100 ;
        RECT 82.400 141.100 82.800 142.800 ;
        RECT 84.600 141.100 85.000 145.300 ;
        RECT 86.200 141.100 86.600 145.800 ;
        RECT 87.800 145.400 88.200 145.800 ;
        RECT 88.500 144.900 88.800 146.800 ;
        RECT 89.100 146.500 89.800 146.900 ;
        RECT 89.500 145.500 89.800 146.500 ;
        RECT 90.200 145.800 90.600 146.600 ;
        RECT 91.000 146.100 91.400 146.600 ;
        RECT 91.800 146.100 92.200 146.200 ;
        RECT 91.000 145.800 92.200 146.100 ;
        RECT 92.600 146.100 93.000 149.900 ;
        RECT 95.300 148.000 95.700 149.500 ;
        RECT 97.400 148.500 97.800 149.500 ;
        RECT 98.800 149.200 99.200 149.900 ;
        RECT 98.200 148.800 99.200 149.200 ;
        RECT 94.900 147.700 95.700 148.000 ;
        RECT 94.900 147.500 95.300 147.700 ;
        RECT 94.900 147.200 95.200 147.500 ;
        RECT 97.500 147.400 97.800 148.500 ;
        RECT 94.200 146.800 95.200 147.200 ;
        RECT 95.700 147.100 97.800 147.400 ;
        RECT 98.800 147.100 99.200 148.800 ;
        RECT 95.700 146.900 96.200 147.100 ;
        RECT 94.200 146.100 94.600 146.200 ;
        RECT 92.600 145.800 94.600 146.100 ;
        RECT 89.500 145.200 91.400 145.500 ;
        RECT 88.500 144.600 89.300 144.900 ;
        RECT 88.900 141.100 89.300 144.600 ;
        RECT 91.100 143.500 91.400 145.200 ;
        RECT 91.000 141.500 91.400 143.500 ;
        RECT 92.600 141.100 93.000 145.800 ;
        RECT 94.200 145.400 94.600 145.800 ;
        RECT 94.900 144.900 95.200 146.800 ;
        RECT 95.500 146.500 96.200 146.900 ;
        RECT 98.300 146.900 99.200 147.100 ;
        RECT 103.200 147.100 103.600 149.900 ;
        RECT 108.000 147.100 108.400 149.900 ;
        RECT 109.400 147.500 109.800 149.900 ;
        RECT 111.600 149.200 112.000 149.900 ;
        RECT 111.000 148.900 112.000 149.200 ;
        RECT 113.800 148.900 114.200 149.900 ;
        RECT 115.900 149.200 116.500 149.900 ;
        RECT 115.800 148.900 116.500 149.200 ;
        RECT 111.000 148.500 111.400 148.900 ;
        RECT 113.800 148.600 114.100 148.900 ;
        RECT 111.800 148.200 112.200 148.600 ;
        RECT 112.700 148.300 114.100 148.600 ;
        RECT 115.800 148.500 116.200 148.900 ;
        RECT 112.700 148.200 113.100 148.300 ;
        RECT 109.800 147.100 110.600 147.200 ;
        RECT 111.900 147.100 112.200 148.200 ;
        RECT 116.700 147.700 117.100 147.800 ;
        RECT 118.200 147.700 118.600 149.900 ;
        RECT 119.100 148.200 119.500 148.600 ;
        RECT 119.000 147.800 119.400 148.200 ;
        RECT 119.800 147.900 120.200 149.900 ;
        RECT 116.700 147.400 118.600 147.700 ;
        RECT 114.700 147.100 115.100 147.200 ;
        RECT 103.200 146.900 104.100 147.100 ;
        RECT 108.000 146.900 108.900 147.100 ;
        RECT 98.300 146.800 99.100 146.900 ;
        RECT 103.300 146.800 104.100 146.900 ;
        RECT 108.100 146.800 108.900 146.900 ;
        RECT 109.800 146.800 115.300 147.100 ;
        RECT 95.900 145.500 96.200 146.500 ;
        RECT 96.600 145.800 97.000 146.600 ;
        RECT 97.400 145.800 97.800 146.600 ;
        RECT 95.900 145.200 97.800 145.500 ;
        RECT 98.300 145.200 98.600 146.800 ;
        RECT 99.400 145.800 100.200 146.200 ;
        RECT 102.200 145.800 103.000 146.200 ;
        RECT 94.900 144.600 95.700 144.900 ;
        RECT 95.300 142.200 95.700 144.600 ;
        RECT 97.500 143.500 97.800 145.200 ;
        RECT 98.200 144.800 98.600 145.200 ;
        RECT 100.600 145.100 101.000 145.600 ;
        RECT 101.400 145.100 101.800 145.600 ;
        RECT 100.600 144.800 101.800 145.100 ;
        RECT 103.800 145.200 104.100 146.800 ;
        RECT 107.000 145.800 107.800 146.200 ;
        RECT 103.800 144.800 104.200 145.200 ;
        RECT 106.200 144.800 106.600 145.600 ;
        RECT 108.600 145.200 108.900 146.800 ;
        RECT 111.300 146.700 111.700 146.800 ;
        RECT 110.500 146.200 110.900 146.300 ;
        RECT 110.500 145.900 113.000 146.200 ;
        RECT 112.600 145.800 113.000 145.900 ;
        RECT 109.400 145.500 112.200 145.600 ;
        RECT 109.400 145.400 112.300 145.500 ;
        RECT 109.400 145.300 114.300 145.400 ;
        RECT 108.600 144.800 109.000 145.200 ;
        RECT 95.300 141.800 96.200 142.200 ;
        RECT 95.300 141.100 95.700 141.800 ;
        RECT 97.400 141.500 97.800 143.500 ;
        RECT 98.300 143.500 98.600 144.800 ;
        RECT 99.000 143.800 99.400 144.600 ;
        RECT 102.200 143.800 102.600 144.200 ;
        RECT 103.000 143.800 103.400 144.600 ;
        RECT 102.200 143.500 102.500 143.800 ;
        RECT 103.800 143.500 104.100 144.800 ;
        RECT 107.800 143.800 108.200 144.600 ;
        RECT 108.600 143.500 108.900 144.800 ;
        RECT 98.300 143.200 100.100 143.500 ;
        RECT 98.300 143.100 98.600 143.200 ;
        RECT 98.200 141.100 98.600 143.100 ;
        RECT 99.800 143.100 100.100 143.200 ;
        RECT 102.200 143.200 104.100 143.500 ;
        RECT 99.800 141.100 100.200 143.100 ;
        RECT 102.200 141.100 102.600 143.200 ;
        RECT 103.800 143.100 104.100 143.200 ;
        RECT 107.100 143.200 108.900 143.500 ;
        RECT 107.100 143.100 107.400 143.200 ;
        RECT 103.800 141.100 104.200 143.100 ;
        RECT 107.000 141.100 107.400 143.100 ;
        RECT 108.600 143.100 108.900 143.200 ;
        RECT 108.600 141.100 109.000 143.100 ;
        RECT 109.400 141.100 109.800 145.300 ;
        RECT 111.900 145.100 114.300 145.300 ;
        RECT 111.000 144.500 113.700 144.800 ;
        RECT 111.000 144.400 111.400 144.500 ;
        RECT 113.300 144.400 113.700 144.500 ;
        RECT 114.000 144.500 114.300 145.100 ;
        RECT 115.000 145.200 115.300 146.800 ;
        RECT 115.800 146.400 116.200 146.500 ;
        RECT 115.800 146.100 117.700 146.400 ;
        RECT 117.300 146.000 117.700 146.100 ;
        RECT 116.500 145.700 116.900 145.800 ;
        RECT 118.200 145.700 118.600 147.400 ;
        RECT 119.900 146.200 120.200 147.900 ;
        RECT 122.200 147.700 122.600 149.900 ;
        RECT 124.300 149.200 124.900 149.900 ;
        RECT 124.300 148.900 125.000 149.200 ;
        RECT 126.600 148.900 127.000 149.900 ;
        RECT 128.800 149.200 129.200 149.900 ;
        RECT 128.800 148.900 129.800 149.200 ;
        RECT 124.600 148.500 125.000 148.900 ;
        RECT 126.700 148.600 127.000 148.900 ;
        RECT 126.700 148.300 128.100 148.600 ;
        RECT 127.700 148.200 128.100 148.300 ;
        RECT 128.600 148.200 129.000 148.600 ;
        RECT 129.400 148.500 129.800 148.900 ;
        RECT 123.700 147.700 124.100 147.800 ;
        RECT 122.200 147.400 124.100 147.700 ;
        RECT 120.600 146.400 121.000 147.200 ;
        RECT 119.000 146.100 119.400 146.200 ;
        RECT 119.800 146.100 120.200 146.200 ;
        RECT 121.400 146.100 121.800 146.200 ;
        RECT 119.000 145.800 120.200 146.100 ;
        RECT 121.000 145.800 121.800 146.100 ;
        RECT 116.500 145.400 118.600 145.700 ;
        RECT 115.000 144.900 116.200 145.200 ;
        RECT 114.700 144.500 115.100 144.600 ;
        RECT 114.000 144.200 115.100 144.500 ;
        RECT 115.900 144.400 116.200 144.900 ;
        RECT 115.900 144.000 116.600 144.400 ;
        RECT 112.700 143.700 113.100 143.800 ;
        RECT 114.100 143.700 114.500 143.800 ;
        RECT 111.000 143.100 111.400 143.500 ;
        RECT 112.700 143.400 114.500 143.700 ;
        RECT 113.800 143.100 114.100 143.400 ;
        RECT 115.800 143.100 116.200 143.500 ;
        RECT 111.000 142.800 112.000 143.100 ;
        RECT 111.600 141.100 112.000 142.800 ;
        RECT 113.800 141.100 114.200 143.100 ;
        RECT 115.900 141.100 116.500 143.100 ;
        RECT 118.200 141.100 118.600 145.400 ;
        RECT 119.100 145.100 119.400 145.800 ;
        RECT 121.000 145.600 121.400 145.800 ;
        RECT 122.200 145.700 122.600 147.400 ;
        RECT 125.700 147.100 126.100 147.200 ;
        RECT 127.000 147.100 127.400 147.200 ;
        RECT 128.600 147.100 128.900 148.200 ;
        RECT 131.000 147.500 131.400 149.900 ;
        RECT 132.100 148.200 132.500 149.900 ;
        RECT 132.100 147.900 133.000 148.200 ;
        RECT 130.200 147.100 131.000 147.200 ;
        RECT 125.500 146.800 131.000 147.100 ;
        RECT 131.800 147.100 132.200 147.200 ;
        RECT 132.600 147.100 133.000 147.900 ;
        RECT 131.800 146.800 133.000 147.100 ;
        RECT 133.400 146.800 133.800 147.600 ;
        RECT 124.600 146.400 125.000 146.500 ;
        RECT 123.100 146.100 125.000 146.400 ;
        RECT 123.100 146.000 123.500 146.100 ;
        RECT 123.900 145.700 124.300 145.800 ;
        RECT 122.200 145.400 124.300 145.700 ;
        RECT 119.000 141.100 119.400 145.100 ;
        RECT 119.800 144.800 121.800 145.100 ;
        RECT 119.800 141.100 120.200 144.800 ;
        RECT 121.400 141.100 121.800 144.800 ;
        RECT 122.200 141.100 122.600 145.400 ;
        RECT 125.500 145.200 125.800 146.800 ;
        RECT 129.100 146.700 129.500 146.800 ;
        RECT 129.900 146.200 130.300 146.300 ;
        RECT 127.000 146.100 127.400 146.200 ;
        RECT 127.800 146.100 130.300 146.200 ;
        RECT 127.000 145.900 130.300 146.100 ;
        RECT 127.000 145.800 128.200 145.900 ;
        RECT 128.600 145.500 131.400 145.600 ;
        RECT 128.500 145.400 131.400 145.500 ;
        RECT 124.600 144.900 125.800 145.200 ;
        RECT 126.500 145.300 131.400 145.400 ;
        RECT 126.500 145.100 128.900 145.300 ;
        RECT 124.600 144.400 124.900 144.900 ;
        RECT 124.200 144.000 124.900 144.400 ;
        RECT 125.700 144.500 126.100 144.600 ;
        RECT 126.500 144.500 126.800 145.100 ;
        RECT 125.700 144.200 126.800 144.500 ;
        RECT 127.100 144.500 129.800 144.800 ;
        RECT 127.100 144.400 127.500 144.500 ;
        RECT 129.400 144.400 129.800 144.500 ;
        RECT 126.300 143.700 126.700 143.800 ;
        RECT 127.700 143.700 128.100 143.800 ;
        RECT 124.600 143.100 125.000 143.500 ;
        RECT 126.300 143.400 128.100 143.700 ;
        RECT 126.700 143.100 127.000 143.400 ;
        RECT 129.400 143.100 129.800 143.500 ;
        RECT 124.300 141.100 124.900 143.100 ;
        RECT 126.600 141.100 127.000 143.100 ;
        RECT 128.800 142.800 129.800 143.100 ;
        RECT 128.800 141.100 129.200 142.800 ;
        RECT 131.000 141.100 131.400 145.300 ;
        RECT 131.800 144.400 132.200 145.200 ;
        RECT 132.600 141.100 133.000 146.800 ;
        RECT 134.200 146.100 134.600 149.900 ;
        RECT 136.600 148.800 137.000 149.900 ;
        RECT 135.800 147.800 136.200 148.600 ;
        RECT 135.000 147.100 135.400 147.600 ;
        RECT 135.800 147.100 136.100 147.800 ;
        RECT 136.700 147.200 137.000 148.800 ;
        RECT 138.200 147.600 138.600 149.900 ;
        RECT 139.800 148.200 140.200 149.900 ;
        RECT 139.800 147.900 140.300 148.200 ;
        RECT 138.200 147.300 139.500 147.600 ;
        RECT 135.000 146.800 136.100 147.100 ;
        RECT 136.600 146.800 137.000 147.200 ;
        RECT 135.000 146.100 135.400 146.200 ;
        RECT 134.200 145.800 135.400 146.100 ;
        RECT 134.200 141.100 134.600 145.800 ;
        RECT 136.700 145.100 137.000 146.800 ;
        RECT 138.300 146.200 138.700 146.600 ;
        RECT 137.400 145.400 137.800 146.200 ;
        RECT 138.200 145.800 138.700 146.200 ;
        RECT 139.200 146.500 139.500 147.300 ;
        RECT 140.000 147.200 140.300 147.900 ;
        RECT 139.800 146.800 140.300 147.200 ;
        RECT 142.000 147.100 142.400 149.900 ;
        RECT 139.200 146.100 139.700 146.500 ;
        RECT 139.200 145.100 139.500 146.100 ;
        RECT 140.000 145.100 140.300 146.800 ;
        RECT 141.500 146.900 142.400 147.100 ;
        RECT 146.400 147.100 146.800 149.900 ;
        RECT 149.600 147.100 150.000 149.900 ;
        RECT 151.000 147.600 151.400 149.900 ;
        RECT 152.600 148.200 153.000 149.900 ;
        RECT 155.500 149.100 155.900 149.900 ;
        RECT 159.500 149.200 159.900 149.900 ;
        RECT 157.400 149.100 157.800 149.200 ;
        RECT 155.500 148.800 157.800 149.100 ;
        RECT 159.500 148.800 160.200 149.200 ;
        RECT 155.500 148.200 155.900 148.800 ;
        RECT 159.500 148.200 159.900 148.800 ;
        RECT 152.600 147.900 153.100 148.200 ;
        RECT 151.000 147.300 152.300 147.600 ;
        RECT 146.400 146.900 147.300 147.100 ;
        RECT 149.600 146.900 150.500 147.100 ;
        RECT 141.500 146.800 142.300 146.900 ;
        RECT 146.500 146.800 147.300 146.900 ;
        RECT 149.700 146.800 150.500 146.900 ;
        RECT 141.500 145.200 141.800 146.800 ;
        RECT 142.600 145.800 143.400 146.200 ;
        RECT 145.400 145.800 146.200 146.200 ;
        RECT 136.600 144.700 137.500 145.100 ;
        RECT 137.100 141.100 137.500 144.700 ;
        RECT 138.200 144.800 139.500 145.100 ;
        RECT 138.200 141.100 138.600 144.800 ;
        RECT 139.800 144.600 140.300 145.100 ;
        RECT 141.400 144.800 141.800 145.200 ;
        RECT 143.800 145.100 144.200 145.600 ;
        RECT 144.600 145.100 145.000 145.600 ;
        RECT 143.800 144.800 145.000 145.100 ;
        RECT 147.000 145.200 147.300 146.800 ;
        RECT 148.600 145.800 149.400 146.200 ;
        RECT 147.000 144.800 147.400 145.200 ;
        RECT 147.800 144.800 148.200 145.600 ;
        RECT 150.200 145.200 150.500 146.800 ;
        RECT 151.100 146.200 151.500 146.600 ;
        RECT 151.000 145.800 151.500 146.200 ;
        RECT 152.000 146.500 152.300 147.300 ;
        RECT 152.800 147.200 153.100 147.900 ;
        RECT 155.000 147.900 155.900 148.200 ;
        RECT 159.000 147.900 159.900 148.200 ;
        RECT 152.600 146.800 153.100 147.200 ;
        RECT 154.200 146.800 154.600 147.600 ;
        RECT 152.000 146.100 152.500 146.500 ;
        RECT 139.800 141.100 140.200 144.600 ;
        RECT 141.500 143.500 141.800 144.800 ;
        RECT 142.200 144.100 142.600 144.600 ;
        RECT 143.000 144.100 143.400 144.200 ;
        RECT 146.200 144.100 146.600 144.600 ;
        RECT 142.200 143.800 146.600 144.100 ;
        RECT 147.000 143.500 147.300 144.800 ;
        RECT 149.400 143.800 149.800 145.200 ;
        RECT 150.200 144.800 150.600 145.200 ;
        RECT 152.000 145.100 152.300 146.100 ;
        RECT 152.800 145.100 153.100 146.800 ;
        RECT 151.000 144.800 152.300 145.100 ;
        RECT 150.200 143.500 150.500 144.800 ;
        RECT 141.500 143.200 143.300 143.500 ;
        RECT 141.500 143.100 141.800 143.200 ;
        RECT 141.400 141.100 141.800 143.100 ;
        RECT 143.000 143.100 143.300 143.200 ;
        RECT 145.500 143.200 147.300 143.500 ;
        RECT 145.500 143.100 145.800 143.200 ;
        RECT 143.000 141.100 143.400 143.100 ;
        RECT 145.400 141.100 145.800 143.100 ;
        RECT 147.000 143.100 147.300 143.200 ;
        RECT 148.700 143.200 150.500 143.500 ;
        RECT 148.700 143.100 149.000 143.200 ;
        RECT 147.000 141.100 147.400 143.100 ;
        RECT 148.600 141.100 149.000 143.100 ;
        RECT 150.200 143.100 150.500 143.200 ;
        RECT 150.200 141.100 150.600 143.100 ;
        RECT 151.000 141.100 151.400 144.800 ;
        RECT 152.600 144.600 153.100 145.100 ;
        RECT 152.600 141.100 153.000 144.600 ;
        RECT 155.000 141.100 155.400 147.900 ;
        RECT 158.200 146.800 158.600 147.600 ;
        RECT 155.800 145.100 156.200 145.200 ;
        RECT 158.200 145.100 158.600 145.200 ;
        RECT 155.800 144.800 158.600 145.100 ;
        RECT 155.800 144.400 156.200 144.800 ;
        RECT 159.000 141.100 159.400 147.900 ;
        RECT 161.200 147.100 161.600 149.900 ;
        RECT 160.700 146.900 161.600 147.100 ;
        RECT 164.600 147.600 165.000 149.900 ;
        RECT 166.200 147.600 166.600 149.900 ;
        RECT 167.800 147.700 168.200 149.900 ;
        RECT 169.900 149.200 170.500 149.900 ;
        RECT 169.900 148.900 170.600 149.200 ;
        RECT 172.200 148.900 172.600 149.900 ;
        RECT 174.400 149.200 174.800 149.900 ;
        RECT 174.400 148.900 175.400 149.200 ;
        RECT 170.200 148.500 170.600 148.900 ;
        RECT 172.300 148.600 172.600 148.900 ;
        RECT 172.300 148.300 173.700 148.600 ;
        RECT 173.300 148.200 173.700 148.300 ;
        RECT 174.200 148.200 174.600 148.600 ;
        RECT 175.000 148.500 175.400 148.900 ;
        RECT 169.300 147.700 169.700 147.800 ;
        RECT 164.600 147.200 166.600 147.600 ;
        RECT 160.700 146.800 161.500 146.900 ;
        RECT 160.700 145.200 161.000 146.800 ;
        RECT 161.400 145.800 162.600 146.200 ;
        RECT 164.600 145.800 165.000 147.200 ;
        RECT 167.000 146.800 167.400 147.600 ;
        RECT 167.800 147.400 169.700 147.700 ;
        RECT 159.800 144.400 160.200 145.200 ;
        RECT 160.600 144.800 161.000 145.200 ;
        RECT 163.000 144.800 163.400 145.600 ;
        RECT 164.600 145.400 166.600 145.800 ;
        RECT 160.700 143.500 161.000 144.800 ;
        RECT 161.400 143.800 161.800 144.600 ;
        RECT 160.700 143.200 162.500 143.500 ;
        RECT 160.700 143.100 161.000 143.200 ;
        RECT 160.600 141.100 161.000 143.100 ;
        RECT 162.200 141.100 162.600 143.200 ;
        RECT 164.600 141.100 165.000 145.400 ;
        RECT 166.200 141.100 166.600 145.400 ;
        RECT 167.800 145.700 168.200 147.400 ;
        RECT 174.200 147.200 174.500 148.200 ;
        RECT 176.600 147.500 177.000 149.900 ;
        RECT 177.400 148.500 177.800 149.500 ;
        RECT 177.400 147.400 177.700 148.500 ;
        RECT 179.500 148.000 179.900 149.500 ;
        RECT 179.500 147.700 180.300 148.000 ;
        RECT 179.900 147.500 180.300 147.700 ;
        RECT 171.300 147.100 171.700 147.200 ;
        RECT 174.200 147.100 174.600 147.200 ;
        RECT 175.800 147.100 176.600 147.200 ;
        RECT 177.400 147.100 179.500 147.400 ;
        RECT 171.100 146.800 176.600 147.100 ;
        RECT 179.000 146.900 179.500 147.100 ;
        RECT 180.000 147.200 180.300 147.500 ;
        RECT 170.200 146.400 170.600 146.500 ;
        RECT 168.700 146.100 170.600 146.400 ;
        RECT 168.700 146.000 169.100 146.100 ;
        RECT 169.500 145.700 169.900 145.800 ;
        RECT 167.800 145.400 169.900 145.700 ;
        RECT 167.800 141.100 168.200 145.400 ;
        RECT 171.100 145.200 171.400 146.800 ;
        RECT 174.700 146.700 175.100 146.800 ;
        RECT 175.500 146.200 175.900 146.300 ;
        RECT 173.400 145.900 175.900 146.200 ;
        RECT 173.400 145.800 173.800 145.900 ;
        RECT 177.400 145.800 177.800 146.600 ;
        RECT 178.200 145.800 178.600 146.600 ;
        RECT 179.000 146.500 179.700 146.900 ;
        RECT 180.000 146.800 181.000 147.200 ;
        RECT 174.200 145.500 177.000 145.600 ;
        RECT 179.000 145.500 179.300 146.500 ;
        RECT 174.100 145.400 177.000 145.500 ;
        RECT 170.200 144.900 171.400 145.200 ;
        RECT 172.100 145.300 177.000 145.400 ;
        RECT 172.100 145.100 174.500 145.300 ;
        RECT 170.200 144.400 170.500 144.900 ;
        RECT 169.800 144.000 170.500 144.400 ;
        RECT 171.300 144.500 171.700 144.600 ;
        RECT 172.100 144.500 172.400 145.100 ;
        RECT 171.300 144.200 172.400 144.500 ;
        RECT 172.700 144.500 175.400 144.800 ;
        RECT 172.700 144.400 173.100 144.500 ;
        RECT 175.000 144.400 175.400 144.500 ;
        RECT 171.900 143.700 172.300 143.800 ;
        RECT 173.300 143.700 173.700 143.800 ;
        RECT 170.200 143.100 170.600 143.500 ;
        RECT 171.900 143.400 173.700 143.700 ;
        RECT 172.300 143.100 172.600 143.400 ;
        RECT 175.000 143.100 175.400 143.500 ;
        RECT 169.900 141.100 170.500 143.100 ;
        RECT 172.200 141.100 172.600 143.100 ;
        RECT 174.400 142.800 175.400 143.100 ;
        RECT 174.400 141.100 174.800 142.800 ;
        RECT 176.600 141.100 177.000 145.300 ;
        RECT 177.400 145.200 179.300 145.500 ;
        RECT 177.400 143.500 177.700 145.200 ;
        RECT 180.000 144.900 180.300 146.800 ;
        RECT 180.600 146.100 181.000 146.200 ;
        RECT 182.200 146.100 182.600 149.900 ;
        RECT 183.000 147.800 183.400 148.600 ;
        RECT 183.800 147.600 184.200 149.900 ;
        RECT 185.400 148.200 185.800 149.900 ;
        RECT 185.400 147.900 185.900 148.200 ;
        RECT 183.800 147.300 185.100 147.600 ;
        RECT 183.900 146.200 184.300 146.600 ;
        RECT 180.600 145.800 182.600 146.100 ;
        RECT 183.800 145.800 184.300 146.200 ;
        RECT 184.800 146.500 185.100 147.300 ;
        RECT 185.600 147.200 185.900 147.900 ;
        RECT 185.400 146.800 185.900 147.200 ;
        RECT 184.800 146.100 185.300 146.500 ;
        RECT 180.600 145.400 181.000 145.800 ;
        RECT 179.500 144.600 180.300 144.900 ;
        RECT 177.400 141.500 177.800 143.500 ;
        RECT 179.500 142.200 179.900 144.600 ;
        RECT 179.500 141.800 180.200 142.200 ;
        RECT 179.500 141.100 179.900 141.800 ;
        RECT 182.200 141.100 182.600 145.800 ;
        RECT 184.800 145.100 185.100 146.100 ;
        RECT 185.600 145.100 185.900 146.800 ;
        RECT 183.800 144.800 185.100 145.100 ;
        RECT 183.800 141.100 184.200 144.800 ;
        RECT 185.400 144.600 185.900 145.100 ;
        RECT 187.000 147.700 187.400 149.900 ;
        RECT 189.100 149.200 189.700 149.900 ;
        RECT 189.100 148.900 189.800 149.200 ;
        RECT 191.400 148.900 191.800 149.900 ;
        RECT 193.600 149.200 194.000 149.900 ;
        RECT 193.600 148.900 194.600 149.200 ;
        RECT 189.400 148.500 189.800 148.900 ;
        RECT 191.500 148.600 191.800 148.900 ;
        RECT 191.500 148.300 192.900 148.600 ;
        RECT 192.500 148.200 192.900 148.300 ;
        RECT 193.400 148.200 193.800 148.600 ;
        RECT 194.200 148.500 194.600 148.900 ;
        RECT 188.500 147.700 188.900 147.800 ;
        RECT 187.000 147.400 188.900 147.700 ;
        RECT 187.000 145.700 187.400 147.400 ;
        RECT 190.500 147.100 190.900 147.200 ;
        RECT 191.800 147.100 192.200 147.200 ;
        RECT 193.400 147.100 193.700 148.200 ;
        RECT 195.800 147.500 196.200 149.900 ;
        RECT 198.500 148.000 198.900 149.500 ;
        RECT 200.600 148.500 201.000 149.500 ;
        RECT 198.100 147.700 198.900 148.000 ;
        RECT 198.100 147.500 198.500 147.700 ;
        RECT 198.100 147.200 198.400 147.500 ;
        RECT 200.700 147.400 201.000 148.500 ;
        RECT 201.400 148.000 201.800 149.900 ;
        RECT 203.000 148.000 203.400 149.900 ;
        RECT 201.400 147.900 203.400 148.000 ;
        RECT 203.800 147.900 204.200 149.900 ;
        RECT 204.600 147.900 205.000 149.900 ;
        RECT 205.400 148.000 205.800 149.900 ;
        RECT 207.000 148.000 207.400 149.900 ;
        RECT 205.400 147.900 207.400 148.000 ;
        RECT 201.500 147.700 203.300 147.900 ;
        RECT 195.000 147.100 195.800 147.200 ;
        RECT 190.300 146.800 195.800 147.100 ;
        RECT 197.400 146.800 198.400 147.200 ;
        RECT 198.900 147.100 201.000 147.400 ;
        RECT 201.800 147.200 202.200 147.400 ;
        RECT 203.800 147.200 204.100 147.900 ;
        RECT 204.700 147.200 205.000 147.900 ;
        RECT 205.500 147.700 207.300 147.900 ;
        RECT 209.400 147.700 209.800 149.900 ;
        RECT 211.500 149.200 212.100 149.900 ;
        RECT 211.500 148.900 212.200 149.200 ;
        RECT 213.800 148.900 214.200 149.900 ;
        RECT 216.000 149.200 216.400 149.900 ;
        RECT 216.000 148.900 217.000 149.200 ;
        RECT 211.800 148.500 212.200 148.900 ;
        RECT 213.900 148.600 214.200 148.900 ;
        RECT 213.900 148.300 215.300 148.600 ;
        RECT 214.900 148.200 215.300 148.300 ;
        RECT 215.800 148.200 216.200 148.600 ;
        RECT 216.600 148.500 217.000 148.900 ;
        RECT 210.900 147.700 211.300 147.800 ;
        RECT 209.400 147.400 211.300 147.700 ;
        RECT 206.600 147.200 207.000 147.400 ;
        RECT 198.900 146.900 199.400 147.100 ;
        RECT 189.400 146.400 189.800 146.500 ;
        RECT 187.900 146.100 189.800 146.400 ;
        RECT 187.900 146.000 188.300 146.100 ;
        RECT 188.700 145.700 189.100 145.800 ;
        RECT 187.000 145.400 189.100 145.700 ;
        RECT 185.400 141.100 185.800 144.600 ;
        RECT 187.000 141.100 187.400 145.400 ;
        RECT 190.300 145.200 190.600 146.800 ;
        RECT 193.900 146.700 194.300 146.800 ;
        RECT 193.400 146.200 193.800 146.300 ;
        RECT 194.700 146.200 195.100 146.300 ;
        RECT 192.600 145.900 195.100 146.200 ;
        RECT 192.600 145.800 193.000 145.900 ;
        RECT 193.400 145.500 196.200 145.600 ;
        RECT 193.300 145.400 196.200 145.500 ;
        RECT 197.400 145.400 197.800 146.200 ;
        RECT 189.400 144.900 190.600 145.200 ;
        RECT 191.300 145.300 196.200 145.400 ;
        RECT 191.300 145.100 193.700 145.300 ;
        RECT 189.400 144.400 189.700 144.900 ;
        RECT 189.000 144.000 189.700 144.400 ;
        RECT 190.500 144.500 190.900 144.600 ;
        RECT 191.300 144.500 191.600 145.100 ;
        RECT 190.500 144.200 191.600 144.500 ;
        RECT 191.900 144.500 194.600 144.800 ;
        RECT 191.900 144.400 192.300 144.500 ;
        RECT 194.200 144.400 194.600 144.500 ;
        RECT 191.100 143.700 191.500 143.800 ;
        RECT 192.500 143.700 192.900 143.800 ;
        RECT 189.400 143.100 189.800 143.500 ;
        RECT 191.100 143.400 192.900 143.700 ;
        RECT 191.500 143.100 191.800 143.400 ;
        RECT 194.200 143.100 194.600 143.500 ;
        RECT 189.100 141.100 189.700 143.100 ;
        RECT 191.400 141.100 191.800 143.100 ;
        RECT 193.600 142.800 194.600 143.100 ;
        RECT 193.600 141.100 194.000 142.800 ;
        RECT 195.800 141.100 196.200 145.300 ;
        RECT 198.100 144.900 198.400 146.800 ;
        RECT 198.700 146.500 199.400 146.900 ;
        RECT 201.400 146.900 202.200 147.200 ;
        RECT 201.400 146.800 201.800 146.900 ;
        RECT 202.900 146.800 204.200 147.200 ;
        RECT 204.600 146.800 205.900 147.200 ;
        RECT 206.600 146.900 207.400 147.200 ;
        RECT 207.000 146.800 207.400 146.900 ;
        RECT 199.100 145.500 199.400 146.500 ;
        RECT 199.800 145.800 200.200 146.600 ;
        RECT 200.600 145.800 201.000 146.600 ;
        RECT 202.200 145.800 202.600 146.600 ;
        RECT 202.900 146.200 203.200 146.800 ;
        RECT 202.900 145.800 203.400 146.200 ;
        RECT 203.800 145.800 204.200 146.200 ;
        RECT 199.100 145.200 201.000 145.500 ;
        RECT 198.100 144.600 198.900 144.900 ;
        RECT 198.500 142.200 198.900 144.600 ;
        RECT 200.700 143.500 201.000 145.200 ;
        RECT 202.900 145.100 203.200 145.800 ;
        RECT 203.800 145.200 204.100 145.800 ;
        RECT 203.800 145.100 204.200 145.200 ;
        RECT 198.200 141.800 198.900 142.200 ;
        RECT 198.500 141.100 198.900 141.800 ;
        RECT 200.600 141.500 201.000 143.500 ;
        RECT 202.700 144.800 203.200 145.100 ;
        RECT 203.500 144.800 204.200 145.100 ;
        RECT 204.600 145.100 205.000 145.200 ;
        RECT 205.600 145.100 205.900 146.800 ;
        RECT 206.200 145.800 206.600 146.600 ;
        RECT 209.400 145.700 209.800 147.400 ;
        RECT 212.900 147.100 213.300 147.200 ;
        RECT 215.800 147.100 216.100 148.200 ;
        RECT 218.200 147.500 218.600 149.900 ;
        RECT 219.000 147.600 219.400 149.900 ;
        RECT 220.600 148.200 221.000 149.900 ;
        RECT 220.600 147.900 221.100 148.200 ;
        RECT 224.100 148.000 224.500 149.500 ;
        RECT 226.200 148.500 226.600 149.500 ;
        RECT 219.000 147.300 220.300 147.600 ;
        RECT 217.400 147.100 218.200 147.200 ;
        RECT 212.700 146.800 218.200 147.100 ;
        RECT 211.800 146.400 212.200 146.500 ;
        RECT 210.300 146.100 212.200 146.400 ;
        RECT 210.300 146.000 210.700 146.100 ;
        RECT 211.100 145.700 211.500 145.800 ;
        RECT 209.400 145.400 211.500 145.700 ;
        RECT 204.600 144.800 205.300 145.100 ;
        RECT 205.600 144.800 206.100 145.100 ;
        RECT 202.700 141.100 203.100 144.800 ;
        RECT 203.500 144.200 203.800 144.800 ;
        RECT 203.400 143.800 203.800 144.200 ;
        RECT 205.000 144.200 205.300 144.800 ;
        RECT 205.000 143.800 205.400 144.200 ;
        RECT 205.700 141.100 206.100 144.800 ;
        RECT 209.400 141.100 209.800 145.400 ;
        RECT 212.700 145.200 213.000 146.800 ;
        RECT 216.300 146.700 216.700 146.800 ;
        RECT 217.100 146.200 217.500 146.300 ;
        RECT 219.100 146.200 219.500 146.600 ;
        RECT 215.000 145.900 217.500 146.200 ;
        RECT 215.000 145.800 215.400 145.900 ;
        RECT 219.000 145.800 219.500 146.200 ;
        RECT 220.000 146.500 220.300 147.300 ;
        RECT 220.800 147.200 221.100 147.900 ;
        RECT 223.700 147.700 224.500 148.000 ;
        RECT 223.700 147.500 224.100 147.700 ;
        RECT 223.700 147.200 224.000 147.500 ;
        RECT 226.300 147.400 226.600 148.500 ;
        RECT 228.300 148.200 228.700 149.900 ;
        RECT 227.800 147.900 228.700 148.200 ;
        RECT 229.400 147.900 229.800 149.900 ;
        RECT 230.200 148.000 230.600 149.900 ;
        RECT 231.800 148.000 232.200 149.900 ;
        RECT 230.200 147.900 232.200 148.000 ;
        RECT 220.600 146.800 221.100 147.200 ;
        RECT 223.000 146.800 224.000 147.200 ;
        RECT 224.500 147.100 226.600 147.400 ;
        RECT 224.500 146.900 225.000 147.100 ;
        RECT 220.000 146.100 220.500 146.500 ;
        RECT 215.800 145.500 218.600 145.600 ;
        RECT 215.700 145.400 218.600 145.500 ;
        RECT 211.800 144.900 213.000 145.200 ;
        RECT 213.700 145.300 218.600 145.400 ;
        RECT 213.700 145.100 216.100 145.300 ;
        RECT 211.800 144.400 212.100 144.900 ;
        RECT 211.400 144.000 212.100 144.400 ;
        RECT 212.900 144.500 213.300 144.600 ;
        RECT 213.700 144.500 214.000 145.100 ;
        RECT 212.900 144.200 214.000 144.500 ;
        RECT 214.300 144.500 217.000 144.800 ;
        RECT 214.300 144.400 214.700 144.500 ;
        RECT 216.600 144.400 217.000 144.500 ;
        RECT 213.500 143.700 213.900 143.800 ;
        RECT 214.900 143.700 215.300 143.800 ;
        RECT 211.800 143.100 212.200 143.500 ;
        RECT 213.500 143.400 215.300 143.700 ;
        RECT 213.900 143.100 214.200 143.400 ;
        RECT 216.600 143.100 217.000 143.500 ;
        RECT 211.500 141.100 212.100 143.100 ;
        RECT 213.800 141.100 214.200 143.100 ;
        RECT 216.000 142.800 217.000 143.100 ;
        RECT 216.000 141.100 216.400 142.800 ;
        RECT 218.200 141.100 218.600 145.300 ;
        RECT 220.000 145.100 220.300 146.100 ;
        RECT 220.800 145.100 221.100 146.800 ;
        RECT 223.000 145.400 223.400 146.200 ;
        RECT 219.000 144.800 220.300 145.100 ;
        RECT 219.000 141.100 219.400 144.800 ;
        RECT 220.600 144.600 221.100 145.100 ;
        RECT 223.700 144.900 224.000 146.800 ;
        RECT 224.300 146.500 225.000 146.900 ;
        RECT 227.000 146.800 227.400 147.600 ;
        RECT 224.700 145.500 225.000 146.500 ;
        RECT 225.400 145.800 225.800 146.600 ;
        RECT 226.200 145.800 226.600 146.600 ;
        RECT 227.800 146.100 228.200 147.900 ;
        RECT 229.500 147.200 229.800 147.900 ;
        RECT 230.300 147.700 232.100 147.900 ;
        RECT 232.600 147.500 233.000 149.900 ;
        RECT 234.800 149.200 235.200 149.900 ;
        RECT 234.200 148.900 235.200 149.200 ;
        RECT 237.000 148.900 237.400 149.900 ;
        RECT 239.100 149.200 239.700 149.900 ;
        RECT 239.000 148.900 239.700 149.200 ;
        RECT 234.200 148.500 234.600 148.900 ;
        RECT 237.000 148.600 237.300 148.900 ;
        RECT 235.000 148.200 235.400 148.600 ;
        RECT 235.900 148.300 237.300 148.600 ;
        RECT 239.000 148.500 239.400 148.900 ;
        RECT 235.900 148.200 236.300 148.300 ;
        RECT 231.400 147.200 231.800 147.400 ;
        RECT 229.400 146.800 230.700 147.200 ;
        RECT 231.400 146.900 232.200 147.200 ;
        RECT 231.800 146.800 232.200 146.900 ;
        RECT 233.000 147.100 233.800 147.200 ;
        RECT 235.100 147.100 235.400 148.200 ;
        RECT 239.900 147.700 240.300 147.800 ;
        RECT 241.400 147.700 241.800 149.900 ;
        RECT 242.200 148.000 242.600 149.900 ;
        RECT 243.800 148.000 244.200 149.900 ;
        RECT 242.200 147.900 244.200 148.000 ;
        RECT 244.600 147.900 245.000 149.900 ;
        RECT 245.700 148.200 246.100 149.900 ;
        RECT 249.100 148.200 249.500 149.900 ;
        RECT 245.700 147.900 246.600 148.200 ;
        RECT 242.300 147.700 244.100 147.900 ;
        RECT 239.900 147.400 241.800 147.700 ;
        RECT 237.900 147.100 238.300 147.200 ;
        RECT 233.000 146.800 238.500 147.100 ;
        RECT 230.400 146.200 230.700 146.800 ;
        RECT 234.500 146.700 234.900 146.800 ;
        RECT 227.800 145.800 229.700 146.100 ;
        RECT 230.200 145.800 230.700 146.200 ;
        RECT 231.000 145.800 231.400 146.600 ;
        RECT 233.700 146.200 234.100 146.300 ;
        RECT 233.700 145.900 236.200 146.200 ;
        RECT 235.800 145.800 236.200 145.900 ;
        RECT 224.700 145.200 226.600 145.500 ;
        RECT 223.700 144.600 224.500 144.900 ;
        RECT 220.600 141.100 221.000 144.600 ;
        RECT 224.100 141.100 224.500 144.600 ;
        RECT 226.300 143.500 226.600 145.200 ;
        RECT 226.200 141.500 226.600 143.500 ;
        RECT 227.800 141.100 228.200 145.800 ;
        RECT 229.400 145.200 229.700 145.800 ;
        RECT 228.600 144.400 229.000 145.200 ;
        RECT 229.400 145.100 229.800 145.200 ;
        RECT 230.400 145.100 230.700 145.800 ;
        RECT 232.600 145.500 235.400 145.600 ;
        RECT 232.600 145.400 235.500 145.500 ;
        RECT 232.600 145.300 237.500 145.400 ;
        RECT 229.400 144.800 230.100 145.100 ;
        RECT 230.400 144.800 230.900 145.100 ;
        RECT 229.800 144.200 230.100 144.800 ;
        RECT 229.800 143.800 230.200 144.200 ;
        RECT 230.500 141.100 230.900 144.800 ;
        RECT 232.600 141.100 233.000 145.300 ;
        RECT 235.100 145.100 237.500 145.300 ;
        RECT 234.200 144.500 236.900 144.800 ;
        RECT 234.200 144.400 234.600 144.500 ;
        RECT 236.500 144.400 236.900 144.500 ;
        RECT 237.200 144.500 237.500 145.100 ;
        RECT 238.200 145.200 238.500 146.800 ;
        RECT 239.000 146.400 239.400 146.500 ;
        RECT 239.000 146.100 240.900 146.400 ;
        RECT 240.500 146.000 240.900 146.100 ;
        RECT 239.700 145.700 240.100 145.800 ;
        RECT 241.400 145.700 241.800 147.400 ;
        RECT 242.600 147.200 243.000 147.400 ;
        RECT 244.600 147.200 244.900 147.900 ;
        RECT 242.200 146.900 243.000 147.200 ;
        RECT 243.700 147.100 245.000 147.200 ;
        RECT 245.400 147.100 245.800 147.200 ;
        RECT 242.200 146.800 242.600 146.900 ;
        RECT 243.700 146.800 245.800 147.100 ;
        RECT 243.000 145.800 243.400 146.600 ;
        RECT 239.700 145.400 241.800 145.700 ;
        RECT 238.200 144.900 239.400 145.200 ;
        RECT 237.900 144.500 238.300 144.600 ;
        RECT 237.200 144.200 238.300 144.500 ;
        RECT 239.100 144.400 239.400 144.900 ;
        RECT 239.100 144.000 239.800 144.400 ;
        RECT 235.900 143.700 236.300 143.800 ;
        RECT 237.300 143.700 237.700 143.800 ;
        RECT 234.200 143.100 234.600 143.500 ;
        RECT 235.900 143.400 237.700 143.700 ;
        RECT 237.000 143.100 237.300 143.400 ;
        RECT 239.000 143.100 239.400 143.500 ;
        RECT 234.200 142.800 235.200 143.100 ;
        RECT 234.800 141.100 235.200 142.800 ;
        RECT 237.000 141.100 237.400 143.100 ;
        RECT 239.100 141.100 239.700 143.100 ;
        RECT 241.400 141.100 241.800 145.400 ;
        RECT 243.700 145.100 244.000 146.800 ;
        RECT 246.200 146.100 246.600 147.900 ;
        RECT 248.600 147.900 249.500 148.200 ;
        RECT 247.000 146.800 247.400 147.600 ;
        RECT 244.600 145.800 246.600 146.100 ;
        RECT 244.600 145.200 244.900 145.800 ;
        RECT 244.600 145.100 245.000 145.200 ;
        RECT 243.500 144.800 244.000 145.100 ;
        RECT 244.300 144.800 245.000 145.100 ;
        RECT 243.500 141.100 243.900 144.800 ;
        RECT 244.300 144.200 244.600 144.800 ;
        RECT 245.400 144.400 245.800 145.200 ;
        RECT 244.200 143.800 244.600 144.200 ;
        RECT 246.200 141.100 246.600 145.800 ;
        RECT 248.600 141.100 249.000 147.900 ;
        RECT 250.200 147.700 250.600 149.900 ;
        RECT 252.300 149.200 252.900 149.900 ;
        RECT 252.300 148.900 253.000 149.200 ;
        RECT 254.600 148.900 255.000 149.900 ;
        RECT 256.800 149.200 257.200 149.900 ;
        RECT 256.800 148.900 257.800 149.200 ;
        RECT 252.600 148.500 253.000 148.900 ;
        RECT 254.700 148.600 255.000 148.900 ;
        RECT 254.700 148.300 256.100 148.600 ;
        RECT 255.700 148.200 256.100 148.300 ;
        RECT 256.600 148.200 257.000 148.600 ;
        RECT 257.400 148.500 257.800 148.900 ;
        RECT 251.700 147.700 252.100 147.800 ;
        RECT 250.200 147.400 252.100 147.700 ;
        RECT 250.200 145.700 250.600 147.400 ;
        RECT 253.700 147.100 254.100 147.200 ;
        RECT 256.600 147.100 256.900 148.200 ;
        RECT 259.000 147.500 259.400 149.900 ;
        RECT 260.600 147.600 261.000 149.900 ;
        RECT 262.200 147.600 262.600 149.900 ;
        RECT 260.600 147.200 262.600 147.600 ;
        RECT 258.200 147.100 259.000 147.200 ;
        RECT 253.500 146.800 259.000 147.100 ;
        RECT 252.600 146.400 253.000 146.500 ;
        RECT 251.100 146.100 253.000 146.400 ;
        RECT 251.100 146.000 251.500 146.100 ;
        RECT 251.900 145.700 252.300 145.800 ;
        RECT 250.200 145.400 252.300 145.700 ;
        RECT 249.400 143.800 249.800 145.200 ;
        RECT 250.200 141.100 250.600 145.400 ;
        RECT 253.500 145.200 253.800 146.800 ;
        RECT 257.100 146.700 257.500 146.800 ;
        RECT 257.900 146.200 258.300 146.300 ;
        RECT 255.800 145.900 258.300 146.200 ;
        RECT 255.800 145.800 256.200 145.900 ;
        RECT 260.600 145.800 261.000 147.200 ;
        RECT 256.600 145.500 259.400 145.600 ;
        RECT 256.500 145.400 259.400 145.500 ;
        RECT 252.600 144.900 253.800 145.200 ;
        RECT 254.500 145.300 259.400 145.400 ;
        RECT 254.500 145.100 256.900 145.300 ;
        RECT 252.600 144.400 252.900 144.900 ;
        RECT 252.200 144.200 252.900 144.400 ;
        RECT 253.700 144.500 254.100 144.600 ;
        RECT 254.500 144.500 254.800 145.100 ;
        RECT 253.700 144.200 254.800 144.500 ;
        RECT 255.100 144.500 257.800 144.800 ;
        RECT 255.100 144.400 255.500 144.500 ;
        RECT 257.400 144.400 257.800 144.500 ;
        RECT 251.800 144.000 252.900 144.200 ;
        RECT 251.800 143.800 252.500 144.000 ;
        RECT 254.300 143.700 254.700 143.800 ;
        RECT 255.700 143.700 256.100 143.800 ;
        RECT 252.600 143.100 253.000 143.500 ;
        RECT 254.300 143.400 256.100 143.700 ;
        RECT 254.700 143.100 255.000 143.400 ;
        RECT 257.400 143.100 257.800 143.500 ;
        RECT 252.300 141.100 252.900 143.100 ;
        RECT 254.600 141.100 255.000 143.100 ;
        RECT 256.800 142.800 257.800 143.100 ;
        RECT 256.800 141.100 257.200 142.800 ;
        RECT 259.000 141.100 259.400 145.300 ;
        RECT 260.600 145.400 262.600 145.800 ;
        RECT 260.600 141.100 261.000 145.400 ;
        RECT 262.200 141.100 262.600 145.400 ;
        RECT 0.600 135.700 1.000 139.900 ;
        RECT 2.800 138.200 3.200 139.900 ;
        RECT 2.200 137.900 3.200 138.200 ;
        RECT 5.000 137.900 5.400 139.900 ;
        RECT 7.100 137.900 7.700 139.900 ;
        RECT 2.200 137.500 2.600 137.900 ;
        RECT 5.000 137.600 5.300 137.900 ;
        RECT 3.900 137.300 5.700 137.600 ;
        RECT 7.000 137.500 7.400 137.900 ;
        RECT 3.900 137.200 4.300 137.300 ;
        RECT 5.300 137.200 5.700 137.300 ;
        RECT 2.200 136.500 2.600 136.600 ;
        RECT 4.500 136.500 4.900 136.600 ;
        RECT 2.200 136.200 4.900 136.500 ;
        RECT 5.200 136.500 6.300 136.800 ;
        RECT 5.200 135.900 5.500 136.500 ;
        RECT 5.900 136.400 6.300 136.500 ;
        RECT 7.100 136.600 7.800 137.000 ;
        RECT 7.100 136.100 7.400 136.600 ;
        RECT 3.100 135.700 5.500 135.900 ;
        RECT 0.600 135.600 5.500 135.700 ;
        RECT 6.200 135.800 7.400 136.100 ;
        RECT 0.600 135.500 3.500 135.600 ;
        RECT 0.600 135.400 3.400 135.500 ;
        RECT 3.800 135.100 4.200 135.200 ;
        RECT 1.700 134.800 4.200 135.100 ;
        RECT 1.700 134.700 2.100 134.800 ;
        RECT 2.500 134.200 2.900 134.300 ;
        RECT 6.200 134.200 6.500 135.800 ;
        RECT 9.400 135.600 9.800 139.900 ;
        RECT 11.500 136.300 11.900 139.900 ;
        RECT 11.000 135.900 11.900 136.300 ;
        RECT 12.600 135.900 13.000 139.900 ;
        RECT 13.400 136.200 13.800 139.900 ;
        RECT 15.000 136.200 15.400 139.900 ;
        RECT 17.700 136.400 18.100 139.900 ;
        RECT 19.800 137.500 20.200 139.500 ;
        RECT 13.400 135.900 15.400 136.200 ;
        RECT 17.300 136.100 18.100 136.400 ;
        RECT 7.700 135.300 9.800 135.600 ;
        RECT 7.700 135.200 8.100 135.300 ;
        RECT 8.500 134.900 8.900 135.000 ;
        RECT 7.000 134.600 8.900 134.900 ;
        RECT 7.000 134.500 7.400 134.600 ;
        RECT 1.000 133.900 6.500 134.200 ;
        RECT 1.000 133.800 1.800 133.900 ;
        RECT 0.600 131.100 1.000 133.500 ;
        RECT 3.100 133.200 3.400 133.900 ;
        RECT 5.900 133.800 6.300 133.900 ;
        RECT 9.400 133.600 9.800 135.300 ;
        RECT 11.100 134.200 11.400 135.900 ;
        RECT 11.800 134.800 12.200 135.600 ;
        RECT 12.700 135.200 13.000 135.900 ;
        RECT 14.600 135.200 15.000 135.400 ;
        RECT 12.600 134.900 13.800 135.200 ;
        RECT 14.600 134.900 15.400 135.200 ;
        RECT 12.600 134.800 13.000 134.900 ;
        RECT 11.000 133.800 11.400 134.200 ;
        RECT 12.600 134.200 12.900 134.800 ;
        RECT 12.600 133.800 13.000 134.200 ;
        RECT 7.900 133.300 9.800 133.600 ;
        RECT 7.900 133.200 8.300 133.300 ;
        RECT 2.200 132.100 2.600 132.500 ;
        RECT 3.000 132.400 3.400 133.200 ;
        RECT 9.400 133.100 9.800 133.300 ;
        RECT 10.200 133.100 10.600 133.200 ;
        RECT 11.100 133.100 11.400 133.800 ;
        RECT 12.600 133.100 13.000 133.200 ;
        RECT 13.500 133.100 13.800 134.900 ;
        RECT 15.000 134.800 15.400 134.900 ;
        RECT 15.800 135.100 16.200 135.200 ;
        RECT 16.600 135.100 17.000 135.600 ;
        RECT 15.800 134.800 17.000 135.100 ;
        RECT 14.200 133.800 14.600 134.600 ;
        RECT 17.300 134.200 17.600 136.100 ;
        RECT 19.900 135.800 20.200 137.500 ;
        RECT 22.500 136.400 22.900 139.900 ;
        RECT 24.600 137.500 25.000 139.500 ;
        RECT 18.300 135.500 20.200 135.800 ;
        RECT 22.100 136.100 22.900 136.400 ;
        RECT 18.300 134.500 18.600 135.500 ;
        RECT 16.600 133.800 17.600 134.200 ;
        RECT 17.900 134.100 18.600 134.500 ;
        RECT 19.000 134.400 19.400 135.200 ;
        RECT 19.800 134.400 20.200 135.200 ;
        RECT 20.600 135.100 21.000 135.200 ;
        RECT 21.400 135.100 21.800 135.600 ;
        RECT 20.600 134.800 21.800 135.100 ;
        RECT 22.100 134.200 22.400 136.100 ;
        RECT 24.700 135.800 25.000 137.500 ;
        RECT 26.200 136.400 26.600 139.900 ;
        RECT 23.100 135.500 25.000 135.800 ;
        RECT 26.100 135.900 26.600 136.400 ;
        RECT 27.800 136.200 28.200 139.900 ;
        RECT 30.500 136.400 30.900 139.900 ;
        RECT 32.600 137.500 33.000 139.500 ;
        RECT 26.900 135.900 28.200 136.200 ;
        RECT 30.100 136.100 30.900 136.400 ;
        RECT 23.100 134.500 23.400 135.500 ;
        RECT 9.400 132.800 10.600 133.100 ;
        RECT 11.000 132.800 13.000 133.100 ;
        RECT 3.900 132.700 4.300 132.800 ;
        RECT 3.900 132.400 5.300 132.700 ;
        RECT 5.000 132.100 5.300 132.400 ;
        RECT 7.000 132.100 7.400 132.500 ;
        RECT 2.200 131.800 3.200 132.100 ;
        RECT 2.800 131.100 3.200 131.800 ;
        RECT 5.000 131.100 5.400 132.100 ;
        RECT 7.000 131.800 7.700 132.100 ;
        RECT 7.100 131.100 7.700 131.800 ;
        RECT 9.400 131.100 9.800 132.800 ;
        RECT 10.200 132.400 10.600 132.800 ;
        RECT 11.100 132.100 11.400 132.800 ;
        RECT 12.700 132.400 13.100 132.800 ;
        RECT 11.000 131.100 11.400 132.100 ;
        RECT 13.400 131.100 13.800 133.100 ;
        RECT 17.300 133.500 17.600 133.800 ;
        RECT 18.100 133.900 18.600 134.100 ;
        RECT 18.100 133.600 20.200 133.900 ;
        RECT 21.400 133.800 22.400 134.200 ;
        RECT 22.700 134.100 23.400 134.500 ;
        RECT 23.800 134.400 24.200 135.200 ;
        RECT 24.600 134.400 25.000 135.200 ;
        RECT 17.300 133.300 17.700 133.500 ;
        RECT 17.300 133.000 18.100 133.300 ;
        RECT 17.700 132.200 18.100 133.000 ;
        RECT 19.900 132.500 20.200 133.600 ;
        RECT 22.100 133.500 22.400 133.800 ;
        RECT 22.900 133.900 23.400 134.100 ;
        RECT 26.100 134.200 26.400 135.900 ;
        RECT 26.900 134.900 27.200 135.900 ;
        RECT 26.700 134.500 27.200 134.900 ;
        RECT 22.900 133.600 25.000 133.900 ;
        RECT 22.100 133.300 22.500 133.500 ;
        RECT 22.100 133.200 22.900 133.300 ;
        RECT 22.100 133.000 23.400 133.200 ;
        RECT 17.700 131.800 18.600 132.200 ;
        RECT 17.700 131.500 18.100 131.800 ;
        RECT 19.800 131.500 20.200 132.500 ;
        RECT 22.500 132.800 23.400 133.000 ;
        RECT 22.500 131.500 22.900 132.800 ;
        RECT 24.700 132.500 25.000 133.600 ;
        RECT 26.100 133.800 26.600 134.200 ;
        RECT 26.100 133.100 26.400 133.800 ;
        RECT 26.900 133.700 27.200 134.500 ;
        RECT 27.700 134.800 28.200 135.200 ;
        RECT 29.400 134.800 29.800 135.600 ;
        RECT 27.700 134.400 28.100 134.800 ;
        RECT 30.100 134.200 30.400 136.100 ;
        RECT 32.700 135.800 33.000 137.500 ;
        RECT 31.100 135.500 33.000 135.800 ;
        RECT 33.400 137.100 33.800 139.900 ;
        RECT 34.200 137.100 34.600 137.200 ;
        RECT 33.400 136.800 34.600 137.100 ;
        RECT 31.100 134.500 31.400 135.500 ;
        RECT 29.400 133.800 30.400 134.200 ;
        RECT 30.700 134.100 31.400 134.500 ;
        RECT 31.800 134.400 32.200 135.200 ;
        RECT 32.600 134.400 33.000 135.200 ;
        RECT 26.900 133.400 28.200 133.700 ;
        RECT 26.100 132.800 26.600 133.100 ;
        RECT 24.600 131.500 25.000 132.500 ;
        RECT 26.200 131.100 26.600 132.800 ;
        RECT 27.800 131.100 28.200 133.400 ;
        RECT 30.100 133.500 30.400 133.800 ;
        RECT 30.900 133.900 31.400 134.100 ;
        RECT 30.900 133.600 33.000 133.900 ;
        RECT 30.100 133.300 30.500 133.500 ;
        RECT 30.100 133.200 30.900 133.300 ;
        RECT 30.100 133.000 31.400 133.200 ;
        RECT 30.500 132.800 31.400 133.000 ;
        RECT 30.500 131.500 30.900 132.800 ;
        RECT 32.700 132.500 33.000 133.600 ;
        RECT 32.600 131.500 33.000 132.500 ;
        RECT 33.400 131.100 33.800 136.800 ;
        RECT 35.000 135.600 35.400 139.900 ;
        RECT 37.100 137.900 37.700 139.900 ;
        RECT 39.400 137.900 39.800 139.900 ;
        RECT 41.600 138.200 42.000 139.900 ;
        RECT 41.600 137.900 42.600 138.200 ;
        RECT 37.400 137.500 37.800 137.900 ;
        RECT 39.500 137.600 39.800 137.900 ;
        RECT 39.100 137.300 40.900 137.600 ;
        RECT 42.200 137.500 42.600 137.900 ;
        RECT 39.100 137.200 39.500 137.300 ;
        RECT 40.500 137.200 40.900 137.300 ;
        RECT 37.000 136.600 37.700 137.000 ;
        RECT 37.400 136.100 37.700 136.600 ;
        RECT 38.500 136.500 39.600 136.800 ;
        RECT 38.500 136.400 38.900 136.500 ;
        RECT 37.400 135.800 38.600 136.100 ;
        RECT 35.000 135.300 37.100 135.600 ;
        RECT 35.000 133.600 35.400 135.300 ;
        RECT 36.700 135.200 37.100 135.300 ;
        RECT 35.900 134.900 36.300 135.000 ;
        RECT 35.900 134.600 37.800 134.900 ;
        RECT 37.400 134.500 37.800 134.600 ;
        RECT 38.300 134.200 38.600 135.800 ;
        RECT 39.300 135.900 39.600 136.500 ;
        RECT 39.900 136.500 40.300 136.600 ;
        RECT 42.200 136.500 42.600 136.600 ;
        RECT 39.900 136.200 42.600 136.500 ;
        RECT 39.300 135.700 41.700 135.900 ;
        RECT 43.800 135.700 44.200 139.900 ;
        RECT 39.300 135.600 44.200 135.700 ;
        RECT 41.300 135.500 44.200 135.600 ;
        RECT 41.400 135.400 44.200 135.500 ;
        RECT 44.600 135.700 45.000 139.900 ;
        RECT 46.800 138.200 47.200 139.900 ;
        RECT 46.200 137.900 47.200 138.200 ;
        RECT 49.000 137.900 49.400 139.900 ;
        RECT 51.100 137.900 51.700 139.900 ;
        RECT 46.200 137.500 46.600 137.900 ;
        RECT 49.000 137.600 49.300 137.900 ;
        RECT 47.900 137.300 49.700 137.600 ;
        RECT 51.000 137.500 51.400 137.900 ;
        RECT 47.900 137.200 48.300 137.300 ;
        RECT 49.300 137.200 49.700 137.300 ;
        RECT 46.200 136.500 46.600 136.600 ;
        RECT 48.500 136.500 48.900 136.600 ;
        RECT 46.200 136.200 48.900 136.500 ;
        RECT 49.200 136.500 50.300 136.800 ;
        RECT 49.200 135.900 49.500 136.500 ;
        RECT 49.900 136.400 50.300 136.500 ;
        RECT 51.100 136.600 51.800 137.000 ;
        RECT 51.100 136.100 51.400 136.600 ;
        RECT 47.100 135.700 49.500 135.900 ;
        RECT 44.600 135.600 49.500 135.700 ;
        RECT 50.200 135.800 51.400 136.100 ;
        RECT 44.600 135.500 47.500 135.600 ;
        RECT 44.600 135.400 47.400 135.500 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 47.800 135.100 48.200 135.200 ;
        RECT 40.600 134.800 43.100 135.100 ;
        RECT 42.700 134.700 43.100 134.800 ;
        RECT 45.700 134.800 48.200 135.100 ;
        RECT 45.700 134.700 46.100 134.800 ;
        RECT 41.900 134.200 42.300 134.300 ;
        RECT 46.500 134.200 46.900 134.300 ;
        RECT 50.200 134.200 50.500 135.800 ;
        RECT 53.400 135.600 53.800 139.900 ;
        RECT 57.100 136.200 57.500 139.900 ;
        RECT 57.800 136.800 58.200 137.200 ;
        RECT 57.900 136.200 58.200 136.800 ;
        RECT 56.600 135.800 57.600 136.200 ;
        RECT 57.900 135.900 58.600 136.200 ;
        RECT 58.200 135.800 58.600 135.900 ;
        RECT 51.700 135.300 53.800 135.600 ;
        RECT 51.700 135.200 52.100 135.300 ;
        RECT 52.500 134.900 52.900 135.000 ;
        RECT 51.000 134.600 52.900 134.900 ;
        RECT 51.000 134.500 51.400 134.600 ;
        RECT 38.300 133.900 43.800 134.200 ;
        RECT 38.500 133.800 38.900 133.900 ;
        RECT 35.000 133.300 36.900 133.600 ;
        RECT 34.200 133.100 34.600 133.200 ;
        RECT 35.000 133.100 35.400 133.300 ;
        RECT 36.500 133.200 36.900 133.300 ;
        RECT 41.400 133.200 41.700 133.900 ;
        RECT 43.000 133.800 43.800 133.900 ;
        RECT 45.000 133.900 50.500 134.200 ;
        RECT 45.000 133.800 45.800 133.900 ;
        RECT 34.200 132.800 35.400 133.100 ;
        RECT 34.200 132.400 34.600 132.800 ;
        RECT 35.000 131.100 35.400 132.800 ;
        RECT 40.500 132.700 40.900 132.800 ;
        RECT 37.400 132.100 37.800 132.500 ;
        RECT 39.500 132.400 40.900 132.700 ;
        RECT 41.400 132.400 41.800 133.200 ;
        RECT 39.500 132.100 39.800 132.400 ;
        RECT 42.200 132.100 42.600 132.500 ;
        RECT 37.100 131.800 37.800 132.100 ;
        RECT 37.100 131.100 37.700 131.800 ;
        RECT 39.400 131.100 39.800 132.100 ;
        RECT 41.600 131.800 42.600 132.100 ;
        RECT 41.600 131.100 42.000 131.800 ;
        RECT 43.800 131.100 44.200 133.500 ;
        RECT 44.600 131.100 45.000 133.500 ;
        RECT 47.100 132.800 47.400 133.900 ;
        RECT 49.900 133.800 50.300 133.900 ;
        RECT 53.400 133.600 53.800 135.300 ;
        RECT 56.600 134.400 57.000 135.200 ;
        RECT 57.300 134.200 57.600 135.800 ;
        RECT 59.800 135.600 60.200 139.900 ;
        RECT 61.400 135.600 61.800 139.900 ;
        RECT 63.000 135.600 63.400 139.900 ;
        RECT 64.600 135.600 65.000 139.900 ;
        RECT 67.000 136.400 67.400 139.900 ;
        RECT 59.000 135.200 60.200 135.600 ;
        RECT 60.700 135.200 61.800 135.600 ;
        RECT 62.300 135.200 63.400 135.600 ;
        RECT 64.100 135.200 65.000 135.600 ;
        RECT 66.900 135.900 67.400 136.400 ;
        RECT 68.600 136.200 69.000 139.900 ;
        RECT 70.200 136.400 70.600 139.900 ;
        RECT 67.700 135.900 69.000 136.200 ;
        RECT 70.100 135.900 70.600 136.400 ;
        RECT 71.800 136.200 72.200 139.900 ;
        RECT 70.900 135.900 72.200 136.200 ;
        RECT 72.600 137.500 73.000 139.500 ;
        RECT 74.700 139.200 75.100 139.900 ;
        RECT 74.700 138.800 75.400 139.200 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 55.800 133.800 56.600 134.100 ;
        RECT 57.300 133.800 58.600 134.200 ;
        RECT 59.000 133.800 59.400 135.200 ;
        RECT 60.700 134.500 61.100 135.200 ;
        RECT 62.300 134.500 62.700 135.200 ;
        RECT 64.100 134.500 64.500 135.200 ;
        RECT 59.800 134.100 61.100 134.500 ;
        RECT 61.500 134.100 62.700 134.500 ;
        RECT 63.200 134.100 64.500 134.500 ;
        RECT 64.900 134.100 65.800 134.500 ;
        RECT 60.700 133.800 61.100 134.100 ;
        RECT 62.300 133.800 62.700 134.100 ;
        RECT 64.100 133.800 64.500 134.100 ;
        RECT 65.400 133.800 65.800 134.100 ;
        RECT 66.900 134.200 67.200 135.900 ;
        RECT 67.700 134.900 68.000 135.900 ;
        RECT 67.500 134.500 68.000 134.900 ;
        RECT 66.900 133.800 67.400 134.200 ;
        RECT 56.200 133.600 56.600 133.800 ;
        RECT 51.900 133.300 53.800 133.600 ;
        RECT 51.900 133.200 52.300 133.300 ;
        RECT 46.200 132.100 46.600 132.500 ;
        RECT 47.000 132.400 47.400 132.800 ;
        RECT 47.900 132.700 48.300 132.800 ;
        RECT 47.900 132.400 49.300 132.700 ;
        RECT 49.000 132.100 49.300 132.400 ;
        RECT 51.000 132.100 51.400 132.500 ;
        RECT 46.200 131.800 47.200 132.100 ;
        RECT 46.800 131.100 47.200 131.800 ;
        RECT 49.000 131.100 49.400 132.100 ;
        RECT 51.000 131.800 51.700 132.100 ;
        RECT 51.100 131.100 51.700 131.800 ;
        RECT 53.400 131.100 53.800 133.300 ;
        RECT 55.900 133.100 57.700 133.300 ;
        RECT 58.200 133.100 58.500 133.800 ;
        RECT 59.000 133.400 60.200 133.800 ;
        RECT 60.700 133.400 61.800 133.800 ;
        RECT 62.300 133.400 63.400 133.800 ;
        RECT 64.100 133.400 65.000 133.800 ;
        RECT 55.800 133.000 57.800 133.100 ;
        RECT 55.800 131.100 56.200 133.000 ;
        RECT 57.400 131.100 57.800 133.000 ;
        RECT 58.200 131.100 58.600 133.100 ;
        RECT 59.800 131.100 60.200 133.400 ;
        RECT 61.400 131.100 61.800 133.400 ;
        RECT 63.000 131.100 63.400 133.400 ;
        RECT 64.600 131.100 65.000 133.400 ;
        RECT 66.900 133.100 67.200 133.800 ;
        RECT 67.700 133.700 68.000 134.500 ;
        RECT 68.500 134.800 69.000 135.200 ;
        RECT 68.500 134.400 68.900 134.800 ;
        RECT 70.100 134.200 70.400 135.900 ;
        RECT 70.900 134.900 71.200 135.900 ;
        RECT 72.600 135.800 72.900 137.500 ;
        RECT 74.700 136.400 75.100 138.800 ;
        RECT 74.700 136.100 75.500 136.400 ;
        RECT 72.600 135.500 74.500 135.800 ;
        RECT 70.700 134.500 71.200 134.900 ;
        RECT 70.100 133.800 70.600 134.200 ;
        RECT 67.700 133.400 69.000 133.700 ;
        RECT 66.900 132.800 67.400 133.100 ;
        RECT 67.000 131.100 67.400 132.800 ;
        RECT 68.600 131.100 69.000 133.400 ;
        RECT 70.100 133.100 70.400 133.800 ;
        RECT 70.900 133.700 71.200 134.500 ;
        RECT 71.700 134.800 72.200 135.200 ;
        RECT 71.700 134.400 72.100 134.800 ;
        RECT 72.600 134.400 73.000 135.200 ;
        RECT 73.400 134.400 73.800 135.200 ;
        RECT 74.200 134.500 74.500 135.500 ;
        RECT 74.200 134.100 74.900 134.500 ;
        RECT 75.200 134.200 75.500 136.100 ;
        RECT 77.400 135.700 77.800 139.900 ;
        RECT 79.600 138.200 80.000 139.900 ;
        RECT 79.000 137.900 80.000 138.200 ;
        RECT 81.800 137.900 82.200 139.900 ;
        RECT 83.900 137.900 84.500 139.900 ;
        RECT 79.000 137.500 79.400 137.900 ;
        RECT 81.800 137.600 82.100 137.900 ;
        RECT 80.700 137.300 82.500 137.600 ;
        RECT 83.800 137.500 84.200 137.900 ;
        RECT 80.700 137.200 81.100 137.300 ;
        RECT 82.100 137.200 82.500 137.300 ;
        RECT 79.000 136.500 79.400 136.600 ;
        RECT 81.300 136.500 81.700 136.600 ;
        RECT 79.000 136.200 81.700 136.500 ;
        RECT 82.000 136.500 83.100 136.800 ;
        RECT 82.000 135.900 82.300 136.500 ;
        RECT 82.700 136.400 83.100 136.500 ;
        RECT 83.900 136.600 84.600 137.000 ;
        RECT 83.900 136.100 84.200 136.600 ;
        RECT 79.900 135.700 82.300 135.900 ;
        RECT 77.400 135.600 82.300 135.700 ;
        RECT 83.000 135.800 84.200 136.100 ;
        RECT 75.800 135.100 76.200 135.600 ;
        RECT 77.400 135.500 80.300 135.600 ;
        RECT 77.400 135.400 80.200 135.500 ;
        RECT 76.600 135.100 77.000 135.200 ;
        RECT 80.600 135.100 81.000 135.200 ;
        RECT 81.400 135.100 81.800 135.200 ;
        RECT 75.800 134.800 77.000 135.100 ;
        RECT 78.500 134.800 81.800 135.100 ;
        RECT 78.500 134.700 78.900 134.800 ;
        RECT 79.300 134.200 79.700 134.300 ;
        RECT 83.000 134.200 83.300 135.800 ;
        RECT 86.200 135.600 86.600 139.900 ;
        RECT 87.400 136.800 87.800 137.200 ;
        RECT 87.400 136.200 87.700 136.800 ;
        RECT 88.100 136.200 88.500 139.900 ;
        RECT 87.000 135.900 87.700 136.200 ;
        RECT 88.000 135.900 88.500 136.200 ;
        RECT 87.000 135.800 87.400 135.900 ;
        RECT 84.500 135.300 86.600 135.600 ;
        RECT 84.500 135.200 84.900 135.300 ;
        RECT 85.300 134.900 85.700 135.000 ;
        RECT 83.800 134.600 85.700 134.900 ;
        RECT 83.800 134.500 84.200 134.600 ;
        RECT 74.200 133.900 74.700 134.100 ;
        RECT 70.900 133.400 72.200 133.700 ;
        RECT 70.100 132.800 70.600 133.100 ;
        RECT 70.200 131.100 70.600 132.800 ;
        RECT 71.800 131.100 72.200 133.400 ;
        RECT 72.600 133.600 74.700 133.900 ;
        RECT 75.200 133.800 76.200 134.200 ;
        RECT 77.800 133.900 83.300 134.200 ;
        RECT 77.800 133.800 78.600 133.900 ;
        RECT 72.600 132.500 72.900 133.600 ;
        RECT 75.200 133.500 75.500 133.800 ;
        RECT 75.100 133.300 75.500 133.500 ;
        RECT 74.700 133.000 75.500 133.300 ;
        RECT 72.600 131.500 73.000 132.500 ;
        RECT 74.700 131.500 75.100 133.000 ;
        RECT 77.400 131.100 77.800 133.500 ;
        RECT 79.900 132.800 80.200 133.900 ;
        RECT 82.700 133.800 83.100 133.900 ;
        RECT 86.200 133.600 86.600 135.300 ;
        RECT 87.000 135.100 87.400 135.200 ;
        RECT 88.000 135.100 88.300 135.900 ;
        RECT 90.200 135.600 90.600 139.900 ;
        RECT 92.300 137.900 92.900 139.900 ;
        RECT 94.600 137.900 95.000 139.900 ;
        RECT 96.800 138.200 97.200 139.900 ;
        RECT 96.800 137.900 97.800 138.200 ;
        RECT 92.600 137.500 93.000 137.900 ;
        RECT 94.700 137.600 95.000 137.900 ;
        RECT 94.300 137.300 96.100 137.600 ;
        RECT 97.400 137.500 97.800 137.900 ;
        RECT 94.300 137.200 94.700 137.300 ;
        RECT 95.700 137.200 96.100 137.300 ;
        RECT 92.200 136.600 92.900 137.000 ;
        RECT 92.600 136.100 92.900 136.600 ;
        RECT 93.700 136.500 94.800 136.800 ;
        RECT 93.700 136.400 94.100 136.500 ;
        RECT 92.600 135.800 93.800 136.100 ;
        RECT 90.200 135.300 92.300 135.600 ;
        RECT 87.000 134.800 88.300 135.100 ;
        RECT 88.000 134.200 88.300 134.800 ;
        RECT 88.600 134.400 89.000 135.200 ;
        RECT 87.000 133.800 88.300 134.200 ;
        RECT 89.400 134.100 89.800 134.200 ;
        RECT 89.000 133.800 89.800 134.100 ;
        RECT 84.700 133.300 86.600 133.600 ;
        RECT 84.700 133.200 85.100 133.300 ;
        RECT 79.000 132.100 79.400 132.500 ;
        RECT 79.800 132.400 80.200 132.800 ;
        RECT 80.700 132.700 81.100 132.800 ;
        RECT 80.700 132.400 82.100 132.700 ;
        RECT 81.800 132.100 82.100 132.400 ;
        RECT 83.800 132.100 84.200 132.500 ;
        RECT 79.000 131.800 80.000 132.100 ;
        RECT 79.600 131.100 80.000 131.800 ;
        RECT 81.800 131.100 82.200 132.100 ;
        RECT 83.800 131.800 84.500 132.100 ;
        RECT 83.900 131.100 84.500 131.800 ;
        RECT 86.200 131.100 86.600 133.300 ;
        RECT 87.100 133.100 87.400 133.800 ;
        RECT 89.000 133.600 89.400 133.800 ;
        RECT 90.200 133.600 90.600 135.300 ;
        RECT 91.900 135.200 92.300 135.300 ;
        RECT 91.100 134.900 91.500 135.000 ;
        RECT 91.100 134.600 93.000 134.900 ;
        RECT 92.600 134.500 93.000 134.600 ;
        RECT 93.500 134.200 93.800 135.800 ;
        RECT 94.500 135.900 94.800 136.500 ;
        RECT 95.100 136.500 95.500 136.600 ;
        RECT 97.400 136.500 97.800 136.600 ;
        RECT 95.100 136.200 97.800 136.500 ;
        RECT 94.500 135.700 96.900 135.900 ;
        RECT 99.000 135.700 99.400 139.900 ;
        RECT 99.800 137.900 100.200 139.900 ;
        RECT 99.900 137.800 100.200 137.900 ;
        RECT 101.400 137.900 101.800 139.900 ;
        RECT 101.400 137.800 101.700 137.900 ;
        RECT 99.900 137.500 101.700 137.800 ;
        RECT 99.900 136.200 100.200 137.500 ;
        RECT 100.600 136.400 101.000 137.200 ;
        RECT 99.800 135.800 100.200 136.200 ;
        RECT 94.500 135.600 99.400 135.700 ;
        RECT 96.500 135.500 99.400 135.600 ;
        RECT 96.600 135.400 99.400 135.500 ;
        RECT 95.800 135.100 96.200 135.200 ;
        RECT 95.800 134.800 98.300 135.100 ;
        RECT 97.900 134.700 98.300 134.800 ;
        RECT 97.100 134.200 97.500 134.300 ;
        RECT 99.900 134.200 100.200 135.800 ;
        RECT 102.200 135.400 102.600 136.200 ;
        RECT 101.000 134.800 101.800 135.200 ;
        RECT 93.500 133.900 99.000 134.200 ;
        RECT 99.900 134.100 100.700 134.200 ;
        RECT 99.900 133.900 100.800 134.100 ;
        RECT 93.700 133.800 94.100 133.900 ;
        RECT 90.200 133.300 92.100 133.600 ;
        RECT 87.900 133.100 89.700 133.300 ;
        RECT 87.000 131.100 87.400 133.100 ;
        RECT 87.800 133.000 89.800 133.100 ;
        RECT 87.800 131.100 88.200 133.000 ;
        RECT 89.400 131.100 89.800 133.000 ;
        RECT 90.200 131.100 90.600 133.300 ;
        RECT 91.700 133.200 92.100 133.300 ;
        RECT 96.600 132.800 96.900 133.900 ;
        RECT 98.200 133.800 99.000 133.900 ;
        RECT 95.700 132.700 96.100 132.800 ;
        RECT 92.600 132.100 93.000 132.500 ;
        RECT 94.700 132.400 96.100 132.700 ;
        RECT 96.600 132.400 97.000 132.800 ;
        RECT 94.700 132.100 95.000 132.400 ;
        RECT 97.400 132.100 97.800 132.500 ;
        RECT 92.300 131.800 93.000 132.100 ;
        RECT 92.300 131.100 92.900 131.800 ;
        RECT 94.600 131.100 95.000 132.100 ;
        RECT 96.800 131.800 97.800 132.100 ;
        RECT 96.800 131.100 97.200 131.800 ;
        RECT 99.000 131.100 99.400 133.500 ;
        RECT 100.400 131.100 100.800 133.900 ;
        RECT 103.000 133.400 103.400 134.200 ;
        RECT 103.800 133.100 104.200 139.900 ;
        RECT 107.000 139.600 109.000 139.900 ;
        RECT 104.600 135.800 105.000 136.600 ;
        RECT 107.000 135.900 107.400 139.600 ;
        RECT 107.800 135.900 108.200 139.300 ;
        RECT 108.600 136.200 109.000 139.600 ;
        RECT 110.200 136.200 110.600 139.900 ;
        RECT 108.600 135.900 110.600 136.200 ;
        RECT 107.900 135.600 108.200 135.900 ;
        RECT 111.000 135.700 111.400 139.900 ;
        RECT 113.200 138.200 113.600 139.900 ;
        RECT 112.600 137.900 113.600 138.200 ;
        RECT 115.400 137.900 115.800 139.900 ;
        RECT 117.500 137.900 118.100 139.900 ;
        RECT 112.600 137.500 113.000 137.900 ;
        RECT 115.400 137.600 115.700 137.900 ;
        RECT 114.300 137.300 116.100 137.600 ;
        RECT 117.400 137.500 117.800 137.900 ;
        RECT 114.300 137.200 114.700 137.300 ;
        RECT 115.700 137.200 116.100 137.300 ;
        RECT 112.600 136.500 113.000 136.600 ;
        RECT 114.900 136.500 115.300 136.600 ;
        RECT 112.600 136.200 115.300 136.500 ;
        RECT 115.600 136.500 116.700 136.800 ;
        RECT 115.600 135.900 115.900 136.500 ;
        RECT 116.300 136.400 116.700 136.500 ;
        RECT 117.500 136.600 118.200 137.000 ;
        RECT 117.500 136.100 117.800 136.600 ;
        RECT 113.500 135.700 115.900 135.900 ;
        RECT 111.000 135.600 115.900 135.700 ;
        RECT 116.600 135.800 117.800 136.100 ;
        RECT 107.000 134.800 107.400 135.600 ;
        RECT 107.900 135.300 108.900 135.600 ;
        RECT 111.000 135.500 113.900 135.600 ;
        RECT 111.000 135.400 113.800 135.500 ;
        RECT 108.600 135.200 108.900 135.300 ;
        RECT 109.800 135.200 110.200 135.400 ;
        RECT 108.600 134.800 109.000 135.200 ;
        RECT 109.800 134.900 110.600 135.200 ;
        RECT 114.200 135.100 114.600 135.200 ;
        RECT 110.200 134.800 110.600 134.900 ;
        RECT 112.100 134.800 114.600 135.100 ;
        RECT 107.900 134.400 108.300 134.800 ;
        RECT 107.900 134.200 108.200 134.400 ;
        RECT 107.800 133.800 108.200 134.200 ;
        RECT 108.600 133.100 108.900 134.800 ;
        RECT 112.100 134.700 112.500 134.800 ;
        RECT 109.400 133.800 109.800 134.600 ;
        RECT 112.900 134.200 113.300 134.300 ;
        RECT 116.600 134.200 116.900 135.800 ;
        RECT 119.800 135.600 120.200 139.900 ;
        RECT 121.900 136.200 122.300 139.900 ;
        RECT 122.600 136.800 123.000 137.200 ;
        RECT 122.700 136.200 123.000 136.800 ;
        RECT 121.900 135.900 122.400 136.200 ;
        RECT 122.700 135.900 123.400 136.200 ;
        RECT 118.100 135.300 120.200 135.600 ;
        RECT 118.100 135.200 118.500 135.300 ;
        RECT 118.900 134.900 119.300 135.000 ;
        RECT 117.400 134.600 119.300 134.900 ;
        RECT 117.400 134.500 117.800 134.600 ;
        RECT 111.400 133.900 116.900 134.200 ;
        RECT 111.400 133.800 112.200 133.900 ;
        RECT 103.800 132.800 104.700 133.100 ;
        RECT 104.300 132.200 104.700 132.800 ;
        RECT 108.300 132.200 109.100 133.100 ;
        RECT 103.800 131.800 104.700 132.200 ;
        RECT 107.800 131.800 109.100 132.200 ;
        RECT 104.300 131.100 104.700 131.800 ;
        RECT 108.300 131.100 109.100 131.800 ;
        RECT 111.000 131.100 111.400 133.500 ;
        RECT 113.500 132.800 113.800 133.900 ;
        RECT 115.000 133.800 115.400 133.900 ;
        RECT 116.300 133.800 116.700 133.900 ;
        RECT 119.800 133.600 120.200 135.300 ;
        RECT 122.100 135.200 122.400 135.900 ;
        RECT 123.000 135.800 123.400 135.900 ;
        RECT 123.800 135.800 124.200 136.600 ;
        RECT 121.400 134.400 121.800 135.200 ;
        RECT 122.100 134.800 122.600 135.200 ;
        RECT 123.000 135.100 123.300 135.800 ;
        RECT 124.600 135.100 125.000 139.900 ;
        RECT 127.000 135.600 127.400 139.900 ;
        RECT 128.600 135.600 129.000 139.900 ;
        RECT 130.200 135.600 130.600 139.900 ;
        RECT 131.800 135.600 132.200 139.900 ;
        RECT 134.200 136.400 134.600 139.900 ;
        RECT 134.100 135.900 134.600 136.400 ;
        RECT 135.800 136.200 136.200 139.900 ;
        RECT 134.900 135.900 136.200 136.200 ;
        RECT 127.000 135.200 127.900 135.600 ;
        RECT 128.600 135.200 129.700 135.600 ;
        RECT 130.200 135.200 131.300 135.600 ;
        RECT 131.800 135.200 133.000 135.600 ;
        RECT 123.000 134.800 125.000 135.100 ;
        RECT 122.100 134.200 122.400 134.800 ;
        RECT 120.600 134.100 121.000 134.200 ;
        RECT 120.600 133.800 121.400 134.100 ;
        RECT 122.100 133.800 123.400 134.200 ;
        RECT 121.000 133.600 121.400 133.800 ;
        RECT 118.300 133.300 120.200 133.600 ;
        RECT 118.300 133.200 118.700 133.300 ;
        RECT 112.600 132.100 113.000 132.500 ;
        RECT 113.400 132.400 113.800 132.800 ;
        RECT 114.300 132.700 114.700 132.800 ;
        RECT 114.300 132.400 115.700 132.700 ;
        RECT 115.400 132.100 115.700 132.400 ;
        RECT 117.400 132.100 117.800 132.500 ;
        RECT 112.600 131.800 113.600 132.100 ;
        RECT 113.200 131.100 113.600 131.800 ;
        RECT 115.400 131.100 115.800 132.100 ;
        RECT 117.400 131.800 118.100 132.100 ;
        RECT 117.500 131.100 118.100 131.800 ;
        RECT 119.800 131.100 120.200 133.300 ;
        RECT 120.700 133.100 122.500 133.300 ;
        RECT 123.000 133.100 123.300 133.800 ;
        RECT 124.600 133.100 125.000 134.800 ;
        RECT 127.500 134.500 127.900 135.200 ;
        RECT 129.300 134.500 129.700 135.200 ;
        RECT 130.900 134.500 131.300 135.200 ;
        RECT 125.400 133.400 125.800 134.200 ;
        RECT 126.200 134.100 127.100 134.500 ;
        RECT 127.500 134.100 128.800 134.500 ;
        RECT 129.300 134.100 130.500 134.500 ;
        RECT 130.900 134.100 132.200 134.500 ;
        RECT 126.200 133.800 126.600 134.100 ;
        RECT 127.500 133.800 127.900 134.100 ;
        RECT 129.300 133.800 129.700 134.100 ;
        RECT 130.900 133.800 131.300 134.100 ;
        RECT 132.600 133.800 133.000 135.200 ;
        RECT 127.000 133.400 127.900 133.800 ;
        RECT 128.600 133.400 129.700 133.800 ;
        RECT 130.200 133.400 131.300 133.800 ;
        RECT 131.800 133.400 133.000 133.800 ;
        RECT 134.100 134.200 134.400 135.900 ;
        RECT 134.900 134.900 135.200 135.900 ;
        RECT 134.700 134.500 135.200 134.900 ;
        RECT 134.100 133.800 134.600 134.200 ;
        RECT 120.600 133.000 122.600 133.100 ;
        RECT 120.600 131.100 121.000 133.000 ;
        RECT 122.200 131.100 122.600 133.000 ;
        RECT 123.000 131.100 123.400 133.100 ;
        RECT 124.100 132.800 125.000 133.100 ;
        RECT 124.100 131.100 124.500 132.800 ;
        RECT 127.000 131.100 127.400 133.400 ;
        RECT 128.600 131.100 129.000 133.400 ;
        RECT 130.200 131.100 130.600 133.400 ;
        RECT 131.800 131.100 132.200 133.400 ;
        RECT 134.100 133.100 134.400 133.800 ;
        RECT 134.900 133.700 135.200 134.500 ;
        RECT 135.700 134.800 136.200 135.200 ;
        RECT 135.700 134.400 136.100 134.800 ;
        RECT 134.900 133.400 136.200 133.700 ;
        RECT 136.600 133.400 137.000 134.200 ;
        RECT 134.100 132.800 134.600 133.100 ;
        RECT 134.200 131.100 134.600 132.800 ;
        RECT 135.800 131.100 136.200 133.400 ;
        RECT 137.400 131.100 137.800 139.900 ;
        RECT 138.200 135.800 138.600 136.600 ;
        RECT 139.000 133.100 139.400 139.900 ;
        RECT 139.800 133.400 140.200 134.200 ;
        RECT 140.600 133.400 141.000 134.200 ;
        RECT 138.500 132.800 139.400 133.100 ;
        RECT 141.400 133.100 141.800 139.900 ;
        RECT 142.200 136.100 142.600 136.600 ;
        RECT 143.000 136.100 143.400 136.600 ;
        RECT 142.200 135.800 143.400 136.100 ;
        RECT 143.800 133.100 144.200 139.900 ;
        RECT 144.600 133.400 145.000 134.200 ;
        RECT 145.400 133.400 145.800 134.200 ;
        RECT 141.400 132.800 142.300 133.100 ;
        RECT 138.500 132.200 138.900 132.800 ;
        RECT 141.900 132.200 142.300 132.800 ;
        RECT 143.300 132.800 144.200 133.100 ;
        RECT 146.200 133.100 146.600 139.900 ;
        RECT 147.000 135.800 147.400 136.600 ;
        RECT 148.100 136.300 148.500 139.900 ;
        RECT 150.500 136.300 150.900 139.900 ;
        RECT 148.100 135.900 149.000 136.300 ;
        RECT 150.500 135.900 151.400 136.300 ;
        RECT 147.800 134.800 148.200 135.600 ;
        RECT 148.600 134.200 148.900 135.900 ;
        RECT 150.200 134.800 150.600 135.600 ;
        RECT 151.000 135.100 151.300 135.900 ;
        RECT 152.600 135.800 153.000 136.600 ;
        RECT 152.600 135.100 152.900 135.800 ;
        RECT 151.000 134.800 152.900 135.100 ;
        RECT 151.000 134.200 151.300 134.800 ;
        RECT 147.800 133.800 148.200 134.200 ;
        RECT 148.600 133.800 149.000 134.200 ;
        RECT 150.200 134.100 150.600 134.200 ;
        RECT 151.000 134.100 151.400 134.200 ;
        RECT 150.200 133.800 151.400 134.100 ;
        RECT 147.800 133.100 148.100 133.800 ;
        RECT 148.600 133.100 148.900 133.800 ;
        RECT 146.200 132.800 147.100 133.100 ;
        RECT 147.800 132.800 148.900 133.100 ;
        RECT 143.300 132.200 143.700 132.800 ;
        RECT 138.500 131.800 139.400 132.200 ;
        RECT 141.900 131.800 142.600 132.200 ;
        RECT 143.300 131.800 144.200 132.200 ;
        RECT 138.500 131.100 138.900 131.800 ;
        RECT 141.900 131.100 142.300 131.800 ;
        RECT 143.300 131.100 143.700 131.800 ;
        RECT 146.700 131.100 147.100 132.800 ;
        RECT 148.600 132.100 148.900 132.800 ;
        RECT 149.400 133.100 149.800 133.200 ;
        RECT 150.200 133.100 150.600 133.200 ;
        RECT 149.400 132.800 150.600 133.100 ;
        RECT 149.400 132.400 149.800 132.800 ;
        RECT 151.000 132.100 151.300 133.800 ;
        RECT 151.800 132.400 152.200 133.200 ;
        RECT 153.400 133.100 153.800 139.900 ;
        RECT 155.000 135.800 155.400 136.600 ;
        RECT 154.200 133.400 154.600 134.200 ;
        RECT 155.800 133.100 156.200 139.900 ;
        RECT 158.200 136.100 158.600 136.200 ;
        RECT 159.000 136.100 159.400 136.600 ;
        RECT 158.200 135.800 159.400 136.100 ;
        RECT 156.600 133.400 157.000 134.200 ;
        RECT 159.800 133.100 160.200 139.900 ;
        RECT 162.700 136.300 163.100 139.900 ;
        RECT 162.200 135.900 163.100 136.300 ;
        RECT 160.600 135.100 161.000 135.200 ;
        RECT 162.300 135.100 162.600 135.900 ;
        RECT 163.800 135.800 164.200 136.600 ;
        RECT 160.600 134.800 162.600 135.100 ;
        RECT 163.000 135.100 163.400 135.600 ;
        RECT 163.800 135.100 164.100 135.800 ;
        RECT 163.000 134.800 164.100 135.100 ;
        RECT 162.300 134.200 162.600 134.800 ;
        RECT 160.600 133.400 161.000 134.200 ;
        RECT 162.200 133.800 162.600 134.200 ;
        RECT 152.900 132.800 153.800 133.100 ;
        RECT 155.300 132.800 156.200 133.100 ;
        RECT 159.300 132.800 160.200 133.100 ;
        RECT 148.600 131.100 149.000 132.100 ;
        RECT 151.000 131.100 151.400 132.100 ;
        RECT 152.900 131.100 153.300 132.800 ;
        RECT 155.300 132.200 155.700 132.800 ;
        RECT 155.000 131.800 155.700 132.200 ;
        RECT 155.300 131.100 155.700 131.800 ;
        RECT 159.300 132.200 159.700 132.800 ;
        RECT 161.400 132.400 161.800 133.200 ;
        RECT 159.300 131.800 160.200 132.200 ;
        RECT 162.300 132.100 162.600 133.800 ;
        RECT 164.600 133.100 165.000 139.900 ;
        RECT 167.500 136.300 167.900 139.900 ;
        RECT 167.000 135.900 167.900 136.300 ;
        RECT 167.100 134.200 167.400 135.900 ;
        RECT 168.600 135.600 169.000 139.900 ;
        RECT 170.700 137.900 171.300 139.900 ;
        RECT 173.000 137.900 173.400 139.900 ;
        RECT 175.200 138.200 175.600 139.900 ;
        RECT 175.200 137.900 176.200 138.200 ;
        RECT 171.000 137.500 171.400 137.900 ;
        RECT 173.100 137.600 173.400 137.900 ;
        RECT 172.700 137.300 174.500 137.600 ;
        RECT 175.800 137.500 176.200 137.900 ;
        RECT 172.700 137.200 173.100 137.300 ;
        RECT 174.100 137.200 174.500 137.300 ;
        RECT 170.600 136.600 171.300 137.000 ;
        RECT 171.000 136.100 171.300 136.600 ;
        RECT 172.100 136.500 173.200 136.800 ;
        RECT 172.100 136.400 172.500 136.500 ;
        RECT 171.000 135.800 172.200 136.100 ;
        RECT 167.800 134.800 168.200 135.600 ;
        RECT 168.600 135.300 170.700 135.600 ;
        RECT 165.400 133.400 165.800 134.200 ;
        RECT 167.000 133.800 167.400 134.200 ;
        RECT 159.300 131.100 159.700 131.800 ;
        RECT 162.200 131.100 162.600 132.100 ;
        RECT 164.100 132.800 165.000 133.100 ;
        RECT 164.100 131.100 164.500 132.800 ;
        RECT 166.200 132.400 166.600 133.200 ;
        RECT 167.100 132.200 167.400 133.800 ;
        RECT 167.000 131.100 167.400 132.200 ;
        RECT 168.600 133.600 169.000 135.300 ;
        RECT 170.300 135.200 170.700 135.300 ;
        RECT 169.500 134.900 169.900 135.000 ;
        RECT 169.500 134.600 171.400 134.900 ;
        RECT 171.000 134.500 171.400 134.600 ;
        RECT 171.900 134.200 172.200 135.800 ;
        RECT 172.900 135.900 173.200 136.500 ;
        RECT 173.500 136.500 173.900 136.600 ;
        RECT 175.800 136.500 176.200 136.600 ;
        RECT 173.500 136.200 176.200 136.500 ;
        RECT 172.900 135.700 175.300 135.900 ;
        RECT 177.400 135.700 177.800 139.900 ;
        RECT 172.900 135.600 177.800 135.700 ;
        RECT 174.900 135.500 177.800 135.600 ;
        RECT 178.200 137.500 178.600 139.500 ;
        RECT 178.200 135.800 178.500 137.500 ;
        RECT 180.300 136.400 180.700 139.900 ;
        RECT 180.300 136.100 181.100 136.400 ;
        RECT 178.200 135.500 180.100 135.800 ;
        RECT 175.000 135.400 177.800 135.500 ;
        RECT 174.200 135.100 174.600 135.200 ;
        RECT 174.200 134.800 176.700 135.100 ;
        RECT 175.000 134.700 175.400 134.800 ;
        RECT 176.300 134.700 176.700 134.800 ;
        RECT 178.200 134.400 178.600 135.200 ;
        RECT 179.000 134.400 179.400 135.200 ;
        RECT 179.800 134.500 180.100 135.500 ;
        RECT 175.500 134.200 175.900 134.300 ;
        RECT 171.900 133.900 177.400 134.200 ;
        RECT 179.800 134.100 180.500 134.500 ;
        RECT 180.800 134.200 181.100 136.100 ;
        RECT 181.400 135.100 181.800 135.600 ;
        RECT 183.000 135.100 183.400 139.900 ;
        RECT 184.600 135.700 185.000 139.900 ;
        RECT 186.800 138.200 187.200 139.900 ;
        RECT 186.200 137.900 187.200 138.200 ;
        RECT 189.000 137.900 189.400 139.900 ;
        RECT 191.100 137.900 191.700 139.900 ;
        RECT 186.200 137.500 186.600 137.900 ;
        RECT 189.000 137.600 189.300 137.900 ;
        RECT 187.900 137.300 189.700 137.600 ;
        RECT 191.000 137.500 191.400 137.900 ;
        RECT 187.900 137.200 188.300 137.300 ;
        RECT 189.300 137.200 189.700 137.300 ;
        RECT 186.200 136.500 186.600 136.600 ;
        RECT 188.500 136.500 188.900 136.600 ;
        RECT 186.200 136.200 188.900 136.500 ;
        RECT 189.200 136.500 190.300 136.800 ;
        RECT 189.200 135.900 189.500 136.500 ;
        RECT 189.900 136.400 190.300 136.500 ;
        RECT 191.100 136.600 191.800 137.000 ;
        RECT 191.100 136.100 191.400 136.600 ;
        RECT 187.100 135.700 189.500 135.900 ;
        RECT 184.600 135.600 189.500 135.700 ;
        RECT 190.200 135.800 191.400 136.100 ;
        RECT 184.600 135.500 187.500 135.600 ;
        RECT 184.600 135.400 187.400 135.500 ;
        RECT 190.200 135.200 190.500 135.800 ;
        RECT 193.400 135.600 193.800 139.900 ;
        RECT 191.700 135.300 193.800 135.600 ;
        RECT 191.700 135.200 192.100 135.300 ;
        RECT 187.800 135.100 188.200 135.200 ;
        RECT 181.400 134.800 183.400 135.100 ;
        RECT 179.800 133.900 180.300 134.100 ;
        RECT 172.100 133.800 172.500 133.900 ;
        RECT 174.200 133.800 174.600 133.900 ;
        RECT 168.600 133.300 170.500 133.600 ;
        RECT 168.600 131.100 169.000 133.300 ;
        RECT 170.100 133.200 170.500 133.300 ;
        RECT 175.000 132.800 175.300 133.900 ;
        RECT 176.600 133.800 177.400 133.900 ;
        RECT 178.200 133.600 180.300 133.900 ;
        RECT 180.800 133.800 181.800 134.200 ;
        RECT 174.100 132.700 174.500 132.800 ;
        RECT 171.000 132.100 171.400 132.500 ;
        RECT 173.100 132.400 174.500 132.700 ;
        RECT 175.000 132.400 175.400 132.800 ;
        RECT 173.100 132.100 173.400 132.400 ;
        RECT 175.800 132.100 176.200 132.500 ;
        RECT 170.700 131.800 171.400 132.100 ;
        RECT 170.700 131.100 171.300 131.800 ;
        RECT 173.000 131.100 173.400 132.100 ;
        RECT 175.200 131.800 176.200 132.100 ;
        RECT 175.200 131.100 175.600 131.800 ;
        RECT 177.400 131.100 177.800 133.500 ;
        RECT 178.200 132.500 178.500 133.600 ;
        RECT 180.800 133.500 181.100 133.800 ;
        RECT 180.700 133.300 181.100 133.500 ;
        RECT 180.300 133.000 181.100 133.300 ;
        RECT 178.200 131.500 178.600 132.500 ;
        RECT 180.300 132.200 180.700 133.000 ;
        RECT 180.300 131.800 181.000 132.200 ;
        RECT 180.300 131.500 180.700 131.800 ;
        RECT 183.000 131.100 183.400 134.800 ;
        RECT 185.700 134.800 188.200 135.100 ;
        RECT 190.200 134.800 190.600 135.200 ;
        RECT 192.500 134.900 192.900 135.000 ;
        RECT 185.700 134.700 186.100 134.800 ;
        RECT 187.000 134.700 187.400 134.800 ;
        RECT 186.500 134.200 186.900 134.300 ;
        RECT 190.200 134.200 190.500 134.800 ;
        RECT 191.000 134.600 192.900 134.900 ;
        RECT 191.000 134.500 191.400 134.600 ;
        RECT 185.000 133.900 190.500 134.200 ;
        RECT 185.000 133.800 185.800 133.900 ;
        RECT 183.800 132.400 184.200 133.200 ;
        RECT 184.600 131.100 185.000 133.500 ;
        RECT 187.100 132.800 187.400 133.900 ;
        RECT 189.900 133.800 190.300 133.900 ;
        RECT 193.400 133.600 193.800 135.300 ;
        RECT 191.900 133.300 193.800 133.600 ;
        RECT 194.200 133.400 194.600 134.200 ;
        RECT 191.900 133.200 192.300 133.300 ;
        RECT 186.200 132.100 186.600 132.500 ;
        RECT 187.000 132.400 187.400 132.800 ;
        RECT 187.900 132.700 188.300 132.800 ;
        RECT 187.900 132.400 189.300 132.700 ;
        RECT 189.000 132.100 189.300 132.400 ;
        RECT 191.000 132.100 191.400 132.500 ;
        RECT 186.200 131.800 187.200 132.100 ;
        RECT 186.800 131.100 187.200 131.800 ;
        RECT 189.000 131.100 189.400 132.100 ;
        RECT 191.000 131.800 191.700 132.100 ;
        RECT 191.100 131.100 191.700 131.800 ;
        RECT 193.400 131.100 193.800 133.300 ;
        RECT 195.000 131.100 195.400 139.900 ;
        RECT 197.700 136.400 198.100 139.900 ;
        RECT 200.600 139.600 202.600 139.900 ;
        RECT 199.800 137.500 200.200 139.500 ;
        RECT 197.300 136.100 198.100 136.400 ;
        RECT 196.600 134.800 197.000 135.600 ;
        RECT 197.300 134.200 197.600 136.100 ;
        RECT 199.900 135.800 200.200 137.500 ;
        RECT 200.600 135.900 201.000 139.600 ;
        RECT 201.400 135.900 201.800 139.300 ;
        RECT 202.200 136.200 202.600 139.600 ;
        RECT 203.800 136.200 204.200 139.900 ;
        RECT 202.200 135.900 204.200 136.200 ;
        RECT 198.300 135.500 200.200 135.800 ;
        RECT 201.500 135.600 201.800 135.900 ;
        RECT 198.300 134.500 198.600 135.500 ;
        RECT 196.600 133.800 197.600 134.200 ;
        RECT 197.900 134.100 198.600 134.500 ;
        RECT 199.000 134.400 199.400 135.200 ;
        RECT 199.800 134.400 200.200 135.200 ;
        RECT 200.600 134.800 201.000 135.600 ;
        RECT 201.500 135.300 202.500 135.600 ;
        RECT 202.200 135.200 202.500 135.300 ;
        RECT 203.400 135.200 203.800 135.400 ;
        RECT 202.200 134.800 202.600 135.200 ;
        RECT 203.400 135.100 204.200 135.200 ;
        RECT 204.600 135.100 205.000 135.200 ;
        RECT 203.400 134.900 205.000 135.100 ;
        RECT 203.800 134.800 205.000 134.900 ;
        RECT 201.500 134.400 201.900 134.800 ;
        RECT 201.500 134.200 201.800 134.400 ;
        RECT 197.300 133.500 197.600 133.800 ;
        RECT 198.100 133.900 198.600 134.100 ;
        RECT 198.100 133.600 200.200 133.900 ;
        RECT 201.400 133.800 201.800 134.200 ;
        RECT 197.300 133.300 197.700 133.500 ;
        RECT 197.300 133.200 198.100 133.300 ;
        RECT 197.300 133.000 198.600 133.200 ;
        RECT 197.700 132.800 198.600 133.000 ;
        RECT 197.700 131.500 198.100 132.800 ;
        RECT 199.900 132.500 200.200 133.600 ;
        RECT 202.200 133.200 202.500 134.800 ;
        RECT 203.000 133.800 203.400 134.600 ;
        RECT 204.600 133.400 205.000 134.200 ;
        RECT 202.200 133.100 202.600 133.200 ;
        RECT 205.400 133.100 205.800 139.900 ;
        RECT 206.200 135.800 206.600 136.600 ;
        RECT 199.800 131.500 200.200 132.500 ;
        RECT 201.900 131.100 202.700 133.100 ;
        RECT 205.400 132.800 206.300 133.100 ;
        RECT 205.900 132.200 206.300 132.800 ;
        RECT 205.400 131.800 206.300 132.200 ;
        RECT 205.900 131.100 206.300 131.800 ;
        RECT 207.000 131.100 207.400 139.900 ;
        RECT 210.200 136.200 210.600 139.900 ;
        RECT 211.800 136.400 212.200 139.900 ;
        RECT 215.300 136.400 215.700 139.900 ;
        RECT 217.400 137.500 217.800 139.500 ;
        RECT 210.200 135.900 211.500 136.200 ;
        RECT 211.800 135.900 212.300 136.400 ;
        RECT 210.200 134.800 210.700 135.200 ;
        RECT 210.300 134.400 210.700 134.800 ;
        RECT 211.200 134.900 211.500 135.900 ;
        RECT 211.200 134.500 211.700 134.900 ;
        RECT 207.800 133.400 208.200 134.200 ;
        RECT 211.200 133.700 211.500 134.500 ;
        RECT 212.000 134.200 212.300 135.900 ;
        RECT 214.900 136.100 215.700 136.400 ;
        RECT 214.200 134.800 214.600 135.600 ;
        RECT 214.900 134.200 215.200 136.100 ;
        RECT 217.500 135.800 217.800 137.500 ;
        RECT 218.200 135.900 218.600 139.900 ;
        RECT 219.000 136.200 219.400 139.900 ;
        RECT 220.600 136.200 221.000 139.900 ;
        RECT 219.000 135.900 221.000 136.200 ;
        RECT 221.700 136.300 222.100 139.900 ;
        RECT 221.700 135.900 222.600 136.300 ;
        RECT 215.900 135.500 217.800 135.800 ;
        RECT 215.900 134.500 216.200 135.500 ;
        RECT 218.300 135.200 218.600 135.900 ;
        RECT 220.200 135.200 220.600 135.400 ;
        RECT 211.800 133.800 212.300 134.200 ;
        RECT 212.600 134.100 213.000 134.200 ;
        RECT 214.200 134.100 215.200 134.200 ;
        RECT 215.500 134.100 216.200 134.500 ;
        RECT 216.600 134.400 217.000 135.200 ;
        RECT 217.400 134.400 217.800 135.200 ;
        RECT 218.200 134.900 219.400 135.200 ;
        RECT 220.200 134.900 221.000 135.200 ;
        RECT 218.200 134.800 218.600 134.900 ;
        RECT 212.600 133.800 215.200 134.100 ;
        RECT 210.200 133.400 211.500 133.700 ;
        RECT 210.200 131.100 210.600 133.400 ;
        RECT 212.000 133.100 212.300 133.800 ;
        RECT 211.800 132.800 212.300 133.100 ;
        RECT 214.900 133.500 215.200 133.800 ;
        RECT 215.700 133.900 216.200 134.100 ;
        RECT 215.700 133.600 217.800 133.900 ;
        RECT 214.900 133.300 215.300 133.500 ;
        RECT 214.900 133.000 215.700 133.300 ;
        RECT 211.800 131.100 212.200 132.800 ;
        RECT 215.300 131.500 215.700 133.000 ;
        RECT 217.500 132.500 217.800 133.600 ;
        RECT 218.200 132.800 218.600 133.200 ;
        RECT 219.100 133.100 219.400 134.900 ;
        RECT 220.600 134.800 221.000 134.900 ;
        RECT 221.400 134.800 221.800 135.600 ;
        RECT 219.800 134.100 220.200 134.600 ;
        RECT 221.400 134.100 221.700 134.800 ;
        RECT 219.800 133.800 221.700 134.100 ;
        RECT 222.200 134.200 222.500 135.900 ;
        RECT 223.800 135.600 224.200 139.900 ;
        RECT 225.900 137.900 226.500 139.900 ;
        RECT 228.200 137.900 228.600 139.900 ;
        RECT 230.400 138.200 230.800 139.900 ;
        RECT 230.400 137.900 231.400 138.200 ;
        RECT 226.200 137.500 226.600 137.900 ;
        RECT 228.300 137.600 228.600 137.900 ;
        RECT 227.900 137.300 229.700 137.600 ;
        RECT 231.000 137.500 231.400 137.900 ;
        RECT 227.900 137.200 228.300 137.300 ;
        RECT 229.300 137.200 229.700 137.300 ;
        RECT 225.800 136.600 226.500 137.000 ;
        RECT 226.200 136.100 226.500 136.600 ;
        RECT 227.300 136.500 228.400 136.800 ;
        RECT 227.300 136.400 227.700 136.500 ;
        RECT 226.200 135.800 227.400 136.100 ;
        RECT 223.800 135.300 225.900 135.600 ;
        RECT 222.200 133.800 222.600 134.200 ;
        RECT 217.400 131.500 217.800 132.500 ;
        RECT 218.300 132.400 218.700 132.800 ;
        RECT 219.000 131.100 219.400 133.100 ;
        RECT 221.400 133.100 221.800 133.200 ;
        RECT 222.200 133.100 222.500 133.800 ;
        RECT 223.800 133.600 224.200 135.300 ;
        RECT 225.500 135.200 225.900 135.300 ;
        RECT 224.700 134.900 225.100 135.000 ;
        RECT 224.700 134.600 226.600 134.900 ;
        RECT 226.200 134.500 226.600 134.600 ;
        RECT 227.100 134.200 227.400 135.800 ;
        RECT 228.100 135.900 228.400 136.500 ;
        RECT 228.700 136.500 229.100 136.600 ;
        RECT 231.000 136.500 231.400 136.600 ;
        RECT 228.700 136.200 231.400 136.500 ;
        RECT 228.100 135.700 230.500 135.900 ;
        RECT 232.600 135.700 233.000 139.900 ;
        RECT 228.100 135.600 233.000 135.700 ;
        RECT 234.200 135.600 234.600 139.900 ;
        RECT 235.800 135.600 236.200 139.900 ;
        RECT 237.400 135.600 237.800 139.900 ;
        RECT 239.000 135.600 239.400 139.900 ;
        RECT 240.600 136.200 241.000 139.900 ;
        RECT 242.200 136.200 242.600 139.900 ;
        RECT 240.600 135.900 242.600 136.200 ;
        RECT 243.000 135.900 243.400 139.900 ;
        RECT 230.100 135.500 233.000 135.600 ;
        RECT 230.200 135.400 233.000 135.500 ;
        RECT 233.400 135.200 234.600 135.600 ;
        RECT 235.100 135.200 236.200 135.600 ;
        RECT 236.700 135.200 237.800 135.600 ;
        RECT 238.500 135.200 239.400 135.600 ;
        RECT 243.000 135.200 243.300 135.900 ;
        RECT 243.800 135.600 244.200 139.900 ;
        RECT 245.900 137.900 246.500 139.900 ;
        RECT 248.200 137.900 248.600 139.900 ;
        RECT 250.400 138.200 250.800 139.900 ;
        RECT 250.400 137.900 251.400 138.200 ;
        RECT 246.200 137.500 246.600 137.900 ;
        RECT 248.300 137.600 248.600 137.900 ;
        RECT 247.900 137.300 249.700 137.600 ;
        RECT 251.000 137.500 251.400 137.900 ;
        RECT 247.900 137.200 248.300 137.300 ;
        RECT 249.300 137.200 249.700 137.300 ;
        RECT 245.800 136.600 246.500 137.000 ;
        RECT 246.200 136.100 246.500 136.600 ;
        RECT 247.300 136.500 248.400 136.800 ;
        RECT 247.300 136.400 247.700 136.500 ;
        RECT 246.200 135.800 247.400 136.100 ;
        RECT 243.800 135.300 245.900 135.600 ;
        RECT 229.400 135.100 229.800 135.200 ;
        RECT 229.400 134.800 231.900 135.100 ;
        RECT 230.200 134.700 230.600 134.800 ;
        RECT 231.500 134.700 231.900 134.800 ;
        RECT 230.700 134.200 231.100 134.300 ;
        RECT 227.100 133.900 232.600 134.200 ;
        RECT 227.300 133.800 227.700 133.900 ;
        RECT 223.800 133.300 225.700 133.600 ;
        RECT 221.400 132.800 222.500 133.100 ;
        RECT 222.200 132.100 222.500 132.800 ;
        RECT 223.000 132.400 223.400 133.200 ;
        RECT 222.200 131.100 222.600 132.100 ;
        RECT 223.800 131.100 224.200 133.300 ;
        RECT 225.300 133.200 225.700 133.300 ;
        RECT 230.200 132.800 230.500 133.900 ;
        RECT 231.800 133.800 232.600 133.900 ;
        RECT 233.400 133.800 233.800 135.200 ;
        RECT 235.100 134.500 235.500 135.200 ;
        RECT 236.700 134.500 237.100 135.200 ;
        RECT 238.500 134.500 238.900 135.200 ;
        RECT 242.200 134.900 243.400 135.200 ;
        RECT 242.200 134.800 242.600 134.900 ;
        RECT 243.000 134.800 243.400 134.900 ;
        RECT 234.200 134.100 235.500 134.500 ;
        RECT 235.900 134.100 237.100 134.500 ;
        RECT 237.600 134.100 238.900 134.500 ;
        RECT 239.300 134.100 240.200 134.500 ;
        RECT 235.100 133.800 235.500 134.100 ;
        RECT 236.700 133.800 237.100 134.100 ;
        RECT 238.500 133.800 238.900 134.100 ;
        RECT 239.800 133.800 240.200 134.100 ;
        RECT 241.400 133.800 241.800 134.600 ;
        RECT 229.300 132.700 229.700 132.800 ;
        RECT 226.200 132.100 226.600 132.500 ;
        RECT 228.300 132.400 229.700 132.700 ;
        RECT 230.200 132.400 230.600 132.800 ;
        RECT 228.300 132.100 228.600 132.400 ;
        RECT 231.000 132.100 231.400 132.500 ;
        RECT 225.900 131.800 226.600 132.100 ;
        RECT 225.900 131.100 226.500 131.800 ;
        RECT 228.200 131.100 228.600 132.100 ;
        RECT 230.400 131.800 231.400 132.100 ;
        RECT 230.400 131.100 230.800 131.800 ;
        RECT 232.600 131.100 233.000 133.500 ;
        RECT 233.400 133.400 234.600 133.800 ;
        RECT 235.100 133.400 236.200 133.800 ;
        RECT 236.700 133.400 237.800 133.800 ;
        RECT 238.500 133.400 239.400 133.800 ;
        RECT 234.200 131.100 234.600 133.400 ;
        RECT 235.800 131.100 236.200 133.400 ;
        RECT 237.400 131.100 237.800 133.400 ;
        RECT 239.000 131.100 239.400 133.400 ;
        RECT 242.200 133.100 242.500 134.800 ;
        RECT 243.800 133.600 244.200 135.300 ;
        RECT 245.500 135.200 245.900 135.300 ;
        RECT 244.700 134.900 245.100 135.000 ;
        RECT 244.700 134.600 246.600 134.900 ;
        RECT 246.200 134.500 246.600 134.600 ;
        RECT 247.100 134.200 247.400 135.800 ;
        RECT 248.100 135.900 248.400 136.500 ;
        RECT 248.700 136.500 249.100 136.600 ;
        RECT 251.000 136.500 251.400 136.600 ;
        RECT 248.700 136.200 251.400 136.500 ;
        RECT 248.100 135.700 250.500 135.900 ;
        RECT 252.600 135.700 253.000 139.900 ;
        RECT 253.400 136.200 253.800 139.900 ;
        RECT 255.000 136.200 255.400 139.900 ;
        RECT 253.400 135.900 255.400 136.200 ;
        RECT 255.800 135.900 256.200 139.900 ;
        RECT 257.900 136.300 258.300 139.900 ;
        RECT 260.300 136.300 260.700 139.900 ;
        RECT 257.400 135.900 258.300 136.300 ;
        RECT 259.800 135.900 260.700 136.300 ;
        RECT 261.400 136.200 261.800 139.900 ;
        RECT 261.400 135.900 262.500 136.200 ;
        RECT 248.100 135.600 253.000 135.700 ;
        RECT 250.100 135.500 253.000 135.600 ;
        RECT 250.200 135.400 253.000 135.500 ;
        RECT 255.800 135.200 256.100 135.900 ;
        RECT 257.400 135.800 257.800 135.900 ;
        RECT 249.400 135.100 249.800 135.200 ;
        RECT 249.400 134.800 251.900 135.100 ;
        RECT 250.200 134.700 250.600 134.800 ;
        RECT 251.500 134.700 251.900 134.800 ;
        RECT 255.000 134.900 256.200 135.200 ;
        RECT 255.000 134.800 255.400 134.900 ;
        RECT 255.800 134.800 256.200 134.900 ;
        RECT 250.700 134.200 251.100 134.300 ;
        RECT 247.100 133.900 252.600 134.200 ;
        RECT 247.300 133.800 247.700 133.900 ;
        RECT 243.800 133.300 245.700 133.600 ;
        RECT 242.200 131.100 242.600 133.100 ;
        RECT 243.000 132.800 243.400 133.200 ;
        RECT 242.900 132.400 243.300 132.800 ;
        RECT 243.800 131.100 244.200 133.300 ;
        RECT 245.300 133.200 245.700 133.300 ;
        RECT 250.200 132.800 250.500 133.900 ;
        RECT 251.800 133.800 252.600 133.900 ;
        RECT 254.200 133.800 254.600 134.600 ;
        RECT 249.300 132.700 249.700 132.800 ;
        RECT 246.200 132.100 246.600 132.500 ;
        RECT 248.300 132.400 249.700 132.700 ;
        RECT 250.200 132.400 250.600 132.800 ;
        RECT 248.300 132.100 248.600 132.400 ;
        RECT 251.000 132.100 251.400 132.500 ;
        RECT 245.900 131.800 246.600 132.100 ;
        RECT 245.900 131.100 246.500 131.800 ;
        RECT 248.200 131.100 248.600 132.100 ;
        RECT 250.400 131.800 251.400 132.100 ;
        RECT 250.400 131.100 250.800 131.800 ;
        RECT 252.600 131.100 253.000 133.500 ;
        RECT 255.000 133.100 255.300 134.800 ;
        RECT 257.500 134.200 257.800 135.800 ;
        RECT 259.900 134.200 260.200 135.900 ;
        RECT 262.200 135.600 262.500 135.900 ;
        RECT 262.200 135.200 262.800 135.600 ;
        RECT 261.400 134.400 261.800 135.200 ;
        RECT 257.400 133.800 257.800 134.200 ;
        RECT 259.000 134.100 259.400 134.200 ;
        RECT 259.800 134.100 260.200 134.200 ;
        RECT 259.000 133.800 260.200 134.100 ;
        RECT 255.000 131.100 255.400 133.100 ;
        RECT 255.800 132.800 256.200 133.200 ;
        RECT 255.700 132.400 256.100 132.800 ;
        RECT 257.500 132.100 257.800 133.800 ;
        RECT 259.900 132.100 260.200 133.800 ;
        RECT 262.200 133.700 262.500 135.200 ;
        RECT 257.400 131.100 257.800 132.100 ;
        RECT 259.800 131.100 260.200 132.100 ;
        RECT 261.400 133.400 262.500 133.700 ;
        RECT 261.400 131.100 261.800 133.400 ;
        RECT 1.400 127.600 1.800 129.900 ;
        RECT 3.000 127.600 3.400 129.900 ;
        RECT 4.600 127.600 5.000 129.900 ;
        RECT 6.200 127.600 6.600 129.900 ;
        RECT 0.600 127.200 1.800 127.600 ;
        RECT 2.300 127.200 3.400 127.600 ;
        RECT 3.900 127.200 5.000 127.600 ;
        RECT 5.700 127.200 6.600 127.600 ;
        RECT 7.800 127.500 8.200 129.900 ;
        RECT 10.000 129.200 10.400 129.900 ;
        RECT 9.400 128.900 10.400 129.200 ;
        RECT 12.200 128.900 12.600 129.900 ;
        RECT 14.300 129.200 14.900 129.900 ;
        RECT 14.200 128.900 14.900 129.200 ;
        RECT 9.400 128.500 9.800 128.900 ;
        RECT 12.200 128.600 12.500 128.900 ;
        RECT 10.200 128.200 10.600 128.600 ;
        RECT 11.100 128.300 12.500 128.600 ;
        RECT 14.200 128.500 14.600 128.900 ;
        RECT 11.100 128.200 11.500 128.300 ;
        RECT 0.600 125.800 1.000 127.200 ;
        RECT 2.300 126.900 2.700 127.200 ;
        RECT 3.900 126.900 4.300 127.200 ;
        RECT 5.700 126.900 6.100 127.200 ;
        RECT 7.000 127.100 7.400 127.200 ;
        RECT 8.200 127.100 9.000 127.200 ;
        RECT 10.300 127.100 10.600 128.200 ;
        RECT 15.100 127.700 15.500 127.800 ;
        RECT 16.600 127.700 17.000 129.900 ;
        RECT 18.700 128.200 19.100 129.900 ;
        RECT 15.100 127.400 17.000 127.700 ;
        RECT 18.200 127.900 19.100 128.200 ;
        RECT 19.800 127.900 20.200 129.900 ;
        RECT 20.600 128.000 21.000 129.900 ;
        RECT 22.200 128.000 22.600 129.900 ;
        RECT 24.900 129.200 25.300 129.500 ;
        RECT 24.900 128.800 25.800 129.200 ;
        RECT 24.900 128.000 25.300 128.800 ;
        RECT 27.000 128.500 27.400 129.500 ;
        RECT 20.600 127.900 22.600 128.000 ;
        RECT 13.100 127.100 13.500 127.200 ;
        RECT 16.600 127.100 17.000 127.400 ;
        RECT 17.400 127.100 17.800 127.600 ;
        RECT 7.000 126.900 13.700 127.100 ;
        RECT 1.400 126.500 2.700 126.900 ;
        RECT 3.100 126.500 4.300 126.900 ;
        RECT 4.800 126.500 6.100 126.900 ;
        RECT 6.500 126.800 13.700 126.900 ;
        RECT 6.500 126.500 7.400 126.800 ;
        RECT 9.700 126.700 10.100 126.800 ;
        RECT 2.300 125.800 2.700 126.500 ;
        RECT 3.900 125.800 4.300 126.500 ;
        RECT 5.700 125.800 6.100 126.500 ;
        RECT 8.900 126.200 9.300 126.300 ;
        RECT 8.900 125.900 11.400 126.200 ;
        RECT 11.000 125.800 11.400 125.900 ;
        RECT 0.600 125.400 1.800 125.800 ;
        RECT 2.300 125.400 3.400 125.800 ;
        RECT 3.900 125.400 5.000 125.800 ;
        RECT 5.700 125.400 6.600 125.800 ;
        RECT 1.400 121.100 1.800 125.400 ;
        RECT 3.000 121.100 3.400 125.400 ;
        RECT 4.600 121.100 5.000 125.400 ;
        RECT 6.200 121.100 6.600 125.400 ;
        RECT 7.800 125.500 10.600 125.600 ;
        RECT 7.800 125.400 10.700 125.500 ;
        RECT 7.800 125.300 12.700 125.400 ;
        RECT 7.800 121.100 8.200 125.300 ;
        RECT 10.300 125.100 12.700 125.300 ;
        RECT 9.400 124.500 12.100 124.800 ;
        RECT 9.400 124.400 9.800 124.500 ;
        RECT 11.700 124.400 12.100 124.500 ;
        RECT 12.400 124.500 12.700 125.100 ;
        RECT 13.400 125.200 13.700 126.800 ;
        RECT 16.600 126.800 17.800 127.100 ;
        RECT 14.200 126.400 14.600 126.500 ;
        RECT 14.200 126.100 16.100 126.400 ;
        RECT 15.700 126.000 16.100 126.100 ;
        RECT 14.900 125.700 15.300 125.800 ;
        RECT 16.600 125.700 17.000 126.800 ;
        RECT 14.900 125.400 17.000 125.700 ;
        RECT 13.400 124.900 14.600 125.200 ;
        RECT 13.100 124.500 13.500 124.600 ;
        RECT 12.400 124.200 13.500 124.500 ;
        RECT 14.300 124.400 14.600 124.900 ;
        RECT 14.300 124.000 15.000 124.400 ;
        RECT 11.100 123.700 11.500 123.800 ;
        RECT 12.500 123.700 12.900 123.800 ;
        RECT 9.400 123.100 9.800 123.500 ;
        RECT 11.100 123.400 12.900 123.700 ;
        RECT 12.200 123.100 12.500 123.400 ;
        RECT 14.200 123.100 14.600 123.500 ;
        RECT 9.400 122.800 10.400 123.100 ;
        RECT 10.000 121.100 10.400 122.800 ;
        RECT 12.200 121.100 12.600 123.100 ;
        RECT 14.300 121.100 14.900 123.100 ;
        RECT 16.600 121.100 17.000 125.400 ;
        RECT 18.200 126.100 18.600 127.900 ;
        RECT 19.900 127.200 20.200 127.900 ;
        RECT 20.700 127.700 22.500 127.900 ;
        RECT 24.500 127.700 25.300 128.000 ;
        RECT 24.500 127.500 24.900 127.700 ;
        RECT 21.800 127.200 22.200 127.400 ;
        RECT 24.500 127.200 24.800 127.500 ;
        RECT 27.100 127.400 27.400 128.500 ;
        RECT 27.800 127.500 28.200 129.900 ;
        RECT 30.000 129.200 30.400 129.900 ;
        RECT 29.400 128.900 30.400 129.200 ;
        RECT 32.200 128.900 32.600 129.900 ;
        RECT 34.300 129.200 34.900 129.900 ;
        RECT 34.200 128.900 34.900 129.200 ;
        RECT 29.400 128.500 29.800 128.900 ;
        RECT 32.200 128.600 32.500 128.900 ;
        RECT 30.200 127.800 30.600 128.600 ;
        RECT 31.100 128.300 32.500 128.600 ;
        RECT 34.200 128.500 34.600 128.900 ;
        RECT 31.100 128.200 31.500 128.300 ;
        RECT 19.000 127.100 19.400 127.200 ;
        RECT 19.800 127.100 21.100 127.200 ;
        RECT 19.000 126.800 21.100 127.100 ;
        RECT 21.800 126.900 22.600 127.200 ;
        RECT 22.200 126.800 22.600 126.900 ;
        RECT 23.800 126.800 24.800 127.200 ;
        RECT 25.300 127.100 27.400 127.400 ;
        RECT 28.200 127.100 29.000 127.200 ;
        RECT 30.300 127.100 30.600 127.800 ;
        RECT 35.100 127.700 35.500 127.800 ;
        RECT 36.600 127.700 37.000 129.900 ;
        RECT 37.400 128.000 37.800 129.900 ;
        RECT 39.000 128.000 39.400 129.900 ;
        RECT 37.400 127.900 39.400 128.000 ;
        RECT 39.800 127.900 40.200 129.900 ;
        RECT 40.900 128.200 41.300 129.900 ;
        RECT 40.900 127.900 41.800 128.200 ;
        RECT 44.500 127.900 45.300 129.900 ;
        RECT 48.900 128.000 49.300 129.500 ;
        RECT 51.000 128.500 51.400 129.500 ;
        RECT 37.500 127.700 39.300 127.900 ;
        RECT 35.100 127.400 37.000 127.700 ;
        RECT 33.100 127.100 33.500 127.200 ;
        RECT 25.300 126.900 25.800 127.100 ;
        RECT 18.200 125.800 20.100 126.100 ;
        RECT 18.200 121.100 18.600 125.800 ;
        RECT 19.800 125.200 20.100 125.800 ;
        RECT 19.000 124.400 19.400 125.200 ;
        RECT 19.800 125.100 20.200 125.200 ;
        RECT 20.800 125.100 21.100 126.800 ;
        RECT 21.400 125.800 21.800 126.600 ;
        RECT 23.000 126.100 23.400 126.200 ;
        RECT 23.800 126.100 24.200 126.200 ;
        RECT 23.000 125.800 24.200 126.100 ;
        RECT 23.800 125.400 24.200 125.800 ;
        RECT 19.800 124.800 20.500 125.100 ;
        RECT 20.800 124.800 21.300 125.100 ;
        RECT 20.200 124.200 20.500 124.800 ;
        RECT 20.200 123.800 20.600 124.200 ;
        RECT 20.900 121.100 21.300 124.800 ;
        RECT 24.500 124.900 24.800 126.800 ;
        RECT 25.100 126.500 25.800 126.900 ;
        RECT 28.200 126.800 33.700 127.100 ;
        RECT 29.700 126.700 30.100 126.800 ;
        RECT 25.500 125.500 25.800 126.500 ;
        RECT 26.200 125.800 26.600 126.600 ;
        RECT 27.000 125.800 27.400 126.600 ;
        RECT 28.900 126.200 29.300 126.300 ;
        RECT 28.900 126.100 31.400 126.200 ;
        RECT 31.800 126.100 32.200 126.200 ;
        RECT 28.900 125.900 32.200 126.100 ;
        RECT 31.000 125.800 32.200 125.900 ;
        RECT 27.800 125.500 30.600 125.600 ;
        RECT 25.500 125.200 27.400 125.500 ;
        RECT 24.500 124.600 25.300 124.900 ;
        RECT 24.900 121.100 25.300 124.600 ;
        RECT 27.100 123.500 27.400 125.200 ;
        RECT 27.000 121.500 27.400 123.500 ;
        RECT 27.800 125.400 30.700 125.500 ;
        RECT 27.800 125.300 32.700 125.400 ;
        RECT 27.800 121.100 28.200 125.300 ;
        RECT 30.300 125.100 32.700 125.300 ;
        RECT 29.400 124.500 32.100 124.800 ;
        RECT 29.400 124.400 29.800 124.500 ;
        RECT 31.700 124.400 32.100 124.500 ;
        RECT 32.400 124.500 32.700 125.100 ;
        RECT 33.400 125.200 33.700 126.800 ;
        RECT 34.200 126.400 34.600 126.500 ;
        RECT 34.200 126.100 36.100 126.400 ;
        RECT 35.700 126.000 36.100 126.100 ;
        RECT 34.900 125.700 35.300 125.800 ;
        RECT 36.600 125.700 37.000 127.400 ;
        RECT 37.800 127.200 38.200 127.400 ;
        RECT 39.800 127.200 40.100 127.900 ;
        RECT 37.400 126.900 38.200 127.200 ;
        RECT 37.400 126.800 37.800 126.900 ;
        RECT 38.900 126.800 40.200 127.200 ;
        RECT 38.200 125.800 38.600 126.600 ;
        RECT 38.900 126.200 39.200 126.800 ;
        RECT 38.900 125.800 39.400 126.200 ;
        RECT 41.400 126.100 41.800 127.900 ;
        RECT 42.200 126.800 42.600 127.600 ;
        RECT 43.800 126.400 44.200 127.200 ;
        RECT 44.700 126.200 45.000 127.900 ;
        RECT 48.500 127.700 49.300 128.000 ;
        RECT 48.500 127.500 48.900 127.700 ;
        RECT 48.500 127.200 48.800 127.500 ;
        RECT 51.100 127.400 51.400 128.500 ;
        RECT 53.700 128.200 54.100 129.500 ;
        RECT 55.800 128.500 56.200 129.500 ;
        RECT 58.500 129.200 58.900 129.900 ;
        RECT 58.200 128.800 58.900 129.200 ;
        RECT 53.700 128.000 54.600 128.200 ;
        RECT 45.400 126.800 45.800 127.200 ;
        RECT 47.800 126.800 48.800 127.200 ;
        RECT 49.300 127.100 51.400 127.400 ;
        RECT 53.300 127.800 54.600 128.000 ;
        RECT 53.300 127.700 54.100 127.800 ;
        RECT 53.300 127.500 53.700 127.700 ;
        RECT 53.300 127.200 53.600 127.500 ;
        RECT 55.900 127.400 56.200 128.500 ;
        RECT 58.500 128.200 58.900 128.800 ;
        RECT 60.600 128.500 61.000 129.500 ;
        RECT 58.500 127.900 59.400 128.200 ;
        RECT 49.300 126.900 49.800 127.100 ;
        RECT 45.400 126.600 45.700 126.800 ;
        RECT 45.300 126.200 45.700 126.600 ;
        RECT 39.800 125.800 41.800 126.100 ;
        RECT 42.200 126.100 42.600 126.200 ;
        RECT 43.000 126.100 43.400 126.200 ;
        RECT 42.200 125.800 43.800 126.100 ;
        RECT 44.600 125.800 45.000 126.200 ;
        RECT 34.900 125.400 37.000 125.700 ;
        RECT 33.400 124.900 34.600 125.200 ;
        RECT 33.100 124.500 33.500 124.600 ;
        RECT 32.400 124.200 33.500 124.500 ;
        RECT 34.300 124.400 34.600 124.900 ;
        RECT 34.300 124.000 35.000 124.400 ;
        RECT 31.100 123.700 31.500 123.800 ;
        RECT 32.500 123.700 32.900 123.800 ;
        RECT 29.400 123.100 29.800 123.500 ;
        RECT 31.100 123.400 32.900 123.700 ;
        RECT 32.200 123.100 32.500 123.400 ;
        RECT 34.200 123.100 34.600 123.500 ;
        RECT 29.400 122.800 30.400 123.100 ;
        RECT 30.000 121.100 30.400 122.800 ;
        RECT 32.200 121.100 32.600 123.100 ;
        RECT 34.300 121.100 34.900 123.100 ;
        RECT 36.600 121.100 37.000 125.400 ;
        RECT 38.900 125.100 39.200 125.800 ;
        RECT 39.800 125.200 40.100 125.800 ;
        RECT 39.800 125.100 40.200 125.200 ;
        RECT 38.700 124.800 39.200 125.100 ;
        RECT 39.500 124.800 40.200 125.100 ;
        RECT 38.700 121.100 39.100 124.800 ;
        RECT 39.500 124.200 39.800 124.800 ;
        RECT 40.600 124.400 41.000 125.200 ;
        RECT 39.400 123.800 39.800 124.200 ;
        RECT 41.400 121.100 41.800 125.800 ;
        RECT 43.400 125.600 43.800 125.800 ;
        RECT 44.700 125.700 45.000 125.800 ;
        RECT 46.200 126.100 46.600 126.200 ;
        RECT 47.000 126.100 47.400 126.200 ;
        RECT 46.200 125.800 47.400 126.100 ;
        RECT 44.700 125.400 45.700 125.700 ;
        RECT 46.200 125.400 46.600 125.800 ;
        RECT 47.800 125.400 48.200 126.200 ;
        RECT 45.400 125.100 45.700 125.400 ;
        RECT 48.500 125.200 48.800 126.800 ;
        RECT 49.100 126.500 49.800 126.900 ;
        RECT 52.600 126.800 53.600 127.200 ;
        RECT 54.100 127.100 56.200 127.400 ;
        RECT 54.100 126.900 54.600 127.100 ;
        RECT 49.500 125.500 49.800 126.500 ;
        RECT 50.200 125.800 50.600 126.600 ;
        RECT 51.000 126.100 51.400 126.600 ;
        RECT 51.800 126.100 52.200 126.200 ;
        RECT 51.000 125.800 52.200 126.100 ;
        RECT 49.500 125.200 51.400 125.500 ;
        RECT 52.600 125.400 53.000 126.200 ;
        RECT 43.000 124.800 45.000 125.100 ;
        RECT 43.000 121.100 43.400 124.800 ;
        RECT 44.600 121.400 45.000 124.800 ;
        RECT 45.400 121.700 45.800 125.100 ;
        RECT 46.200 121.400 46.600 125.100 ;
        RECT 48.500 124.900 49.000 125.200 ;
        RECT 48.500 124.600 49.300 124.900 ;
        RECT 44.600 121.100 46.600 121.400 ;
        RECT 48.900 121.100 49.300 124.600 ;
        RECT 51.100 123.500 51.400 125.200 ;
        RECT 53.300 124.900 53.600 126.800 ;
        RECT 53.900 126.500 54.600 126.900 ;
        RECT 54.300 125.500 54.600 126.500 ;
        RECT 55.000 125.800 55.400 126.600 ;
        RECT 55.800 125.800 56.200 126.600 ;
        RECT 54.300 125.200 56.200 125.500 ;
        RECT 53.300 124.600 54.100 124.900 ;
        RECT 51.000 121.500 51.400 123.500 ;
        RECT 53.700 121.100 54.100 124.600 ;
        RECT 55.900 123.500 56.200 125.200 ;
        RECT 56.600 125.100 57.000 125.200 ;
        RECT 58.200 125.100 58.600 125.200 ;
        RECT 56.600 124.800 58.600 125.100 ;
        RECT 58.200 124.400 58.600 124.800 ;
        RECT 55.800 121.500 56.200 123.500 ;
        RECT 59.000 121.100 59.400 127.900 ;
        RECT 59.800 126.800 60.200 127.600 ;
        RECT 60.600 127.400 60.900 128.500 ;
        RECT 62.700 128.200 63.100 129.500 ;
        RECT 62.200 128.000 63.100 128.200 ;
        RECT 62.200 127.800 63.500 128.000 ;
        RECT 66.700 127.900 67.500 129.900 ;
        RECT 62.700 127.700 63.500 127.800 ;
        RECT 63.100 127.500 63.500 127.700 ;
        RECT 60.600 127.100 62.700 127.400 ;
        RECT 62.200 126.900 62.700 127.100 ;
        RECT 63.200 127.200 63.500 127.500 ;
        RECT 67.000 127.200 67.300 127.900 ;
        RECT 69.400 127.500 69.800 129.900 ;
        RECT 71.600 129.200 72.000 129.900 ;
        RECT 71.000 128.900 72.000 129.200 ;
        RECT 73.800 128.900 74.200 129.900 ;
        RECT 75.900 129.200 76.500 129.900 ;
        RECT 75.800 128.900 76.500 129.200 ;
        RECT 71.000 128.500 71.400 128.900 ;
        RECT 73.800 128.600 74.100 128.900 ;
        RECT 71.800 127.800 72.200 128.600 ;
        RECT 72.700 128.300 74.100 128.600 ;
        RECT 75.800 128.500 76.200 128.900 ;
        RECT 72.700 128.200 73.100 128.300 ;
        RECT 60.600 125.800 61.000 126.600 ;
        RECT 61.400 125.800 61.800 126.600 ;
        RECT 62.200 126.500 62.900 126.900 ;
        RECT 63.200 126.800 64.200 127.200 ;
        RECT 66.200 126.800 66.600 127.200 ;
        RECT 62.200 125.500 62.500 126.500 ;
        RECT 60.600 125.200 62.500 125.500 ;
        RECT 60.600 123.500 60.900 125.200 ;
        RECT 63.200 124.900 63.500 126.800 ;
        RECT 66.300 126.600 66.600 126.800 ;
        RECT 67.000 126.800 67.400 127.200 ;
        RECT 66.300 126.200 66.700 126.600 ;
        RECT 67.000 126.200 67.300 126.800 ;
        RECT 67.800 126.400 68.200 127.200 ;
        RECT 69.800 127.100 70.600 127.200 ;
        RECT 71.900 127.100 72.200 127.800 ;
        RECT 76.700 127.700 77.100 127.800 ;
        RECT 78.200 127.700 78.600 129.900 ;
        RECT 79.000 128.000 79.400 129.900 ;
        RECT 80.600 128.000 81.000 129.900 ;
        RECT 79.000 127.900 81.000 128.000 ;
        RECT 81.400 127.900 81.800 129.900 ;
        RECT 83.500 128.200 83.900 129.900 ;
        RECT 85.900 129.200 86.300 129.900 ;
        RECT 85.400 128.800 86.300 129.200 ;
        RECT 85.900 128.200 86.300 128.800 ;
        RECT 83.000 127.900 83.900 128.200 ;
        RECT 85.400 127.900 86.300 128.200 ;
        RECT 87.000 128.500 87.400 129.500 ;
        RECT 79.100 127.700 80.900 127.900 ;
        RECT 76.700 127.400 78.600 127.700 ;
        RECT 74.700 127.100 75.100 127.200 ;
        RECT 69.800 126.800 75.300 127.100 ;
        RECT 71.300 126.700 71.700 126.800 ;
        RECT 70.500 126.200 70.900 126.300 ;
        RECT 63.800 125.400 64.200 126.200 ;
        RECT 65.400 125.400 65.800 126.200 ;
        RECT 67.000 125.800 67.400 126.200 ;
        RECT 68.600 126.100 69.000 126.200 ;
        RECT 68.200 125.800 69.000 126.100 ;
        RECT 70.500 125.900 73.000 126.200 ;
        RECT 72.600 125.800 73.000 125.900 ;
        RECT 67.000 125.700 67.300 125.800 ;
        RECT 66.300 125.400 67.300 125.700 ;
        RECT 68.200 125.600 68.600 125.800 ;
        RECT 69.400 125.500 72.200 125.600 ;
        RECT 69.400 125.400 72.300 125.500 ;
        RECT 66.300 125.100 66.600 125.400 ;
        RECT 69.400 125.300 74.300 125.400 ;
        RECT 62.700 124.600 63.500 124.900 ;
        RECT 60.600 121.500 61.000 123.500 ;
        RECT 62.700 121.100 63.100 124.600 ;
        RECT 65.400 121.400 65.800 125.100 ;
        RECT 66.200 121.700 66.600 125.100 ;
        RECT 67.000 124.800 69.000 125.100 ;
        RECT 67.000 121.400 67.400 124.800 ;
        RECT 65.400 121.100 67.400 121.400 ;
        RECT 68.600 121.100 69.000 124.800 ;
        RECT 69.400 121.100 69.800 125.300 ;
        RECT 71.900 125.100 74.300 125.300 ;
        RECT 71.000 124.500 73.700 124.800 ;
        RECT 71.000 124.400 71.400 124.500 ;
        RECT 73.300 124.400 73.700 124.500 ;
        RECT 74.000 124.500 74.300 125.100 ;
        RECT 75.000 125.200 75.300 126.800 ;
        RECT 75.800 126.400 76.200 126.500 ;
        RECT 75.800 126.100 77.700 126.400 ;
        RECT 77.300 126.000 77.700 126.100 ;
        RECT 76.500 125.700 76.900 125.800 ;
        RECT 78.200 125.700 78.600 127.400 ;
        RECT 79.400 127.200 79.800 127.400 ;
        RECT 81.400 127.200 81.700 127.900 ;
        RECT 79.000 126.900 79.800 127.200 ;
        RECT 79.000 126.800 79.400 126.900 ;
        RECT 80.500 126.800 81.800 127.200 ;
        RECT 82.200 126.800 82.600 127.600 ;
        RECT 79.800 125.800 80.200 126.600 ;
        RECT 76.500 125.400 78.600 125.700 ;
        RECT 75.000 124.900 76.200 125.200 ;
        RECT 74.700 124.500 75.100 124.600 ;
        RECT 74.000 124.200 75.100 124.500 ;
        RECT 75.900 124.400 76.200 124.900 ;
        RECT 75.900 124.000 76.600 124.400 ;
        RECT 72.700 123.700 73.100 123.800 ;
        RECT 74.100 123.700 74.500 123.800 ;
        RECT 71.000 123.100 71.400 123.500 ;
        RECT 72.700 123.400 74.500 123.700 ;
        RECT 73.800 123.100 74.100 123.400 ;
        RECT 75.800 123.100 76.200 123.500 ;
        RECT 71.000 122.800 72.000 123.100 ;
        RECT 71.600 121.100 72.000 122.800 ;
        RECT 73.800 121.100 74.200 123.100 ;
        RECT 75.900 121.100 76.500 123.100 ;
        RECT 78.200 121.100 78.600 125.400 ;
        RECT 80.500 125.100 80.800 126.800 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 83.000 125.100 83.400 127.900 ;
        RECT 84.600 126.800 85.000 127.600 ;
        RECT 80.300 124.800 80.800 125.100 ;
        RECT 81.100 124.800 83.400 125.100 ;
        RECT 80.300 122.200 80.700 124.800 ;
        RECT 81.100 124.200 81.400 124.800 ;
        RECT 81.000 123.800 81.400 124.200 ;
        RECT 79.800 121.800 80.700 122.200 ;
        RECT 80.300 121.100 80.700 121.800 ;
        RECT 83.000 121.100 83.400 124.800 ;
        RECT 83.800 124.400 84.200 125.200 ;
        RECT 85.400 121.100 85.800 127.900 ;
        RECT 87.000 127.400 87.300 128.500 ;
        RECT 89.100 128.000 89.500 129.500 ;
        RECT 89.100 127.700 89.900 128.000 ;
        RECT 89.500 127.500 89.900 127.700 ;
        RECT 87.000 127.100 89.100 127.400 ;
        RECT 88.600 126.900 89.100 127.100 ;
        RECT 89.600 127.200 89.900 127.500 ;
        RECT 91.800 127.700 92.200 129.900 ;
        RECT 93.900 129.200 94.500 129.900 ;
        RECT 93.900 128.900 94.600 129.200 ;
        RECT 96.200 128.900 96.600 129.900 ;
        RECT 98.400 129.200 98.800 129.900 ;
        RECT 98.400 128.900 99.400 129.200 ;
        RECT 94.200 128.500 94.600 128.900 ;
        RECT 96.300 128.600 96.600 128.900 ;
        RECT 96.300 128.300 97.700 128.600 ;
        RECT 97.300 128.200 97.700 128.300 ;
        RECT 98.200 127.800 98.600 128.600 ;
        RECT 99.000 128.500 99.400 128.900 ;
        RECT 93.300 127.700 93.700 127.800 ;
        RECT 91.800 127.400 93.700 127.700 ;
        RECT 87.000 125.800 87.400 126.600 ;
        RECT 87.800 125.800 88.200 126.600 ;
        RECT 88.600 126.500 89.300 126.900 ;
        RECT 89.600 126.800 90.600 127.200 ;
        RECT 88.600 125.500 88.900 126.500 ;
        RECT 87.000 125.200 88.900 125.500 ;
        RECT 86.200 124.400 86.600 125.200 ;
        RECT 87.000 123.500 87.300 125.200 ;
        RECT 89.600 124.900 89.900 126.800 ;
        RECT 90.200 126.100 90.600 126.200 ;
        RECT 91.800 126.100 92.200 127.400 ;
        RECT 95.300 127.100 95.700 127.200 ;
        RECT 98.200 127.100 98.500 127.800 ;
        RECT 100.600 127.500 101.000 129.900 ;
        RECT 101.400 127.600 101.800 129.900 ;
        RECT 103.000 128.200 103.400 129.900 ;
        RECT 105.900 128.200 106.300 129.900 ;
        RECT 103.000 127.900 103.500 128.200 ;
        RECT 101.400 127.300 102.700 127.600 ;
        RECT 99.800 127.100 100.600 127.200 ;
        RECT 95.100 126.800 100.600 127.100 ;
        RECT 94.200 126.400 94.600 126.500 ;
        RECT 90.200 125.800 92.200 126.100 ;
        RECT 92.700 126.100 94.600 126.400 ;
        RECT 92.700 126.000 93.100 126.100 ;
        RECT 90.200 125.400 90.600 125.800 ;
        RECT 91.800 125.700 92.200 125.800 ;
        RECT 93.500 125.700 93.900 125.800 ;
        RECT 91.800 125.400 93.900 125.700 ;
        RECT 89.100 124.600 89.900 124.900 ;
        RECT 87.000 121.500 87.400 123.500 ;
        RECT 89.100 122.200 89.500 124.600 ;
        RECT 88.600 121.800 89.500 122.200 ;
        RECT 89.100 121.100 89.500 121.800 ;
        RECT 91.800 121.100 92.200 125.400 ;
        RECT 95.100 125.200 95.400 126.800 ;
        RECT 98.700 126.700 99.100 126.800 ;
        RECT 99.500 126.200 99.900 126.300 ;
        RECT 101.500 126.200 101.900 126.600 ;
        RECT 97.400 125.900 99.900 126.200 ;
        RECT 97.400 125.800 97.800 125.900 ;
        RECT 101.400 125.800 101.900 126.200 ;
        RECT 102.400 126.500 102.700 127.300 ;
        RECT 103.200 127.200 103.500 127.900 ;
        RECT 105.400 127.900 106.300 128.200 ;
        RECT 103.000 126.800 103.500 127.200 ;
        RECT 104.600 126.800 105.000 127.600 ;
        RECT 102.400 126.100 102.900 126.500 ;
        RECT 98.200 125.500 101.000 125.600 ;
        RECT 98.100 125.400 101.000 125.500 ;
        RECT 94.200 124.900 95.400 125.200 ;
        RECT 96.100 125.300 101.000 125.400 ;
        RECT 96.100 125.100 98.500 125.300 ;
        RECT 94.200 124.400 94.500 124.900 ;
        RECT 93.800 124.000 94.500 124.400 ;
        RECT 95.300 124.500 95.700 124.600 ;
        RECT 96.100 124.500 96.400 125.100 ;
        RECT 95.300 124.200 96.400 124.500 ;
        RECT 96.700 124.500 99.400 124.800 ;
        RECT 96.700 124.400 97.100 124.500 ;
        RECT 99.000 124.400 99.400 124.500 ;
        RECT 95.900 123.700 96.300 123.800 ;
        RECT 97.300 123.700 97.700 123.800 ;
        RECT 94.200 123.100 94.600 123.500 ;
        RECT 95.900 123.400 97.700 123.700 ;
        RECT 96.300 123.100 96.600 123.400 ;
        RECT 99.000 123.100 99.400 123.500 ;
        RECT 93.900 121.100 94.500 123.100 ;
        RECT 96.200 121.100 96.600 123.100 ;
        RECT 98.400 122.800 99.400 123.100 ;
        RECT 98.400 121.100 98.800 122.800 ;
        RECT 100.600 121.100 101.000 125.300 ;
        RECT 102.400 125.100 102.700 126.100 ;
        RECT 103.200 125.100 103.500 126.800 ;
        RECT 101.400 124.800 102.700 125.100 ;
        RECT 101.400 121.100 101.800 124.800 ;
        RECT 103.000 124.600 103.500 125.100 ;
        RECT 104.600 125.100 105.000 125.200 ;
        RECT 105.400 125.100 105.800 127.900 ;
        RECT 110.400 127.100 110.800 129.900 ;
        RECT 113.100 128.200 113.500 129.900 ;
        RECT 112.600 127.900 113.500 128.200 ;
        RECT 115.500 127.900 116.300 129.900 ;
        RECT 110.400 126.900 111.300 127.100 ;
        RECT 110.500 126.800 111.300 126.900 ;
        RECT 111.800 126.800 112.200 127.600 ;
        RECT 109.400 125.800 110.200 126.200 ;
        RECT 104.600 124.800 105.800 125.100 ;
        RECT 103.000 121.100 103.400 124.600 ;
        RECT 105.400 121.100 105.800 124.800 ;
        RECT 106.200 125.100 106.600 125.200 ;
        RECT 107.800 125.100 108.200 125.200 ;
        RECT 106.200 124.800 108.200 125.100 ;
        RECT 108.600 124.800 109.000 125.600 ;
        RECT 111.000 125.200 111.300 126.800 ;
        RECT 111.000 124.800 111.400 125.200 ;
        RECT 106.200 124.400 106.600 124.800 ;
        RECT 109.400 123.800 109.800 124.200 ;
        RECT 110.200 123.800 110.600 124.600 ;
        RECT 109.400 123.500 109.700 123.800 ;
        RECT 111.000 123.500 111.300 124.800 ;
        RECT 109.400 123.200 111.300 123.500 ;
        RECT 109.400 121.100 109.800 123.200 ;
        RECT 111.000 123.100 111.300 123.200 ;
        RECT 111.000 121.100 111.400 123.100 ;
        RECT 112.600 121.100 113.000 127.900 ;
        RECT 115.000 126.800 115.400 127.200 ;
        RECT 115.100 126.600 115.400 126.800 ;
        RECT 115.100 126.200 115.500 126.600 ;
        RECT 115.800 126.200 116.100 127.900 ;
        RECT 116.600 126.400 117.000 127.200 ;
        RECT 118.800 127.100 119.200 129.900 ;
        RECT 122.200 127.600 122.600 129.900 ;
        RECT 123.800 127.600 124.200 129.900 ;
        RECT 125.400 127.600 125.800 129.900 ;
        RECT 127.000 127.600 127.400 129.900 ;
        RECT 130.400 129.200 130.800 129.900 ;
        RECT 130.200 128.800 130.800 129.200 ;
        RECT 122.200 127.200 123.100 127.600 ;
        RECT 123.800 127.200 124.900 127.600 ;
        RECT 125.400 127.200 126.500 127.600 ;
        RECT 127.000 127.200 128.200 127.600 ;
        RECT 118.300 126.900 119.200 127.100 ;
        RECT 118.300 126.800 119.100 126.900 ;
        RECT 119.800 126.800 120.200 127.200 ;
        RECT 121.400 126.900 121.800 127.200 ;
        RECT 122.700 126.900 123.100 127.200 ;
        RECT 124.500 126.900 124.900 127.200 ;
        RECT 126.100 126.900 126.500 127.200 ;
        RECT 114.200 125.400 114.600 126.200 ;
        RECT 115.800 125.800 116.200 126.200 ;
        RECT 117.400 126.100 117.800 126.200 ;
        RECT 117.000 125.800 117.800 126.100 ;
        RECT 115.800 125.700 116.100 125.800 ;
        RECT 115.100 125.400 116.100 125.700 ;
        RECT 117.000 125.600 117.400 125.800 ;
        RECT 115.100 125.200 115.400 125.400 ;
        RECT 118.300 125.200 118.600 126.800 ;
        RECT 119.800 126.200 120.100 126.800 ;
        RECT 121.400 126.500 122.300 126.900 ;
        RECT 122.700 126.500 124.000 126.900 ;
        RECT 124.500 126.500 125.700 126.900 ;
        RECT 126.100 126.500 127.400 126.900 ;
        RECT 119.400 125.800 120.200 126.200 ;
        RECT 122.700 125.800 123.100 126.500 ;
        RECT 124.500 125.800 124.900 126.500 ;
        RECT 126.100 125.800 126.500 126.500 ;
        RECT 127.800 125.800 128.200 127.200 ;
        RECT 130.400 127.100 130.800 128.800 ;
        RECT 131.800 127.500 132.200 129.900 ;
        RECT 134.000 129.200 134.400 129.900 ;
        RECT 133.400 128.900 134.400 129.200 ;
        RECT 136.200 128.900 136.600 129.900 ;
        RECT 138.300 129.200 138.900 129.900 ;
        RECT 138.200 128.900 138.900 129.200 ;
        RECT 133.400 128.500 133.800 128.900 ;
        RECT 136.200 128.600 136.500 128.900 ;
        RECT 134.200 128.200 134.600 128.600 ;
        RECT 135.100 128.300 136.500 128.600 ;
        RECT 138.200 128.500 138.600 128.900 ;
        RECT 135.100 128.200 135.500 128.300 ;
        RECT 132.200 127.100 133.000 127.200 ;
        RECT 134.300 127.100 134.600 128.200 ;
        RECT 139.100 127.700 139.500 127.800 ;
        RECT 140.600 127.700 141.000 129.900 ;
        RECT 141.400 128.000 141.800 129.900 ;
        RECT 143.000 128.000 143.400 129.900 ;
        RECT 141.400 127.900 143.400 128.000 ;
        RECT 143.800 127.900 144.200 129.900 ;
        RECT 144.900 128.200 145.300 129.900 ;
        RECT 147.000 128.500 147.400 129.500 ;
        RECT 144.900 127.900 145.800 128.200 ;
        RECT 141.500 127.700 143.300 127.900 ;
        RECT 139.100 127.400 141.000 127.700 ;
        RECT 137.100 127.100 137.500 127.200 ;
        RECT 130.400 126.900 131.300 127.100 ;
        RECT 130.500 126.800 131.300 126.900 ;
        RECT 132.200 126.800 137.700 127.100 ;
        RECT 129.400 125.800 130.200 126.200 ;
        RECT 113.400 124.400 113.800 125.200 ;
        RECT 114.200 121.400 114.600 125.100 ;
        RECT 115.000 121.700 115.400 125.200 ;
        RECT 115.800 124.800 117.800 125.100 ;
        RECT 118.200 124.800 118.600 125.200 ;
        RECT 119.800 125.100 120.200 125.200 ;
        RECT 120.600 125.100 121.000 125.600 ;
        RECT 119.800 124.800 121.000 125.100 ;
        RECT 122.200 125.400 123.100 125.800 ;
        RECT 123.800 125.400 124.900 125.800 ;
        RECT 125.400 125.400 126.500 125.800 ;
        RECT 127.000 125.400 128.200 125.800 ;
        RECT 115.800 121.400 116.200 124.800 ;
        RECT 114.200 121.100 116.200 121.400 ;
        RECT 117.400 121.100 117.800 124.800 ;
        RECT 118.300 124.200 118.600 124.800 ;
        RECT 118.200 123.800 118.600 124.200 ;
        RECT 119.000 123.800 119.400 124.600 ;
        RECT 118.300 123.500 118.600 123.800 ;
        RECT 118.300 123.200 120.100 123.500 ;
        RECT 118.300 123.100 118.600 123.200 ;
        RECT 118.200 121.100 118.600 123.100 ;
        RECT 119.800 123.100 120.100 123.200 ;
        RECT 119.800 121.100 120.200 123.100 ;
        RECT 122.200 121.100 122.600 125.400 ;
        RECT 123.800 121.100 124.200 125.400 ;
        RECT 125.400 121.100 125.800 125.400 ;
        RECT 127.000 121.100 127.400 125.400 ;
        RECT 128.600 124.800 129.000 125.600 ;
        RECT 131.000 125.200 131.300 126.800 ;
        RECT 133.700 126.700 134.100 126.800 ;
        RECT 132.900 126.200 133.300 126.300 ;
        RECT 132.900 125.900 135.400 126.200 ;
        RECT 135.000 125.800 135.400 125.900 ;
        RECT 131.800 125.500 134.600 125.600 ;
        RECT 131.800 125.400 134.700 125.500 ;
        RECT 131.800 125.300 136.700 125.400 ;
        RECT 131.000 124.800 131.400 125.200 ;
        RECT 130.200 123.800 130.600 124.600 ;
        RECT 131.000 123.500 131.300 124.800 ;
        RECT 129.500 123.200 131.300 123.500 ;
        RECT 129.500 123.100 129.800 123.200 ;
        RECT 129.400 121.100 129.800 123.100 ;
        RECT 131.000 123.100 131.300 123.200 ;
        RECT 131.000 121.100 131.400 123.100 ;
        RECT 131.800 121.100 132.200 125.300 ;
        RECT 134.300 125.100 136.700 125.300 ;
        RECT 133.400 124.500 136.100 124.800 ;
        RECT 133.400 124.400 133.800 124.500 ;
        RECT 135.700 124.400 136.100 124.500 ;
        RECT 136.400 124.500 136.700 125.100 ;
        RECT 137.400 125.200 137.700 126.800 ;
        RECT 138.200 126.400 138.600 126.500 ;
        RECT 138.200 126.100 140.100 126.400 ;
        RECT 139.700 126.000 140.100 126.100 ;
        RECT 138.900 125.700 139.300 125.800 ;
        RECT 140.600 125.700 141.000 127.400 ;
        RECT 141.800 127.200 142.200 127.400 ;
        RECT 143.800 127.200 144.100 127.900 ;
        RECT 141.400 126.900 142.200 127.200 ;
        RECT 141.400 126.800 141.800 126.900 ;
        RECT 142.900 126.800 144.200 127.200 ;
        RECT 142.200 125.800 142.600 126.600 ;
        RECT 142.900 126.200 143.200 126.800 ;
        RECT 142.900 125.800 143.400 126.200 ;
        RECT 145.400 126.100 145.800 127.900 ;
        RECT 146.200 126.800 146.600 127.600 ;
        RECT 147.000 127.400 147.300 128.500 ;
        RECT 149.100 128.000 149.500 129.500 ;
        RECT 153.700 128.000 154.100 129.500 ;
        RECT 155.800 128.500 156.200 129.500 ;
        RECT 149.100 127.700 149.900 128.000 ;
        RECT 149.500 127.500 149.900 127.700 ;
        RECT 147.000 127.100 149.100 127.400 ;
        RECT 148.600 126.900 149.100 127.100 ;
        RECT 149.600 127.200 149.900 127.500 ;
        RECT 153.300 127.700 154.100 128.000 ;
        RECT 153.300 127.500 153.700 127.700 ;
        RECT 153.300 127.200 153.600 127.500 ;
        RECT 155.900 127.400 156.200 128.500 ;
        RECT 143.800 125.800 145.800 126.100 ;
        RECT 147.000 125.800 147.400 126.600 ;
        RECT 147.800 125.800 148.200 126.600 ;
        RECT 148.600 126.500 149.300 126.900 ;
        RECT 149.600 126.800 150.600 127.200 ;
        RECT 152.600 126.800 153.600 127.200 ;
        RECT 154.100 127.100 156.200 127.400 ;
        RECT 154.100 126.900 154.600 127.100 ;
        RECT 138.900 125.400 141.000 125.700 ;
        RECT 137.400 124.900 138.600 125.200 ;
        RECT 137.100 124.500 137.500 124.600 ;
        RECT 136.400 124.200 137.500 124.500 ;
        RECT 138.300 124.400 138.600 124.900 ;
        RECT 138.300 124.000 139.000 124.400 ;
        RECT 135.100 123.700 135.500 123.800 ;
        RECT 136.500 123.700 136.900 123.800 ;
        RECT 133.400 123.100 133.800 123.500 ;
        RECT 135.100 123.400 136.900 123.700 ;
        RECT 136.200 123.100 136.500 123.400 ;
        RECT 138.200 123.100 138.600 123.500 ;
        RECT 133.400 122.800 134.400 123.100 ;
        RECT 134.000 121.100 134.400 122.800 ;
        RECT 136.200 121.100 136.600 123.100 ;
        RECT 138.300 121.100 138.900 123.100 ;
        RECT 140.600 121.100 141.000 125.400 ;
        RECT 142.900 125.100 143.200 125.800 ;
        RECT 143.800 125.200 144.100 125.800 ;
        RECT 143.800 125.100 144.200 125.200 ;
        RECT 142.700 124.800 143.200 125.100 ;
        RECT 143.500 124.800 144.200 125.100 ;
        RECT 142.700 121.100 143.100 124.800 ;
        RECT 143.500 124.200 143.800 124.800 ;
        RECT 144.600 124.400 145.000 125.200 ;
        RECT 143.400 123.800 143.800 124.200 ;
        RECT 145.400 121.100 145.800 125.800 ;
        RECT 148.600 125.500 148.900 126.500 ;
        RECT 147.000 125.200 148.900 125.500 ;
        RECT 147.000 123.500 147.300 125.200 ;
        RECT 149.600 124.900 149.900 126.800 ;
        RECT 150.200 125.400 150.600 126.200 ;
        RECT 152.600 125.400 153.000 126.200 ;
        RECT 149.100 124.600 149.900 124.900 ;
        RECT 153.300 125.200 153.600 126.800 ;
        RECT 153.900 126.500 154.600 126.900 ;
        RECT 158.200 126.800 158.600 127.600 ;
        RECT 159.000 127.100 159.400 129.900 ;
        RECT 161.100 128.200 161.500 129.900 ;
        RECT 162.500 129.200 162.900 129.900 ;
        RECT 162.200 128.800 162.900 129.200 ;
        RECT 162.500 128.400 162.900 128.800 ;
        RECT 160.600 127.900 161.500 128.200 ;
        RECT 162.200 127.900 162.900 128.400 ;
        RECT 164.600 127.900 165.000 129.900 ;
        RECT 166.200 128.900 166.600 129.900 ;
        RECT 159.800 127.100 160.200 127.600 ;
        RECT 159.000 126.800 160.200 127.100 ;
        RECT 154.300 125.500 154.600 126.500 ;
        RECT 155.000 125.800 155.400 126.600 ;
        RECT 155.800 125.800 156.200 126.600 ;
        RECT 154.300 125.200 156.200 125.500 ;
        RECT 153.300 124.900 153.800 125.200 ;
        RECT 153.300 124.600 154.100 124.900 ;
        RECT 147.000 121.500 147.400 123.500 ;
        RECT 149.100 122.200 149.500 124.600 ;
        RECT 149.100 121.800 149.800 122.200 ;
        RECT 149.100 121.100 149.500 121.800 ;
        RECT 153.700 121.100 154.100 124.600 ;
        RECT 155.900 123.500 156.200 125.200 ;
        RECT 155.800 121.500 156.200 123.500 ;
        RECT 159.000 121.100 159.400 126.800 ;
        RECT 160.600 121.100 161.000 127.900 ;
        RECT 162.200 126.200 162.500 127.900 ;
        RECT 164.600 127.800 164.900 127.900 ;
        RECT 165.400 127.800 165.800 128.600 ;
        RECT 164.000 127.600 164.900 127.800 ;
        RECT 162.800 127.500 164.900 127.600 ;
        RECT 162.800 127.300 164.300 127.500 ;
        RECT 162.800 127.200 163.200 127.300 ;
        RECT 166.300 127.200 166.600 128.900 ;
        RECT 167.800 128.000 168.200 129.900 ;
        RECT 169.400 128.000 169.800 129.900 ;
        RECT 167.800 127.900 169.800 128.000 ;
        RECT 170.200 127.900 170.600 129.900 ;
        RECT 171.800 128.200 172.200 129.900 ;
        RECT 171.700 127.900 172.200 128.200 ;
        RECT 167.900 127.700 169.700 127.900 ;
        RECT 168.200 127.200 168.600 127.400 ;
        RECT 170.200 127.200 170.500 127.900 ;
        RECT 171.700 127.200 172.000 127.900 ;
        RECT 173.400 127.600 173.800 129.900 ;
        RECT 172.500 127.300 173.800 127.600 ;
        RECT 174.200 127.600 174.600 129.900 ;
        RECT 175.800 128.200 176.200 129.900 ;
        RECT 175.800 127.900 176.300 128.200 ;
        RECT 174.200 127.300 175.500 127.600 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 161.400 125.100 161.800 125.200 ;
        RECT 162.200 125.100 162.500 125.800 ;
        RECT 162.900 125.500 163.200 127.200 ;
        RECT 163.600 126.900 164.000 127.000 ;
        RECT 163.600 126.600 164.100 126.900 ;
        RECT 163.800 126.200 164.100 126.600 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 164.600 125.800 165.000 127.200 ;
        RECT 166.200 126.800 166.600 127.200 ;
        RECT 167.000 127.100 167.400 127.200 ;
        RECT 167.800 127.100 168.600 127.200 ;
        RECT 167.000 126.900 168.600 127.100 ;
        RECT 169.300 127.100 170.600 127.200 ;
        RECT 171.000 127.100 171.400 127.200 ;
        RECT 167.000 126.800 168.200 126.900 ;
        RECT 169.300 126.800 171.400 127.100 ;
        RECT 171.700 126.800 172.200 127.200 ;
        RECT 165.400 126.100 165.800 126.200 ;
        RECT 166.300 126.100 166.600 126.800 ;
        RECT 165.400 125.800 166.600 126.100 ;
        RECT 162.900 125.200 164.100 125.500 ;
        RECT 161.400 124.800 162.600 125.100 ;
        RECT 161.400 124.400 161.800 124.800 ;
        RECT 162.200 121.100 162.600 124.800 ;
        RECT 163.800 123.100 164.100 125.200 ;
        RECT 166.300 125.100 166.600 125.800 ;
        RECT 167.000 126.100 167.400 126.200 ;
        RECT 167.000 125.800 168.100 126.100 ;
        RECT 168.600 125.800 169.000 126.600 ;
        RECT 167.000 125.400 167.400 125.800 ;
        RECT 169.300 125.100 169.600 126.800 ;
        RECT 170.200 125.100 170.600 125.200 ;
        RECT 166.200 124.700 167.100 125.100 ;
        RECT 163.800 121.100 164.200 123.100 ;
        RECT 166.700 121.100 167.100 124.700 ;
        RECT 169.100 124.800 169.600 125.100 ;
        RECT 169.900 124.800 170.600 125.100 ;
        RECT 171.700 125.100 172.000 126.800 ;
        RECT 172.500 126.500 172.800 127.300 ;
        RECT 172.300 126.100 172.800 126.500 ;
        RECT 172.500 125.100 172.800 126.100 ;
        RECT 173.300 126.200 173.700 126.600 ;
        RECT 174.300 126.200 174.700 126.600 ;
        RECT 173.300 126.100 173.800 126.200 ;
        RECT 174.200 126.100 174.700 126.200 ;
        RECT 173.300 125.800 174.700 126.100 ;
        RECT 175.200 126.500 175.500 127.300 ;
        RECT 176.000 127.200 176.300 127.900 ;
        RECT 175.800 126.800 176.300 127.200 ;
        RECT 175.200 126.100 175.700 126.500 ;
        RECT 175.200 125.100 175.500 126.100 ;
        RECT 176.000 125.100 176.300 126.800 ;
        RECT 169.100 121.100 169.500 124.800 ;
        RECT 169.900 124.200 170.200 124.800 ;
        RECT 171.700 124.600 172.200 125.100 ;
        RECT 172.500 124.800 173.800 125.100 ;
        RECT 169.800 123.800 170.200 124.200 ;
        RECT 171.800 121.100 172.200 124.600 ;
        RECT 173.400 121.100 173.800 124.800 ;
        RECT 174.200 124.800 175.500 125.100 ;
        RECT 174.200 121.100 174.600 124.800 ;
        RECT 175.800 124.600 176.300 125.100 ;
        RECT 175.800 121.100 176.200 124.600 ;
        RECT 178.200 121.100 178.600 129.900 ;
        RECT 181.400 127.900 181.800 129.900 ;
        RECT 182.100 128.200 182.500 128.600 ;
        RECT 184.300 128.200 184.700 129.900 ;
        RECT 180.600 126.400 181.000 127.200 ;
        RECT 179.000 126.100 179.400 126.200 ;
        RECT 179.800 126.100 180.200 126.200 ;
        RECT 181.400 126.100 181.700 127.900 ;
        RECT 182.200 127.800 182.600 128.200 ;
        RECT 183.800 127.900 184.700 128.200 ;
        RECT 182.200 126.100 182.600 126.200 ;
        RECT 179.000 125.800 180.600 126.100 ;
        RECT 181.400 125.800 182.600 126.100 ;
        RECT 180.200 125.600 180.600 125.800 ;
        RECT 182.200 125.100 182.500 125.800 ;
        RECT 179.800 124.800 181.800 125.100 ;
        RECT 179.800 121.100 180.200 124.800 ;
        RECT 181.400 121.100 181.800 124.800 ;
        RECT 182.200 121.100 182.600 125.100 ;
        RECT 183.800 121.100 184.200 127.900 ;
        RECT 185.400 127.500 185.800 129.900 ;
        RECT 187.600 129.200 188.000 129.900 ;
        RECT 187.000 128.900 188.000 129.200 ;
        RECT 189.800 128.900 190.200 129.900 ;
        RECT 191.900 129.200 192.500 129.900 ;
        RECT 191.800 128.900 192.500 129.200 ;
        RECT 187.000 128.500 187.400 128.900 ;
        RECT 189.800 128.600 190.100 128.900 ;
        RECT 187.800 128.200 188.200 128.600 ;
        RECT 188.700 128.300 190.100 128.600 ;
        RECT 191.800 128.500 192.200 128.900 ;
        RECT 188.700 128.200 189.100 128.300 ;
        RECT 185.800 127.100 186.600 127.200 ;
        RECT 187.900 127.100 188.200 128.200 ;
        RECT 192.700 127.700 193.100 127.800 ;
        RECT 194.200 127.700 194.600 129.900 ;
        RECT 192.700 127.400 194.600 127.700 ;
        RECT 195.800 127.600 196.200 129.900 ;
        RECT 197.400 127.600 197.800 129.900 ;
        RECT 199.000 127.600 199.400 129.900 ;
        RECT 200.600 127.600 201.000 129.900 ;
        RECT 190.700 127.100 191.100 127.200 ;
        RECT 185.800 126.800 191.300 127.100 ;
        RECT 187.300 126.700 187.700 126.800 ;
        RECT 186.500 126.200 186.900 126.300 ;
        RECT 187.800 126.200 188.200 126.300 ;
        RECT 191.000 126.200 191.300 126.800 ;
        RECT 191.800 126.400 192.200 126.500 ;
        RECT 186.500 125.900 189.000 126.200 ;
        RECT 188.600 125.800 189.000 125.900 ;
        RECT 191.000 125.800 191.400 126.200 ;
        RECT 191.800 126.100 193.700 126.400 ;
        RECT 193.300 126.000 193.700 126.100 ;
        RECT 185.400 125.500 188.200 125.600 ;
        RECT 185.400 125.400 188.300 125.500 ;
        RECT 185.400 125.300 190.300 125.400 ;
        RECT 184.600 124.400 185.000 125.200 ;
        RECT 185.400 121.100 185.800 125.300 ;
        RECT 187.900 125.100 190.300 125.300 ;
        RECT 187.000 124.500 189.700 124.800 ;
        RECT 187.000 124.400 187.400 124.500 ;
        RECT 189.300 124.400 189.700 124.500 ;
        RECT 190.000 124.500 190.300 125.100 ;
        RECT 191.000 125.200 191.300 125.800 ;
        RECT 192.500 125.700 192.900 125.800 ;
        RECT 194.200 125.700 194.600 127.400 ;
        RECT 192.500 125.400 194.600 125.700 ;
        RECT 195.000 127.200 196.200 127.600 ;
        RECT 196.700 127.200 197.800 127.600 ;
        RECT 198.300 127.200 199.400 127.600 ;
        RECT 200.100 127.200 201.000 127.600 ;
        RECT 202.200 127.600 202.600 129.900 ;
        RECT 204.600 128.000 205.000 129.900 ;
        RECT 206.200 128.000 206.600 129.900 ;
        RECT 204.600 127.900 206.600 128.000 ;
        RECT 207.000 127.900 207.400 129.900 ;
        RECT 209.400 128.500 209.800 129.500 ;
        RECT 204.700 127.700 206.500 127.900 ;
        RECT 202.200 127.300 203.300 127.600 ;
        RECT 195.000 125.800 195.400 127.200 ;
        RECT 196.700 126.900 197.100 127.200 ;
        RECT 198.300 126.900 198.700 127.200 ;
        RECT 200.100 126.900 200.500 127.200 ;
        RECT 201.400 126.900 201.800 127.200 ;
        RECT 195.800 126.500 197.100 126.900 ;
        RECT 197.500 126.500 198.700 126.900 ;
        RECT 199.200 126.500 200.500 126.900 ;
        RECT 200.900 126.500 201.800 126.900 ;
        RECT 196.700 125.800 197.100 126.500 ;
        RECT 198.300 125.800 198.700 126.500 ;
        RECT 200.100 125.800 200.500 126.500 ;
        RECT 202.200 125.800 202.600 126.600 ;
        RECT 203.000 125.800 203.300 127.300 ;
        RECT 205.000 127.200 205.400 127.400 ;
        RECT 207.000 127.200 207.300 127.900 ;
        RECT 209.400 127.400 209.700 128.500 ;
        RECT 211.500 128.000 211.900 129.500 ;
        RECT 211.500 127.700 212.300 128.000 ;
        RECT 211.900 127.500 212.300 127.700 ;
        RECT 204.600 126.900 205.400 127.200 ;
        RECT 204.600 126.800 205.000 126.900 ;
        RECT 206.100 126.800 207.400 127.200 ;
        RECT 209.400 127.100 211.500 127.400 ;
        RECT 211.000 126.900 211.500 127.100 ;
        RECT 212.000 127.200 212.300 127.500 ;
        RECT 212.000 127.100 213.000 127.200 ;
        RECT 213.400 127.100 213.800 127.200 ;
        RECT 205.400 125.800 205.800 126.600 ;
        RECT 195.000 125.400 196.200 125.800 ;
        RECT 196.700 125.400 197.800 125.800 ;
        RECT 198.300 125.400 199.400 125.800 ;
        RECT 200.100 125.400 201.000 125.800 ;
        RECT 191.000 124.900 192.200 125.200 ;
        RECT 190.700 124.500 191.100 124.600 ;
        RECT 190.000 124.200 191.100 124.500 ;
        RECT 191.900 124.400 192.200 124.900 ;
        RECT 191.900 124.000 192.600 124.400 ;
        RECT 188.700 123.700 189.100 123.800 ;
        RECT 190.100 123.700 190.500 123.800 ;
        RECT 187.000 123.100 187.400 123.500 ;
        RECT 188.700 123.400 190.500 123.700 ;
        RECT 189.800 123.100 190.100 123.400 ;
        RECT 191.800 123.100 192.200 123.500 ;
        RECT 187.000 122.800 188.000 123.100 ;
        RECT 187.600 121.100 188.000 122.800 ;
        RECT 189.800 121.100 190.200 123.100 ;
        RECT 191.900 121.100 192.500 123.100 ;
        RECT 194.200 121.100 194.600 125.400 ;
        RECT 195.800 121.100 196.200 125.400 ;
        RECT 197.400 121.100 197.800 125.400 ;
        RECT 199.000 121.100 199.400 125.400 ;
        RECT 200.600 121.100 201.000 125.400 ;
        RECT 203.000 125.400 203.600 125.800 ;
        RECT 203.000 125.100 203.300 125.400 ;
        RECT 206.100 125.100 206.400 126.800 ;
        RECT 209.400 125.800 209.800 126.600 ;
        RECT 210.200 125.800 210.600 126.600 ;
        RECT 211.000 126.500 211.700 126.900 ;
        RECT 212.000 126.800 213.800 127.100 ;
        RECT 211.000 125.500 211.300 126.500 ;
        RECT 209.400 125.200 211.300 125.500 ;
        RECT 207.000 125.100 207.400 125.200 ;
        RECT 202.200 124.800 203.300 125.100 ;
        RECT 205.900 124.800 206.400 125.100 ;
        RECT 206.700 124.800 207.400 125.100 ;
        RECT 202.200 121.100 202.600 124.800 ;
        RECT 205.900 122.200 206.300 124.800 ;
        RECT 206.700 124.200 207.000 124.800 ;
        RECT 206.600 123.800 207.000 124.200 ;
        RECT 205.400 121.800 206.300 122.200 ;
        RECT 205.900 121.100 206.300 121.800 ;
        RECT 209.400 123.500 209.700 125.200 ;
        RECT 212.000 124.900 212.300 126.800 ;
        RECT 212.600 126.100 213.000 126.200 ;
        RECT 214.200 126.100 214.600 129.900 ;
        RECT 215.000 127.800 215.400 128.600 ;
        RECT 215.800 127.500 216.200 129.900 ;
        RECT 218.000 129.200 218.400 129.900 ;
        RECT 217.400 128.900 218.400 129.200 ;
        RECT 220.200 128.900 220.600 129.900 ;
        RECT 222.300 129.200 222.900 129.900 ;
        RECT 222.200 128.900 222.900 129.200 ;
        RECT 217.400 128.500 217.800 128.900 ;
        RECT 220.200 128.600 220.500 128.900 ;
        RECT 218.200 128.200 218.600 128.600 ;
        RECT 219.100 128.300 220.500 128.600 ;
        RECT 222.200 128.500 222.600 128.900 ;
        RECT 219.100 128.200 219.500 128.300 ;
        RECT 216.200 127.100 217.000 127.200 ;
        RECT 218.300 127.100 218.600 128.200 ;
        RECT 223.100 127.700 223.500 127.800 ;
        RECT 224.600 127.700 225.000 129.900 ;
        RECT 223.100 127.400 225.000 127.700 ;
        RECT 221.100 127.100 221.500 127.200 ;
        RECT 216.200 126.800 221.700 127.100 ;
        RECT 217.700 126.700 218.100 126.800 ;
        RECT 212.600 125.800 214.600 126.100 ;
        RECT 216.900 126.200 217.300 126.300 ;
        RECT 221.400 126.200 221.700 126.800 ;
        RECT 222.200 126.400 222.600 126.500 ;
        RECT 216.900 125.900 219.400 126.200 ;
        RECT 219.000 125.800 219.400 125.900 ;
        RECT 221.400 125.800 221.800 126.200 ;
        RECT 222.200 126.100 224.100 126.400 ;
        RECT 223.700 126.000 224.100 126.100 ;
        RECT 212.600 125.400 213.000 125.800 ;
        RECT 211.500 124.600 212.300 124.900 ;
        RECT 209.400 121.500 209.800 123.500 ;
        RECT 211.500 121.100 211.900 124.600 ;
        RECT 214.200 121.100 214.600 125.800 ;
        RECT 215.800 125.500 218.600 125.600 ;
        RECT 215.800 125.400 218.700 125.500 ;
        RECT 215.800 125.300 220.700 125.400 ;
        RECT 215.800 121.100 216.200 125.300 ;
        RECT 218.300 125.100 220.700 125.300 ;
        RECT 217.400 124.500 220.100 124.800 ;
        RECT 217.400 124.400 217.800 124.500 ;
        RECT 219.700 124.400 220.100 124.500 ;
        RECT 220.400 124.500 220.700 125.100 ;
        RECT 221.400 125.200 221.700 125.800 ;
        RECT 222.900 125.700 223.300 125.800 ;
        RECT 224.600 125.700 225.000 127.400 ;
        RECT 225.400 128.500 225.800 129.500 ;
        RECT 227.500 129.200 227.900 129.500 ;
        RECT 227.000 128.800 227.900 129.200 ;
        RECT 225.400 127.400 225.700 128.500 ;
        RECT 227.500 128.000 227.900 128.800 ;
        RECT 227.500 127.700 228.300 128.000 ;
        RECT 230.200 127.800 230.600 128.600 ;
        RECT 227.900 127.500 228.300 127.700 ;
        RECT 225.400 127.100 227.500 127.400 ;
        RECT 227.000 126.900 227.500 127.100 ;
        RECT 228.000 127.200 228.300 127.500 ;
        RECT 225.400 125.800 225.800 126.600 ;
        RECT 226.200 125.800 226.600 126.600 ;
        RECT 227.000 126.500 227.700 126.900 ;
        RECT 228.000 126.800 229.000 127.200 ;
        RECT 222.900 125.400 225.000 125.700 ;
        RECT 227.000 125.500 227.300 126.500 ;
        RECT 221.400 124.900 222.600 125.200 ;
        RECT 221.100 124.500 221.500 124.600 ;
        RECT 220.400 124.200 221.500 124.500 ;
        RECT 222.300 124.400 222.600 124.900 ;
        RECT 222.300 124.000 223.000 124.400 ;
        RECT 219.100 123.700 219.500 123.800 ;
        RECT 220.500 123.700 220.900 123.800 ;
        RECT 217.400 123.100 217.800 123.500 ;
        RECT 219.100 123.400 220.900 123.700 ;
        RECT 220.200 123.100 220.500 123.400 ;
        RECT 222.200 123.100 222.600 123.500 ;
        RECT 217.400 122.800 218.400 123.100 ;
        RECT 218.000 121.100 218.400 122.800 ;
        RECT 220.200 121.100 220.600 123.100 ;
        RECT 222.300 121.100 222.900 123.100 ;
        RECT 224.600 121.100 225.000 125.400 ;
        RECT 225.400 125.200 227.300 125.500 ;
        RECT 225.400 123.500 225.700 125.200 ;
        RECT 228.000 124.900 228.300 126.800 ;
        RECT 228.600 125.400 229.000 126.200 ;
        RECT 229.400 126.100 229.800 126.200 ;
        RECT 231.000 126.100 231.400 129.900 ;
        RECT 229.400 125.800 231.400 126.100 ;
        RECT 227.500 124.600 228.300 124.900 ;
        RECT 225.400 121.500 225.800 123.500 ;
        RECT 227.500 121.100 227.900 124.600 ;
        RECT 231.000 121.100 231.400 125.800 ;
        RECT 231.800 127.700 232.200 129.900 ;
        RECT 233.900 129.200 234.500 129.900 ;
        RECT 233.900 128.900 234.600 129.200 ;
        RECT 236.200 128.900 236.600 129.900 ;
        RECT 238.400 129.200 238.800 129.900 ;
        RECT 238.400 128.900 239.400 129.200 ;
        RECT 234.200 128.500 234.600 128.900 ;
        RECT 236.300 128.600 236.600 128.900 ;
        RECT 236.300 128.300 237.700 128.600 ;
        RECT 237.300 128.200 237.700 128.300 ;
        RECT 238.200 128.200 238.600 128.600 ;
        RECT 239.000 128.500 239.400 128.900 ;
        RECT 233.300 127.700 233.700 127.800 ;
        RECT 231.800 127.400 233.700 127.700 ;
        RECT 231.800 125.700 232.200 127.400 ;
        RECT 235.300 127.100 235.700 127.200 ;
        RECT 238.200 127.100 238.500 128.200 ;
        RECT 240.600 127.500 241.000 129.900 ;
        RECT 242.200 128.200 242.600 129.900 ;
        RECT 242.100 127.900 242.600 128.200 ;
        RECT 242.100 127.200 242.400 127.900 ;
        RECT 243.800 127.600 244.200 129.900 ;
        RECT 244.600 128.000 245.000 129.900 ;
        RECT 246.200 128.000 246.600 129.900 ;
        RECT 244.600 127.900 246.600 128.000 ;
        RECT 247.000 127.900 247.400 129.900 ;
        RECT 248.100 128.200 248.500 129.900 ;
        RECT 248.100 127.900 249.000 128.200 ;
        RECT 244.700 127.700 246.500 127.900 ;
        RECT 242.900 127.300 244.200 127.600 ;
        RECT 239.800 127.100 240.600 127.200 ;
        RECT 235.100 126.800 240.600 127.100 ;
        RECT 242.100 126.800 242.600 127.200 ;
        RECT 234.200 126.400 234.600 126.500 ;
        RECT 232.700 126.100 234.600 126.400 ;
        RECT 235.100 126.200 235.400 126.800 ;
        RECT 238.700 126.700 239.100 126.800 ;
        RECT 239.500 126.200 239.900 126.300 ;
        RECT 232.700 126.000 233.100 126.100 ;
        RECT 235.000 125.800 235.400 126.200 ;
        RECT 237.400 125.900 239.900 126.200 ;
        RECT 237.400 125.800 237.800 125.900 ;
        RECT 233.500 125.700 233.900 125.800 ;
        RECT 231.800 125.400 233.900 125.700 ;
        RECT 231.800 121.100 232.200 125.400 ;
        RECT 235.100 125.200 235.400 125.800 ;
        RECT 238.200 125.500 241.000 125.600 ;
        RECT 238.100 125.400 241.000 125.500 ;
        RECT 234.200 124.900 235.400 125.200 ;
        RECT 236.100 125.300 241.000 125.400 ;
        RECT 236.100 125.100 238.500 125.300 ;
        RECT 234.200 124.400 234.500 124.900 ;
        RECT 233.800 124.000 234.500 124.400 ;
        RECT 235.300 124.500 235.700 124.600 ;
        RECT 236.100 124.500 236.400 125.100 ;
        RECT 235.300 124.200 236.400 124.500 ;
        RECT 236.700 124.500 239.400 124.800 ;
        RECT 236.700 124.400 237.100 124.500 ;
        RECT 239.000 124.400 239.400 124.500 ;
        RECT 235.900 123.700 236.300 123.800 ;
        RECT 237.300 123.700 237.700 123.800 ;
        RECT 234.200 123.100 234.600 123.500 ;
        RECT 235.900 123.400 237.700 123.700 ;
        RECT 236.300 123.100 236.600 123.400 ;
        RECT 239.000 123.100 239.400 123.500 ;
        RECT 233.900 121.100 234.500 123.100 ;
        RECT 236.200 121.100 236.600 123.100 ;
        RECT 238.400 122.800 239.400 123.100 ;
        RECT 238.400 121.100 238.800 122.800 ;
        RECT 240.600 121.100 241.000 125.300 ;
        RECT 242.100 125.100 242.400 126.800 ;
        RECT 242.900 126.500 243.200 127.300 ;
        RECT 245.000 127.200 245.400 127.400 ;
        RECT 247.000 127.200 247.300 127.900 ;
        RECT 244.600 126.900 245.400 127.200 ;
        RECT 246.100 127.100 247.400 127.200 ;
        RECT 247.800 127.100 248.200 127.200 ;
        RECT 244.600 126.800 245.000 126.900 ;
        RECT 246.100 126.800 248.200 127.100 ;
        RECT 242.700 126.100 243.200 126.500 ;
        RECT 242.900 125.100 243.200 126.100 ;
        RECT 243.700 126.200 244.100 126.600 ;
        RECT 243.700 125.800 244.200 126.200 ;
        RECT 245.400 125.800 245.800 126.600 ;
        RECT 246.100 125.100 246.400 126.800 ;
        RECT 248.600 126.100 249.000 127.900 ;
        RECT 250.200 127.700 250.600 129.900 ;
        RECT 252.300 129.200 252.900 129.900 ;
        RECT 252.300 128.900 253.000 129.200 ;
        RECT 254.600 128.900 255.000 129.900 ;
        RECT 256.800 129.200 257.200 129.900 ;
        RECT 256.800 128.900 257.800 129.200 ;
        RECT 252.600 128.500 253.000 128.900 ;
        RECT 254.700 128.600 255.000 128.900 ;
        RECT 254.700 128.300 256.100 128.600 ;
        RECT 255.700 128.200 256.100 128.300 ;
        RECT 256.600 128.200 257.000 128.600 ;
        RECT 257.400 128.500 257.800 128.900 ;
        RECT 251.700 127.700 252.100 127.800 ;
        RECT 249.400 127.100 249.800 127.600 ;
        RECT 250.200 127.400 252.100 127.700 ;
        RECT 250.200 127.100 250.600 127.400 ;
        RECT 253.700 127.100 254.100 127.200 ;
        RECT 256.600 127.100 256.900 128.200 ;
        RECT 259.000 127.500 259.400 129.900 ;
        RECT 259.800 127.600 260.200 129.900 ;
        RECT 263.000 129.100 263.400 129.200 ;
        RECT 264.000 129.100 264.400 129.900 ;
        RECT 263.000 128.800 264.400 129.100 ;
        RECT 259.800 127.300 260.900 127.600 ;
        RECT 258.200 127.100 259.000 127.200 ;
        RECT 249.400 126.800 250.600 127.100 ;
        RECT 247.000 125.800 249.000 126.100 ;
        RECT 247.000 125.200 247.300 125.800 ;
        RECT 247.000 125.100 247.400 125.200 ;
        RECT 242.100 124.600 242.600 125.100 ;
        RECT 242.900 124.800 244.200 125.100 ;
        RECT 242.200 121.100 242.600 124.600 ;
        RECT 243.800 121.100 244.200 124.800 ;
        RECT 245.900 124.800 246.400 125.100 ;
        RECT 246.700 124.800 247.400 125.100 ;
        RECT 245.900 121.100 246.300 124.800 ;
        RECT 246.700 124.200 247.000 124.800 ;
        RECT 247.800 124.400 248.200 125.200 ;
        RECT 246.600 123.800 247.000 124.200 ;
        RECT 248.600 121.100 249.000 125.800 ;
        RECT 250.200 125.700 250.600 126.800 ;
        RECT 253.500 126.800 259.000 127.100 ;
        RECT 252.600 126.400 253.000 126.500 ;
        RECT 251.100 126.100 253.000 126.400 ;
        RECT 253.500 126.100 253.800 126.800 ;
        RECT 257.100 126.700 257.500 126.800 ;
        RECT 257.900 126.200 258.300 126.300 ;
        RECT 254.200 126.100 254.600 126.200 ;
        RECT 251.100 126.000 251.500 126.100 ;
        RECT 253.400 125.800 254.600 126.100 ;
        RECT 255.800 125.900 258.300 126.200 ;
        RECT 255.800 125.800 256.200 125.900 ;
        RECT 259.800 125.800 260.200 126.600 ;
        RECT 260.600 125.800 260.900 127.300 ;
        RECT 264.000 127.100 264.400 128.800 ;
        RECT 264.000 126.900 264.900 127.100 ;
        RECT 264.100 126.800 264.900 126.900 ;
        RECT 251.900 125.700 252.300 125.800 ;
        RECT 250.200 125.400 252.300 125.700 ;
        RECT 250.200 121.100 250.600 125.400 ;
        RECT 253.500 125.200 253.800 125.800 ;
        RECT 256.600 125.500 259.400 125.600 ;
        RECT 256.500 125.400 259.400 125.500 ;
        RECT 252.600 124.900 253.800 125.200 ;
        RECT 254.500 125.300 259.400 125.400 ;
        RECT 254.500 125.100 256.900 125.300 ;
        RECT 252.600 124.400 252.900 124.900 ;
        RECT 252.200 124.000 252.900 124.400 ;
        RECT 253.700 124.500 254.100 124.600 ;
        RECT 254.500 124.500 254.800 125.100 ;
        RECT 253.700 124.200 254.800 124.500 ;
        RECT 255.100 124.500 257.800 124.800 ;
        RECT 255.100 124.400 255.500 124.500 ;
        RECT 257.400 124.400 257.800 124.500 ;
        RECT 254.300 123.700 254.700 123.800 ;
        RECT 255.700 123.700 256.100 123.800 ;
        RECT 252.600 123.100 253.000 123.500 ;
        RECT 254.300 123.400 256.100 123.700 ;
        RECT 254.700 123.100 255.000 123.400 ;
        RECT 257.400 123.100 257.800 123.500 ;
        RECT 252.300 121.100 252.900 123.100 ;
        RECT 254.600 121.100 255.000 123.100 ;
        RECT 256.800 122.800 257.800 123.100 ;
        RECT 256.800 121.100 257.200 122.800 ;
        RECT 259.000 121.100 259.400 125.300 ;
        RECT 260.600 125.400 261.200 125.800 ;
        RECT 260.600 125.100 260.900 125.400 ;
        RECT 259.800 124.800 260.900 125.100 ;
        RECT 264.600 125.200 264.900 126.800 ;
        RECT 264.600 124.800 265.000 125.200 ;
        RECT 259.800 121.100 260.200 124.800 ;
        RECT 264.600 123.500 264.900 124.800 ;
        RECT 263.100 123.200 264.900 123.500 ;
        RECT 263.100 123.100 263.400 123.200 ;
        RECT 263.000 121.100 263.400 123.100 ;
        RECT 264.600 123.100 264.900 123.200 ;
        RECT 264.600 121.100 265.000 123.100 ;
        RECT 1.400 115.600 1.800 119.900 ;
        RECT 3.000 115.600 3.400 119.900 ;
        RECT 4.600 115.600 5.000 119.900 ;
        RECT 6.200 115.600 6.600 119.900 ;
        RECT 7.800 115.700 8.200 119.900 ;
        RECT 10.000 118.200 10.400 119.900 ;
        RECT 9.400 117.900 10.400 118.200 ;
        RECT 12.200 117.900 12.600 119.900 ;
        RECT 14.300 117.900 14.900 119.900 ;
        RECT 9.400 117.500 9.800 117.900 ;
        RECT 12.200 117.600 12.500 117.900 ;
        RECT 11.100 117.300 12.900 117.600 ;
        RECT 14.200 117.500 14.600 117.900 ;
        RECT 11.100 117.200 11.500 117.300 ;
        RECT 12.500 117.200 12.900 117.300 ;
        RECT 9.400 116.500 9.800 116.600 ;
        RECT 11.700 116.500 12.100 116.600 ;
        RECT 9.400 116.200 12.100 116.500 ;
        RECT 12.400 116.500 13.500 116.800 ;
        RECT 12.400 115.900 12.700 116.500 ;
        RECT 13.100 116.400 13.500 116.500 ;
        RECT 14.300 116.600 15.000 117.000 ;
        RECT 14.300 116.100 14.600 116.600 ;
        RECT 10.300 115.700 12.700 115.900 ;
        RECT 7.800 115.600 12.700 115.700 ;
        RECT 13.400 115.800 14.600 116.100 ;
        RECT 1.400 115.200 2.300 115.600 ;
        RECT 3.000 115.200 4.100 115.600 ;
        RECT 4.600 115.200 5.700 115.600 ;
        RECT 6.200 115.200 7.400 115.600 ;
        RECT 7.800 115.500 10.700 115.600 ;
        RECT 7.800 115.400 10.600 115.500 ;
        RECT 1.900 114.500 2.300 115.200 ;
        RECT 3.700 114.500 4.100 115.200 ;
        RECT 5.300 114.500 5.700 115.200 ;
        RECT 1.900 114.100 3.200 114.500 ;
        RECT 3.700 114.100 4.900 114.500 ;
        RECT 5.300 114.100 6.600 114.500 ;
        RECT 1.900 113.800 2.300 114.100 ;
        RECT 3.700 113.800 4.100 114.100 ;
        RECT 5.300 113.800 5.700 114.100 ;
        RECT 7.000 113.800 7.400 115.200 ;
        RECT 11.000 115.100 11.400 115.200 ;
        RECT 11.800 115.100 12.200 115.200 ;
        RECT 8.900 114.800 12.200 115.100 ;
        RECT 8.900 114.700 9.300 114.800 ;
        RECT 9.700 114.200 10.100 114.300 ;
        RECT 13.400 114.200 13.700 115.800 ;
        RECT 16.600 115.600 17.000 119.900 ;
        RECT 18.700 117.200 19.100 119.900 ;
        RECT 18.200 116.800 19.100 117.200 ;
        RECT 19.400 116.800 19.800 117.200 ;
        RECT 18.700 116.200 19.100 116.800 ;
        RECT 19.500 116.200 19.800 116.800 ;
        RECT 18.700 115.900 19.200 116.200 ;
        RECT 19.500 115.900 20.200 116.200 ;
        RECT 14.900 115.300 17.000 115.600 ;
        RECT 14.900 115.200 15.300 115.300 ;
        RECT 15.700 114.900 16.100 115.000 ;
        RECT 14.200 114.600 16.100 114.900 ;
        RECT 14.200 114.500 14.600 114.600 ;
        RECT 8.200 113.900 13.700 114.200 ;
        RECT 8.200 113.800 9.000 113.900 ;
        RECT 1.400 113.400 2.300 113.800 ;
        RECT 3.000 113.400 4.100 113.800 ;
        RECT 4.600 113.400 5.700 113.800 ;
        RECT 6.200 113.400 7.400 113.800 ;
        RECT 1.400 111.100 1.800 113.400 ;
        RECT 3.000 111.100 3.400 113.400 ;
        RECT 4.600 111.100 5.000 113.400 ;
        RECT 6.200 111.100 6.600 113.400 ;
        RECT 7.800 111.100 8.200 113.500 ;
        RECT 10.300 112.800 10.600 113.900 ;
        RECT 13.100 113.800 13.500 113.900 ;
        RECT 16.600 113.600 17.000 115.300 ;
        RECT 18.200 114.400 18.600 115.200 ;
        RECT 18.900 114.200 19.200 115.900 ;
        RECT 19.800 115.800 20.200 115.900 ;
        RECT 20.600 115.800 21.000 116.600 ;
        RECT 19.800 115.100 20.100 115.800 ;
        RECT 21.400 115.100 21.800 119.900 ;
        RECT 23.000 117.500 23.400 119.500 ;
        RECT 25.100 119.200 25.500 119.900 ;
        RECT 25.100 118.800 25.800 119.200 ;
        RECT 23.000 115.800 23.300 117.500 ;
        RECT 25.100 116.400 25.500 118.800 ;
        RECT 25.100 116.100 25.900 116.400 ;
        RECT 23.000 115.500 24.900 115.800 ;
        RECT 19.800 114.800 21.800 115.100 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 17.400 113.800 18.200 114.100 ;
        RECT 18.900 113.800 20.200 114.200 ;
        RECT 17.800 113.600 18.200 113.800 ;
        RECT 15.100 113.300 17.000 113.600 ;
        RECT 15.100 113.200 15.500 113.300 ;
        RECT 9.400 112.100 9.800 112.500 ;
        RECT 10.200 112.400 10.600 112.800 ;
        RECT 11.100 112.700 11.500 112.800 ;
        RECT 11.100 112.400 12.500 112.700 ;
        RECT 12.200 112.100 12.500 112.400 ;
        RECT 14.200 112.100 14.600 112.500 ;
        RECT 9.400 111.800 10.400 112.100 ;
        RECT 10.000 111.100 10.400 111.800 ;
        RECT 12.200 111.100 12.600 112.100 ;
        RECT 14.200 111.800 14.900 112.100 ;
        RECT 14.300 111.100 14.900 111.800 ;
        RECT 16.600 111.100 17.000 113.300 ;
        RECT 17.500 113.100 19.300 113.300 ;
        RECT 19.800 113.100 20.100 113.800 ;
        RECT 21.400 113.100 21.800 114.800 ;
        RECT 23.000 114.400 23.400 115.200 ;
        RECT 23.800 114.400 24.200 115.200 ;
        RECT 24.600 114.500 24.900 115.500 ;
        RECT 22.200 113.400 22.600 114.200 ;
        RECT 24.600 114.100 25.300 114.500 ;
        RECT 25.600 114.200 25.900 116.100 ;
        RECT 27.800 116.200 28.200 119.900 ;
        RECT 29.400 116.200 29.800 119.900 ;
        RECT 27.800 115.900 29.800 116.200 ;
        RECT 30.200 115.900 30.600 119.900 ;
        RECT 32.300 116.300 32.700 119.900 ;
        RECT 34.200 116.400 34.600 119.900 ;
        RECT 31.800 115.900 32.700 116.300 ;
        RECT 34.100 115.900 34.600 116.400 ;
        RECT 35.800 116.200 36.200 119.900 ;
        RECT 34.900 115.900 36.200 116.200 ;
        RECT 36.600 117.500 37.000 119.500 ;
        RECT 26.200 115.100 26.600 115.600 ;
        RECT 28.200 115.200 28.600 115.400 ;
        RECT 30.200 115.200 30.500 115.900 ;
        RECT 27.000 115.100 27.400 115.200 ;
        RECT 26.200 114.800 27.400 115.100 ;
        RECT 27.800 114.900 28.600 115.200 ;
        RECT 29.400 114.900 30.600 115.200 ;
        RECT 27.800 114.800 28.200 114.900 ;
        RECT 24.600 113.900 25.100 114.100 ;
        RECT 23.000 113.600 25.100 113.900 ;
        RECT 25.600 113.800 26.600 114.200 ;
        RECT 28.600 113.800 29.000 114.600 ;
        RECT 17.400 113.000 19.400 113.100 ;
        RECT 17.400 111.100 17.800 113.000 ;
        RECT 19.000 111.100 19.400 113.000 ;
        RECT 19.800 111.100 20.200 113.100 ;
        RECT 20.900 112.800 21.800 113.100 ;
        RECT 20.900 111.100 21.300 112.800 ;
        RECT 23.000 112.500 23.300 113.600 ;
        RECT 25.600 113.500 25.900 113.800 ;
        RECT 25.500 113.300 25.900 113.500 ;
        RECT 25.100 113.000 25.900 113.300 ;
        RECT 29.400 113.100 29.700 114.900 ;
        RECT 30.200 114.800 30.600 114.900 ;
        RECT 31.900 114.200 32.200 115.900 ;
        RECT 32.600 115.100 33.000 115.600 ;
        RECT 33.400 115.100 33.800 115.200 ;
        RECT 32.600 114.800 33.800 115.100 ;
        RECT 31.800 114.100 32.200 114.200 ;
        RECT 30.200 113.800 32.200 114.100 ;
        RECT 30.200 113.200 30.500 113.800 ;
        RECT 23.000 111.500 23.400 112.500 ;
        RECT 25.100 111.500 25.500 113.000 ;
        RECT 29.400 111.100 29.800 113.100 ;
        RECT 30.200 112.800 30.600 113.200 ;
        RECT 30.100 112.400 30.500 112.800 ;
        RECT 31.000 112.400 31.400 113.200 ;
        RECT 31.900 112.100 32.200 113.800 ;
        RECT 34.100 114.200 34.400 115.900 ;
        RECT 34.900 114.900 35.200 115.900 ;
        RECT 36.600 115.800 36.900 117.500 ;
        RECT 38.700 116.400 39.100 119.900 ;
        RECT 38.700 116.100 39.500 116.400 ;
        RECT 36.600 115.500 38.500 115.800 ;
        RECT 34.700 114.500 35.200 114.900 ;
        RECT 34.100 113.800 34.600 114.200 ;
        RECT 34.100 113.100 34.400 113.800 ;
        RECT 34.900 113.700 35.200 114.500 ;
        RECT 35.700 114.800 36.200 115.200 ;
        RECT 35.700 114.400 36.100 114.800 ;
        RECT 36.600 114.400 37.000 115.200 ;
        RECT 37.400 114.400 37.800 115.200 ;
        RECT 38.200 114.500 38.500 115.500 ;
        RECT 38.200 114.100 38.900 114.500 ;
        RECT 39.200 114.200 39.500 116.100 ;
        RECT 39.800 115.100 40.200 115.600 ;
        RECT 41.400 115.100 41.800 119.900 ;
        RECT 39.800 114.800 41.800 115.100 ;
        RECT 39.200 114.100 40.200 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 38.200 113.900 38.700 114.100 ;
        RECT 34.900 113.400 36.200 113.700 ;
        RECT 34.100 112.800 34.600 113.100 ;
        RECT 31.800 111.100 32.200 112.100 ;
        RECT 34.200 111.100 34.600 112.800 ;
        RECT 35.800 111.100 36.200 113.400 ;
        RECT 36.600 113.600 38.700 113.900 ;
        RECT 39.200 113.800 41.000 114.100 ;
        RECT 36.600 112.500 36.900 113.600 ;
        RECT 39.200 113.500 39.500 113.800 ;
        RECT 39.100 113.300 39.500 113.500 ;
        RECT 38.700 113.000 39.500 113.300 ;
        RECT 36.600 111.500 37.000 112.500 ;
        RECT 38.700 111.500 39.100 113.000 ;
        RECT 41.400 111.100 41.800 114.800 ;
        RECT 43.000 115.600 43.400 119.900 ;
        RECT 45.100 117.900 45.700 119.900 ;
        RECT 47.400 117.900 47.800 119.900 ;
        RECT 49.600 118.200 50.000 119.900 ;
        RECT 49.600 117.900 50.600 118.200 ;
        RECT 45.400 117.500 45.800 117.900 ;
        RECT 47.500 117.600 47.800 117.900 ;
        RECT 47.100 117.300 48.900 117.600 ;
        RECT 50.200 117.500 50.600 117.900 ;
        RECT 47.100 117.200 47.500 117.300 ;
        RECT 48.500 117.200 48.900 117.300 ;
        RECT 45.000 116.600 45.700 117.000 ;
        RECT 45.400 116.100 45.700 116.600 ;
        RECT 46.500 116.500 47.600 116.800 ;
        RECT 46.500 116.400 46.900 116.500 ;
        RECT 45.400 115.800 46.600 116.100 ;
        RECT 43.000 115.300 45.100 115.600 ;
        RECT 43.000 113.600 43.400 115.300 ;
        RECT 44.700 115.200 45.100 115.300 ;
        RECT 43.900 114.900 44.300 115.000 ;
        RECT 43.900 114.600 45.800 114.900 ;
        RECT 45.400 114.500 45.800 114.600 ;
        RECT 46.300 114.200 46.600 115.800 ;
        RECT 47.300 115.900 47.600 116.500 ;
        RECT 47.900 116.500 48.300 116.600 ;
        RECT 50.200 116.500 50.600 116.600 ;
        RECT 47.900 116.200 50.600 116.500 ;
        RECT 47.300 115.700 49.700 115.900 ;
        RECT 51.800 115.700 52.200 119.900 ;
        RECT 52.600 116.200 53.000 119.900 ;
        RECT 54.200 116.200 54.600 119.900 ;
        RECT 52.600 115.900 54.600 116.200 ;
        RECT 55.000 115.900 55.400 119.900 ;
        RECT 57.700 116.300 58.100 119.900 ;
        RECT 57.700 115.900 58.600 116.300 ;
        RECT 47.300 115.600 52.200 115.700 ;
        RECT 49.300 115.500 52.200 115.600 ;
        RECT 49.400 115.400 52.200 115.500 ;
        RECT 53.000 115.200 53.400 115.400 ;
        RECT 55.000 115.200 55.300 115.900 ;
        RECT 48.600 115.100 49.000 115.200 ;
        RECT 48.600 114.800 51.100 115.100 ;
        RECT 52.600 114.900 53.400 115.200 ;
        RECT 54.200 114.900 55.400 115.200 ;
        RECT 52.600 114.800 53.000 114.900 ;
        RECT 50.700 114.700 51.100 114.800 ;
        RECT 49.900 114.200 50.300 114.300 ;
        RECT 46.300 113.900 51.800 114.200 ;
        RECT 46.500 113.800 46.900 113.900 ;
        RECT 49.400 113.800 49.800 113.900 ;
        RECT 51.000 113.800 51.800 113.900 ;
        RECT 53.400 113.800 53.800 114.600 ;
        RECT 43.000 113.300 44.900 113.600 ;
        RECT 42.200 113.100 42.600 113.200 ;
        RECT 43.000 113.100 43.400 113.300 ;
        RECT 44.500 113.200 44.900 113.300 ;
        RECT 42.200 112.800 43.400 113.100 ;
        RECT 49.400 112.800 49.700 113.800 ;
        RECT 42.200 112.400 42.600 112.800 ;
        RECT 43.000 111.100 43.400 112.800 ;
        RECT 48.500 112.700 48.900 112.800 ;
        RECT 45.400 112.100 45.800 112.500 ;
        RECT 47.500 112.400 48.900 112.700 ;
        RECT 49.400 112.400 49.800 112.800 ;
        RECT 47.500 112.100 47.800 112.400 ;
        RECT 50.200 112.100 50.600 112.500 ;
        RECT 45.100 111.800 45.800 112.100 ;
        RECT 45.100 111.100 45.700 111.800 ;
        RECT 47.400 111.100 47.800 112.100 ;
        RECT 49.600 111.800 50.600 112.100 ;
        RECT 49.600 111.100 50.000 111.800 ;
        RECT 51.800 111.100 52.200 113.500 ;
        RECT 54.200 113.100 54.500 114.900 ;
        RECT 55.000 114.800 55.400 114.900 ;
        RECT 57.400 114.800 57.800 115.600 ;
        RECT 58.200 114.200 58.500 115.900 ;
        RECT 59.800 115.700 60.200 119.900 ;
        RECT 62.000 118.200 62.400 119.900 ;
        RECT 61.400 117.900 62.400 118.200 ;
        RECT 64.200 117.900 64.600 119.900 ;
        RECT 66.300 117.900 66.900 119.900 ;
        RECT 61.400 117.500 61.800 117.900 ;
        RECT 64.200 117.600 64.500 117.900 ;
        RECT 63.100 117.300 64.900 117.600 ;
        RECT 66.200 117.500 66.600 117.900 ;
        RECT 63.100 117.200 63.500 117.300 ;
        RECT 64.500 117.200 64.900 117.300 ;
        RECT 61.400 116.500 61.800 116.600 ;
        RECT 63.700 116.500 64.100 116.600 ;
        RECT 61.400 116.200 64.100 116.500 ;
        RECT 64.400 116.500 65.500 116.800 ;
        RECT 64.400 115.900 64.700 116.500 ;
        RECT 65.100 116.400 65.500 116.500 ;
        RECT 66.300 116.600 67.000 117.000 ;
        RECT 66.300 116.100 66.600 116.600 ;
        RECT 62.300 115.700 64.700 115.900 ;
        RECT 59.800 115.600 64.700 115.700 ;
        RECT 65.400 115.800 66.600 116.100 ;
        RECT 59.800 115.500 62.700 115.600 ;
        RECT 59.800 115.400 62.600 115.500 ;
        RECT 63.000 115.100 63.400 115.200 ;
        RECT 64.600 115.100 65.000 115.200 ;
        RECT 60.900 114.800 65.000 115.100 ;
        RECT 60.900 114.700 61.300 114.800 ;
        RECT 61.700 114.200 62.100 114.300 ;
        RECT 65.400 114.200 65.700 115.800 ;
        RECT 68.600 115.600 69.000 119.900 ;
        RECT 70.700 116.200 71.100 119.900 ;
        RECT 71.400 116.800 71.800 117.200 ;
        RECT 71.500 116.200 71.800 116.800 ;
        RECT 70.700 115.900 71.200 116.200 ;
        RECT 71.500 116.100 72.200 116.200 ;
        RECT 73.400 116.100 73.800 119.900 ;
        RECT 75.000 117.500 75.400 119.500 ;
        RECT 77.100 119.200 77.500 119.900 ;
        RECT 76.600 118.800 77.500 119.200 ;
        RECT 71.500 115.900 73.800 116.100 ;
        RECT 66.900 115.300 69.000 115.600 ;
        RECT 66.900 115.200 67.300 115.300 ;
        RECT 67.700 114.900 68.100 115.000 ;
        RECT 66.200 114.600 68.100 114.900 ;
        RECT 66.200 114.500 66.600 114.600 ;
        RECT 58.200 113.800 58.600 114.200 ;
        RECT 60.200 113.900 65.700 114.200 ;
        RECT 60.200 113.800 61.000 113.900 ;
        RECT 55.000 113.100 55.400 113.200 ;
        RECT 58.200 113.100 58.500 113.800 ;
        RECT 54.200 111.100 54.600 113.100 ;
        RECT 55.000 112.800 58.500 113.100 ;
        RECT 54.900 112.400 55.300 112.800 ;
        RECT 58.200 112.100 58.500 112.800 ;
        RECT 59.000 112.400 59.400 113.200 ;
        RECT 58.200 111.100 58.600 112.100 ;
        RECT 59.800 111.100 60.200 113.500 ;
        RECT 62.300 112.800 62.600 113.900 ;
        RECT 65.100 113.800 65.500 113.900 ;
        RECT 68.600 113.600 69.000 115.300 ;
        RECT 70.900 115.200 71.200 115.900 ;
        RECT 71.800 115.800 73.800 115.900 ;
        RECT 74.200 115.800 74.600 116.600 ;
        RECT 75.000 115.800 75.300 117.500 ;
        RECT 77.100 116.400 77.500 118.800 ;
        RECT 79.800 117.500 80.200 119.500 ;
        RECT 77.100 116.100 77.900 116.400 ;
        RECT 70.200 114.400 70.600 115.200 ;
        RECT 70.900 114.800 71.400 115.200 ;
        RECT 70.900 114.200 71.200 114.800 ;
        RECT 69.400 114.100 69.800 114.200 ;
        RECT 69.400 113.800 70.200 114.100 ;
        RECT 70.900 113.800 72.200 114.200 ;
        RECT 69.800 113.600 70.200 113.800 ;
        RECT 67.100 113.300 69.000 113.600 ;
        RECT 67.100 113.200 67.500 113.300 ;
        RECT 61.400 112.100 61.800 112.500 ;
        RECT 62.200 112.400 62.600 112.800 ;
        RECT 63.100 112.700 63.500 112.800 ;
        RECT 63.100 112.400 64.500 112.700 ;
        RECT 64.200 112.100 64.500 112.400 ;
        RECT 66.200 112.100 66.600 112.500 ;
        RECT 61.400 111.800 62.400 112.100 ;
        RECT 62.000 111.100 62.400 111.800 ;
        RECT 64.200 111.100 64.600 112.100 ;
        RECT 66.200 111.800 66.900 112.100 ;
        RECT 66.300 111.100 66.900 111.800 ;
        RECT 68.600 111.100 69.000 113.300 ;
        RECT 69.500 113.100 71.300 113.300 ;
        RECT 71.800 113.100 72.100 113.800 ;
        RECT 72.600 113.400 73.000 114.200 ;
        RECT 73.400 113.100 73.800 115.800 ;
        RECT 75.000 115.500 76.900 115.800 ;
        RECT 75.000 114.400 75.400 115.200 ;
        RECT 75.800 114.400 76.200 115.200 ;
        RECT 76.600 114.500 76.900 115.500 ;
        RECT 76.600 114.100 77.300 114.500 ;
        RECT 77.600 114.200 77.900 116.100 ;
        RECT 79.800 115.800 80.100 117.500 ;
        RECT 81.900 116.400 82.300 119.900 ;
        RECT 85.900 119.200 86.300 119.900 ;
        RECT 85.400 118.800 86.300 119.200 ;
        RECT 81.900 116.100 82.700 116.400 ;
        RECT 78.200 114.800 78.600 115.600 ;
        RECT 79.800 115.500 81.700 115.800 ;
        RECT 79.800 114.400 80.200 115.200 ;
        RECT 80.600 114.400 81.000 115.200 ;
        RECT 81.400 114.500 81.700 115.500 ;
        RECT 76.600 113.900 77.100 114.100 ;
        RECT 75.000 113.600 77.100 113.900 ;
        RECT 77.600 113.800 78.600 114.200 ;
        RECT 81.400 114.100 82.100 114.500 ;
        RECT 82.400 114.200 82.700 116.100 ;
        RECT 85.900 116.200 86.300 118.800 ;
        RECT 86.600 116.800 87.000 117.200 ;
        RECT 86.700 116.200 87.000 116.800 ;
        RECT 85.900 115.900 86.400 116.200 ;
        RECT 86.700 115.900 87.400 116.200 ;
        RECT 83.000 114.800 83.400 115.600 ;
        RECT 85.400 114.400 85.800 115.200 ;
        RECT 86.100 114.200 86.400 115.900 ;
        RECT 87.000 115.800 87.400 115.900 ;
        RECT 87.800 115.800 88.200 116.600 ;
        RECT 87.000 115.100 87.300 115.800 ;
        RECT 88.600 115.100 89.000 119.900 ;
        RECT 90.200 117.500 90.600 119.500 ;
        RECT 92.300 119.200 92.700 119.900 ;
        RECT 92.300 118.800 93.000 119.200 ;
        RECT 90.200 115.800 90.500 117.500 ;
        RECT 92.300 116.400 92.700 118.800 ;
        RECT 92.300 116.100 93.100 116.400 ;
        RECT 90.200 115.500 92.100 115.800 ;
        RECT 87.000 114.800 89.000 115.100 ;
        RECT 81.400 113.900 81.900 114.100 ;
        RECT 69.400 113.000 71.400 113.100 ;
        RECT 69.400 111.100 69.800 113.000 ;
        RECT 71.000 111.100 71.400 113.000 ;
        RECT 71.800 111.100 72.200 113.100 ;
        RECT 73.400 112.800 74.300 113.100 ;
        RECT 73.900 111.100 74.300 112.800 ;
        RECT 75.000 112.500 75.300 113.600 ;
        RECT 77.600 113.500 77.900 113.800 ;
        RECT 77.500 113.300 77.900 113.500 ;
        RECT 77.100 113.000 77.900 113.300 ;
        RECT 79.800 113.600 81.900 113.900 ;
        RECT 82.400 113.800 83.400 114.200 ;
        RECT 84.600 114.100 85.000 114.200 ;
        RECT 84.600 113.800 85.400 114.100 ;
        RECT 86.100 113.800 87.400 114.200 ;
        RECT 75.000 111.500 75.400 112.500 ;
        RECT 77.100 111.500 77.500 113.000 ;
        RECT 79.800 112.500 80.100 113.600 ;
        RECT 82.400 113.500 82.700 113.800 ;
        RECT 85.000 113.600 85.400 113.800 ;
        RECT 82.300 113.300 82.700 113.500 ;
        RECT 81.900 113.000 82.700 113.300 ;
        RECT 84.700 113.100 86.500 113.300 ;
        RECT 87.000 113.100 87.300 113.800 ;
        RECT 88.600 113.100 89.000 114.800 ;
        RECT 90.200 114.400 90.600 115.200 ;
        RECT 91.000 114.400 91.400 115.200 ;
        RECT 91.800 114.500 92.100 115.500 ;
        RECT 89.400 113.400 89.800 114.200 ;
        RECT 91.800 114.100 92.500 114.500 ;
        RECT 92.800 114.200 93.100 116.100 ;
        RECT 95.000 115.600 95.400 119.900 ;
        RECT 97.100 117.900 97.700 119.900 ;
        RECT 99.400 117.900 99.800 119.900 ;
        RECT 101.600 118.200 102.000 119.900 ;
        RECT 101.600 117.900 102.600 118.200 ;
        RECT 97.400 117.500 97.800 117.900 ;
        RECT 99.500 117.600 99.800 117.900 ;
        RECT 99.100 117.300 100.900 117.600 ;
        RECT 102.200 117.500 102.600 117.900 ;
        RECT 99.100 117.200 99.500 117.300 ;
        RECT 100.500 117.200 100.900 117.300 ;
        RECT 97.000 116.600 97.700 117.000 ;
        RECT 97.400 116.100 97.700 116.600 ;
        RECT 98.500 116.500 99.600 116.800 ;
        RECT 98.500 116.400 98.900 116.500 ;
        RECT 97.400 115.800 98.600 116.100 ;
        RECT 93.400 114.800 93.800 115.600 ;
        RECT 95.000 115.300 97.100 115.600 ;
        RECT 91.800 113.900 92.300 114.100 ;
        RECT 90.200 113.600 92.300 113.900 ;
        RECT 92.800 113.800 93.800 114.200 ;
        RECT 84.600 113.000 86.600 113.100 ;
        RECT 81.900 112.800 82.600 113.000 ;
        RECT 79.800 111.500 80.200 112.500 ;
        RECT 81.900 111.500 82.300 112.800 ;
        RECT 84.600 111.100 85.000 113.000 ;
        RECT 86.200 111.100 86.600 113.000 ;
        RECT 87.000 111.100 87.400 113.100 ;
        RECT 88.100 112.800 89.000 113.100 ;
        RECT 88.100 111.100 88.500 112.800 ;
        RECT 90.200 112.500 90.500 113.600 ;
        RECT 92.800 113.500 93.100 113.800 ;
        RECT 92.700 113.300 93.100 113.500 ;
        RECT 92.300 113.000 93.100 113.300 ;
        RECT 95.000 113.600 95.400 115.300 ;
        RECT 96.700 115.200 97.100 115.300 ;
        RECT 95.900 114.900 96.300 115.000 ;
        RECT 95.900 114.600 97.800 114.900 ;
        RECT 97.400 114.500 97.800 114.600 ;
        RECT 98.300 114.200 98.600 115.800 ;
        RECT 99.300 115.900 99.600 116.500 ;
        RECT 99.900 116.500 100.300 116.600 ;
        RECT 102.200 116.500 102.600 116.600 ;
        RECT 99.900 116.200 102.600 116.500 ;
        RECT 99.300 115.700 101.700 115.900 ;
        RECT 103.800 115.700 104.200 119.900 ;
        RECT 99.300 115.600 104.200 115.700 ;
        RECT 101.300 115.500 104.200 115.600 ;
        RECT 101.400 115.400 104.200 115.500 ;
        RECT 106.200 115.700 106.600 119.900 ;
        RECT 108.400 118.200 108.800 119.900 ;
        RECT 107.800 117.900 108.800 118.200 ;
        RECT 110.600 117.900 111.000 119.900 ;
        RECT 112.700 117.900 113.300 119.900 ;
        RECT 107.800 117.500 108.200 117.900 ;
        RECT 110.600 117.600 110.900 117.900 ;
        RECT 109.500 117.300 111.300 117.600 ;
        RECT 112.600 117.500 113.000 117.900 ;
        RECT 109.500 117.200 109.900 117.300 ;
        RECT 110.900 117.200 111.300 117.300 ;
        RECT 107.800 116.500 108.200 116.600 ;
        RECT 110.100 116.500 110.500 116.600 ;
        RECT 107.800 116.200 110.500 116.500 ;
        RECT 110.800 116.500 111.900 116.800 ;
        RECT 110.800 115.900 111.100 116.500 ;
        RECT 111.500 116.400 111.900 116.500 ;
        RECT 112.700 116.600 113.400 117.000 ;
        RECT 112.700 116.100 113.000 116.600 ;
        RECT 108.700 115.700 111.100 115.900 ;
        RECT 106.200 115.600 111.100 115.700 ;
        RECT 111.800 115.800 113.000 116.100 ;
        RECT 106.200 115.500 109.100 115.600 ;
        RECT 106.200 115.400 109.000 115.500 ;
        RECT 100.600 115.100 101.000 115.200 ;
        RECT 109.400 115.100 109.800 115.200 ;
        RECT 111.000 115.100 111.400 115.200 ;
        RECT 100.600 114.800 103.100 115.100 ;
        RECT 101.400 114.700 101.800 114.800 ;
        RECT 102.700 114.700 103.100 114.800 ;
        RECT 107.300 114.800 111.400 115.100 ;
        RECT 107.300 114.700 107.700 114.800 ;
        RECT 101.900 114.200 102.300 114.300 ;
        RECT 108.100 114.200 108.500 114.300 ;
        RECT 111.800 114.200 112.100 115.800 ;
        RECT 115.000 115.600 115.400 119.900 ;
        RECT 113.300 115.300 115.400 115.600 ;
        RECT 115.800 115.700 116.200 119.900 ;
        RECT 118.000 118.200 118.400 119.900 ;
        RECT 117.400 117.900 118.400 118.200 ;
        RECT 120.200 117.900 120.600 119.900 ;
        RECT 122.300 117.900 122.900 119.900 ;
        RECT 117.400 117.500 117.800 117.900 ;
        RECT 120.200 117.600 120.500 117.900 ;
        RECT 119.100 117.300 120.900 117.600 ;
        RECT 122.200 117.500 122.600 117.900 ;
        RECT 119.100 117.200 119.500 117.300 ;
        RECT 120.500 117.200 120.900 117.300 ;
        RECT 122.700 117.000 123.400 117.200 ;
        RECT 122.300 116.800 123.400 117.000 ;
        RECT 117.400 116.500 117.800 116.600 ;
        RECT 119.700 116.500 120.100 116.600 ;
        RECT 117.400 116.200 120.100 116.500 ;
        RECT 120.400 116.500 121.500 116.800 ;
        RECT 120.400 115.900 120.700 116.500 ;
        RECT 121.100 116.400 121.500 116.500 ;
        RECT 122.300 116.600 123.000 116.800 ;
        RECT 122.300 116.100 122.600 116.600 ;
        RECT 118.300 115.700 120.700 115.900 ;
        RECT 115.800 115.600 120.700 115.700 ;
        RECT 121.400 115.800 122.600 116.100 ;
        RECT 115.800 115.500 118.700 115.600 ;
        RECT 115.800 115.400 118.600 115.500 ;
        RECT 113.300 115.200 113.700 115.300 ;
        RECT 114.100 114.900 114.500 115.000 ;
        RECT 112.600 114.600 114.500 114.900 ;
        RECT 112.600 114.500 113.000 114.600 ;
        RECT 98.300 114.100 103.800 114.200 ;
        RECT 106.600 114.100 112.100 114.200 ;
        RECT 98.300 113.900 112.100 114.100 ;
        RECT 98.500 113.800 98.900 113.900 ;
        RECT 95.000 113.300 96.900 113.600 ;
        RECT 90.200 111.500 90.600 112.500 ;
        RECT 92.300 111.500 92.700 113.000 ;
        RECT 95.000 111.100 95.400 113.300 ;
        RECT 96.500 113.200 96.900 113.300 ;
        RECT 101.400 112.800 101.700 113.900 ;
        RECT 103.000 113.800 107.400 113.900 ;
        RECT 100.500 112.700 100.900 112.800 ;
        RECT 97.400 112.100 97.800 112.500 ;
        RECT 99.500 112.400 100.900 112.700 ;
        RECT 101.400 112.400 101.800 112.800 ;
        RECT 99.500 112.100 99.800 112.400 ;
        RECT 102.200 112.100 102.600 112.500 ;
        RECT 97.100 111.800 97.800 112.100 ;
        RECT 97.100 111.100 97.700 111.800 ;
        RECT 99.400 111.100 99.800 112.100 ;
        RECT 101.600 111.800 102.600 112.100 ;
        RECT 101.600 111.100 102.000 111.800 ;
        RECT 103.800 111.100 104.200 113.500 ;
        RECT 106.200 111.100 106.600 113.500 ;
        RECT 108.700 112.800 109.000 113.900 ;
        RECT 109.400 113.800 109.800 113.900 ;
        RECT 111.500 113.800 111.900 113.900 ;
        RECT 115.000 113.600 115.400 115.300 ;
        RECT 121.400 115.200 121.700 115.800 ;
        RECT 124.600 115.600 125.000 119.900 ;
        RECT 126.700 116.200 127.100 119.900 ;
        RECT 127.400 116.800 127.800 117.200 ;
        RECT 127.500 116.200 127.800 116.800 ;
        RECT 129.900 116.200 130.300 119.900 ;
        RECT 130.600 116.800 131.000 117.200 ;
        RECT 130.700 116.200 131.000 116.800 ;
        RECT 126.700 115.900 127.200 116.200 ;
        RECT 127.500 115.900 128.200 116.200 ;
        RECT 129.900 115.900 130.400 116.200 ;
        RECT 130.700 115.900 131.400 116.200 ;
        RECT 122.900 115.300 125.000 115.600 ;
        RECT 122.900 115.200 123.300 115.300 ;
        RECT 119.000 115.100 119.400 115.200 ;
        RECT 116.900 114.800 119.400 115.100 ;
        RECT 121.400 114.800 121.800 115.200 ;
        RECT 123.700 114.900 124.100 115.000 ;
        RECT 116.900 114.700 117.300 114.800 ;
        RECT 117.700 114.200 118.100 114.300 ;
        RECT 121.400 114.200 121.700 114.800 ;
        RECT 122.200 114.600 124.100 114.900 ;
        RECT 122.200 114.500 122.600 114.600 ;
        RECT 116.200 113.900 121.700 114.200 ;
        RECT 116.200 113.800 117.000 113.900 ;
        RECT 113.500 113.300 115.400 113.600 ;
        RECT 113.500 113.200 113.900 113.300 ;
        RECT 107.800 112.100 108.200 112.500 ;
        RECT 108.600 112.400 109.000 112.800 ;
        RECT 109.500 112.700 109.900 112.800 ;
        RECT 109.500 112.400 110.900 112.700 ;
        RECT 110.600 112.100 110.900 112.400 ;
        RECT 112.600 112.100 113.000 112.500 ;
        RECT 107.800 111.800 108.800 112.100 ;
        RECT 108.400 111.100 108.800 111.800 ;
        RECT 110.600 111.100 111.000 112.100 ;
        RECT 112.600 111.800 113.300 112.100 ;
        RECT 112.700 111.100 113.300 111.800 ;
        RECT 115.000 111.100 115.400 113.300 ;
        RECT 115.800 111.100 116.200 113.500 ;
        RECT 118.300 112.800 118.600 113.900 ;
        RECT 121.100 113.800 121.500 113.900 ;
        RECT 124.600 113.600 125.000 115.300 ;
        RECT 126.200 114.400 126.600 115.200 ;
        RECT 126.900 115.100 127.200 115.900 ;
        RECT 127.800 115.800 128.200 115.900 ;
        RECT 128.600 115.100 129.000 115.200 ;
        RECT 126.900 114.800 129.000 115.100 ;
        RECT 126.900 114.200 127.200 114.800 ;
        RECT 129.400 114.400 129.800 115.200 ;
        RECT 130.100 114.200 130.400 115.900 ;
        RECT 131.000 115.800 131.400 115.900 ;
        RECT 131.800 115.800 132.200 116.600 ;
        RECT 131.000 115.100 131.300 115.800 ;
        RECT 132.600 115.100 133.000 119.900 ;
        RECT 134.200 115.700 134.600 119.900 ;
        RECT 136.400 118.200 136.800 119.900 ;
        RECT 135.800 117.900 136.800 118.200 ;
        RECT 138.600 117.900 139.000 119.900 ;
        RECT 140.700 117.900 141.300 119.900 ;
        RECT 135.800 117.500 136.200 117.900 ;
        RECT 138.600 117.600 138.900 117.900 ;
        RECT 137.500 117.300 139.300 117.600 ;
        RECT 140.600 117.500 141.000 117.900 ;
        RECT 137.500 117.200 137.900 117.300 ;
        RECT 138.900 117.200 139.300 117.300 ;
        RECT 135.800 116.500 136.200 116.600 ;
        RECT 138.100 116.500 138.500 116.600 ;
        RECT 135.800 116.200 138.500 116.500 ;
        RECT 138.800 116.500 139.900 116.800 ;
        RECT 138.800 115.900 139.100 116.500 ;
        RECT 139.500 116.400 139.900 116.500 ;
        RECT 140.700 116.600 141.400 117.000 ;
        RECT 140.700 116.100 141.000 116.600 ;
        RECT 136.700 115.700 139.100 115.900 ;
        RECT 134.200 115.600 139.100 115.700 ;
        RECT 139.800 115.800 141.000 116.100 ;
        RECT 134.200 115.500 137.100 115.600 ;
        RECT 134.200 115.400 137.000 115.500 ;
        RECT 137.400 115.100 137.800 115.200 ;
        RECT 131.000 114.800 133.000 115.100 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 125.400 113.800 126.200 114.100 ;
        RECT 126.900 113.800 128.200 114.200 ;
        RECT 128.600 114.100 129.000 114.200 ;
        RECT 130.100 114.100 131.400 114.200 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 128.600 113.800 129.400 114.100 ;
        RECT 130.100 113.800 132.200 114.100 ;
        RECT 125.800 113.600 126.200 113.800 ;
        RECT 123.100 113.300 125.000 113.600 ;
        RECT 123.100 113.200 123.500 113.300 ;
        RECT 117.400 112.100 117.800 112.500 ;
        RECT 118.200 112.400 118.600 112.800 ;
        RECT 119.100 112.700 119.500 112.800 ;
        RECT 119.100 112.400 120.500 112.700 ;
        RECT 120.200 112.100 120.500 112.400 ;
        RECT 122.200 112.100 122.600 112.500 ;
        RECT 117.400 111.800 118.400 112.100 ;
        RECT 118.000 111.100 118.400 111.800 ;
        RECT 120.200 111.100 120.600 112.100 ;
        RECT 122.200 111.800 122.900 112.100 ;
        RECT 122.300 111.100 122.900 111.800 ;
        RECT 124.600 111.100 125.000 113.300 ;
        RECT 125.500 113.100 127.300 113.300 ;
        RECT 127.800 113.100 128.100 113.800 ;
        RECT 129.000 113.600 129.400 113.800 ;
        RECT 128.700 113.100 130.500 113.300 ;
        RECT 131.000 113.100 131.300 113.800 ;
        RECT 132.600 113.100 133.000 114.800 ;
        RECT 135.300 114.800 137.800 115.100 ;
        RECT 135.300 114.700 135.700 114.800 ;
        RECT 136.600 114.700 137.000 114.800 ;
        RECT 136.100 114.200 136.500 114.300 ;
        RECT 139.800 114.200 140.100 115.800 ;
        RECT 143.000 115.600 143.400 119.900 ;
        RECT 145.100 116.300 145.500 119.900 ;
        RECT 147.500 116.300 147.900 119.900 ;
        RECT 148.900 119.200 149.300 119.900 ;
        RECT 148.600 118.800 149.300 119.200 ;
        RECT 144.600 115.900 145.500 116.300 ;
        RECT 147.000 115.900 147.900 116.300 ;
        RECT 148.900 116.300 149.300 118.800 ;
        RECT 151.000 117.500 151.400 119.500 ;
        RECT 153.100 119.200 153.500 119.900 ;
        RECT 152.600 118.800 153.500 119.200 ;
        RECT 148.900 115.900 149.800 116.300 ;
        RECT 141.300 115.300 143.400 115.600 ;
        RECT 141.300 115.200 141.700 115.300 ;
        RECT 142.100 114.900 142.500 115.000 ;
        RECT 140.600 114.600 142.500 114.900 ;
        RECT 140.600 114.500 141.000 114.600 ;
        RECT 133.400 113.400 133.800 114.200 ;
        RECT 134.600 113.900 140.100 114.200 ;
        RECT 134.600 113.800 135.400 113.900 ;
        RECT 125.400 113.000 127.400 113.100 ;
        RECT 125.400 111.100 125.800 113.000 ;
        RECT 127.000 111.100 127.400 113.000 ;
        RECT 127.800 111.100 128.200 113.100 ;
        RECT 128.600 113.000 130.600 113.100 ;
        RECT 128.600 111.100 129.000 113.000 ;
        RECT 130.200 111.100 130.600 113.000 ;
        RECT 131.000 111.100 131.400 113.100 ;
        RECT 132.100 112.800 133.000 113.100 ;
        RECT 132.100 111.100 132.500 112.800 ;
        RECT 134.200 111.100 134.600 113.500 ;
        RECT 136.700 112.800 137.000 113.900 ;
        RECT 138.200 113.800 138.600 113.900 ;
        RECT 139.500 113.800 139.900 113.900 ;
        RECT 143.000 113.600 143.400 115.300 ;
        RECT 144.700 114.200 145.000 115.900 ;
        RECT 147.000 115.800 147.400 115.900 ;
        RECT 145.400 114.800 145.800 115.600 ;
        RECT 147.100 114.200 147.400 115.800 ;
        RECT 147.800 115.100 148.200 115.600 ;
        RECT 148.600 115.100 149.000 115.600 ;
        RECT 147.800 114.800 149.000 115.100 ;
        RECT 144.600 113.800 145.000 114.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 141.500 113.300 143.400 113.600 ;
        RECT 141.500 113.200 141.900 113.300 ;
        RECT 135.800 112.100 136.200 112.500 ;
        RECT 136.600 112.400 137.000 112.800 ;
        RECT 137.500 112.700 137.900 112.800 ;
        RECT 137.500 112.400 138.900 112.700 ;
        RECT 138.600 112.100 138.900 112.400 ;
        RECT 140.600 112.100 141.000 112.500 ;
        RECT 135.800 111.800 136.800 112.100 ;
        RECT 136.400 111.100 136.800 111.800 ;
        RECT 138.600 111.100 139.000 112.100 ;
        RECT 140.600 111.800 141.300 112.100 ;
        RECT 140.700 111.100 141.300 111.800 ;
        RECT 143.000 111.100 143.400 113.300 ;
        RECT 143.800 112.400 144.200 113.200 ;
        RECT 144.700 112.200 145.000 113.800 ;
        RECT 146.200 112.400 146.600 113.200 ;
        RECT 144.600 111.100 145.000 112.200 ;
        RECT 147.100 112.100 147.400 113.800 ;
        RECT 147.000 111.100 147.400 112.100 ;
        RECT 149.400 114.200 149.700 115.900 ;
        RECT 151.000 115.800 151.300 117.500 ;
        RECT 153.100 116.400 153.500 118.800 ;
        RECT 153.100 116.100 153.900 116.400 ;
        RECT 151.000 115.500 152.900 115.800 ;
        RECT 151.000 114.400 151.400 115.200 ;
        RECT 151.800 114.400 152.200 115.200 ;
        RECT 152.600 114.500 152.900 115.500 ;
        RECT 149.400 113.800 149.800 114.200 ;
        RECT 152.600 114.100 153.300 114.500 ;
        RECT 153.600 114.200 153.900 116.100 ;
        RECT 154.200 115.100 154.600 115.600 ;
        RECT 156.600 115.100 157.000 119.900 ;
        RECT 160.200 116.800 160.600 117.200 ;
        RECT 157.400 115.800 157.800 116.600 ;
        RECT 160.200 116.200 160.500 116.800 ;
        RECT 160.900 116.200 161.300 119.900 ;
        RECT 159.800 115.900 160.500 116.200 ;
        RECT 160.800 115.900 161.300 116.200 ;
        RECT 159.800 115.800 160.200 115.900 ;
        RECT 159.800 115.100 160.100 115.800 ;
        RECT 154.200 114.800 155.300 115.100 ;
        RECT 152.600 113.900 153.100 114.100 ;
        RECT 149.400 112.100 149.700 113.800 ;
        RECT 151.000 113.600 153.100 113.900 ;
        RECT 153.600 113.800 154.600 114.200 ;
        RECT 155.000 114.100 155.300 114.800 ;
        RECT 156.600 114.800 160.100 115.100 ;
        RECT 155.800 114.100 156.200 114.200 ;
        RECT 155.000 113.800 156.200 114.100 ;
        RECT 150.200 112.400 150.600 113.200 ;
        RECT 151.000 112.500 151.300 113.600 ;
        RECT 153.600 113.500 153.900 113.800 ;
        RECT 153.500 113.300 153.900 113.500 ;
        RECT 155.800 113.400 156.200 113.800 ;
        RECT 153.100 113.000 153.900 113.300 ;
        RECT 156.600 113.100 157.000 114.800 ;
        RECT 160.800 114.200 161.100 115.900 ;
        RECT 163.000 115.600 163.400 119.900 ;
        RECT 165.100 117.900 165.700 119.900 ;
        RECT 167.400 117.900 167.800 119.900 ;
        RECT 169.600 118.200 170.000 119.900 ;
        RECT 169.600 117.900 170.600 118.200 ;
        RECT 165.400 117.500 165.800 117.900 ;
        RECT 167.500 117.600 167.800 117.900 ;
        RECT 167.100 117.300 168.900 117.600 ;
        RECT 170.200 117.500 170.600 117.900 ;
        RECT 167.100 117.200 167.500 117.300 ;
        RECT 168.500 117.200 168.900 117.300 ;
        RECT 165.000 116.600 165.700 117.000 ;
        RECT 165.400 116.100 165.700 116.600 ;
        RECT 166.500 116.500 167.600 116.800 ;
        RECT 166.500 116.400 166.900 116.500 ;
        RECT 165.400 115.800 166.600 116.100 ;
        RECT 163.000 115.300 165.100 115.600 ;
        RECT 161.400 114.400 161.800 115.200 ;
        RECT 159.800 113.800 161.100 114.200 ;
        RECT 162.200 114.100 162.600 114.200 ;
        RECT 161.800 113.800 162.600 114.100 ;
        RECT 159.900 113.100 160.200 113.800 ;
        RECT 161.800 113.600 162.200 113.800 ;
        RECT 163.000 113.600 163.400 115.300 ;
        RECT 164.700 115.200 165.100 115.300 ;
        RECT 163.900 114.900 164.300 115.000 ;
        RECT 163.900 114.600 165.800 114.900 ;
        RECT 165.400 114.500 165.800 114.600 ;
        RECT 166.300 114.200 166.600 115.800 ;
        RECT 167.300 115.900 167.600 116.500 ;
        RECT 167.900 116.500 168.300 116.600 ;
        RECT 170.200 116.500 170.600 116.600 ;
        RECT 167.900 116.200 170.600 116.500 ;
        RECT 167.300 115.700 169.700 115.900 ;
        RECT 171.800 115.700 172.200 119.900 ;
        RECT 167.300 115.600 172.200 115.700 ;
        RECT 173.400 115.600 173.800 119.900 ;
        RECT 175.000 115.600 175.400 119.900 ;
        RECT 176.600 115.600 177.000 119.900 ;
        RECT 178.200 115.600 178.600 119.900 ;
        RECT 169.300 115.500 172.200 115.600 ;
        RECT 169.400 115.400 172.200 115.500 ;
        RECT 172.600 115.200 173.800 115.600 ;
        RECT 174.300 115.200 175.400 115.600 ;
        RECT 175.900 115.200 177.000 115.600 ;
        RECT 177.700 115.200 178.600 115.600 ;
        RECT 180.600 115.600 181.000 119.900 ;
        RECT 182.200 115.600 182.600 119.900 ;
        RECT 183.800 115.600 184.200 119.900 ;
        RECT 185.400 115.600 185.800 119.900 ;
        RECT 180.600 115.200 181.500 115.600 ;
        RECT 182.200 115.200 183.300 115.600 ;
        RECT 183.800 115.200 184.900 115.600 ;
        RECT 185.400 115.200 186.600 115.600 ;
        RECT 167.800 115.100 168.200 115.200 ;
        RECT 168.600 115.100 169.000 115.200 ;
        RECT 167.800 114.800 171.100 115.100 ;
        RECT 170.700 114.700 171.100 114.800 ;
        RECT 169.900 114.200 170.300 114.300 ;
        RECT 166.300 113.900 171.800 114.200 ;
        RECT 166.500 113.800 166.900 113.900 ;
        RECT 163.000 113.300 164.900 113.600 ;
        RECT 160.700 113.100 162.500 113.300 ;
        RECT 149.400 111.100 149.800 112.100 ;
        RECT 151.000 111.500 151.400 112.500 ;
        RECT 153.100 111.500 153.500 113.000 ;
        RECT 156.600 112.800 157.500 113.100 ;
        RECT 157.100 111.100 157.500 112.800 ;
        RECT 159.800 111.100 160.200 113.100 ;
        RECT 160.600 113.000 162.600 113.100 ;
        RECT 160.600 111.100 161.000 113.000 ;
        RECT 162.200 111.100 162.600 113.000 ;
        RECT 163.000 111.100 163.400 113.300 ;
        RECT 164.500 113.200 164.900 113.300 ;
        RECT 169.400 112.800 169.700 113.900 ;
        RECT 171.000 113.800 171.800 113.900 ;
        RECT 172.600 113.800 173.000 115.200 ;
        RECT 174.300 114.500 174.700 115.200 ;
        RECT 175.900 114.500 176.300 115.200 ;
        RECT 177.700 114.500 178.100 115.200 ;
        RECT 181.100 114.500 181.500 115.200 ;
        RECT 182.900 114.500 183.300 115.200 ;
        RECT 184.500 114.500 184.900 115.200 ;
        RECT 173.400 114.100 174.700 114.500 ;
        RECT 175.100 114.100 176.300 114.500 ;
        RECT 176.800 114.100 178.100 114.500 ;
        RECT 178.500 114.100 179.400 114.500 ;
        RECT 179.800 114.100 180.700 114.500 ;
        RECT 181.100 114.100 182.400 114.500 ;
        RECT 182.900 114.100 184.100 114.500 ;
        RECT 184.500 114.100 185.800 114.500 ;
        RECT 174.300 113.800 174.700 114.100 ;
        RECT 175.900 113.800 176.300 114.100 ;
        RECT 177.700 113.800 178.100 114.100 ;
        RECT 179.000 113.800 180.200 114.100 ;
        RECT 181.100 113.800 181.500 114.100 ;
        RECT 182.900 113.800 183.300 114.100 ;
        RECT 184.500 113.800 184.900 114.100 ;
        RECT 186.200 113.800 186.600 115.200 ;
        RECT 168.500 112.700 168.900 112.800 ;
        RECT 165.400 112.100 165.800 112.500 ;
        RECT 167.500 112.400 168.900 112.700 ;
        RECT 169.400 112.400 169.800 112.800 ;
        RECT 167.500 112.100 167.800 112.400 ;
        RECT 170.200 112.100 170.600 112.500 ;
        RECT 165.100 111.800 165.800 112.100 ;
        RECT 165.100 111.100 165.700 111.800 ;
        RECT 167.400 111.100 167.800 112.100 ;
        RECT 169.600 111.800 170.600 112.100 ;
        RECT 169.600 111.100 170.000 111.800 ;
        RECT 171.800 111.100 172.200 113.500 ;
        RECT 172.600 113.400 173.800 113.800 ;
        RECT 174.300 113.400 175.400 113.800 ;
        RECT 175.900 113.400 177.000 113.800 ;
        RECT 177.700 113.400 178.600 113.800 ;
        RECT 173.400 111.100 173.800 113.400 ;
        RECT 175.000 111.100 175.400 113.400 ;
        RECT 176.600 111.100 177.000 113.400 ;
        RECT 178.200 111.100 178.600 113.400 ;
        RECT 180.600 113.400 181.500 113.800 ;
        RECT 182.200 113.400 183.300 113.800 ;
        RECT 183.800 113.400 184.900 113.800 ;
        RECT 185.400 113.400 186.600 113.800 ;
        RECT 187.000 113.400 187.400 114.200 ;
        RECT 180.600 111.100 181.000 113.400 ;
        RECT 182.200 111.100 182.600 113.400 ;
        RECT 183.800 111.100 184.200 113.400 ;
        RECT 185.400 111.100 185.800 113.400 ;
        RECT 187.800 111.100 188.200 119.900 ;
        RECT 188.600 115.600 189.000 119.900 ;
        RECT 190.700 117.900 191.300 119.900 ;
        RECT 193.000 117.900 193.400 119.900 ;
        RECT 195.200 118.200 195.600 119.900 ;
        RECT 195.200 117.900 196.200 118.200 ;
        RECT 191.000 117.500 191.400 117.900 ;
        RECT 193.100 117.600 193.400 117.900 ;
        RECT 192.700 117.300 194.500 117.600 ;
        RECT 195.800 117.500 196.200 117.900 ;
        RECT 192.700 117.200 193.100 117.300 ;
        RECT 194.100 117.200 194.500 117.300 ;
        RECT 190.600 116.600 191.300 117.000 ;
        RECT 191.000 116.100 191.300 116.600 ;
        RECT 192.100 116.500 193.200 116.800 ;
        RECT 192.100 116.400 192.500 116.500 ;
        RECT 191.000 115.800 192.200 116.100 ;
        RECT 188.600 115.300 190.700 115.600 ;
        RECT 188.600 113.600 189.000 115.300 ;
        RECT 190.300 115.200 190.700 115.300 ;
        RECT 191.900 115.200 192.200 115.800 ;
        RECT 192.900 115.900 193.200 116.500 ;
        RECT 193.500 116.500 193.900 116.600 ;
        RECT 195.800 116.500 196.200 116.600 ;
        RECT 193.500 116.200 196.200 116.500 ;
        RECT 192.900 115.700 195.300 115.900 ;
        RECT 197.400 115.700 197.800 119.900 ;
        RECT 199.000 116.400 199.400 119.900 ;
        RECT 192.900 115.600 197.800 115.700 ;
        RECT 194.900 115.500 197.800 115.600 ;
        RECT 195.000 115.400 197.800 115.500 ;
        RECT 198.900 115.900 199.400 116.400 ;
        RECT 200.600 116.200 201.000 119.900 ;
        RECT 202.200 116.400 202.600 119.900 ;
        RECT 199.700 115.900 201.000 116.200 ;
        RECT 202.100 115.900 202.600 116.400 ;
        RECT 203.800 116.200 204.200 119.900 ;
        RECT 206.500 119.200 206.900 119.900 ;
        RECT 206.200 118.800 206.900 119.200 ;
        RECT 206.500 116.400 206.900 118.800 ;
        RECT 208.600 117.500 209.000 119.500 ;
        RECT 202.900 115.900 204.200 116.200 ;
        RECT 206.100 116.100 206.900 116.400 ;
        RECT 189.500 114.900 189.900 115.000 ;
        RECT 189.500 114.600 191.400 114.900 ;
        RECT 191.800 114.800 192.200 115.200 ;
        RECT 194.200 115.100 194.600 115.200 ;
        RECT 194.200 114.800 196.700 115.100 ;
        RECT 191.000 114.500 191.400 114.600 ;
        RECT 191.900 114.200 192.200 114.800 ;
        RECT 195.000 114.700 195.400 114.800 ;
        RECT 196.300 114.700 196.700 114.800 ;
        RECT 195.500 114.200 195.900 114.300 ;
        RECT 198.900 114.200 199.200 115.900 ;
        RECT 199.700 114.900 200.000 115.900 ;
        RECT 199.500 114.500 200.000 114.900 ;
        RECT 191.900 113.900 197.400 114.200 ;
        RECT 192.100 113.800 192.500 113.900 ;
        RECT 188.600 113.300 190.500 113.600 ;
        RECT 188.600 111.100 189.000 113.300 ;
        RECT 190.100 113.200 190.500 113.300 ;
        RECT 195.000 112.800 195.300 113.900 ;
        RECT 196.600 113.800 197.400 113.900 ;
        RECT 198.900 113.800 199.400 114.200 ;
        RECT 194.100 112.700 194.500 112.800 ;
        RECT 191.000 112.100 191.400 112.500 ;
        RECT 193.100 112.400 194.500 112.700 ;
        RECT 195.000 112.400 195.400 112.800 ;
        RECT 193.100 112.100 193.400 112.400 ;
        RECT 195.800 112.100 196.200 112.500 ;
        RECT 190.700 111.800 191.400 112.100 ;
        RECT 190.700 111.100 191.300 111.800 ;
        RECT 193.000 111.100 193.400 112.100 ;
        RECT 195.200 111.800 196.200 112.100 ;
        RECT 195.200 111.100 195.600 111.800 ;
        RECT 197.400 111.100 197.800 113.500 ;
        RECT 198.900 113.100 199.200 113.800 ;
        RECT 199.700 113.700 200.000 114.500 ;
        RECT 200.500 115.100 201.000 115.200 ;
        RECT 201.400 115.100 201.800 115.200 ;
        RECT 200.500 114.800 201.800 115.100 ;
        RECT 200.500 114.400 200.900 114.800 ;
        RECT 202.100 114.200 202.400 115.900 ;
        RECT 202.900 114.900 203.200 115.900 ;
        RECT 202.700 114.500 203.200 114.900 ;
        RECT 202.100 113.800 202.600 114.200 ;
        RECT 199.700 113.400 201.000 113.700 ;
        RECT 198.900 112.800 199.400 113.100 ;
        RECT 199.000 111.100 199.400 112.800 ;
        RECT 200.600 111.100 201.000 113.400 ;
        RECT 202.100 113.100 202.400 113.800 ;
        RECT 202.900 113.700 203.200 114.500 ;
        RECT 203.700 114.800 204.200 115.200 ;
        RECT 205.400 114.800 205.800 115.600 ;
        RECT 203.700 114.400 204.100 114.800 ;
        RECT 206.100 114.200 206.400 116.100 ;
        RECT 208.700 115.800 209.000 117.500 ;
        RECT 207.100 115.500 209.000 115.800 ;
        RECT 207.100 114.500 207.400 115.500 ;
        RECT 205.400 113.800 206.400 114.200 ;
        RECT 206.700 114.100 207.400 114.500 ;
        RECT 207.800 114.400 208.200 115.200 ;
        RECT 208.600 114.400 209.000 115.200 ;
        RECT 211.000 115.100 211.400 115.200 ;
        RECT 211.800 115.100 212.200 119.900 ;
        RECT 212.600 115.800 213.000 116.600 ;
        RECT 214.700 116.300 215.100 119.900 ;
        RECT 214.200 115.900 215.100 116.300 ;
        RECT 215.800 115.900 216.200 119.900 ;
        RECT 216.600 116.200 217.000 119.900 ;
        RECT 218.200 116.200 218.600 119.900 ;
        RECT 216.600 115.900 218.600 116.200 ;
        RECT 211.000 114.800 212.200 115.100 ;
        RECT 202.900 113.400 204.200 113.700 ;
        RECT 202.100 112.800 202.600 113.100 ;
        RECT 202.200 111.100 202.600 112.800 ;
        RECT 203.800 111.100 204.200 113.400 ;
        RECT 206.100 113.500 206.400 113.800 ;
        RECT 206.900 113.900 207.400 114.100 ;
        RECT 210.200 114.100 210.600 114.200 ;
        RECT 211.000 114.100 211.400 114.200 ;
        RECT 206.900 113.600 209.000 113.900 ;
        RECT 210.200 113.800 211.400 114.100 ;
        RECT 206.100 113.300 206.500 113.500 ;
        RECT 206.100 113.000 206.900 113.300 ;
        RECT 206.500 111.500 206.900 113.000 ;
        RECT 208.700 112.500 209.000 113.600 ;
        RECT 211.000 113.400 211.400 113.800 ;
        RECT 211.800 113.100 212.200 114.800 ;
        RECT 214.300 114.200 214.600 115.900 ;
        RECT 215.000 114.800 215.400 115.600 ;
        RECT 215.900 115.200 216.200 115.900 ;
        RECT 219.000 115.700 219.400 119.900 ;
        RECT 221.200 118.200 221.600 119.900 ;
        RECT 220.600 117.900 221.600 118.200 ;
        RECT 223.400 117.900 223.800 119.900 ;
        RECT 225.500 117.900 226.100 119.900 ;
        RECT 220.600 117.500 221.000 117.900 ;
        RECT 223.400 117.600 223.700 117.900 ;
        RECT 222.300 117.300 224.100 117.600 ;
        RECT 225.400 117.500 225.800 117.900 ;
        RECT 222.300 117.200 222.700 117.300 ;
        RECT 223.700 117.200 224.100 117.300 ;
        RECT 227.800 117.100 228.200 119.900 ;
        RECT 228.600 117.100 229.000 117.200 ;
        RECT 220.600 116.500 221.000 116.600 ;
        RECT 222.900 116.500 223.300 116.600 ;
        RECT 220.600 116.200 223.300 116.500 ;
        RECT 223.600 116.500 224.700 116.800 ;
        RECT 223.600 115.900 223.900 116.500 ;
        RECT 224.300 116.400 224.700 116.500 ;
        RECT 225.500 116.600 226.200 117.000 ;
        RECT 227.800 116.800 229.000 117.100 ;
        RECT 225.500 116.100 225.800 116.600 ;
        RECT 221.500 115.700 223.900 115.900 ;
        RECT 219.000 115.600 223.900 115.700 ;
        RECT 224.600 115.800 225.800 116.100 ;
        RECT 219.000 115.500 221.900 115.600 ;
        RECT 219.000 115.400 221.800 115.500 ;
        RECT 217.800 115.200 218.200 115.400 ;
        RECT 215.800 114.900 217.000 115.200 ;
        RECT 217.800 114.900 218.600 115.200 ;
        RECT 222.200 115.100 222.600 115.200 ;
        RECT 215.800 114.800 216.200 114.900 ;
        RECT 214.200 113.800 214.600 114.200 ;
        RECT 211.800 112.800 212.700 113.100 ;
        RECT 208.600 111.500 209.000 112.500 ;
        RECT 212.300 111.100 212.700 112.800 ;
        RECT 213.400 112.400 213.800 113.200 ;
        RECT 214.300 113.100 214.600 113.800 ;
        RECT 215.800 113.100 216.200 113.200 ;
        RECT 216.700 113.100 217.000 114.900 ;
        RECT 218.200 114.800 218.600 114.900 ;
        RECT 220.100 114.800 222.600 115.100 ;
        RECT 220.100 114.700 220.500 114.800 ;
        RECT 217.400 113.800 217.800 114.600 ;
        RECT 220.900 114.200 221.300 114.300 ;
        RECT 224.600 114.200 224.900 115.800 ;
        RECT 227.800 115.600 228.200 116.800 ;
        RECT 226.100 115.300 228.200 115.600 ;
        RECT 226.100 115.200 226.500 115.300 ;
        RECT 226.900 114.900 227.300 115.000 ;
        RECT 225.400 114.600 227.300 114.900 ;
        RECT 225.400 114.500 225.800 114.600 ;
        RECT 219.400 113.900 224.900 114.200 ;
        RECT 219.400 113.800 220.200 113.900 ;
        RECT 214.200 112.800 216.200 113.100 ;
        RECT 214.300 112.100 214.600 112.800 ;
        RECT 215.900 112.400 216.300 112.800 ;
        RECT 214.200 111.100 214.600 112.100 ;
        RECT 216.600 111.100 217.000 113.100 ;
        RECT 219.000 111.100 219.400 113.500 ;
        RECT 221.500 113.200 221.800 113.900 ;
        RECT 224.300 113.800 224.700 113.900 ;
        RECT 227.800 113.600 228.200 115.300 ;
        RECT 229.400 115.100 229.800 119.900 ;
        RECT 231.400 116.800 231.800 117.200 ;
        RECT 230.200 115.800 230.600 116.600 ;
        RECT 231.400 116.200 231.700 116.800 ;
        RECT 232.100 116.200 232.500 119.900 ;
        RECT 231.000 115.900 231.700 116.200 ;
        RECT 232.000 115.900 232.500 116.200 ;
        RECT 234.200 116.200 234.600 119.900 ;
        RECT 235.800 116.200 236.200 119.900 ;
        RECT 234.200 115.900 236.200 116.200 ;
        RECT 236.600 115.900 237.000 119.900 ;
        RECT 237.400 116.200 237.800 119.900 ;
        RECT 239.000 116.400 239.400 119.900 ;
        RECT 237.400 115.900 238.700 116.200 ;
        RECT 239.000 115.900 239.500 116.400 ;
        RECT 241.900 116.300 242.300 119.900 ;
        RECT 241.400 115.900 242.300 116.300 ;
        RECT 243.000 116.200 243.400 119.900 ;
        RECT 244.600 116.200 245.000 119.900 ;
        RECT 243.000 115.900 245.000 116.200 ;
        RECT 231.000 115.800 231.400 115.900 ;
        RECT 231.000 115.100 231.300 115.800 ;
        RECT 229.400 114.800 231.300 115.100 ;
        RECT 226.300 113.300 228.200 113.600 ;
        RECT 228.600 113.400 229.000 114.200 ;
        RECT 226.300 113.200 226.700 113.300 ;
        RECT 220.600 112.100 221.000 112.500 ;
        RECT 221.400 112.400 221.800 113.200 ;
        RECT 222.300 112.700 222.700 112.800 ;
        RECT 222.300 112.400 223.700 112.700 ;
        RECT 223.400 112.100 223.700 112.400 ;
        RECT 225.400 112.100 225.800 112.500 ;
        RECT 220.600 111.800 221.600 112.100 ;
        RECT 221.200 111.100 221.600 111.800 ;
        RECT 223.400 111.100 223.800 112.100 ;
        RECT 225.400 111.800 226.100 112.100 ;
        RECT 225.500 111.100 226.100 111.800 ;
        RECT 227.800 111.100 228.200 113.300 ;
        RECT 229.400 113.100 229.800 114.800 ;
        RECT 232.000 114.200 232.300 115.900 ;
        RECT 236.600 115.200 236.900 115.900 ;
        RECT 232.600 114.400 233.000 115.200 ;
        RECT 235.800 114.900 237.000 115.200 ;
        RECT 230.200 114.100 230.600 114.200 ;
        RECT 231.000 114.100 232.300 114.200 ;
        RECT 233.400 114.100 233.800 114.200 ;
        RECT 230.200 113.800 232.300 114.100 ;
        RECT 233.000 113.800 233.800 114.100 ;
        RECT 235.000 113.800 235.400 114.600 ;
        RECT 231.100 113.100 231.400 113.800 ;
        RECT 233.000 113.600 233.400 113.800 ;
        RECT 231.900 113.100 233.700 113.300 ;
        RECT 235.800 113.200 236.100 114.900 ;
        RECT 236.600 114.800 237.000 114.900 ;
        RECT 237.400 114.800 237.900 115.200 ;
        RECT 237.500 114.400 237.900 114.800 ;
        RECT 238.400 114.900 238.700 115.900 ;
        RECT 238.400 114.500 238.900 114.900 ;
        RECT 238.400 113.700 238.700 114.500 ;
        RECT 239.200 114.200 239.500 115.900 ;
        RECT 241.500 114.200 241.800 115.900 ;
        RECT 245.400 115.800 245.800 119.900 ;
        RECT 243.400 115.200 243.800 115.400 ;
        RECT 245.400 115.200 245.700 115.800 ;
        RECT 246.200 115.600 246.600 119.900 ;
        RECT 248.300 117.900 248.900 119.900 ;
        RECT 250.600 117.900 251.000 119.900 ;
        RECT 252.800 118.200 253.200 119.900 ;
        RECT 252.800 117.900 253.800 118.200 ;
        RECT 248.600 117.500 249.000 117.900 ;
        RECT 250.700 117.600 251.000 117.900 ;
        RECT 250.300 117.300 252.100 117.600 ;
        RECT 253.400 117.500 253.800 117.900 ;
        RECT 250.300 117.200 250.700 117.300 ;
        RECT 251.700 117.200 252.100 117.300 ;
        RECT 248.200 116.600 248.900 117.000 ;
        RECT 248.600 116.100 248.900 116.600 ;
        RECT 249.700 116.500 250.800 116.800 ;
        RECT 249.700 116.400 250.100 116.500 ;
        RECT 248.600 115.800 249.800 116.100 ;
        RECT 246.200 115.300 248.300 115.600 ;
        RECT 243.000 114.900 243.800 115.200 ;
        RECT 244.600 114.900 245.800 115.200 ;
        RECT 243.000 114.800 243.400 114.900 ;
        RECT 239.000 113.800 239.500 114.200 ;
        RECT 241.400 113.800 241.800 114.200 ;
        RECT 243.800 113.800 244.200 114.600 ;
        RECT 237.400 113.400 238.700 113.700 ;
        RECT 229.400 112.800 230.300 113.100 ;
        RECT 229.900 111.100 230.300 112.800 ;
        RECT 231.000 111.100 231.400 113.100 ;
        RECT 231.800 113.000 233.800 113.100 ;
        RECT 231.800 111.100 232.200 113.000 ;
        RECT 233.400 111.100 233.800 113.000 ;
        RECT 235.800 111.100 236.200 113.200 ;
        RECT 236.600 112.800 237.000 113.200 ;
        RECT 236.500 112.400 236.900 112.800 ;
        RECT 237.400 111.100 237.800 113.400 ;
        RECT 239.200 113.100 239.500 113.800 ;
        RECT 241.500 113.100 241.800 113.800 ;
        RECT 242.200 113.100 242.600 113.200 ;
        RECT 239.000 112.800 239.500 113.100 ;
        RECT 241.400 112.800 242.600 113.100 ;
        RECT 244.600 113.100 244.900 114.900 ;
        RECT 245.400 114.800 245.800 114.900 ;
        RECT 246.200 113.600 246.600 115.300 ;
        RECT 247.900 115.200 248.300 115.300 ;
        RECT 247.100 114.900 247.500 115.000 ;
        RECT 247.100 114.600 249.000 114.900 ;
        RECT 248.600 114.500 249.000 114.600 ;
        RECT 249.500 114.200 249.800 115.800 ;
        RECT 250.500 115.900 250.800 116.500 ;
        RECT 251.100 116.500 251.500 116.600 ;
        RECT 253.400 116.500 253.800 116.600 ;
        RECT 251.100 116.200 253.800 116.500 ;
        RECT 250.500 115.700 252.900 115.900 ;
        RECT 255.000 115.700 255.400 119.900 ;
        RECT 250.500 115.600 255.400 115.700 ;
        RECT 252.500 115.500 255.400 115.600 ;
        RECT 252.600 115.400 255.400 115.500 ;
        RECT 255.800 115.700 256.200 119.900 ;
        RECT 258.000 118.200 258.400 119.900 ;
        RECT 257.400 117.900 258.400 118.200 ;
        RECT 260.200 117.900 260.600 119.900 ;
        RECT 262.300 117.900 262.900 119.900 ;
        RECT 257.400 117.500 257.800 117.900 ;
        RECT 260.200 117.600 260.500 117.900 ;
        RECT 259.100 117.300 260.900 117.600 ;
        RECT 262.200 117.500 262.600 117.900 ;
        RECT 259.100 117.200 259.500 117.300 ;
        RECT 260.500 117.200 260.900 117.300 ;
        RECT 257.400 116.500 257.800 116.600 ;
        RECT 259.700 116.500 260.100 116.600 ;
        RECT 257.400 116.200 260.100 116.500 ;
        RECT 260.400 116.500 261.500 116.800 ;
        RECT 260.400 115.900 260.700 116.500 ;
        RECT 261.100 116.400 261.500 116.500 ;
        RECT 262.300 116.600 263.000 117.000 ;
        RECT 262.300 116.100 262.600 116.600 ;
        RECT 258.300 115.700 260.700 115.900 ;
        RECT 255.800 115.600 260.700 115.700 ;
        RECT 261.400 115.800 262.600 116.100 ;
        RECT 255.800 115.500 258.700 115.600 ;
        RECT 255.800 115.400 258.600 115.500 ;
        RECT 251.800 115.100 252.200 115.200 ;
        RECT 259.000 115.100 259.400 115.200 ;
        RECT 251.800 114.800 254.300 115.100 ;
        RECT 253.900 114.700 254.300 114.800 ;
        RECT 256.900 114.800 259.400 115.100 ;
        RECT 256.900 114.700 257.300 114.800 ;
        RECT 258.200 114.700 258.600 114.800 ;
        RECT 253.100 114.200 253.500 114.300 ;
        RECT 257.700 114.200 258.100 114.300 ;
        RECT 261.400 114.200 261.700 115.800 ;
        RECT 264.600 115.600 265.000 119.900 ;
        RECT 262.900 115.300 265.000 115.600 ;
        RECT 262.900 115.200 263.300 115.300 ;
        RECT 263.700 114.900 264.100 115.000 ;
        RECT 262.200 114.600 264.100 114.900 ;
        RECT 262.200 114.500 262.600 114.600 ;
        RECT 249.500 113.900 255.000 114.200 ;
        RECT 249.700 113.800 250.100 113.900 ;
        RECT 246.200 113.300 248.100 113.600 ;
        RECT 239.000 111.100 239.400 112.800 ;
        RECT 241.500 112.100 241.800 112.800 ;
        RECT 241.400 111.100 241.800 112.100 ;
        RECT 244.600 111.100 245.000 113.100 ;
        RECT 245.400 112.800 245.800 113.200 ;
        RECT 245.300 112.400 245.700 112.800 ;
        RECT 246.200 111.100 246.600 113.300 ;
        RECT 247.700 113.200 248.100 113.300 ;
        RECT 252.600 112.800 252.900 113.900 ;
        RECT 254.200 113.800 255.000 113.900 ;
        RECT 256.200 113.900 261.700 114.200 ;
        RECT 256.200 113.800 257.000 113.900 ;
        RECT 251.700 112.700 252.100 112.800 ;
        RECT 248.600 112.100 249.000 112.500 ;
        RECT 250.700 112.400 252.100 112.700 ;
        RECT 252.600 112.400 253.000 112.800 ;
        RECT 250.700 112.100 251.000 112.400 ;
        RECT 253.400 112.100 253.800 112.500 ;
        RECT 248.300 111.800 249.000 112.100 ;
        RECT 248.300 111.100 248.900 111.800 ;
        RECT 250.600 111.100 251.000 112.100 ;
        RECT 252.800 111.800 253.800 112.100 ;
        RECT 252.800 111.100 253.200 111.800 ;
        RECT 255.000 111.100 255.400 113.500 ;
        RECT 255.800 111.100 256.200 113.500 ;
        RECT 258.300 112.800 258.600 113.900 ;
        RECT 261.100 113.800 261.500 113.900 ;
        RECT 264.600 113.600 265.000 115.300 ;
        RECT 263.100 113.300 265.000 113.600 ;
        RECT 263.100 113.200 263.500 113.300 ;
        RECT 257.400 112.100 257.800 112.500 ;
        RECT 258.200 112.400 258.600 112.800 ;
        RECT 259.100 112.700 259.500 112.800 ;
        RECT 259.100 112.400 260.500 112.700 ;
        RECT 260.200 112.100 260.500 112.400 ;
        RECT 262.200 112.100 262.600 112.500 ;
        RECT 257.400 111.800 258.400 112.100 ;
        RECT 258.000 111.100 258.400 111.800 ;
        RECT 260.200 111.100 260.600 112.100 ;
        RECT 262.200 111.800 262.900 112.100 ;
        RECT 262.300 111.100 262.900 111.800 ;
        RECT 264.600 111.100 265.000 113.300 ;
        RECT 1.400 107.600 1.800 109.900 ;
        RECT 3.000 107.600 3.400 109.900 ;
        RECT 1.400 107.200 3.400 107.600 ;
        RECT 4.600 107.500 5.000 109.900 ;
        RECT 6.800 109.200 7.200 109.900 ;
        RECT 6.200 108.900 7.200 109.200 ;
        RECT 9.000 108.900 9.400 109.900 ;
        RECT 11.100 109.200 11.700 109.900 ;
        RECT 11.000 108.900 11.700 109.200 ;
        RECT 6.200 108.500 6.600 108.900 ;
        RECT 9.000 108.600 9.300 108.900 ;
        RECT 7.000 107.800 7.400 108.600 ;
        RECT 7.900 108.300 9.300 108.600 ;
        RECT 11.000 108.500 11.400 108.900 ;
        RECT 7.900 108.200 8.300 108.300 ;
        RECT 3.000 105.800 3.400 107.200 ;
        RECT 5.000 107.100 5.800 107.200 ;
        RECT 7.100 107.100 7.400 107.800 ;
        RECT 11.900 107.700 12.300 107.800 ;
        RECT 13.400 107.700 13.800 109.900 ;
        RECT 11.900 107.400 13.800 107.700 ;
        RECT 8.600 107.100 9.000 107.200 ;
        RECT 9.900 107.100 10.300 107.200 ;
        RECT 5.000 106.800 10.500 107.100 ;
        RECT 6.500 106.700 6.900 106.800 ;
        RECT 5.700 106.200 6.100 106.300 ;
        RECT 5.700 105.900 8.200 106.200 ;
        RECT 7.800 105.800 8.200 105.900 ;
        RECT 1.400 105.400 3.400 105.800 ;
        RECT 1.400 101.100 1.800 105.400 ;
        RECT 3.000 101.100 3.400 105.400 ;
        RECT 4.600 105.500 7.400 105.600 ;
        RECT 4.600 105.400 7.500 105.500 ;
        RECT 4.600 105.300 9.500 105.400 ;
        RECT 4.600 101.100 5.000 105.300 ;
        RECT 7.100 105.100 9.500 105.300 ;
        RECT 6.200 104.500 8.900 104.800 ;
        RECT 6.200 104.400 6.600 104.500 ;
        RECT 8.500 104.400 8.900 104.500 ;
        RECT 9.200 104.500 9.500 105.100 ;
        RECT 10.200 105.200 10.500 106.800 ;
        RECT 11.000 106.400 11.400 106.500 ;
        RECT 11.000 106.100 12.900 106.400 ;
        RECT 12.500 106.000 12.900 106.100 ;
        RECT 11.700 105.700 12.100 105.800 ;
        RECT 13.400 105.700 13.800 107.400 ;
        RECT 15.800 107.900 16.200 109.900 ;
        RECT 18.200 108.900 18.600 109.900 ;
        RECT 16.500 108.200 16.900 108.600 ;
        RECT 16.600 108.100 17.000 108.200 ;
        RECT 18.200 108.100 18.500 108.900 ;
        RECT 15.000 106.400 15.400 107.200 ;
        RECT 15.800 106.200 16.100 107.900 ;
        RECT 16.600 107.800 18.500 108.100 ;
        RECT 19.000 107.800 19.400 108.600 ;
        RECT 18.200 107.200 18.500 107.800 ;
        RECT 19.800 107.500 20.200 109.900 ;
        RECT 22.000 109.200 22.400 109.900 ;
        RECT 21.400 108.900 22.400 109.200 ;
        RECT 24.200 108.900 24.600 109.900 ;
        RECT 26.300 109.200 26.900 109.900 ;
        RECT 26.200 108.900 26.900 109.200 ;
        RECT 21.400 108.500 21.800 108.900 ;
        RECT 24.200 108.600 24.500 108.900 ;
        RECT 22.200 108.200 22.600 108.600 ;
        RECT 23.100 108.300 24.500 108.600 ;
        RECT 26.200 108.500 26.600 108.900 ;
        RECT 23.100 108.200 23.500 108.300 ;
        RECT 18.200 106.800 18.600 107.200 ;
        RECT 20.200 107.100 21.000 107.200 ;
        RECT 22.300 107.100 22.600 108.200 ;
        RECT 27.100 107.700 27.500 107.800 ;
        RECT 28.600 107.700 29.000 109.900 ;
        RECT 27.100 107.400 29.000 107.700 ;
        RECT 25.100 107.100 25.500 107.200 ;
        RECT 20.200 106.800 25.700 107.100 ;
        RECT 14.200 106.100 14.600 106.200 ;
        RECT 15.800 106.100 16.200 106.200 ;
        RECT 16.600 106.100 17.000 106.200 ;
        RECT 14.200 105.800 15.000 106.100 ;
        RECT 15.800 105.800 17.000 106.100 ;
        RECT 11.700 105.400 13.800 105.700 ;
        RECT 14.600 105.600 15.000 105.800 ;
        RECT 10.200 104.900 11.400 105.200 ;
        RECT 9.900 104.500 10.300 104.600 ;
        RECT 9.200 104.200 10.300 104.500 ;
        RECT 11.100 104.400 11.400 104.900 ;
        RECT 11.100 104.000 11.800 104.400 ;
        RECT 7.900 103.700 8.300 103.800 ;
        RECT 9.300 103.700 9.700 103.800 ;
        RECT 6.200 103.100 6.600 103.500 ;
        RECT 7.900 103.400 9.700 103.700 ;
        RECT 9.000 103.100 9.300 103.400 ;
        RECT 11.000 103.100 11.400 103.500 ;
        RECT 6.200 102.800 7.200 103.100 ;
        RECT 6.800 101.100 7.200 102.800 ;
        RECT 9.000 101.100 9.400 103.100 ;
        RECT 11.100 101.100 11.700 103.100 ;
        RECT 13.400 101.100 13.800 105.400 ;
        RECT 16.600 105.100 16.900 105.800 ;
        RECT 17.400 105.400 17.800 106.200 ;
        RECT 18.200 105.100 18.500 106.800 ;
        RECT 21.700 106.700 22.100 106.800 ;
        RECT 20.900 106.200 21.300 106.300 ;
        RECT 20.900 106.100 23.400 106.200 ;
        RECT 24.600 106.100 25.000 106.200 ;
        RECT 20.900 105.900 25.000 106.100 ;
        RECT 23.000 105.800 25.000 105.900 ;
        RECT 19.800 105.500 22.600 105.600 ;
        RECT 19.800 105.400 22.700 105.500 ;
        RECT 19.800 105.300 24.700 105.400 ;
        RECT 14.200 104.800 16.200 105.100 ;
        RECT 14.200 101.100 14.600 104.800 ;
        RECT 15.800 101.100 16.200 104.800 ;
        RECT 16.600 101.100 17.000 105.100 ;
        RECT 17.700 104.700 18.600 105.100 ;
        RECT 17.700 101.100 18.100 104.700 ;
        RECT 19.800 101.100 20.200 105.300 ;
        RECT 22.300 105.100 24.700 105.300 ;
        RECT 21.400 104.500 24.100 104.800 ;
        RECT 21.400 104.400 21.800 104.500 ;
        RECT 23.700 104.400 24.100 104.500 ;
        RECT 24.400 104.500 24.700 105.100 ;
        RECT 25.400 105.200 25.700 106.800 ;
        RECT 26.200 106.400 26.600 106.500 ;
        RECT 26.200 106.100 28.100 106.400 ;
        RECT 27.700 106.000 28.100 106.100 ;
        RECT 26.900 105.700 27.300 105.800 ;
        RECT 28.600 105.700 29.000 107.400 ;
        RECT 29.400 108.500 29.800 109.500 ;
        RECT 29.400 107.400 29.700 108.500 ;
        RECT 31.500 108.000 31.900 109.500 ;
        RECT 31.500 107.700 32.300 108.000 ;
        RECT 34.200 107.800 34.600 108.600 ;
        RECT 31.900 107.500 32.300 107.700 ;
        RECT 29.400 107.100 31.500 107.400 ;
        RECT 31.000 106.900 31.500 107.100 ;
        RECT 32.000 107.200 32.300 107.500 ;
        RECT 32.000 107.100 33.000 107.200 ;
        RECT 33.400 107.100 33.800 107.200 ;
        RECT 29.400 105.800 29.800 106.600 ;
        RECT 30.200 105.800 30.600 106.600 ;
        RECT 31.000 106.500 31.700 106.900 ;
        RECT 32.000 106.800 33.800 107.100 ;
        RECT 26.900 105.400 29.000 105.700 ;
        RECT 31.000 105.500 31.300 106.500 ;
        RECT 25.400 104.900 26.600 105.200 ;
        RECT 25.100 104.500 25.500 104.600 ;
        RECT 24.400 104.200 25.500 104.500 ;
        RECT 26.300 104.400 26.600 104.900 ;
        RECT 26.300 104.000 27.000 104.400 ;
        RECT 23.100 103.700 23.500 103.800 ;
        RECT 24.500 103.700 24.900 103.800 ;
        RECT 21.400 103.100 21.800 103.500 ;
        RECT 23.100 103.400 24.900 103.700 ;
        RECT 24.200 103.100 24.500 103.400 ;
        RECT 26.200 103.100 26.600 103.500 ;
        RECT 21.400 102.800 22.400 103.100 ;
        RECT 22.000 101.100 22.400 102.800 ;
        RECT 24.200 101.100 24.600 103.100 ;
        RECT 26.300 101.100 26.900 103.100 ;
        RECT 28.600 101.100 29.000 105.400 ;
        RECT 29.400 105.200 31.300 105.500 ;
        RECT 29.400 103.500 29.700 105.200 ;
        RECT 32.000 104.900 32.300 106.800 ;
        RECT 32.600 106.100 33.000 106.200 ;
        RECT 34.200 106.100 34.600 106.200 ;
        RECT 32.600 105.800 34.600 106.100 ;
        RECT 35.000 106.100 35.400 109.900 ;
        RECT 37.700 108.000 38.100 109.500 ;
        RECT 39.800 108.500 40.200 109.500 ;
        RECT 42.500 109.200 42.900 109.500 ;
        RECT 42.200 108.800 42.900 109.200 ;
        RECT 37.300 107.700 38.100 108.000 ;
        RECT 37.300 107.500 37.700 107.700 ;
        RECT 37.300 107.200 37.600 107.500 ;
        RECT 39.900 107.400 40.200 108.500 ;
        RECT 42.500 108.000 42.900 108.800 ;
        RECT 44.600 108.500 45.000 109.500 ;
        RECT 36.600 106.800 37.600 107.200 ;
        RECT 38.100 107.100 40.200 107.400 ;
        RECT 42.100 107.700 42.900 108.000 ;
        RECT 42.100 107.500 42.500 107.700 ;
        RECT 42.100 107.200 42.400 107.500 ;
        RECT 44.700 107.400 45.000 108.500 ;
        RECT 38.100 106.900 38.600 107.100 ;
        RECT 36.600 106.100 37.000 106.200 ;
        RECT 35.000 105.800 37.000 106.100 ;
        RECT 32.600 105.400 33.000 105.800 ;
        RECT 31.500 104.600 32.300 104.900 ;
        RECT 29.400 101.500 29.800 103.500 ;
        RECT 31.500 101.100 31.900 104.600 ;
        RECT 35.000 101.100 35.400 105.800 ;
        RECT 36.600 105.400 37.000 105.800 ;
        RECT 37.300 105.200 37.600 106.800 ;
        RECT 37.900 106.500 38.600 106.900 ;
        RECT 41.400 106.800 42.400 107.200 ;
        RECT 42.900 107.100 45.000 107.400 ;
        RECT 45.400 107.700 45.800 109.900 ;
        RECT 47.500 109.200 48.100 109.900 ;
        RECT 47.500 108.900 48.200 109.200 ;
        RECT 49.800 108.900 50.200 109.900 ;
        RECT 52.000 109.200 52.400 109.900 ;
        RECT 52.000 108.900 53.000 109.200 ;
        RECT 47.800 108.500 48.200 108.900 ;
        RECT 49.900 108.600 50.200 108.900 ;
        RECT 49.900 108.300 51.300 108.600 ;
        RECT 50.900 108.200 51.300 108.300 ;
        RECT 51.800 108.200 52.200 108.600 ;
        RECT 52.600 108.500 53.000 108.900 ;
        RECT 46.900 107.700 47.300 107.800 ;
        RECT 45.400 107.400 47.300 107.700 ;
        RECT 42.900 106.900 43.400 107.100 ;
        RECT 38.300 105.500 38.600 106.500 ;
        RECT 39.000 105.800 39.400 106.600 ;
        RECT 39.800 105.800 40.200 106.600 ;
        RECT 38.300 105.200 40.200 105.500 ;
        RECT 41.400 105.400 41.800 106.200 ;
        RECT 37.300 104.900 37.800 105.200 ;
        RECT 37.300 104.600 38.100 104.900 ;
        RECT 37.700 101.100 38.100 104.600 ;
        RECT 39.900 103.500 40.200 105.200 ;
        RECT 42.100 104.900 42.400 106.800 ;
        RECT 42.700 106.500 43.400 106.900 ;
        RECT 43.100 105.500 43.400 106.500 ;
        RECT 43.800 105.800 44.200 106.600 ;
        RECT 44.600 105.800 45.000 106.600 ;
        RECT 45.400 105.700 45.800 107.400 ;
        RECT 48.900 107.100 49.300 107.200 ;
        RECT 51.000 107.100 51.400 107.200 ;
        RECT 51.800 107.100 52.100 108.200 ;
        RECT 54.200 107.500 54.600 109.900 ;
        RECT 57.400 108.200 57.800 109.900 ;
        RECT 57.300 107.900 57.800 108.200 ;
        RECT 57.300 107.200 57.600 107.900 ;
        RECT 59.000 107.600 59.400 109.900 ;
        RECT 58.100 107.300 59.400 107.600 ;
        RECT 59.800 107.500 60.200 109.900 ;
        RECT 62.000 109.200 62.400 109.900 ;
        RECT 61.400 108.900 62.400 109.200 ;
        RECT 64.200 108.900 64.600 109.900 ;
        RECT 66.300 109.200 66.900 109.900 ;
        RECT 66.200 108.900 66.900 109.200 ;
        RECT 61.400 108.500 61.800 108.900 ;
        RECT 64.200 108.600 64.500 108.900 ;
        RECT 62.200 108.200 62.600 108.600 ;
        RECT 63.100 108.300 64.500 108.600 ;
        RECT 66.200 108.500 66.600 108.900 ;
        RECT 63.100 108.200 63.500 108.300 ;
        RECT 53.400 107.100 54.200 107.200 ;
        RECT 48.700 106.800 54.200 107.100 ;
        RECT 55.000 107.100 55.400 107.200 ;
        RECT 57.300 107.100 57.800 107.200 ;
        RECT 55.000 106.800 57.800 107.100 ;
        RECT 47.800 106.400 48.200 106.500 ;
        RECT 46.300 106.100 48.200 106.400 ;
        RECT 46.300 106.000 46.700 106.100 ;
        RECT 47.100 105.700 47.500 105.800 ;
        RECT 43.100 105.200 45.000 105.500 ;
        RECT 42.100 104.600 42.900 104.900 ;
        RECT 39.800 101.500 40.200 103.500 ;
        RECT 42.500 101.100 42.900 104.600 ;
        RECT 44.700 103.500 45.000 105.200 ;
        RECT 44.600 101.500 45.000 103.500 ;
        RECT 45.400 105.400 47.500 105.700 ;
        RECT 45.400 101.100 45.800 105.400 ;
        RECT 48.700 105.200 49.000 106.800 ;
        RECT 52.300 106.700 52.700 106.800 ;
        RECT 53.100 106.200 53.500 106.300 ;
        RECT 51.000 105.900 53.500 106.200 ;
        RECT 51.000 105.800 51.400 105.900 ;
        RECT 51.800 105.500 54.600 105.600 ;
        RECT 51.700 105.400 54.600 105.500 ;
        RECT 47.800 104.900 49.000 105.200 ;
        RECT 49.700 105.300 54.600 105.400 ;
        RECT 49.700 105.100 52.100 105.300 ;
        RECT 47.800 104.400 48.100 104.900 ;
        RECT 47.400 104.000 48.100 104.400 ;
        RECT 48.900 104.500 49.300 104.600 ;
        RECT 49.700 104.500 50.000 105.100 ;
        RECT 48.900 104.200 50.000 104.500 ;
        RECT 50.300 104.500 53.000 104.800 ;
        RECT 50.300 104.400 50.700 104.500 ;
        RECT 52.600 104.400 53.000 104.500 ;
        RECT 49.500 103.700 49.900 103.800 ;
        RECT 50.900 103.700 51.300 103.800 ;
        RECT 47.800 103.100 48.200 103.500 ;
        RECT 49.500 103.400 51.300 103.700 ;
        RECT 49.900 103.100 50.200 103.400 ;
        RECT 52.600 103.100 53.000 103.500 ;
        RECT 47.500 101.100 48.100 103.100 ;
        RECT 49.800 101.100 50.200 103.100 ;
        RECT 52.000 102.800 53.000 103.100 ;
        RECT 52.000 101.100 52.400 102.800 ;
        RECT 54.200 101.100 54.600 105.300 ;
        RECT 57.300 105.100 57.600 106.800 ;
        RECT 58.100 106.500 58.400 107.300 ;
        RECT 60.200 107.100 61.000 107.200 ;
        RECT 62.300 107.100 62.600 108.200 ;
        RECT 67.100 107.700 67.500 107.800 ;
        RECT 68.600 107.700 69.000 109.900 ;
        RECT 69.400 108.000 69.800 109.900 ;
        RECT 71.000 108.000 71.400 109.900 ;
        RECT 69.400 107.900 71.400 108.000 ;
        RECT 71.800 107.900 72.200 109.900 ;
        RECT 72.900 108.200 73.300 109.900 ;
        RECT 72.900 107.900 73.800 108.200 ;
        RECT 69.500 107.700 71.300 107.900 ;
        RECT 67.100 107.400 69.000 107.700 ;
        RECT 65.100 107.100 65.500 107.200 ;
        RECT 60.200 106.800 65.700 107.100 ;
        RECT 61.700 106.700 62.100 106.800 ;
        RECT 57.900 106.100 58.400 106.500 ;
        RECT 58.100 105.100 58.400 106.100 ;
        RECT 58.900 106.200 59.300 106.600 ;
        RECT 60.900 106.200 61.300 106.300 ;
        RECT 62.200 106.200 62.600 106.300 ;
        RECT 65.400 106.200 65.700 106.800 ;
        RECT 66.200 106.400 66.600 106.500 ;
        RECT 58.900 105.800 59.400 106.200 ;
        RECT 60.900 105.900 63.400 106.200 ;
        RECT 63.000 105.800 63.400 105.900 ;
        RECT 65.400 105.800 65.800 106.200 ;
        RECT 66.200 106.100 68.100 106.400 ;
        RECT 67.700 106.000 68.100 106.100 ;
        RECT 59.800 105.500 62.600 105.600 ;
        RECT 59.800 105.400 62.700 105.500 ;
        RECT 59.800 105.300 64.700 105.400 ;
        RECT 57.300 104.600 57.800 105.100 ;
        RECT 58.100 104.800 59.400 105.100 ;
        RECT 57.400 101.100 57.800 104.600 ;
        RECT 59.000 101.100 59.400 104.800 ;
        RECT 59.800 101.100 60.200 105.300 ;
        RECT 62.300 105.100 64.700 105.300 ;
        RECT 61.400 104.500 64.100 104.800 ;
        RECT 61.400 104.400 61.800 104.500 ;
        RECT 63.700 104.400 64.100 104.500 ;
        RECT 64.400 104.500 64.700 105.100 ;
        RECT 65.400 105.200 65.700 105.800 ;
        RECT 66.900 105.700 67.300 105.800 ;
        RECT 68.600 105.700 69.000 107.400 ;
        RECT 69.800 107.200 70.200 107.400 ;
        RECT 71.800 107.200 72.100 107.900 ;
        RECT 69.400 106.900 70.200 107.200 ;
        RECT 70.900 107.100 72.200 107.200 ;
        RECT 72.600 107.100 73.000 107.200 ;
        RECT 69.400 106.800 69.800 106.900 ;
        RECT 70.900 106.800 73.000 107.100 ;
        RECT 70.200 105.800 70.600 106.600 ;
        RECT 66.900 105.400 69.000 105.700 ;
        RECT 65.400 104.900 66.600 105.200 ;
        RECT 65.100 104.500 65.500 104.600 ;
        RECT 64.400 104.200 65.500 104.500 ;
        RECT 66.300 104.400 66.600 104.900 ;
        RECT 66.300 104.000 67.000 104.400 ;
        RECT 63.100 103.700 63.500 103.800 ;
        RECT 64.500 103.700 64.900 103.800 ;
        RECT 61.400 103.100 61.800 103.500 ;
        RECT 63.100 103.400 64.900 103.700 ;
        RECT 64.200 103.100 64.500 103.400 ;
        RECT 66.200 103.100 66.600 103.500 ;
        RECT 61.400 102.800 62.400 103.100 ;
        RECT 62.000 101.100 62.400 102.800 ;
        RECT 64.200 101.100 64.600 103.100 ;
        RECT 66.300 101.100 66.900 103.100 ;
        RECT 68.600 101.100 69.000 105.400 ;
        RECT 70.900 105.100 71.200 106.800 ;
        RECT 73.400 106.100 73.800 107.900 ;
        RECT 74.200 106.800 74.600 107.600 ;
        RECT 75.000 107.500 75.400 109.900 ;
        RECT 77.200 109.200 77.600 109.900 ;
        RECT 76.600 108.900 77.600 109.200 ;
        RECT 79.400 108.900 79.800 109.900 ;
        RECT 81.500 109.200 82.100 109.900 ;
        RECT 81.400 108.900 82.100 109.200 ;
        RECT 76.600 108.500 77.000 108.900 ;
        RECT 79.400 108.600 79.700 108.900 ;
        RECT 77.400 108.200 77.800 108.600 ;
        RECT 78.300 108.300 79.700 108.600 ;
        RECT 81.400 108.500 81.800 108.900 ;
        RECT 78.300 108.200 78.700 108.300 ;
        RECT 75.400 107.100 76.200 107.200 ;
        RECT 77.500 107.100 77.800 108.200 ;
        RECT 82.300 107.700 82.700 107.800 ;
        RECT 83.800 107.700 84.200 109.900 ;
        RECT 85.400 108.900 85.800 109.900 ;
        RECT 84.600 107.800 85.000 108.600 ;
        RECT 85.500 108.100 85.800 108.900 ;
        RECT 87.100 108.200 87.500 108.600 ;
        RECT 87.000 108.100 87.400 108.200 ;
        RECT 85.400 107.800 87.400 108.100 ;
        RECT 87.800 107.900 88.200 109.900 ;
        RECT 82.300 107.400 84.200 107.700 ;
        RECT 80.300 107.100 80.700 107.200 ;
        RECT 75.400 106.800 80.900 107.100 ;
        RECT 76.900 106.700 77.300 106.800 ;
        RECT 71.800 105.800 73.800 106.100 ;
        RECT 76.100 106.200 76.500 106.300 ;
        RECT 77.400 106.200 77.800 106.300 ;
        RECT 80.600 106.200 80.900 106.800 ;
        RECT 81.400 106.400 81.800 106.500 ;
        RECT 76.100 105.900 78.600 106.200 ;
        RECT 78.200 105.800 78.600 105.900 ;
        RECT 80.600 105.800 81.000 106.200 ;
        RECT 81.400 106.100 83.300 106.400 ;
        RECT 82.900 106.000 83.300 106.100 ;
        RECT 71.800 105.200 72.100 105.800 ;
        RECT 71.800 105.100 72.200 105.200 ;
        RECT 70.700 104.800 71.200 105.100 ;
        RECT 71.500 104.800 72.200 105.100 ;
        RECT 70.700 101.100 71.100 104.800 ;
        RECT 71.500 104.200 71.800 104.800 ;
        RECT 72.600 104.400 73.000 105.200 ;
        RECT 71.400 103.800 71.800 104.200 ;
        RECT 73.400 101.100 73.800 105.800 ;
        RECT 75.000 105.500 77.800 105.600 ;
        RECT 75.000 105.400 77.900 105.500 ;
        RECT 75.000 105.300 79.900 105.400 ;
        RECT 75.000 101.100 75.400 105.300 ;
        RECT 77.500 105.100 79.900 105.300 ;
        RECT 76.600 104.500 79.300 104.800 ;
        RECT 76.600 104.400 77.000 104.500 ;
        RECT 78.900 104.400 79.300 104.500 ;
        RECT 79.600 104.500 79.900 105.100 ;
        RECT 80.600 105.200 80.900 105.800 ;
        RECT 82.100 105.700 82.500 105.800 ;
        RECT 83.800 105.700 84.200 107.400 ;
        RECT 85.500 107.200 85.800 107.800 ;
        RECT 85.400 106.800 85.800 107.200 ;
        RECT 82.100 105.400 84.200 105.700 ;
        RECT 80.600 104.900 81.800 105.200 ;
        RECT 80.300 104.500 80.700 104.600 ;
        RECT 79.600 104.200 80.700 104.500 ;
        RECT 81.500 104.400 81.800 104.900 ;
        RECT 81.500 104.000 82.200 104.400 ;
        RECT 78.300 103.700 78.700 103.800 ;
        RECT 79.700 103.700 80.100 103.800 ;
        RECT 76.600 103.100 77.000 103.500 ;
        RECT 78.300 103.400 80.100 103.700 ;
        RECT 79.400 103.100 79.700 103.400 ;
        RECT 81.400 103.100 81.800 103.500 ;
        RECT 76.600 102.800 77.600 103.100 ;
        RECT 77.200 101.100 77.600 102.800 ;
        RECT 79.400 101.100 79.800 103.100 ;
        RECT 81.500 101.100 82.100 103.100 ;
        RECT 83.800 101.100 84.200 105.400 ;
        RECT 85.500 105.100 85.800 106.800 ;
        RECT 87.900 106.200 88.200 107.900 ;
        RECT 90.200 107.500 90.600 109.900 ;
        RECT 92.400 109.200 92.800 109.900 ;
        RECT 91.800 108.900 92.800 109.200 ;
        RECT 94.600 108.900 95.000 109.900 ;
        RECT 96.700 109.200 97.300 109.900 ;
        RECT 96.600 108.900 97.300 109.200 ;
        RECT 91.800 108.500 92.200 108.900 ;
        RECT 94.600 108.600 94.900 108.900 ;
        RECT 92.600 108.200 93.000 108.600 ;
        RECT 93.500 108.300 94.900 108.600 ;
        RECT 96.600 108.500 97.000 108.900 ;
        RECT 93.500 108.200 93.900 108.300 ;
        RECT 92.700 107.200 93.000 108.200 ;
        RECT 97.500 107.700 97.900 107.800 ;
        RECT 99.000 107.700 99.400 109.900 ;
        RECT 100.600 108.200 101.000 109.900 ;
        RECT 97.500 107.400 99.400 107.700 ;
        RECT 88.600 106.400 89.000 107.200 ;
        RECT 90.600 107.100 91.400 107.200 ;
        RECT 92.600 107.100 93.000 107.200 ;
        RECT 95.500 107.100 95.900 107.200 ;
        RECT 90.600 106.800 96.100 107.100 ;
        RECT 92.100 106.700 92.500 106.800 ;
        RECT 91.300 106.200 91.700 106.300 ;
        RECT 86.200 105.400 86.600 106.200 ;
        RECT 87.000 106.100 87.400 106.200 ;
        RECT 87.800 106.100 88.200 106.200 ;
        RECT 89.400 106.100 89.800 106.200 ;
        RECT 87.000 105.800 88.200 106.100 ;
        RECT 89.000 105.800 89.800 106.100 ;
        RECT 91.300 105.900 93.800 106.200 ;
        RECT 93.400 105.800 93.800 105.900 ;
        RECT 87.100 105.100 87.400 105.800 ;
        RECT 89.000 105.600 89.400 105.800 ;
        RECT 90.200 105.500 93.000 105.600 ;
        RECT 90.200 105.400 93.100 105.500 ;
        RECT 90.200 105.300 95.100 105.400 ;
        RECT 85.400 104.700 86.300 105.100 ;
        RECT 85.900 101.100 86.300 104.700 ;
        RECT 87.000 101.100 87.400 105.100 ;
        RECT 87.800 104.800 89.800 105.100 ;
        RECT 87.800 101.100 88.200 104.800 ;
        RECT 89.400 101.100 89.800 104.800 ;
        RECT 90.200 101.100 90.600 105.300 ;
        RECT 92.700 105.100 95.100 105.300 ;
        RECT 91.800 104.500 94.500 104.800 ;
        RECT 91.800 104.400 92.200 104.500 ;
        RECT 94.100 104.400 94.500 104.500 ;
        RECT 94.800 104.500 95.100 105.100 ;
        RECT 95.800 105.200 96.100 106.800 ;
        RECT 96.600 106.400 97.000 106.500 ;
        RECT 96.600 106.100 98.500 106.400 ;
        RECT 98.100 106.000 98.500 106.100 ;
        RECT 97.300 105.700 97.700 105.800 ;
        RECT 99.000 105.700 99.400 107.400 ;
        RECT 100.500 107.900 101.000 108.200 ;
        RECT 100.500 107.200 100.800 107.900 ;
        RECT 102.200 107.600 102.600 109.900 ;
        RECT 101.300 107.300 102.600 107.600 ;
        RECT 104.600 107.900 105.000 109.900 ;
        RECT 108.600 108.900 109.000 109.900 ;
        RECT 105.300 108.200 105.700 108.600 ;
        RECT 99.800 107.100 100.200 107.200 ;
        RECT 100.500 107.100 101.000 107.200 ;
        RECT 99.800 106.800 101.000 107.100 ;
        RECT 97.300 105.400 99.400 105.700 ;
        RECT 95.800 104.900 97.000 105.200 ;
        RECT 95.500 104.500 95.900 104.600 ;
        RECT 94.800 104.200 95.900 104.500 ;
        RECT 96.700 104.400 97.000 104.900 ;
        RECT 96.700 104.000 97.400 104.400 ;
        RECT 93.500 103.700 93.900 103.800 ;
        RECT 94.900 103.700 95.300 103.800 ;
        RECT 91.800 103.100 92.200 103.500 ;
        RECT 93.500 103.400 95.300 103.700 ;
        RECT 94.600 103.100 94.900 103.400 ;
        RECT 96.600 103.100 97.000 103.500 ;
        RECT 91.800 102.800 92.800 103.100 ;
        RECT 92.400 101.100 92.800 102.800 ;
        RECT 94.600 101.100 95.000 103.100 ;
        RECT 96.700 101.100 97.300 103.100 ;
        RECT 99.000 101.100 99.400 105.400 ;
        RECT 100.500 105.100 100.800 106.800 ;
        RECT 101.300 106.500 101.600 107.300 ;
        RECT 101.100 106.100 101.600 106.500 ;
        RECT 101.300 105.100 101.600 106.100 ;
        RECT 102.100 106.200 102.500 106.600 ;
        RECT 103.800 106.400 104.200 107.200 ;
        RECT 102.100 105.800 102.600 106.200 ;
        RECT 103.000 106.100 103.400 106.200 ;
        RECT 104.600 106.100 104.900 107.900 ;
        RECT 105.400 107.800 105.800 108.200 ;
        RECT 106.200 108.100 106.600 108.200 ;
        RECT 107.800 108.100 108.200 108.600 ;
        RECT 106.200 107.800 108.200 108.100 ;
        RECT 105.400 107.100 105.700 107.800 ;
        RECT 108.700 107.200 109.000 108.900 ;
        RECT 108.600 107.100 109.000 107.200 ;
        RECT 110.200 108.500 110.600 109.500 ;
        RECT 112.300 109.200 112.700 109.500 ;
        RECT 112.300 108.800 113.000 109.200 ;
        RECT 110.200 107.400 110.500 108.500 ;
        RECT 112.300 108.000 112.700 108.800 ;
        RECT 112.300 107.700 113.100 108.000 ;
        RECT 112.700 107.500 113.100 107.700 ;
        RECT 110.200 107.100 112.300 107.400 ;
        RECT 105.400 106.800 109.000 107.100 ;
        RECT 105.400 106.100 105.800 106.200 ;
        RECT 103.000 105.800 103.800 106.100 ;
        RECT 104.600 105.800 105.800 106.100 ;
        RECT 103.400 105.600 103.800 105.800 ;
        RECT 105.400 105.100 105.700 105.800 ;
        RECT 108.700 105.100 109.000 106.800 ;
        RECT 111.800 106.900 112.300 107.100 ;
        RECT 112.800 107.200 113.100 107.500 ;
        RECT 109.400 105.400 109.800 106.200 ;
        RECT 110.200 105.800 110.600 106.600 ;
        RECT 111.000 105.800 111.400 106.600 ;
        RECT 111.800 106.500 112.500 106.900 ;
        RECT 112.800 106.800 113.800 107.200 ;
        RECT 111.800 105.500 112.100 106.500 ;
        RECT 110.200 105.200 112.100 105.500 ;
        RECT 100.500 104.600 101.000 105.100 ;
        RECT 101.300 104.800 102.600 105.100 ;
        RECT 100.600 101.100 101.000 104.600 ;
        RECT 102.200 101.100 102.600 104.800 ;
        RECT 103.000 104.800 105.000 105.100 ;
        RECT 103.000 101.100 103.400 104.800 ;
        RECT 104.600 101.100 105.000 104.800 ;
        RECT 105.400 101.100 105.800 105.100 ;
        RECT 108.600 104.700 109.500 105.100 ;
        RECT 109.100 101.100 109.500 104.700 ;
        RECT 110.200 103.500 110.500 105.200 ;
        RECT 112.800 104.900 113.100 106.800 ;
        RECT 113.400 106.100 113.800 106.200 ;
        RECT 115.000 106.100 115.400 109.900 ;
        RECT 115.800 107.800 116.200 108.600 ;
        RECT 117.400 107.600 117.800 109.900 ;
        RECT 119.000 107.600 119.400 109.900 ;
        RECT 120.600 107.600 121.000 109.900 ;
        RECT 122.200 107.600 122.600 109.900 ;
        RECT 124.600 108.200 125.000 109.900 ;
        RECT 113.400 105.800 115.400 106.100 ;
        RECT 113.400 105.400 113.800 105.800 ;
        RECT 112.300 104.600 113.100 104.900 ;
        RECT 110.200 101.500 110.600 103.500 ;
        RECT 112.300 101.100 112.700 104.600 ;
        RECT 115.000 101.100 115.400 105.800 ;
        RECT 116.600 107.200 117.800 107.600 ;
        RECT 118.300 107.200 119.400 107.600 ;
        RECT 119.900 107.200 121.000 107.600 ;
        RECT 121.700 107.200 122.600 107.600 ;
        RECT 124.500 107.900 125.000 108.200 ;
        RECT 124.500 107.200 124.800 107.900 ;
        RECT 126.200 107.600 126.600 109.900 ;
        RECT 127.300 109.200 127.700 109.900 ;
        RECT 127.000 108.800 127.700 109.200 ;
        RECT 127.300 108.200 127.700 108.800 ;
        RECT 129.400 108.500 129.800 109.500 ;
        RECT 127.300 107.900 128.200 108.200 ;
        RECT 125.300 107.300 126.600 107.600 ;
        RECT 116.600 105.800 117.000 107.200 ;
        RECT 118.300 106.900 118.700 107.200 ;
        RECT 119.900 106.900 120.300 107.200 ;
        RECT 121.700 106.900 122.100 107.200 ;
        RECT 123.000 106.900 123.400 107.200 ;
        RECT 117.400 106.500 118.700 106.900 ;
        RECT 119.100 106.500 120.300 106.900 ;
        RECT 120.800 106.500 122.100 106.900 ;
        RECT 122.500 106.500 123.400 106.900 ;
        RECT 124.500 106.800 125.000 107.200 ;
        RECT 118.300 105.800 118.700 106.500 ;
        RECT 119.900 105.800 120.300 106.500 ;
        RECT 121.700 105.800 122.100 106.500 ;
        RECT 116.600 105.400 117.800 105.800 ;
        RECT 118.300 105.400 119.400 105.800 ;
        RECT 119.900 105.400 121.000 105.800 ;
        RECT 121.700 105.400 122.600 105.800 ;
        RECT 117.400 101.100 117.800 105.400 ;
        RECT 119.000 101.100 119.400 105.400 ;
        RECT 120.600 101.100 121.000 105.400 ;
        RECT 122.200 101.100 122.600 105.400 ;
        RECT 124.500 105.100 124.800 106.800 ;
        RECT 125.300 106.500 125.600 107.300 ;
        RECT 125.100 106.100 125.600 106.500 ;
        RECT 125.300 105.100 125.600 106.100 ;
        RECT 126.100 106.200 126.500 106.600 ;
        RECT 126.100 105.800 126.600 106.200 ;
        RECT 124.500 104.600 125.000 105.100 ;
        RECT 125.300 104.800 126.600 105.100 ;
        RECT 124.600 101.100 125.000 104.600 ;
        RECT 126.200 101.100 126.600 104.800 ;
        RECT 127.000 104.400 127.400 105.200 ;
        RECT 127.800 101.100 128.200 107.900 ;
        RECT 128.600 106.800 129.000 107.600 ;
        RECT 129.400 107.400 129.700 108.500 ;
        RECT 131.500 108.000 131.900 109.500 ;
        RECT 134.200 108.500 134.600 109.500 ;
        RECT 131.500 107.700 132.300 108.000 ;
        RECT 131.900 107.500 132.300 107.700 ;
        RECT 129.400 107.100 131.500 107.400 ;
        RECT 131.000 106.900 131.500 107.100 ;
        RECT 132.000 107.200 132.300 107.500 ;
        RECT 134.200 107.400 134.500 108.500 ;
        RECT 136.300 108.000 136.700 109.500 ;
        RECT 136.300 107.700 137.100 108.000 ;
        RECT 136.700 107.500 137.100 107.700 ;
        RECT 129.400 105.800 129.800 106.600 ;
        RECT 130.200 105.800 130.600 106.600 ;
        RECT 131.000 106.500 131.700 106.900 ;
        RECT 132.000 106.800 133.000 107.200 ;
        RECT 134.200 107.100 136.300 107.400 ;
        RECT 135.800 106.900 136.300 107.100 ;
        RECT 136.800 107.200 137.100 107.500 ;
        RECT 139.800 107.600 140.200 109.900 ;
        RECT 141.400 107.600 141.800 109.900 ;
        RECT 143.800 108.800 144.200 109.900 ;
        RECT 143.000 107.800 143.400 108.600 ;
        RECT 139.800 107.200 141.800 107.600 ;
        RECT 136.800 107.100 137.800 107.200 ;
        RECT 138.200 107.100 138.600 107.200 ;
        RECT 131.000 105.500 131.300 106.500 ;
        RECT 129.400 105.200 131.300 105.500 ;
        RECT 132.000 105.200 132.300 106.800 ;
        RECT 132.600 105.400 133.000 106.200 ;
        RECT 134.200 105.800 134.600 106.600 ;
        RECT 135.000 105.800 135.400 106.600 ;
        RECT 135.800 106.500 136.500 106.900 ;
        RECT 136.800 106.800 138.600 107.100 ;
        RECT 135.800 105.500 136.100 106.500 ;
        RECT 129.400 103.500 129.700 105.200 ;
        RECT 131.800 104.900 132.300 105.200 ;
        RECT 131.500 104.600 132.300 104.900 ;
        RECT 134.200 105.200 136.100 105.500 ;
        RECT 129.400 101.500 129.800 103.500 ;
        RECT 131.500 101.100 131.900 104.600 ;
        RECT 134.200 103.500 134.500 105.200 ;
        RECT 136.800 104.900 137.100 106.800 ;
        RECT 137.400 105.400 137.800 106.200 ;
        RECT 139.800 105.800 140.200 107.200 ;
        RECT 142.200 107.100 142.600 107.600 ;
        RECT 143.000 107.200 143.300 107.800 ;
        RECT 143.900 107.200 144.200 108.800 ;
        RECT 143.000 107.100 143.400 107.200 ;
        RECT 142.200 106.800 143.400 107.100 ;
        RECT 143.800 106.800 144.200 107.200 ;
        RECT 139.800 105.400 141.800 105.800 ;
        RECT 136.300 104.600 137.100 104.900 ;
        RECT 134.200 101.500 134.600 103.500 ;
        RECT 136.300 101.100 136.700 104.600 ;
        RECT 139.800 101.100 140.200 105.400 ;
        RECT 141.400 101.100 141.800 105.400 ;
        RECT 143.900 105.100 144.200 106.800 ;
        RECT 145.400 107.900 145.800 109.900 ;
        RECT 147.000 108.900 147.400 109.900 ;
        RECT 149.400 108.900 149.800 109.900 ;
        RECT 145.400 106.200 145.700 107.900 ;
        RECT 147.000 107.800 147.300 108.900 ;
        RECT 147.800 108.100 148.200 108.600 ;
        RECT 148.600 108.100 149.000 108.200 ;
        RECT 147.800 107.800 149.000 108.100 ;
        RECT 146.100 107.500 147.300 107.800 ;
        RECT 144.600 105.400 145.000 106.200 ;
        RECT 145.400 105.800 145.800 106.200 ;
        RECT 146.100 106.000 146.400 107.500 ;
        RECT 149.400 107.200 149.700 108.900 ;
        RECT 150.200 107.800 150.600 108.600 ;
        RECT 151.000 107.600 151.400 109.900 ;
        RECT 152.600 108.200 153.000 109.900 ;
        RECT 152.600 107.900 153.100 108.200 ;
        RECT 156.100 108.000 156.500 109.500 ;
        RECT 158.200 108.500 158.600 109.500 ;
        RECT 151.000 107.300 152.300 107.600 ;
        RECT 146.900 106.800 147.400 107.200 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 146.800 106.400 147.200 106.800 ;
        RECT 145.400 105.200 145.700 105.800 ;
        RECT 146.100 105.700 146.500 106.000 ;
        RECT 146.100 105.600 148.200 105.700 ;
        RECT 146.200 105.400 148.200 105.600 ;
        RECT 148.600 105.400 149.000 106.200 ;
        RECT 145.400 105.100 145.800 105.200 ;
        RECT 143.800 104.700 144.700 105.100 ;
        RECT 145.400 104.800 146.100 105.100 ;
        RECT 144.300 101.100 144.700 104.700 ;
        RECT 145.700 101.100 146.100 104.800 ;
        RECT 147.800 101.100 148.200 105.400 ;
        RECT 149.400 105.100 149.700 106.800 ;
        RECT 151.100 106.200 151.500 106.600 ;
        RECT 150.200 106.100 150.600 106.200 ;
        RECT 151.000 106.100 151.500 106.200 ;
        RECT 150.200 105.800 151.500 106.100 ;
        RECT 152.000 106.500 152.300 107.300 ;
        RECT 152.800 107.200 153.100 107.900 ;
        RECT 155.700 107.700 156.500 108.000 ;
        RECT 155.700 107.500 156.100 107.700 ;
        RECT 155.700 107.200 156.000 107.500 ;
        RECT 158.300 107.400 158.600 108.500 ;
        RECT 162.100 107.900 162.900 109.900 ;
        RECT 165.900 109.200 166.300 109.900 ;
        RECT 165.900 108.800 166.600 109.200 ;
        RECT 165.900 108.200 166.300 108.800 ;
        RECT 165.400 107.900 166.300 108.200 ;
        RECT 168.500 107.900 169.300 109.900 ;
        RECT 152.600 106.800 153.100 107.200 ;
        RECT 155.000 106.800 156.000 107.200 ;
        RECT 156.500 107.100 158.600 107.400 ;
        RECT 156.500 106.900 157.000 107.100 ;
        RECT 152.000 106.100 152.500 106.500 ;
        RECT 152.000 105.100 152.300 106.100 ;
        RECT 152.800 105.100 153.100 106.800 ;
        RECT 155.700 106.200 156.000 106.800 ;
        RECT 156.300 106.500 157.000 106.900 ;
        RECT 154.200 106.100 154.600 106.200 ;
        RECT 155.000 106.100 155.400 106.200 ;
        RECT 154.200 105.800 155.400 106.100 ;
        RECT 155.000 105.400 155.400 105.800 ;
        RECT 155.700 105.800 156.200 106.200 ;
        RECT 148.900 104.700 149.800 105.100 ;
        RECT 151.000 104.800 152.300 105.100 ;
        RECT 148.900 102.200 149.300 104.700 ;
        RECT 148.600 101.800 149.300 102.200 ;
        RECT 148.900 101.100 149.300 101.800 ;
        RECT 151.000 101.100 151.400 104.800 ;
        RECT 152.600 104.600 153.100 105.100 ;
        RECT 155.700 104.900 156.000 105.800 ;
        RECT 156.700 105.500 157.000 106.500 ;
        RECT 157.400 105.800 157.800 106.600 ;
        RECT 158.200 106.100 158.600 106.600 ;
        RECT 161.400 106.400 161.800 107.200 ;
        RECT 162.300 106.200 162.600 107.900 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 164.600 106.800 165.000 107.600 ;
        RECT 163.000 106.600 163.300 106.800 ;
        RECT 162.900 106.200 163.300 106.600 ;
        RECT 159.000 106.100 159.400 106.200 ;
        RECT 158.200 105.800 159.400 106.100 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 160.600 105.800 161.400 106.100 ;
        RECT 162.200 105.800 162.600 106.200 ;
        RECT 161.000 105.600 161.400 105.800 ;
        RECT 162.300 105.700 162.600 105.800 ;
        RECT 156.700 105.200 158.600 105.500 ;
        RECT 162.300 105.400 163.300 105.700 ;
        RECT 163.800 105.400 164.200 106.200 ;
        RECT 155.700 104.600 156.500 104.900 ;
        RECT 152.600 101.100 153.000 104.600 ;
        RECT 156.100 101.100 156.500 104.600 ;
        RECT 158.300 103.500 158.600 105.200 ;
        RECT 163.000 105.200 163.300 105.400 ;
        RECT 158.200 101.500 158.600 103.500 ;
        RECT 160.600 104.800 162.600 105.100 ;
        RECT 160.600 101.100 161.000 104.800 ;
        RECT 162.200 101.400 162.600 104.800 ;
        RECT 163.000 101.700 163.400 105.200 ;
        RECT 163.800 101.400 164.200 105.100 ;
        RECT 162.200 101.100 164.200 101.400 ;
        RECT 165.400 101.100 165.800 107.900 ;
        RECT 167.800 106.400 168.200 107.200 ;
        RECT 168.700 106.200 169.000 107.900 ;
        RECT 171.000 107.700 171.400 109.900 ;
        RECT 173.100 109.200 173.700 109.900 ;
        RECT 173.100 108.900 173.800 109.200 ;
        RECT 175.400 108.900 175.800 109.900 ;
        RECT 177.600 109.200 178.000 109.900 ;
        RECT 177.600 108.900 178.600 109.200 ;
        RECT 173.400 108.500 173.800 108.900 ;
        RECT 175.500 108.600 175.800 108.900 ;
        RECT 175.500 108.300 176.900 108.600 ;
        RECT 176.500 108.200 176.900 108.300 ;
        RECT 177.400 108.200 177.800 108.600 ;
        RECT 178.200 108.500 178.600 108.900 ;
        RECT 172.500 107.700 172.900 107.800 ;
        RECT 171.000 107.400 172.900 107.700 ;
        RECT 169.400 106.800 169.800 107.200 ;
        RECT 169.400 106.600 169.700 106.800 ;
        RECT 169.300 106.200 169.700 106.600 ;
        RECT 167.000 106.100 167.400 106.200 ;
        RECT 167.000 105.800 167.800 106.100 ;
        RECT 168.600 105.800 169.000 106.200 ;
        RECT 167.400 105.600 167.800 105.800 ;
        RECT 168.700 105.700 169.000 105.800 ;
        RECT 168.700 105.400 169.700 105.700 ;
        RECT 170.200 105.400 170.600 106.200 ;
        RECT 171.000 105.700 171.400 107.400 ;
        RECT 174.500 107.100 174.900 107.200 ;
        RECT 177.400 107.100 177.700 108.200 ;
        RECT 179.800 107.500 180.200 109.900 ;
        RECT 181.900 108.200 182.300 109.900 ;
        RECT 181.400 107.900 182.300 108.200 ;
        RECT 183.000 107.900 183.400 109.900 ;
        RECT 183.800 108.000 184.200 109.900 ;
        RECT 185.400 108.000 185.800 109.900 ;
        RECT 183.800 107.900 185.800 108.000 ;
        RECT 187.800 107.900 188.200 109.900 ;
        RECT 190.200 108.900 190.600 109.900 ;
        RECT 188.500 108.200 188.900 108.600 ;
        RECT 188.600 108.100 189.000 108.200 ;
        RECT 190.200 108.100 190.500 108.900 ;
        RECT 179.000 107.100 179.800 107.200 ;
        RECT 174.300 106.800 179.800 107.100 ;
        RECT 180.600 106.800 181.000 107.600 ;
        RECT 173.400 106.400 173.800 106.500 ;
        RECT 171.900 106.100 173.800 106.400 ;
        RECT 171.900 106.000 172.300 106.100 ;
        RECT 172.700 105.700 173.100 105.800 ;
        RECT 171.000 105.400 173.100 105.700 ;
        RECT 166.200 104.400 166.600 105.200 ;
        RECT 169.400 105.100 169.700 105.400 ;
        RECT 167.000 104.800 169.000 105.100 ;
        RECT 167.000 101.100 167.400 104.800 ;
        RECT 168.600 101.400 169.000 104.800 ;
        RECT 169.400 101.700 169.800 105.100 ;
        RECT 170.200 101.400 170.600 105.100 ;
        RECT 168.600 101.100 170.600 101.400 ;
        RECT 171.000 101.100 171.400 105.400 ;
        RECT 174.300 105.200 174.600 106.800 ;
        RECT 177.900 106.700 178.300 106.800 ;
        RECT 177.400 106.200 177.800 106.300 ;
        RECT 178.700 106.200 179.100 106.300 ;
        RECT 176.600 105.900 179.100 106.200 ;
        RECT 181.400 106.100 181.800 107.900 ;
        RECT 183.100 107.200 183.400 107.900 ;
        RECT 183.900 107.700 185.700 107.900 ;
        RECT 185.000 107.200 185.400 107.400 ;
        RECT 183.000 106.800 184.300 107.200 ;
        RECT 185.000 107.100 185.800 107.200 ;
        RECT 185.000 106.900 186.500 107.100 ;
        RECT 185.400 106.800 186.500 106.900 ;
        RECT 176.600 105.800 177.000 105.900 ;
        RECT 181.400 105.800 183.300 106.100 ;
        RECT 177.400 105.500 180.200 105.600 ;
        RECT 177.300 105.400 180.200 105.500 ;
        RECT 173.400 104.900 174.600 105.200 ;
        RECT 175.300 105.300 180.200 105.400 ;
        RECT 175.300 105.100 177.700 105.300 ;
        RECT 173.400 104.400 173.700 104.900 ;
        RECT 173.000 104.000 173.700 104.400 ;
        RECT 174.500 104.500 174.900 104.600 ;
        RECT 175.300 104.500 175.600 105.100 ;
        RECT 174.500 104.200 175.600 104.500 ;
        RECT 175.900 104.500 178.600 104.800 ;
        RECT 175.900 104.400 176.300 104.500 ;
        RECT 178.200 104.400 178.600 104.500 ;
        RECT 175.100 103.700 175.500 103.800 ;
        RECT 176.500 103.700 176.900 103.800 ;
        RECT 173.400 103.100 173.800 103.500 ;
        RECT 175.100 103.400 176.900 103.700 ;
        RECT 175.500 103.100 175.800 103.400 ;
        RECT 178.200 103.100 178.600 103.500 ;
        RECT 173.100 101.100 173.700 103.100 ;
        RECT 175.400 101.100 175.800 103.100 ;
        RECT 177.600 102.800 178.600 103.100 ;
        RECT 177.600 101.100 178.000 102.800 ;
        RECT 179.800 101.100 180.200 105.300 ;
        RECT 181.400 101.100 181.800 105.800 ;
        RECT 183.000 105.200 183.300 105.800 ;
        RECT 182.200 104.400 182.600 105.200 ;
        RECT 183.000 105.100 183.400 105.200 ;
        RECT 184.000 105.100 184.300 106.800 ;
        RECT 184.600 105.800 185.000 106.600 ;
        RECT 186.200 106.200 186.500 106.800 ;
        RECT 187.000 106.400 187.400 107.200 ;
        RECT 186.200 106.100 186.600 106.200 ;
        RECT 187.800 106.100 188.100 107.900 ;
        RECT 188.600 107.800 190.500 108.100 ;
        RECT 191.000 108.100 191.400 108.600 ;
        RECT 191.800 108.100 192.200 109.900 ;
        RECT 193.900 109.200 194.500 109.900 ;
        RECT 193.900 108.900 194.600 109.200 ;
        RECT 196.200 108.900 196.600 109.900 ;
        RECT 198.400 109.200 198.800 109.900 ;
        RECT 198.400 108.900 199.400 109.200 ;
        RECT 194.200 108.500 194.600 108.900 ;
        RECT 196.300 108.600 196.600 108.900 ;
        RECT 196.300 108.300 197.700 108.600 ;
        RECT 197.300 108.200 197.700 108.300 ;
        RECT 198.200 108.200 198.600 108.600 ;
        RECT 199.000 108.500 199.400 108.900 ;
        RECT 191.000 107.800 192.200 108.100 ;
        RECT 190.200 107.200 190.500 107.800 ;
        RECT 191.800 107.700 192.200 107.800 ;
        RECT 193.300 107.700 193.700 107.800 ;
        RECT 191.800 107.400 193.700 107.700 ;
        RECT 188.600 106.800 189.000 107.200 ;
        RECT 190.200 106.800 190.600 107.200 ;
        RECT 188.600 106.200 188.900 106.800 ;
        RECT 188.600 106.100 189.000 106.200 ;
        RECT 186.200 105.800 187.000 106.100 ;
        RECT 187.800 105.800 189.000 106.100 ;
        RECT 186.600 105.600 187.000 105.800 ;
        RECT 188.600 105.100 188.900 105.800 ;
        RECT 189.400 105.400 189.800 106.200 ;
        RECT 190.200 105.100 190.500 106.800 ;
        RECT 191.800 105.700 192.200 107.400 ;
        RECT 195.300 107.100 195.700 107.200 ;
        RECT 198.200 107.100 198.500 108.200 ;
        RECT 200.600 107.500 201.000 109.900 ;
        RECT 201.400 107.600 201.800 109.900 ;
        RECT 203.000 108.200 203.400 109.900 ;
        RECT 205.900 109.200 206.300 109.900 ;
        RECT 205.400 108.800 206.300 109.200 ;
        RECT 207.800 108.900 208.200 109.900 ;
        RECT 211.800 108.900 212.200 109.900 ;
        RECT 205.900 108.200 206.300 108.800 ;
        RECT 203.000 107.900 203.500 108.200 ;
        RECT 201.400 107.300 202.700 107.600 ;
        RECT 199.800 107.100 200.600 107.200 ;
        RECT 195.100 106.800 200.600 107.100 ;
        RECT 194.200 106.400 194.600 106.500 ;
        RECT 192.700 106.100 194.600 106.400 ;
        RECT 192.700 106.000 193.100 106.100 ;
        RECT 193.500 105.700 193.900 105.800 ;
        RECT 191.800 105.400 193.900 105.700 ;
        RECT 183.000 104.800 183.700 105.100 ;
        RECT 184.000 104.800 184.500 105.100 ;
        RECT 183.400 104.200 183.700 104.800 ;
        RECT 183.400 103.800 183.800 104.200 ;
        RECT 184.100 101.100 184.500 104.800 ;
        RECT 186.200 104.800 188.200 105.100 ;
        RECT 186.200 101.100 186.600 104.800 ;
        RECT 187.800 101.100 188.200 104.800 ;
        RECT 188.600 101.100 189.000 105.100 ;
        RECT 189.700 104.700 190.600 105.100 ;
        RECT 189.700 101.100 190.100 104.700 ;
        RECT 191.800 101.100 192.200 105.400 ;
        RECT 195.100 105.200 195.400 106.800 ;
        RECT 198.700 106.700 199.100 106.800 ;
        RECT 199.500 106.200 199.900 106.300 ;
        RECT 201.500 106.200 201.900 106.600 ;
        RECT 197.400 105.900 199.900 106.200 ;
        RECT 197.400 105.800 197.800 105.900 ;
        RECT 201.400 105.800 201.900 106.200 ;
        RECT 202.400 106.500 202.700 107.300 ;
        RECT 203.200 107.200 203.500 107.900 ;
        RECT 205.400 107.900 206.300 108.200 ;
        RECT 203.000 106.800 203.500 107.200 ;
        RECT 204.600 106.800 205.000 107.600 ;
        RECT 202.400 106.100 202.900 106.500 ;
        RECT 198.200 105.500 201.000 105.600 ;
        RECT 198.100 105.400 201.000 105.500 ;
        RECT 194.200 104.900 195.400 105.200 ;
        RECT 196.100 105.300 201.000 105.400 ;
        RECT 196.100 105.100 198.500 105.300 ;
        RECT 194.200 104.400 194.500 104.900 ;
        RECT 193.800 104.000 194.500 104.400 ;
        RECT 195.300 104.500 195.700 104.600 ;
        RECT 196.100 104.500 196.400 105.100 ;
        RECT 195.300 104.200 196.400 104.500 ;
        RECT 196.700 104.500 199.400 104.800 ;
        RECT 196.700 104.400 197.100 104.500 ;
        RECT 199.000 104.400 199.400 104.500 ;
        RECT 195.900 103.700 196.300 103.800 ;
        RECT 197.300 103.700 197.700 103.800 ;
        RECT 194.200 103.100 194.600 103.500 ;
        RECT 195.900 103.400 197.700 103.700 ;
        RECT 196.300 103.100 196.600 103.400 ;
        RECT 199.000 103.100 199.400 103.500 ;
        RECT 193.900 101.100 194.500 103.100 ;
        RECT 196.200 101.100 196.600 103.100 ;
        RECT 198.400 102.800 199.400 103.100 ;
        RECT 198.400 101.100 198.800 102.800 ;
        RECT 200.600 101.100 201.000 105.300 ;
        RECT 202.400 105.100 202.700 106.100 ;
        RECT 203.200 105.100 203.500 106.800 ;
        RECT 201.400 104.800 202.700 105.100 ;
        RECT 201.400 101.100 201.800 104.800 ;
        RECT 203.000 104.600 203.500 105.100 ;
        RECT 203.000 101.100 203.400 104.600 ;
        RECT 205.400 101.100 205.800 107.900 ;
        RECT 207.000 107.800 207.400 108.600 ;
        RECT 207.900 107.200 208.200 108.900 ;
        RECT 210.200 108.100 210.600 108.200 ;
        RECT 211.000 108.100 211.400 108.600 ;
        RECT 210.200 107.800 211.400 108.100 ;
        RECT 211.900 107.200 212.200 108.900 ;
        RECT 213.400 107.700 213.800 109.900 ;
        RECT 215.500 109.200 216.100 109.900 ;
        RECT 215.500 108.900 216.200 109.200 ;
        RECT 217.800 108.900 218.200 109.900 ;
        RECT 220.000 109.200 220.400 109.900 ;
        RECT 220.000 108.900 221.000 109.200 ;
        RECT 215.800 108.500 216.200 108.900 ;
        RECT 217.900 108.600 218.200 108.900 ;
        RECT 217.900 108.300 219.300 108.600 ;
        RECT 218.900 108.200 219.300 108.300 ;
        RECT 219.800 108.200 220.200 108.600 ;
        RECT 220.600 108.500 221.000 108.900 ;
        RECT 214.900 107.700 215.300 107.800 ;
        RECT 213.400 107.400 215.300 107.700 ;
        RECT 207.800 106.800 208.200 107.200 ;
        RECT 211.800 106.800 212.200 107.200 ;
        RECT 206.200 105.800 206.600 106.200 ;
        RECT 206.200 105.200 206.500 105.800 ;
        RECT 206.200 104.400 206.600 105.200 ;
        RECT 207.900 105.100 208.200 106.800 ;
        RECT 208.600 105.400 209.000 106.200 ;
        RECT 211.900 105.100 212.200 106.800 ;
        RECT 212.600 106.800 213.000 107.200 ;
        RECT 212.600 106.200 212.900 106.800 ;
        RECT 212.600 105.400 213.000 106.200 ;
        RECT 213.400 105.700 213.800 107.400 ;
        RECT 216.900 107.100 217.300 107.200 ;
        RECT 218.200 107.100 218.600 107.200 ;
        RECT 219.800 107.100 220.100 108.200 ;
        RECT 222.200 107.500 222.600 109.900 ;
        RECT 223.300 109.200 223.700 109.900 ;
        RECT 223.000 108.800 223.700 109.200 ;
        RECT 226.200 108.900 226.600 109.900 ;
        RECT 223.300 108.200 223.700 108.800 ;
        RECT 223.300 107.900 224.200 108.200 ;
        RECT 221.400 107.100 222.200 107.200 ;
        RECT 216.700 106.800 222.200 107.100 ;
        RECT 215.800 106.400 216.200 106.500 ;
        RECT 214.300 106.100 216.200 106.400 ;
        RECT 214.300 106.000 214.700 106.100 ;
        RECT 215.100 105.700 215.500 105.800 ;
        RECT 213.400 105.400 215.500 105.700 ;
        RECT 207.800 104.700 208.700 105.100 ;
        RECT 211.800 104.700 212.700 105.100 ;
        RECT 208.300 102.200 208.700 104.700 ;
        RECT 212.300 102.200 212.700 104.700 ;
        RECT 208.300 101.800 209.000 102.200 ;
        RECT 211.800 101.800 212.700 102.200 ;
        RECT 208.300 101.100 208.700 101.800 ;
        RECT 212.300 101.100 212.700 101.800 ;
        RECT 213.400 101.100 213.800 105.400 ;
        RECT 216.700 105.200 217.000 106.800 ;
        RECT 220.300 106.700 220.700 106.800 ;
        RECT 221.100 106.200 221.500 106.300 ;
        RECT 217.400 106.100 217.800 106.200 ;
        RECT 219.000 106.100 221.500 106.200 ;
        RECT 217.400 105.900 221.500 106.100 ;
        RECT 217.400 105.800 219.400 105.900 ;
        RECT 219.800 105.500 222.600 105.600 ;
        RECT 219.700 105.400 222.600 105.500 ;
        RECT 215.800 104.900 217.000 105.200 ;
        RECT 217.700 105.300 222.600 105.400 ;
        RECT 217.700 105.100 220.100 105.300 ;
        RECT 215.800 104.400 216.100 104.900 ;
        RECT 215.400 104.000 216.100 104.400 ;
        RECT 216.900 104.500 217.300 104.600 ;
        RECT 217.700 104.500 218.000 105.100 ;
        RECT 216.900 104.200 218.000 104.500 ;
        RECT 218.300 104.500 221.000 104.800 ;
        RECT 218.300 104.400 218.700 104.500 ;
        RECT 220.600 104.400 221.000 104.500 ;
        RECT 217.500 103.700 217.900 103.800 ;
        RECT 218.900 103.700 219.300 103.800 ;
        RECT 215.800 103.100 216.200 103.500 ;
        RECT 217.500 103.400 219.300 103.700 ;
        RECT 217.900 103.100 218.200 103.400 ;
        RECT 220.600 103.100 221.000 103.500 ;
        RECT 215.500 101.100 216.100 103.100 ;
        RECT 217.800 101.100 218.200 103.100 ;
        RECT 220.000 102.800 221.000 103.100 ;
        RECT 220.000 101.100 220.400 102.800 ;
        RECT 222.200 101.100 222.600 105.300 ;
        RECT 223.000 104.400 223.400 105.200 ;
        RECT 223.800 101.100 224.200 107.900 ;
        RECT 225.400 107.800 225.800 108.600 ;
        RECT 224.600 107.100 225.000 107.600 ;
        RECT 225.400 107.100 225.700 107.800 ;
        RECT 226.300 107.200 226.600 108.900 ;
        RECT 229.100 108.200 229.500 109.900 ;
        RECT 231.500 109.200 231.900 109.900 ;
        RECT 231.000 108.800 231.900 109.200 ;
        RECT 231.500 108.200 231.900 108.800 ;
        RECT 228.600 107.900 229.500 108.200 ;
        RECT 231.000 107.900 231.900 108.200 ;
        RECT 224.600 106.800 225.700 107.100 ;
        RECT 226.200 106.800 226.600 107.200 ;
        RECT 227.800 106.800 228.200 107.600 ;
        RECT 226.300 105.200 226.600 106.800 ;
        RECT 227.000 105.400 227.400 106.200 ;
        RECT 226.200 105.100 226.600 105.200 ;
        RECT 226.200 104.700 227.100 105.100 ;
        RECT 226.700 101.100 227.100 104.700 ;
        RECT 228.600 101.100 229.000 107.900 ;
        RECT 230.200 106.800 230.600 107.600 ;
        RECT 229.400 104.400 229.800 105.200 ;
        RECT 231.000 101.100 231.400 107.900 ;
        RECT 232.600 107.700 233.000 109.900 ;
        RECT 234.700 109.200 235.300 109.900 ;
        RECT 234.700 108.900 235.400 109.200 ;
        RECT 237.000 108.900 237.400 109.900 ;
        RECT 239.200 109.200 239.600 109.900 ;
        RECT 239.200 108.900 240.200 109.200 ;
        RECT 235.000 108.500 235.400 108.900 ;
        RECT 237.100 108.600 237.400 108.900 ;
        RECT 237.100 108.300 238.500 108.600 ;
        RECT 238.100 108.200 238.500 108.300 ;
        RECT 239.000 108.200 239.400 108.600 ;
        RECT 239.800 108.500 240.200 108.900 ;
        RECT 234.100 107.700 234.500 107.800 ;
        RECT 232.600 107.400 234.500 107.700 ;
        RECT 232.600 105.700 233.000 107.400 ;
        RECT 236.100 107.100 236.500 107.200 ;
        RECT 238.200 107.100 238.600 107.200 ;
        RECT 239.000 107.100 239.300 108.200 ;
        RECT 241.400 107.500 241.800 109.900 ;
        RECT 243.800 107.900 244.200 109.900 ;
        RECT 244.500 108.200 244.900 108.600 ;
        RECT 240.600 107.100 241.400 107.200 ;
        RECT 235.900 106.800 241.400 107.100 ;
        RECT 235.000 106.400 235.400 106.500 ;
        RECT 233.500 106.100 235.400 106.400 ;
        RECT 233.500 106.000 233.900 106.100 ;
        RECT 234.300 105.700 234.700 105.800 ;
        RECT 232.600 105.400 234.700 105.700 ;
        RECT 231.800 104.400 232.200 105.200 ;
        RECT 232.600 101.100 233.000 105.400 ;
        RECT 235.900 105.200 236.200 106.800 ;
        RECT 239.500 106.700 239.900 106.800 ;
        RECT 243.000 106.400 243.400 107.200 ;
        RECT 239.000 106.200 239.400 106.300 ;
        RECT 240.300 106.200 240.700 106.300 ;
        RECT 238.200 105.900 240.700 106.200 ;
        RECT 243.800 106.200 244.100 107.900 ;
        RECT 244.600 107.800 245.000 108.200 ;
        RECT 246.200 107.600 246.600 109.900 ;
        RECT 247.800 107.600 248.200 109.900 ;
        RECT 249.400 107.600 249.800 109.900 ;
        RECT 251.000 107.600 251.400 109.900 ;
        RECT 245.400 107.200 246.600 107.600 ;
        RECT 247.100 107.200 248.200 107.600 ;
        RECT 248.700 107.200 249.800 107.600 ;
        RECT 250.500 107.200 251.400 107.600 ;
        RECT 252.600 107.500 253.000 109.900 ;
        RECT 254.800 109.200 255.200 109.900 ;
        RECT 254.200 108.900 255.200 109.200 ;
        RECT 257.000 108.900 257.400 109.900 ;
        RECT 259.100 109.200 259.700 109.900 ;
        RECT 259.000 108.900 259.700 109.200 ;
        RECT 254.200 108.500 254.600 108.900 ;
        RECT 257.000 108.600 257.300 108.900 ;
        RECT 255.000 108.200 255.400 108.600 ;
        RECT 255.900 108.300 257.300 108.600 ;
        RECT 259.000 108.500 259.400 108.900 ;
        RECT 255.900 108.200 256.300 108.300 ;
        RECT 243.800 106.100 244.200 106.200 ;
        RECT 244.600 106.100 245.000 106.200 ;
        RECT 238.200 105.800 238.600 105.900 ;
        RECT 243.800 105.800 245.000 106.100 ;
        RECT 245.400 105.800 245.800 107.200 ;
        RECT 247.100 106.900 247.500 107.200 ;
        RECT 248.700 106.900 249.100 107.200 ;
        RECT 250.500 106.900 250.900 107.200 ;
        RECT 251.800 106.900 252.200 107.200 ;
        RECT 246.200 106.500 247.500 106.900 ;
        RECT 247.900 106.500 249.100 106.900 ;
        RECT 249.600 106.500 250.900 106.900 ;
        RECT 251.300 106.500 252.200 106.900 ;
        RECT 253.000 107.100 253.800 107.200 ;
        RECT 255.100 107.100 255.400 108.200 ;
        RECT 259.900 107.700 260.300 107.800 ;
        RECT 261.400 107.700 261.800 109.900 ;
        RECT 263.000 108.900 263.400 109.900 ;
        RECT 259.900 107.400 261.800 107.700 ;
        RECT 257.900 107.100 258.300 107.200 ;
        RECT 253.000 106.800 258.500 107.100 ;
        RECT 260.600 106.800 261.000 107.400 ;
        RECT 254.500 106.700 254.900 106.800 ;
        RECT 247.100 105.800 247.500 106.500 ;
        RECT 248.700 105.800 249.100 106.500 ;
        RECT 250.500 105.800 250.900 106.500 ;
        RECT 253.700 106.200 254.100 106.300 ;
        RECT 253.700 105.900 256.200 106.200 ;
        RECT 255.800 105.800 256.200 105.900 ;
        RECT 239.000 105.500 241.800 105.600 ;
        RECT 238.900 105.400 241.800 105.500 ;
        RECT 235.000 104.900 236.200 105.200 ;
        RECT 236.900 105.300 241.800 105.400 ;
        RECT 236.900 105.100 239.300 105.300 ;
        RECT 235.000 104.400 235.300 104.900 ;
        RECT 234.600 104.000 235.300 104.400 ;
        RECT 236.100 104.500 236.500 104.600 ;
        RECT 236.900 104.500 237.200 105.100 ;
        RECT 236.100 104.200 237.200 104.500 ;
        RECT 237.500 104.500 240.200 104.800 ;
        RECT 237.500 104.400 237.900 104.500 ;
        RECT 239.800 104.400 240.200 104.500 ;
        RECT 236.700 103.700 237.100 103.800 ;
        RECT 238.100 103.700 238.500 103.800 ;
        RECT 235.000 103.100 235.400 103.500 ;
        RECT 236.700 103.400 238.500 103.700 ;
        RECT 237.100 103.100 237.400 103.400 ;
        RECT 239.800 103.100 240.200 103.500 ;
        RECT 234.700 101.100 235.300 103.100 ;
        RECT 237.000 101.100 237.400 103.100 ;
        RECT 239.200 102.800 240.200 103.100 ;
        RECT 239.200 101.100 239.600 102.800 ;
        RECT 241.400 101.100 241.800 105.300 ;
        RECT 244.600 105.100 244.900 105.800 ;
        RECT 245.400 105.400 246.600 105.800 ;
        RECT 247.100 105.400 248.200 105.800 ;
        RECT 248.700 105.400 249.800 105.800 ;
        RECT 250.500 105.400 251.400 105.800 ;
        RECT 242.200 104.800 244.200 105.100 ;
        RECT 242.200 101.100 242.600 104.800 ;
        RECT 243.800 101.100 244.200 104.800 ;
        RECT 244.600 101.100 245.000 105.100 ;
        RECT 246.200 101.100 246.600 105.400 ;
        RECT 247.800 101.100 248.200 105.400 ;
        RECT 249.400 101.100 249.800 105.400 ;
        RECT 251.000 101.100 251.400 105.400 ;
        RECT 252.600 105.500 255.400 105.600 ;
        RECT 252.600 105.400 255.500 105.500 ;
        RECT 252.600 105.300 257.500 105.400 ;
        RECT 252.600 101.100 253.000 105.300 ;
        RECT 255.100 105.100 257.500 105.300 ;
        RECT 254.200 104.500 256.900 104.800 ;
        RECT 254.200 104.400 254.600 104.500 ;
        RECT 256.500 104.400 256.900 104.500 ;
        RECT 257.200 104.500 257.500 105.100 ;
        RECT 258.200 105.200 258.500 106.800 ;
        RECT 259.000 106.400 259.400 106.500 ;
        RECT 259.000 106.100 260.900 106.400 ;
        RECT 260.500 106.000 260.900 106.100 ;
        RECT 259.700 105.700 260.100 105.800 ;
        RECT 261.400 105.700 261.800 107.400 ;
        RECT 263.100 107.200 263.400 108.900 ;
        RECT 262.200 106.800 262.600 107.200 ;
        RECT 263.000 106.800 263.400 107.200 ;
        RECT 262.200 106.100 262.500 106.800 ;
        RECT 263.100 106.100 263.400 106.800 ;
        RECT 262.200 105.800 263.400 106.100 ;
        RECT 259.700 105.400 261.800 105.700 ;
        RECT 258.200 104.900 259.400 105.200 ;
        RECT 257.900 104.500 258.300 104.600 ;
        RECT 257.200 104.200 258.300 104.500 ;
        RECT 259.100 104.400 259.400 104.900 ;
        RECT 259.100 104.000 259.800 104.400 ;
        RECT 255.900 103.700 256.300 103.800 ;
        RECT 257.300 103.700 257.700 103.800 ;
        RECT 254.200 103.100 254.600 103.500 ;
        RECT 255.900 103.400 257.700 103.700 ;
        RECT 257.000 103.100 257.300 103.400 ;
        RECT 259.000 103.100 259.400 103.500 ;
        RECT 254.200 102.800 255.200 103.100 ;
        RECT 254.800 101.100 255.200 102.800 ;
        RECT 257.000 101.100 257.400 103.100 ;
        RECT 259.100 101.100 259.700 103.100 ;
        RECT 261.400 101.100 261.800 105.400 ;
        RECT 263.100 105.100 263.400 105.800 ;
        RECT 263.000 104.700 263.900 105.100 ;
        RECT 263.500 101.100 263.900 104.700 ;
        RECT 0.600 95.700 1.000 99.900 ;
        RECT 2.800 98.200 3.200 99.900 ;
        RECT 2.200 97.900 3.200 98.200 ;
        RECT 5.000 97.900 5.400 99.900 ;
        RECT 7.100 97.900 7.700 99.900 ;
        RECT 2.200 97.500 2.600 97.900 ;
        RECT 5.000 97.600 5.300 97.900 ;
        RECT 3.900 97.300 5.700 97.600 ;
        RECT 7.000 97.500 7.400 97.900 ;
        RECT 3.900 97.200 4.300 97.300 ;
        RECT 5.300 97.200 5.700 97.300 ;
        RECT 2.200 96.500 2.600 96.600 ;
        RECT 4.500 96.500 4.900 96.600 ;
        RECT 2.200 96.200 4.900 96.500 ;
        RECT 5.200 96.500 6.300 96.800 ;
        RECT 5.200 95.900 5.500 96.500 ;
        RECT 5.900 96.400 6.300 96.500 ;
        RECT 7.100 96.600 7.800 97.000 ;
        RECT 7.100 96.100 7.400 96.600 ;
        RECT 3.100 95.700 5.500 95.900 ;
        RECT 0.600 95.600 5.500 95.700 ;
        RECT 6.200 95.800 7.400 96.100 ;
        RECT 0.600 95.500 3.500 95.600 ;
        RECT 0.600 95.400 3.400 95.500 ;
        RECT 3.800 95.100 4.200 95.200 ;
        RECT 5.400 95.100 5.800 95.200 ;
        RECT 1.700 94.800 5.800 95.100 ;
        RECT 1.700 94.700 2.100 94.800 ;
        RECT 2.500 94.200 2.900 94.300 ;
        RECT 6.200 94.200 6.500 95.800 ;
        RECT 9.400 95.600 9.800 99.900 ;
        RECT 7.700 95.300 9.800 95.600 ;
        RECT 7.700 95.200 8.100 95.300 ;
        RECT 8.500 94.900 8.900 95.000 ;
        RECT 7.000 94.600 8.900 94.900 ;
        RECT 7.000 94.500 7.400 94.600 ;
        RECT 1.000 93.900 6.500 94.200 ;
        RECT 9.400 94.100 9.800 95.300 ;
        RECT 11.000 95.100 11.400 99.900 ;
        RECT 13.000 96.800 13.400 97.200 ;
        RECT 11.800 95.800 12.200 96.600 ;
        RECT 13.000 96.200 13.300 96.800 ;
        RECT 13.700 96.200 14.100 99.900 ;
        RECT 12.600 95.900 13.300 96.200 ;
        RECT 13.600 95.900 14.100 96.200 ;
        RECT 15.800 97.500 16.200 99.500 ;
        RECT 17.900 99.200 18.300 99.900 ;
        RECT 17.900 98.800 18.600 99.200 ;
        RECT 12.600 95.800 13.000 95.900 ;
        RECT 12.600 95.100 12.900 95.800 ;
        RECT 11.000 94.800 12.900 95.100 ;
        RECT 10.200 94.100 10.600 94.200 ;
        RECT 1.000 93.800 1.800 93.900 ;
        RECT 3.000 93.800 3.400 93.900 ;
        RECT 5.900 93.800 6.300 93.900 ;
        RECT 9.400 93.800 10.600 94.100 ;
        RECT 0.600 91.100 1.000 93.500 ;
        RECT 3.100 92.800 3.400 93.800 ;
        RECT 9.400 93.600 9.800 93.800 ;
        RECT 7.900 93.300 9.800 93.600 ;
        RECT 10.200 93.400 10.600 93.800 ;
        RECT 7.900 93.200 8.300 93.300 ;
        RECT 2.200 92.100 2.600 92.500 ;
        RECT 3.000 92.400 3.400 92.800 ;
        RECT 3.900 92.700 4.300 92.800 ;
        RECT 3.900 92.400 5.300 92.700 ;
        RECT 5.000 92.100 5.300 92.400 ;
        RECT 7.000 92.100 7.400 92.500 ;
        RECT 2.200 91.800 3.200 92.100 ;
        RECT 2.800 91.100 3.200 91.800 ;
        RECT 5.000 91.100 5.400 92.100 ;
        RECT 7.000 91.800 7.700 92.100 ;
        RECT 7.100 91.100 7.700 91.800 ;
        RECT 9.400 91.100 9.800 93.300 ;
        RECT 11.000 93.100 11.400 94.800 ;
        RECT 13.600 94.200 13.900 95.900 ;
        RECT 15.800 95.800 16.100 97.500 ;
        RECT 17.900 96.400 18.300 98.800 ;
        RECT 17.900 96.100 18.700 96.400 ;
        RECT 15.800 95.500 17.700 95.800 ;
        RECT 14.200 94.400 14.600 95.200 ;
        RECT 15.800 94.400 16.200 95.200 ;
        RECT 16.600 94.400 17.000 95.200 ;
        RECT 17.400 94.500 17.700 95.500 ;
        RECT 12.600 93.800 13.900 94.200 ;
        RECT 15.000 94.100 15.400 94.200 ;
        RECT 14.600 93.800 15.400 94.100 ;
        RECT 17.400 94.100 18.100 94.500 ;
        RECT 18.400 94.200 18.700 96.100 ;
        RECT 19.000 95.100 19.400 95.600 ;
        RECT 19.000 94.800 20.100 95.100 ;
        RECT 19.800 94.200 20.100 94.800 ;
        RECT 17.400 93.900 17.900 94.100 ;
        RECT 12.700 93.100 13.000 93.800 ;
        RECT 14.600 93.600 15.000 93.800 ;
        RECT 15.800 93.600 17.900 93.900 ;
        RECT 18.400 93.800 19.400 94.200 ;
        RECT 19.800 94.100 20.200 94.200 ;
        RECT 20.600 94.100 21.000 94.200 ;
        RECT 19.800 93.800 21.000 94.100 ;
        RECT 13.500 93.100 15.300 93.300 ;
        RECT 11.000 92.800 11.900 93.100 ;
        RECT 11.500 91.100 11.900 92.800 ;
        RECT 12.600 91.100 13.000 93.100 ;
        RECT 13.400 93.000 15.400 93.100 ;
        RECT 13.400 91.100 13.800 93.000 ;
        RECT 15.000 91.100 15.400 93.000 ;
        RECT 15.800 92.500 16.100 93.600 ;
        RECT 18.400 93.500 18.700 93.800 ;
        RECT 18.300 93.300 18.700 93.500 ;
        RECT 20.600 93.400 21.000 93.800 ;
        RECT 17.900 93.000 18.700 93.300 ;
        RECT 21.400 93.100 21.800 99.900 ;
        RECT 22.200 95.800 22.600 96.600 ;
        RECT 23.000 95.700 23.400 99.900 ;
        RECT 25.200 98.200 25.600 99.900 ;
        RECT 24.600 97.900 25.600 98.200 ;
        RECT 27.400 97.900 27.800 99.900 ;
        RECT 29.500 97.900 30.100 99.900 ;
        RECT 24.600 97.500 25.000 97.900 ;
        RECT 27.400 97.600 27.700 97.900 ;
        RECT 26.300 97.300 28.100 97.600 ;
        RECT 29.400 97.500 29.800 97.900 ;
        RECT 26.300 97.200 26.700 97.300 ;
        RECT 27.700 97.200 28.100 97.300 ;
        RECT 31.800 97.100 32.200 99.900 ;
        RECT 32.600 97.100 33.000 97.200 ;
        RECT 24.600 96.500 25.000 96.600 ;
        RECT 26.900 96.500 27.300 96.600 ;
        RECT 24.600 96.200 27.300 96.500 ;
        RECT 27.600 96.500 28.700 96.800 ;
        RECT 27.600 95.900 27.900 96.500 ;
        RECT 28.300 96.400 28.700 96.500 ;
        RECT 29.500 96.600 30.200 97.000 ;
        RECT 31.800 96.800 33.000 97.100 ;
        RECT 29.500 96.100 29.800 96.600 ;
        RECT 25.500 95.700 27.900 95.900 ;
        RECT 23.000 95.600 27.900 95.700 ;
        RECT 28.600 95.800 29.800 96.100 ;
        RECT 23.000 95.500 25.900 95.600 ;
        RECT 23.000 95.400 25.800 95.500 ;
        RECT 26.200 95.100 26.600 95.200 ;
        RECT 24.100 94.800 26.600 95.100 ;
        RECT 24.100 94.700 24.500 94.800 ;
        RECT 24.900 94.200 25.300 94.300 ;
        RECT 28.600 94.200 28.900 95.800 ;
        RECT 31.800 95.600 32.200 96.800 ;
        RECT 30.100 95.300 32.200 95.600 ;
        RECT 30.100 95.200 30.500 95.300 ;
        RECT 30.900 94.900 31.300 95.000 ;
        RECT 29.400 94.600 31.300 94.900 ;
        RECT 29.400 94.500 29.800 94.600 ;
        RECT 23.400 93.900 28.900 94.200 ;
        RECT 23.400 93.800 24.200 93.900 ;
        RECT 15.800 91.500 16.200 92.500 ;
        RECT 17.900 91.500 18.300 93.000 ;
        RECT 21.400 92.800 22.300 93.100 ;
        RECT 21.900 92.200 22.300 92.800 ;
        RECT 21.400 91.800 22.300 92.200 ;
        RECT 21.900 91.100 22.300 91.800 ;
        RECT 23.000 91.100 23.400 93.500 ;
        RECT 25.500 92.800 25.800 93.900 ;
        RECT 28.300 93.800 28.700 93.900 ;
        RECT 31.800 93.600 32.200 95.300 ;
        RECT 33.400 95.100 33.800 99.900 ;
        RECT 35.400 96.800 35.800 97.200 ;
        RECT 34.200 95.800 34.600 96.600 ;
        RECT 35.400 96.200 35.700 96.800 ;
        RECT 36.100 96.200 36.500 99.900 ;
        RECT 39.500 96.300 39.900 99.900 ;
        RECT 42.500 99.200 42.900 99.900 ;
        RECT 42.500 98.800 43.400 99.200 ;
        RECT 42.500 96.400 42.900 98.800 ;
        RECT 44.600 97.500 45.000 99.500 ;
        RECT 35.000 95.900 35.700 96.200 ;
        RECT 36.000 95.900 36.500 96.200 ;
        RECT 39.000 95.900 39.900 96.300 ;
        RECT 42.100 96.100 42.900 96.400 ;
        RECT 35.000 95.800 35.400 95.900 ;
        RECT 35.000 95.100 35.300 95.800 ;
        RECT 33.400 94.800 35.300 95.100 ;
        RECT 30.300 93.300 32.200 93.600 ;
        RECT 32.600 93.400 33.000 94.200 ;
        RECT 30.300 93.200 30.700 93.300 ;
        RECT 24.600 92.100 25.000 92.500 ;
        RECT 25.400 92.400 25.800 92.800 ;
        RECT 26.300 92.700 26.700 92.800 ;
        RECT 26.300 92.400 27.700 92.700 ;
        RECT 27.400 92.100 27.700 92.400 ;
        RECT 29.400 92.100 29.800 92.500 ;
        RECT 24.600 91.800 25.600 92.100 ;
        RECT 25.200 91.100 25.600 91.800 ;
        RECT 27.400 91.100 27.800 92.100 ;
        RECT 29.400 91.800 30.100 92.100 ;
        RECT 29.500 91.100 30.100 91.800 ;
        RECT 31.800 91.100 32.200 93.300 ;
        RECT 33.400 93.100 33.800 94.800 ;
        RECT 36.000 94.200 36.300 95.900 ;
        RECT 36.600 94.400 37.000 95.200 ;
        RECT 39.100 94.200 39.400 95.900 ;
        RECT 39.800 95.100 40.200 95.600 ;
        RECT 40.600 95.100 41.000 95.200 ;
        RECT 39.800 94.800 41.000 95.100 ;
        RECT 41.400 94.800 41.800 95.600 ;
        RECT 42.100 94.200 42.400 96.100 ;
        RECT 44.700 95.800 45.000 97.500 ;
        RECT 46.700 96.200 47.100 99.900 ;
        RECT 47.400 96.800 47.800 97.200 ;
        RECT 47.500 96.200 47.800 96.800 ;
        RECT 46.700 95.900 47.200 96.200 ;
        RECT 47.500 95.900 48.200 96.200 ;
        RECT 43.100 95.500 45.000 95.800 ;
        RECT 43.100 94.500 43.400 95.500 ;
        RECT 35.000 93.800 36.300 94.200 ;
        RECT 37.400 94.100 37.800 94.200 ;
        RECT 38.200 94.100 38.600 94.200 ;
        RECT 37.000 93.800 38.600 94.100 ;
        RECT 39.000 93.800 39.400 94.200 ;
        RECT 41.400 93.800 42.400 94.200 ;
        RECT 42.700 94.100 43.400 94.500 ;
        RECT 43.800 94.400 44.200 95.200 ;
        RECT 44.600 94.400 45.000 95.200 ;
        RECT 46.200 94.400 46.600 95.200 ;
        RECT 46.900 94.200 47.200 95.900 ;
        RECT 47.800 95.800 48.200 95.900 ;
        RECT 48.600 95.800 49.000 96.600 ;
        RECT 47.800 95.100 48.100 95.800 ;
        RECT 49.400 95.100 49.800 99.900 ;
        RECT 47.800 94.800 49.800 95.100 ;
        RECT 35.100 93.100 35.400 93.800 ;
        RECT 37.000 93.600 37.400 93.800 ;
        RECT 35.900 93.100 37.700 93.300 ;
        RECT 33.400 92.800 34.300 93.100 ;
        RECT 33.900 91.100 34.300 92.800 ;
        RECT 35.000 91.100 35.400 93.100 ;
        RECT 35.800 93.000 37.800 93.100 ;
        RECT 35.800 91.100 36.200 93.000 ;
        RECT 37.400 91.100 37.800 93.000 ;
        RECT 38.200 92.400 38.600 93.200 ;
        RECT 39.100 92.200 39.400 93.800 ;
        RECT 42.100 93.500 42.400 93.800 ;
        RECT 42.900 93.900 43.400 94.100 ;
        RECT 45.400 94.100 45.800 94.200 ;
        RECT 46.900 94.100 48.200 94.200 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 42.900 93.600 45.000 93.900 ;
        RECT 45.400 93.800 46.200 94.100 ;
        RECT 46.900 93.800 49.000 94.100 ;
        RECT 45.800 93.600 46.200 93.800 ;
        RECT 42.100 93.300 42.500 93.500 ;
        RECT 42.100 93.000 42.900 93.300 ;
        RECT 39.000 91.100 39.400 92.200 ;
        RECT 42.500 91.500 42.900 93.000 ;
        RECT 44.700 92.500 45.000 93.600 ;
        RECT 45.500 93.100 47.300 93.300 ;
        RECT 47.800 93.100 48.100 93.800 ;
        RECT 49.400 93.100 49.800 94.800 ;
        RECT 52.600 95.600 53.000 99.900 ;
        RECT 54.700 97.900 55.300 99.900 ;
        RECT 57.000 97.900 57.400 99.900 ;
        RECT 59.200 98.200 59.600 99.900 ;
        RECT 59.200 97.900 60.200 98.200 ;
        RECT 55.000 97.500 55.400 97.900 ;
        RECT 57.100 97.600 57.400 97.900 ;
        RECT 56.700 97.300 58.500 97.600 ;
        RECT 59.800 97.500 60.200 97.900 ;
        RECT 56.700 97.200 57.100 97.300 ;
        RECT 58.100 97.200 58.500 97.300 ;
        RECT 54.600 96.600 55.300 97.000 ;
        RECT 55.000 96.100 55.300 96.600 ;
        RECT 56.100 96.500 57.200 96.800 ;
        RECT 56.100 96.400 56.500 96.500 ;
        RECT 55.000 95.800 56.200 96.100 ;
        RECT 52.600 95.300 54.700 95.600 ;
        RECT 50.200 94.100 50.600 94.200 ;
        RECT 51.800 94.100 52.200 94.200 ;
        RECT 50.200 93.800 52.200 94.100 ;
        RECT 50.200 93.400 50.600 93.800 ;
        RECT 52.600 93.600 53.000 95.300 ;
        RECT 54.300 95.200 54.700 95.300 ;
        RECT 53.500 94.900 53.900 95.000 ;
        RECT 53.500 94.600 55.400 94.900 ;
        RECT 55.000 94.500 55.400 94.600 ;
        RECT 55.900 94.200 56.200 95.800 ;
        RECT 56.900 95.900 57.200 96.500 ;
        RECT 57.500 96.500 57.900 96.600 ;
        RECT 59.800 96.500 60.200 96.600 ;
        RECT 57.500 96.200 60.200 96.500 ;
        RECT 56.900 95.700 59.300 95.900 ;
        RECT 61.400 95.700 61.800 99.900 ;
        RECT 62.600 96.800 63.000 97.200 ;
        RECT 62.600 96.200 62.900 96.800 ;
        RECT 63.300 96.200 63.700 99.900 ;
        RECT 62.200 95.900 62.900 96.200 ;
        RECT 62.200 95.800 62.600 95.900 ;
        RECT 63.200 95.800 64.200 96.200 ;
        RECT 56.900 95.600 61.800 95.700 ;
        RECT 58.900 95.500 61.800 95.600 ;
        RECT 59.000 95.400 61.800 95.500 ;
        RECT 58.200 95.100 58.600 95.200 ;
        RECT 58.200 94.800 60.700 95.100 ;
        RECT 60.300 94.700 60.700 94.800 ;
        RECT 59.500 94.200 59.900 94.300 ;
        RECT 63.200 94.200 63.500 95.800 ;
        RECT 65.400 95.600 65.800 99.900 ;
        RECT 67.500 97.900 68.100 99.900 ;
        RECT 69.800 97.900 70.200 99.900 ;
        RECT 72.000 98.200 72.400 99.900 ;
        RECT 72.000 97.900 73.000 98.200 ;
        RECT 67.800 97.500 68.200 97.900 ;
        RECT 69.900 97.600 70.200 97.900 ;
        RECT 69.500 97.300 71.300 97.600 ;
        RECT 72.600 97.500 73.000 97.900 ;
        RECT 69.500 97.200 69.900 97.300 ;
        RECT 70.900 97.200 71.300 97.300 ;
        RECT 67.000 97.000 67.700 97.200 ;
        RECT 67.000 96.800 68.100 97.000 ;
        RECT 67.400 96.600 68.100 96.800 ;
        RECT 67.800 96.100 68.100 96.600 ;
        RECT 68.900 96.500 70.000 96.800 ;
        RECT 68.900 96.400 69.300 96.500 ;
        RECT 67.800 95.800 69.000 96.100 ;
        RECT 65.400 95.300 67.500 95.600 ;
        RECT 63.800 94.400 64.200 95.200 ;
        RECT 55.900 93.900 61.400 94.200 ;
        RECT 56.100 93.800 56.500 93.900 ;
        RECT 44.600 91.500 45.000 92.500 ;
        RECT 45.400 93.000 47.400 93.100 ;
        RECT 45.400 91.100 45.800 93.000 ;
        RECT 47.000 91.100 47.400 93.000 ;
        RECT 47.800 91.100 48.200 93.100 ;
        RECT 48.900 92.800 49.800 93.100 ;
        RECT 52.600 93.300 54.500 93.600 ;
        RECT 48.900 91.100 49.300 92.800 ;
        RECT 51.800 92.100 52.200 92.200 ;
        RECT 52.600 92.100 53.000 93.300 ;
        RECT 54.100 93.200 54.500 93.300 ;
        RECT 59.000 92.800 59.300 93.900 ;
        RECT 60.600 93.800 61.400 93.900 ;
        RECT 62.200 93.800 63.500 94.200 ;
        RECT 64.600 94.100 65.000 94.200 ;
        RECT 64.200 93.800 65.000 94.100 ;
        RECT 58.100 92.700 58.500 92.800 ;
        RECT 55.000 92.100 55.400 92.500 ;
        RECT 57.100 92.400 58.500 92.700 ;
        RECT 59.000 92.400 59.400 92.800 ;
        RECT 57.100 92.100 57.400 92.400 ;
        RECT 59.800 92.100 60.200 92.500 ;
        RECT 51.800 91.800 53.000 92.100 ;
        RECT 52.600 91.100 53.000 91.800 ;
        RECT 54.700 91.800 55.400 92.100 ;
        RECT 54.700 91.100 55.300 91.800 ;
        RECT 57.000 91.100 57.400 92.100 ;
        RECT 59.200 91.800 60.200 92.100 ;
        RECT 59.200 91.100 59.600 91.800 ;
        RECT 61.400 91.100 61.800 93.500 ;
        RECT 62.300 93.100 62.600 93.800 ;
        RECT 64.200 93.600 64.600 93.800 ;
        RECT 65.400 93.600 65.800 95.300 ;
        RECT 67.100 95.200 67.500 95.300 ;
        RECT 66.300 94.900 66.700 95.000 ;
        RECT 66.300 94.600 68.200 94.900 ;
        RECT 67.800 94.500 68.200 94.600 ;
        RECT 68.700 94.200 69.000 95.800 ;
        RECT 69.700 95.900 70.000 96.500 ;
        RECT 70.300 96.500 70.700 96.600 ;
        RECT 72.600 96.500 73.000 96.600 ;
        RECT 70.300 96.200 73.000 96.500 ;
        RECT 69.700 95.700 72.100 95.900 ;
        RECT 74.200 95.700 74.600 99.900 ;
        RECT 69.700 95.600 74.600 95.700 ;
        RECT 75.800 95.600 76.200 99.900 ;
        RECT 77.400 95.600 77.800 99.900 ;
        RECT 79.000 95.600 79.400 99.900 ;
        RECT 80.600 95.600 81.000 99.900 ;
        RECT 71.700 95.500 74.600 95.600 ;
        RECT 71.800 95.400 74.600 95.500 ;
        RECT 75.000 95.200 76.200 95.600 ;
        RECT 76.700 95.200 77.800 95.600 ;
        RECT 78.300 95.200 79.400 95.600 ;
        RECT 80.100 95.200 81.000 95.600 ;
        RECT 82.200 97.500 82.600 99.500 ;
        RECT 82.200 95.800 82.500 97.500 ;
        RECT 84.300 96.400 84.700 99.900 ;
        RECT 88.900 96.400 89.300 99.900 ;
        RECT 91.000 97.500 91.400 99.500 ;
        RECT 84.300 96.100 85.100 96.400 ;
        RECT 82.200 95.500 84.100 95.800 ;
        RECT 71.000 95.100 71.400 95.200 ;
        RECT 71.000 94.800 73.500 95.100 ;
        RECT 73.100 94.700 73.500 94.800 ;
        RECT 72.300 94.200 72.700 94.300 ;
        RECT 68.700 93.900 74.200 94.200 ;
        RECT 68.900 93.800 69.300 93.900 ;
        RECT 65.400 93.300 67.300 93.600 ;
        RECT 63.100 93.100 64.900 93.300 ;
        RECT 62.200 91.100 62.600 93.100 ;
        RECT 63.000 93.000 65.000 93.100 ;
        RECT 63.000 91.100 63.400 93.000 ;
        RECT 64.600 91.100 65.000 93.000 ;
        RECT 65.400 91.100 65.800 93.300 ;
        RECT 66.900 93.200 67.300 93.300 ;
        RECT 71.800 92.800 72.100 93.900 ;
        RECT 73.400 93.800 74.200 93.900 ;
        RECT 75.000 93.800 75.400 95.200 ;
        RECT 76.700 94.500 77.100 95.200 ;
        RECT 78.300 94.500 78.700 95.200 ;
        RECT 80.100 94.500 80.500 95.200 ;
        RECT 75.800 94.100 77.100 94.500 ;
        RECT 77.500 94.100 78.700 94.500 ;
        RECT 79.200 94.100 80.500 94.500 ;
        RECT 80.900 94.100 81.800 94.500 ;
        RECT 82.200 94.400 82.600 95.200 ;
        RECT 83.000 94.400 83.400 95.200 ;
        RECT 83.800 94.500 84.100 95.500 ;
        RECT 76.700 93.800 77.100 94.100 ;
        RECT 78.300 93.800 78.700 94.100 ;
        RECT 80.100 93.800 80.500 94.100 ;
        RECT 81.400 93.800 81.800 94.100 ;
        RECT 83.800 94.100 84.500 94.500 ;
        RECT 84.800 94.200 85.100 96.100 ;
        RECT 88.500 96.100 89.300 96.400 ;
        RECT 85.400 95.100 85.800 95.600 ;
        RECT 85.400 94.800 86.500 95.100 ;
        RECT 87.800 94.800 88.200 95.600 ;
        RECT 83.800 93.900 84.300 94.100 ;
        RECT 70.900 92.700 71.300 92.800 ;
        RECT 67.800 92.100 68.200 92.500 ;
        RECT 69.900 92.400 71.300 92.700 ;
        RECT 71.800 92.400 72.200 92.800 ;
        RECT 69.900 92.100 70.200 92.400 ;
        RECT 72.600 92.100 73.000 92.500 ;
        RECT 67.500 91.800 68.200 92.100 ;
        RECT 67.500 91.100 68.100 91.800 ;
        RECT 69.800 91.100 70.200 92.100 ;
        RECT 72.000 91.800 73.000 92.100 ;
        RECT 72.000 91.100 72.400 91.800 ;
        RECT 74.200 91.100 74.600 93.500 ;
        RECT 75.000 93.400 76.200 93.800 ;
        RECT 76.700 93.400 77.800 93.800 ;
        RECT 78.300 93.400 79.400 93.800 ;
        RECT 80.100 93.400 81.000 93.800 ;
        RECT 75.800 91.100 76.200 93.400 ;
        RECT 77.400 91.100 77.800 93.400 ;
        RECT 79.000 91.100 79.400 93.400 ;
        RECT 80.600 91.100 81.000 93.400 ;
        RECT 82.200 93.600 84.300 93.900 ;
        RECT 84.800 93.800 85.800 94.200 ;
        RECT 86.200 94.100 86.500 94.800 ;
        RECT 88.500 94.200 88.800 96.100 ;
        RECT 91.100 95.800 91.400 97.500 ;
        RECT 89.500 95.500 91.400 95.800 ;
        RECT 91.800 97.500 92.200 99.500 ;
        RECT 91.800 95.800 92.100 97.500 ;
        RECT 93.900 96.400 94.300 99.900 ;
        RECT 93.900 96.100 94.700 96.400 ;
        RECT 91.800 95.500 93.700 95.800 ;
        RECT 89.500 94.500 89.800 95.500 ;
        RECT 87.800 94.100 88.800 94.200 ;
        RECT 89.100 94.100 89.800 94.500 ;
        RECT 90.200 94.400 90.600 95.200 ;
        RECT 91.000 94.400 91.400 95.200 ;
        RECT 91.800 94.400 92.200 95.200 ;
        RECT 92.600 94.400 93.000 95.200 ;
        RECT 93.400 94.500 93.700 95.500 ;
        RECT 86.200 93.800 88.800 94.100 ;
        RECT 82.200 92.500 82.500 93.600 ;
        RECT 84.800 93.500 85.100 93.800 ;
        RECT 84.700 93.300 85.100 93.500 ;
        RECT 84.300 93.000 85.100 93.300 ;
        RECT 88.500 93.500 88.800 93.800 ;
        RECT 89.300 93.900 89.800 94.100 ;
        RECT 93.400 94.100 94.100 94.500 ;
        RECT 94.400 94.200 94.700 96.100 ;
        RECT 95.000 95.100 95.400 95.600 ;
        RECT 96.600 95.100 97.000 99.900 ;
        RECT 95.000 94.800 97.000 95.100 ;
        RECT 94.400 94.100 95.400 94.200 ;
        RECT 95.800 94.100 96.200 94.200 ;
        RECT 93.400 93.900 93.900 94.100 ;
        RECT 89.300 93.600 91.400 93.900 ;
        RECT 88.500 93.300 88.900 93.500 ;
        RECT 88.500 93.000 89.300 93.300 ;
        RECT 82.200 91.500 82.600 92.500 ;
        RECT 84.300 92.200 84.700 93.000 ;
        RECT 83.800 91.800 84.700 92.200 ;
        RECT 84.300 91.500 84.700 91.800 ;
        RECT 88.900 91.500 89.300 93.000 ;
        RECT 91.100 92.500 91.400 93.600 ;
        RECT 91.000 91.500 91.400 92.500 ;
        RECT 91.800 93.600 93.900 93.900 ;
        RECT 94.400 93.800 96.200 94.100 ;
        RECT 91.800 92.500 92.100 93.600 ;
        RECT 94.400 93.500 94.700 93.800 ;
        RECT 94.300 93.300 94.700 93.500 ;
        RECT 93.900 93.000 94.700 93.300 ;
        RECT 91.800 91.500 92.200 92.500 ;
        RECT 93.900 91.500 94.300 93.000 ;
        RECT 96.600 91.100 97.000 94.800 ;
        RECT 98.200 95.600 98.600 99.900 ;
        RECT 100.300 97.900 100.900 99.900 ;
        RECT 102.600 97.900 103.000 99.900 ;
        RECT 104.800 98.200 105.200 99.900 ;
        RECT 104.800 97.900 105.800 98.200 ;
        RECT 100.600 97.500 101.000 97.900 ;
        RECT 102.700 97.600 103.000 97.900 ;
        RECT 102.300 97.300 104.100 97.600 ;
        RECT 105.400 97.500 105.800 97.900 ;
        RECT 102.300 97.200 102.700 97.300 ;
        RECT 103.700 97.200 104.100 97.300 ;
        RECT 100.200 96.600 100.900 97.000 ;
        RECT 100.600 96.100 100.900 96.600 ;
        RECT 101.700 96.500 102.800 96.800 ;
        RECT 101.700 96.400 102.100 96.500 ;
        RECT 100.600 95.800 101.800 96.100 ;
        RECT 98.200 95.300 100.300 95.600 ;
        RECT 97.400 93.800 97.800 94.200 ;
        RECT 97.400 93.200 97.700 93.800 ;
        RECT 98.200 93.600 98.600 95.300 ;
        RECT 99.900 95.200 100.300 95.300 ;
        RECT 99.100 94.900 99.500 95.000 ;
        RECT 99.100 94.600 101.000 94.900 ;
        RECT 100.600 94.500 101.000 94.600 ;
        RECT 101.500 94.200 101.800 95.800 ;
        RECT 102.500 95.900 102.800 96.500 ;
        RECT 103.100 96.500 103.500 96.600 ;
        RECT 105.400 96.500 105.800 96.600 ;
        RECT 103.100 96.200 105.800 96.500 ;
        RECT 102.500 95.700 104.900 95.900 ;
        RECT 107.000 95.700 107.400 99.900 ;
        RECT 102.500 95.600 107.400 95.700 ;
        RECT 104.500 95.500 107.400 95.600 ;
        RECT 109.400 97.500 109.800 99.500 ;
        RECT 109.400 95.800 109.700 97.500 ;
        RECT 111.500 96.400 111.900 99.900 ;
        RECT 111.500 96.100 112.300 96.400 ;
        RECT 109.400 95.500 111.300 95.800 ;
        RECT 104.600 95.400 107.400 95.500 ;
        RECT 103.800 95.100 104.200 95.200 ;
        RECT 108.600 95.100 109.000 95.200 ;
        RECT 109.400 95.100 109.800 95.200 ;
        RECT 103.800 94.800 106.300 95.100 ;
        RECT 108.600 94.800 109.800 95.100 ;
        RECT 105.900 94.700 106.300 94.800 ;
        RECT 109.400 94.400 109.800 94.800 ;
        RECT 110.200 94.400 110.600 95.200 ;
        RECT 111.000 94.500 111.300 95.500 ;
        RECT 105.100 94.200 105.500 94.300 ;
        RECT 101.400 93.900 107.000 94.200 ;
        RECT 111.000 94.100 111.700 94.500 ;
        RECT 112.000 94.200 112.300 96.100 ;
        RECT 112.600 95.100 113.000 95.600 ;
        RECT 114.200 95.100 114.600 99.900 ;
        RECT 115.800 95.700 116.200 99.900 ;
        RECT 118.000 98.200 118.400 99.900 ;
        RECT 117.400 97.900 118.400 98.200 ;
        RECT 120.200 97.900 120.600 99.900 ;
        RECT 122.300 97.900 122.900 99.900 ;
        RECT 117.400 97.500 117.800 97.900 ;
        RECT 120.200 97.600 120.500 97.900 ;
        RECT 119.100 97.300 120.900 97.600 ;
        RECT 122.200 97.500 122.600 97.900 ;
        RECT 119.100 97.200 119.500 97.300 ;
        RECT 120.500 97.200 120.900 97.300 ;
        RECT 117.400 96.500 117.800 96.600 ;
        RECT 119.700 96.500 120.100 96.600 ;
        RECT 117.400 96.200 120.100 96.500 ;
        RECT 120.400 96.500 121.500 96.800 ;
        RECT 120.400 95.900 120.700 96.500 ;
        RECT 121.100 96.400 121.500 96.500 ;
        RECT 122.300 96.600 123.000 97.000 ;
        RECT 122.300 96.100 122.600 96.600 ;
        RECT 118.300 95.700 120.700 95.900 ;
        RECT 115.800 95.600 120.700 95.700 ;
        RECT 121.400 95.800 122.600 96.100 ;
        RECT 115.800 95.500 118.700 95.600 ;
        RECT 115.800 95.400 118.600 95.500 ;
        RECT 119.000 95.100 119.400 95.200 ;
        RECT 112.600 94.800 114.600 95.100 ;
        RECT 112.000 94.100 113.000 94.200 ;
        RECT 113.400 94.100 113.800 94.200 ;
        RECT 111.000 93.900 111.500 94.100 ;
        RECT 101.400 93.800 102.100 93.900 ;
        RECT 98.200 93.300 100.100 93.600 ;
        RECT 97.400 93.100 97.800 93.200 ;
        RECT 98.200 93.100 98.600 93.300 ;
        RECT 99.700 93.200 100.100 93.300 ;
        RECT 97.400 92.800 98.600 93.100 ;
        RECT 104.600 92.800 104.900 93.900 ;
        RECT 106.200 93.800 107.000 93.900 ;
        RECT 109.400 93.600 111.500 93.900 ;
        RECT 112.000 93.800 113.800 94.100 ;
        RECT 97.400 92.400 97.800 92.800 ;
        RECT 98.200 91.100 98.600 92.800 ;
        RECT 103.700 92.700 104.100 92.800 ;
        RECT 100.600 92.100 101.000 92.500 ;
        RECT 102.700 92.400 104.100 92.700 ;
        RECT 104.600 92.400 105.000 92.800 ;
        RECT 102.700 92.100 103.000 92.400 ;
        RECT 105.400 92.100 105.800 92.500 ;
        RECT 100.300 91.800 101.000 92.100 ;
        RECT 100.300 91.100 100.900 91.800 ;
        RECT 102.600 91.100 103.000 92.100 ;
        RECT 104.800 91.800 105.800 92.100 ;
        RECT 104.800 91.100 105.200 91.800 ;
        RECT 107.000 91.100 107.400 93.500 ;
        RECT 109.400 92.500 109.700 93.600 ;
        RECT 112.000 93.500 112.300 93.800 ;
        RECT 111.900 93.300 112.300 93.500 ;
        RECT 111.500 93.000 112.300 93.300 ;
        RECT 109.400 91.500 109.800 92.500 ;
        RECT 111.500 91.500 111.900 93.000 ;
        RECT 114.200 91.100 114.600 94.800 ;
        RECT 116.900 94.800 119.400 95.100 ;
        RECT 116.900 94.700 117.300 94.800 ;
        RECT 118.200 94.700 118.600 94.800 ;
        RECT 117.700 94.200 118.100 94.300 ;
        RECT 121.400 94.200 121.700 95.800 ;
        RECT 124.600 95.600 125.000 99.900 ;
        RECT 122.900 95.300 125.000 95.600 ;
        RECT 122.900 95.200 123.300 95.300 ;
        RECT 123.700 94.900 124.100 95.000 ;
        RECT 122.200 94.600 124.100 94.900 ;
        RECT 122.200 94.500 122.600 94.600 ;
        RECT 116.200 93.900 121.700 94.200 ;
        RECT 116.200 93.800 117.000 93.900 ;
        RECT 115.000 92.400 115.400 93.200 ;
        RECT 115.800 91.100 116.200 93.500 ;
        RECT 118.300 92.800 118.600 93.900 ;
        RECT 119.800 93.800 120.200 93.900 ;
        RECT 121.100 93.800 121.500 93.900 ;
        RECT 124.600 93.600 125.000 95.300 ;
        RECT 123.100 93.300 125.000 93.600 ;
        RECT 123.100 93.200 123.500 93.300 ;
        RECT 117.400 92.100 117.800 92.500 ;
        RECT 118.200 92.400 118.600 92.800 ;
        RECT 119.100 92.700 119.500 92.800 ;
        RECT 119.100 92.400 120.500 92.700 ;
        RECT 120.200 92.100 120.500 92.400 ;
        RECT 122.200 92.100 122.600 92.500 ;
        RECT 117.400 91.800 118.400 92.100 ;
        RECT 118.000 91.100 118.400 91.800 ;
        RECT 120.200 91.100 120.600 92.100 ;
        RECT 122.200 91.800 122.900 92.100 ;
        RECT 122.300 91.100 122.900 91.800 ;
        RECT 124.600 91.100 125.000 93.300 ;
        RECT 125.400 92.400 125.800 93.200 ;
        RECT 126.200 93.100 126.600 99.900 ;
        RECT 128.300 96.300 128.700 99.900 ;
        RECT 127.800 95.900 128.700 96.300 ;
        RECT 129.400 97.500 129.800 99.500 ;
        RECT 131.500 99.200 131.900 99.900 ;
        RECT 131.500 98.800 132.200 99.200 ;
        RECT 127.000 95.100 127.400 95.200 ;
        RECT 127.900 95.100 128.200 95.900 ;
        RECT 129.400 95.800 129.700 97.500 ;
        RECT 131.500 96.400 131.900 98.800 ;
        RECT 131.500 96.100 132.300 96.400 ;
        RECT 127.000 94.800 128.200 95.100 ;
        RECT 128.600 94.800 129.000 95.600 ;
        RECT 129.400 95.500 131.300 95.800 ;
        RECT 127.900 94.200 128.200 94.800 ;
        RECT 129.400 94.400 129.800 95.200 ;
        RECT 130.200 94.400 130.600 95.200 ;
        RECT 131.000 94.500 131.300 95.500 ;
        RECT 127.800 93.800 128.200 94.200 ;
        RECT 131.000 94.100 131.700 94.500 ;
        RECT 132.000 94.200 132.300 96.100 ;
        RECT 134.200 96.200 134.600 99.900 ;
        RECT 135.800 96.400 136.200 99.900 ;
        RECT 134.200 95.900 135.500 96.200 ;
        RECT 135.800 95.900 136.300 96.400 ;
        RECT 137.400 96.200 137.800 99.900 ;
        RECT 139.000 96.200 139.400 99.900 ;
        RECT 137.400 95.900 139.400 96.200 ;
        RECT 139.800 95.900 140.200 99.900 ;
        RECT 132.600 94.800 133.000 95.600 ;
        RECT 134.200 94.800 134.700 95.200 ;
        RECT 134.300 94.400 134.700 94.800 ;
        RECT 135.200 94.900 135.500 95.900 ;
        RECT 135.200 94.500 135.700 94.900 ;
        RECT 131.000 93.900 131.500 94.100 ;
        RECT 127.000 93.100 127.400 93.200 ;
        RECT 126.200 92.800 127.400 93.100 ;
        RECT 126.200 91.100 126.600 92.800 ;
        RECT 127.000 92.400 127.400 92.800 ;
        RECT 127.900 92.100 128.200 93.800 ;
        RECT 127.800 91.100 128.200 92.100 ;
        RECT 129.400 93.600 131.500 93.900 ;
        RECT 132.000 93.800 133.000 94.200 ;
        RECT 129.400 92.500 129.700 93.600 ;
        RECT 132.000 93.500 132.300 93.800 ;
        RECT 135.200 93.700 135.500 94.500 ;
        RECT 136.000 94.200 136.300 95.900 ;
        RECT 137.800 95.200 138.200 95.400 ;
        RECT 139.800 95.200 140.100 95.900 ;
        RECT 140.600 95.700 141.000 99.900 ;
        RECT 142.800 98.200 143.200 99.900 ;
        RECT 142.200 97.900 143.200 98.200 ;
        RECT 145.000 97.900 145.400 99.900 ;
        RECT 147.100 97.900 147.700 99.900 ;
        RECT 142.200 97.500 142.600 97.900 ;
        RECT 145.000 97.600 145.300 97.900 ;
        RECT 143.900 97.300 145.700 97.600 ;
        RECT 147.000 97.500 147.400 97.900 ;
        RECT 143.900 97.200 144.300 97.300 ;
        RECT 145.300 97.200 145.700 97.300 ;
        RECT 142.200 96.500 142.600 96.600 ;
        RECT 144.500 96.500 144.900 96.600 ;
        RECT 142.200 96.200 144.900 96.500 ;
        RECT 145.200 96.500 146.300 96.800 ;
        RECT 145.200 95.900 145.500 96.500 ;
        RECT 145.900 96.400 146.300 96.500 ;
        RECT 147.100 96.600 147.800 97.000 ;
        RECT 147.100 96.100 147.400 96.600 ;
        RECT 143.100 95.700 145.500 95.900 ;
        RECT 140.600 95.600 145.500 95.700 ;
        RECT 146.200 95.800 147.400 96.100 ;
        RECT 140.600 95.500 143.500 95.600 ;
        RECT 140.600 95.400 143.400 95.500 ;
        RECT 137.400 94.900 138.200 95.200 ;
        RECT 139.000 94.900 140.200 95.200 ;
        RECT 143.800 95.100 144.200 95.200 ;
        RECT 137.400 94.800 137.800 94.900 ;
        RECT 135.800 93.800 136.300 94.200 ;
        RECT 138.200 93.800 138.600 94.600 ;
        RECT 131.900 93.300 132.300 93.500 ;
        RECT 131.500 93.000 132.300 93.300 ;
        RECT 134.200 93.400 135.500 93.700 ;
        RECT 129.400 91.500 129.800 92.500 ;
        RECT 131.500 91.500 131.900 93.000 ;
        RECT 134.200 91.100 134.600 93.400 ;
        RECT 136.000 93.100 136.300 93.800 ;
        RECT 135.800 92.800 136.300 93.100 ;
        RECT 139.000 93.100 139.300 94.900 ;
        RECT 139.800 94.800 140.200 94.900 ;
        RECT 141.700 94.800 144.200 95.100 ;
        RECT 141.700 94.700 142.100 94.800 ;
        RECT 143.000 94.700 143.400 94.800 ;
        RECT 142.500 94.200 142.900 94.300 ;
        RECT 146.200 94.200 146.500 95.800 ;
        RECT 149.400 95.600 149.800 99.900 ;
        RECT 151.500 96.300 151.900 99.900 ;
        RECT 154.500 99.200 154.900 99.900 ;
        RECT 154.500 98.800 155.400 99.200 ;
        RECT 154.500 96.400 154.900 98.800 ;
        RECT 156.600 97.500 157.000 99.500 ;
        RECT 151.000 95.900 151.900 96.300 ;
        RECT 154.100 96.100 154.900 96.400 ;
        RECT 151.000 95.800 151.400 95.900 ;
        RECT 147.700 95.300 149.800 95.600 ;
        RECT 147.700 95.200 148.100 95.300 ;
        RECT 148.500 94.900 148.900 95.000 ;
        RECT 147.000 94.600 148.900 94.900 ;
        RECT 147.000 94.500 147.400 94.600 ;
        RECT 141.000 93.900 146.500 94.200 ;
        RECT 141.000 93.800 141.800 93.900 ;
        RECT 135.800 91.100 136.200 92.800 ;
        RECT 139.000 91.100 139.400 93.100 ;
        RECT 139.800 92.800 140.200 93.200 ;
        RECT 139.700 92.400 140.100 92.800 ;
        RECT 140.600 91.100 141.000 93.500 ;
        RECT 143.100 93.200 143.400 93.900 ;
        RECT 145.900 93.800 146.300 93.900 ;
        RECT 149.400 93.600 149.800 95.300 ;
        RECT 151.100 94.200 151.400 95.800 ;
        RECT 151.800 94.800 152.200 95.600 ;
        RECT 153.400 95.100 153.800 95.600 ;
        RECT 152.600 94.800 153.800 95.100 ;
        RECT 151.000 93.800 151.400 94.200 ;
        RECT 152.600 94.200 152.900 94.800 ;
        RECT 154.100 94.200 154.400 96.100 ;
        RECT 156.700 95.800 157.000 97.500 ;
        RECT 155.100 95.500 157.000 95.800 ;
        RECT 155.100 94.500 155.400 95.500 ;
        RECT 152.600 93.800 153.000 94.200 ;
        RECT 153.400 93.800 154.400 94.200 ;
        RECT 154.700 94.100 155.400 94.500 ;
        RECT 155.800 94.400 156.200 95.200 ;
        RECT 156.600 95.100 157.000 95.200 ;
        RECT 158.200 95.100 158.600 95.200 ;
        RECT 156.600 94.800 158.600 95.100 ;
        RECT 156.600 94.400 157.000 94.800 ;
        RECT 147.900 93.300 149.800 93.600 ;
        RECT 147.900 93.200 148.300 93.300 ;
        RECT 142.200 92.100 142.600 92.500 ;
        RECT 143.000 92.400 143.400 93.200 ;
        RECT 143.900 92.700 144.300 92.800 ;
        RECT 143.900 92.400 145.300 92.700 ;
        RECT 145.000 92.100 145.300 92.400 ;
        RECT 147.000 92.100 147.400 92.500 ;
        RECT 142.200 91.800 143.200 92.100 ;
        RECT 142.800 91.100 143.200 91.800 ;
        RECT 145.000 91.100 145.400 92.100 ;
        RECT 147.000 91.800 147.700 92.100 ;
        RECT 147.100 91.100 147.700 91.800 ;
        RECT 149.400 91.100 149.800 93.300 ;
        RECT 150.200 92.400 150.600 93.200 ;
        RECT 151.100 92.100 151.400 93.800 ;
        RECT 154.100 93.500 154.400 93.800 ;
        RECT 154.900 93.900 155.400 94.100 ;
        RECT 157.400 94.100 157.800 94.200 ;
        RECT 159.000 94.100 159.400 94.200 ;
        RECT 154.900 93.600 157.000 93.900 ;
        RECT 157.400 93.800 159.400 94.100 ;
        RECT 154.100 93.300 154.500 93.500 ;
        RECT 154.100 93.000 154.900 93.300 ;
        RECT 151.000 91.100 151.400 92.100 ;
        RECT 154.500 91.500 154.900 93.000 ;
        RECT 156.700 92.500 157.000 93.600 ;
        RECT 159.000 93.400 159.400 93.800 ;
        RECT 159.800 93.100 160.200 99.900 ;
        RECT 160.600 95.800 161.000 96.600 ;
        RECT 161.400 95.700 161.800 99.900 ;
        RECT 163.600 98.200 164.000 99.900 ;
        RECT 163.000 97.900 164.000 98.200 ;
        RECT 165.800 97.900 166.200 99.900 ;
        RECT 167.900 97.900 168.500 99.900 ;
        RECT 163.000 97.500 163.400 97.900 ;
        RECT 165.800 97.600 166.100 97.900 ;
        RECT 164.700 97.300 166.500 97.600 ;
        RECT 167.800 97.500 168.200 97.900 ;
        RECT 164.700 97.200 165.100 97.300 ;
        RECT 166.100 97.200 166.500 97.300 ;
        RECT 163.000 96.500 163.400 96.600 ;
        RECT 165.300 96.500 165.700 96.600 ;
        RECT 163.000 96.200 165.700 96.500 ;
        RECT 166.000 96.500 167.100 96.800 ;
        RECT 166.000 95.900 166.300 96.500 ;
        RECT 166.700 96.400 167.100 96.500 ;
        RECT 167.900 96.600 168.600 97.000 ;
        RECT 167.900 96.100 168.200 96.600 ;
        RECT 163.900 95.700 166.300 95.900 ;
        RECT 161.400 95.600 166.300 95.700 ;
        RECT 167.000 95.800 168.200 96.100 ;
        RECT 161.400 95.500 164.300 95.600 ;
        RECT 161.400 95.400 164.200 95.500 ;
        RECT 164.600 95.100 165.000 95.200 ;
        RECT 162.500 94.800 165.000 95.100 ;
        RECT 162.500 94.700 162.900 94.800 ;
        RECT 163.300 94.200 163.700 94.300 ;
        RECT 167.000 94.200 167.300 95.800 ;
        RECT 170.200 95.600 170.600 99.900 ;
        RECT 168.500 95.300 170.600 95.600 ;
        RECT 168.500 95.200 168.900 95.300 ;
        RECT 169.300 94.900 169.700 95.000 ;
        RECT 167.800 94.600 169.700 94.900 ;
        RECT 167.800 94.500 168.200 94.600 ;
        RECT 161.800 93.900 167.300 94.200 ;
        RECT 170.200 94.100 170.600 95.300 ;
        RECT 171.800 95.100 172.200 99.900 ;
        RECT 173.800 96.800 174.200 97.200 ;
        RECT 172.600 95.800 173.000 96.600 ;
        RECT 173.800 96.200 174.100 96.800 ;
        RECT 174.500 96.200 174.900 99.900 ;
        RECT 178.500 99.200 178.900 99.900 ;
        RECT 178.200 98.800 178.900 99.200 ;
        RECT 178.500 96.400 178.900 98.800 ;
        RECT 180.600 97.500 181.000 99.500 ;
        RECT 183.300 99.200 183.700 99.900 ;
        RECT 183.000 98.800 183.700 99.200 ;
        RECT 173.400 95.900 174.100 96.200 ;
        RECT 174.400 95.900 174.900 96.200 ;
        RECT 178.100 96.100 178.900 96.400 ;
        RECT 173.400 95.800 173.800 95.900 ;
        RECT 173.400 95.100 173.700 95.800 ;
        RECT 171.800 94.800 173.700 95.100 ;
        RECT 171.000 94.100 171.400 94.200 ;
        RECT 161.800 93.800 162.600 93.900 ;
        RECT 159.800 92.800 160.700 93.100 ;
        RECT 156.600 91.500 157.000 92.500 ;
        RECT 160.300 92.200 160.700 92.800 ;
        RECT 160.300 91.800 161.000 92.200 ;
        RECT 160.300 91.100 160.700 91.800 ;
        RECT 161.400 91.100 161.800 93.500 ;
        RECT 163.900 93.200 164.200 93.900 ;
        RECT 166.700 93.800 167.100 93.900 ;
        RECT 170.200 93.800 171.400 94.100 ;
        RECT 170.200 93.600 170.600 93.800 ;
        RECT 163.000 92.100 163.400 92.500 ;
        RECT 163.800 92.400 164.200 93.200 ;
        RECT 168.600 93.300 170.600 93.600 ;
        RECT 171.000 93.400 171.400 93.800 ;
        RECT 168.600 93.200 169.100 93.300 ;
        RECT 168.600 92.800 169.000 93.200 ;
        RECT 164.700 92.700 165.100 92.800 ;
        RECT 164.700 92.400 166.100 92.700 ;
        RECT 165.800 92.100 166.100 92.400 ;
        RECT 167.800 92.100 168.200 92.500 ;
        RECT 163.000 91.800 164.000 92.100 ;
        RECT 163.600 91.100 164.000 91.800 ;
        RECT 165.800 91.100 166.200 92.100 ;
        RECT 167.800 91.800 168.500 92.100 ;
        RECT 167.900 91.100 168.500 91.800 ;
        RECT 170.200 91.100 170.600 93.300 ;
        RECT 171.800 93.100 172.200 94.800 ;
        RECT 174.400 94.200 174.700 95.900 ;
        RECT 175.000 94.400 175.400 95.200 ;
        RECT 177.400 94.800 177.800 95.600 ;
        RECT 178.100 94.200 178.400 96.100 ;
        RECT 180.700 95.800 181.000 97.500 ;
        RECT 183.300 96.400 183.700 98.800 ;
        RECT 185.400 97.500 185.800 99.500 ;
        RECT 179.100 95.500 181.000 95.800 ;
        RECT 182.900 96.100 183.700 96.400 ;
        RECT 179.100 94.500 179.400 95.500 ;
        RECT 172.600 94.100 173.000 94.200 ;
        RECT 173.400 94.100 174.700 94.200 ;
        RECT 175.800 94.100 176.200 94.200 ;
        RECT 176.600 94.100 177.000 94.200 ;
        RECT 172.600 93.800 174.700 94.100 ;
        RECT 175.400 93.800 177.000 94.100 ;
        RECT 177.400 93.800 178.400 94.200 ;
        RECT 178.700 94.100 179.400 94.500 ;
        RECT 179.800 94.400 180.200 95.200 ;
        RECT 180.600 94.400 181.000 95.200 ;
        RECT 182.200 94.800 182.600 95.600 ;
        RECT 182.900 94.200 183.200 96.100 ;
        RECT 185.500 95.800 185.800 97.500 ;
        RECT 188.100 96.400 188.500 99.900 ;
        RECT 190.200 97.500 190.600 99.500 ;
        RECT 183.900 95.500 185.800 95.800 ;
        RECT 187.700 96.100 188.500 96.400 ;
        RECT 183.900 94.500 184.200 95.500 ;
        RECT 173.500 93.100 173.800 93.800 ;
        RECT 175.400 93.600 175.800 93.800 ;
        RECT 178.100 93.500 178.400 93.800 ;
        RECT 178.900 93.900 179.400 94.100 ;
        RECT 178.900 93.600 181.000 93.900 ;
        RECT 182.200 93.800 183.200 94.200 ;
        RECT 183.500 94.100 184.200 94.500 ;
        RECT 184.600 94.400 185.000 95.200 ;
        RECT 185.400 94.400 185.800 95.200 ;
        RECT 187.000 94.800 187.400 95.600 ;
        RECT 187.700 94.200 188.000 96.100 ;
        RECT 190.300 95.800 190.600 97.500 ;
        RECT 188.700 95.500 190.600 95.800 ;
        RECT 188.700 94.500 189.000 95.500 ;
        RECT 178.100 93.300 178.500 93.500 ;
        RECT 174.300 93.100 176.100 93.300 ;
        RECT 171.800 92.800 172.700 93.100 ;
        RECT 172.300 91.100 172.700 92.800 ;
        RECT 173.400 91.100 173.800 93.100 ;
        RECT 174.200 93.000 176.200 93.100 ;
        RECT 178.100 93.000 178.900 93.300 ;
        RECT 174.200 91.100 174.600 93.000 ;
        RECT 175.800 91.100 176.200 93.000 ;
        RECT 178.500 91.500 178.900 93.000 ;
        RECT 180.700 92.500 181.000 93.600 ;
        RECT 182.900 93.500 183.200 93.800 ;
        RECT 183.700 93.900 184.200 94.100 ;
        RECT 186.200 94.100 186.600 94.200 ;
        RECT 187.000 94.100 188.000 94.200 ;
        RECT 188.300 94.100 189.000 94.500 ;
        RECT 189.400 94.400 189.800 95.200 ;
        RECT 190.200 94.400 190.600 95.200 ;
        RECT 191.000 94.800 191.400 95.200 ;
        RECT 183.700 93.600 185.800 93.900 ;
        RECT 186.200 93.800 188.000 94.100 ;
        RECT 182.900 93.300 183.300 93.500 ;
        RECT 182.900 93.000 183.700 93.300 ;
        RECT 180.600 91.500 181.000 92.500 ;
        RECT 183.300 91.500 183.700 93.000 ;
        RECT 185.500 92.500 185.800 93.600 ;
        RECT 187.700 93.500 188.000 93.800 ;
        RECT 188.500 93.900 189.000 94.100 ;
        RECT 191.000 94.200 191.300 94.800 ;
        RECT 188.500 93.600 190.600 93.900 ;
        RECT 187.700 93.300 188.100 93.500 ;
        RECT 187.700 93.000 188.500 93.300 ;
        RECT 185.400 91.500 185.800 92.500 ;
        RECT 188.100 91.500 188.500 93.000 ;
        RECT 190.300 92.500 190.600 93.600 ;
        RECT 191.000 93.400 191.400 94.200 ;
        RECT 191.800 93.100 192.200 99.900 ;
        RECT 192.600 95.800 193.000 96.600 ;
        RECT 194.200 96.400 194.600 99.900 ;
        RECT 194.100 95.900 194.600 96.400 ;
        RECT 195.800 96.200 196.200 99.900 ;
        RECT 197.400 96.400 197.800 99.900 ;
        RECT 194.900 95.900 196.200 96.200 ;
        RECT 197.300 95.900 197.800 96.400 ;
        RECT 199.000 96.200 199.400 99.900 ;
        RECT 200.600 96.400 201.000 99.900 ;
        RECT 198.100 95.900 199.400 96.200 ;
        RECT 200.500 95.900 201.000 96.400 ;
        RECT 202.200 96.200 202.600 99.900 ;
        RECT 201.300 95.900 202.600 96.200 ;
        RECT 203.000 96.200 203.400 99.900 ;
        RECT 204.600 96.400 205.000 99.900 ;
        RECT 203.000 95.900 204.300 96.200 ;
        RECT 204.600 95.900 205.100 96.400 ;
        RECT 194.100 94.200 194.400 95.900 ;
        RECT 194.900 94.900 195.200 95.900 ;
        RECT 194.700 94.500 195.200 94.900 ;
        RECT 194.100 93.800 194.600 94.200 ;
        RECT 194.100 93.100 194.400 93.800 ;
        RECT 194.900 93.700 195.200 94.500 ;
        RECT 195.700 94.800 196.200 95.200 ;
        RECT 195.700 94.400 196.100 94.800 ;
        RECT 197.300 94.200 197.600 95.900 ;
        RECT 198.100 94.900 198.400 95.900 ;
        RECT 197.900 94.500 198.400 94.900 ;
        RECT 197.300 93.800 197.800 94.200 ;
        RECT 194.900 93.400 196.200 93.700 ;
        RECT 191.800 92.800 192.700 93.100 ;
        RECT 194.100 92.800 194.600 93.100 ;
        RECT 190.200 91.500 190.600 92.500 ;
        RECT 192.300 92.200 192.700 92.800 ;
        RECT 191.800 91.800 192.700 92.200 ;
        RECT 192.300 91.100 192.700 91.800 ;
        RECT 194.200 91.100 194.600 92.800 ;
        RECT 195.800 91.100 196.200 93.400 ;
        RECT 197.300 93.100 197.600 93.800 ;
        RECT 198.100 93.700 198.400 94.500 ;
        RECT 198.900 94.800 199.400 95.200 ;
        RECT 198.900 94.400 199.300 94.800 ;
        RECT 200.500 94.200 200.800 95.900 ;
        RECT 201.300 94.900 201.600 95.900 ;
        RECT 201.100 94.500 201.600 94.900 ;
        RECT 200.500 93.800 201.000 94.200 ;
        RECT 198.100 93.400 199.400 93.700 ;
        RECT 197.300 92.800 197.800 93.100 ;
        RECT 197.400 91.100 197.800 92.800 ;
        RECT 199.000 91.100 199.400 93.400 ;
        RECT 200.500 93.100 200.800 93.800 ;
        RECT 201.300 93.700 201.600 94.500 ;
        RECT 202.100 95.100 202.600 95.200 ;
        RECT 203.000 95.100 203.500 95.200 ;
        RECT 202.100 94.800 203.500 95.100 ;
        RECT 202.100 94.400 202.500 94.800 ;
        RECT 203.100 94.400 203.500 94.800 ;
        RECT 204.000 94.900 204.300 95.900 ;
        RECT 204.000 94.500 204.500 94.900 ;
        RECT 204.000 93.700 204.300 94.500 ;
        RECT 204.800 94.200 205.100 95.900 ;
        RECT 204.600 93.800 205.100 94.200 ;
        RECT 201.300 93.400 202.600 93.700 ;
        RECT 200.500 92.800 201.000 93.100 ;
        RECT 200.600 91.100 201.000 92.800 ;
        RECT 202.200 91.100 202.600 93.400 ;
        RECT 203.000 93.400 204.300 93.700 ;
        RECT 203.000 91.100 203.400 93.400 ;
        RECT 204.800 93.100 205.100 93.800 ;
        RECT 204.600 92.800 205.100 93.100 ;
        RECT 207.800 95.600 208.200 99.900 ;
        RECT 209.900 97.900 210.500 99.900 ;
        RECT 212.200 97.900 212.600 99.900 ;
        RECT 214.400 98.200 214.800 99.900 ;
        RECT 214.400 97.900 215.400 98.200 ;
        RECT 210.200 97.500 210.600 97.900 ;
        RECT 212.300 97.600 212.600 97.900 ;
        RECT 211.900 97.300 213.700 97.600 ;
        RECT 215.000 97.500 215.400 97.900 ;
        RECT 211.900 97.200 212.300 97.300 ;
        RECT 213.300 97.200 213.700 97.300 ;
        RECT 209.800 96.600 210.500 97.000 ;
        RECT 210.200 96.100 210.500 96.600 ;
        RECT 211.300 96.500 212.400 96.800 ;
        RECT 211.300 96.400 211.700 96.500 ;
        RECT 210.200 95.800 211.400 96.100 ;
        RECT 207.800 95.300 209.900 95.600 ;
        RECT 207.800 93.600 208.200 95.300 ;
        RECT 209.500 95.200 209.900 95.300 ;
        RECT 208.700 94.900 209.100 95.000 ;
        RECT 208.700 94.600 210.600 94.900 ;
        RECT 210.200 94.500 210.600 94.600 ;
        RECT 211.100 94.200 211.400 95.800 ;
        RECT 212.100 95.900 212.400 96.500 ;
        RECT 212.700 96.500 213.100 96.600 ;
        RECT 215.000 96.500 215.400 96.600 ;
        RECT 212.700 96.200 215.400 96.500 ;
        RECT 212.100 95.700 214.500 95.900 ;
        RECT 216.600 95.700 217.000 99.900 ;
        RECT 212.100 95.600 217.000 95.700 ;
        RECT 214.100 95.500 217.000 95.600 ;
        RECT 214.200 95.400 217.000 95.500 ;
        RECT 213.400 95.100 213.800 95.200 ;
        RECT 213.400 94.800 215.900 95.100 ;
        RECT 214.200 94.700 214.600 94.800 ;
        RECT 215.500 94.700 215.900 94.800 ;
        RECT 214.700 94.200 215.100 94.300 ;
        RECT 211.100 93.900 216.600 94.200 ;
        RECT 211.300 93.800 211.700 93.900 ;
        RECT 207.800 93.300 209.700 93.600 ;
        RECT 204.600 91.100 205.000 92.800 ;
        RECT 207.800 91.100 208.200 93.300 ;
        RECT 209.300 93.200 209.700 93.300 ;
        RECT 214.200 92.800 214.500 93.900 ;
        RECT 215.800 93.800 216.600 93.900 ;
        RECT 213.300 92.700 213.700 92.800 ;
        RECT 210.200 92.100 210.600 92.500 ;
        RECT 212.300 92.400 213.700 92.700 ;
        RECT 214.200 92.400 214.600 92.800 ;
        RECT 212.300 92.100 212.600 92.400 ;
        RECT 215.000 92.100 215.400 92.500 ;
        RECT 209.900 91.800 210.600 92.100 ;
        RECT 209.900 91.100 210.500 91.800 ;
        RECT 212.200 91.100 212.600 92.100 ;
        RECT 214.400 91.800 215.400 92.100 ;
        RECT 214.400 91.100 214.800 91.800 ;
        RECT 216.600 91.100 217.000 93.500 ;
        RECT 218.200 93.100 218.600 99.900 ;
        RECT 219.000 95.800 219.400 97.200 ;
        RECT 219.800 95.700 220.200 99.900 ;
        RECT 222.000 98.200 222.400 99.900 ;
        RECT 221.400 97.900 222.400 98.200 ;
        RECT 224.200 97.900 224.600 99.900 ;
        RECT 226.300 97.900 226.900 99.900 ;
        RECT 221.400 97.500 221.800 97.900 ;
        RECT 224.200 97.600 224.500 97.900 ;
        RECT 223.100 97.300 224.900 97.600 ;
        RECT 226.200 97.500 226.600 97.900 ;
        RECT 223.100 97.200 223.500 97.300 ;
        RECT 224.500 97.200 224.900 97.300 ;
        RECT 221.400 96.500 221.800 96.600 ;
        RECT 223.700 96.500 224.100 96.600 ;
        RECT 221.400 96.200 224.100 96.500 ;
        RECT 224.400 96.500 225.500 96.800 ;
        RECT 224.400 95.900 224.700 96.500 ;
        RECT 225.100 96.400 225.500 96.500 ;
        RECT 226.300 96.600 227.000 97.000 ;
        RECT 226.300 96.100 226.600 96.600 ;
        RECT 222.300 95.700 224.700 95.900 ;
        RECT 219.800 95.600 224.700 95.700 ;
        RECT 225.400 95.800 226.600 96.100 ;
        RECT 219.800 95.500 222.700 95.600 ;
        RECT 219.800 95.400 222.600 95.500 ;
        RECT 223.000 95.100 223.400 95.200 ;
        RECT 220.900 94.800 223.400 95.100 ;
        RECT 220.900 94.700 221.300 94.800 ;
        RECT 221.700 94.200 222.100 94.300 ;
        RECT 225.400 94.200 225.700 95.800 ;
        RECT 228.600 95.600 229.000 99.900 ;
        RECT 230.200 96.400 230.600 99.900 ;
        RECT 226.900 95.300 229.000 95.600 ;
        RECT 226.900 95.200 227.300 95.300 ;
        RECT 227.700 94.900 228.100 95.000 ;
        RECT 226.200 94.600 228.100 94.900 ;
        RECT 226.200 94.500 226.600 94.600 ;
        RECT 220.200 93.900 225.700 94.200 ;
        RECT 220.200 93.800 221.000 93.900 ;
        RECT 218.200 92.800 219.100 93.100 ;
        RECT 218.700 92.200 219.100 92.800 ;
        RECT 218.200 91.800 219.100 92.200 ;
        RECT 218.700 91.100 219.100 91.800 ;
        RECT 219.800 91.100 220.200 93.500 ;
        RECT 222.300 93.200 222.600 93.900 ;
        RECT 225.100 93.800 225.500 93.900 ;
        RECT 228.600 93.600 229.000 95.300 ;
        RECT 227.100 93.300 229.000 93.600 ;
        RECT 227.100 93.200 227.500 93.300 ;
        RECT 221.400 92.100 221.800 92.500 ;
        RECT 222.200 92.400 222.600 93.200 ;
        RECT 223.100 92.700 223.500 92.800 ;
        RECT 223.100 92.400 224.500 92.700 ;
        RECT 224.200 92.100 224.500 92.400 ;
        RECT 226.200 92.100 226.600 92.500 ;
        RECT 221.400 91.800 222.400 92.100 ;
        RECT 222.000 91.100 222.400 91.800 ;
        RECT 224.200 91.100 224.600 92.100 ;
        RECT 226.200 91.800 226.900 92.100 ;
        RECT 226.300 91.100 226.900 91.800 ;
        RECT 228.600 91.100 229.000 93.300 ;
        RECT 230.100 95.900 230.600 96.400 ;
        RECT 231.800 96.200 232.200 99.900 ;
        RECT 230.900 95.900 232.200 96.200 ;
        RECT 232.600 95.900 233.000 99.900 ;
        RECT 233.400 96.200 233.800 99.900 ;
        RECT 235.000 96.200 235.400 99.900 ;
        RECT 233.400 95.900 235.400 96.200 ;
        RECT 230.100 94.200 230.400 95.900 ;
        RECT 230.900 94.900 231.200 95.900 ;
        RECT 232.700 95.200 233.000 95.900 ;
        RECT 234.600 95.200 235.000 95.400 ;
        RECT 230.700 94.500 231.200 94.900 ;
        RECT 230.100 93.800 230.600 94.200 ;
        RECT 230.100 93.100 230.400 93.800 ;
        RECT 230.900 93.700 231.200 94.500 ;
        RECT 231.700 94.800 232.200 95.200 ;
        RECT 232.600 94.900 233.800 95.200 ;
        RECT 234.600 95.100 235.400 95.200 ;
        RECT 236.600 95.100 237.000 99.900 ;
        RECT 237.400 95.800 237.800 96.600 ;
        RECT 234.600 94.900 237.000 95.100 ;
        RECT 232.600 94.800 233.000 94.900 ;
        RECT 231.700 94.400 232.100 94.800 ;
        RECT 230.900 93.400 232.200 93.700 ;
        RECT 230.100 92.800 230.600 93.100 ;
        RECT 230.200 91.100 230.600 92.800 ;
        RECT 231.800 91.100 232.200 93.400 ;
        RECT 232.600 92.800 233.000 93.200 ;
        RECT 233.500 93.100 233.800 94.900 ;
        RECT 235.000 94.800 237.000 94.900 ;
        RECT 234.200 93.800 234.600 94.600 ;
        RECT 232.700 92.400 233.100 92.800 ;
        RECT 233.400 91.100 233.800 93.100 ;
        RECT 236.600 93.100 237.000 94.800 ;
        RECT 236.600 92.800 237.500 93.100 ;
        RECT 237.100 91.100 237.500 92.800 ;
        RECT 238.200 91.100 238.600 99.900 ;
        RECT 239.800 95.600 240.200 99.900 ;
        RECT 241.900 97.900 242.500 99.900 ;
        RECT 244.200 97.900 244.600 99.900 ;
        RECT 246.400 98.200 246.800 99.900 ;
        RECT 246.400 97.900 247.400 98.200 ;
        RECT 242.200 97.500 242.600 97.900 ;
        RECT 244.300 97.600 244.600 97.900 ;
        RECT 243.900 97.300 245.700 97.600 ;
        RECT 247.000 97.500 247.400 97.900 ;
        RECT 243.900 97.200 244.300 97.300 ;
        RECT 245.300 97.200 245.700 97.300 ;
        RECT 241.800 96.600 242.500 97.000 ;
        RECT 242.200 96.100 242.500 96.600 ;
        RECT 243.300 96.500 244.400 96.800 ;
        RECT 243.300 96.400 243.700 96.500 ;
        RECT 242.200 95.800 243.400 96.100 ;
        RECT 239.800 95.300 241.900 95.600 ;
        RECT 239.800 93.600 240.200 95.300 ;
        RECT 241.500 95.200 241.900 95.300 ;
        RECT 243.100 95.200 243.400 95.800 ;
        RECT 244.100 95.900 244.400 96.500 ;
        RECT 244.700 96.500 245.100 96.600 ;
        RECT 247.000 96.500 247.400 96.600 ;
        RECT 244.700 96.200 247.400 96.500 ;
        RECT 244.100 95.700 246.500 95.900 ;
        RECT 248.600 95.700 249.000 99.900 ;
        RECT 244.100 95.600 249.000 95.700 ;
        RECT 246.100 95.500 249.000 95.600 ;
        RECT 246.200 95.400 249.000 95.500 ;
        RECT 240.700 94.900 241.100 95.000 ;
        RECT 240.700 94.600 242.600 94.900 ;
        RECT 243.000 94.800 243.400 95.200 ;
        RECT 245.400 95.100 245.800 95.200 ;
        RECT 245.400 94.800 247.900 95.100 ;
        RECT 242.200 94.500 242.600 94.600 ;
        RECT 243.100 94.200 243.400 94.800 ;
        RECT 246.200 94.700 246.600 94.800 ;
        RECT 247.500 94.700 247.900 94.800 ;
        RECT 246.700 94.200 247.100 94.300 ;
        RECT 243.100 93.900 248.600 94.200 ;
        RECT 243.300 93.800 243.700 93.900 ;
        RECT 239.800 93.300 241.700 93.600 ;
        RECT 239.000 93.100 239.400 93.200 ;
        RECT 239.800 93.100 240.200 93.300 ;
        RECT 241.300 93.200 241.700 93.300 ;
        RECT 239.000 92.800 240.200 93.100 ;
        RECT 246.200 92.800 246.500 93.900 ;
        RECT 247.800 93.800 248.600 93.900 ;
        RECT 239.000 92.400 239.400 92.800 ;
        RECT 239.800 91.100 240.200 92.800 ;
        RECT 245.300 92.700 245.700 92.800 ;
        RECT 242.200 92.100 242.600 92.500 ;
        RECT 244.300 92.400 245.700 92.700 ;
        RECT 246.200 92.400 246.600 92.800 ;
        RECT 244.300 92.100 244.600 92.400 ;
        RECT 247.000 92.100 247.400 92.500 ;
        RECT 241.900 91.800 242.600 92.100 ;
        RECT 241.900 91.100 242.500 91.800 ;
        RECT 244.200 91.100 244.600 92.100 ;
        RECT 246.400 91.800 247.400 92.100 ;
        RECT 246.400 91.100 246.800 91.800 ;
        RECT 248.600 91.100 249.000 93.500 ;
        RECT 249.400 93.400 249.800 94.200 ;
        RECT 250.200 93.100 250.600 99.900 ;
        RECT 251.000 95.800 251.400 96.600 ;
        RECT 251.800 96.200 252.200 99.900 ;
        RECT 253.400 96.200 253.800 99.900 ;
        RECT 251.800 95.900 253.800 96.200 ;
        RECT 254.200 95.900 254.600 99.900 ;
        RECT 255.000 96.200 255.400 99.900 ;
        RECT 258.700 96.300 259.100 99.900 ;
        RECT 255.000 95.900 256.100 96.200 ;
        RECT 258.200 95.900 259.100 96.300 ;
        RECT 254.200 95.200 254.500 95.900 ;
        RECT 255.800 95.600 256.100 95.900 ;
        RECT 255.800 95.200 256.400 95.600 ;
        RECT 253.400 94.900 254.600 95.200 ;
        RECT 251.000 94.100 251.400 94.200 ;
        RECT 252.600 94.100 253.000 94.600 ;
        RECT 251.000 93.800 253.000 94.100 ;
        RECT 253.400 93.200 253.700 94.900 ;
        RECT 254.200 94.800 254.600 94.900 ;
        RECT 255.000 94.400 255.400 95.200 ;
        RECT 255.800 93.700 256.100 95.200 ;
        RECT 258.300 94.200 258.600 95.900 ;
        RECT 258.200 93.800 258.600 94.200 ;
        RECT 255.000 93.400 256.100 93.700 ;
        RECT 250.200 92.800 251.100 93.100 ;
        RECT 250.700 92.200 251.100 92.800 ;
        RECT 250.700 91.800 251.400 92.200 ;
        RECT 250.700 91.100 251.100 91.800 ;
        RECT 253.400 91.100 253.800 93.200 ;
        RECT 254.200 92.800 254.600 93.200 ;
        RECT 254.100 92.400 254.500 92.800 ;
        RECT 255.000 91.100 255.400 93.400 ;
        RECT 258.300 93.100 258.600 93.800 ;
        RECT 259.000 93.100 259.400 93.200 ;
        RECT 258.200 92.800 259.400 93.100 ;
        RECT 260.600 93.100 261.000 99.900 ;
        RECT 261.400 95.800 261.800 97.200 ;
        RECT 262.200 96.200 262.600 99.900 ;
        RECT 262.200 95.900 263.300 96.200 ;
        RECT 263.000 95.600 263.300 95.900 ;
        RECT 263.000 95.200 263.600 95.600 ;
        RECT 262.200 94.400 262.600 95.200 ;
        RECT 263.000 93.700 263.300 95.200 ;
        RECT 262.200 93.400 263.300 93.700 ;
        RECT 260.600 92.800 261.500 93.100 ;
        RECT 258.300 92.100 258.600 92.800 ;
        RECT 261.100 92.200 261.500 92.800 ;
        RECT 258.200 91.100 258.600 92.100 ;
        RECT 260.600 91.800 261.500 92.200 ;
        RECT 261.100 91.100 261.500 91.800 ;
        RECT 262.200 91.100 262.600 93.400 ;
        RECT 0.600 87.500 1.000 89.900 ;
        RECT 2.800 89.200 3.200 89.900 ;
        RECT 2.200 88.900 3.200 89.200 ;
        RECT 5.000 88.900 5.400 89.900 ;
        RECT 7.100 89.200 7.700 89.900 ;
        RECT 7.000 88.900 7.700 89.200 ;
        RECT 2.200 88.500 2.600 88.900 ;
        RECT 5.000 88.600 5.300 88.900 ;
        RECT 3.000 88.200 3.400 88.600 ;
        RECT 3.900 88.300 5.300 88.600 ;
        RECT 7.000 88.500 7.400 88.900 ;
        RECT 3.900 88.200 4.300 88.300 ;
        RECT 1.000 87.100 1.800 87.200 ;
        RECT 3.100 87.100 3.400 88.200 ;
        RECT 9.400 88.100 9.800 89.900 ;
        RECT 10.200 88.100 10.600 88.600 ;
        RECT 9.400 87.800 10.600 88.100 ;
        RECT 7.900 87.700 8.300 87.800 ;
        RECT 9.400 87.700 9.800 87.800 ;
        RECT 7.900 87.400 9.800 87.700 ;
        RECT 5.900 87.100 6.300 87.200 ;
        RECT 1.000 86.800 6.500 87.100 ;
        RECT 2.500 86.700 2.900 86.800 ;
        RECT 1.700 86.200 2.100 86.300 ;
        RECT 1.700 85.900 4.200 86.200 ;
        RECT 3.800 85.800 4.200 85.900 ;
        RECT 0.600 85.500 3.400 85.600 ;
        RECT 0.600 85.400 3.500 85.500 ;
        RECT 0.600 85.300 5.500 85.400 ;
        RECT 0.600 81.100 1.000 85.300 ;
        RECT 3.100 85.100 5.500 85.300 ;
        RECT 2.200 84.500 4.900 84.800 ;
        RECT 2.200 84.400 2.600 84.500 ;
        RECT 4.500 84.400 4.900 84.500 ;
        RECT 5.200 84.500 5.500 85.100 ;
        RECT 6.200 85.200 6.500 86.800 ;
        RECT 7.000 86.400 7.400 86.500 ;
        RECT 7.000 86.100 8.900 86.400 ;
        RECT 8.500 86.000 8.900 86.100 ;
        RECT 7.700 85.700 8.100 85.800 ;
        RECT 9.400 85.700 9.800 87.400 ;
        RECT 7.700 85.400 9.800 85.700 ;
        RECT 6.200 84.900 7.400 85.200 ;
        RECT 5.900 84.500 6.300 84.600 ;
        RECT 5.200 84.200 6.300 84.500 ;
        RECT 7.100 84.400 7.400 84.900 ;
        RECT 7.100 84.000 7.800 84.400 ;
        RECT 3.900 83.700 4.300 83.800 ;
        RECT 5.300 83.700 5.700 83.800 ;
        RECT 2.200 83.100 2.600 83.500 ;
        RECT 3.900 83.400 5.700 83.700 ;
        RECT 5.000 83.100 5.300 83.400 ;
        RECT 7.000 83.100 7.400 83.500 ;
        RECT 2.200 82.800 3.200 83.100 ;
        RECT 2.800 81.100 3.200 82.800 ;
        RECT 5.000 81.100 5.400 83.100 ;
        RECT 7.100 81.100 7.700 83.100 ;
        RECT 9.400 81.100 9.800 85.400 ;
        RECT 11.000 86.100 11.400 89.900 ;
        RECT 13.700 88.000 14.100 89.500 ;
        RECT 15.800 88.500 16.200 89.500 ;
        RECT 13.300 87.700 14.100 88.000 ;
        RECT 13.300 87.500 13.700 87.700 ;
        RECT 13.300 87.200 13.600 87.500 ;
        RECT 15.900 87.400 16.200 88.500 ;
        RECT 11.800 87.100 12.200 87.200 ;
        RECT 12.600 87.100 13.600 87.200 ;
        RECT 11.800 86.800 13.600 87.100 ;
        RECT 14.100 87.100 16.200 87.400 ;
        RECT 16.600 87.700 17.000 89.900 ;
        RECT 18.700 89.200 19.300 89.900 ;
        RECT 18.700 88.900 19.400 89.200 ;
        RECT 21.000 88.900 21.400 89.900 ;
        RECT 23.200 89.200 23.600 89.900 ;
        RECT 23.200 88.900 24.200 89.200 ;
        RECT 19.000 88.500 19.400 88.900 ;
        RECT 21.100 88.600 21.400 88.900 ;
        RECT 21.100 88.300 22.500 88.600 ;
        RECT 22.100 88.200 22.500 88.300 ;
        RECT 23.000 88.200 23.400 88.600 ;
        RECT 23.800 88.500 24.200 88.900 ;
        RECT 18.100 87.700 18.500 87.800 ;
        RECT 16.600 87.400 18.500 87.700 ;
        RECT 14.100 86.900 14.600 87.100 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 11.000 85.800 13.000 86.100 ;
        RECT 11.000 81.100 11.400 85.800 ;
        RECT 12.600 85.400 13.000 85.800 ;
        RECT 13.300 84.900 13.600 86.800 ;
        RECT 13.900 86.500 14.600 86.900 ;
        RECT 14.300 85.500 14.600 86.500 ;
        RECT 15.000 85.800 15.400 86.600 ;
        RECT 15.800 85.800 16.200 86.600 ;
        RECT 16.600 85.700 17.000 87.400 ;
        RECT 20.100 87.100 20.500 87.200 ;
        RECT 23.000 87.100 23.300 88.200 ;
        RECT 25.400 87.500 25.800 89.900 ;
        RECT 26.200 87.900 26.600 89.900 ;
        RECT 27.000 88.000 27.400 89.900 ;
        RECT 28.600 88.000 29.000 89.900 ;
        RECT 27.000 87.900 29.000 88.000 ;
        RECT 26.300 87.200 26.600 87.900 ;
        RECT 27.100 87.700 28.900 87.900 ;
        RECT 29.400 87.500 29.800 89.900 ;
        RECT 31.600 89.200 32.000 89.900 ;
        RECT 31.000 88.900 32.000 89.200 ;
        RECT 33.800 88.900 34.200 89.900 ;
        RECT 35.900 89.200 36.500 89.900 ;
        RECT 35.800 88.900 36.500 89.200 ;
        RECT 31.000 88.500 31.400 88.900 ;
        RECT 33.800 88.600 34.100 88.900 ;
        RECT 31.800 88.200 32.200 88.600 ;
        RECT 32.700 88.300 34.100 88.600 ;
        RECT 35.800 88.500 36.200 88.900 ;
        RECT 32.700 88.200 33.100 88.300 ;
        RECT 28.200 87.200 28.600 87.400 ;
        RECT 31.900 87.200 32.200 88.200 ;
        RECT 36.700 87.700 37.100 87.800 ;
        RECT 38.200 87.700 38.600 89.900 ;
        RECT 39.100 88.200 39.500 88.600 ;
        RECT 39.000 87.800 39.400 88.200 ;
        RECT 39.800 87.900 40.200 89.900 ;
        RECT 44.100 88.000 44.500 89.500 ;
        RECT 46.200 88.500 46.600 89.500 ;
        RECT 36.700 87.400 38.600 87.700 ;
        RECT 24.600 87.100 25.400 87.200 ;
        RECT 19.900 86.800 25.400 87.100 ;
        RECT 26.200 86.800 27.500 87.200 ;
        RECT 28.200 86.900 29.000 87.200 ;
        RECT 28.600 86.800 29.000 86.900 ;
        RECT 29.800 87.100 30.600 87.200 ;
        RECT 31.800 87.100 32.200 87.200 ;
        RECT 34.700 87.100 35.100 87.200 ;
        RECT 29.800 86.800 35.300 87.100 ;
        RECT 19.000 86.400 19.400 86.500 ;
        RECT 17.500 86.100 19.400 86.400 ;
        RECT 17.500 86.000 17.900 86.100 ;
        RECT 18.300 85.700 18.700 85.800 ;
        RECT 14.300 85.200 16.200 85.500 ;
        RECT 13.300 84.600 14.100 84.900 ;
        RECT 13.700 81.100 14.100 84.600 ;
        RECT 15.900 83.500 16.200 85.200 ;
        RECT 15.800 81.500 16.200 83.500 ;
        RECT 16.600 85.400 18.700 85.700 ;
        RECT 16.600 81.100 17.000 85.400 ;
        RECT 19.900 85.200 20.200 86.800 ;
        RECT 23.500 86.700 23.900 86.800 ;
        RECT 24.300 86.200 24.700 86.300 ;
        RECT 22.200 85.900 24.700 86.200 ;
        RECT 22.200 85.800 22.600 85.900 ;
        RECT 23.000 85.500 25.800 85.600 ;
        RECT 22.900 85.400 25.800 85.500 ;
        RECT 19.000 84.900 20.200 85.200 ;
        RECT 20.900 85.300 25.800 85.400 ;
        RECT 20.900 85.100 23.300 85.300 ;
        RECT 19.000 84.400 19.300 84.900 ;
        RECT 18.600 84.000 19.300 84.400 ;
        RECT 20.100 84.500 20.500 84.600 ;
        RECT 20.900 84.500 21.200 85.100 ;
        RECT 20.100 84.200 21.200 84.500 ;
        RECT 21.500 84.500 24.200 84.800 ;
        RECT 21.500 84.400 21.900 84.500 ;
        RECT 23.800 84.400 24.200 84.500 ;
        RECT 20.700 83.700 21.100 83.800 ;
        RECT 22.100 83.700 22.500 83.800 ;
        RECT 19.000 83.100 19.400 83.500 ;
        RECT 20.700 83.400 22.500 83.700 ;
        RECT 21.100 83.100 21.400 83.400 ;
        RECT 23.800 83.100 24.200 83.500 ;
        RECT 18.700 81.100 19.300 83.100 ;
        RECT 21.000 81.100 21.400 83.100 ;
        RECT 23.200 82.800 24.200 83.100 ;
        RECT 23.200 81.100 23.600 82.800 ;
        RECT 25.400 81.100 25.800 85.300 ;
        RECT 26.200 85.100 26.600 85.200 ;
        RECT 27.200 85.100 27.500 86.800 ;
        RECT 31.300 86.700 31.700 86.800 ;
        RECT 27.800 85.800 28.200 86.600 ;
        RECT 30.500 86.200 30.900 86.300 ;
        RECT 30.500 86.100 33.000 86.200 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 30.500 85.900 33.800 86.100 ;
        RECT 32.600 85.800 33.800 85.900 ;
        RECT 29.400 85.500 32.200 85.600 ;
        RECT 29.400 85.400 32.300 85.500 ;
        RECT 29.400 85.300 34.300 85.400 ;
        RECT 26.200 84.800 26.900 85.100 ;
        RECT 27.200 84.800 27.700 85.100 ;
        RECT 26.600 84.200 26.900 84.800 ;
        RECT 26.600 83.800 27.000 84.200 ;
        RECT 27.300 81.100 27.700 84.800 ;
        RECT 29.400 81.100 29.800 85.300 ;
        RECT 31.900 85.100 34.300 85.300 ;
        RECT 31.000 84.500 33.700 84.800 ;
        RECT 31.000 84.400 31.400 84.500 ;
        RECT 33.300 84.400 33.700 84.500 ;
        RECT 34.000 84.500 34.300 85.100 ;
        RECT 35.000 85.200 35.300 86.800 ;
        RECT 35.800 86.400 36.200 86.500 ;
        RECT 35.800 86.100 37.700 86.400 ;
        RECT 37.300 86.000 37.700 86.100 ;
        RECT 36.500 85.700 36.900 85.800 ;
        RECT 38.200 85.700 38.600 87.400 ;
        RECT 39.000 86.100 39.400 86.200 ;
        RECT 39.900 86.100 40.200 87.900 ;
        RECT 43.700 87.700 44.500 88.000 ;
        RECT 43.700 87.500 44.100 87.700 ;
        RECT 43.700 87.200 44.000 87.500 ;
        RECT 46.300 87.400 46.600 88.500 ;
        RECT 40.600 86.400 41.000 87.200 ;
        RECT 43.000 86.800 44.000 87.200 ;
        RECT 44.500 87.100 46.600 87.400 ;
        RECT 47.000 88.500 47.400 89.500 ;
        RECT 49.100 89.200 49.500 89.500 ;
        RECT 49.100 88.800 49.800 89.200 ;
        RECT 47.000 87.400 47.300 88.500 ;
        RECT 49.100 88.000 49.500 88.800 ;
        RECT 53.700 88.000 54.100 89.500 ;
        RECT 55.800 88.500 56.200 89.500 ;
        RECT 49.100 87.700 49.900 88.000 ;
        RECT 49.500 87.500 49.900 87.700 ;
        RECT 47.000 87.100 49.100 87.400 ;
        RECT 44.500 86.900 45.000 87.100 ;
        RECT 41.400 86.100 41.800 86.200 ;
        RECT 39.000 85.800 40.200 86.100 ;
        RECT 41.000 85.800 41.800 86.100 ;
        RECT 42.200 86.100 42.600 86.200 ;
        RECT 43.000 86.100 43.400 86.200 ;
        RECT 42.200 85.800 43.400 86.100 ;
        RECT 36.500 85.400 38.600 85.700 ;
        RECT 35.000 84.900 36.200 85.200 ;
        RECT 34.700 84.500 35.100 84.600 ;
        RECT 34.000 84.200 35.100 84.500 ;
        RECT 35.900 84.400 36.200 84.900 ;
        RECT 35.900 84.000 36.600 84.400 ;
        RECT 32.700 83.700 33.100 83.800 ;
        RECT 34.100 83.700 34.500 83.800 ;
        RECT 31.000 83.100 31.400 83.500 ;
        RECT 32.700 83.400 34.500 83.700 ;
        RECT 33.800 83.100 34.100 83.400 ;
        RECT 35.800 83.100 36.200 83.500 ;
        RECT 31.000 82.800 32.000 83.100 ;
        RECT 31.600 81.100 32.000 82.800 ;
        RECT 33.800 81.100 34.200 83.100 ;
        RECT 35.900 81.100 36.500 83.100 ;
        RECT 38.200 81.100 38.600 85.400 ;
        RECT 39.100 85.100 39.400 85.800 ;
        RECT 41.000 85.600 41.400 85.800 ;
        RECT 43.000 85.400 43.400 85.800 ;
        RECT 43.700 85.200 44.000 86.800 ;
        RECT 44.300 86.500 45.000 86.900 ;
        RECT 48.600 86.900 49.100 87.100 ;
        RECT 49.600 87.200 49.900 87.500 ;
        RECT 53.300 87.700 54.100 88.000 ;
        RECT 53.300 87.500 53.700 87.700 ;
        RECT 53.300 87.200 53.600 87.500 ;
        RECT 55.900 87.400 56.200 88.500 ;
        RECT 59.500 89.200 59.900 89.900 ;
        RECT 59.500 88.800 60.200 89.200 ;
        RECT 59.500 88.200 59.900 88.800 ;
        RECT 59.000 87.900 59.900 88.200 ;
        RECT 44.700 85.500 45.000 86.500 ;
        RECT 45.400 85.800 45.800 86.600 ;
        RECT 46.200 85.800 46.600 86.600 ;
        RECT 47.000 85.800 47.400 86.600 ;
        RECT 47.800 85.800 48.200 86.600 ;
        RECT 48.600 86.500 49.300 86.900 ;
        RECT 49.600 86.800 50.600 87.200 ;
        RECT 52.600 87.100 53.600 87.200 ;
        RECT 51.000 86.800 53.600 87.100 ;
        RECT 54.100 87.100 56.200 87.400 ;
        RECT 57.400 87.100 57.800 87.200 ;
        RECT 58.200 87.100 58.600 87.600 ;
        RECT 54.100 86.900 54.600 87.100 ;
        RECT 48.600 85.500 48.900 86.500 ;
        RECT 44.700 85.200 46.600 85.500 ;
        RECT 39.000 81.100 39.400 85.100 ;
        RECT 39.800 84.800 41.800 85.100 ;
        RECT 39.800 81.100 40.200 84.800 ;
        RECT 41.400 81.100 41.800 84.800 ;
        RECT 43.700 84.900 44.200 85.200 ;
        RECT 43.700 84.600 44.500 84.900 ;
        RECT 44.100 81.100 44.500 84.600 ;
        RECT 46.300 83.500 46.600 85.200 ;
        RECT 46.200 81.500 46.600 83.500 ;
        RECT 47.000 85.200 48.900 85.500 ;
        RECT 47.000 83.500 47.300 85.200 ;
        RECT 49.600 84.900 49.900 86.800 ;
        RECT 50.200 86.100 50.600 86.200 ;
        RECT 51.000 86.100 51.300 86.800 ;
        RECT 50.200 85.800 51.300 86.100 ;
        RECT 50.200 85.400 50.600 85.800 ;
        RECT 52.600 85.400 53.000 86.200 ;
        RECT 49.100 84.600 49.900 84.900 ;
        RECT 53.300 84.900 53.600 86.800 ;
        RECT 53.900 86.500 54.600 86.900 ;
        RECT 57.400 86.800 58.600 87.100 ;
        RECT 54.300 85.500 54.600 86.500 ;
        RECT 55.000 85.800 55.400 86.600 ;
        RECT 55.800 86.100 56.200 86.600 ;
        RECT 56.600 86.100 57.000 86.200 ;
        RECT 55.800 85.800 57.000 86.100 ;
        RECT 54.300 85.200 56.200 85.500 ;
        RECT 53.300 84.600 54.100 84.900 ;
        RECT 47.000 81.500 47.400 83.500 ;
        RECT 49.100 81.100 49.500 84.600 ;
        RECT 53.700 81.100 54.100 84.600 ;
        RECT 55.900 83.500 56.200 85.200 ;
        RECT 55.800 81.500 56.200 83.500 ;
        RECT 59.000 81.100 59.400 87.900 ;
        RECT 60.600 87.700 61.000 89.900 ;
        RECT 62.700 89.200 63.300 89.900 ;
        RECT 62.700 88.900 63.400 89.200 ;
        RECT 65.000 88.900 65.400 89.900 ;
        RECT 67.200 89.200 67.600 89.900 ;
        RECT 67.200 88.900 68.200 89.200 ;
        RECT 63.000 88.500 63.400 88.900 ;
        RECT 65.100 88.600 65.400 88.900 ;
        RECT 65.100 88.300 66.500 88.600 ;
        RECT 66.100 88.200 66.500 88.300 ;
        RECT 67.000 88.200 67.400 88.600 ;
        RECT 67.800 88.500 68.200 88.900 ;
        RECT 62.100 87.700 62.500 87.800 ;
        RECT 60.600 87.400 62.500 87.700 ;
        RECT 60.600 85.700 61.000 87.400 ;
        RECT 64.100 87.100 64.500 87.200 ;
        RECT 67.000 87.100 67.300 88.200 ;
        RECT 69.400 87.500 69.800 89.900 ;
        RECT 70.500 88.200 70.900 89.900 ;
        RECT 70.500 87.900 71.400 88.200 ;
        RECT 72.600 87.900 73.000 89.900 ;
        RECT 73.400 88.000 73.800 89.900 ;
        RECT 75.000 88.000 75.400 89.900 ;
        RECT 73.400 87.900 75.400 88.000 ;
        RECT 77.100 87.900 77.900 89.900 ;
        RECT 81.700 89.200 82.100 89.500 ;
        RECT 81.700 88.800 82.600 89.200 ;
        RECT 81.700 88.000 82.100 88.800 ;
        RECT 83.800 88.500 84.200 89.500 ;
        RECT 68.600 87.100 69.400 87.200 ;
        RECT 63.900 86.800 69.400 87.100 ;
        RECT 63.000 86.400 63.400 86.500 ;
        RECT 61.500 86.100 63.400 86.400 ;
        RECT 63.900 86.200 64.200 86.800 ;
        RECT 67.500 86.700 67.900 86.800 ;
        RECT 67.000 86.200 67.400 86.300 ;
        RECT 68.300 86.200 68.700 86.300 ;
        RECT 61.500 86.000 61.900 86.100 ;
        RECT 63.800 85.800 64.200 86.200 ;
        RECT 66.200 85.900 68.700 86.200 ;
        RECT 66.200 85.800 66.600 85.900 ;
        RECT 62.300 85.700 62.700 85.800 ;
        RECT 60.600 85.400 62.700 85.700 ;
        RECT 59.800 84.400 60.200 85.200 ;
        RECT 60.600 81.100 61.000 85.400 ;
        RECT 63.900 85.200 64.200 85.800 ;
        RECT 67.000 85.500 69.800 85.600 ;
        RECT 66.900 85.400 69.800 85.500 ;
        RECT 63.000 84.900 64.200 85.200 ;
        RECT 64.900 85.300 69.800 85.400 ;
        RECT 64.900 85.100 67.300 85.300 ;
        RECT 63.000 84.400 63.300 84.900 ;
        RECT 62.600 84.000 63.300 84.400 ;
        RECT 64.100 84.500 64.500 84.600 ;
        RECT 64.900 84.500 65.200 85.100 ;
        RECT 64.100 84.200 65.200 84.500 ;
        RECT 65.500 84.500 68.200 84.800 ;
        RECT 65.500 84.400 65.900 84.500 ;
        RECT 67.800 84.400 68.200 84.500 ;
        RECT 64.700 83.700 65.100 83.800 ;
        RECT 66.100 83.700 66.500 83.800 ;
        RECT 63.000 83.100 63.400 83.500 ;
        RECT 64.700 83.400 66.500 83.700 ;
        RECT 65.100 83.100 65.400 83.400 ;
        RECT 67.800 83.100 68.200 83.500 ;
        RECT 62.700 81.100 63.300 83.100 ;
        RECT 65.000 81.100 65.400 83.100 ;
        RECT 67.200 82.800 68.200 83.100 ;
        RECT 67.200 81.100 67.600 82.800 ;
        RECT 69.400 81.100 69.800 85.300 ;
        RECT 70.200 84.400 70.600 85.200 ;
        RECT 71.000 85.100 71.400 87.900 ;
        RECT 71.800 86.800 72.200 87.600 ;
        RECT 72.700 87.200 73.000 87.900 ;
        RECT 73.500 87.700 75.300 87.900 ;
        RECT 74.600 87.200 75.000 87.400 ;
        RECT 72.600 86.800 73.900 87.200 ;
        RECT 74.600 86.900 75.400 87.200 ;
        RECT 75.000 86.800 75.400 86.900 ;
        RECT 76.600 86.800 77.000 87.200 ;
        RECT 72.600 85.100 73.000 85.200 ;
        RECT 73.600 85.100 73.900 86.800 ;
        RECT 76.700 86.600 77.000 86.800 ;
        RECT 74.200 85.800 74.600 86.600 ;
        RECT 76.700 86.200 77.100 86.600 ;
        RECT 77.400 86.200 77.700 87.900 ;
        RECT 81.300 87.700 82.100 88.000 ;
        RECT 81.300 87.500 81.700 87.700 ;
        RECT 81.300 87.200 81.600 87.500 ;
        RECT 83.900 87.400 84.200 88.500 ;
        RECT 78.200 86.400 78.600 87.200 ;
        RECT 80.600 86.800 81.600 87.200 ;
        RECT 82.100 87.100 84.200 87.400 ;
        RECT 85.400 87.600 85.800 89.900 ;
        RECT 87.000 87.600 87.400 89.900 ;
        RECT 88.600 87.600 89.000 89.900 ;
        RECT 90.200 87.600 90.600 89.900 ;
        RECT 91.800 87.800 92.200 88.600 ;
        RECT 85.400 87.200 86.300 87.600 ;
        RECT 87.000 87.200 88.100 87.600 ;
        RECT 88.600 87.200 89.700 87.600 ;
        RECT 90.200 87.200 91.400 87.600 ;
        RECT 82.100 86.900 82.600 87.100 ;
        RECT 75.800 85.400 76.200 86.200 ;
        RECT 77.400 85.800 77.800 86.200 ;
        RECT 79.000 86.100 79.400 86.200 ;
        RECT 78.600 85.800 79.400 86.100 ;
        RECT 79.800 86.100 80.200 86.200 ;
        RECT 80.600 86.100 81.000 86.200 ;
        RECT 79.800 85.800 81.000 86.100 ;
        RECT 77.400 85.700 77.700 85.800 ;
        RECT 76.700 85.400 77.700 85.700 ;
        RECT 78.600 85.600 79.000 85.800 ;
        RECT 80.600 85.400 81.000 85.800 ;
        RECT 76.700 85.100 77.000 85.400 ;
        RECT 71.000 84.800 73.300 85.100 ;
        RECT 73.600 84.800 74.100 85.100 ;
        RECT 71.000 81.100 71.400 84.800 ;
        RECT 73.000 84.200 73.300 84.800 ;
        RECT 73.000 83.800 73.400 84.200 ;
        RECT 73.700 81.100 74.100 84.800 ;
        RECT 75.800 81.400 76.200 85.100 ;
        RECT 76.600 81.700 77.000 85.100 ;
        RECT 77.400 84.800 79.400 85.100 ;
        RECT 77.400 81.400 77.800 84.800 ;
        RECT 75.800 81.100 77.800 81.400 ;
        RECT 79.000 81.100 79.400 84.800 ;
        RECT 81.300 84.900 81.600 86.800 ;
        RECT 81.900 86.500 82.600 86.900 ;
        RECT 85.900 86.900 86.300 87.200 ;
        RECT 87.700 86.900 88.100 87.200 ;
        RECT 89.300 86.900 89.700 87.200 ;
        RECT 82.300 85.500 82.600 86.500 ;
        RECT 83.000 85.800 83.400 86.600 ;
        RECT 83.800 85.800 84.200 86.600 ;
        RECT 85.900 86.500 87.200 86.900 ;
        RECT 87.700 86.500 88.900 86.900 ;
        RECT 89.300 86.500 90.600 86.900 ;
        RECT 85.900 85.800 86.300 86.500 ;
        RECT 87.700 85.800 88.100 86.500 ;
        RECT 89.300 85.800 89.700 86.500 ;
        RECT 91.000 85.800 91.400 87.200 ;
        RECT 82.300 85.200 84.200 85.500 ;
        RECT 81.300 84.600 82.100 84.900 ;
        RECT 81.700 81.100 82.100 84.600 ;
        RECT 83.900 83.500 84.200 85.200 ;
        RECT 83.800 81.500 84.200 83.500 ;
        RECT 85.400 85.400 86.300 85.800 ;
        RECT 87.000 85.400 88.100 85.800 ;
        RECT 88.600 85.400 89.700 85.800 ;
        RECT 90.200 85.400 91.400 85.800 ;
        RECT 85.400 81.100 85.800 85.400 ;
        RECT 87.000 81.100 87.400 85.400 ;
        RECT 88.600 81.100 89.000 85.400 ;
        RECT 90.200 81.100 90.600 85.400 ;
        RECT 91.800 85.100 92.200 85.200 ;
        RECT 92.600 85.100 93.000 89.900 ;
        RECT 91.800 84.800 93.000 85.100 ;
        RECT 92.600 81.100 93.000 84.800 ;
        RECT 93.400 87.700 93.800 89.900 ;
        RECT 95.500 89.200 96.100 89.900 ;
        RECT 95.500 88.900 96.200 89.200 ;
        RECT 97.800 88.900 98.200 89.900 ;
        RECT 100.000 89.200 100.400 89.900 ;
        RECT 100.000 88.900 101.000 89.200 ;
        RECT 95.800 88.500 96.200 88.900 ;
        RECT 97.900 88.600 98.200 88.900 ;
        RECT 97.900 88.300 99.300 88.600 ;
        RECT 98.900 88.200 99.300 88.300 ;
        RECT 99.800 88.200 100.200 88.600 ;
        RECT 100.600 88.500 101.000 88.900 ;
        RECT 94.900 87.700 95.300 87.800 ;
        RECT 93.400 87.400 95.300 87.700 ;
        RECT 93.400 85.700 93.800 87.400 ;
        RECT 96.900 87.100 97.300 87.200 ;
        RECT 99.000 87.100 99.400 87.200 ;
        RECT 99.800 87.100 100.100 88.200 ;
        RECT 102.200 87.500 102.600 89.900 ;
        RECT 103.000 88.500 103.400 89.500 ;
        RECT 103.000 87.400 103.300 88.500 ;
        RECT 105.100 88.200 105.500 89.500 ;
        RECT 104.600 88.000 105.500 88.200 ;
        RECT 104.600 87.800 105.900 88.000 ;
        RECT 105.100 87.700 105.900 87.800 ;
        RECT 105.500 87.500 105.900 87.700 ;
        RECT 109.400 87.500 109.800 89.900 ;
        RECT 111.600 89.200 112.000 89.900 ;
        RECT 111.000 88.900 112.000 89.200 ;
        RECT 113.800 88.900 114.200 89.900 ;
        RECT 115.900 89.200 116.500 89.900 ;
        RECT 115.800 88.900 116.500 89.200 ;
        RECT 111.000 88.500 111.400 88.900 ;
        RECT 113.800 88.600 114.100 88.900 ;
        RECT 111.800 88.200 112.200 88.600 ;
        RECT 112.700 88.300 114.100 88.600 ;
        RECT 115.800 88.500 116.200 88.900 ;
        RECT 112.700 88.200 113.100 88.300 ;
        RECT 101.400 87.100 102.200 87.200 ;
        RECT 103.000 87.100 105.100 87.400 ;
        RECT 96.700 86.800 102.200 87.100 ;
        RECT 104.600 86.900 105.100 87.100 ;
        RECT 105.600 87.200 105.900 87.500 ;
        RECT 95.800 86.400 96.200 86.500 ;
        RECT 94.300 86.100 96.200 86.400 ;
        RECT 94.300 86.000 94.700 86.100 ;
        RECT 95.100 85.700 95.500 85.800 ;
        RECT 93.400 85.400 95.500 85.700 ;
        RECT 93.400 81.100 93.800 85.400 ;
        RECT 96.700 85.200 97.000 86.800 ;
        RECT 100.300 86.700 100.700 86.800 ;
        RECT 99.800 86.200 100.200 86.300 ;
        RECT 101.100 86.200 101.500 86.300 ;
        RECT 99.000 85.900 101.500 86.200 ;
        RECT 99.000 85.800 99.400 85.900 ;
        RECT 103.000 85.800 103.400 86.600 ;
        RECT 103.800 85.800 104.200 86.600 ;
        RECT 104.600 86.500 105.300 86.900 ;
        RECT 105.600 86.800 106.600 87.200 ;
        RECT 109.800 87.100 110.600 87.200 ;
        RECT 111.900 87.100 112.200 88.200 ;
        RECT 118.200 88.100 118.600 89.900 ;
        RECT 119.000 88.100 119.400 88.600 ;
        RECT 118.200 87.800 119.400 88.100 ;
        RECT 116.700 87.700 117.100 87.800 ;
        RECT 118.200 87.700 118.600 87.800 ;
        RECT 116.700 87.400 118.600 87.700 ;
        RECT 114.700 87.100 115.100 87.200 ;
        RECT 109.800 86.800 115.300 87.100 ;
        RECT 99.800 85.500 102.600 85.600 ;
        RECT 104.600 85.500 104.900 86.500 ;
        RECT 99.700 85.400 102.600 85.500 ;
        RECT 95.800 84.900 97.000 85.200 ;
        RECT 97.700 85.300 102.600 85.400 ;
        RECT 97.700 85.100 100.100 85.300 ;
        RECT 95.800 84.400 96.100 84.900 ;
        RECT 95.400 84.000 96.100 84.400 ;
        RECT 96.900 84.500 97.300 84.600 ;
        RECT 97.700 84.500 98.000 85.100 ;
        RECT 96.900 84.200 98.000 84.500 ;
        RECT 98.300 84.500 101.000 84.800 ;
        RECT 98.300 84.400 98.700 84.500 ;
        RECT 100.600 84.400 101.000 84.500 ;
        RECT 97.500 83.700 97.900 83.800 ;
        RECT 98.900 83.700 99.300 83.800 ;
        RECT 95.800 83.100 96.200 83.500 ;
        RECT 97.500 83.400 99.300 83.700 ;
        RECT 97.900 83.100 98.200 83.400 ;
        RECT 100.600 83.100 101.000 83.500 ;
        RECT 95.500 81.100 96.100 83.100 ;
        RECT 97.800 81.100 98.200 83.100 ;
        RECT 100.000 82.800 101.000 83.100 ;
        RECT 100.000 81.100 100.400 82.800 ;
        RECT 102.200 81.100 102.600 85.300 ;
        RECT 103.000 85.200 104.900 85.500 ;
        RECT 103.000 83.500 103.300 85.200 ;
        RECT 105.600 84.900 105.900 86.800 ;
        RECT 111.300 86.700 111.700 86.800 ;
        RECT 110.500 86.200 110.900 86.300 ;
        RECT 106.200 85.400 106.600 86.200 ;
        RECT 110.500 85.900 113.000 86.200 ;
        RECT 112.600 85.800 113.000 85.900 ;
        RECT 109.400 85.500 112.200 85.600 ;
        RECT 109.400 85.400 112.300 85.500 ;
        RECT 105.100 84.600 105.900 84.900 ;
        RECT 109.400 85.300 114.300 85.400 ;
        RECT 103.000 81.500 103.400 83.500 ;
        RECT 105.100 81.100 105.500 84.600 ;
        RECT 109.400 81.100 109.800 85.300 ;
        RECT 111.900 85.100 114.300 85.300 ;
        RECT 111.000 84.500 113.700 84.800 ;
        RECT 111.000 84.400 111.400 84.500 ;
        RECT 113.300 84.400 113.700 84.500 ;
        RECT 114.000 84.500 114.300 85.100 ;
        RECT 115.000 85.200 115.300 86.800 ;
        RECT 115.800 86.400 116.200 86.500 ;
        RECT 115.800 86.100 117.700 86.400 ;
        RECT 117.300 86.000 117.700 86.100 ;
        RECT 116.500 85.700 116.900 85.800 ;
        RECT 118.200 85.700 118.600 87.400 ;
        RECT 116.500 85.400 118.600 85.700 ;
        RECT 115.000 84.900 116.200 85.200 ;
        RECT 114.700 84.500 115.100 84.600 ;
        RECT 114.000 84.200 115.100 84.500 ;
        RECT 115.900 84.400 116.200 84.900 ;
        RECT 115.900 84.000 116.600 84.400 ;
        RECT 112.700 83.700 113.100 83.800 ;
        RECT 114.100 83.700 114.500 83.800 ;
        RECT 111.000 83.100 111.400 83.500 ;
        RECT 112.700 83.400 114.500 83.700 ;
        RECT 113.800 83.100 114.100 83.400 ;
        RECT 115.800 83.100 116.200 83.500 ;
        RECT 111.000 82.800 112.000 83.100 ;
        RECT 111.600 81.100 112.000 82.800 ;
        RECT 113.800 81.100 114.200 83.100 ;
        RECT 115.900 81.100 116.500 83.100 ;
        RECT 118.200 81.100 118.600 85.400 ;
        RECT 119.800 86.100 120.200 89.900 ;
        RECT 122.500 88.000 122.900 89.500 ;
        RECT 124.600 88.500 125.000 89.500 ;
        RECT 122.100 87.700 122.900 88.000 ;
        RECT 122.100 87.500 122.500 87.700 ;
        RECT 122.100 87.200 122.400 87.500 ;
        RECT 124.700 87.400 125.000 88.500 ;
        RECT 125.400 87.500 125.800 89.900 ;
        RECT 127.600 89.200 128.000 89.900 ;
        RECT 127.000 88.900 128.000 89.200 ;
        RECT 129.800 88.900 130.200 89.900 ;
        RECT 131.900 89.200 132.500 89.900 ;
        RECT 131.800 88.900 132.500 89.200 ;
        RECT 127.000 88.500 127.400 88.900 ;
        RECT 129.800 88.600 130.100 88.900 ;
        RECT 127.800 87.800 128.200 88.600 ;
        RECT 128.700 88.300 130.100 88.600 ;
        RECT 131.800 88.500 132.200 88.900 ;
        RECT 128.700 88.200 129.100 88.300 ;
        RECT 134.200 88.100 134.600 89.900 ;
        RECT 135.000 88.100 135.400 88.600 ;
        RECT 134.200 87.800 135.400 88.100 ;
        RECT 120.600 87.100 121.000 87.200 ;
        RECT 121.400 87.100 122.400 87.200 ;
        RECT 120.600 86.800 122.400 87.100 ;
        RECT 122.900 87.100 125.000 87.400 ;
        RECT 125.800 87.100 126.600 87.200 ;
        RECT 127.900 87.100 128.200 87.800 ;
        RECT 132.700 87.700 133.100 87.800 ;
        RECT 134.200 87.700 134.600 87.800 ;
        RECT 132.700 87.400 134.600 87.700 ;
        RECT 130.700 87.100 131.100 87.200 ;
        RECT 122.900 86.900 123.400 87.100 ;
        RECT 121.400 86.100 121.800 86.200 ;
        RECT 119.800 85.800 121.800 86.100 ;
        RECT 119.800 81.100 120.200 85.800 ;
        RECT 121.400 85.400 121.800 85.800 ;
        RECT 122.100 84.900 122.400 86.800 ;
        RECT 122.700 86.500 123.400 86.900 ;
        RECT 125.800 86.800 131.300 87.100 ;
        RECT 127.300 86.700 127.700 86.800 ;
        RECT 123.100 85.500 123.400 86.500 ;
        RECT 123.800 85.800 124.200 86.600 ;
        RECT 124.600 85.800 125.000 86.600 ;
        RECT 126.500 86.200 126.900 86.300 ;
        RECT 126.500 85.900 129.000 86.200 ;
        RECT 128.600 85.800 129.000 85.900 ;
        RECT 125.400 85.500 128.200 85.600 ;
        RECT 123.100 85.200 125.000 85.500 ;
        RECT 122.100 84.600 122.900 84.900 ;
        RECT 122.500 81.100 122.900 84.600 ;
        RECT 124.700 83.500 125.000 85.200 ;
        RECT 124.600 81.500 125.000 83.500 ;
        RECT 125.400 85.400 128.300 85.500 ;
        RECT 125.400 85.300 130.300 85.400 ;
        RECT 125.400 81.100 125.800 85.300 ;
        RECT 127.900 85.100 130.300 85.300 ;
        RECT 127.000 84.500 129.700 84.800 ;
        RECT 127.000 84.400 127.400 84.500 ;
        RECT 129.300 84.400 129.700 84.500 ;
        RECT 130.000 84.500 130.300 85.100 ;
        RECT 131.000 85.200 131.300 86.800 ;
        RECT 131.800 86.400 132.200 86.500 ;
        RECT 131.800 86.100 133.700 86.400 ;
        RECT 133.300 86.000 133.700 86.100 ;
        RECT 132.500 85.700 132.900 85.800 ;
        RECT 134.200 85.700 134.600 87.400 ;
        RECT 135.000 87.200 135.300 87.800 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 132.500 85.400 134.600 85.700 ;
        RECT 131.000 84.900 132.200 85.200 ;
        RECT 130.700 84.500 131.100 84.600 ;
        RECT 130.000 84.200 131.100 84.500 ;
        RECT 131.900 84.400 132.200 84.900 ;
        RECT 131.900 84.000 132.600 84.400 ;
        RECT 128.700 83.700 129.100 83.800 ;
        RECT 130.100 83.700 130.500 83.800 ;
        RECT 127.000 83.100 127.400 83.500 ;
        RECT 128.700 83.400 130.500 83.700 ;
        RECT 129.800 83.100 130.100 83.400 ;
        RECT 131.800 83.100 132.200 83.500 ;
        RECT 127.000 82.800 128.000 83.100 ;
        RECT 127.600 81.100 128.000 82.800 ;
        RECT 129.800 81.100 130.200 83.100 ;
        RECT 131.900 81.100 132.500 83.100 ;
        RECT 134.200 81.100 134.600 85.400 ;
        RECT 135.800 86.100 136.200 89.900 ;
        RECT 138.500 88.000 138.900 89.500 ;
        RECT 140.600 88.500 141.000 89.500 ;
        RECT 138.100 87.700 138.900 88.000 ;
        RECT 138.100 87.500 138.500 87.700 ;
        RECT 138.100 87.200 138.400 87.500 ;
        RECT 140.700 87.400 141.000 88.500 ;
        RECT 143.300 88.000 143.700 89.500 ;
        RECT 145.400 88.500 145.800 89.500 ;
        RECT 136.600 87.100 137.000 87.200 ;
        RECT 137.400 87.100 138.400 87.200 ;
        RECT 136.600 86.800 138.400 87.100 ;
        RECT 138.900 87.100 141.000 87.400 ;
        RECT 142.900 87.700 143.700 88.000 ;
        RECT 142.900 87.500 143.300 87.700 ;
        RECT 142.900 87.200 143.200 87.500 ;
        RECT 145.500 87.400 145.800 88.500 ;
        RECT 146.200 87.900 146.600 89.900 ;
        RECT 148.300 89.200 148.700 89.900 ;
        RECT 148.300 88.800 149.000 89.200 ;
        RECT 148.300 88.400 148.700 88.800 ;
        RECT 148.300 87.900 149.000 88.400 ;
        RECT 146.300 87.800 146.600 87.900 ;
        RECT 146.300 87.600 147.200 87.800 ;
        RECT 146.300 87.500 148.400 87.600 ;
        RECT 138.900 86.900 139.400 87.100 ;
        RECT 137.400 86.100 137.800 86.200 ;
        RECT 135.800 85.800 137.800 86.100 ;
        RECT 135.800 81.100 136.200 85.800 ;
        RECT 137.400 85.400 137.800 85.800 ;
        RECT 138.100 84.900 138.400 86.800 ;
        RECT 138.700 86.500 139.400 86.900 ;
        RECT 142.200 86.800 143.200 87.200 ;
        RECT 143.700 87.100 145.800 87.400 ;
        RECT 146.900 87.300 148.400 87.500 ;
        RECT 148.000 87.200 148.400 87.300 ;
        RECT 143.700 86.900 144.200 87.100 ;
        RECT 139.100 85.500 139.400 86.500 ;
        RECT 139.800 85.800 140.200 86.600 ;
        RECT 140.600 86.100 141.000 86.600 ;
        RECT 141.400 86.100 141.800 86.200 ;
        RECT 140.600 85.800 141.800 86.100 ;
        RECT 139.100 85.200 141.000 85.500 ;
        RECT 142.200 85.400 142.600 86.200 ;
        RECT 138.100 84.600 138.900 84.900 ;
        RECT 138.500 81.100 138.900 84.600 ;
        RECT 140.700 83.500 141.000 85.200 ;
        RECT 142.900 84.900 143.200 86.800 ;
        RECT 143.500 86.500 144.200 86.900 ;
        RECT 143.900 85.500 144.200 86.500 ;
        RECT 144.600 85.800 145.000 86.600 ;
        RECT 145.400 85.800 145.800 86.600 ;
        RECT 146.200 86.400 146.600 87.200 ;
        RECT 147.200 86.900 147.600 87.000 ;
        RECT 147.100 86.600 147.600 86.900 ;
        RECT 147.100 86.200 147.400 86.600 ;
        RECT 147.000 85.800 147.400 86.200 ;
        RECT 148.000 85.500 148.300 87.200 ;
        RECT 148.700 86.200 149.000 87.900 ;
        RECT 149.400 86.800 149.800 87.600 ;
        RECT 148.600 85.800 149.000 86.200 ;
        RECT 143.900 85.200 145.800 85.500 ;
        RECT 142.900 84.600 143.700 84.900 ;
        RECT 140.600 81.500 141.000 83.500 ;
        RECT 143.300 82.200 143.700 84.600 ;
        RECT 145.500 83.500 145.800 85.200 ;
        RECT 143.000 81.800 143.700 82.200 ;
        RECT 143.300 81.100 143.700 81.800 ;
        RECT 145.400 81.500 145.800 83.500 ;
        RECT 147.100 85.200 148.300 85.500 ;
        RECT 147.100 83.100 147.400 85.200 ;
        RECT 148.700 85.100 149.000 85.800 ;
        RECT 147.000 81.100 147.400 83.100 ;
        RECT 148.600 81.100 149.000 85.100 ;
        RECT 150.200 81.100 150.600 89.900 ;
        RECT 151.000 87.700 151.400 89.900 ;
        RECT 153.100 89.200 153.700 89.900 ;
        RECT 153.100 88.900 153.800 89.200 ;
        RECT 155.400 88.900 155.800 89.900 ;
        RECT 157.600 89.200 158.000 89.900 ;
        RECT 157.600 88.900 158.600 89.200 ;
        RECT 153.400 88.500 153.800 88.900 ;
        RECT 155.500 88.600 155.800 88.900 ;
        RECT 155.500 88.300 156.900 88.600 ;
        RECT 156.500 88.200 156.900 88.300 ;
        RECT 157.400 88.200 157.800 88.600 ;
        RECT 158.200 88.500 158.600 88.900 ;
        RECT 152.500 87.700 152.900 87.800 ;
        RECT 151.000 87.400 152.900 87.700 ;
        RECT 151.000 85.700 151.400 87.400 ;
        RECT 154.500 87.100 154.900 87.200 ;
        RECT 157.400 87.100 157.700 88.200 ;
        RECT 159.800 87.500 160.200 89.900 ;
        RECT 161.400 87.800 161.800 88.200 ;
        RECT 162.200 87.900 162.600 89.900 ;
        RECT 163.000 88.000 163.400 89.900 ;
        RECT 164.600 88.000 165.000 89.900 ;
        RECT 167.300 89.200 167.700 89.500 ;
        RECT 167.300 88.800 168.200 89.200 ;
        RECT 167.300 88.000 167.700 88.800 ;
        RECT 169.400 88.500 169.800 89.500 ;
        RECT 163.000 87.900 165.000 88.000 ;
        RECT 159.000 87.100 159.800 87.200 ;
        RECT 154.300 86.800 159.800 87.100 ;
        RECT 161.400 87.100 161.700 87.800 ;
        RECT 162.300 87.200 162.600 87.900 ;
        RECT 163.100 87.700 164.900 87.900 ;
        RECT 166.900 87.700 167.700 88.000 ;
        RECT 166.900 87.500 167.300 87.700 ;
        RECT 164.200 87.200 164.600 87.400 ;
        RECT 166.900 87.200 167.200 87.500 ;
        RECT 169.500 87.400 169.800 88.500 ;
        RECT 170.200 87.500 170.600 89.900 ;
        RECT 172.400 89.200 172.800 89.900 ;
        RECT 171.800 88.900 172.800 89.200 ;
        RECT 174.600 88.900 175.000 89.900 ;
        RECT 176.700 89.200 177.300 89.900 ;
        RECT 176.600 88.900 177.300 89.200 ;
        RECT 171.800 88.500 172.200 88.900 ;
        RECT 174.600 88.600 174.900 88.900 ;
        RECT 172.600 88.200 173.000 88.600 ;
        RECT 173.500 88.300 174.900 88.600 ;
        RECT 176.600 88.500 177.000 88.900 ;
        RECT 173.500 88.200 173.900 88.300 ;
        RECT 162.200 87.100 163.500 87.200 ;
        RECT 161.400 86.800 163.500 87.100 ;
        RECT 164.200 86.900 165.000 87.200 ;
        RECT 164.600 86.800 165.000 86.900 ;
        RECT 166.200 86.800 167.200 87.200 ;
        RECT 167.700 87.100 169.800 87.400 ;
        RECT 170.600 87.100 171.400 87.200 ;
        RECT 172.700 87.100 173.000 88.200 ;
        RECT 177.500 87.700 177.900 87.800 ;
        RECT 179.000 87.700 179.400 89.900 ;
        RECT 179.800 87.900 180.200 89.900 ;
        RECT 180.600 88.000 181.000 89.900 ;
        RECT 182.200 88.000 182.600 89.900 ;
        RECT 180.600 87.900 182.600 88.000 ;
        RECT 183.000 87.900 183.400 89.900 ;
        RECT 183.800 88.000 184.200 89.900 ;
        RECT 185.400 88.000 185.800 89.900 ;
        RECT 183.800 87.900 185.800 88.000 ;
        RECT 186.200 88.000 186.600 89.900 ;
        RECT 187.800 88.000 188.200 89.900 ;
        RECT 186.200 87.900 188.200 88.000 ;
        RECT 177.500 87.400 179.400 87.700 ;
        RECT 173.400 87.100 173.800 87.200 ;
        RECT 175.500 87.100 175.900 87.200 ;
        RECT 167.700 86.900 168.200 87.100 ;
        RECT 153.400 86.400 153.800 86.500 ;
        RECT 151.900 86.100 153.800 86.400 ;
        RECT 154.300 86.200 154.600 86.800 ;
        RECT 157.900 86.700 158.300 86.800 ;
        RECT 157.400 86.200 157.800 86.300 ;
        RECT 158.700 86.200 159.100 86.300 ;
        RECT 151.900 86.000 152.300 86.100 ;
        RECT 154.200 85.800 154.600 86.200 ;
        RECT 156.600 85.900 159.100 86.200 ;
        RECT 156.600 85.800 157.000 85.900 ;
        RECT 152.700 85.700 153.100 85.800 ;
        RECT 151.000 85.400 153.100 85.700 ;
        RECT 151.000 81.100 151.400 85.400 ;
        RECT 154.300 85.200 154.600 85.800 ;
        RECT 157.400 85.500 160.200 85.600 ;
        RECT 157.300 85.400 160.200 85.500 ;
        RECT 153.400 84.900 154.600 85.200 ;
        RECT 155.300 85.300 160.200 85.400 ;
        RECT 155.300 85.100 157.700 85.300 ;
        RECT 153.400 84.400 153.700 84.900 ;
        RECT 153.000 84.000 153.700 84.400 ;
        RECT 154.500 84.500 154.900 84.600 ;
        RECT 155.300 84.500 155.600 85.100 ;
        RECT 154.500 84.200 155.600 84.500 ;
        RECT 155.900 84.500 158.600 84.800 ;
        RECT 155.900 84.400 156.300 84.500 ;
        RECT 158.200 84.400 158.600 84.500 ;
        RECT 155.100 83.700 155.500 83.800 ;
        RECT 156.500 83.700 156.900 83.800 ;
        RECT 153.400 83.100 153.800 83.500 ;
        RECT 155.100 83.400 156.900 83.700 ;
        RECT 155.500 83.100 155.800 83.400 ;
        RECT 158.200 83.100 158.600 83.500 ;
        RECT 153.100 81.100 153.700 83.100 ;
        RECT 155.400 81.100 155.800 83.100 ;
        RECT 157.600 82.800 158.600 83.100 ;
        RECT 157.600 81.100 158.000 82.800 ;
        RECT 159.800 81.100 160.200 85.300 ;
        RECT 160.600 85.100 161.000 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 163.200 85.100 163.500 86.800 ;
        RECT 163.800 85.800 164.200 86.600 ;
        RECT 164.600 86.100 165.000 86.200 ;
        RECT 166.200 86.100 166.600 86.200 ;
        RECT 164.600 85.800 166.600 86.100 ;
        RECT 166.200 85.400 166.600 85.800 ;
        RECT 160.600 84.800 162.900 85.100 ;
        RECT 163.200 84.800 163.700 85.100 ;
        RECT 162.600 84.200 162.900 84.800 ;
        RECT 162.600 83.800 163.000 84.200 ;
        RECT 163.300 81.100 163.700 84.800 ;
        RECT 166.900 84.900 167.200 86.800 ;
        RECT 167.500 86.500 168.200 86.900 ;
        RECT 170.600 86.800 176.100 87.100 ;
        RECT 172.100 86.700 172.500 86.800 ;
        RECT 167.900 85.500 168.200 86.500 ;
        RECT 168.600 85.800 169.000 86.600 ;
        RECT 169.400 85.800 169.800 86.600 ;
        RECT 171.300 86.200 171.700 86.300 ;
        RECT 171.300 86.100 173.800 86.200 ;
        RECT 175.000 86.100 175.400 86.200 ;
        RECT 171.300 85.900 175.400 86.100 ;
        RECT 173.400 85.800 175.400 85.900 ;
        RECT 170.200 85.500 173.000 85.600 ;
        RECT 167.900 85.200 169.800 85.500 ;
        RECT 166.900 84.600 167.700 84.900 ;
        RECT 167.300 81.100 167.700 84.600 ;
        RECT 169.500 83.500 169.800 85.200 ;
        RECT 169.400 81.500 169.800 83.500 ;
        RECT 170.200 85.400 173.100 85.500 ;
        RECT 170.200 85.300 175.100 85.400 ;
        RECT 170.200 81.100 170.600 85.300 ;
        RECT 172.700 85.100 175.100 85.300 ;
        RECT 171.800 84.500 174.500 84.800 ;
        RECT 171.800 84.400 172.200 84.500 ;
        RECT 174.100 84.400 174.500 84.500 ;
        RECT 174.800 84.500 175.100 85.100 ;
        RECT 175.800 85.200 176.100 86.800 ;
        RECT 176.600 86.400 177.000 86.500 ;
        RECT 176.600 86.100 178.500 86.400 ;
        RECT 178.100 86.000 178.500 86.100 ;
        RECT 177.300 85.700 177.700 85.800 ;
        RECT 179.000 85.700 179.400 87.400 ;
        RECT 179.900 87.200 180.200 87.900 ;
        RECT 180.700 87.700 182.500 87.900 ;
        RECT 181.800 87.200 182.200 87.400 ;
        RECT 183.100 87.200 183.400 87.900 ;
        RECT 183.900 87.700 185.700 87.900 ;
        RECT 186.300 87.700 188.100 87.900 ;
        RECT 188.600 87.800 189.000 89.900 ;
        RECT 185.000 87.200 185.400 87.400 ;
        RECT 186.600 87.200 187.000 87.400 ;
        RECT 188.600 87.200 188.900 87.800 ;
        RECT 189.400 87.700 189.800 89.900 ;
        RECT 191.500 89.200 192.100 89.900 ;
        RECT 191.500 88.900 192.200 89.200 ;
        RECT 193.800 88.900 194.200 89.900 ;
        RECT 196.000 89.200 196.400 89.900 ;
        RECT 196.000 88.900 197.000 89.200 ;
        RECT 191.800 88.500 192.200 88.900 ;
        RECT 193.900 88.600 194.200 88.900 ;
        RECT 193.900 88.300 195.300 88.600 ;
        RECT 194.900 88.200 195.300 88.300 ;
        RECT 195.800 88.200 196.200 88.600 ;
        RECT 196.600 88.500 197.000 88.900 ;
        RECT 190.900 87.700 191.300 87.800 ;
        RECT 189.400 87.400 191.300 87.700 ;
        RECT 179.800 86.800 181.100 87.200 ;
        RECT 181.800 86.900 182.600 87.200 ;
        RECT 182.200 86.800 182.600 86.900 ;
        RECT 183.000 86.800 184.300 87.200 ;
        RECT 185.000 86.900 185.800 87.200 ;
        RECT 185.400 86.800 185.800 86.900 ;
        RECT 186.200 86.900 187.000 87.200 ;
        RECT 186.200 86.800 186.600 86.900 ;
        RECT 187.700 86.800 189.000 87.200 ;
        RECT 177.300 85.400 179.400 85.700 ;
        RECT 175.800 84.900 177.000 85.200 ;
        RECT 175.500 84.500 175.900 84.600 ;
        RECT 174.800 84.200 175.900 84.500 ;
        RECT 176.700 84.400 177.000 84.900 ;
        RECT 179.000 85.100 179.400 85.400 ;
        RECT 179.800 85.100 180.200 85.200 ;
        RECT 180.800 85.100 181.100 86.800 ;
        RECT 181.400 86.100 181.800 86.600 ;
        RECT 182.200 86.100 182.600 86.200 ;
        RECT 181.400 85.800 182.600 86.100 ;
        RECT 183.000 85.100 183.400 85.200 ;
        RECT 184.000 85.100 184.300 86.800 ;
        RECT 184.600 86.100 185.000 86.600 ;
        RECT 186.200 86.100 186.500 86.800 ;
        RECT 184.600 85.800 186.500 86.100 ;
        RECT 187.000 85.800 187.400 86.600 ;
        RECT 187.700 85.100 188.000 86.800 ;
        RECT 189.400 85.700 189.800 87.400 ;
        RECT 192.900 87.100 193.300 87.200 ;
        RECT 195.800 87.100 196.100 88.200 ;
        RECT 198.200 87.500 198.600 89.900 ;
        RECT 199.800 87.600 200.200 89.900 ;
        RECT 201.400 87.600 201.800 89.900 ;
        RECT 203.000 87.600 203.400 89.900 ;
        RECT 204.600 87.600 205.000 89.900 ;
        RECT 207.000 87.600 207.400 89.900 ;
        RECT 208.600 87.600 209.000 89.900 ;
        RECT 211.800 87.900 212.200 89.900 ;
        RECT 212.600 88.000 213.000 89.900 ;
        RECT 214.200 88.000 214.600 89.900 ;
        RECT 212.600 87.900 214.600 88.000 ;
        RECT 215.000 87.900 215.400 89.900 ;
        RECT 215.800 88.000 216.200 89.900 ;
        RECT 217.400 88.000 217.800 89.900 ;
        RECT 215.800 87.900 217.800 88.000 ;
        RECT 219.800 87.900 220.200 89.900 ;
        RECT 220.500 88.200 220.900 88.600 ;
        RECT 199.000 87.200 200.200 87.600 ;
        RECT 200.700 87.200 201.800 87.600 ;
        RECT 202.300 87.200 203.400 87.600 ;
        RECT 204.100 87.200 205.000 87.600 ;
        RECT 197.400 87.100 198.200 87.200 ;
        RECT 192.700 86.800 198.200 87.100 ;
        RECT 191.800 86.400 192.200 86.500 ;
        RECT 190.300 86.100 192.200 86.400 ;
        RECT 190.300 86.000 190.700 86.100 ;
        RECT 191.100 85.700 191.500 85.800 ;
        RECT 189.400 85.400 191.500 85.700 ;
        RECT 188.600 85.100 189.000 85.200 ;
        RECT 179.000 84.800 180.500 85.100 ;
        RECT 180.800 84.800 181.300 85.100 ;
        RECT 183.000 84.800 183.700 85.100 ;
        RECT 184.000 84.800 184.500 85.100 ;
        RECT 176.700 84.000 177.400 84.400 ;
        RECT 173.500 83.700 173.900 83.800 ;
        RECT 174.900 83.700 175.300 83.800 ;
        RECT 171.800 83.100 172.200 83.500 ;
        RECT 173.500 83.400 175.300 83.700 ;
        RECT 174.600 83.100 174.900 83.400 ;
        RECT 176.600 83.100 177.000 83.500 ;
        RECT 171.800 82.800 172.800 83.100 ;
        RECT 172.400 81.100 172.800 82.800 ;
        RECT 174.600 81.100 175.000 83.100 ;
        RECT 176.700 81.100 177.300 83.100 ;
        RECT 179.000 81.100 179.400 84.800 ;
        RECT 180.200 84.200 180.500 84.800 ;
        RECT 180.900 84.200 181.300 84.800 ;
        RECT 183.400 84.200 183.700 84.800 ;
        RECT 180.200 83.800 180.600 84.200 ;
        RECT 180.900 83.800 181.800 84.200 ;
        RECT 183.400 83.800 183.800 84.200 ;
        RECT 180.900 81.100 181.300 83.800 ;
        RECT 184.100 81.100 184.500 84.800 ;
        RECT 187.500 84.800 188.000 85.100 ;
        RECT 188.300 84.800 189.000 85.100 ;
        RECT 187.500 81.100 187.900 84.800 ;
        RECT 188.300 84.200 188.600 84.800 ;
        RECT 188.200 83.800 188.600 84.200 ;
        RECT 189.400 81.100 189.800 85.400 ;
        RECT 192.700 85.200 193.000 86.800 ;
        RECT 196.300 86.700 196.700 86.800 ;
        RECT 197.100 86.200 197.500 86.300 ;
        RECT 195.000 85.900 197.500 86.200 ;
        RECT 195.000 85.800 195.400 85.900 ;
        RECT 199.000 85.800 199.400 87.200 ;
        RECT 200.700 86.900 201.100 87.200 ;
        RECT 202.300 86.900 202.700 87.200 ;
        RECT 204.100 86.900 204.500 87.200 ;
        RECT 205.400 86.900 205.800 87.200 ;
        RECT 199.800 86.500 201.100 86.900 ;
        RECT 201.500 86.500 202.700 86.900 ;
        RECT 203.200 86.500 204.500 86.900 ;
        RECT 204.900 86.500 205.800 86.900 ;
        RECT 206.200 86.800 206.600 87.600 ;
        RECT 207.000 87.200 209.000 87.600 ;
        RECT 211.900 87.200 212.200 87.900 ;
        RECT 212.700 87.700 214.500 87.900 ;
        RECT 213.800 87.200 214.200 87.400 ;
        RECT 215.100 87.200 215.400 87.900 ;
        RECT 215.900 87.700 217.700 87.900 ;
        RECT 217.000 87.200 217.400 87.400 ;
        RECT 200.700 85.800 201.100 86.500 ;
        RECT 202.300 85.800 202.700 86.500 ;
        RECT 204.100 85.800 204.500 86.500 ;
        RECT 205.400 86.100 205.800 86.200 ;
        RECT 205.400 85.800 207.400 86.100 ;
        RECT 208.600 85.800 209.000 87.200 ;
        RECT 211.800 86.800 213.100 87.200 ;
        RECT 213.800 86.900 214.600 87.200 ;
        RECT 214.200 86.800 214.600 86.900 ;
        RECT 215.000 86.800 216.300 87.200 ;
        RECT 217.000 86.900 217.800 87.200 ;
        RECT 217.400 86.800 217.800 86.900 ;
        RECT 195.800 85.500 198.600 85.600 ;
        RECT 195.700 85.400 198.600 85.500 ;
        RECT 199.000 85.400 200.200 85.800 ;
        RECT 200.700 85.400 201.800 85.800 ;
        RECT 202.300 85.400 203.400 85.800 ;
        RECT 204.100 85.400 205.000 85.800 ;
        RECT 191.800 84.900 193.000 85.200 ;
        RECT 193.700 85.300 198.600 85.400 ;
        RECT 193.700 85.100 196.100 85.300 ;
        RECT 191.800 84.400 192.100 84.900 ;
        RECT 191.400 84.000 192.100 84.400 ;
        RECT 192.900 84.500 193.300 84.600 ;
        RECT 193.700 84.500 194.000 85.100 ;
        RECT 192.900 84.200 194.000 84.500 ;
        RECT 194.300 84.500 197.000 84.800 ;
        RECT 194.300 84.400 194.700 84.500 ;
        RECT 196.600 84.400 197.000 84.500 ;
        RECT 193.500 83.700 193.900 83.800 ;
        RECT 194.900 83.700 195.300 83.800 ;
        RECT 191.800 83.100 192.200 83.500 ;
        RECT 193.500 83.400 195.300 83.700 ;
        RECT 193.900 83.100 194.200 83.400 ;
        RECT 196.600 83.100 197.000 83.500 ;
        RECT 191.500 81.100 192.100 83.100 ;
        RECT 193.800 81.100 194.200 83.100 ;
        RECT 196.000 82.800 197.000 83.100 ;
        RECT 196.000 81.100 196.400 82.800 ;
        RECT 198.200 81.100 198.600 85.300 ;
        RECT 199.800 81.100 200.200 85.400 ;
        RECT 201.400 81.100 201.800 85.400 ;
        RECT 203.000 81.100 203.400 85.400 ;
        RECT 204.600 81.100 205.000 85.400 ;
        RECT 207.000 85.400 209.000 85.800 ;
        RECT 207.000 81.100 207.400 85.400 ;
        RECT 208.600 81.100 209.000 85.400 ;
        RECT 211.800 85.100 212.200 85.200 ;
        RECT 212.800 85.100 213.100 86.800 ;
        RECT 213.400 85.800 213.800 86.600 ;
        RECT 215.000 85.100 215.400 85.200 ;
        RECT 216.000 85.100 216.300 86.800 ;
        RECT 216.600 85.800 217.000 86.600 ;
        RECT 219.000 86.400 219.400 87.200 ;
        RECT 218.200 86.100 218.600 86.200 ;
        RECT 219.800 86.100 220.100 87.900 ;
        RECT 220.600 87.800 221.000 88.200 ;
        RECT 221.400 87.900 221.800 89.900 ;
        RECT 222.200 88.000 222.600 89.900 ;
        RECT 223.800 88.000 224.200 89.900 ;
        RECT 225.400 88.200 225.800 89.900 ;
        RECT 222.200 87.900 224.200 88.000 ;
        RECT 225.300 87.900 225.800 88.200 ;
        RECT 221.500 87.200 221.800 87.900 ;
        RECT 222.300 87.700 224.100 87.900 ;
        RECT 223.400 87.200 223.800 87.400 ;
        RECT 225.300 87.200 225.600 87.900 ;
        RECT 227.000 87.600 227.400 89.900 ;
        RECT 227.800 88.000 228.200 89.900 ;
        RECT 229.400 88.000 229.800 89.900 ;
        RECT 227.800 87.900 229.800 88.000 ;
        RECT 230.200 87.900 230.600 89.900 ;
        RECT 227.900 87.700 229.700 87.900 ;
        RECT 226.100 87.300 227.400 87.600 ;
        RECT 221.400 86.800 222.700 87.200 ;
        RECT 223.400 86.900 224.200 87.200 ;
        RECT 223.800 86.800 224.200 86.900 ;
        RECT 225.300 86.800 225.800 87.200 ;
        RECT 220.600 86.100 221.000 86.200 ;
        RECT 218.200 85.800 219.000 86.100 ;
        RECT 219.800 85.800 221.000 86.100 ;
        RECT 218.600 85.600 219.000 85.800 ;
        RECT 220.600 85.100 220.900 85.800 ;
        RECT 221.400 85.100 221.800 85.200 ;
        RECT 222.400 85.100 222.700 86.800 ;
        RECT 223.000 85.800 223.400 86.600 ;
        RECT 225.300 85.100 225.600 86.800 ;
        RECT 226.100 86.500 226.400 87.300 ;
        RECT 228.200 87.200 228.600 87.400 ;
        RECT 230.200 87.200 230.500 87.900 ;
        RECT 231.000 87.500 231.400 89.900 ;
        RECT 233.200 89.200 233.600 89.900 ;
        RECT 232.600 88.900 233.600 89.200 ;
        RECT 235.400 88.900 235.800 89.900 ;
        RECT 237.500 89.200 238.100 89.900 ;
        RECT 237.400 88.900 238.100 89.200 ;
        RECT 232.600 88.500 233.000 88.900 ;
        RECT 235.400 88.600 235.700 88.900 ;
        RECT 233.400 88.200 233.800 88.600 ;
        RECT 234.300 88.300 235.700 88.600 ;
        RECT 237.400 88.500 237.800 88.900 ;
        RECT 234.300 88.200 234.700 88.300 ;
        RECT 227.800 86.900 228.600 87.200 ;
        RECT 227.800 86.800 228.200 86.900 ;
        RECT 229.300 86.800 230.600 87.200 ;
        RECT 231.400 87.100 232.200 87.200 ;
        RECT 233.500 87.100 233.800 88.200 ;
        RECT 238.300 87.700 238.700 87.800 ;
        RECT 239.800 87.700 240.200 89.900 ;
        RECT 238.300 87.400 240.200 87.700 ;
        RECT 241.400 87.600 241.800 89.900 ;
        RECT 243.000 87.600 243.400 89.900 ;
        RECT 244.600 87.600 245.000 89.900 ;
        RECT 246.200 87.600 246.600 89.900 ;
        RECT 236.300 87.100 236.700 87.200 ;
        RECT 231.400 86.800 236.900 87.100 ;
        RECT 225.900 86.100 226.400 86.500 ;
        RECT 226.100 85.100 226.400 86.100 ;
        RECT 226.900 86.200 227.300 86.600 ;
        RECT 226.900 85.800 227.400 86.200 ;
        RECT 228.600 85.800 229.000 86.600 ;
        RECT 229.300 86.200 229.600 86.800 ;
        RECT 232.900 86.700 233.300 86.800 ;
        RECT 232.100 86.200 232.500 86.300 ;
        RECT 233.400 86.200 233.800 86.300 ;
        RECT 229.300 85.800 229.800 86.200 ;
        RECT 232.100 85.900 234.600 86.200 ;
        RECT 234.200 85.800 234.600 85.900 ;
        RECT 229.300 85.100 229.600 85.800 ;
        RECT 231.000 85.500 233.800 85.600 ;
        RECT 231.000 85.400 233.900 85.500 ;
        RECT 231.000 85.300 235.900 85.400 ;
        RECT 230.200 85.100 230.600 85.200 ;
        RECT 211.800 84.800 212.500 85.100 ;
        RECT 212.800 84.800 213.300 85.100 ;
        RECT 215.000 84.800 215.700 85.100 ;
        RECT 216.000 84.800 216.500 85.100 ;
        RECT 212.200 84.200 212.500 84.800 ;
        RECT 212.900 84.200 213.300 84.800 ;
        RECT 215.400 84.200 215.700 84.800 ;
        RECT 212.200 83.800 212.600 84.200 ;
        RECT 212.900 83.800 213.800 84.200 ;
        RECT 215.400 83.800 215.800 84.200 ;
        RECT 212.900 81.100 213.300 83.800 ;
        RECT 216.100 81.100 216.500 84.800 ;
        RECT 218.200 84.800 220.200 85.100 ;
        RECT 218.200 81.100 218.600 84.800 ;
        RECT 219.800 81.100 220.200 84.800 ;
        RECT 220.600 81.100 221.000 85.100 ;
        RECT 221.400 84.800 222.100 85.100 ;
        RECT 222.400 84.800 222.900 85.100 ;
        RECT 221.800 84.200 222.100 84.800 ;
        RECT 221.800 83.800 222.200 84.200 ;
        RECT 222.500 82.200 222.900 84.800 ;
        RECT 225.300 84.600 225.800 85.100 ;
        RECT 226.100 84.800 227.400 85.100 ;
        RECT 222.500 81.800 223.400 82.200 ;
        RECT 222.500 81.100 222.900 81.800 ;
        RECT 225.400 81.100 225.800 84.600 ;
        RECT 227.000 81.100 227.400 84.800 ;
        RECT 229.100 84.800 229.600 85.100 ;
        RECT 229.900 84.800 230.600 85.100 ;
        RECT 229.100 81.100 229.500 84.800 ;
        RECT 229.900 84.200 230.200 84.800 ;
        RECT 229.800 83.800 230.200 84.200 ;
        RECT 231.000 81.100 231.400 85.300 ;
        RECT 233.500 85.100 235.900 85.300 ;
        RECT 232.600 84.500 235.300 84.800 ;
        RECT 232.600 84.400 233.000 84.500 ;
        RECT 234.900 84.400 235.300 84.500 ;
        RECT 235.600 84.500 235.900 85.100 ;
        RECT 236.600 85.200 236.900 86.800 ;
        RECT 237.400 86.400 237.800 86.500 ;
        RECT 237.400 86.100 239.300 86.400 ;
        RECT 238.900 86.000 239.300 86.100 ;
        RECT 238.100 85.700 238.500 85.800 ;
        RECT 239.800 85.700 240.200 87.400 ;
        RECT 238.100 85.400 240.200 85.700 ;
        RECT 240.600 87.200 241.800 87.600 ;
        RECT 242.300 87.200 243.400 87.600 ;
        RECT 243.900 87.200 245.000 87.600 ;
        RECT 245.700 87.200 246.600 87.600 ;
        RECT 248.600 87.600 249.000 89.900 ;
        RECT 250.200 87.600 250.600 89.900 ;
        RECT 251.800 87.600 252.200 89.900 ;
        RECT 253.400 87.600 253.800 89.900 ;
        RECT 255.100 88.200 255.500 88.600 ;
        RECT 255.000 87.800 255.400 88.200 ;
        RECT 255.800 87.900 256.200 89.900 ;
        RECT 248.600 87.200 249.500 87.600 ;
        RECT 250.200 87.200 251.300 87.600 ;
        RECT 251.800 87.200 252.900 87.600 ;
        RECT 253.400 87.200 254.600 87.600 ;
        RECT 240.600 85.800 241.000 87.200 ;
        RECT 242.300 86.900 242.700 87.200 ;
        RECT 243.900 86.900 244.300 87.200 ;
        RECT 245.700 86.900 246.100 87.200 ;
        RECT 247.000 86.900 247.400 87.200 ;
        RECT 241.400 86.500 242.700 86.900 ;
        RECT 243.100 86.500 244.300 86.900 ;
        RECT 244.800 86.500 246.100 86.900 ;
        RECT 246.500 86.500 247.400 86.900 ;
        RECT 249.100 86.900 249.500 87.200 ;
        RECT 250.900 86.900 251.300 87.200 ;
        RECT 252.500 86.900 252.900 87.200 ;
        RECT 249.100 86.500 250.400 86.900 ;
        RECT 250.900 86.500 252.100 86.900 ;
        RECT 252.500 86.500 253.800 86.900 ;
        RECT 242.300 85.800 242.700 86.500 ;
        RECT 243.900 85.800 244.300 86.500 ;
        RECT 245.700 85.800 246.100 86.500 ;
        RECT 249.100 85.800 249.500 86.500 ;
        RECT 250.900 85.800 251.300 86.500 ;
        RECT 252.500 85.800 252.900 86.500 ;
        RECT 254.200 85.800 254.600 87.200 ;
        RECT 255.000 86.100 255.400 86.200 ;
        RECT 255.900 86.100 256.200 87.900 ;
        RECT 259.000 87.600 259.400 89.900 ;
        RECT 260.600 87.600 261.000 89.900 ;
        RECT 262.200 87.600 262.600 89.900 ;
        RECT 263.800 87.600 264.200 89.900 ;
        RECT 259.000 87.200 259.900 87.600 ;
        RECT 260.600 87.200 261.700 87.600 ;
        RECT 262.200 87.200 263.300 87.600 ;
        RECT 263.800 87.200 265.000 87.600 ;
        RECT 256.600 86.400 257.000 87.200 ;
        RECT 258.200 86.900 258.600 87.200 ;
        RECT 259.500 86.900 259.900 87.200 ;
        RECT 261.300 86.900 261.700 87.200 ;
        RECT 262.900 86.900 263.300 87.200 ;
        RECT 258.200 86.500 259.100 86.900 ;
        RECT 259.500 86.500 260.800 86.900 ;
        RECT 261.300 86.500 262.500 86.900 ;
        RECT 262.900 86.500 264.200 86.900 ;
        RECT 257.400 86.100 257.800 86.200 ;
        RECT 255.000 85.800 256.200 86.100 ;
        RECT 257.000 85.800 257.800 86.100 ;
        RECT 259.500 85.800 259.900 86.500 ;
        RECT 261.300 85.800 261.700 86.500 ;
        RECT 262.900 85.800 263.300 86.500 ;
        RECT 264.600 85.800 265.000 87.200 ;
        RECT 240.600 85.400 241.800 85.800 ;
        RECT 242.300 85.400 243.400 85.800 ;
        RECT 243.900 85.400 245.000 85.800 ;
        RECT 245.700 85.400 246.600 85.800 ;
        RECT 236.600 84.900 237.800 85.200 ;
        RECT 236.300 84.500 236.700 84.600 ;
        RECT 235.600 84.200 236.700 84.500 ;
        RECT 237.500 84.400 237.800 84.900 ;
        RECT 237.500 84.200 238.200 84.400 ;
        RECT 237.500 84.000 238.600 84.200 ;
        RECT 237.900 83.800 238.600 84.000 ;
        RECT 234.300 83.700 234.700 83.800 ;
        RECT 235.700 83.700 236.100 83.800 ;
        RECT 232.600 83.100 233.000 83.500 ;
        RECT 234.300 83.400 236.100 83.700 ;
        RECT 235.400 83.100 235.700 83.400 ;
        RECT 237.400 83.100 237.800 83.500 ;
        RECT 232.600 82.800 233.600 83.100 ;
        RECT 233.200 81.100 233.600 82.800 ;
        RECT 235.400 81.100 235.800 83.100 ;
        RECT 237.500 81.100 238.100 83.100 ;
        RECT 239.800 81.100 240.200 85.400 ;
        RECT 241.400 81.100 241.800 85.400 ;
        RECT 243.000 81.100 243.400 85.400 ;
        RECT 244.600 81.100 245.000 85.400 ;
        RECT 246.200 81.100 246.600 85.400 ;
        RECT 248.600 85.400 249.500 85.800 ;
        RECT 250.200 85.400 251.300 85.800 ;
        RECT 251.800 85.400 252.900 85.800 ;
        RECT 253.400 85.400 254.600 85.800 ;
        RECT 248.600 81.100 249.000 85.400 ;
        RECT 250.200 81.100 250.600 85.400 ;
        RECT 251.800 81.100 252.200 85.400 ;
        RECT 253.400 81.100 253.800 85.400 ;
        RECT 255.100 85.100 255.400 85.800 ;
        RECT 257.000 85.600 257.400 85.800 ;
        RECT 259.000 85.400 259.900 85.800 ;
        RECT 260.600 85.400 261.700 85.800 ;
        RECT 262.200 85.400 263.300 85.800 ;
        RECT 263.800 85.400 265.000 85.800 ;
        RECT 255.000 81.100 255.400 85.100 ;
        RECT 255.800 84.800 257.800 85.100 ;
        RECT 255.800 81.100 256.200 84.800 ;
        RECT 257.400 81.100 257.800 84.800 ;
        RECT 259.000 81.100 259.400 85.400 ;
        RECT 260.600 81.100 261.000 85.400 ;
        RECT 262.200 81.100 262.600 85.400 ;
        RECT 263.800 81.100 264.200 85.400 ;
        RECT 0.600 75.700 1.000 79.900 ;
        RECT 2.800 78.200 3.200 79.900 ;
        RECT 2.200 77.900 3.200 78.200 ;
        RECT 5.000 77.900 5.400 79.900 ;
        RECT 7.100 77.900 7.700 79.900 ;
        RECT 2.200 77.500 2.600 77.900 ;
        RECT 5.000 77.600 5.300 77.900 ;
        RECT 3.900 77.300 5.700 77.600 ;
        RECT 7.000 77.500 7.400 77.900 ;
        RECT 3.900 77.200 4.300 77.300 ;
        RECT 5.300 77.200 5.700 77.300 ;
        RECT 9.400 77.100 9.800 79.900 ;
        RECT 10.200 77.100 10.600 77.200 ;
        RECT 2.200 76.500 2.600 76.600 ;
        RECT 4.500 76.500 4.900 76.600 ;
        RECT 2.200 76.200 4.900 76.500 ;
        RECT 5.200 76.500 6.300 76.800 ;
        RECT 5.200 75.900 5.500 76.500 ;
        RECT 5.900 76.400 6.300 76.500 ;
        RECT 7.100 76.600 7.800 77.000 ;
        RECT 9.400 76.800 10.600 77.100 ;
        RECT 7.100 76.100 7.400 76.600 ;
        RECT 3.100 75.700 5.500 75.900 ;
        RECT 0.600 75.600 5.500 75.700 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 0.600 75.500 3.500 75.600 ;
        RECT 0.600 75.400 3.400 75.500 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 1.700 74.800 4.200 75.100 ;
        RECT 1.700 74.700 2.100 74.800 ;
        RECT 2.500 74.200 2.900 74.300 ;
        RECT 6.200 74.200 6.500 75.800 ;
        RECT 9.400 75.600 9.800 76.800 ;
        RECT 7.700 75.300 9.800 75.600 ;
        RECT 7.700 75.200 8.100 75.300 ;
        RECT 8.500 74.900 8.900 75.000 ;
        RECT 7.000 74.600 8.900 74.900 ;
        RECT 7.000 74.500 7.400 74.600 ;
        RECT 1.000 73.900 6.500 74.200 ;
        RECT 1.000 73.800 1.800 73.900 ;
        RECT 0.600 71.100 1.000 73.500 ;
        RECT 3.100 72.800 3.400 73.900 ;
        RECT 5.900 73.800 6.300 73.900 ;
        RECT 9.400 73.600 9.800 75.300 ;
        RECT 11.000 75.100 11.400 79.900 ;
        RECT 13.000 76.800 13.400 77.200 ;
        RECT 11.800 75.800 12.200 76.600 ;
        RECT 13.000 76.200 13.300 76.800 ;
        RECT 13.700 76.200 14.100 79.900 ;
        RECT 12.600 75.900 13.300 76.200 ;
        RECT 13.600 75.900 14.100 76.200 ;
        RECT 12.600 75.800 13.000 75.900 ;
        RECT 12.600 75.100 12.900 75.800 ;
        RECT 11.000 74.800 12.900 75.100 ;
        RECT 7.900 73.300 9.800 73.600 ;
        RECT 10.200 73.400 10.600 74.200 ;
        RECT 7.900 73.200 8.300 73.300 ;
        RECT 2.200 72.100 2.600 72.500 ;
        RECT 3.000 72.400 3.400 72.800 ;
        RECT 3.900 72.700 4.300 72.800 ;
        RECT 3.900 72.400 5.300 72.700 ;
        RECT 5.000 72.100 5.300 72.400 ;
        RECT 7.000 72.100 7.400 72.500 ;
        RECT 2.200 71.800 3.200 72.100 ;
        RECT 2.800 71.100 3.200 71.800 ;
        RECT 5.000 71.100 5.400 72.100 ;
        RECT 7.000 71.800 7.700 72.100 ;
        RECT 7.100 71.100 7.700 71.800 ;
        RECT 9.400 71.100 9.800 73.300 ;
        RECT 11.000 73.100 11.400 74.800 ;
        RECT 13.600 74.200 13.900 75.900 ;
        RECT 15.800 75.700 16.200 79.900 ;
        RECT 18.000 78.200 18.400 79.900 ;
        RECT 17.400 77.900 18.400 78.200 ;
        RECT 20.200 77.900 20.600 79.900 ;
        RECT 22.300 77.900 22.900 79.900 ;
        RECT 17.400 77.500 17.800 77.900 ;
        RECT 20.200 77.600 20.500 77.900 ;
        RECT 19.100 77.300 20.900 77.600 ;
        RECT 22.200 77.500 22.600 77.900 ;
        RECT 19.100 77.200 19.500 77.300 ;
        RECT 20.500 77.200 20.900 77.300 ;
        RECT 17.400 76.500 17.800 76.600 ;
        RECT 19.700 76.500 20.100 76.600 ;
        RECT 17.400 76.200 20.100 76.500 ;
        RECT 20.400 76.500 21.500 76.800 ;
        RECT 20.400 75.900 20.700 76.500 ;
        RECT 21.100 76.400 21.500 76.500 ;
        RECT 22.300 76.600 23.000 77.000 ;
        RECT 22.300 76.100 22.600 76.600 ;
        RECT 18.300 75.700 20.700 75.900 ;
        RECT 15.800 75.600 20.700 75.700 ;
        RECT 21.400 75.800 22.600 76.100 ;
        RECT 15.800 75.500 18.700 75.600 ;
        RECT 15.800 75.400 18.600 75.500 ;
        RECT 14.200 74.400 14.600 75.200 ;
        RECT 19.000 75.100 19.400 75.200 ;
        RECT 16.900 74.800 19.400 75.100 ;
        RECT 16.900 74.700 17.300 74.800 ;
        RECT 17.700 74.200 18.100 74.300 ;
        RECT 21.400 74.200 21.700 75.800 ;
        RECT 24.600 75.600 25.000 79.900 ;
        RECT 25.700 76.300 26.100 79.900 ;
        RECT 25.700 75.900 26.600 76.300 ;
        RECT 27.800 75.900 28.200 79.900 ;
        RECT 28.600 76.200 29.000 79.900 ;
        RECT 30.200 76.200 30.600 79.900 ;
        RECT 28.600 75.900 30.600 76.200 ;
        RECT 22.900 75.300 25.000 75.600 ;
        RECT 22.900 75.200 23.300 75.300 ;
        RECT 23.700 74.900 24.100 75.000 ;
        RECT 22.200 74.600 24.100 74.900 ;
        RECT 22.200 74.500 22.600 74.600 ;
        RECT 11.800 74.100 12.200 74.200 ;
        RECT 12.600 74.100 13.900 74.200 ;
        RECT 15.000 74.100 15.400 74.200 ;
        RECT 11.800 73.800 13.900 74.100 ;
        RECT 14.600 73.800 15.400 74.100 ;
        RECT 16.200 73.900 21.700 74.200 ;
        RECT 16.200 73.800 17.000 73.900 ;
        RECT 12.700 73.100 13.000 73.800 ;
        RECT 14.600 73.600 15.000 73.800 ;
        RECT 13.500 73.100 15.300 73.300 ;
        RECT 11.000 72.800 11.900 73.100 ;
        RECT 11.500 71.100 11.900 72.800 ;
        RECT 12.600 71.100 13.000 73.100 ;
        RECT 13.400 73.000 15.400 73.100 ;
        RECT 13.400 71.100 13.800 73.000 ;
        RECT 15.000 71.100 15.400 73.000 ;
        RECT 15.800 71.100 16.200 73.500 ;
        RECT 18.300 73.200 18.600 73.900 ;
        RECT 21.100 73.800 21.500 73.900 ;
        RECT 24.600 73.600 25.000 75.300 ;
        RECT 25.400 74.800 25.800 75.600 ;
        RECT 23.100 73.300 25.000 73.600 ;
        RECT 23.100 73.200 23.500 73.300 ;
        RECT 17.400 72.100 17.800 72.500 ;
        RECT 18.200 72.400 18.600 73.200 ;
        RECT 19.100 72.700 19.500 72.800 ;
        RECT 19.100 72.400 20.500 72.700 ;
        RECT 20.200 72.100 20.500 72.400 ;
        RECT 22.200 72.100 22.600 72.500 ;
        RECT 17.400 71.800 18.400 72.100 ;
        RECT 18.000 71.100 18.400 71.800 ;
        RECT 20.200 71.100 20.600 72.100 ;
        RECT 22.200 71.800 22.900 72.100 ;
        RECT 22.300 71.100 22.900 71.800 ;
        RECT 24.600 71.100 25.000 73.300 ;
        RECT 26.200 74.200 26.500 75.900 ;
        RECT 27.900 75.200 28.200 75.900 ;
        RECT 31.000 75.700 31.400 79.900 ;
        RECT 33.200 78.200 33.600 79.900 ;
        RECT 32.600 77.900 33.600 78.200 ;
        RECT 35.400 77.900 35.800 79.900 ;
        RECT 37.500 77.900 38.100 79.900 ;
        RECT 32.600 77.500 33.000 77.900 ;
        RECT 35.400 77.600 35.700 77.900 ;
        RECT 34.300 77.300 36.100 77.600 ;
        RECT 37.400 77.500 37.800 77.900 ;
        RECT 34.300 77.200 34.700 77.300 ;
        RECT 35.700 77.200 36.100 77.300 ;
        RECT 32.600 76.500 33.000 76.600 ;
        RECT 34.900 76.500 35.300 76.600 ;
        RECT 32.600 76.200 35.300 76.500 ;
        RECT 35.600 76.500 36.700 76.800 ;
        RECT 35.600 75.900 35.900 76.500 ;
        RECT 36.300 76.400 36.700 76.500 ;
        RECT 37.500 76.600 38.200 77.000 ;
        RECT 37.500 76.100 37.800 76.600 ;
        RECT 33.500 75.700 35.900 75.900 ;
        RECT 31.000 75.600 35.900 75.700 ;
        RECT 36.600 75.800 37.800 76.100 ;
        RECT 31.000 75.500 33.900 75.600 ;
        RECT 31.000 75.400 33.800 75.500 ;
        RECT 29.800 75.200 30.200 75.400 ;
        RECT 27.800 74.900 29.000 75.200 ;
        RECT 29.800 74.900 30.600 75.200 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 27.800 74.800 28.200 74.900 ;
        RECT 26.200 74.100 26.600 74.200 ;
        RECT 26.200 73.800 28.100 74.100 ;
        RECT 26.200 72.100 26.500 73.800 ;
        RECT 27.800 73.200 28.100 73.800 ;
        RECT 28.700 73.200 29.000 74.900 ;
        RECT 30.200 74.800 30.600 74.900 ;
        RECT 32.100 74.800 36.200 75.100 ;
        RECT 32.100 74.700 32.500 74.800 ;
        RECT 29.400 73.800 29.800 74.600 ;
        RECT 32.900 74.200 33.300 74.300 ;
        RECT 36.600 74.200 36.900 75.800 ;
        RECT 39.800 75.600 40.200 79.900 ;
        RECT 38.100 75.300 40.200 75.600 ;
        RECT 40.600 77.500 41.000 79.500 ;
        RECT 40.600 75.800 40.900 77.500 ;
        RECT 42.700 76.400 43.100 79.900 ;
        RECT 42.700 76.100 43.500 76.400 ;
        RECT 40.600 75.500 42.500 75.800 ;
        RECT 38.100 75.200 38.500 75.300 ;
        RECT 38.900 74.900 39.300 75.000 ;
        RECT 37.400 74.600 39.300 74.900 ;
        RECT 37.400 74.500 37.800 74.600 ;
        RECT 31.400 73.900 36.900 74.200 ;
        RECT 31.400 73.800 32.200 73.900 ;
        RECT 27.000 72.400 27.400 73.200 ;
        RECT 27.800 72.800 28.200 73.200 ;
        RECT 27.900 72.400 28.300 72.800 ;
        RECT 26.200 71.100 26.600 72.100 ;
        RECT 28.600 71.100 29.000 73.200 ;
        RECT 31.000 71.100 31.400 73.500 ;
        RECT 33.500 73.200 33.800 73.900 ;
        RECT 36.300 73.800 36.700 73.900 ;
        RECT 39.800 73.600 40.200 75.300 ;
        RECT 40.600 74.400 41.000 75.200 ;
        RECT 41.400 74.400 41.800 75.200 ;
        RECT 42.200 74.500 42.500 75.500 ;
        RECT 42.200 74.100 42.900 74.500 ;
        RECT 43.200 74.200 43.500 76.100 ;
        RECT 43.800 75.100 44.200 75.600 ;
        RECT 45.400 75.100 45.800 79.900 ;
        RECT 43.800 74.800 45.800 75.100 ;
        RECT 43.200 74.100 44.200 74.200 ;
        RECT 44.600 74.100 45.000 74.200 ;
        RECT 42.200 73.900 42.700 74.100 ;
        RECT 38.300 73.300 40.200 73.600 ;
        RECT 38.300 73.200 38.700 73.300 ;
        RECT 32.600 72.100 33.000 72.500 ;
        RECT 33.400 72.400 33.800 73.200 ;
        RECT 34.300 72.700 34.700 72.800 ;
        RECT 34.300 72.400 35.700 72.700 ;
        RECT 35.400 72.100 35.700 72.400 ;
        RECT 37.400 72.100 37.800 72.500 ;
        RECT 32.600 71.800 33.600 72.100 ;
        RECT 33.200 71.100 33.600 71.800 ;
        RECT 35.400 71.100 35.800 72.100 ;
        RECT 37.400 71.800 38.100 72.100 ;
        RECT 37.500 71.100 38.100 71.800 ;
        RECT 39.800 71.100 40.200 73.300 ;
        RECT 40.600 73.600 42.700 73.900 ;
        RECT 43.200 73.800 45.000 74.100 ;
        RECT 40.600 72.500 40.900 73.600 ;
        RECT 43.200 73.500 43.500 73.800 ;
        RECT 43.100 73.300 43.500 73.500 ;
        RECT 42.700 73.000 43.500 73.300 ;
        RECT 40.600 71.500 41.000 72.500 ;
        RECT 42.700 71.500 43.100 73.000 ;
        RECT 45.400 71.100 45.800 74.800 ;
        RECT 47.000 75.600 47.400 79.900 ;
        RECT 49.100 77.900 49.700 79.900 ;
        RECT 51.400 77.900 51.800 79.900 ;
        RECT 53.600 78.200 54.000 79.900 ;
        RECT 53.600 77.900 54.600 78.200 ;
        RECT 49.400 77.500 49.800 77.900 ;
        RECT 51.500 77.600 51.800 77.900 ;
        RECT 51.100 77.300 52.900 77.600 ;
        RECT 54.200 77.500 54.600 77.900 ;
        RECT 51.100 77.200 51.500 77.300 ;
        RECT 52.500 77.200 52.900 77.300 ;
        RECT 49.000 76.600 49.700 77.000 ;
        RECT 49.400 76.100 49.700 76.600 ;
        RECT 50.500 76.500 51.600 76.800 ;
        RECT 50.500 76.400 50.900 76.500 ;
        RECT 49.400 75.800 50.600 76.100 ;
        RECT 47.000 75.300 49.100 75.600 ;
        RECT 47.000 73.600 47.400 75.300 ;
        RECT 48.700 75.200 49.100 75.300 ;
        RECT 47.900 74.900 48.300 75.000 ;
        RECT 47.900 74.600 49.800 74.900 ;
        RECT 49.400 74.500 49.800 74.600 ;
        RECT 50.300 74.200 50.600 75.800 ;
        RECT 51.300 75.900 51.600 76.500 ;
        RECT 51.900 76.500 52.300 76.600 ;
        RECT 54.200 76.500 54.600 76.600 ;
        RECT 51.900 76.200 54.600 76.500 ;
        RECT 51.300 75.700 53.700 75.900 ;
        RECT 55.800 75.700 56.200 79.900 ;
        RECT 51.300 75.600 56.200 75.700 ;
        RECT 53.300 75.500 56.200 75.600 ;
        RECT 53.400 75.400 56.200 75.500 ;
        RECT 58.200 75.600 58.600 79.900 ;
        RECT 60.300 77.900 60.900 79.900 ;
        RECT 62.600 77.900 63.000 79.900 ;
        RECT 64.800 78.200 65.200 79.900 ;
        RECT 64.800 77.900 65.800 78.200 ;
        RECT 60.600 77.500 61.000 77.900 ;
        RECT 62.700 77.600 63.000 77.900 ;
        RECT 62.300 77.300 64.100 77.600 ;
        RECT 65.400 77.500 65.800 77.900 ;
        RECT 62.300 77.200 62.700 77.300 ;
        RECT 63.700 77.200 64.100 77.300 ;
        RECT 60.200 76.600 60.900 77.000 ;
        RECT 60.600 76.100 60.900 76.600 ;
        RECT 61.700 76.500 62.800 76.800 ;
        RECT 61.700 76.400 62.100 76.500 ;
        RECT 60.600 75.800 61.800 76.100 ;
        RECT 58.200 75.300 60.300 75.600 ;
        RECT 52.600 75.100 53.000 75.200 ;
        RECT 52.600 74.800 55.100 75.100 ;
        RECT 54.700 74.700 55.100 74.800 ;
        RECT 53.900 74.200 54.300 74.300 ;
        RECT 50.300 74.100 55.800 74.200 ;
        RECT 57.400 74.100 57.800 74.200 ;
        RECT 50.300 73.900 57.800 74.100 ;
        RECT 50.500 73.800 50.900 73.900 ;
        RECT 52.600 73.800 53.000 73.900 ;
        RECT 47.000 73.300 48.900 73.600 ;
        RECT 46.200 73.100 46.600 73.200 ;
        RECT 47.000 73.100 47.400 73.300 ;
        RECT 48.500 73.200 48.900 73.300 ;
        RECT 46.200 72.800 47.400 73.100 ;
        RECT 53.400 72.800 53.700 73.900 ;
        RECT 55.000 73.800 57.800 73.900 ;
        RECT 58.200 73.600 58.600 75.300 ;
        RECT 59.900 75.200 60.300 75.300 ;
        RECT 59.100 74.900 59.500 75.000 ;
        RECT 59.100 74.600 61.000 74.900 ;
        RECT 60.600 74.500 61.000 74.600 ;
        RECT 61.500 74.200 61.800 75.800 ;
        RECT 62.500 75.900 62.800 76.500 ;
        RECT 63.100 76.500 63.500 76.600 ;
        RECT 65.400 76.500 65.800 76.600 ;
        RECT 63.100 76.200 65.800 76.500 ;
        RECT 62.500 75.700 64.900 75.900 ;
        RECT 67.000 75.700 67.400 79.900 ;
        RECT 62.500 75.600 67.400 75.700 ;
        RECT 64.500 75.500 67.400 75.600 ;
        RECT 64.600 75.400 67.400 75.500 ;
        RECT 63.800 75.100 64.200 75.200 ;
        RECT 68.600 75.100 69.000 79.900 ;
        RECT 70.600 76.800 71.000 77.200 ;
        RECT 69.400 75.800 69.800 76.600 ;
        RECT 70.600 76.200 70.900 76.800 ;
        RECT 71.300 76.200 71.700 79.900 ;
        RECT 70.200 75.900 70.900 76.200 ;
        RECT 71.200 75.900 71.700 76.200 ;
        RECT 73.400 77.500 73.800 79.500 ;
        RECT 70.200 75.800 70.600 75.900 ;
        RECT 70.200 75.100 70.500 75.800 ;
        RECT 63.800 74.800 66.300 75.100 ;
        RECT 65.900 74.700 66.300 74.800 ;
        RECT 68.600 74.800 70.500 75.100 ;
        RECT 65.100 74.200 65.500 74.300 ;
        RECT 61.500 73.900 67.000 74.200 ;
        RECT 61.700 73.800 62.100 73.900 ;
        RECT 46.200 72.400 46.600 72.800 ;
        RECT 47.000 71.100 47.400 72.800 ;
        RECT 52.500 72.700 52.900 72.800 ;
        RECT 49.400 72.100 49.800 72.500 ;
        RECT 51.500 72.400 52.900 72.700 ;
        RECT 53.400 72.400 53.800 72.800 ;
        RECT 51.500 72.100 51.800 72.400 ;
        RECT 54.200 72.100 54.600 72.500 ;
        RECT 49.100 71.800 49.800 72.100 ;
        RECT 49.100 71.100 49.700 71.800 ;
        RECT 51.400 71.100 51.800 72.100 ;
        RECT 53.600 71.800 54.600 72.100 ;
        RECT 53.600 71.100 54.000 71.800 ;
        RECT 55.800 71.100 56.200 73.500 ;
        RECT 58.200 73.300 60.100 73.600 ;
        RECT 58.200 71.100 58.600 73.300 ;
        RECT 59.700 73.200 60.100 73.300 ;
        RECT 64.600 72.800 64.900 73.900 ;
        RECT 66.200 73.800 67.000 73.900 ;
        RECT 63.700 72.700 64.100 72.800 ;
        RECT 60.600 72.100 61.000 72.500 ;
        RECT 62.700 72.400 64.100 72.700 ;
        RECT 64.600 72.400 65.000 72.800 ;
        RECT 62.700 72.100 63.000 72.400 ;
        RECT 65.400 72.100 65.800 72.500 ;
        RECT 60.300 71.800 61.000 72.100 ;
        RECT 60.300 71.100 60.900 71.800 ;
        RECT 62.600 71.100 63.000 72.100 ;
        RECT 64.800 71.800 65.800 72.100 ;
        RECT 64.800 71.100 65.200 71.800 ;
        RECT 67.000 71.100 67.400 73.500 ;
        RECT 67.800 73.400 68.200 74.200 ;
        RECT 68.600 73.100 69.000 74.800 ;
        RECT 71.200 74.200 71.500 75.900 ;
        RECT 73.400 75.800 73.700 77.500 ;
        RECT 75.500 76.400 75.900 79.900 ;
        RECT 75.500 76.100 76.300 76.400 ;
        RECT 73.400 75.500 75.300 75.800 ;
        RECT 71.800 74.400 72.200 75.200 ;
        RECT 73.400 74.400 73.800 75.200 ;
        RECT 74.200 74.400 74.600 75.200 ;
        RECT 75.000 74.500 75.300 75.500 ;
        RECT 70.200 73.800 71.500 74.200 ;
        RECT 72.600 74.100 73.000 74.200 ;
        RECT 72.200 73.800 73.000 74.100 ;
        RECT 75.000 74.100 75.700 74.500 ;
        RECT 76.000 74.200 76.300 76.100 ;
        RECT 76.600 75.100 77.000 75.600 ;
        RECT 78.200 75.100 78.600 79.900 ;
        RECT 76.600 74.800 78.600 75.100 ;
        RECT 76.000 74.100 77.000 74.200 ;
        RECT 77.400 74.100 77.800 74.200 ;
        RECT 75.000 73.900 75.500 74.100 ;
        RECT 70.300 73.200 70.600 73.800 ;
        RECT 72.200 73.600 72.600 73.800 ;
        RECT 73.400 73.600 75.500 73.900 ;
        RECT 76.000 73.800 77.800 74.100 ;
        RECT 68.600 72.800 69.500 73.100 ;
        RECT 69.100 71.100 69.500 72.800 ;
        RECT 70.200 71.100 70.600 73.200 ;
        RECT 71.100 73.100 72.900 73.300 ;
        RECT 71.000 73.000 73.000 73.100 ;
        RECT 71.000 71.100 71.400 73.000 ;
        RECT 72.600 71.100 73.000 73.000 ;
        RECT 73.400 72.500 73.700 73.600 ;
        RECT 76.000 73.500 76.300 73.800 ;
        RECT 75.900 73.300 76.300 73.500 ;
        RECT 75.500 73.000 76.300 73.300 ;
        RECT 73.400 71.500 73.800 72.500 ;
        RECT 75.500 71.500 75.900 73.000 ;
        RECT 78.200 71.100 78.600 74.800 ;
        RECT 79.800 75.600 80.200 79.900 ;
        RECT 81.900 77.900 82.500 79.900 ;
        RECT 84.200 77.900 84.600 79.900 ;
        RECT 86.400 78.200 86.800 79.900 ;
        RECT 86.400 77.900 87.400 78.200 ;
        RECT 82.200 77.500 82.600 77.900 ;
        RECT 84.300 77.600 84.600 77.900 ;
        RECT 83.900 77.300 85.700 77.600 ;
        RECT 87.000 77.500 87.400 77.900 ;
        RECT 83.900 77.200 84.300 77.300 ;
        RECT 85.300 77.200 85.700 77.300 ;
        RECT 81.800 76.600 82.500 77.000 ;
        RECT 82.200 76.100 82.500 76.600 ;
        RECT 83.300 76.500 84.400 76.800 ;
        RECT 83.300 76.400 83.700 76.500 ;
        RECT 82.200 75.800 83.400 76.100 ;
        RECT 79.800 75.300 81.900 75.600 ;
        RECT 79.800 73.600 80.200 75.300 ;
        RECT 81.500 75.200 81.900 75.300 ;
        RECT 80.700 74.900 81.100 75.000 ;
        RECT 80.700 74.600 82.600 74.900 ;
        RECT 82.200 74.500 82.600 74.600 ;
        RECT 83.100 74.200 83.400 75.800 ;
        RECT 84.100 75.900 84.400 76.500 ;
        RECT 84.700 76.500 85.100 76.600 ;
        RECT 87.000 76.500 87.400 76.600 ;
        RECT 84.700 76.200 87.400 76.500 ;
        RECT 84.100 75.700 86.500 75.900 ;
        RECT 88.600 75.700 89.000 79.900 ;
        RECT 89.400 76.800 89.800 77.200 ;
        RECT 89.400 76.100 89.700 76.800 ;
        RECT 90.200 76.100 90.600 79.900 ;
        RECT 89.400 75.800 90.600 76.100 ;
        RECT 91.000 75.800 91.400 76.600 ;
        RECT 91.800 75.900 92.200 79.900 ;
        RECT 93.400 77.900 93.800 79.900 ;
        RECT 84.100 75.600 89.000 75.700 ;
        RECT 86.100 75.500 89.000 75.600 ;
        RECT 86.200 75.400 89.000 75.500 ;
        RECT 85.400 75.100 85.800 75.200 ;
        RECT 85.400 74.800 87.900 75.100 ;
        RECT 87.500 74.700 87.900 74.800 ;
        RECT 86.700 74.200 87.100 74.300 ;
        RECT 83.100 73.900 88.600 74.200 ;
        RECT 83.300 73.800 83.700 73.900 ;
        RECT 79.800 73.300 81.700 73.600 ;
        RECT 79.000 73.100 79.400 73.200 ;
        RECT 79.800 73.100 80.200 73.300 ;
        RECT 81.300 73.200 81.700 73.300 ;
        RECT 79.000 72.800 80.200 73.100 ;
        RECT 86.200 72.800 86.500 73.900 ;
        RECT 87.800 73.800 88.600 73.900 ;
        RECT 79.000 72.400 79.400 72.800 ;
        RECT 79.800 71.100 80.200 72.800 ;
        RECT 85.300 72.700 85.700 72.800 ;
        RECT 82.200 72.100 82.600 72.500 ;
        RECT 84.300 72.400 85.700 72.700 ;
        RECT 86.200 72.400 86.600 72.800 ;
        RECT 84.300 72.100 84.600 72.400 ;
        RECT 87.000 72.100 87.400 72.500 ;
        RECT 81.900 71.800 82.600 72.100 ;
        RECT 81.900 71.100 82.500 71.800 ;
        RECT 84.200 71.100 84.600 72.100 ;
        RECT 86.400 71.800 87.400 72.100 ;
        RECT 86.400 71.100 86.800 71.800 ;
        RECT 88.600 71.100 89.000 73.500 ;
        RECT 89.400 73.400 89.800 74.200 ;
        RECT 90.200 73.100 90.600 75.800 ;
        RECT 91.800 75.200 92.100 75.900 ;
        RECT 93.400 75.800 93.700 77.900 ;
        RECT 95.000 76.100 95.400 76.200 ;
        RECT 95.800 76.100 96.200 79.900 ;
        RECT 95.000 75.800 96.200 76.100 ;
        RECT 96.600 75.800 97.000 76.600 ;
        RECT 98.200 76.400 98.600 79.900 ;
        RECT 98.100 75.900 98.600 76.400 ;
        RECT 99.800 76.200 100.200 79.900 ;
        RECT 98.900 75.900 100.200 76.200 ;
        RECT 100.600 76.200 101.000 79.900 ;
        RECT 102.200 76.400 102.600 79.900 ;
        RECT 100.600 75.900 101.900 76.200 ;
        RECT 102.200 75.900 102.700 76.400 ;
        RECT 105.100 76.200 105.500 79.900 ;
        RECT 105.800 76.800 106.200 77.200 ;
        RECT 105.900 76.200 106.200 76.800 ;
        RECT 105.100 75.900 105.600 76.200 ;
        RECT 105.900 75.900 106.600 76.200 ;
        RECT 92.500 75.500 93.700 75.800 ;
        RECT 91.800 74.800 92.200 75.200 ;
        RECT 91.800 73.100 92.100 74.800 ;
        RECT 92.500 73.800 92.800 75.500 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 93.400 74.400 93.700 74.800 ;
        RECT 93.200 74.100 93.700 74.400 ;
        RECT 93.200 74.000 93.600 74.100 ;
        RECT 94.200 73.800 94.600 75.200 ;
        RECT 92.400 73.700 92.800 73.800 ;
        RECT 92.400 73.500 93.900 73.700 ;
        RECT 92.400 73.400 94.500 73.500 ;
        RECT 95.000 73.400 95.400 74.200 ;
        RECT 93.600 73.200 94.500 73.400 ;
        RECT 94.200 73.100 94.500 73.200 ;
        RECT 95.800 73.100 96.200 75.800 ;
        RECT 98.100 74.200 98.400 75.900 ;
        RECT 98.900 74.900 99.200 75.900 ;
        RECT 98.700 74.500 99.200 74.900 ;
        RECT 98.100 73.800 98.600 74.200 ;
        RECT 98.100 73.100 98.400 73.800 ;
        RECT 98.900 73.700 99.200 74.500 ;
        RECT 99.700 75.100 100.200 75.200 ;
        RECT 100.600 75.100 101.100 75.200 ;
        RECT 99.700 74.800 101.100 75.100 ;
        RECT 99.700 74.400 100.100 74.800 ;
        RECT 100.700 74.400 101.100 74.800 ;
        RECT 101.600 74.900 101.900 75.900 ;
        RECT 101.600 74.500 102.100 74.900 ;
        RECT 101.600 73.700 101.900 74.500 ;
        RECT 102.400 74.200 102.700 75.900 ;
        RECT 104.600 74.400 105.000 75.200 ;
        RECT 105.300 74.200 105.600 75.900 ;
        RECT 106.200 75.800 106.600 75.900 ;
        RECT 108.600 75.800 109.000 76.600 ;
        RECT 106.200 75.100 106.500 75.800 ;
        RECT 109.400 75.100 109.800 79.900 ;
        RECT 111.000 75.700 111.400 79.900 ;
        RECT 113.200 78.200 113.600 79.900 ;
        RECT 112.600 77.900 113.600 78.200 ;
        RECT 115.400 77.900 115.800 79.900 ;
        RECT 117.500 77.900 118.100 79.900 ;
        RECT 112.600 77.500 113.000 77.900 ;
        RECT 115.400 77.600 115.700 77.900 ;
        RECT 114.300 77.300 116.100 77.600 ;
        RECT 117.400 77.500 117.800 77.900 ;
        RECT 114.300 77.200 114.700 77.300 ;
        RECT 115.700 77.200 116.100 77.300 ;
        RECT 112.600 76.500 113.000 76.600 ;
        RECT 114.900 76.500 115.300 76.600 ;
        RECT 112.600 76.200 115.300 76.500 ;
        RECT 115.600 76.500 116.700 76.800 ;
        RECT 115.600 75.900 115.900 76.500 ;
        RECT 116.300 76.400 116.700 76.500 ;
        RECT 117.500 76.600 118.200 77.000 ;
        RECT 117.500 76.100 117.800 76.600 ;
        RECT 113.500 75.700 115.900 75.900 ;
        RECT 111.000 75.600 115.900 75.700 ;
        RECT 116.600 75.800 117.800 76.100 ;
        RECT 111.000 75.500 113.900 75.600 ;
        RECT 111.000 75.400 113.800 75.500 ;
        RECT 116.600 75.200 116.900 75.800 ;
        RECT 119.800 75.600 120.200 79.900 ;
        RECT 121.400 75.600 121.800 79.900 ;
        RECT 123.000 75.600 123.400 79.900 ;
        RECT 124.600 75.600 125.000 79.900 ;
        RECT 126.200 75.600 126.600 79.900 ;
        RECT 127.800 77.100 128.200 77.200 ;
        RECT 128.600 77.100 129.000 79.900 ;
        RECT 127.800 76.800 129.000 77.100 ;
        RECT 118.100 75.300 120.200 75.600 ;
        RECT 118.100 75.200 118.500 75.300 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 106.200 74.800 109.800 75.100 ;
        RECT 102.200 74.100 102.700 74.200 ;
        RECT 103.800 74.100 104.200 74.200 ;
        RECT 102.200 73.800 104.600 74.100 ;
        RECT 105.300 73.800 106.600 74.200 ;
        RECT 98.900 73.400 100.200 73.700 ;
        RECT 90.200 72.800 91.100 73.100 ;
        RECT 90.700 71.100 91.100 72.800 ;
        RECT 91.800 72.600 92.500 73.100 ;
        RECT 92.100 72.200 92.500 72.600 ;
        RECT 91.800 71.800 92.500 72.200 ;
        RECT 92.100 71.100 92.500 71.800 ;
        RECT 94.200 71.100 94.600 73.100 ;
        RECT 95.800 72.800 96.700 73.100 ;
        RECT 98.100 72.800 98.600 73.100 ;
        RECT 96.300 71.100 96.700 72.800 ;
        RECT 98.200 71.100 98.600 72.800 ;
        RECT 99.800 71.100 100.200 73.400 ;
        RECT 100.600 73.400 101.900 73.700 ;
        RECT 100.600 71.100 101.000 73.400 ;
        RECT 102.400 73.100 102.700 73.800 ;
        RECT 104.200 73.600 104.600 73.800 ;
        RECT 103.900 73.100 105.700 73.300 ;
        RECT 106.200 73.100 106.500 73.800 ;
        RECT 109.400 73.100 109.800 74.800 ;
        RECT 112.100 74.800 114.600 75.100 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 118.900 74.900 119.300 75.000 ;
        RECT 112.100 74.700 112.500 74.800 ;
        RECT 113.400 74.700 113.800 74.800 ;
        RECT 112.900 74.200 113.300 74.300 ;
        RECT 116.600 74.200 116.900 74.800 ;
        RECT 117.400 74.600 119.300 74.900 ;
        RECT 117.400 74.500 117.800 74.600 ;
        RECT 110.200 73.400 110.600 74.200 ;
        RECT 111.400 73.900 116.900 74.200 ;
        RECT 111.400 73.800 112.200 73.900 ;
        RECT 102.200 72.800 102.700 73.100 ;
        RECT 103.800 73.000 105.800 73.100 ;
        RECT 102.200 71.100 102.600 72.800 ;
        RECT 103.800 71.100 104.200 73.000 ;
        RECT 105.400 71.100 105.800 73.000 ;
        RECT 106.200 71.100 106.600 73.100 ;
        RECT 108.900 72.800 109.800 73.100 ;
        RECT 108.900 71.100 109.300 72.800 ;
        RECT 111.000 71.100 111.400 73.500 ;
        RECT 113.500 72.800 113.800 73.900 ;
        RECT 116.300 73.800 116.700 73.900 ;
        RECT 119.800 73.600 120.200 75.300 ;
        RECT 118.300 73.300 120.200 73.600 ;
        RECT 120.600 75.200 121.800 75.600 ;
        RECT 122.300 75.200 123.400 75.600 ;
        RECT 123.900 75.200 125.000 75.600 ;
        RECT 125.700 75.200 126.600 75.600 ;
        RECT 120.600 73.800 121.000 75.200 ;
        RECT 122.300 74.500 122.700 75.200 ;
        RECT 123.900 74.500 124.300 75.200 ;
        RECT 125.700 74.500 126.100 75.200 ;
        RECT 127.000 75.100 127.400 75.200 ;
        RECT 127.000 74.800 128.100 75.100 ;
        RECT 121.400 74.100 122.700 74.500 ;
        RECT 123.100 74.100 124.300 74.500 ;
        RECT 124.800 74.100 126.100 74.500 ;
        RECT 126.500 74.100 127.400 74.500 ;
        RECT 122.300 73.800 122.700 74.100 ;
        RECT 123.900 73.800 124.300 74.100 ;
        RECT 125.700 73.800 126.100 74.100 ;
        RECT 127.000 73.800 127.400 74.100 ;
        RECT 127.800 74.200 128.100 74.800 ;
        RECT 120.600 73.400 121.800 73.800 ;
        RECT 122.300 73.400 123.400 73.800 ;
        RECT 123.900 73.400 125.000 73.800 ;
        RECT 125.700 73.400 126.600 73.800 ;
        RECT 127.800 73.400 128.200 74.200 ;
        RECT 118.300 73.200 118.700 73.300 ;
        RECT 112.600 72.100 113.000 72.500 ;
        RECT 113.400 72.400 113.800 72.800 ;
        RECT 114.300 72.700 114.700 72.800 ;
        RECT 114.300 72.400 115.700 72.700 ;
        RECT 115.400 72.100 115.700 72.400 ;
        RECT 117.400 72.100 117.800 72.500 ;
        RECT 112.600 71.800 113.600 72.100 ;
        RECT 113.200 71.100 113.600 71.800 ;
        RECT 115.400 71.100 115.800 72.100 ;
        RECT 117.400 71.800 118.100 72.100 ;
        RECT 117.500 71.100 118.100 71.800 ;
        RECT 119.800 71.100 120.200 73.300 ;
        RECT 121.400 71.100 121.800 73.400 ;
        RECT 123.000 71.100 123.400 73.400 ;
        RECT 124.600 71.100 125.000 73.400 ;
        RECT 126.200 71.100 126.600 73.400 ;
        RECT 128.600 73.100 129.000 76.800 ;
        RECT 129.400 75.800 129.800 76.600 ;
        RECT 130.200 75.700 130.600 79.900 ;
        RECT 132.400 78.200 132.800 79.900 ;
        RECT 131.800 77.900 132.800 78.200 ;
        RECT 134.600 77.900 135.000 79.900 ;
        RECT 136.700 77.900 137.300 79.900 ;
        RECT 131.800 77.500 132.200 77.900 ;
        RECT 134.600 77.600 134.900 77.900 ;
        RECT 133.500 77.300 135.300 77.600 ;
        RECT 136.600 77.500 137.000 77.900 ;
        RECT 133.500 77.200 133.900 77.300 ;
        RECT 134.900 77.200 135.300 77.300 ;
        RECT 131.800 76.500 132.200 76.600 ;
        RECT 134.100 76.500 134.500 76.600 ;
        RECT 131.800 76.200 134.500 76.500 ;
        RECT 134.800 76.500 135.900 76.800 ;
        RECT 134.800 75.900 135.100 76.500 ;
        RECT 135.500 76.400 135.900 76.500 ;
        RECT 136.700 76.600 137.400 77.000 ;
        RECT 136.700 76.100 137.000 76.600 ;
        RECT 132.700 75.700 135.100 75.900 ;
        RECT 130.200 75.600 135.100 75.700 ;
        RECT 135.800 75.800 137.000 76.100 ;
        RECT 130.200 75.500 133.100 75.600 ;
        RECT 130.200 75.400 133.000 75.500 ;
        RECT 133.400 75.100 133.800 75.200 ;
        RECT 131.300 74.800 133.800 75.100 ;
        RECT 131.300 74.700 131.700 74.800 ;
        RECT 132.100 74.200 132.500 74.300 ;
        RECT 135.800 74.200 136.100 75.800 ;
        RECT 139.000 75.600 139.400 79.900 ;
        RECT 141.100 76.300 141.500 79.900 ;
        RECT 140.600 75.900 141.500 76.300 ;
        RECT 142.200 77.500 142.600 79.500 ;
        RECT 144.300 79.200 144.700 79.900 ;
        RECT 144.300 78.800 145.000 79.200 ;
        RECT 137.300 75.300 139.400 75.600 ;
        RECT 137.300 75.200 137.700 75.300 ;
        RECT 138.100 74.900 138.500 75.000 ;
        RECT 136.600 74.600 138.500 74.900 ;
        RECT 136.600 74.500 137.000 74.600 ;
        RECT 130.600 73.900 136.100 74.200 ;
        RECT 130.600 73.800 131.400 73.900 ;
        RECT 128.600 72.800 129.500 73.100 ;
        RECT 129.100 71.100 129.500 72.800 ;
        RECT 130.200 71.100 130.600 73.500 ;
        RECT 132.700 73.200 133.000 73.900 ;
        RECT 135.500 73.800 135.900 73.900 ;
        RECT 139.000 73.600 139.400 75.300 ;
        RECT 140.700 74.200 141.000 75.900 ;
        RECT 142.200 75.800 142.500 77.500 ;
        RECT 144.300 76.400 144.700 78.800 ;
        RECT 144.300 76.100 145.100 76.400 ;
        RECT 141.400 74.800 141.800 75.600 ;
        RECT 142.200 75.500 144.100 75.800 ;
        RECT 142.200 74.400 142.600 75.200 ;
        RECT 143.000 74.400 143.400 75.200 ;
        RECT 143.800 74.500 144.100 75.500 ;
        RECT 140.600 73.800 141.000 74.200 ;
        RECT 143.800 74.100 144.500 74.500 ;
        RECT 144.800 74.200 145.100 76.100 ;
        RECT 147.000 75.700 147.400 79.900 ;
        RECT 149.200 78.200 149.600 79.900 ;
        RECT 148.600 77.900 149.600 78.200 ;
        RECT 151.400 77.900 151.800 79.900 ;
        RECT 153.500 77.900 154.100 79.900 ;
        RECT 148.600 77.500 149.000 77.900 ;
        RECT 151.400 77.600 151.700 77.900 ;
        RECT 150.300 77.300 152.100 77.600 ;
        RECT 153.400 77.500 153.800 77.900 ;
        RECT 150.300 77.200 150.700 77.300 ;
        RECT 151.700 77.200 152.100 77.300 ;
        RECT 148.600 76.500 149.000 76.600 ;
        RECT 150.900 76.500 151.300 76.600 ;
        RECT 148.600 76.200 151.300 76.500 ;
        RECT 151.600 76.500 152.700 76.800 ;
        RECT 151.600 75.900 151.900 76.500 ;
        RECT 152.300 76.400 152.700 76.500 ;
        RECT 153.500 76.600 154.200 77.000 ;
        RECT 153.500 76.100 153.800 76.600 ;
        RECT 149.500 75.700 151.900 75.900 ;
        RECT 147.000 75.600 151.900 75.700 ;
        RECT 152.600 75.800 153.800 76.100 ;
        RECT 145.400 74.800 145.800 75.600 ;
        RECT 147.000 75.500 149.900 75.600 ;
        RECT 147.000 75.400 149.800 75.500 ;
        RECT 150.200 75.100 150.600 75.200 ;
        RECT 151.000 75.100 151.400 75.200 ;
        RECT 148.100 74.800 151.400 75.100 ;
        RECT 148.100 74.700 148.500 74.800 ;
        RECT 148.900 74.200 149.300 74.300 ;
        RECT 152.600 74.200 152.900 75.800 ;
        RECT 155.800 75.600 156.200 79.900 ;
        RECT 154.100 75.300 156.200 75.600 ;
        RECT 154.100 75.200 154.500 75.300 ;
        RECT 154.900 74.900 155.300 75.000 ;
        RECT 153.400 74.600 155.300 74.900 ;
        RECT 153.400 74.500 153.800 74.600 ;
        RECT 143.800 73.900 144.300 74.100 ;
        RECT 137.500 73.300 139.400 73.600 ;
        RECT 137.500 73.200 137.900 73.300 ;
        RECT 131.800 72.100 132.200 72.500 ;
        RECT 132.600 72.400 133.000 73.200 ;
        RECT 139.000 73.100 139.400 73.300 ;
        RECT 139.800 73.100 140.200 73.200 ;
        RECT 139.000 72.800 140.200 73.100 ;
        RECT 133.500 72.700 133.900 72.800 ;
        RECT 133.500 72.400 134.900 72.700 ;
        RECT 134.600 72.100 134.900 72.400 ;
        RECT 136.600 72.100 137.000 72.500 ;
        RECT 131.800 71.800 132.800 72.100 ;
        RECT 132.400 71.100 132.800 71.800 ;
        RECT 134.600 71.100 135.000 72.100 ;
        RECT 136.600 71.800 137.300 72.100 ;
        RECT 136.700 71.100 137.300 71.800 ;
        RECT 139.000 71.100 139.400 72.800 ;
        RECT 139.800 72.400 140.200 72.800 ;
        RECT 140.700 72.200 141.000 73.800 ;
        RECT 140.600 71.100 141.000 72.200 ;
        RECT 142.200 73.600 144.300 73.900 ;
        RECT 144.800 73.800 145.800 74.200 ;
        RECT 147.400 73.900 152.900 74.200 ;
        RECT 147.400 73.800 148.200 73.900 ;
        RECT 142.200 72.500 142.500 73.600 ;
        RECT 144.800 73.500 145.100 73.800 ;
        RECT 144.700 73.300 145.100 73.500 ;
        RECT 144.300 73.000 145.100 73.300 ;
        RECT 142.200 71.500 142.600 72.500 ;
        RECT 144.300 71.500 144.700 73.000 ;
        RECT 147.000 71.100 147.400 73.500 ;
        RECT 149.500 72.800 149.800 73.900 ;
        RECT 152.300 73.800 152.700 73.900 ;
        RECT 155.800 73.600 156.200 75.300 ;
        RECT 154.300 73.300 156.200 73.600 ;
        RECT 158.200 73.400 158.600 74.200 ;
        RECT 154.300 73.200 154.700 73.300 ;
        RECT 148.600 72.100 149.000 72.500 ;
        RECT 149.400 72.400 149.800 72.800 ;
        RECT 150.300 72.700 150.700 72.800 ;
        RECT 150.300 72.400 151.700 72.700 ;
        RECT 151.400 72.100 151.700 72.400 ;
        RECT 153.400 72.100 153.800 72.500 ;
        RECT 148.600 71.800 149.600 72.100 ;
        RECT 149.200 71.100 149.600 71.800 ;
        RECT 151.400 71.100 151.800 72.100 ;
        RECT 153.400 71.800 154.100 72.100 ;
        RECT 153.500 71.100 154.100 71.800 ;
        RECT 155.800 71.100 156.200 73.300 ;
        RECT 159.000 73.100 159.400 79.900 ;
        RECT 161.400 77.900 161.800 79.900 ;
        RECT 159.800 75.800 160.200 76.600 ;
        RECT 161.500 75.800 161.800 77.900 ;
        RECT 163.000 75.900 163.400 79.900 ;
        RECT 164.900 79.200 165.300 79.900 ;
        RECT 164.900 78.800 165.800 79.200 ;
        RECT 164.200 76.800 164.600 77.200 ;
        RECT 164.200 76.200 164.500 76.800 ;
        RECT 164.900 76.200 165.300 78.800 ;
        RECT 168.900 76.400 169.300 79.900 ;
        RECT 171.000 77.500 171.400 79.500 ;
        RECT 161.500 75.500 162.700 75.800 ;
        RECT 161.400 74.800 161.800 75.200 ;
        RECT 159.800 74.100 160.200 74.200 ;
        RECT 160.600 74.100 161.000 74.600 ;
        RECT 161.500 74.400 161.800 74.800 ;
        RECT 159.800 73.800 161.000 74.100 ;
        RECT 161.400 74.000 162.000 74.400 ;
        RECT 162.400 73.800 162.700 75.500 ;
        RECT 163.100 75.200 163.400 75.900 ;
        RECT 163.800 75.900 164.500 76.200 ;
        RECT 164.800 75.900 165.300 76.200 ;
        RECT 168.500 76.100 169.300 76.400 ;
        RECT 163.800 75.800 164.200 75.900 ;
        RECT 163.000 74.800 163.400 75.200 ;
        RECT 162.400 73.700 162.800 73.800 ;
        RECT 161.300 73.500 162.800 73.700 ;
        RECT 160.700 73.400 162.800 73.500 ;
        RECT 160.700 73.200 161.600 73.400 ;
        RECT 160.700 73.100 161.000 73.200 ;
        RECT 163.100 73.100 163.400 74.800 ;
        RECT 164.800 74.200 165.100 75.900 ;
        RECT 165.400 74.400 165.800 75.200 ;
        RECT 167.000 75.100 167.400 75.200 ;
        RECT 167.800 75.100 168.200 75.600 ;
        RECT 167.000 74.800 168.200 75.100 ;
        RECT 168.500 74.200 168.800 76.100 ;
        RECT 171.100 75.800 171.400 77.500 ;
        RECT 169.500 75.500 171.400 75.800 ;
        RECT 171.800 77.500 172.200 79.500 ;
        RECT 171.800 75.800 172.100 77.500 ;
        RECT 173.900 76.400 174.300 79.900 ;
        RECT 173.900 76.100 174.700 76.400 ;
        RECT 171.800 75.500 173.700 75.800 ;
        RECT 169.500 74.500 169.800 75.500 ;
        RECT 163.800 73.800 165.100 74.200 ;
        RECT 166.200 74.100 166.600 74.200 ;
        RECT 165.800 73.800 166.600 74.100 ;
        RECT 167.800 73.800 168.800 74.200 ;
        RECT 169.100 74.100 169.800 74.500 ;
        RECT 170.200 74.400 170.600 75.200 ;
        RECT 171.000 74.400 171.400 75.200 ;
        RECT 171.800 74.400 172.200 75.200 ;
        RECT 172.600 74.400 173.000 75.200 ;
        RECT 173.400 74.500 173.700 75.500 ;
        RECT 163.900 73.100 164.200 73.800 ;
        RECT 165.800 73.600 166.200 73.800 ;
        RECT 168.500 73.500 168.800 73.800 ;
        RECT 169.300 73.900 169.800 74.100 ;
        RECT 173.400 74.100 174.100 74.500 ;
        RECT 174.400 74.200 174.700 76.100 ;
        RECT 176.600 75.600 177.000 79.900 ;
        RECT 178.700 77.900 179.300 79.900 ;
        RECT 181.000 77.900 181.400 79.900 ;
        RECT 183.200 78.200 183.600 79.900 ;
        RECT 183.200 77.900 184.200 78.200 ;
        RECT 179.000 77.500 179.400 77.900 ;
        RECT 181.100 77.600 181.400 77.900 ;
        RECT 180.700 77.300 182.500 77.600 ;
        RECT 183.800 77.500 184.200 77.900 ;
        RECT 180.700 77.200 181.100 77.300 ;
        RECT 182.100 77.200 182.500 77.300 ;
        RECT 178.600 76.600 179.300 77.000 ;
        RECT 179.000 76.100 179.300 76.600 ;
        RECT 180.100 76.500 181.200 76.800 ;
        RECT 180.100 76.400 180.500 76.500 ;
        RECT 179.000 75.800 180.200 76.100 ;
        RECT 175.000 75.100 175.400 75.600 ;
        RECT 176.600 75.300 178.700 75.600 ;
        RECT 176.600 75.100 177.000 75.300 ;
        RECT 178.300 75.200 178.700 75.300 ;
        RECT 175.000 74.800 177.000 75.100 ;
        RECT 173.400 73.900 173.900 74.100 ;
        RECT 169.300 73.600 171.400 73.900 ;
        RECT 168.500 73.300 168.900 73.500 ;
        RECT 164.700 73.100 166.500 73.300 ;
        RECT 159.000 72.800 159.900 73.100 ;
        RECT 159.500 71.100 159.900 72.800 ;
        RECT 160.600 71.100 161.000 73.100 ;
        RECT 162.700 72.600 163.400 73.100 ;
        RECT 162.700 71.100 163.100 72.600 ;
        RECT 163.800 71.100 164.200 73.100 ;
        RECT 164.600 73.000 166.600 73.100 ;
        RECT 168.500 73.000 169.300 73.300 ;
        RECT 164.600 71.100 165.000 73.000 ;
        RECT 166.200 71.100 166.600 73.000 ;
        RECT 168.900 71.500 169.300 73.000 ;
        RECT 171.100 72.500 171.400 73.600 ;
        RECT 171.000 71.500 171.400 72.500 ;
        RECT 171.800 73.600 173.900 73.900 ;
        RECT 174.400 73.800 175.400 74.200 ;
        RECT 171.800 72.500 172.100 73.600 ;
        RECT 174.400 73.500 174.700 73.800 ;
        RECT 174.300 73.300 174.700 73.500 ;
        RECT 173.900 73.000 174.700 73.300 ;
        RECT 176.600 73.600 177.000 74.800 ;
        RECT 177.500 74.900 177.900 75.000 ;
        RECT 177.500 74.600 179.400 74.900 ;
        RECT 179.000 74.500 179.400 74.600 ;
        RECT 179.900 74.200 180.200 75.800 ;
        RECT 180.900 75.900 181.200 76.500 ;
        RECT 181.500 76.500 181.900 76.600 ;
        RECT 183.800 76.500 184.200 76.600 ;
        RECT 181.500 76.200 184.200 76.500 ;
        RECT 180.900 75.700 183.300 75.900 ;
        RECT 185.400 75.700 185.800 79.900 ;
        RECT 187.500 76.300 187.900 79.900 ;
        RECT 187.000 75.900 187.900 76.300 ;
        RECT 188.600 75.900 189.000 79.900 ;
        RECT 189.400 76.200 189.800 79.900 ;
        RECT 191.000 76.200 191.400 79.900 ;
        RECT 193.700 76.400 194.100 79.900 ;
        RECT 195.800 77.500 196.200 79.500 ;
        RECT 189.400 75.900 191.400 76.200 ;
        RECT 193.300 76.100 194.100 76.400 ;
        RECT 180.900 75.600 185.800 75.700 ;
        RECT 182.900 75.500 185.800 75.600 ;
        RECT 183.000 75.400 185.800 75.500 ;
        RECT 182.200 75.100 182.600 75.200 ;
        RECT 182.200 74.800 184.700 75.100 ;
        RECT 183.000 74.700 183.400 74.800 ;
        RECT 184.300 74.700 184.700 74.800 ;
        RECT 183.500 74.200 183.900 74.300 ;
        RECT 187.100 74.200 187.400 75.900 ;
        RECT 187.800 74.800 188.200 75.600 ;
        RECT 188.700 75.200 189.000 75.900 ;
        RECT 190.600 75.200 191.000 75.400 ;
        RECT 188.600 74.900 189.800 75.200 ;
        RECT 190.600 74.900 191.400 75.200 ;
        RECT 188.600 74.800 189.000 74.900 ;
        RECT 189.500 74.200 189.800 74.900 ;
        RECT 191.000 74.800 191.400 74.900 ;
        RECT 191.800 75.100 192.200 75.200 ;
        RECT 192.600 75.100 193.000 75.600 ;
        RECT 191.800 74.800 193.000 75.100 ;
        RECT 178.200 73.600 178.600 74.200 ;
        RECT 179.900 73.900 185.400 74.200 ;
        RECT 180.100 73.800 180.500 73.900 ;
        RECT 176.600 73.300 178.600 73.600 ;
        RECT 171.800 71.500 172.200 72.500 ;
        RECT 173.900 72.200 174.300 73.000 ;
        RECT 173.400 71.800 174.300 72.200 ;
        RECT 173.900 71.500 174.300 71.800 ;
        RECT 176.600 71.100 177.000 73.300 ;
        RECT 178.100 73.200 178.500 73.300 ;
        RECT 183.000 72.800 183.300 73.900 ;
        RECT 184.600 73.800 185.400 73.900 ;
        RECT 187.000 73.800 187.400 74.200 ;
        RECT 189.400 73.800 189.800 74.200 ;
        RECT 190.200 73.800 190.600 74.600 ;
        RECT 193.300 74.200 193.600 76.100 ;
        RECT 195.900 75.800 196.200 77.500 ;
        RECT 197.700 79.200 198.100 79.900 ;
        RECT 197.700 78.800 198.600 79.200 ;
        RECT 197.000 76.800 197.400 77.200 ;
        RECT 197.000 76.200 197.300 76.800 ;
        RECT 197.700 76.200 198.100 78.800 ;
        RECT 196.600 75.900 197.300 76.200 ;
        RECT 197.600 75.900 198.100 76.200 ;
        RECT 196.600 75.800 197.000 75.900 ;
        RECT 194.300 75.500 196.200 75.800 ;
        RECT 194.300 74.500 194.600 75.500 ;
        RECT 192.600 73.800 193.600 74.200 ;
        RECT 193.900 74.100 194.600 74.500 ;
        RECT 195.000 74.400 195.400 75.200 ;
        RECT 195.800 74.400 196.200 75.200 ;
        RECT 197.600 74.200 197.900 75.900 ;
        RECT 200.600 75.600 201.000 79.900 ;
        RECT 202.200 75.600 202.600 79.900 ;
        RECT 203.800 75.600 204.200 79.900 ;
        RECT 205.400 75.600 205.800 79.900 ;
        RECT 209.700 78.200 210.100 79.900 ;
        RECT 209.700 77.800 210.600 78.200 ;
        RECT 209.000 76.800 209.400 77.200 ;
        RECT 209.000 76.200 209.300 76.800 ;
        RECT 209.700 76.200 210.100 77.800 ;
        RECT 208.600 75.900 209.300 76.200 ;
        RECT 209.600 75.900 210.100 76.200 ;
        RECT 208.600 75.800 209.000 75.900 ;
        RECT 199.800 75.200 201.000 75.600 ;
        RECT 201.500 75.200 202.600 75.600 ;
        RECT 203.100 75.200 204.200 75.600 ;
        RECT 204.900 75.200 205.800 75.600 ;
        RECT 198.200 74.400 198.600 75.200 ;
        RECT 182.100 72.700 182.500 72.800 ;
        RECT 179.000 72.100 179.400 72.500 ;
        RECT 181.100 72.400 182.500 72.700 ;
        RECT 183.000 72.400 183.400 72.800 ;
        RECT 181.100 72.100 181.400 72.400 ;
        RECT 183.800 72.100 184.200 72.500 ;
        RECT 178.700 71.800 179.400 72.100 ;
        RECT 178.700 71.100 179.300 71.800 ;
        RECT 181.000 71.100 181.400 72.100 ;
        RECT 183.200 71.800 184.200 72.100 ;
        RECT 183.200 71.100 183.600 71.800 ;
        RECT 185.400 71.100 185.800 73.500 ;
        RECT 186.200 72.400 186.600 73.200 ;
        RECT 187.100 73.100 187.400 73.800 ;
        RECT 188.600 73.100 189.000 73.200 ;
        RECT 189.500 73.100 189.800 73.800 ;
        RECT 187.000 72.800 189.000 73.100 ;
        RECT 187.100 72.100 187.400 72.800 ;
        RECT 188.700 72.400 189.100 72.800 ;
        RECT 187.000 71.100 187.400 72.100 ;
        RECT 189.400 71.100 189.800 73.100 ;
        RECT 193.300 73.500 193.600 73.800 ;
        RECT 194.100 73.900 194.600 74.100 ;
        RECT 194.100 73.600 196.200 73.900 ;
        RECT 196.600 73.800 197.900 74.200 ;
        RECT 199.000 74.100 199.400 74.200 ;
        RECT 198.600 73.800 199.400 74.100 ;
        RECT 199.800 73.800 200.200 75.200 ;
        RECT 201.500 74.500 201.900 75.200 ;
        RECT 203.100 74.500 203.500 75.200 ;
        RECT 204.900 74.500 205.300 75.200 ;
        RECT 200.600 74.100 201.900 74.500 ;
        RECT 202.300 74.100 203.500 74.500 ;
        RECT 204.000 74.100 205.300 74.500 ;
        RECT 209.600 74.200 209.900 75.900 ;
        RECT 211.800 75.700 212.200 79.900 ;
        RECT 214.000 78.200 214.400 79.900 ;
        RECT 213.400 77.900 214.400 78.200 ;
        RECT 216.200 77.900 216.600 79.900 ;
        RECT 218.300 77.900 218.900 79.900 ;
        RECT 213.400 77.500 213.800 77.900 ;
        RECT 216.200 77.600 216.500 77.900 ;
        RECT 215.100 77.300 216.900 77.600 ;
        RECT 218.200 77.500 218.600 77.900 ;
        RECT 215.100 77.200 215.500 77.300 ;
        RECT 216.500 77.200 216.900 77.300 ;
        RECT 213.400 76.500 213.800 76.600 ;
        RECT 215.700 76.500 216.100 76.600 ;
        RECT 213.400 76.200 216.100 76.500 ;
        RECT 216.400 76.500 217.500 76.800 ;
        RECT 216.400 75.900 216.700 76.500 ;
        RECT 217.100 76.400 217.500 76.500 ;
        RECT 218.300 76.600 219.000 77.000 ;
        RECT 218.300 76.100 218.600 76.600 ;
        RECT 214.300 75.700 216.700 75.900 ;
        RECT 211.800 75.600 216.700 75.700 ;
        RECT 217.400 75.800 218.600 76.100 ;
        RECT 211.800 75.500 214.700 75.600 ;
        RECT 211.800 75.400 214.600 75.500 ;
        RECT 210.200 74.400 210.600 75.200 ;
        RECT 215.000 75.100 215.400 75.200 ;
        RECT 215.800 75.100 216.200 75.200 ;
        RECT 212.900 74.800 216.200 75.100 ;
        RECT 212.900 74.700 213.300 74.800 ;
        RECT 213.700 74.200 214.100 74.300 ;
        RECT 217.400 74.200 217.700 75.800 ;
        RECT 220.600 75.600 221.000 79.900 ;
        RECT 221.800 76.800 222.200 77.200 ;
        RECT 221.800 76.200 222.100 76.800 ;
        RECT 222.500 76.200 222.900 79.900 ;
        RECT 221.400 75.900 222.100 76.200 ;
        RECT 222.400 75.900 222.900 76.200 ;
        RECT 221.400 75.800 221.800 75.900 ;
        RECT 218.900 75.300 221.000 75.600 ;
        RECT 218.900 75.200 219.300 75.300 ;
        RECT 219.700 74.900 220.100 75.000 ;
        RECT 218.200 74.600 220.100 74.900 ;
        RECT 218.200 74.500 218.600 74.600 ;
        RECT 201.500 73.800 201.900 74.100 ;
        RECT 203.100 73.800 203.500 74.100 ;
        RECT 204.900 73.800 205.300 74.100 ;
        RECT 208.600 73.800 209.900 74.200 ;
        RECT 211.000 74.100 211.400 74.200 ;
        RECT 210.600 73.800 211.400 74.100 ;
        RECT 212.200 73.900 217.700 74.200 ;
        RECT 212.200 73.800 213.000 73.900 ;
        RECT 193.300 73.300 193.700 73.500 ;
        RECT 193.300 73.000 194.100 73.300 ;
        RECT 193.700 71.500 194.100 73.000 ;
        RECT 195.900 72.500 196.200 73.600 ;
        RECT 196.700 73.100 197.000 73.800 ;
        RECT 198.600 73.600 199.000 73.800 ;
        RECT 199.800 73.400 201.000 73.800 ;
        RECT 201.500 73.400 202.600 73.800 ;
        RECT 203.100 73.400 204.200 73.800 ;
        RECT 204.900 73.400 205.800 73.800 ;
        RECT 197.500 73.100 199.300 73.300 ;
        RECT 195.800 71.500 196.200 72.500 ;
        RECT 196.600 71.100 197.000 73.100 ;
        RECT 197.400 73.000 199.400 73.100 ;
        RECT 197.400 71.100 197.800 73.000 ;
        RECT 199.000 71.100 199.400 73.000 ;
        RECT 200.600 71.100 201.000 73.400 ;
        RECT 202.200 71.100 202.600 73.400 ;
        RECT 203.800 71.100 204.200 73.400 ;
        RECT 205.400 71.100 205.800 73.400 ;
        RECT 208.700 73.100 209.000 73.800 ;
        RECT 210.600 73.600 211.000 73.800 ;
        RECT 209.500 73.100 211.300 73.300 ;
        RECT 208.600 71.100 209.000 73.100 ;
        RECT 209.400 73.000 211.400 73.100 ;
        RECT 209.400 71.100 209.800 73.000 ;
        RECT 211.000 71.100 211.400 73.000 ;
        RECT 211.800 71.100 212.200 73.500 ;
        RECT 214.300 72.800 214.600 73.900 ;
        RECT 217.100 73.800 217.500 73.900 ;
        RECT 220.600 73.600 221.000 75.300 ;
        RECT 221.400 75.100 221.800 75.200 ;
        RECT 222.400 75.100 222.700 75.900 ;
        RECT 221.400 74.800 222.700 75.100 ;
        RECT 222.400 74.200 222.700 74.800 ;
        RECT 223.000 74.400 223.400 75.200 ;
        RECT 225.400 75.100 225.800 79.900 ;
        RECT 226.200 75.800 226.600 76.600 ;
        RECT 228.300 76.200 228.700 79.900 ;
        RECT 231.300 77.200 231.700 79.900 ;
        RECT 229.000 76.800 229.400 77.200 ;
        RECT 229.100 76.200 229.400 76.800 ;
        RECT 230.600 76.800 231.000 77.200 ;
        RECT 231.300 76.800 232.200 77.200 ;
        RECT 230.600 76.200 230.900 76.800 ;
        RECT 231.300 76.200 231.700 76.800 ;
        RECT 228.300 75.900 228.800 76.200 ;
        RECT 229.100 75.900 229.800 76.200 ;
        RECT 227.000 75.100 227.400 75.200 ;
        RECT 225.400 74.800 227.400 75.100 ;
        RECT 221.400 73.800 222.700 74.200 ;
        RECT 223.800 74.100 224.200 74.200 ;
        RECT 223.400 73.800 224.200 74.100 ;
        RECT 219.100 73.300 221.000 73.600 ;
        RECT 219.100 73.200 219.500 73.300 ;
        RECT 213.400 72.100 213.800 72.500 ;
        RECT 214.200 72.400 214.600 72.800 ;
        RECT 215.100 72.700 215.500 72.800 ;
        RECT 215.100 72.400 216.500 72.700 ;
        RECT 216.200 72.100 216.500 72.400 ;
        RECT 218.200 72.100 218.600 72.500 ;
        RECT 213.400 71.800 214.400 72.100 ;
        RECT 214.000 71.100 214.400 71.800 ;
        RECT 216.200 71.100 216.600 72.100 ;
        RECT 218.200 71.800 218.900 72.100 ;
        RECT 218.300 71.100 218.900 71.800 ;
        RECT 220.600 71.100 221.000 73.300 ;
        RECT 221.500 73.100 221.800 73.800 ;
        RECT 223.400 73.600 223.800 73.800 ;
        RECT 224.600 73.400 225.000 74.200 ;
        RECT 222.300 73.100 224.100 73.300 ;
        RECT 225.400 73.100 225.800 74.800 ;
        RECT 227.800 74.400 228.200 75.200 ;
        RECT 228.500 74.200 228.800 75.900 ;
        RECT 229.400 75.800 229.800 75.900 ;
        RECT 230.200 75.900 230.900 76.200 ;
        RECT 231.200 75.900 231.700 76.200 ;
        RECT 230.200 75.800 230.600 75.900 ;
        RECT 231.200 74.200 231.500 75.900 ;
        RECT 233.400 75.600 233.800 79.900 ;
        RECT 235.500 77.900 236.100 79.900 ;
        RECT 237.800 77.900 238.200 79.900 ;
        RECT 240.000 78.200 240.400 79.900 ;
        RECT 240.000 77.900 241.000 78.200 ;
        RECT 235.800 77.500 236.200 77.900 ;
        RECT 237.900 77.600 238.200 77.900 ;
        RECT 237.500 77.300 239.300 77.600 ;
        RECT 240.600 77.500 241.000 77.900 ;
        RECT 237.500 77.200 237.900 77.300 ;
        RECT 238.900 77.200 239.300 77.300 ;
        RECT 235.400 76.600 236.100 77.000 ;
        RECT 235.800 76.100 236.100 76.600 ;
        RECT 236.900 76.500 238.000 76.800 ;
        RECT 236.900 76.400 237.300 76.500 ;
        RECT 235.800 75.800 237.000 76.100 ;
        RECT 233.400 75.300 235.500 75.600 ;
        RECT 231.800 74.400 232.200 75.200 ;
        RECT 226.200 74.100 226.600 74.200 ;
        RECT 227.000 74.100 227.400 74.200 ;
        RECT 226.200 73.800 227.800 74.100 ;
        RECT 228.500 73.800 229.800 74.200 ;
        RECT 230.200 73.800 231.500 74.200 ;
        RECT 232.600 74.100 233.000 74.200 ;
        RECT 232.200 73.800 233.000 74.100 ;
        RECT 227.400 73.600 227.800 73.800 ;
        RECT 227.100 73.100 228.900 73.300 ;
        RECT 229.400 73.100 229.700 73.800 ;
        RECT 230.300 73.100 230.600 73.800 ;
        RECT 232.200 73.600 232.600 73.800 ;
        RECT 233.400 73.600 233.800 75.300 ;
        RECT 235.100 75.200 235.500 75.300 ;
        RECT 234.300 74.900 234.700 75.000 ;
        RECT 234.300 74.600 236.200 74.900 ;
        RECT 235.800 74.500 236.200 74.600 ;
        RECT 236.700 74.200 237.000 75.800 ;
        RECT 237.700 75.900 238.000 76.500 ;
        RECT 238.300 76.500 238.700 76.600 ;
        RECT 240.600 76.500 241.000 76.600 ;
        RECT 238.300 76.200 241.000 76.500 ;
        RECT 237.700 75.700 240.100 75.900 ;
        RECT 242.200 75.700 242.600 79.900 ;
        RECT 243.000 76.200 243.400 79.900 ;
        RECT 244.600 76.200 245.000 79.900 ;
        RECT 243.000 75.900 245.000 76.200 ;
        RECT 245.400 75.900 245.800 79.900 ;
        RECT 237.700 75.600 242.600 75.700 ;
        RECT 239.700 75.500 242.600 75.600 ;
        RECT 239.800 75.400 242.600 75.500 ;
        RECT 243.400 75.200 243.800 75.400 ;
        RECT 245.400 75.200 245.700 75.900 ;
        RECT 246.200 75.600 246.600 79.900 ;
        RECT 248.300 77.900 248.900 79.900 ;
        RECT 250.600 77.900 251.000 79.900 ;
        RECT 252.800 78.200 253.200 79.900 ;
        RECT 252.800 77.900 253.800 78.200 ;
        RECT 248.600 77.500 249.000 77.900 ;
        RECT 250.700 77.600 251.000 77.900 ;
        RECT 250.300 77.300 252.100 77.600 ;
        RECT 253.400 77.500 253.800 77.900 ;
        RECT 250.300 77.200 250.700 77.300 ;
        RECT 251.700 77.200 252.100 77.300 ;
        RECT 248.200 76.600 248.900 77.000 ;
        RECT 248.600 76.100 248.900 76.600 ;
        RECT 249.700 76.500 250.800 76.800 ;
        RECT 249.700 76.400 250.100 76.500 ;
        RECT 248.600 75.800 249.800 76.100 ;
        RECT 246.200 75.300 248.300 75.600 ;
        RECT 238.200 75.100 238.600 75.200 ;
        RECT 239.000 75.100 239.400 75.200 ;
        RECT 238.200 74.800 241.500 75.100 ;
        RECT 243.000 74.900 243.800 75.200 ;
        RECT 244.600 74.900 245.800 75.200 ;
        RECT 243.000 74.800 243.400 74.900 ;
        RECT 241.100 74.700 241.500 74.800 ;
        RECT 240.300 74.200 240.700 74.300 ;
        RECT 236.700 73.900 242.200 74.200 ;
        RECT 236.900 73.800 237.300 73.900 ;
        RECT 233.400 73.300 235.300 73.600 ;
        RECT 231.100 73.100 232.900 73.300 ;
        RECT 221.400 71.100 221.800 73.100 ;
        RECT 222.200 73.000 224.200 73.100 ;
        RECT 222.200 71.100 222.600 73.000 ;
        RECT 223.800 71.100 224.200 73.000 ;
        RECT 225.400 72.800 226.300 73.100 ;
        RECT 225.900 71.100 226.300 72.800 ;
        RECT 227.000 73.000 229.000 73.100 ;
        RECT 227.000 71.100 227.400 73.000 ;
        RECT 228.600 71.100 229.000 73.000 ;
        RECT 229.400 71.100 229.800 73.100 ;
        RECT 230.200 71.100 230.600 73.100 ;
        RECT 231.000 73.000 233.000 73.100 ;
        RECT 231.000 71.100 231.400 73.000 ;
        RECT 232.600 71.100 233.000 73.000 ;
        RECT 233.400 71.100 233.800 73.300 ;
        RECT 234.900 73.200 235.300 73.300 ;
        RECT 239.800 72.800 240.100 73.900 ;
        RECT 241.400 73.800 242.200 73.900 ;
        RECT 243.800 73.800 244.200 74.600 ;
        RECT 238.900 72.700 239.300 72.800 ;
        RECT 235.800 72.100 236.200 72.500 ;
        RECT 237.900 72.400 239.300 72.700 ;
        RECT 239.800 72.400 240.200 72.800 ;
        RECT 237.900 72.100 238.200 72.400 ;
        RECT 240.600 72.100 241.000 72.500 ;
        RECT 235.500 71.800 236.200 72.100 ;
        RECT 235.500 71.100 236.100 71.800 ;
        RECT 237.800 71.100 238.200 72.100 ;
        RECT 240.000 71.800 241.000 72.100 ;
        RECT 240.000 71.100 240.400 71.800 ;
        RECT 242.200 71.100 242.600 73.500 ;
        RECT 244.600 73.100 244.900 74.900 ;
        RECT 245.400 74.800 245.800 74.900 ;
        RECT 245.400 74.200 245.700 74.800 ;
        RECT 245.400 73.800 245.800 74.200 ;
        RECT 246.200 73.600 246.600 75.300 ;
        RECT 247.900 75.200 248.300 75.300 ;
        RECT 247.100 74.900 247.500 75.000 ;
        RECT 247.100 74.600 249.000 74.900 ;
        RECT 248.600 74.500 249.000 74.600 ;
        RECT 249.500 74.200 249.800 75.800 ;
        RECT 250.500 75.900 250.800 76.500 ;
        RECT 251.100 76.500 251.500 76.600 ;
        RECT 253.400 76.500 253.800 76.600 ;
        RECT 251.100 76.200 253.800 76.500 ;
        RECT 250.500 75.700 252.900 75.900 ;
        RECT 255.000 75.700 255.400 79.900 ;
        RECT 250.500 75.600 255.400 75.700 ;
        RECT 252.500 75.500 255.400 75.600 ;
        RECT 252.600 75.400 255.400 75.500 ;
        RECT 255.800 75.600 256.200 79.900 ;
        RECT 257.900 77.900 258.500 79.900 ;
        RECT 260.200 77.900 260.600 79.900 ;
        RECT 262.400 78.200 262.800 79.900 ;
        RECT 262.400 77.900 263.400 78.200 ;
        RECT 258.200 77.500 258.600 77.900 ;
        RECT 260.300 77.600 260.600 77.900 ;
        RECT 259.900 77.300 261.700 77.600 ;
        RECT 263.000 77.500 263.400 77.900 ;
        RECT 259.900 77.200 260.300 77.300 ;
        RECT 261.300 77.200 261.700 77.300 ;
        RECT 257.800 76.600 258.500 77.000 ;
        RECT 258.200 76.100 258.500 76.600 ;
        RECT 259.300 76.500 260.400 76.800 ;
        RECT 259.300 76.400 259.700 76.500 ;
        RECT 258.200 75.800 259.400 76.100 ;
        RECT 255.800 75.300 257.900 75.600 ;
        RECT 250.200 75.100 250.600 75.200 ;
        RECT 251.800 75.100 252.200 75.200 ;
        RECT 250.200 74.800 254.300 75.100 ;
        RECT 253.900 74.700 254.300 74.800 ;
        RECT 253.100 74.200 253.500 74.300 ;
        RECT 249.500 73.900 255.000 74.200 ;
        RECT 249.700 73.800 250.100 73.900 ;
        RECT 252.600 73.800 253.000 73.900 ;
        RECT 254.200 73.800 255.000 73.900 ;
        RECT 246.200 73.300 248.100 73.600 ;
        RECT 244.600 71.100 245.000 73.100 ;
        RECT 245.400 72.800 245.800 73.200 ;
        RECT 245.300 72.400 245.700 72.800 ;
        RECT 246.200 71.100 246.600 73.300 ;
        RECT 247.700 73.200 248.100 73.300 ;
        RECT 252.600 72.800 252.900 73.800 ;
        RECT 255.800 73.600 256.200 75.300 ;
        RECT 257.500 75.200 257.900 75.300 ;
        RECT 256.700 74.900 257.100 75.000 ;
        RECT 256.700 74.600 258.600 74.900 ;
        RECT 258.200 74.500 258.600 74.600 ;
        RECT 259.100 74.200 259.400 75.800 ;
        RECT 260.100 75.900 260.400 76.500 ;
        RECT 260.700 76.500 261.100 76.600 ;
        RECT 263.000 76.500 263.400 76.600 ;
        RECT 260.700 76.200 263.400 76.500 ;
        RECT 260.100 75.700 262.500 75.900 ;
        RECT 264.600 75.700 265.000 79.900 ;
        RECT 260.100 75.600 265.000 75.700 ;
        RECT 262.100 75.500 265.000 75.600 ;
        RECT 262.200 75.400 265.000 75.500 ;
        RECT 261.400 75.100 261.800 75.200 ;
        RECT 261.400 74.800 263.900 75.100 ;
        RECT 263.500 74.700 263.900 74.800 ;
        RECT 262.700 74.200 263.100 74.300 ;
        RECT 259.100 73.900 264.600 74.200 ;
        RECT 259.300 73.800 259.700 73.900 ;
        RECT 251.700 72.700 252.100 72.800 ;
        RECT 248.600 72.100 249.000 72.500 ;
        RECT 250.700 72.400 252.100 72.700 ;
        RECT 252.600 72.400 253.000 72.800 ;
        RECT 250.700 72.100 251.000 72.400 ;
        RECT 253.400 72.100 253.800 72.500 ;
        RECT 248.300 71.800 249.000 72.100 ;
        RECT 248.300 71.100 248.900 71.800 ;
        RECT 250.600 71.100 251.000 72.100 ;
        RECT 252.800 71.800 253.800 72.100 ;
        RECT 252.800 71.100 253.200 71.800 ;
        RECT 255.000 71.100 255.400 73.500 ;
        RECT 255.800 73.300 257.700 73.600 ;
        RECT 255.800 71.100 256.200 73.300 ;
        RECT 257.300 73.200 257.700 73.300 ;
        RECT 262.200 72.800 262.500 73.900 ;
        RECT 263.800 73.800 264.600 73.900 ;
        RECT 261.300 72.700 261.700 72.800 ;
        RECT 258.200 72.100 258.600 72.500 ;
        RECT 260.300 72.400 261.700 72.700 ;
        RECT 262.200 72.400 262.600 72.800 ;
        RECT 260.300 72.100 260.600 72.400 ;
        RECT 263.000 72.100 263.400 72.500 ;
        RECT 257.900 71.800 258.600 72.100 ;
        RECT 257.900 71.100 258.500 71.800 ;
        RECT 260.200 71.100 260.600 72.100 ;
        RECT 262.400 71.800 263.400 72.100 ;
        RECT 262.400 71.100 262.800 71.800 ;
        RECT 264.600 71.100 265.000 73.500 ;
        RECT 1.400 67.600 1.800 69.900 ;
        RECT 3.000 67.600 3.400 69.900 ;
        RECT 4.600 67.600 5.000 69.900 ;
        RECT 6.200 67.600 6.600 69.900 ;
        RECT 0.600 67.200 1.800 67.600 ;
        RECT 2.300 67.200 3.400 67.600 ;
        RECT 3.900 67.200 5.000 67.600 ;
        RECT 5.700 67.200 6.600 67.600 ;
        RECT 8.600 67.600 9.000 69.900 ;
        RECT 10.200 67.600 10.600 69.900 ;
        RECT 11.800 67.600 12.200 69.900 ;
        RECT 13.400 67.600 13.800 69.900 ;
        RECT 8.600 67.200 9.500 67.600 ;
        RECT 10.200 67.200 11.300 67.600 ;
        RECT 11.800 67.200 12.900 67.600 ;
        RECT 13.400 67.200 14.600 67.600 ;
        RECT 15.000 67.500 15.400 69.900 ;
        RECT 17.200 69.200 17.600 69.900 ;
        RECT 16.600 68.900 17.600 69.200 ;
        RECT 19.400 68.900 19.800 69.900 ;
        RECT 21.500 69.200 22.100 69.900 ;
        RECT 21.400 68.900 22.100 69.200 ;
        RECT 16.600 68.500 17.000 68.900 ;
        RECT 19.400 68.600 19.700 68.900 ;
        RECT 17.400 68.200 17.800 68.600 ;
        RECT 18.300 68.300 19.700 68.600 ;
        RECT 21.400 68.500 21.800 68.900 ;
        RECT 18.300 68.200 18.700 68.300 ;
        RECT 0.600 65.800 1.000 67.200 ;
        RECT 2.300 66.900 2.700 67.200 ;
        RECT 3.900 66.900 4.300 67.200 ;
        RECT 5.700 66.900 6.100 67.200 ;
        RECT 1.400 66.500 2.700 66.900 ;
        RECT 3.100 66.500 4.300 66.900 ;
        RECT 4.800 66.500 6.100 66.900 ;
        RECT 7.800 66.900 8.200 67.200 ;
        RECT 9.100 66.900 9.500 67.200 ;
        RECT 10.900 66.900 11.300 67.200 ;
        RECT 12.500 66.900 12.900 67.200 ;
        RECT 7.800 66.500 8.700 66.900 ;
        RECT 9.100 66.500 10.400 66.900 ;
        RECT 10.900 66.500 12.100 66.900 ;
        RECT 12.500 66.500 13.800 66.900 ;
        RECT 2.300 65.800 2.700 66.500 ;
        RECT 3.900 65.800 4.300 66.500 ;
        RECT 5.700 65.800 6.100 66.500 ;
        RECT 9.100 65.800 9.500 66.500 ;
        RECT 10.900 65.800 11.300 66.500 ;
        RECT 12.500 65.800 12.900 66.500 ;
        RECT 14.200 65.800 14.600 67.200 ;
        RECT 15.400 67.100 16.200 67.200 ;
        RECT 17.500 67.100 17.800 68.200 ;
        RECT 22.300 67.700 22.700 67.800 ;
        RECT 23.800 67.700 24.200 69.900 ;
        RECT 22.300 67.400 24.200 67.700 ;
        RECT 18.200 67.100 18.600 67.200 ;
        RECT 20.300 67.100 20.700 67.200 ;
        RECT 15.400 66.800 20.900 67.100 ;
        RECT 16.900 66.700 17.300 66.800 ;
        RECT 16.100 66.200 16.500 66.300 ;
        RECT 20.600 66.200 20.900 66.800 ;
        RECT 21.400 66.400 21.800 66.500 ;
        RECT 16.100 66.100 18.600 66.200 ;
        RECT 19.800 66.100 20.200 66.200 ;
        RECT 16.100 65.900 20.200 66.100 ;
        RECT 18.200 65.800 20.200 65.900 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 21.400 66.100 23.300 66.400 ;
        RECT 22.900 66.000 23.300 66.100 ;
        RECT 0.600 65.400 1.800 65.800 ;
        RECT 2.300 65.400 3.400 65.800 ;
        RECT 3.900 65.400 5.000 65.800 ;
        RECT 5.700 65.400 6.600 65.800 ;
        RECT 1.400 61.100 1.800 65.400 ;
        RECT 3.000 61.100 3.400 65.400 ;
        RECT 4.600 61.100 5.000 65.400 ;
        RECT 6.200 61.100 6.600 65.400 ;
        RECT 8.600 65.400 9.500 65.800 ;
        RECT 10.200 65.400 11.300 65.800 ;
        RECT 11.800 65.400 12.900 65.800 ;
        RECT 13.400 65.400 14.600 65.800 ;
        RECT 15.000 65.500 17.800 65.600 ;
        RECT 15.000 65.400 17.900 65.500 ;
        RECT 8.600 61.100 9.000 65.400 ;
        RECT 10.200 61.100 10.600 65.400 ;
        RECT 11.800 61.100 12.200 65.400 ;
        RECT 13.400 61.100 13.800 65.400 ;
        RECT 15.000 65.300 19.900 65.400 ;
        RECT 15.000 61.100 15.400 65.300 ;
        RECT 17.500 65.100 19.900 65.300 ;
        RECT 16.600 64.500 19.300 64.800 ;
        RECT 16.600 64.400 17.000 64.500 ;
        RECT 18.900 64.400 19.300 64.500 ;
        RECT 19.600 64.500 19.900 65.100 ;
        RECT 20.600 65.200 20.900 65.800 ;
        RECT 22.100 65.700 22.500 65.800 ;
        RECT 23.800 65.700 24.200 67.400 ;
        RECT 26.200 67.900 26.600 69.900 ;
        RECT 28.600 68.900 29.000 69.900 ;
        RECT 26.900 68.200 27.300 68.600 ;
        RECT 27.000 68.100 27.400 68.200 ;
        RECT 28.600 68.100 28.900 68.900 ;
        RECT 25.400 66.400 25.800 67.200 ;
        RECT 24.600 66.100 25.000 66.200 ;
        RECT 26.200 66.100 26.500 67.900 ;
        RECT 27.000 67.800 28.900 68.100 ;
        RECT 29.400 67.800 29.800 68.600 ;
        RECT 32.100 68.000 32.500 69.500 ;
        RECT 34.200 68.500 34.600 69.500 ;
        RECT 28.600 67.200 28.900 67.800 ;
        RECT 31.700 67.700 32.500 68.000 ;
        RECT 31.700 67.500 32.100 67.700 ;
        RECT 31.700 67.200 32.000 67.500 ;
        RECT 34.300 67.400 34.600 68.500 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 31.000 66.800 32.000 67.200 ;
        RECT 32.500 67.100 34.600 67.400 ;
        RECT 35.000 68.500 35.400 69.500 ;
        RECT 37.100 69.200 37.500 69.500 ;
        RECT 37.100 68.800 37.800 69.200 ;
        RECT 35.000 67.400 35.300 68.500 ;
        RECT 37.100 68.000 37.500 68.800 ;
        RECT 37.100 67.700 37.900 68.000 ;
        RECT 37.500 67.500 37.900 67.700 ;
        RECT 35.000 67.100 37.100 67.400 ;
        RECT 32.500 66.900 33.000 67.100 ;
        RECT 27.000 66.100 27.400 66.200 ;
        RECT 24.600 65.800 25.400 66.100 ;
        RECT 26.200 65.800 27.400 66.100 ;
        RECT 22.100 65.400 24.200 65.700 ;
        RECT 25.000 65.600 25.400 65.800 ;
        RECT 20.600 64.900 21.800 65.200 ;
        RECT 20.300 64.500 20.700 64.600 ;
        RECT 19.600 64.200 20.700 64.500 ;
        RECT 21.500 64.400 21.800 64.900 ;
        RECT 21.500 64.000 22.200 64.400 ;
        RECT 18.300 63.700 18.700 63.800 ;
        RECT 19.700 63.700 20.100 63.800 ;
        RECT 16.600 63.100 17.000 63.500 ;
        RECT 18.300 63.400 20.100 63.700 ;
        RECT 19.400 63.100 19.700 63.400 ;
        RECT 21.400 63.100 21.800 63.500 ;
        RECT 16.600 62.800 17.600 63.100 ;
        RECT 17.200 61.100 17.600 62.800 ;
        RECT 19.400 61.100 19.800 63.100 ;
        RECT 21.500 61.100 22.100 63.100 ;
        RECT 23.800 61.100 24.200 65.400 ;
        RECT 27.000 65.100 27.300 65.800 ;
        RECT 27.800 65.400 28.200 66.200 ;
        RECT 28.600 65.100 28.900 66.800 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 31.000 66.100 31.400 66.200 ;
        RECT 29.400 65.800 31.400 66.100 ;
        RECT 31.000 65.400 31.400 65.800 ;
        RECT 24.600 64.800 26.600 65.100 ;
        RECT 24.600 61.100 25.000 64.800 ;
        RECT 26.200 61.100 26.600 64.800 ;
        RECT 27.000 61.100 27.400 65.100 ;
        RECT 28.100 64.700 29.000 65.100 ;
        RECT 31.700 64.900 32.000 66.800 ;
        RECT 32.300 66.500 33.000 66.900 ;
        RECT 36.600 66.900 37.100 67.100 ;
        RECT 37.600 67.200 37.900 67.500 ;
        RECT 32.700 65.500 33.000 66.500 ;
        RECT 33.400 65.800 33.800 66.600 ;
        RECT 34.200 65.800 34.600 66.600 ;
        RECT 35.000 65.800 35.400 66.600 ;
        RECT 35.800 65.800 36.200 66.600 ;
        RECT 36.600 66.500 37.300 66.900 ;
        RECT 37.600 66.800 38.600 67.200 ;
        RECT 36.600 65.500 36.900 66.500 ;
        RECT 32.700 65.200 34.600 65.500 ;
        RECT 28.100 61.100 28.500 64.700 ;
        RECT 31.700 64.600 32.500 64.900 ;
        RECT 32.100 63.200 32.500 64.600 ;
        RECT 34.300 63.500 34.600 65.200 ;
        RECT 32.100 62.800 33.000 63.200 ;
        RECT 32.100 61.100 32.500 62.800 ;
        RECT 34.200 61.500 34.600 63.500 ;
        RECT 35.000 65.200 36.900 65.500 ;
        RECT 35.000 63.500 35.300 65.200 ;
        RECT 37.600 64.900 37.900 66.800 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 39.800 66.100 40.200 69.900 ;
        RECT 40.600 67.800 41.000 68.600 ;
        RECT 43.300 68.000 43.700 69.500 ;
        RECT 45.400 68.500 45.800 69.500 ;
        RECT 42.900 67.700 43.700 68.000 ;
        RECT 42.900 67.500 43.300 67.700 ;
        RECT 42.900 67.200 43.200 67.500 ;
        RECT 45.500 67.400 45.800 68.500 ;
        RECT 48.100 68.000 48.500 69.500 ;
        RECT 50.200 68.500 50.600 69.500 ;
        RECT 42.200 66.800 43.200 67.200 ;
        RECT 43.700 67.100 45.800 67.400 ;
        RECT 47.700 67.700 48.500 68.000 ;
        RECT 47.700 67.500 48.100 67.700 ;
        RECT 47.700 67.200 48.000 67.500 ;
        RECT 50.300 67.400 50.600 68.500 ;
        RECT 52.500 69.200 53.300 69.900 ;
        RECT 52.500 68.800 53.800 69.200 ;
        RECT 52.500 67.900 53.300 68.800 ;
        RECT 56.600 68.500 57.000 69.500 ;
        RECT 58.700 69.200 59.100 69.500 ;
        RECT 58.200 68.800 59.100 69.200 ;
        RECT 43.700 66.900 44.200 67.100 ;
        RECT 38.200 65.800 40.200 66.100 ;
        RECT 38.200 65.400 38.600 65.800 ;
        RECT 37.100 64.600 37.900 64.900 ;
        RECT 35.000 61.500 35.400 63.500 ;
        RECT 37.100 61.100 37.500 64.600 ;
        RECT 39.800 61.100 40.200 65.800 ;
        RECT 42.200 65.400 42.600 66.200 ;
        RECT 42.900 64.900 43.200 66.800 ;
        RECT 43.500 66.500 44.200 66.900 ;
        RECT 47.000 66.800 48.000 67.200 ;
        RECT 48.500 67.100 50.600 67.400 ;
        RECT 48.500 66.900 49.000 67.100 ;
        RECT 43.900 65.500 44.200 66.500 ;
        RECT 44.600 65.800 45.000 66.600 ;
        RECT 45.400 65.800 45.800 66.600 ;
        RECT 43.900 65.200 45.800 65.500 ;
        RECT 47.000 65.400 47.400 66.200 ;
        RECT 42.900 64.600 43.700 64.900 ;
        RECT 43.300 64.200 43.700 64.600 ;
        RECT 43.300 63.800 44.200 64.200 ;
        RECT 43.300 61.100 43.700 63.800 ;
        RECT 45.500 63.500 45.800 65.200 ;
        RECT 47.700 64.900 48.000 66.800 ;
        RECT 48.300 66.500 49.000 66.900 ;
        RECT 48.700 65.500 49.000 66.500 ;
        RECT 49.400 65.800 49.800 66.600 ;
        RECT 50.200 65.800 50.600 66.600 ;
        RECT 51.800 66.400 52.200 67.200 ;
        RECT 52.700 66.200 53.000 67.900 ;
        RECT 56.600 67.400 56.900 68.500 ;
        RECT 58.700 68.000 59.100 68.800 ;
        RECT 63.300 68.000 63.700 69.500 ;
        RECT 65.400 68.500 65.800 69.500 ;
        RECT 58.700 67.700 59.500 68.000 ;
        RECT 59.100 67.500 59.500 67.700 ;
        RECT 53.400 67.100 53.800 67.200 ;
        RECT 54.200 67.100 54.600 67.200 ;
        RECT 56.600 67.100 58.700 67.400 ;
        RECT 53.400 66.800 54.600 67.100 ;
        RECT 58.200 66.900 58.700 67.100 ;
        RECT 59.200 67.200 59.500 67.500 ;
        RECT 62.900 67.700 63.700 68.000 ;
        RECT 62.900 67.500 63.300 67.700 ;
        RECT 62.900 67.200 63.200 67.500 ;
        RECT 65.500 67.400 65.800 68.500 ;
        RECT 53.400 66.600 53.700 66.800 ;
        RECT 53.300 66.200 53.700 66.600 ;
        RECT 51.000 66.100 51.400 66.200 ;
        RECT 51.000 65.800 51.800 66.100 ;
        RECT 52.600 65.800 53.000 66.200 ;
        RECT 51.400 65.600 51.800 65.800 ;
        RECT 52.700 65.700 53.000 65.800 ;
        RECT 48.700 65.200 50.600 65.500 ;
        RECT 52.700 65.400 53.700 65.700 ;
        RECT 54.200 65.400 54.600 66.200 ;
        RECT 56.600 65.800 57.000 66.600 ;
        RECT 57.400 65.800 57.800 66.600 ;
        RECT 58.200 66.500 58.900 66.900 ;
        RECT 59.200 66.800 60.200 67.200 ;
        RECT 62.200 67.100 63.200 67.200 ;
        RECT 60.600 66.800 63.200 67.100 ;
        RECT 63.700 67.100 65.800 67.400 ;
        RECT 66.200 68.500 66.600 69.500 ;
        RECT 66.200 67.400 66.500 68.500 ;
        RECT 68.300 68.000 68.700 69.500 ;
        RECT 71.000 68.500 71.400 69.500 ;
        RECT 68.300 67.700 69.100 68.000 ;
        RECT 68.700 67.500 69.100 67.700 ;
        RECT 66.200 67.100 68.300 67.400 ;
        RECT 63.700 66.900 64.200 67.100 ;
        RECT 58.200 65.500 58.500 66.500 ;
        RECT 47.700 64.600 48.500 64.900 ;
        RECT 45.400 61.500 45.800 63.500 ;
        RECT 48.100 64.200 48.500 64.600 ;
        RECT 48.100 63.800 49.000 64.200 ;
        RECT 48.100 61.100 48.500 63.800 ;
        RECT 50.300 63.500 50.600 65.200 ;
        RECT 53.400 65.100 53.700 65.400 ;
        RECT 56.600 65.200 58.500 65.500 ;
        RECT 50.200 61.500 50.600 63.500 ;
        RECT 51.000 64.800 53.000 65.100 ;
        RECT 51.000 61.100 51.400 64.800 ;
        RECT 52.600 61.400 53.000 64.800 ;
        RECT 53.400 61.700 53.800 65.100 ;
        RECT 54.200 61.400 54.600 65.100 ;
        RECT 56.600 63.500 56.900 65.200 ;
        RECT 59.200 64.900 59.500 66.800 ;
        RECT 59.800 66.100 60.200 66.200 ;
        RECT 60.600 66.100 60.900 66.800 ;
        RECT 59.800 65.800 60.900 66.100 ;
        RECT 59.800 65.400 60.200 65.800 ;
        RECT 62.200 65.400 62.600 66.200 ;
        RECT 58.700 64.600 59.500 64.900 ;
        RECT 62.900 64.900 63.200 66.800 ;
        RECT 63.500 66.500 64.200 66.900 ;
        RECT 67.800 66.900 68.300 67.100 ;
        RECT 68.800 67.200 69.100 67.500 ;
        RECT 71.000 67.400 71.300 68.500 ;
        RECT 73.100 68.000 73.500 69.500 ;
        RECT 73.100 67.700 73.900 68.000 ;
        RECT 77.300 67.900 78.100 69.900 ;
        RECT 73.500 67.500 73.900 67.700 ;
        RECT 68.800 67.100 69.800 67.200 ;
        RECT 70.200 67.100 70.600 67.200 ;
        RECT 71.000 67.100 73.100 67.400 ;
        RECT 63.900 65.500 64.200 66.500 ;
        RECT 64.600 65.800 65.000 66.600 ;
        RECT 65.400 65.800 65.800 66.600 ;
        RECT 66.200 65.800 66.600 66.600 ;
        RECT 67.000 65.800 67.400 66.600 ;
        RECT 67.800 66.500 68.500 66.900 ;
        RECT 68.800 66.800 70.600 67.100 ;
        RECT 72.600 66.900 73.100 67.100 ;
        RECT 73.600 67.200 73.900 67.500 ;
        RECT 73.600 67.100 74.600 67.200 ;
        RECT 67.800 65.500 68.100 66.500 ;
        RECT 63.900 65.200 65.800 65.500 ;
        RECT 62.900 64.600 63.700 64.900 ;
        RECT 56.600 61.500 57.000 63.500 ;
        RECT 52.600 61.100 54.600 61.400 ;
        RECT 58.700 61.100 59.100 64.600 ;
        RECT 63.300 61.100 63.700 64.600 ;
        RECT 65.500 63.500 65.800 65.200 ;
        RECT 65.400 61.500 65.800 63.500 ;
        RECT 66.200 65.200 68.100 65.500 ;
        RECT 66.200 63.500 66.500 65.200 ;
        RECT 68.800 64.900 69.100 66.800 ;
        RECT 69.400 65.400 69.800 66.200 ;
        RECT 71.000 65.800 71.400 66.600 ;
        RECT 71.800 65.800 72.200 66.600 ;
        RECT 72.600 66.500 73.300 66.900 ;
        RECT 73.600 66.800 76.100 67.100 ;
        RECT 72.600 65.500 72.900 66.500 ;
        RECT 68.300 64.600 69.100 64.900 ;
        RECT 71.000 65.200 72.900 65.500 ;
        RECT 66.200 61.500 66.600 63.500 ;
        RECT 68.300 61.100 68.700 64.600 ;
        RECT 71.000 63.500 71.300 65.200 ;
        RECT 73.600 64.900 73.900 66.800 ;
        RECT 75.800 66.200 76.100 66.800 ;
        RECT 76.600 66.400 77.000 67.200 ;
        RECT 77.500 66.200 77.800 67.900 ;
        RECT 79.800 67.500 80.200 69.900 ;
        RECT 82.000 69.200 82.400 69.900 ;
        RECT 81.400 68.900 82.400 69.200 ;
        RECT 84.200 68.900 84.600 69.900 ;
        RECT 86.300 69.200 86.900 69.900 ;
        RECT 86.200 68.900 86.900 69.200 ;
        RECT 81.400 68.500 81.800 68.900 ;
        RECT 84.200 68.600 84.500 68.900 ;
        RECT 82.200 68.200 82.600 68.600 ;
        RECT 83.100 68.300 84.500 68.600 ;
        RECT 86.200 68.500 86.600 68.900 ;
        RECT 83.100 68.200 83.500 68.300 ;
        RECT 78.200 66.800 78.600 67.200 ;
        RECT 80.200 67.100 81.000 67.200 ;
        RECT 82.300 67.100 82.600 68.200 ;
        RECT 87.100 67.700 87.500 67.800 ;
        RECT 88.600 67.700 89.000 69.900 ;
        RECT 87.100 67.400 89.000 67.700 ;
        RECT 85.100 67.100 85.500 67.200 ;
        RECT 80.200 66.800 85.700 67.100 ;
        RECT 78.200 66.600 78.500 66.800 ;
        RECT 81.700 66.700 82.100 66.800 ;
        RECT 78.100 66.200 78.500 66.600 ;
        RECT 80.900 66.200 81.300 66.300 ;
        RECT 74.200 65.400 74.600 66.200 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 75.800 65.800 76.600 66.100 ;
        RECT 77.400 65.800 77.800 66.200 ;
        RECT 76.200 65.600 76.600 65.800 ;
        RECT 77.500 65.700 77.800 65.800 ;
        RECT 77.500 65.400 78.500 65.700 ;
        RECT 79.000 65.400 79.400 66.200 ;
        RECT 80.900 65.900 83.400 66.200 ;
        RECT 83.000 65.800 83.400 65.900 ;
        RECT 79.800 65.500 82.600 65.600 ;
        RECT 79.800 65.400 82.700 65.500 ;
        RECT 78.200 65.100 78.500 65.400 ;
        RECT 79.800 65.300 84.700 65.400 ;
        RECT 73.100 64.600 73.900 64.900 ;
        RECT 75.800 64.800 77.800 65.100 ;
        RECT 71.000 61.500 71.400 63.500 ;
        RECT 73.100 61.100 73.500 64.600 ;
        RECT 75.800 61.100 76.200 64.800 ;
        RECT 77.400 61.400 77.800 64.800 ;
        RECT 78.200 61.700 78.600 65.100 ;
        RECT 79.000 61.400 79.400 65.100 ;
        RECT 77.400 61.100 79.400 61.400 ;
        RECT 79.800 61.100 80.200 65.300 ;
        RECT 82.300 65.100 84.700 65.300 ;
        RECT 81.400 64.500 84.100 64.800 ;
        RECT 81.400 64.400 81.800 64.500 ;
        RECT 83.700 64.400 84.100 64.500 ;
        RECT 84.400 64.500 84.700 65.100 ;
        RECT 85.400 65.200 85.700 66.800 ;
        RECT 86.200 66.400 86.600 66.500 ;
        RECT 86.200 66.100 88.100 66.400 ;
        RECT 87.700 66.000 88.100 66.100 ;
        RECT 86.900 65.700 87.300 65.800 ;
        RECT 88.600 65.700 89.000 67.400 ;
        RECT 89.400 68.500 89.800 69.500 ;
        RECT 89.400 67.400 89.700 68.500 ;
        RECT 91.500 68.200 91.900 69.500 ;
        RECT 91.000 68.000 91.900 68.200 ;
        RECT 91.000 67.800 92.300 68.000 ;
        RECT 91.500 67.700 92.300 67.800 ;
        RECT 91.900 67.500 92.300 67.700 ;
        RECT 89.400 67.100 91.500 67.400 ;
        RECT 91.000 66.900 91.500 67.100 ;
        RECT 92.000 67.200 92.300 67.500 ;
        RECT 89.400 65.800 89.800 66.600 ;
        RECT 90.200 65.800 90.600 66.600 ;
        RECT 91.000 66.500 91.700 66.900 ;
        RECT 92.000 66.800 93.000 67.200 ;
        RECT 86.900 65.400 89.000 65.700 ;
        RECT 91.000 65.500 91.300 66.500 ;
        RECT 85.400 64.900 86.600 65.200 ;
        RECT 85.100 64.500 85.500 64.600 ;
        RECT 84.400 64.200 85.500 64.500 ;
        RECT 86.300 64.400 86.600 64.900 ;
        RECT 86.300 64.000 87.000 64.400 ;
        RECT 83.100 63.700 83.500 63.800 ;
        RECT 84.500 63.700 84.900 63.800 ;
        RECT 81.400 63.100 81.800 63.500 ;
        RECT 83.100 63.400 84.900 63.700 ;
        RECT 84.200 63.100 84.500 63.400 ;
        RECT 86.200 63.100 86.600 63.500 ;
        RECT 81.400 62.800 82.400 63.100 ;
        RECT 82.000 61.100 82.400 62.800 ;
        RECT 84.200 61.100 84.600 63.100 ;
        RECT 86.300 61.100 86.900 63.100 ;
        RECT 88.600 61.100 89.000 65.400 ;
        RECT 89.400 65.200 91.300 65.500 ;
        RECT 89.400 63.500 89.700 65.200 ;
        RECT 92.000 64.900 92.300 66.800 ;
        RECT 92.600 66.100 93.000 66.200 ;
        RECT 94.200 66.100 94.600 69.900 ;
        RECT 97.100 69.200 97.900 69.900 ;
        RECT 96.600 68.800 97.900 69.200 ;
        RECT 95.000 67.800 95.400 68.600 ;
        RECT 97.100 67.900 97.900 68.800 ;
        RECT 101.700 68.000 102.100 69.500 ;
        RECT 103.800 68.500 104.200 69.500 ;
        RECT 95.000 67.100 95.400 67.200 ;
        RECT 96.600 67.100 97.000 67.200 ;
        RECT 95.000 66.800 97.000 67.100 ;
        RECT 96.700 66.600 97.000 66.800 ;
        RECT 96.700 66.200 97.100 66.600 ;
        RECT 97.400 66.200 97.700 67.900 ;
        RECT 101.300 67.700 102.100 68.000 ;
        RECT 101.300 67.500 101.700 67.700 ;
        RECT 101.300 67.200 101.600 67.500 ;
        RECT 103.900 67.400 104.200 68.500 ;
        RECT 98.200 66.400 98.600 67.200 ;
        RECT 100.600 67.100 101.600 67.200 ;
        RECT 99.000 66.800 101.600 67.100 ;
        RECT 102.100 67.100 104.200 67.400 ;
        RECT 106.200 68.500 106.600 69.500 ;
        RECT 106.200 67.400 106.500 68.500 ;
        RECT 108.300 68.000 108.700 69.500 ;
        RECT 111.300 68.200 111.700 69.900 ;
        RECT 113.400 68.500 113.800 69.500 ;
        RECT 108.300 67.700 109.100 68.000 ;
        RECT 111.300 67.900 112.200 68.200 ;
        RECT 108.700 67.500 109.100 67.700 ;
        RECT 106.200 67.100 108.300 67.400 ;
        RECT 102.100 66.900 102.600 67.100 ;
        RECT 99.000 66.200 99.300 66.800 ;
        RECT 92.600 65.800 94.600 66.100 ;
        RECT 92.600 65.400 93.000 65.800 ;
        RECT 91.500 64.600 92.300 64.900 ;
        RECT 89.400 61.500 89.800 63.500 ;
        RECT 91.500 61.100 91.900 64.600 ;
        RECT 94.200 61.100 94.600 65.800 ;
        RECT 95.800 65.400 96.200 66.200 ;
        RECT 97.400 65.800 97.800 66.200 ;
        RECT 99.000 66.100 99.400 66.200 ;
        RECT 98.600 65.800 99.400 66.100 ;
        RECT 97.400 65.700 97.700 65.800 ;
        RECT 96.700 65.400 97.700 65.700 ;
        RECT 98.600 65.600 99.000 65.800 ;
        RECT 100.600 65.400 101.000 66.200 ;
        RECT 96.700 65.100 97.000 65.400 ;
        RECT 95.800 61.400 96.200 65.100 ;
        RECT 96.600 61.700 97.000 65.100 ;
        RECT 97.400 64.800 99.400 65.100 ;
        RECT 97.400 61.400 97.800 64.800 ;
        RECT 95.800 61.100 97.800 61.400 ;
        RECT 99.000 61.100 99.400 64.800 ;
        RECT 101.300 64.900 101.600 66.800 ;
        RECT 101.900 66.500 102.600 66.900 ;
        RECT 107.800 66.900 108.300 67.100 ;
        RECT 108.800 67.200 109.100 67.500 ;
        RECT 108.800 67.100 109.800 67.200 ;
        RECT 111.000 67.100 111.400 67.200 ;
        RECT 102.300 65.500 102.600 66.500 ;
        RECT 103.000 65.800 103.400 66.600 ;
        RECT 103.800 65.800 104.200 66.600 ;
        RECT 106.200 65.800 106.600 66.600 ;
        RECT 107.000 65.800 107.400 66.600 ;
        RECT 107.800 66.500 108.500 66.900 ;
        RECT 108.800 66.800 111.400 67.100 ;
        RECT 107.800 65.500 108.100 66.500 ;
        RECT 102.300 65.200 104.200 65.500 ;
        RECT 101.300 64.600 102.100 64.900 ;
        RECT 101.700 61.100 102.100 64.600 ;
        RECT 103.900 63.500 104.200 65.200 ;
        RECT 103.800 61.500 104.200 63.500 ;
        RECT 106.200 65.200 108.100 65.500 ;
        RECT 106.200 63.500 106.500 65.200 ;
        RECT 108.800 64.900 109.100 66.800 ;
        RECT 109.400 66.100 109.800 66.200 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 109.400 65.800 110.600 66.100 ;
        RECT 109.400 65.400 109.800 65.800 ;
        RECT 108.300 64.600 109.100 64.900 ;
        RECT 106.200 61.500 106.600 63.500 ;
        RECT 108.300 61.100 108.700 64.600 ;
        RECT 111.000 64.400 111.400 65.200 ;
        RECT 111.800 61.100 112.200 67.900 ;
        RECT 112.600 66.800 113.000 67.600 ;
        RECT 113.400 67.400 113.700 68.500 ;
        RECT 115.500 68.000 115.900 69.500 ;
        RECT 118.200 68.500 118.600 69.500 ;
        RECT 115.500 67.700 116.300 68.000 ;
        RECT 115.900 67.500 116.300 67.700 ;
        RECT 113.400 67.100 115.500 67.400 ;
        RECT 115.000 66.900 115.500 67.100 ;
        RECT 116.000 67.200 116.300 67.500 ;
        RECT 118.200 67.400 118.500 68.500 ;
        RECT 120.300 68.000 120.700 69.500 ;
        RECT 124.300 69.200 124.700 69.900 ;
        RECT 124.300 68.800 125.000 69.200 ;
        RECT 124.300 68.200 124.700 68.800 ;
        RECT 120.300 67.700 121.100 68.000 ;
        RECT 120.700 67.500 121.100 67.700 ;
        RECT 123.800 67.900 124.700 68.200 ;
        RECT 126.700 67.900 127.500 69.900 ;
        RECT 130.700 69.200 131.500 69.900 ;
        RECT 130.200 68.800 131.500 69.200 ;
        RECT 130.700 67.900 131.500 68.800 ;
        RECT 135.300 68.000 135.700 69.500 ;
        RECT 137.400 68.500 137.800 69.500 ;
        RECT 116.000 67.100 117.000 67.200 ;
        RECT 117.400 67.100 117.800 67.200 ;
        RECT 118.200 67.100 120.300 67.400 ;
        RECT 113.400 65.800 113.800 66.600 ;
        RECT 114.200 65.800 114.600 66.600 ;
        RECT 115.000 66.500 115.700 66.900 ;
        RECT 116.000 66.800 117.800 67.100 ;
        RECT 119.800 66.900 120.300 67.100 ;
        RECT 120.800 67.200 121.100 67.500 ;
        RECT 120.800 67.100 121.800 67.200 ;
        RECT 122.200 67.100 122.600 67.200 ;
        RECT 115.000 65.500 115.300 66.500 ;
        RECT 113.400 65.200 115.300 65.500 ;
        RECT 113.400 63.500 113.700 65.200 ;
        RECT 116.000 64.900 116.300 66.800 ;
        RECT 116.600 65.400 117.000 66.200 ;
        RECT 118.200 65.800 118.600 66.600 ;
        RECT 119.000 65.800 119.400 66.600 ;
        RECT 119.800 66.500 120.500 66.900 ;
        RECT 120.800 66.800 122.600 67.100 ;
        RECT 123.000 66.800 123.400 67.600 ;
        RECT 119.800 65.500 120.100 66.500 ;
        RECT 115.500 64.600 116.300 64.900 ;
        RECT 118.200 65.200 120.100 65.500 ;
        RECT 113.400 61.500 113.800 63.500 ;
        RECT 115.500 61.100 115.900 64.600 ;
        RECT 118.200 63.500 118.500 65.200 ;
        RECT 120.800 64.900 121.100 66.800 ;
        RECT 121.400 65.400 121.800 66.200 ;
        RECT 120.300 64.600 121.100 64.900 ;
        RECT 118.200 61.500 118.600 63.500 ;
        RECT 120.300 61.100 120.700 64.600 ;
        RECT 123.800 61.100 124.200 67.900 ;
        RECT 126.200 66.800 126.600 67.200 ;
        RECT 126.300 66.600 126.600 66.800 ;
        RECT 126.300 66.200 126.700 66.600 ;
        RECT 127.000 66.200 127.300 67.900 ;
        RECT 127.800 66.400 128.200 67.200 ;
        RECT 129.400 67.100 129.800 67.200 ;
        RECT 130.200 67.100 130.600 67.200 ;
        RECT 129.400 66.800 130.600 67.100 ;
        RECT 130.300 66.600 130.600 66.800 ;
        RECT 130.300 66.200 130.700 66.600 ;
        RECT 131.000 66.200 131.300 67.900 ;
        RECT 134.900 67.700 135.700 68.000 ;
        RECT 134.900 67.500 135.300 67.700 ;
        RECT 134.900 67.200 135.200 67.500 ;
        RECT 137.500 67.400 137.800 68.500 ;
        RECT 131.800 66.400 132.200 67.200 ;
        RECT 134.200 67.100 135.200 67.200 ;
        RECT 132.600 66.800 135.200 67.100 ;
        RECT 135.700 67.100 137.800 67.400 ;
        RECT 139.800 67.900 140.200 69.900 ;
        RECT 140.500 68.200 140.900 68.600 ;
        RECT 135.700 66.900 136.200 67.100 ;
        RECT 132.600 66.200 132.900 66.800 ;
        RECT 125.400 65.400 125.800 66.200 ;
        RECT 127.000 65.800 127.400 66.200 ;
        RECT 128.600 66.100 129.000 66.200 ;
        RECT 128.200 65.800 129.000 66.100 ;
        RECT 127.000 65.700 127.300 65.800 ;
        RECT 126.300 65.400 127.300 65.700 ;
        RECT 128.200 65.600 128.600 65.800 ;
        RECT 129.400 65.400 129.800 66.200 ;
        RECT 131.000 65.800 131.400 66.200 ;
        RECT 132.600 66.100 133.000 66.200 ;
        RECT 132.200 65.800 133.000 66.100 ;
        RECT 131.000 65.700 131.300 65.800 ;
        RECT 130.300 65.400 131.300 65.700 ;
        RECT 132.200 65.600 132.600 65.800 ;
        RECT 134.200 65.400 134.600 66.200 ;
        RECT 124.600 64.400 125.000 65.200 ;
        RECT 126.300 65.100 126.600 65.400 ;
        RECT 130.300 65.100 130.600 65.400 ;
        RECT 125.400 61.400 125.800 65.100 ;
        RECT 126.200 61.700 126.600 65.100 ;
        RECT 127.000 64.800 129.000 65.100 ;
        RECT 127.000 61.400 127.400 64.800 ;
        RECT 125.400 61.100 127.400 61.400 ;
        RECT 128.600 61.100 129.000 64.800 ;
        RECT 129.400 61.400 129.800 65.100 ;
        RECT 130.200 61.700 130.600 65.100 ;
        RECT 131.000 64.800 133.000 65.100 ;
        RECT 131.000 61.400 131.400 64.800 ;
        RECT 129.400 61.100 131.400 61.400 ;
        RECT 132.600 61.100 133.000 64.800 ;
        RECT 134.900 64.900 135.200 66.800 ;
        RECT 135.500 66.500 136.200 66.900 ;
        RECT 135.900 65.500 136.200 66.500 ;
        RECT 136.600 65.800 137.000 66.600 ;
        RECT 137.400 65.800 137.800 66.600 ;
        RECT 139.000 66.400 139.400 67.200 ;
        RECT 138.200 66.100 138.600 66.200 ;
        RECT 139.800 66.100 140.100 67.900 ;
        RECT 140.600 67.800 141.000 68.200 ;
        RECT 142.200 67.600 142.600 69.900 ;
        RECT 143.800 67.600 144.200 69.900 ;
        RECT 145.400 67.600 145.800 69.900 ;
        RECT 147.000 67.600 147.400 69.900 ;
        RECT 148.600 68.000 149.000 69.900 ;
        RECT 150.200 68.000 150.600 69.900 ;
        RECT 148.600 67.900 150.600 68.000 ;
        RECT 151.000 67.900 151.400 69.900 ;
        RECT 153.700 68.000 154.100 69.500 ;
        RECT 155.800 68.500 156.200 69.500 ;
        RECT 148.700 67.700 150.500 67.900 ;
        RECT 141.400 67.200 142.600 67.600 ;
        RECT 143.100 67.200 144.200 67.600 ;
        RECT 144.700 67.200 145.800 67.600 ;
        RECT 146.500 67.200 147.400 67.600 ;
        RECT 149.000 67.200 149.400 67.400 ;
        RECT 151.000 67.200 151.300 67.900 ;
        RECT 153.300 67.700 154.100 68.000 ;
        RECT 153.300 67.500 153.700 67.700 ;
        RECT 153.300 67.200 153.600 67.500 ;
        RECT 155.900 67.400 156.200 68.500 ;
        RECT 158.500 68.200 158.900 69.900 ;
        RECT 157.400 68.100 157.800 68.200 ;
        RECT 158.500 68.100 159.400 68.200 ;
        RECT 157.400 67.800 159.400 68.100 ;
        RECT 161.900 67.900 162.700 69.900 ;
        RECT 165.900 69.200 166.300 69.900 ;
        RECT 165.400 68.800 166.300 69.200 ;
        RECT 165.900 68.200 166.300 68.800 ;
        RECT 165.400 67.900 166.300 68.200 ;
        RECT 168.500 67.900 169.300 69.900 ;
        RECT 140.600 66.100 141.000 66.200 ;
        RECT 138.200 65.800 139.000 66.100 ;
        RECT 139.800 65.800 141.000 66.100 ;
        RECT 141.400 65.800 141.800 67.200 ;
        RECT 143.100 66.900 143.500 67.200 ;
        RECT 144.700 66.900 145.100 67.200 ;
        RECT 146.500 66.900 146.900 67.200 ;
        RECT 142.200 66.500 143.500 66.900 ;
        RECT 143.900 66.500 145.100 66.900 ;
        RECT 145.600 66.500 146.900 66.900 ;
        RECT 148.600 66.900 149.400 67.200 ;
        RECT 148.600 66.800 149.000 66.900 ;
        RECT 150.100 66.800 151.400 67.200 ;
        RECT 152.600 67.100 153.600 67.200 ;
        RECT 151.800 66.800 153.600 67.100 ;
        RECT 154.100 67.100 156.200 67.400 ;
        RECT 154.100 66.900 154.600 67.100 ;
        RECT 143.100 65.800 143.500 66.500 ;
        RECT 144.700 65.800 145.100 66.500 ;
        RECT 146.500 65.800 146.900 66.500 ;
        RECT 149.400 65.800 149.800 66.600 ;
        RECT 138.600 65.600 139.000 65.800 ;
        RECT 135.900 65.200 137.800 65.500 ;
        RECT 134.900 64.600 135.700 64.900 ;
        RECT 135.300 61.100 135.700 64.600 ;
        RECT 137.500 63.500 137.800 65.200 ;
        RECT 140.600 65.100 140.900 65.800 ;
        RECT 141.400 65.400 142.600 65.800 ;
        RECT 143.100 65.400 144.200 65.800 ;
        RECT 144.700 65.400 145.800 65.800 ;
        RECT 146.500 65.400 147.400 65.800 ;
        RECT 137.400 61.500 137.800 63.500 ;
        RECT 138.200 64.800 140.200 65.100 ;
        RECT 138.200 61.100 138.600 64.800 ;
        RECT 139.800 61.100 140.200 64.800 ;
        RECT 140.600 61.100 141.000 65.100 ;
        RECT 142.200 61.100 142.600 65.400 ;
        RECT 143.800 61.100 144.200 65.400 ;
        RECT 145.400 61.100 145.800 65.400 ;
        RECT 147.000 61.100 147.400 65.400 ;
        RECT 150.100 65.100 150.400 66.800 ;
        RECT 151.800 66.200 152.100 66.800 ;
        RECT 151.800 65.800 152.200 66.200 ;
        RECT 152.600 65.400 153.000 66.200 ;
        RECT 151.000 65.100 151.400 65.200 ;
        RECT 149.900 64.800 150.400 65.100 ;
        RECT 150.700 64.800 151.400 65.100 ;
        RECT 153.300 64.900 153.600 66.800 ;
        RECT 153.900 66.500 154.600 66.900 ;
        RECT 154.300 65.500 154.600 66.500 ;
        RECT 155.000 65.800 155.400 66.600 ;
        RECT 155.800 65.800 156.200 66.600 ;
        RECT 154.300 65.200 156.200 65.500 ;
        RECT 149.900 61.100 150.300 64.800 ;
        RECT 150.700 64.200 151.000 64.800 ;
        RECT 153.300 64.600 154.100 64.900 ;
        RECT 150.600 63.800 151.000 64.200 ;
        RECT 153.700 61.100 154.100 64.600 ;
        RECT 155.900 63.500 156.200 65.200 ;
        RECT 158.200 64.400 158.600 65.200 ;
        RECT 155.800 61.500 156.200 63.500 ;
        RECT 159.000 61.100 159.400 67.800 ;
        RECT 159.800 67.100 160.200 67.600 ;
        RECT 162.200 67.200 162.500 67.900 ;
        RECT 160.600 67.100 161.000 67.200 ;
        RECT 159.800 66.800 161.000 67.100 ;
        RECT 161.400 66.800 161.800 67.200 ;
        RECT 161.500 66.600 161.800 66.800 ;
        RECT 162.200 66.800 162.600 67.200 ;
        RECT 161.500 66.200 161.900 66.600 ;
        RECT 162.200 66.200 162.500 66.800 ;
        RECT 163.000 66.400 163.400 67.200 ;
        RECT 164.600 66.800 165.000 67.600 ;
        RECT 159.800 66.100 160.200 66.200 ;
        RECT 160.600 66.100 161.000 66.200 ;
        RECT 159.800 65.800 161.000 66.100 ;
        RECT 160.600 65.400 161.000 65.800 ;
        RECT 162.200 65.800 162.600 66.200 ;
        RECT 163.800 66.100 164.200 66.200 ;
        RECT 163.400 65.800 164.200 66.100 ;
        RECT 162.200 65.700 162.500 65.800 ;
        RECT 161.500 65.400 162.500 65.700 ;
        RECT 163.400 65.600 163.800 65.800 ;
        RECT 161.500 65.100 161.800 65.400 ;
        RECT 160.600 61.400 161.000 65.100 ;
        RECT 161.400 61.700 161.800 65.100 ;
        RECT 162.200 64.800 164.200 65.100 ;
        RECT 162.200 61.400 162.600 64.800 ;
        RECT 160.600 61.100 162.600 61.400 ;
        RECT 163.800 61.100 164.200 64.800 ;
        RECT 165.400 61.100 165.800 67.900 ;
        RECT 167.800 66.400 168.200 67.200 ;
        RECT 168.700 66.200 169.000 67.900 ;
        RECT 171.000 67.700 171.400 69.900 ;
        RECT 173.100 69.200 173.700 69.900 ;
        RECT 173.100 68.900 173.800 69.200 ;
        RECT 175.400 68.900 175.800 69.900 ;
        RECT 177.600 69.200 178.000 69.900 ;
        RECT 177.600 68.900 178.600 69.200 ;
        RECT 173.400 68.500 173.800 68.900 ;
        RECT 175.500 68.600 175.800 68.900 ;
        RECT 175.500 68.300 176.900 68.600 ;
        RECT 176.500 68.200 176.900 68.300 ;
        RECT 177.400 68.200 177.800 68.600 ;
        RECT 178.200 68.500 178.600 68.900 ;
        RECT 172.500 67.700 172.900 67.800 ;
        RECT 171.000 67.400 172.900 67.700 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 169.400 66.600 169.700 66.800 ;
        RECT 169.300 66.200 169.700 66.600 ;
        RECT 167.000 66.100 167.400 66.200 ;
        RECT 167.000 65.800 167.800 66.100 ;
        RECT 168.600 65.800 169.000 66.200 ;
        RECT 167.400 65.600 167.800 65.800 ;
        RECT 168.700 65.700 169.000 65.800 ;
        RECT 168.700 65.400 169.700 65.700 ;
        RECT 170.200 65.400 170.600 66.200 ;
        RECT 171.000 65.700 171.400 67.400 ;
        RECT 174.500 67.100 174.900 67.200 ;
        RECT 177.400 67.100 177.700 68.200 ;
        RECT 179.800 67.500 180.200 69.900 ;
        RECT 181.900 68.200 182.300 69.900 ;
        RECT 181.400 67.900 182.300 68.200 ;
        RECT 183.000 67.900 183.400 69.900 ;
        RECT 183.800 68.000 184.200 69.900 ;
        RECT 185.400 68.000 185.800 69.900 ;
        RECT 187.000 68.200 187.400 69.900 ;
        RECT 183.800 67.900 185.800 68.000 ;
        RECT 186.900 67.900 187.400 68.200 ;
        RECT 179.000 67.100 179.800 67.200 ;
        RECT 174.300 66.800 179.800 67.100 ;
        RECT 180.600 66.800 181.000 67.600 ;
        RECT 173.400 66.400 173.800 66.500 ;
        RECT 171.900 66.100 173.800 66.400 ;
        RECT 174.300 66.200 174.600 66.800 ;
        RECT 177.900 66.700 178.300 66.800 ;
        RECT 177.400 66.200 177.800 66.300 ;
        RECT 178.700 66.200 179.100 66.300 ;
        RECT 171.900 66.000 172.300 66.100 ;
        RECT 174.200 65.800 174.600 66.200 ;
        RECT 176.600 65.900 179.100 66.200 ;
        RECT 181.400 66.100 181.800 67.900 ;
        RECT 183.100 67.200 183.400 67.900 ;
        RECT 183.900 67.700 185.700 67.900 ;
        RECT 185.000 67.200 185.400 67.400 ;
        RECT 186.900 67.200 187.200 67.900 ;
        RECT 188.600 67.600 189.000 69.900 ;
        RECT 187.700 67.300 189.000 67.600 ;
        RECT 190.200 67.600 190.600 69.900 ;
        RECT 191.800 67.600 192.200 69.900 ;
        RECT 193.400 67.600 193.800 69.900 ;
        RECT 195.000 67.600 195.400 69.900 ;
        RECT 198.100 67.900 198.900 69.900 ;
        RECT 200.900 69.200 201.300 69.900 ;
        RECT 200.600 68.800 201.300 69.200 ;
        RECT 200.900 68.200 201.300 68.800 ;
        RECT 204.300 68.200 205.100 69.900 ;
        RECT 200.900 67.900 201.800 68.200 ;
        RECT 183.000 66.800 184.300 67.200 ;
        RECT 185.000 67.100 185.800 67.200 ;
        RECT 186.900 67.100 187.400 67.200 ;
        RECT 185.000 66.900 187.400 67.100 ;
        RECT 185.400 66.800 187.400 66.900 ;
        RECT 176.600 65.800 177.000 65.900 ;
        RECT 181.400 65.800 183.300 66.100 ;
        RECT 172.700 65.700 173.100 65.800 ;
        RECT 171.000 65.400 173.100 65.700 ;
        RECT 166.200 64.400 166.600 65.200 ;
        RECT 169.400 65.100 169.700 65.400 ;
        RECT 167.000 64.800 169.000 65.100 ;
        RECT 167.000 61.100 167.400 64.800 ;
        RECT 168.600 61.400 169.000 64.800 ;
        RECT 169.400 61.700 169.800 65.100 ;
        RECT 170.200 61.400 170.600 65.100 ;
        RECT 168.600 61.100 170.600 61.400 ;
        RECT 171.000 61.100 171.400 65.400 ;
        RECT 174.300 65.200 174.600 65.800 ;
        RECT 177.400 65.500 180.200 65.600 ;
        RECT 177.300 65.400 180.200 65.500 ;
        RECT 173.400 64.900 174.600 65.200 ;
        RECT 175.300 65.300 180.200 65.400 ;
        RECT 175.300 65.100 177.700 65.300 ;
        RECT 173.400 64.400 173.700 64.900 ;
        RECT 173.000 64.000 173.700 64.400 ;
        RECT 174.500 64.500 174.900 64.600 ;
        RECT 175.300 64.500 175.600 65.100 ;
        RECT 174.500 64.200 175.600 64.500 ;
        RECT 175.900 64.500 178.600 64.800 ;
        RECT 175.900 64.400 176.300 64.500 ;
        RECT 178.200 64.400 178.600 64.500 ;
        RECT 175.100 63.700 175.500 63.800 ;
        RECT 176.500 63.700 176.900 63.800 ;
        RECT 173.400 63.100 173.800 63.500 ;
        RECT 175.100 63.400 176.900 63.700 ;
        RECT 175.500 63.100 175.800 63.400 ;
        RECT 178.200 63.100 178.600 63.500 ;
        RECT 173.100 61.100 173.700 63.100 ;
        RECT 175.400 61.100 175.800 63.100 ;
        RECT 177.600 62.800 178.600 63.100 ;
        RECT 177.600 61.100 178.000 62.800 ;
        RECT 179.800 61.100 180.200 65.300 ;
        RECT 181.400 61.100 181.800 65.800 ;
        RECT 183.000 65.200 183.300 65.800 ;
        RECT 182.200 64.400 182.600 65.200 ;
        RECT 183.000 65.100 183.400 65.200 ;
        RECT 184.000 65.100 184.300 66.800 ;
        RECT 184.600 65.800 185.000 66.600 ;
        RECT 186.900 65.100 187.200 66.800 ;
        RECT 187.700 66.500 188.000 67.300 ;
        RECT 190.200 67.200 191.100 67.600 ;
        RECT 191.800 67.200 192.900 67.600 ;
        RECT 193.400 67.200 194.500 67.600 ;
        RECT 195.000 67.200 196.200 67.600 ;
        RECT 189.400 66.900 189.800 67.200 ;
        RECT 190.700 66.900 191.100 67.200 ;
        RECT 192.500 66.900 192.900 67.200 ;
        RECT 194.100 66.900 194.500 67.200 ;
        RECT 187.500 66.100 188.000 66.500 ;
        RECT 187.700 65.100 188.000 66.100 ;
        RECT 188.500 66.200 188.900 66.600 ;
        RECT 189.400 66.500 190.300 66.900 ;
        RECT 190.700 66.500 192.000 66.900 ;
        RECT 192.500 66.500 193.700 66.900 ;
        RECT 194.100 66.500 195.400 66.900 ;
        RECT 188.500 65.800 189.000 66.200 ;
        RECT 190.700 65.800 191.100 66.500 ;
        RECT 192.500 65.800 192.900 66.500 ;
        RECT 194.100 65.800 194.500 66.500 ;
        RECT 195.800 65.800 196.200 67.200 ;
        RECT 197.400 66.400 197.800 67.200 ;
        RECT 198.300 66.200 198.600 67.900 ;
        RECT 199.000 67.100 199.400 67.200 ;
        RECT 200.600 67.100 201.000 67.200 ;
        RECT 199.000 66.800 201.000 67.100 ;
        RECT 199.000 66.600 199.300 66.800 ;
        RECT 198.900 66.200 199.300 66.600 ;
        RECT 196.600 66.100 197.000 66.200 ;
        RECT 196.600 65.800 197.400 66.100 ;
        RECT 198.200 65.800 198.600 66.200 ;
        RECT 190.200 65.400 191.100 65.800 ;
        RECT 191.800 65.400 192.900 65.800 ;
        RECT 193.400 65.400 194.500 65.800 ;
        RECT 195.000 65.400 196.200 65.800 ;
        RECT 197.000 65.600 197.400 65.800 ;
        RECT 198.300 65.700 198.600 65.800 ;
        RECT 198.300 65.400 199.300 65.700 ;
        RECT 199.800 65.400 200.200 66.200 ;
        RECT 183.000 64.800 183.700 65.100 ;
        RECT 184.000 64.800 184.500 65.100 ;
        RECT 183.400 64.200 183.700 64.800 ;
        RECT 183.400 63.800 183.800 64.200 ;
        RECT 184.100 61.100 184.500 64.800 ;
        RECT 186.900 64.600 187.400 65.100 ;
        RECT 187.700 64.800 189.000 65.100 ;
        RECT 187.000 61.100 187.400 64.600 ;
        RECT 188.600 61.100 189.000 64.800 ;
        RECT 190.200 61.100 190.600 65.400 ;
        RECT 191.800 61.100 192.200 65.400 ;
        RECT 193.400 61.100 193.800 65.400 ;
        RECT 195.000 61.100 195.400 65.400 ;
        RECT 199.000 65.200 199.300 65.400 ;
        RECT 196.600 64.800 198.600 65.100 ;
        RECT 196.600 61.100 197.000 64.800 ;
        RECT 198.200 61.400 198.600 64.800 ;
        RECT 199.000 61.700 199.400 65.200 ;
        RECT 199.800 61.400 200.200 65.100 ;
        RECT 200.600 64.400 201.000 65.200 ;
        RECT 198.200 61.100 200.200 61.400 ;
        RECT 201.400 61.100 201.800 67.900 ;
        RECT 203.800 67.900 205.100 68.200 ;
        RECT 210.100 67.900 210.900 69.900 ;
        RECT 212.900 69.200 213.300 69.900 ;
        RECT 212.600 68.800 213.300 69.200 ;
        RECT 212.900 68.200 213.300 68.800 ;
        RECT 216.300 68.200 217.100 69.900 ;
        RECT 212.900 67.900 213.800 68.200 ;
        RECT 203.800 67.800 204.900 67.900 ;
        RECT 202.200 67.100 202.600 67.600 ;
        RECT 203.000 67.100 203.400 67.200 ;
        RECT 202.200 66.800 203.400 67.100 ;
        RECT 203.800 66.800 204.200 67.200 ;
        RECT 203.900 66.600 204.200 66.800 ;
        RECT 203.900 66.200 204.300 66.600 ;
        RECT 204.600 66.200 204.900 67.800 ;
        RECT 205.400 66.400 205.800 67.200 ;
        RECT 207.000 67.100 207.400 67.200 ;
        RECT 209.400 67.100 209.800 67.200 ;
        RECT 207.000 66.800 209.800 67.100 ;
        RECT 209.400 66.400 209.800 66.800 ;
        RECT 210.300 66.200 210.600 67.900 ;
        RECT 211.000 66.800 211.400 67.200 ;
        RECT 211.000 66.600 211.300 66.800 ;
        RECT 210.900 66.200 211.300 66.600 ;
        RECT 203.000 65.400 203.400 66.200 ;
        RECT 204.600 65.800 205.000 66.200 ;
        RECT 206.200 66.100 206.600 66.200 ;
        RECT 207.800 66.100 208.200 66.200 ;
        RECT 205.800 65.800 208.200 66.100 ;
        RECT 208.600 66.100 209.000 66.200 ;
        RECT 208.600 65.800 209.400 66.100 ;
        RECT 210.200 65.800 210.600 66.200 ;
        RECT 204.600 65.700 204.900 65.800 ;
        RECT 203.900 65.400 204.900 65.700 ;
        RECT 205.800 65.600 206.200 65.800 ;
        RECT 209.000 65.600 209.400 65.800 ;
        RECT 210.300 65.700 210.600 65.800 ;
        RECT 210.300 65.400 211.300 65.700 ;
        RECT 211.800 65.400 212.200 66.200 ;
        RECT 203.900 65.100 204.200 65.400 ;
        RECT 211.000 65.100 211.300 65.400 ;
        RECT 203.000 61.400 203.400 65.100 ;
        RECT 203.800 61.700 204.200 65.100 ;
        RECT 204.600 64.800 206.600 65.100 ;
        RECT 204.600 61.400 205.000 64.800 ;
        RECT 203.000 61.100 205.000 61.400 ;
        RECT 206.200 61.100 206.600 64.800 ;
        RECT 208.600 64.800 210.600 65.100 ;
        RECT 208.600 61.100 209.000 64.800 ;
        RECT 210.200 61.400 210.600 64.800 ;
        RECT 211.000 61.700 211.400 65.100 ;
        RECT 211.800 61.400 212.200 65.100 ;
        RECT 212.600 64.400 213.000 65.200 ;
        RECT 210.200 61.100 212.200 61.400 ;
        RECT 213.400 61.100 213.800 67.900 ;
        RECT 215.800 67.900 217.100 68.200 ;
        RECT 220.900 68.000 221.300 69.500 ;
        RECT 223.000 68.500 223.400 69.500 ;
        RECT 215.800 67.800 216.900 67.900 ;
        RECT 214.200 67.100 214.600 67.600 ;
        RECT 215.000 67.100 215.400 67.200 ;
        RECT 214.200 66.800 215.400 67.100 ;
        RECT 215.800 66.800 216.200 67.200 ;
        RECT 215.900 66.600 216.200 66.800 ;
        RECT 215.900 66.200 216.300 66.600 ;
        RECT 216.600 66.200 216.900 67.800 ;
        RECT 220.500 67.700 221.300 68.000 ;
        RECT 220.500 67.500 220.900 67.700 ;
        RECT 220.500 67.200 220.800 67.500 ;
        RECT 223.100 67.400 223.400 68.500 ;
        RECT 217.400 66.400 217.800 67.200 ;
        RECT 219.800 67.100 220.800 67.200 ;
        RECT 218.200 66.800 220.800 67.100 ;
        RECT 221.300 67.100 223.400 67.400 ;
        RECT 223.800 68.500 224.200 69.500 ;
        RECT 223.800 67.400 224.100 68.500 ;
        RECT 225.900 68.200 226.300 69.500 ;
        RECT 225.400 68.000 226.300 68.200 ;
        RECT 225.400 67.800 226.700 68.000 ;
        RECT 225.900 67.700 226.700 67.800 ;
        RECT 226.300 67.500 226.700 67.700 ;
        RECT 228.600 67.500 229.000 69.900 ;
        RECT 230.800 69.200 231.200 69.900 ;
        RECT 230.200 68.900 231.200 69.200 ;
        RECT 233.000 68.900 233.400 69.900 ;
        RECT 235.100 69.200 235.700 69.900 ;
        RECT 235.000 68.900 235.700 69.200 ;
        RECT 230.200 68.500 230.600 68.900 ;
        RECT 233.000 68.600 233.300 68.900 ;
        RECT 231.000 67.800 231.400 68.600 ;
        RECT 231.900 68.300 233.300 68.600 ;
        RECT 235.000 68.500 235.400 68.900 ;
        RECT 231.900 68.200 232.300 68.300 ;
        RECT 234.200 68.100 234.600 68.200 ;
        RECT 234.200 67.800 236.200 68.100 ;
        RECT 223.800 67.100 225.900 67.400 ;
        RECT 221.300 66.900 221.800 67.100 ;
        RECT 218.200 66.200 218.500 66.800 ;
        RECT 215.000 65.400 215.400 66.200 ;
        RECT 216.600 65.800 217.000 66.200 ;
        RECT 218.200 66.100 218.600 66.200 ;
        RECT 217.800 65.800 218.600 66.100 ;
        RECT 219.000 66.100 219.400 66.200 ;
        RECT 219.800 66.100 220.200 66.200 ;
        RECT 219.000 65.800 220.200 66.100 ;
        RECT 216.600 65.700 216.900 65.800 ;
        RECT 215.900 65.400 216.900 65.700 ;
        RECT 217.800 65.600 218.200 65.800 ;
        RECT 219.800 65.400 220.200 65.800 ;
        RECT 215.900 65.100 216.200 65.400 ;
        RECT 215.000 61.400 215.400 65.100 ;
        RECT 215.800 61.700 216.200 65.100 ;
        RECT 216.600 64.800 218.600 65.100 ;
        RECT 216.600 61.400 217.000 64.800 ;
        RECT 215.000 61.100 217.000 61.400 ;
        RECT 218.200 61.100 218.600 64.800 ;
        RECT 220.500 64.900 220.800 66.800 ;
        RECT 221.100 66.500 221.800 66.900 ;
        RECT 225.400 66.900 225.900 67.100 ;
        RECT 226.400 67.200 226.700 67.500 ;
        RECT 221.500 65.500 221.800 66.500 ;
        RECT 222.200 65.800 222.600 66.600 ;
        RECT 223.000 66.100 223.400 66.600 ;
        RECT 223.800 66.100 224.200 66.600 ;
        RECT 223.000 65.800 224.200 66.100 ;
        RECT 224.600 65.800 225.000 66.600 ;
        RECT 225.400 66.500 226.100 66.900 ;
        RECT 226.400 66.800 227.400 67.200 ;
        RECT 229.000 67.100 229.800 67.200 ;
        RECT 231.100 67.100 231.400 67.800 ;
        RECT 235.800 67.700 236.300 67.800 ;
        RECT 237.400 67.700 237.800 69.900 ;
        RECT 240.100 68.000 240.500 69.500 ;
        RECT 242.200 68.500 242.600 69.500 ;
        RECT 235.800 67.400 237.800 67.700 ;
        RECT 233.900 67.100 234.300 67.200 ;
        RECT 229.000 66.800 234.500 67.100 ;
        RECT 225.400 65.500 225.700 66.500 ;
        RECT 221.500 65.200 223.400 65.500 ;
        RECT 220.500 64.600 221.300 64.900 ;
        RECT 220.900 61.100 221.300 64.600 ;
        RECT 223.100 63.500 223.400 65.200 ;
        RECT 223.000 61.500 223.400 63.500 ;
        RECT 223.800 65.200 225.700 65.500 ;
        RECT 223.800 63.500 224.100 65.200 ;
        RECT 226.400 64.900 226.700 66.800 ;
        RECT 230.500 66.700 230.900 66.800 ;
        RECT 229.700 66.200 230.100 66.300 ;
        RECT 227.000 66.100 227.400 66.200 ;
        RECT 227.800 66.100 228.200 66.200 ;
        RECT 227.000 65.800 228.200 66.100 ;
        RECT 229.700 65.900 232.200 66.200 ;
        RECT 231.800 65.800 232.200 65.900 ;
        RECT 233.400 66.100 233.800 66.200 ;
        RECT 234.200 66.100 234.500 66.800 ;
        RECT 235.000 66.400 235.400 66.500 ;
        RECT 235.000 66.100 236.900 66.400 ;
        RECT 233.400 65.800 234.500 66.100 ;
        RECT 236.500 66.000 236.900 66.100 ;
        RECT 237.400 66.100 237.800 67.400 ;
        RECT 239.700 67.700 240.500 68.000 ;
        RECT 239.700 67.500 240.100 67.700 ;
        RECT 239.700 67.200 240.000 67.500 ;
        RECT 242.300 67.400 242.600 68.500 ;
        RECT 238.200 67.100 238.600 67.200 ;
        RECT 239.000 67.100 240.000 67.200 ;
        RECT 238.200 66.800 240.000 67.100 ;
        RECT 240.500 67.100 242.600 67.400 ;
        RECT 243.000 68.500 243.400 69.500 ;
        RECT 243.000 67.400 243.300 68.500 ;
        RECT 245.100 68.200 245.500 69.500 ;
        RECT 244.600 68.000 245.500 68.200 ;
        RECT 247.800 68.500 248.200 69.500 ;
        RECT 244.600 67.800 245.900 68.000 ;
        RECT 245.100 67.700 245.900 67.800 ;
        RECT 245.500 67.500 245.900 67.700 ;
        RECT 243.000 67.100 245.100 67.400 ;
        RECT 240.500 66.900 241.000 67.100 ;
        RECT 239.000 66.100 239.400 66.200 ;
        RECT 237.400 65.800 239.400 66.100 ;
        RECT 227.000 65.400 227.400 65.800 ;
        RECT 228.600 65.500 231.400 65.600 ;
        RECT 228.600 65.400 231.500 65.500 ;
        RECT 225.900 64.600 226.700 64.900 ;
        RECT 228.600 65.300 233.500 65.400 ;
        RECT 223.800 61.500 224.200 63.500 ;
        RECT 225.900 61.100 226.300 64.600 ;
        RECT 228.600 61.100 229.000 65.300 ;
        RECT 231.100 65.100 233.500 65.300 ;
        RECT 230.200 64.500 232.900 64.800 ;
        RECT 230.200 64.400 230.600 64.500 ;
        RECT 232.500 64.400 232.900 64.500 ;
        RECT 233.200 64.500 233.500 65.100 ;
        RECT 234.200 65.200 234.500 65.800 ;
        RECT 235.700 65.700 236.100 65.800 ;
        RECT 237.400 65.700 237.800 65.800 ;
        RECT 235.700 65.400 237.800 65.700 ;
        RECT 239.000 65.400 239.400 65.800 ;
        RECT 234.200 64.900 235.400 65.200 ;
        RECT 233.900 64.500 234.300 64.600 ;
        RECT 233.200 64.200 234.300 64.500 ;
        RECT 235.100 64.400 235.400 64.900 ;
        RECT 235.100 64.000 235.800 64.400 ;
        RECT 231.900 63.700 232.300 63.800 ;
        RECT 233.300 63.700 233.700 63.800 ;
        RECT 230.200 63.100 230.600 63.500 ;
        RECT 231.900 63.400 233.700 63.700 ;
        RECT 233.000 63.100 233.300 63.400 ;
        RECT 235.000 63.100 235.400 63.500 ;
        RECT 230.200 62.800 231.200 63.100 ;
        RECT 230.800 61.100 231.200 62.800 ;
        RECT 233.000 61.100 233.400 63.100 ;
        RECT 235.100 61.100 235.700 63.100 ;
        RECT 237.400 61.100 237.800 65.400 ;
        RECT 239.700 64.900 240.000 66.800 ;
        RECT 240.300 66.500 241.000 66.900 ;
        RECT 244.600 66.900 245.100 67.100 ;
        RECT 245.600 67.200 245.900 67.500 ;
        RECT 247.800 67.400 248.100 68.500 ;
        RECT 249.900 68.000 250.300 69.500 ;
        RECT 249.900 67.700 250.700 68.000 ;
        RECT 252.600 67.900 253.000 69.900 ;
        RECT 253.400 68.000 253.800 69.900 ;
        RECT 255.000 68.000 255.400 69.900 ;
        RECT 253.400 67.900 255.400 68.000 ;
        RECT 250.300 67.500 250.700 67.700 ;
        RECT 240.700 65.500 241.000 66.500 ;
        RECT 241.400 65.800 241.800 66.600 ;
        RECT 242.200 65.800 242.600 66.600 ;
        RECT 243.000 65.800 243.400 66.600 ;
        RECT 243.800 65.800 244.200 66.600 ;
        RECT 244.600 66.500 245.300 66.900 ;
        RECT 245.600 66.800 246.600 67.200 ;
        RECT 247.800 67.100 249.900 67.400 ;
        RECT 249.400 66.900 249.900 67.100 ;
        RECT 250.400 67.200 250.700 67.500 ;
        RECT 252.700 67.200 253.000 67.900 ;
        RECT 253.500 67.700 255.300 67.900 ;
        RECT 255.800 67.700 256.200 69.900 ;
        RECT 257.900 69.200 258.500 69.900 ;
        RECT 257.900 68.900 258.600 69.200 ;
        RECT 260.200 68.900 260.600 69.900 ;
        RECT 262.400 69.200 262.800 69.900 ;
        RECT 262.400 68.900 263.400 69.200 ;
        RECT 258.200 68.500 258.600 68.900 ;
        RECT 260.300 68.600 260.600 68.900 ;
        RECT 260.300 68.300 261.700 68.600 ;
        RECT 261.300 68.200 261.700 68.300 ;
        RECT 262.200 68.200 262.600 68.600 ;
        RECT 263.000 68.500 263.400 68.900 ;
        RECT 257.300 67.700 257.700 67.800 ;
        RECT 255.800 67.400 257.700 67.700 ;
        RECT 254.600 67.200 255.000 67.400 ;
        RECT 244.600 65.500 244.900 66.500 ;
        RECT 240.700 65.200 242.600 65.500 ;
        RECT 239.700 64.600 240.500 64.900 ;
        RECT 240.100 61.100 240.500 64.600 ;
        RECT 242.300 63.500 242.600 65.200 ;
        RECT 242.200 61.500 242.600 63.500 ;
        RECT 243.000 65.200 244.900 65.500 ;
        RECT 243.000 63.500 243.300 65.200 ;
        RECT 245.600 64.900 245.900 66.800 ;
        RECT 246.200 65.400 246.600 66.200 ;
        RECT 247.800 65.800 248.200 66.600 ;
        RECT 248.600 65.800 249.000 66.600 ;
        RECT 249.400 66.500 250.100 66.900 ;
        RECT 250.400 66.800 251.400 67.200 ;
        RECT 252.600 66.800 253.900 67.200 ;
        RECT 254.600 66.900 255.400 67.200 ;
        RECT 255.000 66.800 255.400 66.900 ;
        RECT 249.400 65.500 249.700 66.500 ;
        RECT 245.100 64.600 245.900 64.900 ;
        RECT 247.800 65.200 249.700 65.500 ;
        RECT 250.400 65.200 250.700 66.800 ;
        RECT 251.000 65.400 251.400 66.200 ;
        RECT 253.600 65.200 253.900 66.800 ;
        RECT 254.200 65.800 254.600 66.600 ;
        RECT 255.800 65.700 256.200 67.400 ;
        RECT 262.200 67.200 262.500 68.200 ;
        RECT 264.600 67.500 265.000 69.900 ;
        RECT 259.300 67.100 259.700 67.200 ;
        RECT 262.200 67.100 262.600 67.200 ;
        RECT 263.800 67.100 264.600 67.200 ;
        RECT 259.100 66.800 264.600 67.100 ;
        RECT 258.200 66.400 258.600 66.500 ;
        RECT 256.700 66.100 258.600 66.400 ;
        RECT 256.700 66.000 257.100 66.100 ;
        RECT 257.500 65.700 257.900 65.800 ;
        RECT 255.800 65.400 257.900 65.700 ;
        RECT 243.000 61.500 243.400 63.500 ;
        RECT 245.100 61.100 245.500 64.600 ;
        RECT 247.800 63.500 248.100 65.200 ;
        RECT 250.200 64.900 250.700 65.200 ;
        RECT 249.900 64.600 250.700 64.900 ;
        RECT 252.600 65.100 253.000 65.200 ;
        RECT 252.600 64.800 253.300 65.100 ;
        RECT 253.600 64.800 254.600 65.200 ;
        RECT 247.800 61.500 248.200 63.500 ;
        RECT 249.900 61.100 250.300 64.600 ;
        RECT 253.000 64.200 253.300 64.800 ;
        RECT 253.000 63.800 253.400 64.200 ;
        RECT 253.700 61.100 254.100 64.800 ;
        RECT 255.800 61.100 256.200 65.400 ;
        RECT 259.100 65.200 259.400 66.800 ;
        RECT 262.700 66.700 263.100 66.800 ;
        RECT 263.500 66.200 263.900 66.300 ;
        RECT 260.600 66.100 261.000 66.200 ;
        RECT 261.400 66.100 263.900 66.200 ;
        RECT 260.600 65.900 263.900 66.100 ;
        RECT 260.600 65.800 261.800 65.900 ;
        RECT 262.200 65.500 265.000 65.600 ;
        RECT 262.100 65.400 265.000 65.500 ;
        RECT 258.200 64.900 259.400 65.200 ;
        RECT 260.100 65.300 265.000 65.400 ;
        RECT 260.100 65.100 262.500 65.300 ;
        RECT 258.200 64.400 258.500 64.900 ;
        RECT 257.800 64.000 258.500 64.400 ;
        RECT 259.300 64.500 259.700 64.600 ;
        RECT 260.100 64.500 260.400 65.100 ;
        RECT 259.300 64.200 260.400 64.500 ;
        RECT 260.700 64.500 263.400 64.800 ;
        RECT 260.700 64.400 261.100 64.500 ;
        RECT 263.000 64.400 263.400 64.500 ;
        RECT 259.900 63.700 260.300 63.800 ;
        RECT 261.300 63.700 261.700 63.800 ;
        RECT 258.200 63.100 258.600 63.500 ;
        RECT 259.900 63.400 261.700 63.700 ;
        RECT 260.300 63.100 260.600 63.400 ;
        RECT 263.000 63.100 263.400 63.500 ;
        RECT 257.900 61.100 258.500 63.100 ;
        RECT 260.200 61.100 260.600 63.100 ;
        RECT 262.400 62.800 263.400 63.100 ;
        RECT 262.400 61.100 262.800 62.800 ;
        RECT 264.600 61.100 265.000 65.300 ;
        RECT 1.400 55.600 1.800 59.900 ;
        RECT 3.000 55.600 3.400 59.900 ;
        RECT 4.600 55.600 5.000 59.900 ;
        RECT 6.200 55.600 6.600 59.900 ;
        RECT 8.600 55.600 9.000 59.900 ;
        RECT 10.200 55.600 10.600 59.900 ;
        RECT 11.800 55.600 12.200 59.900 ;
        RECT 13.400 55.600 13.800 59.900 ;
        RECT 15.000 57.500 15.400 59.500 ;
        RECT 17.100 59.200 17.500 59.900 ;
        RECT 17.100 58.800 17.800 59.200 ;
        RECT 15.000 55.800 15.300 57.500 ;
        RECT 17.100 56.400 17.500 58.800 ;
        RECT 17.100 56.100 17.900 56.400 ;
        RECT 1.400 55.200 2.300 55.600 ;
        RECT 3.000 55.200 4.100 55.600 ;
        RECT 4.600 55.200 5.700 55.600 ;
        RECT 6.200 55.200 7.400 55.600 ;
        RECT 8.600 55.200 9.500 55.600 ;
        RECT 10.200 55.200 11.300 55.600 ;
        RECT 11.800 55.200 12.900 55.600 ;
        RECT 13.400 55.200 14.600 55.600 ;
        RECT 15.000 55.500 16.900 55.800 ;
        RECT 1.900 54.500 2.300 55.200 ;
        RECT 3.700 54.500 4.100 55.200 ;
        RECT 5.300 54.500 5.700 55.200 ;
        RECT 0.600 54.100 1.500 54.500 ;
        RECT 1.900 54.100 3.200 54.500 ;
        RECT 3.700 54.100 4.900 54.500 ;
        RECT 5.300 54.100 6.600 54.500 ;
        RECT 0.600 53.800 1.000 54.100 ;
        RECT 1.900 53.800 2.300 54.100 ;
        RECT 3.700 53.800 4.100 54.100 ;
        RECT 5.300 53.800 5.700 54.100 ;
        RECT 7.000 53.800 7.400 55.200 ;
        RECT 9.100 54.500 9.500 55.200 ;
        RECT 10.900 54.500 11.300 55.200 ;
        RECT 12.500 54.500 12.900 55.200 ;
        RECT 7.800 54.100 8.700 54.500 ;
        RECT 9.100 54.100 10.400 54.500 ;
        RECT 10.900 54.100 12.100 54.500 ;
        RECT 12.500 54.100 13.800 54.500 ;
        RECT 7.800 53.800 8.200 54.100 ;
        RECT 9.100 53.800 9.500 54.100 ;
        RECT 10.900 53.800 11.300 54.100 ;
        RECT 12.500 53.800 12.900 54.100 ;
        RECT 14.200 53.800 14.600 55.200 ;
        RECT 15.000 54.400 15.400 55.200 ;
        RECT 15.800 54.400 16.200 55.200 ;
        RECT 16.600 54.500 16.900 55.500 ;
        RECT 16.600 54.100 17.300 54.500 ;
        RECT 17.600 54.200 17.900 56.100 ;
        RECT 19.800 55.700 20.200 59.900 ;
        RECT 22.000 58.200 22.400 59.900 ;
        RECT 21.400 57.900 22.400 58.200 ;
        RECT 24.200 57.900 24.600 59.900 ;
        RECT 26.300 57.900 26.900 59.900 ;
        RECT 21.400 57.500 21.800 57.900 ;
        RECT 24.200 57.600 24.500 57.900 ;
        RECT 23.100 57.300 24.900 57.600 ;
        RECT 26.200 57.500 26.600 57.900 ;
        RECT 23.100 57.200 23.500 57.300 ;
        RECT 24.500 57.200 24.900 57.300 ;
        RECT 21.400 56.500 21.800 56.600 ;
        RECT 23.700 56.500 24.100 56.600 ;
        RECT 21.400 56.200 24.100 56.500 ;
        RECT 24.400 56.500 25.500 56.800 ;
        RECT 24.400 55.900 24.700 56.500 ;
        RECT 25.100 56.400 25.500 56.500 ;
        RECT 26.300 56.600 27.000 57.000 ;
        RECT 26.300 56.100 26.600 56.600 ;
        RECT 22.300 55.700 24.700 55.900 ;
        RECT 19.800 55.600 24.700 55.700 ;
        RECT 25.400 55.800 26.600 56.100 ;
        RECT 18.200 54.800 18.600 55.600 ;
        RECT 19.800 55.500 22.700 55.600 ;
        RECT 19.800 55.400 22.600 55.500 ;
        RECT 23.000 55.100 23.400 55.200 ;
        RECT 20.900 54.800 23.400 55.100 ;
        RECT 20.900 54.700 21.300 54.800 ;
        RECT 21.700 54.200 22.100 54.300 ;
        RECT 25.400 54.200 25.700 55.800 ;
        RECT 28.600 55.600 29.000 59.900 ;
        RECT 26.900 55.300 29.000 55.600 ;
        RECT 29.400 57.500 29.800 59.500 ;
        RECT 29.400 55.800 29.700 57.500 ;
        RECT 31.500 56.400 31.900 59.900 ;
        RECT 31.500 56.100 32.300 56.400 ;
        RECT 29.400 55.500 31.300 55.800 ;
        RECT 26.900 55.200 27.300 55.300 ;
        RECT 27.700 54.900 28.100 55.000 ;
        RECT 26.200 54.600 28.100 54.900 ;
        RECT 26.200 54.500 26.600 54.600 ;
        RECT 16.600 53.900 17.100 54.100 ;
        RECT 1.400 53.400 2.300 53.800 ;
        RECT 3.000 53.400 4.100 53.800 ;
        RECT 4.600 53.400 5.700 53.800 ;
        RECT 6.200 53.400 7.400 53.800 ;
        RECT 8.600 53.400 9.500 53.800 ;
        RECT 10.200 53.400 11.300 53.800 ;
        RECT 11.800 53.400 12.900 53.800 ;
        RECT 13.400 53.400 14.600 53.800 ;
        RECT 15.000 53.600 17.100 53.900 ;
        RECT 17.600 53.800 18.600 54.200 ;
        RECT 20.200 53.900 25.700 54.200 ;
        RECT 20.200 53.800 21.000 53.900 ;
        RECT 1.400 51.100 1.800 53.400 ;
        RECT 3.000 51.100 3.400 53.400 ;
        RECT 4.600 51.100 5.000 53.400 ;
        RECT 6.200 51.100 6.600 53.400 ;
        RECT 8.600 51.100 9.000 53.400 ;
        RECT 10.200 51.100 10.600 53.400 ;
        RECT 11.800 51.100 12.200 53.400 ;
        RECT 13.400 51.100 13.800 53.400 ;
        RECT 15.000 52.500 15.300 53.600 ;
        RECT 17.600 53.500 17.900 53.800 ;
        RECT 17.500 53.300 17.900 53.500 ;
        RECT 17.100 53.000 17.900 53.300 ;
        RECT 15.000 51.500 15.400 52.500 ;
        RECT 17.100 51.500 17.500 53.000 ;
        RECT 19.800 51.100 20.200 53.500 ;
        RECT 22.300 52.800 22.600 53.900 ;
        RECT 25.100 53.800 25.500 53.900 ;
        RECT 28.600 53.600 29.000 55.300 ;
        RECT 29.400 54.400 29.800 55.200 ;
        RECT 30.200 54.400 30.600 55.200 ;
        RECT 31.000 54.500 31.300 55.500 ;
        RECT 31.000 54.100 31.700 54.500 ;
        RECT 32.000 54.200 32.300 56.100 ;
        RECT 32.600 55.100 33.000 55.600 ;
        RECT 34.200 55.100 34.600 59.900 ;
        RECT 32.600 54.800 34.600 55.100 ;
        RECT 31.000 53.900 31.500 54.100 ;
        RECT 27.100 53.300 29.000 53.600 ;
        RECT 27.100 53.200 27.500 53.300 ;
        RECT 21.400 52.100 21.800 52.500 ;
        RECT 22.200 52.400 22.600 52.800 ;
        RECT 23.100 52.700 23.500 52.800 ;
        RECT 23.100 52.400 24.500 52.700 ;
        RECT 24.200 52.100 24.500 52.400 ;
        RECT 26.200 52.100 26.600 52.500 ;
        RECT 21.400 51.800 22.400 52.100 ;
        RECT 22.000 51.100 22.400 51.800 ;
        RECT 24.200 51.100 24.600 52.100 ;
        RECT 26.200 51.800 26.900 52.100 ;
        RECT 26.300 51.100 26.900 51.800 ;
        RECT 28.600 51.100 29.000 53.300 ;
        RECT 29.400 53.600 31.500 53.900 ;
        RECT 32.000 53.800 33.000 54.200 ;
        RECT 29.400 52.500 29.700 53.600 ;
        RECT 32.000 53.500 32.300 53.800 ;
        RECT 31.900 53.300 32.300 53.500 ;
        RECT 31.500 53.200 32.300 53.300 ;
        RECT 31.000 53.000 32.300 53.200 ;
        RECT 31.000 52.800 31.900 53.000 ;
        RECT 29.400 51.500 29.800 52.500 ;
        RECT 31.500 51.500 31.900 52.800 ;
        RECT 34.200 51.100 34.600 54.800 ;
        RECT 36.600 55.100 37.000 59.900 ;
        RECT 39.300 56.400 39.700 59.900 ;
        RECT 41.400 57.500 41.800 59.500 ;
        RECT 38.900 56.100 39.700 56.400 ;
        RECT 38.200 55.100 38.600 55.600 ;
        RECT 36.600 54.800 38.600 55.100 ;
        RECT 35.000 52.400 35.400 53.200 ;
        RECT 35.800 52.400 36.200 53.200 ;
        RECT 36.600 51.100 37.000 54.800 ;
        RECT 38.900 54.200 39.200 56.100 ;
        RECT 41.500 55.800 41.800 57.500 ;
        RECT 39.900 55.500 41.800 55.800 ;
        RECT 42.200 57.500 42.600 59.500 ;
        RECT 44.300 59.200 44.700 59.900 ;
        RECT 44.300 58.800 45.000 59.200 ;
        RECT 42.200 55.800 42.500 57.500 ;
        RECT 44.300 56.400 44.700 58.800 ;
        RECT 44.300 56.100 45.100 56.400 ;
        RECT 42.200 55.500 44.100 55.800 ;
        RECT 39.900 54.500 40.200 55.500 ;
        RECT 38.200 53.800 39.200 54.200 ;
        RECT 39.500 54.100 40.200 54.500 ;
        RECT 40.600 54.400 41.000 55.200 ;
        RECT 41.400 54.400 41.800 55.200 ;
        RECT 42.200 54.400 42.600 55.200 ;
        RECT 43.000 54.400 43.400 55.200 ;
        RECT 43.800 54.500 44.100 55.500 ;
        RECT 38.900 53.500 39.200 53.800 ;
        RECT 39.700 53.900 40.200 54.100 ;
        RECT 43.800 54.100 44.500 54.500 ;
        RECT 44.800 54.200 45.100 56.100 ;
        RECT 47.000 55.700 47.400 59.900 ;
        RECT 49.200 58.200 49.600 59.900 ;
        RECT 48.600 57.900 49.600 58.200 ;
        RECT 51.400 57.900 51.800 59.900 ;
        RECT 53.500 57.900 54.100 59.900 ;
        RECT 48.600 57.500 49.000 57.900 ;
        RECT 51.400 57.600 51.700 57.900 ;
        RECT 50.300 57.300 52.100 57.600 ;
        RECT 53.400 57.500 53.800 57.900 ;
        RECT 50.300 57.200 50.700 57.300 ;
        RECT 51.700 57.200 52.100 57.300 ;
        RECT 48.600 56.500 49.000 56.600 ;
        RECT 50.900 56.500 51.300 56.600 ;
        RECT 48.600 56.200 51.300 56.500 ;
        RECT 51.600 56.500 52.700 56.800 ;
        RECT 51.600 55.900 51.900 56.500 ;
        RECT 52.300 56.400 52.700 56.500 ;
        RECT 53.500 56.600 54.200 57.000 ;
        RECT 53.500 56.100 53.800 56.600 ;
        RECT 49.500 55.700 51.900 55.900 ;
        RECT 47.000 55.600 51.900 55.700 ;
        RECT 52.600 55.800 53.800 56.100 ;
        RECT 45.400 55.100 45.800 55.600 ;
        RECT 47.000 55.500 49.900 55.600 ;
        RECT 47.000 55.400 49.800 55.500 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 50.200 55.100 50.600 55.200 ;
        RECT 51.000 55.100 51.400 55.200 ;
        RECT 45.400 54.800 46.600 55.100 ;
        RECT 48.100 54.800 51.400 55.100 ;
        RECT 48.100 54.700 48.500 54.800 ;
        RECT 48.900 54.200 49.300 54.300 ;
        RECT 52.600 54.200 52.900 55.800 ;
        RECT 55.800 55.600 56.200 59.900 ;
        RECT 58.200 56.200 58.600 59.900 ;
        RECT 59.800 56.200 60.200 59.900 ;
        RECT 58.200 55.900 60.200 56.200 ;
        RECT 54.100 55.300 56.200 55.600 ;
        RECT 60.600 55.800 61.000 59.900 ;
        RECT 62.700 56.300 63.100 59.900 ;
        RECT 65.700 59.200 66.100 59.900 ;
        RECT 65.700 58.800 66.600 59.200 ;
        RECT 65.700 56.400 66.100 58.800 ;
        RECT 67.800 57.500 68.200 59.500 ;
        RECT 62.200 55.900 63.100 56.300 ;
        RECT 65.300 56.100 66.100 56.400 ;
        RECT 54.100 55.200 54.500 55.300 ;
        RECT 54.900 54.900 55.300 55.000 ;
        RECT 53.400 54.600 55.300 54.900 ;
        RECT 53.400 54.500 53.800 54.600 ;
        RECT 43.800 53.900 44.300 54.100 ;
        RECT 39.700 53.600 41.800 53.900 ;
        RECT 38.900 53.300 39.300 53.500 ;
        RECT 38.900 53.000 39.700 53.300 ;
        RECT 39.300 51.500 39.700 53.000 ;
        RECT 41.500 52.500 41.800 53.600 ;
        RECT 41.400 51.500 41.800 52.500 ;
        RECT 42.200 53.600 44.300 53.900 ;
        RECT 44.800 53.800 45.800 54.200 ;
        RECT 47.400 53.900 52.900 54.200 ;
        RECT 47.400 53.800 48.200 53.900 ;
        RECT 42.200 52.500 42.500 53.600 ;
        RECT 44.800 53.500 45.100 53.800 ;
        RECT 44.700 53.300 45.100 53.500 ;
        RECT 44.300 53.000 45.100 53.300 ;
        RECT 42.200 51.500 42.600 52.500 ;
        RECT 44.300 51.500 44.700 53.000 ;
        RECT 47.000 51.100 47.400 53.500 ;
        RECT 49.500 52.800 49.800 53.900 ;
        RECT 50.200 53.800 50.600 53.900 ;
        RECT 52.300 53.800 52.700 53.900 ;
        RECT 55.800 53.600 56.200 55.300 ;
        RECT 58.600 55.200 59.000 55.400 ;
        RECT 60.600 55.200 60.900 55.800 ;
        RECT 57.400 55.100 57.800 55.200 ;
        RECT 58.200 55.100 59.000 55.200 ;
        RECT 57.400 54.900 59.000 55.100 ;
        RECT 59.800 54.900 61.000 55.200 ;
        RECT 57.400 54.800 58.600 54.900 ;
        RECT 59.000 53.800 59.400 54.600 ;
        RECT 54.300 53.300 56.200 53.600 ;
        RECT 54.300 53.200 54.700 53.300 ;
        RECT 48.600 52.100 49.000 52.500 ;
        RECT 49.400 52.400 49.800 52.800 ;
        RECT 50.300 52.700 50.700 52.800 ;
        RECT 50.300 52.400 51.700 52.700 ;
        RECT 51.400 52.100 51.700 52.400 ;
        RECT 53.400 52.100 53.800 52.500 ;
        RECT 48.600 51.800 49.600 52.100 ;
        RECT 49.200 51.100 49.600 51.800 ;
        RECT 51.400 51.100 51.800 52.100 ;
        RECT 53.400 51.800 54.100 52.100 ;
        RECT 53.500 51.100 54.100 51.800 ;
        RECT 55.800 51.100 56.200 53.300 ;
        RECT 59.800 53.100 60.100 54.900 ;
        RECT 60.600 54.800 61.000 54.900 ;
        RECT 62.300 54.200 62.600 55.900 ;
        RECT 63.000 54.800 63.400 55.600 ;
        RECT 63.800 55.100 64.200 55.200 ;
        RECT 64.600 55.100 65.000 55.600 ;
        RECT 63.800 54.800 65.000 55.100 ;
        RECT 65.300 54.200 65.600 56.100 ;
        RECT 67.900 55.800 68.200 57.500 ;
        RECT 69.900 56.200 70.300 59.900 ;
        RECT 70.600 56.800 71.000 57.200 ;
        RECT 70.700 56.200 71.000 56.800 ;
        RECT 69.900 55.900 70.400 56.200 ;
        RECT 70.700 56.100 71.400 56.200 ;
        RECT 72.600 56.100 73.000 59.900 ;
        RECT 70.700 55.900 73.000 56.100 ;
        RECT 66.300 55.500 68.200 55.800 ;
        RECT 66.300 54.500 66.600 55.500 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 60.600 53.800 62.600 54.100 ;
        RECT 64.600 53.800 65.600 54.200 ;
        RECT 65.900 54.100 66.600 54.500 ;
        RECT 67.000 54.400 67.400 55.200 ;
        RECT 67.800 54.400 68.200 55.200 ;
        RECT 69.400 54.400 69.800 55.200 ;
        RECT 70.100 54.200 70.400 55.900 ;
        RECT 71.000 55.800 73.000 55.900 ;
        RECT 73.400 55.800 73.800 56.600 ;
        RECT 71.800 54.800 72.200 55.200 ;
        RECT 71.800 54.200 72.100 54.800 ;
        RECT 60.600 53.200 60.900 53.800 ;
        RECT 59.800 51.100 60.200 53.100 ;
        RECT 60.600 52.800 61.000 53.200 ;
        RECT 60.500 52.400 60.900 52.800 ;
        RECT 61.400 52.400 61.800 53.200 ;
        RECT 62.300 52.100 62.600 53.800 ;
        RECT 65.300 53.500 65.600 53.800 ;
        RECT 66.100 53.900 66.600 54.100 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 66.100 53.600 68.200 53.900 ;
        RECT 68.600 53.800 69.400 54.100 ;
        RECT 70.100 53.800 71.400 54.200 ;
        RECT 69.000 53.600 69.400 53.800 ;
        RECT 65.300 53.300 65.700 53.500 ;
        RECT 65.300 53.000 66.100 53.300 ;
        RECT 62.200 51.100 62.600 52.100 ;
        RECT 65.700 51.500 66.100 53.000 ;
        RECT 67.900 52.500 68.200 53.600 ;
        RECT 68.700 53.100 70.500 53.300 ;
        RECT 71.000 53.100 71.300 53.800 ;
        RECT 71.800 53.400 72.200 54.200 ;
        RECT 72.600 53.100 73.000 55.800 ;
        RECT 74.200 55.600 74.600 59.900 ;
        RECT 76.300 57.900 76.900 59.900 ;
        RECT 78.600 57.900 79.000 59.900 ;
        RECT 80.800 58.200 81.200 59.900 ;
        RECT 80.800 57.900 81.800 58.200 ;
        RECT 76.600 57.500 77.000 57.900 ;
        RECT 78.700 57.600 79.000 57.900 ;
        RECT 78.300 57.300 80.100 57.600 ;
        RECT 81.400 57.500 81.800 57.900 ;
        RECT 78.300 57.200 78.700 57.300 ;
        RECT 79.700 57.200 80.100 57.300 ;
        RECT 76.200 56.600 76.900 57.000 ;
        RECT 76.600 56.100 76.900 56.600 ;
        RECT 77.700 56.500 78.800 56.800 ;
        RECT 77.700 56.400 78.100 56.500 ;
        RECT 76.600 55.800 77.800 56.100 ;
        RECT 74.200 55.300 76.300 55.600 ;
        RECT 74.200 53.600 74.600 55.300 ;
        RECT 75.900 55.200 76.300 55.300 ;
        RECT 75.100 54.900 75.500 55.000 ;
        RECT 75.100 54.600 77.000 54.900 ;
        RECT 76.600 54.500 77.000 54.600 ;
        RECT 77.500 54.200 77.800 55.800 ;
        RECT 78.500 55.900 78.800 56.500 ;
        RECT 79.100 56.500 79.500 56.600 ;
        RECT 81.400 56.500 81.800 56.600 ;
        RECT 79.100 56.200 81.800 56.500 ;
        RECT 78.500 55.700 80.900 55.900 ;
        RECT 83.000 55.700 83.400 59.900 ;
        RECT 85.100 56.200 85.500 59.900 ;
        RECT 85.800 56.800 86.200 57.200 ;
        RECT 85.900 56.200 86.200 56.800 ;
        RECT 85.100 55.900 85.600 56.200 ;
        RECT 85.900 56.100 86.600 56.200 ;
        RECT 87.800 56.100 88.200 59.900 ;
        RECT 89.400 57.500 89.800 59.500 ;
        RECT 91.500 59.200 91.900 59.900 ;
        RECT 91.500 58.800 92.200 59.200 ;
        RECT 85.900 55.900 88.200 56.100 ;
        RECT 78.500 55.600 83.400 55.700 ;
        RECT 80.500 55.500 83.400 55.600 ;
        RECT 80.600 55.400 83.400 55.500 ;
        RECT 85.300 55.200 85.600 55.900 ;
        RECT 86.200 55.800 88.200 55.900 ;
        RECT 88.600 55.800 89.000 56.600 ;
        RECT 89.400 55.800 89.700 57.500 ;
        RECT 91.500 56.400 91.900 58.800 ;
        RECT 94.200 57.500 94.600 59.500 ;
        RECT 96.300 59.200 96.700 59.900 ;
        RECT 96.300 58.800 97.000 59.200 ;
        RECT 91.500 56.100 92.300 56.400 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 83.800 55.100 84.200 55.200 ;
        RECT 84.600 55.100 85.000 55.200 ;
        RECT 79.800 54.800 82.300 55.100 ;
        RECT 83.800 54.800 85.000 55.100 ;
        RECT 80.600 54.700 81.000 54.800 ;
        RECT 81.900 54.700 82.300 54.800 ;
        RECT 84.600 54.400 85.000 54.800 ;
        RECT 85.300 54.800 85.800 55.200 ;
        RECT 81.100 54.200 81.500 54.300 ;
        RECT 85.300 54.200 85.600 54.800 ;
        RECT 77.500 53.900 83.000 54.200 ;
        RECT 77.700 53.800 78.100 53.900 ;
        RECT 79.800 53.800 80.200 53.900 ;
        RECT 74.200 53.300 76.100 53.600 ;
        RECT 67.800 51.500 68.200 52.500 ;
        RECT 68.600 53.000 70.600 53.100 ;
        RECT 68.600 51.100 69.000 53.000 ;
        RECT 70.200 51.100 70.600 53.000 ;
        RECT 71.000 51.100 71.400 53.100 ;
        RECT 72.600 52.800 73.500 53.100 ;
        RECT 73.100 51.100 73.500 52.800 ;
        RECT 74.200 51.100 74.600 53.300 ;
        RECT 75.700 53.200 76.100 53.300 ;
        RECT 80.600 52.800 80.900 53.900 ;
        RECT 82.200 53.800 83.000 53.900 ;
        RECT 83.800 54.100 84.200 54.200 ;
        RECT 83.800 53.800 84.600 54.100 ;
        RECT 85.300 53.800 86.600 54.200 ;
        RECT 84.200 53.600 84.600 53.800 ;
        RECT 79.700 52.700 80.100 52.800 ;
        RECT 76.600 52.100 77.000 52.500 ;
        RECT 78.700 52.400 80.100 52.700 ;
        RECT 80.600 52.400 81.000 52.800 ;
        RECT 78.700 52.100 79.000 52.400 ;
        RECT 81.400 52.100 81.800 52.500 ;
        RECT 76.300 51.800 77.000 52.100 ;
        RECT 76.300 51.100 76.900 51.800 ;
        RECT 78.600 51.100 79.000 52.100 ;
        RECT 80.800 51.800 81.800 52.100 ;
        RECT 80.800 51.100 81.200 51.800 ;
        RECT 83.000 51.100 83.400 53.500 ;
        RECT 83.900 53.100 85.700 53.300 ;
        RECT 86.200 53.100 86.500 53.800 ;
        RECT 87.000 53.400 87.400 54.200 ;
        RECT 87.800 53.100 88.200 55.800 ;
        RECT 89.400 55.500 91.300 55.800 ;
        RECT 89.400 54.400 89.800 55.200 ;
        RECT 90.200 54.400 90.600 55.200 ;
        RECT 91.000 54.500 91.300 55.500 ;
        RECT 91.000 54.100 91.700 54.500 ;
        RECT 92.000 54.200 92.300 56.100 ;
        RECT 94.200 55.800 94.500 57.500 ;
        RECT 96.300 56.400 96.700 58.800 ;
        RECT 96.300 56.100 97.100 56.400 ;
        RECT 92.600 54.800 93.000 55.600 ;
        RECT 94.200 55.500 96.100 55.800 ;
        RECT 94.200 54.400 94.600 55.200 ;
        RECT 95.000 54.400 95.400 55.200 ;
        RECT 95.800 54.500 96.100 55.500 ;
        RECT 91.000 53.900 91.500 54.100 ;
        RECT 89.400 53.600 91.500 53.900 ;
        RECT 92.000 53.800 93.000 54.200 ;
        RECT 95.800 54.100 96.500 54.500 ;
        RECT 96.800 54.200 97.100 56.100 ;
        RECT 99.000 55.700 99.400 59.900 ;
        RECT 101.200 58.200 101.600 59.900 ;
        RECT 100.600 57.900 101.600 58.200 ;
        RECT 103.400 57.900 103.800 59.900 ;
        RECT 105.500 57.900 106.100 59.900 ;
        RECT 100.600 57.500 101.000 57.900 ;
        RECT 103.400 57.600 103.700 57.900 ;
        RECT 102.300 57.300 104.100 57.600 ;
        RECT 105.400 57.500 105.800 57.900 ;
        RECT 102.300 57.200 102.700 57.300 ;
        RECT 103.700 57.200 104.100 57.300 ;
        RECT 100.600 56.500 101.000 56.600 ;
        RECT 102.900 56.500 103.300 56.600 ;
        RECT 100.600 56.200 103.300 56.500 ;
        RECT 103.600 56.500 104.700 56.800 ;
        RECT 103.600 55.900 103.900 56.500 ;
        RECT 104.300 56.400 104.700 56.500 ;
        RECT 105.500 56.600 106.200 57.000 ;
        RECT 105.500 56.100 105.800 56.600 ;
        RECT 101.500 55.700 103.900 55.900 ;
        RECT 99.000 55.600 103.900 55.700 ;
        RECT 104.600 55.800 105.800 56.100 ;
        RECT 97.400 55.100 97.800 55.600 ;
        RECT 99.000 55.500 101.900 55.600 ;
        RECT 99.000 55.400 101.800 55.500 ;
        RECT 98.200 55.100 98.600 55.200 ;
        RECT 102.200 55.100 102.600 55.200 ;
        RECT 97.400 54.800 98.600 55.100 ;
        RECT 100.100 54.800 102.600 55.100 ;
        RECT 100.100 54.700 100.500 54.800 ;
        RECT 100.900 54.200 101.300 54.300 ;
        RECT 104.600 54.200 104.900 55.800 ;
        RECT 107.800 55.600 108.200 59.900 ;
        RECT 110.600 56.800 111.000 57.200 ;
        RECT 110.600 56.200 110.900 56.800 ;
        RECT 111.300 56.200 111.700 59.900 ;
        RECT 114.700 56.300 115.100 59.900 ;
        RECT 110.200 55.900 110.900 56.200 ;
        RECT 111.200 55.900 111.700 56.200 ;
        RECT 114.200 55.900 115.100 56.300 ;
        RECT 115.800 55.900 116.200 59.900 ;
        RECT 116.600 56.200 117.000 59.900 ;
        RECT 118.200 56.200 118.600 59.900 ;
        RECT 116.600 55.900 118.600 56.200 ;
        RECT 110.200 55.800 110.600 55.900 ;
        RECT 106.100 55.300 108.200 55.600 ;
        RECT 106.100 55.200 106.500 55.300 ;
        RECT 106.900 54.900 107.300 55.000 ;
        RECT 105.400 54.600 107.300 54.900 ;
        RECT 105.400 54.500 105.800 54.600 ;
        RECT 95.800 53.900 96.300 54.100 ;
        RECT 83.800 53.000 85.800 53.100 ;
        RECT 83.800 51.100 84.200 53.000 ;
        RECT 85.400 51.100 85.800 53.000 ;
        RECT 86.200 51.100 86.600 53.100 ;
        RECT 87.800 52.800 88.700 53.100 ;
        RECT 88.300 51.100 88.700 52.800 ;
        RECT 89.400 52.500 89.700 53.600 ;
        RECT 92.000 53.500 92.300 53.800 ;
        RECT 91.900 53.300 92.300 53.500 ;
        RECT 91.500 53.000 92.300 53.300 ;
        RECT 94.200 53.600 96.300 53.900 ;
        RECT 96.800 53.800 97.800 54.200 ;
        RECT 99.400 53.900 105.000 54.200 ;
        RECT 99.400 53.800 100.200 53.900 ;
        RECT 101.400 53.800 101.800 53.900 ;
        RECT 104.300 53.800 105.000 53.900 ;
        RECT 89.400 51.500 89.800 52.500 ;
        RECT 91.500 51.500 91.900 53.000 ;
        RECT 94.200 52.500 94.500 53.600 ;
        RECT 96.800 53.500 97.100 53.800 ;
        RECT 96.700 53.300 97.100 53.500 ;
        RECT 96.300 53.000 97.100 53.300 ;
        RECT 94.200 51.500 94.600 52.500 ;
        RECT 96.300 51.500 96.700 53.000 ;
        RECT 99.000 51.100 99.400 53.500 ;
        RECT 101.500 52.800 101.800 53.800 ;
        RECT 107.800 53.600 108.200 55.300 ;
        RECT 109.400 55.100 109.800 55.200 ;
        RECT 111.200 55.100 111.500 55.900 ;
        RECT 109.400 54.800 111.500 55.100 ;
        RECT 111.200 54.200 111.500 54.800 ;
        RECT 111.800 54.400 112.200 55.200 ;
        RECT 114.300 54.200 114.600 55.900 ;
        RECT 115.000 54.800 115.400 55.600 ;
        RECT 115.900 55.200 116.200 55.900 ;
        RECT 119.000 55.700 119.400 59.900 ;
        RECT 121.200 58.200 121.600 59.900 ;
        RECT 120.600 57.900 121.600 58.200 ;
        RECT 123.400 57.900 123.800 59.900 ;
        RECT 125.500 57.900 126.100 59.900 ;
        RECT 120.600 57.500 121.000 57.900 ;
        RECT 123.400 57.600 123.700 57.900 ;
        RECT 122.300 57.300 124.100 57.600 ;
        RECT 125.400 57.500 125.800 57.900 ;
        RECT 122.300 57.200 122.700 57.300 ;
        RECT 123.700 57.200 124.100 57.300 ;
        RECT 120.600 56.500 121.000 56.600 ;
        RECT 122.900 56.500 123.300 56.600 ;
        RECT 120.600 56.200 123.300 56.500 ;
        RECT 123.600 56.500 124.700 56.800 ;
        RECT 123.600 55.900 123.900 56.500 ;
        RECT 124.300 56.400 124.700 56.500 ;
        RECT 125.500 56.600 126.200 57.000 ;
        RECT 125.500 56.100 125.800 56.600 ;
        RECT 121.500 55.700 123.900 55.900 ;
        RECT 119.000 55.600 123.900 55.700 ;
        RECT 124.600 55.800 125.800 56.100 ;
        RECT 119.000 55.500 121.900 55.600 ;
        RECT 119.000 55.400 121.800 55.500 ;
        RECT 117.800 55.200 118.200 55.400 ;
        RECT 115.800 54.900 117.000 55.200 ;
        RECT 117.800 54.900 118.600 55.200 ;
        RECT 122.200 55.100 122.600 55.200 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 115.800 54.800 116.200 54.900 ;
        RECT 110.200 53.800 111.500 54.200 ;
        RECT 112.600 54.100 113.000 54.200 ;
        RECT 113.400 54.100 113.800 54.200 ;
        RECT 112.200 53.800 113.800 54.100 ;
        RECT 114.200 53.800 114.600 54.200 ;
        RECT 106.300 53.300 108.200 53.600 ;
        RECT 106.300 53.200 106.700 53.300 ;
        RECT 100.600 52.100 101.000 52.500 ;
        RECT 101.400 52.400 101.800 52.800 ;
        RECT 102.300 52.700 102.700 52.800 ;
        RECT 102.300 52.400 103.700 52.700 ;
        RECT 103.400 52.100 103.700 52.400 ;
        RECT 105.400 52.100 105.800 52.500 ;
        RECT 100.600 51.800 101.600 52.100 ;
        RECT 101.200 51.100 101.600 51.800 ;
        RECT 103.400 51.100 103.800 52.100 ;
        RECT 105.400 51.800 106.100 52.100 ;
        RECT 105.500 51.100 106.100 51.800 ;
        RECT 107.800 51.100 108.200 53.300 ;
        RECT 110.300 53.100 110.600 53.800 ;
        RECT 112.200 53.600 112.600 53.800 ;
        RECT 111.100 53.100 112.900 53.300 ;
        RECT 110.200 51.100 110.600 53.100 ;
        RECT 111.000 53.000 113.000 53.100 ;
        RECT 111.000 51.100 111.400 53.000 ;
        RECT 112.600 51.100 113.000 53.000 ;
        RECT 113.400 52.400 113.800 53.200 ;
        RECT 114.300 53.100 114.600 53.800 ;
        RECT 115.800 53.100 116.200 53.200 ;
        RECT 116.700 53.100 117.000 54.900 ;
        RECT 118.200 54.800 118.600 54.900 ;
        RECT 120.100 54.800 123.400 55.100 ;
        RECT 120.100 54.700 120.500 54.800 ;
        RECT 117.400 53.800 117.800 54.600 ;
        RECT 120.900 54.200 121.300 54.300 ;
        RECT 124.600 54.200 124.900 55.800 ;
        RECT 127.800 55.600 128.200 59.900 ;
        RECT 126.100 55.300 128.200 55.600 ;
        RECT 126.100 55.200 126.500 55.300 ;
        RECT 126.900 54.900 127.300 55.000 ;
        RECT 125.400 54.600 127.300 54.900 ;
        RECT 125.400 54.500 125.800 54.600 ;
        RECT 119.400 53.900 124.900 54.200 ;
        RECT 127.800 54.100 128.200 55.300 ;
        RECT 129.400 55.100 129.800 59.900 ;
        RECT 131.400 56.800 131.800 57.200 ;
        RECT 130.200 55.800 130.600 56.600 ;
        RECT 131.400 56.200 131.700 56.800 ;
        RECT 132.100 56.200 132.500 59.900 ;
        RECT 136.100 59.200 136.500 59.900 ;
        RECT 136.100 58.800 137.000 59.200 ;
        RECT 136.100 56.400 136.500 58.800 ;
        RECT 138.200 57.500 138.600 59.500 ;
        RECT 131.000 55.900 131.700 56.200 ;
        RECT 132.000 55.900 132.500 56.200 ;
        RECT 135.700 56.100 136.500 56.400 ;
        RECT 131.000 55.800 131.400 55.900 ;
        RECT 131.000 55.100 131.300 55.800 ;
        RECT 132.000 55.200 132.300 55.900 ;
        RECT 129.400 54.800 131.300 55.100 ;
        RECT 131.800 54.800 132.300 55.200 ;
        RECT 128.600 54.100 129.000 54.200 ;
        RECT 119.400 53.800 120.200 53.900 ;
        RECT 114.200 52.800 116.200 53.100 ;
        RECT 114.300 52.100 114.600 52.800 ;
        RECT 115.900 52.400 116.300 52.800 ;
        RECT 114.200 51.100 114.600 52.100 ;
        RECT 116.600 51.100 117.000 53.100 ;
        RECT 119.000 51.100 119.400 53.500 ;
        RECT 121.500 52.800 121.800 53.900 ;
        RECT 124.300 53.800 124.700 53.900 ;
        RECT 127.800 53.800 129.000 54.100 ;
        RECT 127.800 53.600 128.200 53.800 ;
        RECT 126.300 53.300 128.200 53.600 ;
        RECT 128.600 53.400 129.000 53.800 ;
        RECT 126.300 53.200 126.700 53.300 ;
        RECT 120.600 52.100 121.000 52.500 ;
        RECT 121.400 52.400 121.800 52.800 ;
        RECT 122.300 52.700 122.700 52.800 ;
        RECT 122.300 52.400 123.700 52.700 ;
        RECT 123.400 52.100 123.700 52.400 ;
        RECT 125.400 52.100 125.800 52.500 ;
        RECT 120.600 51.800 121.600 52.100 ;
        RECT 121.200 51.100 121.600 51.800 ;
        RECT 123.400 51.100 123.800 52.100 ;
        RECT 125.400 51.800 126.100 52.100 ;
        RECT 125.500 51.100 126.100 51.800 ;
        RECT 127.800 51.100 128.200 53.300 ;
        RECT 129.400 53.100 129.800 54.800 ;
        RECT 132.000 54.200 132.300 54.800 ;
        RECT 132.600 54.400 133.000 55.200 ;
        RECT 135.000 54.800 135.400 55.600 ;
        RECT 135.700 54.200 136.000 56.100 ;
        RECT 138.300 55.800 138.600 57.500 ;
        RECT 136.700 55.500 138.600 55.800 ;
        RECT 139.000 57.500 139.400 59.500 ;
        RECT 141.100 59.200 141.500 59.900 ;
        RECT 141.100 58.800 141.800 59.200 ;
        RECT 139.000 55.800 139.300 57.500 ;
        RECT 141.100 56.400 141.500 58.800 ;
        RECT 143.800 57.500 144.200 59.500 ;
        RECT 145.900 59.200 146.300 59.900 ;
        RECT 145.400 58.800 146.300 59.200 ;
        RECT 141.100 56.100 141.900 56.400 ;
        RECT 139.000 55.500 140.900 55.800 ;
        RECT 136.700 54.500 137.000 55.500 ;
        RECT 131.000 53.800 132.300 54.200 ;
        RECT 133.400 54.100 133.800 54.200 ;
        RECT 133.000 53.800 133.800 54.100 ;
        RECT 135.000 53.800 136.000 54.200 ;
        RECT 136.300 54.100 137.000 54.500 ;
        RECT 137.400 54.400 137.800 55.200 ;
        RECT 138.200 54.400 138.600 55.200 ;
        RECT 139.000 54.400 139.400 55.200 ;
        RECT 139.800 54.400 140.200 55.200 ;
        RECT 140.600 54.500 140.900 55.500 ;
        RECT 131.100 53.100 131.400 53.800 ;
        RECT 133.000 53.600 133.400 53.800 ;
        RECT 135.700 53.500 136.000 53.800 ;
        RECT 136.500 53.900 137.000 54.100 ;
        RECT 140.600 54.100 141.300 54.500 ;
        RECT 141.600 54.200 141.900 56.100 ;
        RECT 143.800 55.800 144.100 57.500 ;
        RECT 145.900 56.400 146.300 58.800 ;
        RECT 145.900 56.100 146.700 56.400 ;
        RECT 142.200 54.800 142.600 55.600 ;
        RECT 143.800 55.500 145.700 55.800 ;
        RECT 143.000 55.100 143.400 55.200 ;
        RECT 143.800 55.100 144.200 55.200 ;
        RECT 143.000 54.800 144.200 55.100 ;
        RECT 143.800 54.400 144.200 54.800 ;
        RECT 144.600 54.400 145.000 55.200 ;
        RECT 145.400 54.500 145.700 55.500 ;
        RECT 140.600 53.900 141.100 54.100 ;
        RECT 136.500 53.600 138.600 53.900 ;
        RECT 135.700 53.300 136.100 53.500 ;
        RECT 131.900 53.100 133.700 53.300 ;
        RECT 129.400 52.800 130.300 53.100 ;
        RECT 129.900 51.100 130.300 52.800 ;
        RECT 131.000 51.100 131.400 53.100 ;
        RECT 131.800 53.000 133.800 53.100 ;
        RECT 135.700 53.000 136.500 53.300 ;
        RECT 131.800 51.100 132.200 53.000 ;
        RECT 133.400 51.100 133.800 53.000 ;
        RECT 136.100 51.500 136.500 53.000 ;
        RECT 138.300 52.500 138.600 53.600 ;
        RECT 138.200 51.500 138.600 52.500 ;
        RECT 139.000 53.600 141.100 53.900 ;
        RECT 141.600 53.800 142.600 54.200 ;
        RECT 145.400 54.100 146.100 54.500 ;
        RECT 146.400 54.200 146.700 56.100 ;
        RECT 148.600 55.700 149.000 59.900 ;
        RECT 150.800 58.200 151.200 59.900 ;
        RECT 150.200 57.900 151.200 58.200 ;
        RECT 153.000 57.900 153.400 59.900 ;
        RECT 155.100 57.900 155.700 59.900 ;
        RECT 150.200 57.500 150.600 57.900 ;
        RECT 153.000 57.600 153.300 57.900 ;
        RECT 151.900 57.300 153.700 57.600 ;
        RECT 155.000 57.500 155.400 57.900 ;
        RECT 151.900 57.200 152.300 57.300 ;
        RECT 153.300 57.200 153.700 57.300 ;
        RECT 150.200 56.500 150.600 56.600 ;
        RECT 152.500 56.500 152.900 56.600 ;
        RECT 150.200 56.200 152.900 56.500 ;
        RECT 153.200 56.500 154.300 56.800 ;
        RECT 153.200 55.900 153.500 56.500 ;
        RECT 153.900 56.400 154.300 56.500 ;
        RECT 155.100 56.600 155.800 57.000 ;
        RECT 155.100 56.100 155.400 56.600 ;
        RECT 151.100 55.700 153.500 55.900 ;
        RECT 148.600 55.600 153.500 55.700 ;
        RECT 154.200 55.800 155.400 56.100 ;
        RECT 147.000 54.800 147.400 55.600 ;
        RECT 148.600 55.500 151.500 55.600 ;
        RECT 148.600 55.400 151.400 55.500 ;
        RECT 151.800 55.100 152.200 55.200 ;
        RECT 149.700 54.800 152.200 55.100 ;
        RECT 149.700 54.700 150.100 54.800 ;
        RECT 150.500 54.200 150.900 54.300 ;
        RECT 154.200 54.200 154.500 55.800 ;
        RECT 157.400 55.600 157.800 59.900 ;
        RECT 161.100 56.200 161.500 59.900 ;
        RECT 161.800 56.800 162.200 57.200 ;
        RECT 161.900 56.200 162.200 56.800 ;
        RECT 161.100 55.900 161.600 56.200 ;
        RECT 161.900 55.900 162.600 56.200 ;
        RECT 155.700 55.300 157.800 55.600 ;
        RECT 155.700 55.200 156.100 55.300 ;
        RECT 156.500 54.900 156.900 55.000 ;
        RECT 155.000 54.600 156.900 54.900 ;
        RECT 155.000 54.500 155.400 54.600 ;
        RECT 145.400 53.900 145.900 54.100 ;
        RECT 139.000 52.500 139.300 53.600 ;
        RECT 141.600 53.500 141.900 53.800 ;
        RECT 141.500 53.300 141.900 53.500 ;
        RECT 141.100 53.000 141.900 53.300 ;
        RECT 143.800 53.600 145.900 53.900 ;
        RECT 146.400 53.800 147.400 54.200 ;
        RECT 149.000 53.900 154.500 54.200 ;
        RECT 149.000 53.800 149.800 53.900 ;
        RECT 139.000 51.500 139.400 52.500 ;
        RECT 141.100 51.500 141.500 53.000 ;
        RECT 143.800 52.500 144.100 53.600 ;
        RECT 146.400 53.500 146.700 53.800 ;
        RECT 146.300 53.300 146.700 53.500 ;
        RECT 145.900 53.000 146.700 53.300 ;
        RECT 143.800 51.500 144.200 52.500 ;
        RECT 145.900 51.500 146.300 53.000 ;
        RECT 148.600 51.100 149.000 53.500 ;
        RECT 151.100 52.800 151.400 53.900 ;
        RECT 153.900 53.800 154.300 53.900 ;
        RECT 157.400 53.600 157.800 55.300 ;
        RECT 161.300 55.200 161.600 55.900 ;
        RECT 162.200 55.800 162.600 55.900 ;
        RECT 163.000 55.800 163.400 56.600 ;
        RECT 160.600 54.400 161.000 55.200 ;
        RECT 161.300 54.800 161.800 55.200 ;
        RECT 162.200 55.100 162.500 55.800 ;
        RECT 163.800 55.100 164.200 59.900 ;
        RECT 167.300 59.200 167.700 59.900 ;
        RECT 167.000 58.800 167.700 59.200 ;
        RECT 167.300 56.400 167.700 58.800 ;
        RECT 169.400 57.500 169.800 59.500 ;
        RECT 172.100 59.200 172.500 59.900 ;
        RECT 171.800 58.800 172.500 59.200 ;
        RECT 166.900 56.100 167.700 56.400 ;
        RECT 166.200 55.100 166.600 55.600 ;
        RECT 162.200 54.800 164.200 55.100 ;
        RECT 161.300 54.200 161.600 54.800 ;
        RECT 159.800 54.100 160.200 54.200 ;
        RECT 159.800 53.800 160.600 54.100 ;
        RECT 161.300 53.800 162.600 54.200 ;
        RECT 160.200 53.600 160.600 53.800 ;
        RECT 155.900 53.300 157.800 53.600 ;
        RECT 155.900 53.200 156.300 53.300 ;
        RECT 150.200 52.100 150.600 52.500 ;
        RECT 151.000 52.400 151.400 52.800 ;
        RECT 151.900 52.700 152.300 52.800 ;
        RECT 151.900 52.400 153.300 52.700 ;
        RECT 153.000 52.100 153.300 52.400 ;
        RECT 155.000 52.100 155.400 52.500 ;
        RECT 150.200 51.800 151.200 52.100 ;
        RECT 150.800 51.100 151.200 51.800 ;
        RECT 153.000 51.100 153.400 52.100 ;
        RECT 155.000 51.800 155.700 52.100 ;
        RECT 155.100 51.100 155.700 51.800 ;
        RECT 157.400 51.100 157.800 53.300 ;
        RECT 159.900 53.100 161.700 53.300 ;
        RECT 162.200 53.100 162.500 53.800 ;
        RECT 163.800 53.100 164.200 54.800 ;
        RECT 165.400 54.800 166.600 55.100 ;
        RECT 164.600 54.100 165.000 54.200 ;
        RECT 165.400 54.100 165.700 54.800 ;
        RECT 166.900 54.200 167.200 56.100 ;
        RECT 169.500 55.800 169.800 57.500 ;
        RECT 172.100 56.400 172.500 58.800 ;
        RECT 174.200 57.500 174.600 59.500 ;
        RECT 167.900 55.500 169.800 55.800 ;
        RECT 171.700 56.100 172.500 56.400 ;
        RECT 167.900 54.500 168.200 55.500 ;
        RECT 164.600 53.800 165.700 54.100 ;
        RECT 166.200 53.800 167.200 54.200 ;
        RECT 167.500 54.100 168.200 54.500 ;
        RECT 168.600 54.400 169.000 55.200 ;
        RECT 169.400 54.400 169.800 55.200 ;
        RECT 170.200 55.100 170.600 55.200 ;
        RECT 171.000 55.100 171.400 55.600 ;
        RECT 170.200 54.800 171.400 55.100 ;
        RECT 171.700 54.200 172.000 56.100 ;
        RECT 174.300 55.800 174.600 57.500 ;
        RECT 176.300 56.300 176.700 59.900 ;
        RECT 175.800 55.900 176.700 56.300 ;
        RECT 177.400 55.900 177.800 59.900 ;
        RECT 178.200 56.200 178.600 59.900 ;
        RECT 179.800 56.200 180.200 59.900 ;
        RECT 178.200 55.900 180.200 56.200 ;
        RECT 172.700 55.500 174.600 55.800 ;
        RECT 172.700 54.500 173.000 55.500 ;
        RECT 164.600 53.400 165.000 53.800 ;
        RECT 166.900 53.500 167.200 53.800 ;
        RECT 167.700 53.900 168.200 54.100 ;
        RECT 167.700 53.600 169.800 53.900 ;
        RECT 171.000 53.800 172.000 54.200 ;
        RECT 172.300 54.100 173.000 54.500 ;
        RECT 173.400 54.400 173.800 55.200 ;
        RECT 174.200 54.400 174.600 55.200 ;
        RECT 175.900 54.200 176.200 55.900 ;
        RECT 176.600 54.800 177.000 55.600 ;
        RECT 177.500 55.200 177.800 55.900 ;
        RECT 180.600 55.600 181.000 59.900 ;
        RECT 182.700 57.900 183.300 59.900 ;
        RECT 185.000 57.900 185.400 59.900 ;
        RECT 187.200 58.200 187.600 59.900 ;
        RECT 187.200 57.900 188.200 58.200 ;
        RECT 183.000 57.500 183.400 57.900 ;
        RECT 185.100 57.600 185.400 57.900 ;
        RECT 184.700 57.300 186.500 57.600 ;
        RECT 187.800 57.500 188.200 57.900 ;
        RECT 184.700 57.200 185.100 57.300 ;
        RECT 186.100 57.200 186.500 57.300 ;
        RECT 182.600 56.600 183.300 57.000 ;
        RECT 183.000 56.100 183.300 56.600 ;
        RECT 184.100 56.500 185.200 56.800 ;
        RECT 184.100 56.400 184.500 56.500 ;
        RECT 183.000 55.800 184.200 56.100 ;
        RECT 179.400 55.200 179.800 55.400 ;
        RECT 180.600 55.300 182.700 55.600 ;
        RECT 177.400 54.900 178.600 55.200 ;
        RECT 179.400 54.900 180.200 55.200 ;
        RECT 177.400 54.800 177.800 54.900 ;
        RECT 178.200 54.800 178.600 54.900 ;
        RECT 179.800 54.800 180.200 54.900 ;
        RECT 159.800 53.000 161.800 53.100 ;
        RECT 159.800 51.100 160.200 53.000 ;
        RECT 161.400 51.100 161.800 53.000 ;
        RECT 162.200 51.100 162.600 53.100 ;
        RECT 163.300 52.800 164.200 53.100 ;
        RECT 166.900 53.300 167.300 53.500 ;
        RECT 166.900 53.000 167.700 53.300 ;
        RECT 163.300 51.100 163.700 52.800 ;
        RECT 167.300 51.500 167.700 53.000 ;
        RECT 169.500 52.500 169.800 53.600 ;
        RECT 171.700 53.500 172.000 53.800 ;
        RECT 172.500 53.900 173.000 54.100 ;
        RECT 172.500 53.600 174.600 53.900 ;
        RECT 175.800 53.800 176.200 54.200 ;
        RECT 171.700 53.300 172.100 53.500 ;
        RECT 171.700 53.000 172.500 53.300 ;
        RECT 169.400 51.500 169.800 52.500 ;
        RECT 172.100 51.500 172.500 53.000 ;
        RECT 174.300 52.500 174.600 53.600 ;
        RECT 174.200 51.500 174.600 52.500 ;
        RECT 175.000 52.400 175.400 53.200 ;
        RECT 175.900 53.100 176.200 53.800 ;
        RECT 177.400 53.100 177.800 53.200 ;
        RECT 178.300 53.100 178.600 54.800 ;
        RECT 179.000 53.800 179.400 54.600 ;
        RECT 175.800 52.800 177.800 53.100 ;
        RECT 175.900 52.100 176.200 52.800 ;
        RECT 177.500 52.400 177.900 52.800 ;
        RECT 175.800 51.100 176.200 52.100 ;
        RECT 178.200 51.100 178.600 53.100 ;
        RECT 180.600 53.600 181.000 55.300 ;
        RECT 182.300 55.200 182.700 55.300 ;
        RECT 181.500 54.900 181.900 55.000 ;
        RECT 181.500 54.600 183.400 54.900 ;
        RECT 183.000 54.500 183.400 54.600 ;
        RECT 183.900 54.200 184.200 55.800 ;
        RECT 184.900 55.900 185.200 56.500 ;
        RECT 185.500 56.500 185.900 56.600 ;
        RECT 187.800 56.500 188.200 56.600 ;
        RECT 185.500 56.200 188.200 56.500 ;
        RECT 184.900 55.700 187.300 55.900 ;
        RECT 189.400 55.700 189.800 59.900 ;
        RECT 184.900 55.600 189.800 55.700 ;
        RECT 186.900 55.500 189.800 55.600 ;
        RECT 190.200 57.500 190.600 59.500 ;
        RECT 190.200 55.800 190.500 57.500 ;
        RECT 192.300 56.400 192.700 59.900 ;
        RECT 192.300 56.100 193.100 56.400 ;
        RECT 190.200 55.500 192.100 55.800 ;
        RECT 187.000 55.400 189.800 55.500 ;
        RECT 185.400 55.100 185.800 55.200 ;
        RECT 186.200 55.100 186.600 55.200 ;
        RECT 185.400 54.800 188.700 55.100 ;
        RECT 188.300 54.700 188.700 54.800 ;
        RECT 190.200 54.400 190.600 55.200 ;
        RECT 191.000 54.400 191.400 55.200 ;
        RECT 191.800 54.500 192.100 55.500 ;
        RECT 187.500 54.200 187.900 54.300 ;
        RECT 183.900 53.900 189.400 54.200 ;
        RECT 191.800 54.100 192.500 54.500 ;
        RECT 192.800 54.200 193.100 56.100 ;
        RECT 193.400 55.100 193.800 55.600 ;
        RECT 195.000 55.100 195.400 59.900 ;
        RECT 196.600 57.500 197.000 59.500 ;
        RECT 196.600 55.800 196.900 57.500 ;
        RECT 198.700 56.400 199.100 59.900 ;
        RECT 201.400 57.500 201.800 59.500 ;
        RECT 203.500 59.200 203.900 59.900 ;
        RECT 203.500 58.800 204.200 59.200 ;
        RECT 198.700 56.100 199.500 56.400 ;
        RECT 199.000 55.800 199.500 56.100 ;
        RECT 196.600 55.500 198.500 55.800 ;
        RECT 193.400 54.800 195.400 55.100 ;
        RECT 191.800 53.900 192.300 54.100 ;
        RECT 184.100 53.800 184.500 53.900 ;
        RECT 185.400 53.800 185.800 53.900 ;
        RECT 180.600 53.300 182.500 53.600 ;
        RECT 180.600 51.100 181.000 53.300 ;
        RECT 182.100 53.200 182.500 53.300 ;
        RECT 187.000 52.800 187.300 53.900 ;
        RECT 188.600 53.800 189.400 53.900 ;
        RECT 190.200 53.600 192.300 53.900 ;
        RECT 192.800 53.800 193.800 54.200 ;
        RECT 186.100 52.700 186.500 52.800 ;
        RECT 183.000 52.100 183.400 52.500 ;
        RECT 185.100 52.400 186.500 52.700 ;
        RECT 187.000 52.400 187.400 52.800 ;
        RECT 185.100 52.100 185.400 52.400 ;
        RECT 187.800 52.100 188.200 52.500 ;
        RECT 182.700 51.800 183.400 52.100 ;
        RECT 182.700 51.100 183.300 51.800 ;
        RECT 185.000 51.100 185.400 52.100 ;
        RECT 187.200 51.800 188.200 52.100 ;
        RECT 187.200 51.100 187.600 51.800 ;
        RECT 189.400 51.100 189.800 53.500 ;
        RECT 190.200 52.500 190.500 53.600 ;
        RECT 192.800 53.500 193.100 53.800 ;
        RECT 192.700 53.300 193.100 53.500 ;
        RECT 192.300 53.000 193.100 53.300 ;
        RECT 190.200 51.500 190.600 52.500 ;
        RECT 192.300 52.200 192.700 53.000 ;
        RECT 191.800 51.800 192.700 52.200 ;
        RECT 192.300 51.500 192.700 51.800 ;
        RECT 195.000 51.100 195.400 54.800 ;
        RECT 196.600 54.400 197.000 55.200 ;
        RECT 197.400 54.400 197.800 55.200 ;
        RECT 198.200 54.500 198.500 55.500 ;
        RECT 198.200 54.100 198.900 54.500 ;
        RECT 199.200 54.200 199.500 55.800 ;
        RECT 201.400 55.800 201.700 57.500 ;
        RECT 203.500 56.400 203.900 58.800 ;
        RECT 203.500 56.100 204.300 56.400 ;
        RECT 199.800 54.800 200.200 55.600 ;
        RECT 201.400 55.500 203.300 55.800 ;
        RECT 201.400 54.400 201.800 55.200 ;
        RECT 202.200 54.400 202.600 55.200 ;
        RECT 203.000 54.500 203.300 55.500 ;
        RECT 198.200 53.900 198.700 54.100 ;
        RECT 196.600 53.600 198.700 53.900 ;
        RECT 199.200 53.800 200.200 54.200 ;
        RECT 203.000 54.100 203.700 54.500 ;
        RECT 204.000 54.200 204.300 56.100 ;
        RECT 207.500 56.200 207.900 59.900 ;
        RECT 208.200 56.800 208.600 57.200 ;
        RECT 208.300 56.200 208.600 56.800 ;
        RECT 207.500 55.900 208.000 56.200 ;
        RECT 208.300 55.900 209.000 56.200 ;
        RECT 204.600 54.800 205.000 55.600 ;
        RECT 206.200 55.100 206.600 55.200 ;
        RECT 207.000 55.100 207.400 55.200 ;
        RECT 206.200 54.800 207.400 55.100 ;
        RECT 207.000 54.400 207.400 54.800 ;
        RECT 207.700 55.100 208.000 55.900 ;
        RECT 208.600 55.800 209.000 55.900 ;
        RECT 211.000 55.700 211.400 59.900 ;
        RECT 213.200 58.200 213.600 59.900 ;
        RECT 212.600 57.900 213.600 58.200 ;
        RECT 215.400 57.900 215.800 59.900 ;
        RECT 217.500 57.900 218.100 59.900 ;
        RECT 212.600 57.500 213.000 57.900 ;
        RECT 215.400 57.600 215.700 57.900 ;
        RECT 214.300 57.300 216.100 57.600 ;
        RECT 217.400 57.500 217.800 57.900 ;
        RECT 214.300 57.200 214.700 57.300 ;
        RECT 215.700 57.200 216.100 57.300 ;
        RECT 212.600 56.500 213.000 56.600 ;
        RECT 214.900 56.500 215.300 56.600 ;
        RECT 212.600 56.200 215.300 56.500 ;
        RECT 215.600 56.500 216.700 56.800 ;
        RECT 215.600 55.900 215.900 56.500 ;
        RECT 216.300 56.400 216.700 56.500 ;
        RECT 217.500 56.600 218.200 57.000 ;
        RECT 217.500 56.100 217.800 56.600 ;
        RECT 213.500 55.700 215.900 55.900 ;
        RECT 211.000 55.600 215.900 55.700 ;
        RECT 216.600 55.800 217.800 56.100 ;
        RECT 211.000 55.500 213.900 55.600 ;
        RECT 211.000 55.400 213.800 55.500 ;
        RECT 209.400 55.100 209.800 55.200 ;
        RECT 214.200 55.100 214.600 55.200 ;
        RECT 207.700 54.800 209.800 55.100 ;
        RECT 212.100 54.800 214.600 55.100 ;
        RECT 207.700 54.200 208.000 54.800 ;
        RECT 212.100 54.700 212.500 54.800 ;
        RECT 213.400 54.700 213.800 54.800 ;
        RECT 212.900 54.200 213.300 54.300 ;
        RECT 216.600 54.200 216.900 55.800 ;
        RECT 219.800 55.600 220.200 59.900 ;
        RECT 222.500 59.200 222.900 59.900 ;
        RECT 222.200 58.800 222.900 59.200 ;
        RECT 222.500 56.400 222.900 58.800 ;
        RECT 224.600 57.500 225.000 59.500 ;
        RECT 222.100 56.100 222.900 56.400 ;
        RECT 218.100 55.300 220.200 55.600 ;
        RECT 218.100 55.200 218.500 55.300 ;
        RECT 218.900 54.900 219.300 55.000 ;
        RECT 217.400 54.600 219.300 54.900 ;
        RECT 217.400 54.500 217.800 54.600 ;
        RECT 203.000 53.900 203.500 54.100 ;
        RECT 195.800 52.400 196.200 53.200 ;
        RECT 196.600 52.500 196.900 53.600 ;
        RECT 199.200 53.500 199.500 53.800 ;
        RECT 199.100 53.300 199.500 53.500 ;
        RECT 198.700 53.000 199.500 53.300 ;
        RECT 201.400 53.600 203.500 53.900 ;
        RECT 204.000 53.800 205.000 54.200 ;
        RECT 205.400 54.100 205.800 54.200 ;
        RECT 206.200 54.100 206.600 54.200 ;
        RECT 205.400 53.800 207.000 54.100 ;
        RECT 207.700 53.800 209.000 54.200 ;
        RECT 211.400 53.900 216.900 54.200 ;
        RECT 211.400 53.800 212.200 53.900 ;
        RECT 196.600 51.500 197.000 52.500 ;
        RECT 198.700 51.500 199.100 53.000 ;
        RECT 201.400 52.500 201.700 53.600 ;
        RECT 204.000 53.500 204.300 53.800 ;
        RECT 206.600 53.600 207.000 53.800 ;
        RECT 203.900 53.300 204.300 53.500 ;
        RECT 203.500 53.000 204.300 53.300 ;
        RECT 206.300 53.100 208.100 53.300 ;
        RECT 208.600 53.100 208.900 53.800 ;
        RECT 206.200 53.000 208.200 53.100 ;
        RECT 201.400 51.500 201.800 52.500 ;
        RECT 203.500 51.500 203.900 53.000 ;
        RECT 206.200 51.100 206.600 53.000 ;
        RECT 207.800 51.100 208.200 53.000 ;
        RECT 208.600 51.100 209.000 53.100 ;
        RECT 211.000 51.100 211.400 53.500 ;
        RECT 213.500 52.800 213.800 53.900 ;
        RECT 216.300 53.800 216.700 53.900 ;
        RECT 219.800 53.600 220.200 55.300 ;
        RECT 220.600 55.100 221.000 55.200 ;
        RECT 221.400 55.100 221.800 55.600 ;
        RECT 220.600 54.800 221.800 55.100 ;
        RECT 222.100 54.200 222.400 56.100 ;
        RECT 224.700 55.800 225.000 57.500 ;
        RECT 223.100 55.500 225.000 55.800 ;
        RECT 225.400 57.500 225.800 59.500 ;
        RECT 227.500 59.200 227.900 59.900 ;
        RECT 227.000 58.800 227.900 59.200 ;
        RECT 225.400 55.800 225.700 57.500 ;
        RECT 227.500 56.400 227.900 58.800 ;
        RECT 230.200 57.500 230.600 59.500 ;
        RECT 227.500 56.100 228.300 56.400 ;
        RECT 225.400 55.500 227.300 55.800 ;
        RECT 223.100 54.500 223.400 55.500 ;
        RECT 221.400 53.800 222.400 54.200 ;
        RECT 222.700 54.100 223.400 54.500 ;
        RECT 223.800 54.400 224.200 55.200 ;
        RECT 224.600 54.400 225.000 55.200 ;
        RECT 225.400 54.400 225.800 55.200 ;
        RECT 226.200 54.400 226.600 55.200 ;
        RECT 227.000 54.500 227.300 55.500 ;
        RECT 218.300 53.300 220.200 53.600 ;
        RECT 218.300 53.200 218.700 53.300 ;
        RECT 212.600 52.100 213.000 52.500 ;
        RECT 213.400 52.400 213.800 52.800 ;
        RECT 214.300 52.700 214.700 52.800 ;
        RECT 214.300 52.400 215.700 52.700 ;
        RECT 215.400 52.100 215.700 52.400 ;
        RECT 217.400 52.100 217.800 52.500 ;
        RECT 212.600 51.800 213.600 52.100 ;
        RECT 213.200 51.100 213.600 51.800 ;
        RECT 215.400 51.100 215.800 52.100 ;
        RECT 217.400 51.800 218.100 52.100 ;
        RECT 217.500 51.100 218.100 51.800 ;
        RECT 219.800 51.100 220.200 53.300 ;
        RECT 222.100 53.500 222.400 53.800 ;
        RECT 222.900 53.900 223.400 54.100 ;
        RECT 227.000 54.100 227.700 54.500 ;
        RECT 228.000 54.200 228.300 56.100 ;
        RECT 230.200 55.800 230.500 57.500 ;
        RECT 232.300 56.400 232.700 59.900 ;
        RECT 232.300 56.100 233.100 56.400 ;
        RECT 228.600 54.800 229.000 55.600 ;
        RECT 230.200 55.500 232.100 55.800 ;
        RECT 229.400 55.100 229.800 55.200 ;
        RECT 230.200 55.100 230.600 55.200 ;
        RECT 229.400 54.800 230.600 55.100 ;
        RECT 230.200 54.400 230.600 54.800 ;
        RECT 231.000 54.400 231.400 55.200 ;
        RECT 231.800 54.500 232.100 55.500 ;
        RECT 227.000 53.900 227.500 54.100 ;
        RECT 222.900 53.600 225.000 53.900 ;
        RECT 222.100 53.300 222.500 53.500 ;
        RECT 222.100 53.000 222.900 53.300 ;
        RECT 222.500 51.500 222.900 53.000 ;
        RECT 224.700 52.500 225.000 53.600 ;
        RECT 224.600 51.500 225.000 52.500 ;
        RECT 225.400 53.600 227.500 53.900 ;
        RECT 228.000 53.800 229.000 54.200 ;
        RECT 231.800 54.100 232.500 54.500 ;
        RECT 232.800 54.200 233.100 56.100 ;
        RECT 236.300 56.200 236.700 59.900 ;
        RECT 237.000 56.800 237.400 57.200 ;
        RECT 237.100 56.200 237.400 56.800 ;
        RECT 236.300 55.900 236.800 56.200 ;
        RECT 237.100 55.900 237.800 56.200 ;
        RECT 233.400 55.100 233.800 55.600 ;
        RECT 236.500 55.200 236.800 55.900 ;
        RECT 237.400 55.800 237.800 55.900 ;
        RECT 238.200 55.700 238.600 59.900 ;
        RECT 240.400 58.200 240.800 59.900 ;
        RECT 239.800 57.900 240.800 58.200 ;
        RECT 242.600 57.900 243.000 59.900 ;
        RECT 244.700 57.900 245.300 59.900 ;
        RECT 239.800 57.500 240.200 57.900 ;
        RECT 242.600 57.600 242.900 57.900 ;
        RECT 241.500 57.300 243.300 57.600 ;
        RECT 244.600 57.500 245.000 57.900 ;
        RECT 241.500 57.200 241.900 57.300 ;
        RECT 242.900 57.200 243.300 57.300 ;
        RECT 239.800 56.500 240.200 56.600 ;
        RECT 242.100 56.500 242.500 56.600 ;
        RECT 239.800 56.200 242.500 56.500 ;
        RECT 242.800 56.500 243.900 56.800 ;
        RECT 242.800 55.900 243.100 56.500 ;
        RECT 243.500 56.400 243.900 56.500 ;
        RECT 244.700 56.600 245.400 57.000 ;
        RECT 244.700 56.100 245.000 56.600 ;
        RECT 240.700 55.700 243.100 55.900 ;
        RECT 238.200 55.600 243.100 55.700 ;
        RECT 243.800 55.800 245.000 56.100 ;
        RECT 238.200 55.500 241.100 55.600 ;
        RECT 238.200 55.400 241.000 55.500 ;
        RECT 235.000 55.100 235.400 55.200 ;
        RECT 233.400 54.800 235.400 55.100 ;
        RECT 235.800 54.400 236.200 55.200 ;
        RECT 236.500 54.800 237.000 55.200 ;
        RECT 241.400 55.100 241.800 55.200 ;
        RECT 239.300 54.800 241.800 55.100 ;
        RECT 236.500 54.200 236.800 54.800 ;
        RECT 239.300 54.700 239.700 54.800 ;
        RECT 240.600 54.700 241.000 54.800 ;
        RECT 240.100 54.200 240.500 54.300 ;
        RECT 243.800 54.200 244.100 55.800 ;
        RECT 247.000 55.600 247.400 59.900 ;
        RECT 249.100 56.200 249.500 59.900 ;
        RECT 249.800 56.800 250.200 57.200 ;
        RECT 249.900 56.200 250.200 56.800 ;
        RECT 249.100 55.900 249.600 56.200 ;
        RECT 249.900 55.900 250.600 56.200 ;
        RECT 245.300 55.300 247.400 55.600 ;
        RECT 245.300 55.200 245.700 55.300 ;
        RECT 246.100 54.900 246.500 55.000 ;
        RECT 244.600 54.600 246.500 54.900 ;
        RECT 244.600 54.500 245.000 54.600 ;
        RECT 231.800 53.900 232.300 54.100 ;
        RECT 225.400 52.500 225.700 53.600 ;
        RECT 228.000 53.500 228.300 53.800 ;
        RECT 227.900 53.300 228.300 53.500 ;
        RECT 227.500 53.000 228.300 53.300 ;
        RECT 230.200 53.600 232.300 53.900 ;
        RECT 232.800 53.800 233.800 54.200 ;
        RECT 234.200 54.100 234.600 54.200 ;
        RECT 235.000 54.100 235.400 54.200 ;
        RECT 234.200 53.800 235.800 54.100 ;
        RECT 236.500 53.800 237.800 54.200 ;
        RECT 238.600 53.900 244.100 54.200 ;
        RECT 238.600 53.800 239.400 53.900 ;
        RECT 225.400 51.500 225.800 52.500 ;
        RECT 227.500 51.500 227.900 53.000 ;
        RECT 230.200 52.500 230.500 53.600 ;
        RECT 232.800 53.500 233.100 53.800 ;
        RECT 235.400 53.600 235.800 53.800 ;
        RECT 232.700 53.300 233.100 53.500 ;
        RECT 232.300 53.200 233.100 53.300 ;
        RECT 231.800 53.000 233.100 53.200 ;
        RECT 235.100 53.100 236.900 53.300 ;
        RECT 237.400 53.100 237.700 53.800 ;
        RECT 235.000 53.000 237.000 53.100 ;
        RECT 231.800 52.800 232.700 53.000 ;
        RECT 230.200 51.500 230.600 52.500 ;
        RECT 232.300 51.500 232.700 52.800 ;
        RECT 235.000 51.100 235.400 53.000 ;
        RECT 236.600 51.100 237.000 53.000 ;
        RECT 237.400 51.100 237.800 53.100 ;
        RECT 238.200 51.100 238.600 53.500 ;
        RECT 240.700 52.800 241.000 53.900 ;
        RECT 243.500 53.800 243.900 53.900 ;
        RECT 247.000 53.600 247.400 55.300 ;
        RECT 248.600 54.400 249.000 55.200 ;
        RECT 249.300 54.200 249.600 55.900 ;
        RECT 250.200 55.800 250.600 55.900 ;
        RECT 251.000 55.800 251.400 56.600 ;
        RECT 250.200 55.100 250.500 55.800 ;
        RECT 251.800 55.100 252.200 59.900 ;
        RECT 253.400 57.500 253.800 59.500 ;
        RECT 255.500 59.200 255.900 59.900 ;
        RECT 255.500 58.800 256.200 59.200 ;
        RECT 253.400 55.800 253.700 57.500 ;
        RECT 255.500 56.400 255.900 58.800 ;
        RECT 258.200 57.100 258.600 57.200 ;
        RECT 259.000 57.100 259.400 59.900 ;
        RECT 261.900 59.200 262.300 59.900 ;
        RECT 261.400 58.800 262.300 59.200 ;
        RECT 258.200 56.800 259.400 57.100 ;
        RECT 255.500 56.100 256.300 56.400 ;
        RECT 253.400 55.500 255.300 55.800 ;
        RECT 250.200 54.800 252.200 55.100 ;
        RECT 247.800 54.100 248.200 54.200 ;
        RECT 247.800 53.800 248.600 54.100 ;
        RECT 249.300 53.800 250.600 54.200 ;
        RECT 248.200 53.600 248.600 53.800 ;
        RECT 245.500 53.300 247.400 53.600 ;
        RECT 245.500 53.200 245.900 53.300 ;
        RECT 239.800 52.100 240.200 52.500 ;
        RECT 240.600 52.400 241.000 52.800 ;
        RECT 241.500 52.700 241.900 52.800 ;
        RECT 241.500 52.400 242.900 52.700 ;
        RECT 242.600 52.100 242.900 52.400 ;
        RECT 244.600 52.100 245.000 52.500 ;
        RECT 239.800 51.800 240.800 52.100 ;
        RECT 240.400 51.100 240.800 51.800 ;
        RECT 242.600 51.100 243.000 52.100 ;
        RECT 244.600 51.800 245.300 52.100 ;
        RECT 244.700 51.100 245.300 51.800 ;
        RECT 247.000 51.100 247.400 53.300 ;
        RECT 247.900 53.100 249.700 53.300 ;
        RECT 250.200 53.100 250.500 53.800 ;
        RECT 251.800 53.100 252.200 54.800 ;
        RECT 253.400 54.400 253.800 55.200 ;
        RECT 254.200 54.400 254.600 55.200 ;
        RECT 255.000 54.500 255.300 55.500 ;
        RECT 252.600 53.400 253.000 54.200 ;
        RECT 255.000 54.100 255.700 54.500 ;
        RECT 256.000 54.200 256.300 56.100 ;
        RECT 256.600 54.800 257.000 55.600 ;
        RECT 255.000 53.900 255.500 54.100 ;
        RECT 253.400 53.600 255.500 53.900 ;
        RECT 256.000 53.800 257.000 54.200 ;
        RECT 257.400 54.100 257.800 54.200 ;
        RECT 258.200 54.100 258.600 54.200 ;
        RECT 257.400 53.800 258.600 54.100 ;
        RECT 247.800 53.000 249.800 53.100 ;
        RECT 247.800 51.100 248.200 53.000 ;
        RECT 249.400 51.100 249.800 53.000 ;
        RECT 250.200 51.100 250.600 53.100 ;
        RECT 251.300 52.800 252.200 53.100 ;
        RECT 251.300 51.100 251.700 52.800 ;
        RECT 253.400 52.500 253.700 53.600 ;
        RECT 256.000 53.500 256.300 53.800 ;
        RECT 255.900 53.300 256.300 53.500 ;
        RECT 258.200 53.400 258.600 53.800 ;
        RECT 255.500 53.000 256.300 53.300 ;
        RECT 259.000 53.100 259.400 56.800 ;
        RECT 259.800 55.800 260.200 56.600 ;
        RECT 261.900 56.200 262.300 58.800 ;
        RECT 262.600 56.800 263.000 57.200 ;
        RECT 262.700 56.200 263.000 56.800 ;
        RECT 261.900 55.900 262.400 56.200 ;
        RECT 262.700 55.900 263.400 56.200 ;
        RECT 259.800 55.100 260.100 55.800 ;
        RECT 261.400 55.100 261.800 55.200 ;
        RECT 259.800 54.800 261.800 55.100 ;
        RECT 261.400 54.400 261.800 54.800 ;
        RECT 262.100 54.200 262.400 55.900 ;
        RECT 263.000 55.800 263.400 55.900 ;
        RECT 260.600 54.100 261.000 54.200 ;
        RECT 260.600 53.800 261.400 54.100 ;
        RECT 262.100 53.800 263.400 54.200 ;
        RECT 261.000 53.600 261.400 53.800 ;
        RECT 260.700 53.100 262.500 53.300 ;
        RECT 263.000 53.100 263.300 53.800 ;
        RECT 253.400 51.500 253.800 52.500 ;
        RECT 255.500 51.500 255.900 53.000 ;
        RECT 259.000 52.800 259.900 53.100 ;
        RECT 259.500 51.100 259.900 52.800 ;
        RECT 260.600 53.000 262.600 53.100 ;
        RECT 260.600 51.100 261.000 53.000 ;
        RECT 262.200 51.100 262.600 53.000 ;
        RECT 263.000 51.100 263.400 53.100 ;
        RECT 0.600 47.500 1.000 49.900 ;
        RECT 2.800 49.200 3.200 49.900 ;
        RECT 2.200 48.900 3.200 49.200 ;
        RECT 5.000 48.900 5.400 49.900 ;
        RECT 7.100 49.200 7.700 49.900 ;
        RECT 7.000 48.900 7.700 49.200 ;
        RECT 2.200 48.500 2.600 48.900 ;
        RECT 5.000 48.600 5.300 48.900 ;
        RECT 3.000 48.200 3.400 48.600 ;
        RECT 3.900 48.300 5.300 48.600 ;
        RECT 7.000 48.500 7.400 48.900 ;
        RECT 3.900 48.200 4.300 48.300 ;
        RECT 1.000 47.100 1.800 47.200 ;
        RECT 3.100 47.100 3.400 48.200 ;
        RECT 9.400 48.100 9.800 49.900 ;
        RECT 10.200 48.100 10.600 48.600 ;
        RECT 9.400 47.800 10.600 48.100 ;
        RECT 7.900 47.700 8.300 47.800 ;
        RECT 9.400 47.700 9.800 47.800 ;
        RECT 7.900 47.400 9.800 47.700 ;
        RECT 5.900 47.100 6.300 47.200 ;
        RECT 1.000 46.800 6.500 47.100 ;
        RECT 2.500 46.700 2.900 46.800 ;
        RECT 1.700 46.200 2.100 46.300 ;
        RECT 1.700 45.900 4.200 46.200 ;
        RECT 3.800 45.800 4.200 45.900 ;
        RECT 5.400 46.100 5.800 46.200 ;
        RECT 6.200 46.100 6.500 46.800 ;
        RECT 7.000 46.400 7.400 46.500 ;
        RECT 7.000 46.100 8.900 46.400 ;
        RECT 5.400 45.800 6.500 46.100 ;
        RECT 8.500 46.000 8.900 46.100 ;
        RECT 0.600 45.500 3.400 45.600 ;
        RECT 0.600 45.400 3.500 45.500 ;
        RECT 0.600 45.300 5.500 45.400 ;
        RECT 0.600 41.100 1.000 45.300 ;
        RECT 3.100 45.100 5.500 45.300 ;
        RECT 2.200 44.500 4.900 44.800 ;
        RECT 2.200 44.400 2.600 44.500 ;
        RECT 4.500 44.400 4.900 44.500 ;
        RECT 5.200 44.500 5.500 45.100 ;
        RECT 6.200 45.200 6.500 45.800 ;
        RECT 7.700 45.700 8.100 45.800 ;
        RECT 9.400 45.700 9.800 47.400 ;
        RECT 7.700 45.400 9.800 45.700 ;
        RECT 6.200 44.900 7.400 45.200 ;
        RECT 5.900 44.500 6.300 44.600 ;
        RECT 5.200 44.200 6.300 44.500 ;
        RECT 7.100 44.400 7.400 44.900 ;
        RECT 7.100 44.200 7.800 44.400 ;
        RECT 7.100 44.000 8.200 44.200 ;
        RECT 7.500 43.800 8.200 44.000 ;
        RECT 3.900 43.700 4.300 43.800 ;
        RECT 5.300 43.700 5.700 43.800 ;
        RECT 2.200 43.100 2.600 43.500 ;
        RECT 3.900 43.400 5.700 43.700 ;
        RECT 5.000 43.100 5.300 43.400 ;
        RECT 7.000 43.100 7.400 43.500 ;
        RECT 2.200 42.800 3.200 43.100 ;
        RECT 2.800 41.100 3.200 42.800 ;
        RECT 5.000 41.100 5.400 43.100 ;
        RECT 7.100 41.100 7.700 43.100 ;
        RECT 9.400 41.100 9.800 45.400 ;
        RECT 11.000 46.100 11.400 49.900 ;
        RECT 13.700 48.000 14.100 49.500 ;
        RECT 15.800 48.500 16.200 49.500 ;
        RECT 13.300 47.700 14.100 48.000 ;
        RECT 13.300 47.500 13.700 47.700 ;
        RECT 13.300 47.200 13.600 47.500 ;
        RECT 15.900 47.400 16.200 48.500 ;
        RECT 11.800 47.100 12.200 47.200 ;
        RECT 12.600 47.100 13.600 47.200 ;
        RECT 11.800 46.800 13.600 47.100 ;
        RECT 14.100 47.100 16.200 47.400 ;
        RECT 16.600 47.700 17.000 49.900 ;
        RECT 18.700 49.200 19.300 49.900 ;
        RECT 18.700 48.900 19.400 49.200 ;
        RECT 21.000 48.900 21.400 49.900 ;
        RECT 23.200 49.200 23.600 49.900 ;
        RECT 23.200 48.900 24.200 49.200 ;
        RECT 19.000 48.500 19.400 48.900 ;
        RECT 21.100 48.600 21.400 48.900 ;
        RECT 21.100 48.300 22.500 48.600 ;
        RECT 22.100 48.200 22.500 48.300 ;
        RECT 23.000 48.200 23.400 48.600 ;
        RECT 23.800 48.500 24.200 48.900 ;
        RECT 18.100 47.700 18.500 47.800 ;
        RECT 16.600 47.400 18.500 47.700 ;
        RECT 14.100 46.900 14.600 47.100 ;
        RECT 12.600 46.100 13.000 46.200 ;
        RECT 11.000 45.800 13.000 46.100 ;
        RECT 11.000 41.100 11.400 45.800 ;
        RECT 12.600 45.400 13.000 45.800 ;
        RECT 13.300 44.900 13.600 46.800 ;
        RECT 13.900 46.500 14.600 46.900 ;
        RECT 14.300 45.500 14.600 46.500 ;
        RECT 15.000 45.800 15.400 46.600 ;
        RECT 15.800 45.800 16.200 46.600 ;
        RECT 16.600 45.700 17.000 47.400 ;
        RECT 20.100 47.100 20.500 47.200 ;
        RECT 23.000 47.100 23.300 48.200 ;
        RECT 25.400 47.500 25.800 49.900 ;
        RECT 26.200 47.800 26.600 48.600 ;
        RECT 24.600 47.100 25.400 47.200 ;
        RECT 19.900 46.800 26.500 47.100 ;
        RECT 19.000 46.400 19.400 46.500 ;
        RECT 17.500 46.100 19.400 46.400 ;
        RECT 19.900 46.100 20.200 46.800 ;
        RECT 23.500 46.700 23.900 46.800 ;
        RECT 23.000 46.200 23.400 46.300 ;
        RECT 24.300 46.200 24.700 46.300 ;
        RECT 20.600 46.100 21.000 46.200 ;
        RECT 17.500 46.000 17.900 46.100 ;
        RECT 19.800 45.800 21.000 46.100 ;
        RECT 22.200 45.900 24.700 46.200 ;
        RECT 26.200 46.200 26.500 46.800 ;
        RECT 22.200 45.800 22.600 45.900 ;
        RECT 26.200 45.800 26.600 46.200 ;
        RECT 27.000 46.100 27.400 49.900 ;
        RECT 29.700 48.000 30.100 49.500 ;
        RECT 31.800 48.500 32.200 49.500 ;
        RECT 29.300 47.700 30.100 48.000 ;
        RECT 29.300 47.500 29.700 47.700 ;
        RECT 29.300 47.200 29.600 47.500 ;
        RECT 31.900 47.400 32.200 48.500 ;
        RECT 27.800 47.100 28.200 47.200 ;
        RECT 28.600 47.100 29.600 47.200 ;
        RECT 27.800 46.800 29.600 47.100 ;
        RECT 30.100 47.100 32.200 47.400 ;
        RECT 32.600 47.700 33.000 49.900 ;
        RECT 34.700 49.200 35.300 49.900 ;
        RECT 34.700 48.900 35.400 49.200 ;
        RECT 37.000 48.900 37.400 49.900 ;
        RECT 39.200 49.200 39.600 49.900 ;
        RECT 39.200 48.900 40.200 49.200 ;
        RECT 35.000 48.500 35.400 48.900 ;
        RECT 37.100 48.600 37.400 48.900 ;
        RECT 37.100 48.300 38.500 48.600 ;
        RECT 38.100 48.200 38.500 48.300 ;
        RECT 39.000 47.800 39.400 48.600 ;
        RECT 39.800 48.500 40.200 48.900 ;
        RECT 34.100 47.700 34.500 47.800 ;
        RECT 32.600 47.400 34.500 47.700 ;
        RECT 30.100 46.900 30.600 47.100 ;
        RECT 28.600 46.100 29.000 46.200 ;
        RECT 27.000 45.800 29.000 46.100 ;
        RECT 18.300 45.700 18.700 45.800 ;
        RECT 14.300 45.200 16.200 45.500 ;
        RECT 13.300 44.600 14.100 44.900 ;
        RECT 13.700 41.100 14.100 44.600 ;
        RECT 15.900 43.500 16.200 45.200 ;
        RECT 15.800 41.500 16.200 43.500 ;
        RECT 16.600 45.400 18.700 45.700 ;
        RECT 16.600 41.100 17.000 45.400 ;
        RECT 19.900 45.200 20.200 45.800 ;
        RECT 23.000 45.500 25.800 45.600 ;
        RECT 22.900 45.400 25.800 45.500 ;
        RECT 19.000 44.900 20.200 45.200 ;
        RECT 20.900 45.300 25.800 45.400 ;
        RECT 20.900 45.100 23.300 45.300 ;
        RECT 19.000 44.400 19.300 44.900 ;
        RECT 18.600 44.000 19.300 44.400 ;
        RECT 20.100 44.500 20.500 44.600 ;
        RECT 20.900 44.500 21.200 45.100 ;
        RECT 20.100 44.200 21.200 44.500 ;
        RECT 21.500 44.500 24.200 44.800 ;
        RECT 21.500 44.400 21.900 44.500 ;
        RECT 23.800 44.400 24.200 44.500 ;
        RECT 20.700 43.700 21.100 43.800 ;
        RECT 22.100 43.700 22.500 43.800 ;
        RECT 19.000 43.100 19.400 43.500 ;
        RECT 20.700 43.400 22.500 43.700 ;
        RECT 21.100 43.100 21.400 43.400 ;
        RECT 23.800 43.100 24.200 43.500 ;
        RECT 18.700 41.100 19.300 43.100 ;
        RECT 21.000 41.100 21.400 43.100 ;
        RECT 23.200 42.800 24.200 43.100 ;
        RECT 23.200 41.100 23.600 42.800 ;
        RECT 25.400 41.100 25.800 45.300 ;
        RECT 27.000 41.100 27.400 45.800 ;
        RECT 28.600 45.400 29.000 45.800 ;
        RECT 29.300 44.900 29.600 46.800 ;
        RECT 29.900 46.500 30.600 46.900 ;
        RECT 30.300 45.500 30.600 46.500 ;
        RECT 31.000 45.800 31.400 46.600 ;
        RECT 31.800 45.800 32.200 46.600 ;
        RECT 32.600 45.700 33.000 47.400 ;
        RECT 36.100 47.100 36.500 47.200 ;
        RECT 39.000 47.100 39.300 47.800 ;
        RECT 41.400 47.500 41.800 49.900 ;
        RECT 42.200 47.700 42.600 49.900 ;
        RECT 44.300 49.200 44.900 49.900 ;
        RECT 44.300 48.900 45.000 49.200 ;
        RECT 46.600 48.900 47.000 49.900 ;
        RECT 48.800 49.200 49.200 49.900 ;
        RECT 48.800 48.900 49.800 49.200 ;
        RECT 44.600 48.500 45.000 48.900 ;
        RECT 46.700 48.600 47.000 48.900 ;
        RECT 46.700 48.300 48.100 48.600 ;
        RECT 47.700 48.200 48.100 48.300 ;
        RECT 48.600 48.200 49.000 48.600 ;
        RECT 49.400 48.500 49.800 48.900 ;
        RECT 43.700 47.700 44.100 47.800 ;
        RECT 42.200 47.400 44.100 47.700 ;
        RECT 40.600 47.100 41.400 47.200 ;
        RECT 35.900 46.800 41.400 47.100 ;
        RECT 35.000 46.400 35.400 46.500 ;
        RECT 33.500 46.100 35.400 46.400 ;
        RECT 33.500 46.000 33.900 46.100 ;
        RECT 34.300 45.700 34.700 45.800 ;
        RECT 30.300 45.200 32.200 45.500 ;
        RECT 29.300 44.600 30.100 44.900 ;
        RECT 29.700 41.100 30.100 44.600 ;
        RECT 31.900 43.500 32.200 45.200 ;
        RECT 31.800 41.500 32.200 43.500 ;
        RECT 32.600 45.400 34.700 45.700 ;
        RECT 32.600 41.100 33.000 45.400 ;
        RECT 35.900 45.200 36.200 46.800 ;
        RECT 39.500 46.700 39.900 46.800 ;
        RECT 40.300 46.200 40.700 46.300 ;
        RECT 38.200 45.900 40.700 46.200 ;
        RECT 38.200 45.800 38.600 45.900 ;
        RECT 42.200 45.700 42.600 47.400 ;
        RECT 45.700 47.100 46.100 47.200 ;
        RECT 48.600 47.100 48.900 48.200 ;
        RECT 51.000 47.500 51.400 49.900 ;
        RECT 53.100 48.200 53.500 49.900 ;
        RECT 52.600 47.900 53.500 48.200 ;
        RECT 55.800 47.900 56.200 49.900 ;
        RECT 56.600 48.000 57.000 49.900 ;
        RECT 58.200 48.000 58.600 49.900 ;
        RECT 59.800 48.200 60.200 49.900 ;
        RECT 56.600 47.900 58.600 48.000 ;
        RECT 59.700 47.900 60.200 48.200 ;
        RECT 50.200 47.100 51.000 47.200 ;
        RECT 45.500 46.800 51.000 47.100 ;
        RECT 51.800 46.800 52.200 47.600 ;
        RECT 44.600 46.400 45.000 46.500 ;
        RECT 43.100 46.100 45.000 46.400 ;
        RECT 43.100 46.000 43.500 46.100 ;
        RECT 43.900 45.700 44.300 45.800 ;
        RECT 39.000 45.500 41.800 45.600 ;
        RECT 38.900 45.400 41.800 45.500 ;
        RECT 35.000 44.900 36.200 45.200 ;
        RECT 36.900 45.300 41.800 45.400 ;
        RECT 36.900 45.100 39.300 45.300 ;
        RECT 35.000 44.400 35.300 44.900 ;
        RECT 34.600 44.000 35.300 44.400 ;
        RECT 36.100 44.500 36.500 44.600 ;
        RECT 36.900 44.500 37.200 45.100 ;
        RECT 36.100 44.200 37.200 44.500 ;
        RECT 37.500 44.500 40.200 44.800 ;
        RECT 37.500 44.400 37.900 44.500 ;
        RECT 39.800 44.400 40.200 44.500 ;
        RECT 36.700 43.700 37.100 43.800 ;
        RECT 38.100 43.700 38.500 43.800 ;
        RECT 35.000 43.100 35.400 43.500 ;
        RECT 36.700 43.400 38.500 43.700 ;
        RECT 37.100 43.100 37.400 43.400 ;
        RECT 39.800 43.100 40.200 43.500 ;
        RECT 34.700 41.100 35.300 43.100 ;
        RECT 37.000 41.100 37.400 43.100 ;
        RECT 39.200 42.800 40.200 43.100 ;
        RECT 39.200 41.100 39.600 42.800 ;
        RECT 41.400 41.100 41.800 45.300 ;
        RECT 42.200 45.400 44.300 45.700 ;
        RECT 42.200 41.100 42.600 45.400 ;
        RECT 45.500 45.200 45.800 46.800 ;
        RECT 49.100 46.700 49.500 46.800 ;
        RECT 48.600 46.200 49.000 46.300 ;
        RECT 49.900 46.200 50.300 46.300 ;
        RECT 47.800 45.900 50.300 46.200 ;
        RECT 52.600 46.100 53.000 47.900 ;
        RECT 55.900 47.200 56.200 47.900 ;
        RECT 56.700 47.700 58.500 47.900 ;
        RECT 57.800 47.200 58.200 47.400 ;
        RECT 59.700 47.200 60.000 47.900 ;
        RECT 61.400 47.600 61.800 49.900 ;
        RECT 60.500 47.300 61.800 47.600 ;
        RECT 62.200 47.700 62.600 49.900 ;
        RECT 64.300 49.200 64.900 49.900 ;
        RECT 64.300 48.900 65.000 49.200 ;
        RECT 66.600 48.900 67.000 49.900 ;
        RECT 68.800 49.200 69.200 49.900 ;
        RECT 68.800 48.900 69.800 49.200 ;
        RECT 64.600 48.500 65.000 48.900 ;
        RECT 66.700 48.600 67.000 48.900 ;
        RECT 66.700 48.300 68.100 48.600 ;
        RECT 67.700 48.200 68.100 48.300 ;
        RECT 68.600 48.200 69.000 48.600 ;
        RECT 69.400 48.500 69.800 48.900 ;
        RECT 63.700 47.700 64.100 47.800 ;
        RECT 62.200 47.400 64.100 47.700 ;
        RECT 54.200 47.100 54.600 47.200 ;
        RECT 55.800 47.100 57.100 47.200 ;
        RECT 54.200 46.800 57.100 47.100 ;
        RECT 57.800 46.900 58.600 47.200 ;
        RECT 58.200 46.800 58.600 46.900 ;
        RECT 59.700 46.800 60.200 47.200 ;
        RECT 47.800 45.800 48.200 45.900 ;
        RECT 52.600 45.800 56.100 46.100 ;
        RECT 48.600 45.500 51.400 45.600 ;
        RECT 48.500 45.400 51.400 45.500 ;
        RECT 44.600 44.900 45.800 45.200 ;
        RECT 46.500 45.300 51.400 45.400 ;
        RECT 46.500 45.100 48.900 45.300 ;
        RECT 44.600 44.400 44.900 44.900 ;
        RECT 44.200 44.000 44.900 44.400 ;
        RECT 45.700 44.500 46.100 44.600 ;
        RECT 46.500 44.500 46.800 45.100 ;
        RECT 45.700 44.200 46.800 44.500 ;
        RECT 47.100 44.500 49.800 44.800 ;
        RECT 47.100 44.400 47.500 44.500 ;
        RECT 49.400 44.400 49.800 44.500 ;
        RECT 46.300 43.700 46.700 43.800 ;
        RECT 47.700 43.700 48.100 43.800 ;
        RECT 44.600 43.100 45.000 43.500 ;
        RECT 46.300 43.400 48.100 43.700 ;
        RECT 46.700 43.100 47.000 43.400 ;
        RECT 49.400 43.100 49.800 43.500 ;
        RECT 44.300 41.100 44.900 43.100 ;
        RECT 46.600 41.100 47.000 43.100 ;
        RECT 48.800 42.800 49.800 43.100 ;
        RECT 48.800 41.100 49.200 42.800 ;
        RECT 51.000 41.100 51.400 45.300 ;
        RECT 52.600 41.100 53.000 45.800 ;
        RECT 55.800 45.200 56.100 45.800 ;
        RECT 53.400 44.400 53.800 45.200 ;
        RECT 55.800 45.100 56.200 45.200 ;
        RECT 56.800 45.100 57.100 46.800 ;
        RECT 57.400 45.800 57.800 46.600 ;
        RECT 59.700 45.100 60.000 46.800 ;
        RECT 60.500 46.500 60.800 47.300 ;
        RECT 60.300 46.100 60.800 46.500 ;
        RECT 60.500 45.100 60.800 46.100 ;
        RECT 61.300 46.200 61.700 46.600 ;
        RECT 61.300 45.800 61.800 46.200 ;
        RECT 62.200 45.700 62.600 47.400 ;
        RECT 65.700 47.100 66.100 47.200 ;
        RECT 68.600 47.100 68.900 48.200 ;
        RECT 71.000 47.500 71.400 49.900 ;
        RECT 71.800 47.700 72.200 49.900 ;
        RECT 73.900 49.200 74.500 49.900 ;
        RECT 73.900 48.900 74.600 49.200 ;
        RECT 76.200 48.900 76.600 49.900 ;
        RECT 78.400 49.200 78.800 49.900 ;
        RECT 78.400 48.900 79.400 49.200 ;
        RECT 74.200 48.500 74.600 48.900 ;
        RECT 76.300 48.600 76.600 48.900 ;
        RECT 76.300 48.300 77.700 48.600 ;
        RECT 77.300 48.200 77.700 48.300 ;
        RECT 78.200 48.200 78.600 48.600 ;
        RECT 79.000 48.500 79.400 48.900 ;
        RECT 73.300 47.700 73.700 47.800 ;
        RECT 71.800 47.400 73.700 47.700 ;
        RECT 70.200 47.100 71.000 47.200 ;
        RECT 65.500 46.800 71.000 47.100 ;
        RECT 64.600 46.400 65.000 46.500 ;
        RECT 63.100 46.100 65.000 46.400 ;
        RECT 63.100 46.000 63.500 46.100 ;
        RECT 63.900 45.700 64.300 45.800 ;
        RECT 62.200 45.400 64.300 45.700 ;
        RECT 55.800 44.800 56.500 45.100 ;
        RECT 56.800 44.800 57.300 45.100 ;
        RECT 56.200 44.200 56.500 44.800 ;
        RECT 56.200 43.800 56.600 44.200 ;
        RECT 56.900 41.100 57.300 44.800 ;
        RECT 59.700 44.600 60.200 45.100 ;
        RECT 60.500 44.800 61.800 45.100 ;
        RECT 59.800 41.100 60.200 44.600 ;
        RECT 61.400 41.100 61.800 44.800 ;
        RECT 62.200 41.100 62.600 45.400 ;
        RECT 65.500 45.200 65.800 46.800 ;
        RECT 69.100 46.700 69.500 46.800 ;
        RECT 68.600 46.200 69.000 46.300 ;
        RECT 69.900 46.200 70.300 46.300 ;
        RECT 67.800 45.900 70.300 46.200 ;
        RECT 67.800 45.800 68.200 45.900 ;
        RECT 71.800 45.700 72.200 47.400 ;
        RECT 75.300 47.100 75.700 47.200 ;
        RECT 78.200 47.100 78.500 48.200 ;
        RECT 80.600 47.500 81.000 49.900 ;
        RECT 81.400 48.000 81.800 49.900 ;
        RECT 83.000 48.000 83.400 49.900 ;
        RECT 81.400 47.900 83.400 48.000 ;
        RECT 83.800 47.900 84.200 49.900 ;
        RECT 84.900 48.200 85.300 49.900 ;
        RECT 84.900 47.900 85.800 48.200 ;
        RECT 81.500 47.700 83.300 47.900 ;
        RECT 81.800 47.200 82.200 47.400 ;
        RECT 83.800 47.200 84.100 47.900 ;
        RECT 79.800 47.100 80.600 47.200 ;
        RECT 75.100 46.800 80.600 47.100 ;
        RECT 81.400 46.900 82.200 47.200 ;
        RECT 81.400 46.800 81.800 46.900 ;
        RECT 82.900 46.800 84.200 47.200 ;
        RECT 74.200 46.400 74.600 46.500 ;
        RECT 72.700 46.100 74.600 46.400 ;
        RECT 72.700 46.000 73.100 46.100 ;
        RECT 73.500 45.700 73.900 45.800 ;
        RECT 68.600 45.500 71.400 45.600 ;
        RECT 68.500 45.400 71.400 45.500 ;
        RECT 64.600 44.900 65.800 45.200 ;
        RECT 66.500 45.300 71.400 45.400 ;
        RECT 66.500 45.100 68.900 45.300 ;
        RECT 64.600 44.400 64.900 44.900 ;
        RECT 64.200 44.000 64.900 44.400 ;
        RECT 65.700 44.500 66.100 44.600 ;
        RECT 66.500 44.500 66.800 45.100 ;
        RECT 65.700 44.200 66.800 44.500 ;
        RECT 67.100 44.500 69.800 44.800 ;
        RECT 67.100 44.400 67.500 44.500 ;
        RECT 69.400 44.400 69.800 44.500 ;
        RECT 66.300 43.700 66.700 43.800 ;
        RECT 67.700 43.700 68.100 43.800 ;
        RECT 64.600 43.100 65.000 43.500 ;
        RECT 66.300 43.400 68.100 43.700 ;
        RECT 66.700 43.100 67.000 43.400 ;
        RECT 69.400 43.100 69.800 43.500 ;
        RECT 64.300 41.100 64.900 43.100 ;
        RECT 66.600 41.100 67.000 43.100 ;
        RECT 68.800 42.800 69.800 43.100 ;
        RECT 68.800 41.100 69.200 42.800 ;
        RECT 71.000 41.100 71.400 45.300 ;
        RECT 71.800 45.400 73.900 45.700 ;
        RECT 71.800 41.100 72.200 45.400 ;
        RECT 75.100 45.200 75.400 46.800 ;
        RECT 78.700 46.700 79.100 46.800 ;
        RECT 78.200 46.200 78.600 46.300 ;
        RECT 79.500 46.200 79.900 46.300 ;
        RECT 77.400 45.900 79.900 46.200 ;
        RECT 77.400 45.800 77.800 45.900 ;
        RECT 82.200 45.800 82.600 46.600 ;
        RECT 78.200 45.500 81.000 45.600 ;
        RECT 78.100 45.400 81.000 45.500 ;
        RECT 74.200 44.900 75.400 45.200 ;
        RECT 76.100 45.300 81.000 45.400 ;
        RECT 76.100 45.100 78.500 45.300 ;
        RECT 74.200 44.400 74.500 44.900 ;
        RECT 73.800 44.000 74.500 44.400 ;
        RECT 75.300 44.500 75.700 44.600 ;
        RECT 76.100 44.500 76.400 45.100 ;
        RECT 75.300 44.200 76.400 44.500 ;
        RECT 76.700 44.500 79.400 44.800 ;
        RECT 76.700 44.400 77.100 44.500 ;
        RECT 79.000 44.400 79.400 44.500 ;
        RECT 75.900 43.700 76.300 43.800 ;
        RECT 77.300 43.700 77.700 43.800 ;
        RECT 74.200 43.100 74.600 43.500 ;
        RECT 75.900 43.400 77.700 43.700 ;
        RECT 76.300 43.100 76.600 43.400 ;
        RECT 79.000 43.100 79.400 43.500 ;
        RECT 73.900 41.100 74.500 43.100 ;
        RECT 76.200 41.100 76.600 43.100 ;
        RECT 78.400 42.800 79.400 43.100 ;
        RECT 78.400 41.100 78.800 42.800 ;
        RECT 80.600 41.100 81.000 45.300 ;
        RECT 82.900 45.200 83.200 46.800 ;
        RECT 85.400 46.100 85.800 47.900 ;
        RECT 86.200 46.800 86.600 47.600 ;
        RECT 87.000 47.500 87.400 49.900 ;
        RECT 89.200 49.200 89.600 49.900 ;
        RECT 88.600 48.900 89.600 49.200 ;
        RECT 91.400 48.900 91.800 49.900 ;
        RECT 93.500 49.200 94.100 49.900 ;
        RECT 93.400 48.900 94.100 49.200 ;
        RECT 88.600 48.500 89.000 48.900 ;
        RECT 91.400 48.600 91.700 48.900 ;
        RECT 89.400 48.200 89.800 48.600 ;
        RECT 90.300 48.300 91.700 48.600 ;
        RECT 93.400 48.500 93.800 48.900 ;
        RECT 90.300 48.200 90.700 48.300 ;
        RECT 87.400 47.100 88.200 47.200 ;
        RECT 89.500 47.100 89.800 48.200 ;
        RECT 94.300 47.700 94.700 47.800 ;
        RECT 95.800 47.700 96.200 49.900 ;
        RECT 97.900 48.200 98.300 49.900 ;
        RECT 94.300 47.400 96.200 47.700 ;
        RECT 97.400 47.900 98.300 48.200 ;
        RECT 92.300 47.100 92.700 47.200 ;
        RECT 87.400 46.800 92.900 47.100 ;
        RECT 95.000 46.800 95.400 47.400 ;
        RECT 95.800 47.100 96.200 47.400 ;
        RECT 96.600 47.100 97.000 47.600 ;
        RECT 95.800 46.800 97.000 47.100 ;
        RECT 88.900 46.700 89.300 46.800 ;
        RECT 82.200 44.800 83.200 45.200 ;
        RECT 83.800 45.800 85.800 46.100 ;
        RECT 88.100 46.200 88.500 46.300 ;
        RECT 92.600 46.200 92.900 46.800 ;
        RECT 93.400 46.400 93.800 46.500 ;
        RECT 88.100 45.900 90.600 46.200 ;
        RECT 90.200 45.800 90.600 45.900 ;
        RECT 92.600 45.800 93.000 46.200 ;
        RECT 93.400 46.100 95.300 46.400 ;
        RECT 94.900 46.000 95.300 46.100 ;
        RECT 83.800 45.200 84.100 45.800 ;
        RECT 83.800 45.100 84.200 45.200 ;
        RECT 83.500 44.800 84.200 45.100 ;
        RECT 82.700 41.100 83.100 44.800 ;
        RECT 83.500 44.200 83.800 44.800 ;
        RECT 84.600 44.400 85.000 45.200 ;
        RECT 83.400 43.800 83.800 44.200 ;
        RECT 85.400 41.100 85.800 45.800 ;
        RECT 87.000 45.500 89.800 45.600 ;
        RECT 87.000 45.400 89.900 45.500 ;
        RECT 87.000 45.300 91.900 45.400 ;
        RECT 87.000 41.100 87.400 45.300 ;
        RECT 89.500 45.100 91.900 45.300 ;
        RECT 88.600 44.500 91.300 44.800 ;
        RECT 88.600 44.400 89.000 44.500 ;
        RECT 90.900 44.400 91.300 44.500 ;
        RECT 91.600 44.500 91.900 45.100 ;
        RECT 92.600 45.200 92.900 45.800 ;
        RECT 94.100 45.700 94.500 45.800 ;
        RECT 95.800 45.700 96.200 46.800 ;
        RECT 94.100 45.400 96.200 45.700 ;
        RECT 92.600 44.900 93.800 45.200 ;
        RECT 92.300 44.500 92.700 44.600 ;
        RECT 91.600 44.200 92.700 44.500 ;
        RECT 93.500 44.400 93.800 44.900 ;
        RECT 93.500 44.000 94.200 44.400 ;
        RECT 90.300 43.700 90.700 43.800 ;
        RECT 91.700 43.700 92.100 43.800 ;
        RECT 88.600 43.100 89.000 43.500 ;
        RECT 90.300 43.400 92.100 43.700 ;
        RECT 91.400 43.100 91.700 43.400 ;
        RECT 93.400 43.100 93.800 43.500 ;
        RECT 88.600 42.800 89.600 43.100 ;
        RECT 89.200 41.100 89.600 42.800 ;
        RECT 91.400 41.100 91.800 43.100 ;
        RECT 93.500 41.100 94.100 43.100 ;
        RECT 95.800 41.100 96.200 45.400 ;
        RECT 97.400 46.100 97.800 47.900 ;
        RECT 99.000 47.800 99.400 49.900 ;
        RECT 99.800 48.000 100.200 49.900 ;
        RECT 101.400 48.000 101.800 49.900 ;
        RECT 99.800 47.900 101.800 48.000 ;
        RECT 99.100 47.200 99.400 47.800 ;
        RECT 99.900 47.700 101.700 47.900 ;
        RECT 103.800 47.700 104.200 49.900 ;
        RECT 105.900 49.200 106.500 49.900 ;
        RECT 105.900 48.900 106.600 49.200 ;
        RECT 108.200 48.900 108.600 49.900 ;
        RECT 110.400 49.200 110.800 49.900 ;
        RECT 110.400 48.900 111.400 49.200 ;
        RECT 106.200 48.500 106.600 48.900 ;
        RECT 108.300 48.600 108.600 48.900 ;
        RECT 108.300 48.300 109.700 48.600 ;
        RECT 109.300 48.200 109.700 48.300 ;
        RECT 110.200 48.200 110.600 48.600 ;
        RECT 111.000 48.500 111.400 48.900 ;
        RECT 105.300 47.700 105.700 47.800 ;
        RECT 103.800 47.400 105.700 47.700 ;
        RECT 101.000 47.200 101.400 47.400 ;
        RECT 99.000 46.800 100.300 47.200 ;
        RECT 101.000 46.900 101.800 47.200 ;
        RECT 101.400 46.800 101.800 46.900 ;
        RECT 97.400 45.800 99.300 46.100 ;
        RECT 97.400 41.100 97.800 45.800 ;
        RECT 99.000 45.200 99.300 45.800 ;
        RECT 98.200 44.400 98.600 45.200 ;
        RECT 99.000 45.100 99.400 45.200 ;
        RECT 100.000 45.100 100.300 46.800 ;
        RECT 100.600 46.100 101.000 46.600 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 100.600 45.800 103.400 46.100 ;
        RECT 103.800 45.700 104.200 47.400 ;
        RECT 110.200 47.200 110.500 48.200 ;
        RECT 112.600 47.500 113.000 49.900 ;
        RECT 113.400 47.500 113.800 49.900 ;
        RECT 115.600 49.200 116.000 49.900 ;
        RECT 115.000 48.900 116.000 49.200 ;
        RECT 117.800 48.900 118.200 49.900 ;
        RECT 119.900 49.200 120.500 49.900 ;
        RECT 119.800 48.900 120.500 49.200 ;
        RECT 115.000 48.500 115.400 48.900 ;
        RECT 117.800 48.600 118.100 48.900 ;
        RECT 115.800 48.200 116.200 48.600 ;
        RECT 116.700 48.300 118.100 48.600 ;
        RECT 119.800 48.500 120.200 48.900 ;
        RECT 116.700 48.200 117.100 48.300 ;
        RECT 107.300 47.100 107.700 47.200 ;
        RECT 110.200 47.100 110.600 47.200 ;
        RECT 111.800 47.100 112.600 47.200 ;
        RECT 107.100 46.800 112.600 47.100 ;
        RECT 113.800 47.100 114.600 47.200 ;
        RECT 115.900 47.100 116.200 48.200 ;
        RECT 120.700 47.700 121.100 47.800 ;
        RECT 122.200 47.700 122.600 49.900 ;
        RECT 123.000 47.900 123.400 49.900 ;
        RECT 123.800 48.000 124.200 49.900 ;
        RECT 125.400 48.000 125.800 49.900 ;
        RECT 123.800 47.900 125.800 48.000 ;
        RECT 126.200 47.900 126.600 49.900 ;
        RECT 127.000 48.000 127.400 49.900 ;
        RECT 128.600 48.000 129.000 49.900 ;
        RECT 127.000 47.900 129.000 48.000 ;
        RECT 120.700 47.400 122.600 47.700 ;
        RECT 118.700 47.100 119.100 47.200 ;
        RECT 113.800 46.800 119.300 47.100 ;
        RECT 106.200 46.400 106.600 46.500 ;
        RECT 104.700 46.100 106.600 46.400 ;
        RECT 104.700 46.000 105.100 46.100 ;
        RECT 105.500 45.700 105.900 45.800 ;
        RECT 103.800 45.400 105.900 45.700 ;
        RECT 99.000 44.800 99.700 45.100 ;
        RECT 100.000 44.800 100.500 45.100 ;
        RECT 99.400 44.200 99.700 44.800 ;
        RECT 99.400 43.800 99.800 44.200 ;
        RECT 100.100 41.100 100.500 44.800 ;
        RECT 103.800 41.100 104.200 45.400 ;
        RECT 107.100 45.200 107.400 46.800 ;
        RECT 110.700 46.700 111.100 46.800 ;
        RECT 115.300 46.700 115.700 46.800 ;
        RECT 111.500 46.200 111.900 46.300 ;
        RECT 109.400 45.900 111.900 46.200 ;
        RECT 114.500 46.200 114.900 46.300 ;
        RECT 114.500 46.100 117.000 46.200 ;
        RECT 117.400 46.100 117.800 46.200 ;
        RECT 114.500 45.900 117.800 46.100 ;
        RECT 109.400 45.800 109.800 45.900 ;
        RECT 116.600 45.800 117.800 45.900 ;
        RECT 110.200 45.500 113.000 45.600 ;
        RECT 110.100 45.400 113.000 45.500 ;
        RECT 106.200 44.900 107.400 45.200 ;
        RECT 108.100 45.300 113.000 45.400 ;
        RECT 108.100 45.100 110.500 45.300 ;
        RECT 106.200 44.400 106.500 44.900 ;
        RECT 105.800 44.000 106.500 44.400 ;
        RECT 107.300 44.500 107.700 44.600 ;
        RECT 108.100 44.500 108.400 45.100 ;
        RECT 107.300 44.200 108.400 44.500 ;
        RECT 108.700 44.500 111.400 44.800 ;
        RECT 108.700 44.400 109.100 44.500 ;
        RECT 111.000 44.400 111.400 44.500 ;
        RECT 107.900 43.700 108.300 43.800 ;
        RECT 109.300 43.700 109.700 43.800 ;
        RECT 106.200 43.100 106.600 43.500 ;
        RECT 107.900 43.400 109.700 43.700 ;
        RECT 108.300 43.100 108.600 43.400 ;
        RECT 111.000 43.100 111.400 43.500 ;
        RECT 105.900 41.100 106.500 43.100 ;
        RECT 108.200 41.100 108.600 43.100 ;
        RECT 110.400 42.800 111.400 43.100 ;
        RECT 110.400 41.100 110.800 42.800 ;
        RECT 112.600 41.100 113.000 45.300 ;
        RECT 113.400 45.500 116.200 45.600 ;
        RECT 113.400 45.400 116.300 45.500 ;
        RECT 113.400 45.300 118.300 45.400 ;
        RECT 113.400 41.100 113.800 45.300 ;
        RECT 115.900 45.100 118.300 45.300 ;
        RECT 115.000 44.500 117.700 44.800 ;
        RECT 115.000 44.400 115.400 44.500 ;
        RECT 117.300 44.400 117.700 44.500 ;
        RECT 118.000 44.500 118.300 45.100 ;
        RECT 119.000 45.200 119.300 46.800 ;
        RECT 119.800 46.400 120.200 46.500 ;
        RECT 119.800 46.100 121.700 46.400 ;
        RECT 121.300 46.000 121.700 46.100 ;
        RECT 120.500 45.700 120.900 45.800 ;
        RECT 122.200 45.700 122.600 47.400 ;
        RECT 123.100 47.200 123.400 47.900 ;
        RECT 123.900 47.700 125.700 47.900 ;
        RECT 125.000 47.200 125.400 47.400 ;
        RECT 126.300 47.200 126.600 47.900 ;
        RECT 127.100 47.700 128.900 47.900 ;
        RECT 129.400 47.500 129.800 49.900 ;
        RECT 131.600 49.200 132.000 49.900 ;
        RECT 131.000 48.900 132.000 49.200 ;
        RECT 133.800 48.900 134.200 49.900 ;
        RECT 135.900 49.200 136.500 49.900 ;
        RECT 135.800 48.900 136.500 49.200 ;
        RECT 131.000 48.500 131.400 48.900 ;
        RECT 133.800 48.600 134.100 48.900 ;
        RECT 131.800 47.800 132.200 48.600 ;
        RECT 132.700 48.300 134.100 48.600 ;
        RECT 135.800 48.500 136.200 48.900 ;
        RECT 132.700 48.200 133.100 48.300 ;
        RECT 128.200 47.200 128.600 47.400 ;
        RECT 123.000 46.800 124.300 47.200 ;
        RECT 125.000 46.900 125.800 47.200 ;
        RECT 125.400 46.800 125.800 46.900 ;
        RECT 126.200 46.800 127.500 47.200 ;
        RECT 128.200 46.900 129.000 47.200 ;
        RECT 128.600 46.800 129.000 46.900 ;
        RECT 129.800 47.100 130.600 47.200 ;
        RECT 131.900 47.100 132.200 47.800 ;
        RECT 136.700 47.700 137.100 47.800 ;
        RECT 138.200 47.700 138.600 49.900 ;
        RECT 139.000 48.000 139.400 49.900 ;
        RECT 140.600 48.000 141.000 49.900 ;
        RECT 139.000 47.900 141.000 48.000 ;
        RECT 141.400 47.900 141.800 49.900 ;
        RECT 142.200 47.900 142.600 49.900 ;
        RECT 143.000 48.000 143.400 49.900 ;
        RECT 144.600 48.000 145.000 49.900 ;
        RECT 143.000 47.900 145.000 48.000 ;
        RECT 145.400 48.500 145.800 49.500 ;
        RECT 139.100 47.700 140.900 47.900 ;
        RECT 136.700 47.400 138.600 47.700 ;
        RECT 134.700 47.100 135.100 47.200 ;
        RECT 129.800 46.800 135.300 47.100 ;
        RECT 120.500 45.400 122.600 45.700 ;
        RECT 119.000 44.900 120.200 45.200 ;
        RECT 118.700 44.500 119.100 44.600 ;
        RECT 118.000 44.200 119.100 44.500 ;
        RECT 119.900 44.400 120.200 44.900 ;
        RECT 119.900 44.000 120.600 44.400 ;
        RECT 116.700 43.700 117.100 43.800 ;
        RECT 118.100 43.700 118.500 43.800 ;
        RECT 115.000 43.100 115.400 43.500 ;
        RECT 116.700 43.400 118.500 43.700 ;
        RECT 117.800 43.100 118.100 43.400 ;
        RECT 119.800 43.100 120.200 43.500 ;
        RECT 115.000 42.800 116.000 43.100 ;
        RECT 115.600 41.100 116.000 42.800 ;
        RECT 117.800 41.100 118.200 43.100 ;
        RECT 119.900 41.100 120.500 43.100 ;
        RECT 122.200 41.100 122.600 45.400 ;
        RECT 123.000 45.100 123.400 45.200 ;
        RECT 124.000 45.100 124.300 46.800 ;
        RECT 124.600 45.800 125.000 46.600 ;
        RECT 126.200 45.100 126.600 45.200 ;
        RECT 127.200 45.100 127.500 46.800 ;
        RECT 131.300 46.700 131.700 46.800 ;
        RECT 127.800 45.800 128.200 46.600 ;
        RECT 130.500 46.200 130.900 46.300 ;
        RECT 130.500 45.900 133.000 46.200 ;
        RECT 132.600 45.800 133.000 45.900 ;
        RECT 129.400 45.500 132.200 45.600 ;
        RECT 129.400 45.400 132.300 45.500 ;
        RECT 129.400 45.300 134.300 45.400 ;
        RECT 123.000 44.800 123.700 45.100 ;
        RECT 124.000 44.800 124.500 45.100 ;
        RECT 126.200 44.800 126.900 45.100 ;
        RECT 127.200 44.800 127.700 45.100 ;
        RECT 123.400 44.200 123.700 44.800 ;
        RECT 123.400 43.800 123.800 44.200 ;
        RECT 124.100 41.100 124.500 44.800 ;
        RECT 126.600 44.200 126.900 44.800 ;
        RECT 126.200 43.800 127.000 44.200 ;
        RECT 127.300 41.100 127.700 44.800 ;
        RECT 129.400 41.100 129.800 45.300 ;
        RECT 131.900 45.100 134.300 45.300 ;
        RECT 131.000 44.500 133.700 44.800 ;
        RECT 131.000 44.400 131.400 44.500 ;
        RECT 133.300 44.400 133.700 44.500 ;
        RECT 134.000 44.500 134.300 45.100 ;
        RECT 135.000 45.200 135.300 46.800 ;
        RECT 135.800 46.400 136.200 46.500 ;
        RECT 135.800 46.100 137.700 46.400 ;
        RECT 137.300 46.000 137.700 46.100 ;
        RECT 136.500 45.700 136.900 45.800 ;
        RECT 138.200 45.700 138.600 47.400 ;
        RECT 139.400 47.200 139.800 47.400 ;
        RECT 141.400 47.200 141.700 47.900 ;
        RECT 142.300 47.200 142.600 47.900 ;
        RECT 143.100 47.700 144.900 47.900 ;
        RECT 145.400 47.400 145.700 48.500 ;
        RECT 147.500 48.000 147.900 49.500 ;
        RECT 147.500 47.700 148.300 48.000 ;
        RECT 147.900 47.500 148.300 47.700 ;
        RECT 144.200 47.200 144.600 47.400 ;
        RECT 139.000 46.900 139.800 47.200 ;
        RECT 139.000 46.800 139.400 46.900 ;
        RECT 140.500 46.800 141.800 47.200 ;
        RECT 142.200 46.800 143.500 47.200 ;
        RECT 144.200 46.900 145.000 47.200 ;
        RECT 145.400 47.100 147.500 47.400 ;
        RECT 144.600 46.800 145.000 46.900 ;
        RECT 147.000 46.900 147.500 47.100 ;
        RECT 148.000 47.200 148.300 47.500 ;
        RECT 139.800 45.800 140.200 46.600 ;
        RECT 136.500 45.400 138.600 45.700 ;
        RECT 135.000 44.900 136.200 45.200 ;
        RECT 134.700 44.500 135.100 44.600 ;
        RECT 134.000 44.200 135.100 44.500 ;
        RECT 135.900 44.400 136.200 44.900 ;
        RECT 135.900 44.000 136.600 44.400 ;
        RECT 132.700 43.700 133.100 43.800 ;
        RECT 134.100 43.700 134.500 43.800 ;
        RECT 131.000 43.100 131.400 43.500 ;
        RECT 132.700 43.400 134.500 43.700 ;
        RECT 133.800 43.100 134.100 43.400 ;
        RECT 135.800 43.100 136.200 43.500 ;
        RECT 131.000 42.800 132.000 43.100 ;
        RECT 131.600 41.100 132.000 42.800 ;
        RECT 133.800 41.100 134.200 43.100 ;
        RECT 135.900 41.100 136.500 43.100 ;
        RECT 138.200 41.100 138.600 45.400 ;
        RECT 140.500 45.100 140.800 46.800 ;
        RECT 143.200 46.100 143.500 46.800 ;
        RECT 141.400 45.800 143.500 46.100 ;
        RECT 143.800 45.800 144.200 46.600 ;
        RECT 145.400 45.800 145.800 46.600 ;
        RECT 146.200 45.800 146.600 46.600 ;
        RECT 147.000 46.500 147.700 46.900 ;
        RECT 148.000 46.800 149.000 47.200 ;
        RECT 141.400 45.200 141.700 45.800 ;
        RECT 141.400 45.100 141.800 45.200 ;
        RECT 140.300 44.800 140.800 45.100 ;
        RECT 141.100 44.800 141.800 45.100 ;
        RECT 142.200 45.100 142.600 45.200 ;
        RECT 143.200 45.100 143.500 45.800 ;
        RECT 147.000 45.500 147.300 46.500 ;
        RECT 145.400 45.200 147.300 45.500 ;
        RECT 142.200 44.800 142.900 45.100 ;
        RECT 143.200 44.800 143.700 45.100 ;
        RECT 140.300 43.200 140.700 44.800 ;
        RECT 141.100 44.200 141.400 44.800 ;
        RECT 141.000 43.800 141.400 44.200 ;
        RECT 142.600 44.200 142.900 44.800 ;
        RECT 142.600 43.800 143.000 44.200 ;
        RECT 139.800 42.800 140.700 43.200 ;
        RECT 140.300 41.100 140.700 42.800 ;
        RECT 143.300 41.100 143.700 44.800 ;
        RECT 145.400 43.500 145.700 45.200 ;
        RECT 148.000 44.900 148.300 46.800 ;
        RECT 148.600 46.100 149.000 46.200 ;
        RECT 150.200 46.100 150.600 49.900 ;
        RECT 151.000 47.800 151.400 48.600 ;
        RECT 153.100 48.200 153.500 49.900 ;
        RECT 152.600 47.900 153.500 48.200 ;
        RECT 154.200 47.900 154.600 49.900 ;
        RECT 155.000 48.000 155.400 49.900 ;
        RECT 156.600 48.000 157.000 49.900 ;
        RECT 155.000 47.900 157.000 48.000 ;
        RECT 151.800 46.800 152.200 47.600 ;
        RECT 148.600 45.800 150.600 46.100 ;
        RECT 148.600 45.400 149.000 45.800 ;
        RECT 147.500 44.600 148.300 44.900 ;
        RECT 145.400 41.500 145.800 43.500 ;
        RECT 147.500 42.200 147.900 44.600 ;
        RECT 147.000 41.800 147.900 42.200 ;
        RECT 147.500 41.100 147.900 41.800 ;
        RECT 150.200 41.100 150.600 45.800 ;
        RECT 152.600 46.100 153.000 47.900 ;
        RECT 154.300 47.200 154.600 47.900 ;
        RECT 155.100 47.700 156.900 47.900 ;
        RECT 159.000 47.700 159.400 49.900 ;
        RECT 161.100 49.200 161.700 49.900 ;
        RECT 161.100 48.900 161.800 49.200 ;
        RECT 163.400 48.900 163.800 49.900 ;
        RECT 165.600 49.200 166.000 49.900 ;
        RECT 165.600 48.900 166.600 49.200 ;
        RECT 161.400 48.500 161.800 48.900 ;
        RECT 163.500 48.600 163.800 48.900 ;
        RECT 163.500 48.300 164.900 48.600 ;
        RECT 164.500 48.200 164.900 48.300 ;
        RECT 165.400 48.200 165.800 48.600 ;
        RECT 166.200 48.500 166.600 48.900 ;
        RECT 160.500 47.700 160.900 47.800 ;
        RECT 159.000 47.400 160.900 47.700 ;
        RECT 156.200 47.200 156.600 47.400 ;
        RECT 154.200 46.800 155.500 47.200 ;
        RECT 156.200 46.900 157.000 47.200 ;
        RECT 156.600 46.800 157.000 46.900 ;
        RECT 152.600 45.800 154.500 46.100 ;
        RECT 152.600 41.100 153.000 45.800 ;
        RECT 154.200 45.200 154.500 45.800 ;
        RECT 155.200 45.200 155.500 46.800 ;
        RECT 155.800 45.800 156.200 46.600 ;
        RECT 159.000 45.700 159.400 47.400 ;
        RECT 162.500 47.100 162.900 47.200 ;
        RECT 165.400 47.100 165.700 48.200 ;
        RECT 167.800 47.500 168.200 49.900 ;
        RECT 168.600 47.600 169.000 49.900 ;
        RECT 170.200 48.200 170.600 49.900 ;
        RECT 170.200 47.900 170.700 48.200 ;
        RECT 171.800 48.000 172.200 49.900 ;
        RECT 173.400 48.000 173.800 49.900 ;
        RECT 171.800 47.900 173.800 48.000 ;
        RECT 174.200 47.900 174.600 49.900 ;
        RECT 175.300 48.200 175.700 49.900 ;
        RECT 175.300 47.900 176.200 48.200 ;
        RECT 168.600 47.300 169.900 47.600 ;
        RECT 167.000 47.100 167.800 47.200 ;
        RECT 162.300 46.800 167.800 47.100 ;
        RECT 161.400 46.400 161.800 46.500 ;
        RECT 159.900 46.100 161.800 46.400 ;
        RECT 159.900 46.000 160.300 46.100 ;
        RECT 160.700 45.700 161.100 45.800 ;
        RECT 159.000 45.400 161.100 45.700 ;
        RECT 153.400 44.400 153.800 45.200 ;
        RECT 154.200 45.100 154.600 45.200 ;
        RECT 154.200 44.800 154.900 45.100 ;
        RECT 155.200 44.800 156.200 45.200 ;
        RECT 154.600 44.200 154.900 44.800 ;
        RECT 154.600 43.800 155.000 44.200 ;
        RECT 155.300 41.100 155.700 44.800 ;
        RECT 159.000 41.100 159.400 45.400 ;
        RECT 162.300 45.200 162.600 46.800 ;
        RECT 165.900 46.700 166.300 46.800 ;
        RECT 166.700 46.200 167.100 46.300 ;
        RECT 168.700 46.200 169.100 46.600 ;
        RECT 164.600 45.900 167.100 46.200 ;
        RECT 164.600 45.800 165.000 45.900 ;
        RECT 168.600 45.800 169.100 46.200 ;
        RECT 169.600 46.500 169.900 47.300 ;
        RECT 170.400 47.200 170.700 47.900 ;
        RECT 171.900 47.700 173.700 47.900 ;
        RECT 172.200 47.200 172.600 47.400 ;
        RECT 174.200 47.200 174.500 47.900 ;
        RECT 170.200 46.800 170.700 47.200 ;
        RECT 171.800 46.900 172.600 47.200 ;
        RECT 173.300 47.100 174.600 47.200 ;
        RECT 175.000 47.100 175.400 47.200 ;
        RECT 171.800 46.800 172.200 46.900 ;
        RECT 173.300 46.800 175.400 47.100 ;
        RECT 169.600 46.100 170.100 46.500 ;
        RECT 165.400 45.500 168.200 45.600 ;
        RECT 165.300 45.400 168.200 45.500 ;
        RECT 161.400 44.900 162.600 45.200 ;
        RECT 163.300 45.300 168.200 45.400 ;
        RECT 163.300 45.100 165.700 45.300 ;
        RECT 161.400 44.400 161.700 44.900 ;
        RECT 161.000 44.000 161.700 44.400 ;
        RECT 162.500 44.500 162.900 44.600 ;
        RECT 163.300 44.500 163.600 45.100 ;
        RECT 162.500 44.200 163.600 44.500 ;
        RECT 163.900 44.500 166.600 44.800 ;
        RECT 163.900 44.400 164.300 44.500 ;
        RECT 166.200 44.400 166.600 44.500 ;
        RECT 163.100 43.700 163.500 43.800 ;
        RECT 164.500 43.700 164.900 43.800 ;
        RECT 161.400 43.100 161.800 43.500 ;
        RECT 163.100 43.400 164.900 43.700 ;
        RECT 163.500 43.100 163.800 43.400 ;
        RECT 166.200 43.100 166.600 43.500 ;
        RECT 161.100 41.100 161.700 43.100 ;
        RECT 163.400 41.100 163.800 43.100 ;
        RECT 165.600 42.800 166.600 43.100 ;
        RECT 165.600 41.100 166.000 42.800 ;
        RECT 167.800 41.100 168.200 45.300 ;
        RECT 169.600 45.100 169.900 46.100 ;
        RECT 170.400 45.100 170.700 46.800 ;
        RECT 172.600 45.800 173.000 46.600 ;
        RECT 173.300 45.100 173.600 46.800 ;
        RECT 175.800 46.100 176.200 47.900 ;
        RECT 177.400 47.700 177.800 49.900 ;
        RECT 179.500 49.200 180.100 49.900 ;
        RECT 179.500 48.900 180.200 49.200 ;
        RECT 181.800 48.900 182.200 49.900 ;
        RECT 184.000 49.200 184.400 49.900 ;
        RECT 184.000 48.900 185.000 49.200 ;
        RECT 179.800 48.500 180.200 48.900 ;
        RECT 181.900 48.600 182.200 48.900 ;
        RECT 181.900 48.300 183.300 48.600 ;
        RECT 182.900 48.200 183.300 48.300 ;
        RECT 183.800 48.200 184.200 48.600 ;
        RECT 184.600 48.500 185.000 48.900 ;
        RECT 178.900 47.700 179.300 47.800 ;
        RECT 176.600 47.100 177.000 47.600 ;
        RECT 177.400 47.400 179.300 47.700 ;
        RECT 177.400 47.100 177.800 47.400 ;
        RECT 180.900 47.100 181.300 47.200 ;
        RECT 183.800 47.100 184.100 48.200 ;
        RECT 186.200 47.500 186.600 49.900 ;
        RECT 187.000 47.500 187.400 49.900 ;
        RECT 189.200 49.200 189.600 49.900 ;
        RECT 188.600 48.900 189.600 49.200 ;
        RECT 191.400 48.900 191.800 49.900 ;
        RECT 193.500 49.200 194.100 49.900 ;
        RECT 193.400 48.900 194.100 49.200 ;
        RECT 188.600 48.500 189.000 48.900 ;
        RECT 191.400 48.600 191.700 48.900 ;
        RECT 189.400 48.200 189.800 48.600 ;
        RECT 190.300 48.300 191.700 48.600 ;
        RECT 193.400 48.500 193.800 48.900 ;
        RECT 190.300 48.200 190.700 48.300 ;
        RECT 185.400 47.100 186.200 47.200 ;
        RECT 176.600 46.800 177.800 47.100 ;
        RECT 174.200 45.800 176.200 46.100 ;
        RECT 174.200 45.200 174.500 45.800 ;
        RECT 174.200 45.100 174.600 45.200 ;
        RECT 168.600 44.800 169.900 45.100 ;
        RECT 168.600 41.100 169.000 44.800 ;
        RECT 170.200 44.600 170.700 45.100 ;
        RECT 173.100 44.800 173.600 45.100 ;
        RECT 173.900 44.800 174.600 45.100 ;
        RECT 170.200 41.100 170.600 44.600 ;
        RECT 173.100 41.100 173.500 44.800 ;
        RECT 173.900 44.200 174.200 44.800 ;
        RECT 175.000 44.400 175.400 45.200 ;
        RECT 173.800 43.800 174.200 44.200 ;
        RECT 175.800 41.100 176.200 45.800 ;
        RECT 177.400 45.700 177.800 46.800 ;
        RECT 180.700 46.800 186.200 47.100 ;
        RECT 187.400 47.100 188.200 47.200 ;
        RECT 189.500 47.100 189.800 48.200 ;
        RECT 194.300 47.700 194.700 47.800 ;
        RECT 195.800 47.700 196.200 49.900 ;
        RECT 194.300 47.400 196.200 47.700 ;
        RECT 196.600 47.500 197.000 49.900 ;
        RECT 198.800 49.200 199.200 49.900 ;
        RECT 198.200 48.900 199.200 49.200 ;
        RECT 201.000 48.900 201.400 49.900 ;
        RECT 203.100 49.200 203.700 49.900 ;
        RECT 203.000 48.900 203.700 49.200 ;
        RECT 198.200 48.500 198.600 48.900 ;
        RECT 201.000 48.600 201.300 48.900 ;
        RECT 199.000 48.200 199.400 48.600 ;
        RECT 199.900 48.300 201.300 48.600 ;
        RECT 203.000 48.500 203.400 48.900 ;
        RECT 199.900 48.200 200.300 48.300 ;
        RECT 192.300 47.100 192.700 47.200 ;
        RECT 187.400 46.800 192.900 47.100 ;
        RECT 179.800 46.400 180.200 46.500 ;
        RECT 178.300 46.100 180.200 46.400 ;
        RECT 178.300 46.000 178.700 46.100 ;
        RECT 179.100 45.700 179.500 45.800 ;
        RECT 177.400 45.400 179.500 45.700 ;
        RECT 177.400 41.100 177.800 45.400 ;
        RECT 180.700 45.200 181.000 46.800 ;
        RECT 184.300 46.700 184.700 46.800 ;
        RECT 188.900 46.700 189.300 46.800 ;
        RECT 185.100 46.200 185.500 46.300 ;
        RECT 183.000 45.900 185.500 46.200 ;
        RECT 188.100 46.200 188.500 46.300 ;
        RECT 188.100 46.100 190.600 46.200 ;
        RECT 191.800 46.100 192.200 46.200 ;
        RECT 188.100 45.900 192.200 46.100 ;
        RECT 183.000 45.800 183.400 45.900 ;
        RECT 190.200 45.800 192.200 45.900 ;
        RECT 183.800 45.500 186.600 45.600 ;
        RECT 183.700 45.400 186.600 45.500 ;
        RECT 179.800 44.900 181.000 45.200 ;
        RECT 181.700 45.300 186.600 45.400 ;
        RECT 181.700 45.100 184.100 45.300 ;
        RECT 179.800 44.400 180.100 44.900 ;
        RECT 179.400 44.000 180.100 44.400 ;
        RECT 180.900 44.500 181.300 44.600 ;
        RECT 181.700 44.500 182.000 45.100 ;
        RECT 180.900 44.200 182.000 44.500 ;
        RECT 182.300 44.500 185.000 44.800 ;
        RECT 182.300 44.400 182.700 44.500 ;
        RECT 184.600 44.400 185.000 44.500 ;
        RECT 181.500 43.700 181.900 43.800 ;
        RECT 182.900 43.700 183.300 43.800 ;
        RECT 179.800 43.100 180.200 43.500 ;
        RECT 181.500 43.400 183.300 43.700 ;
        RECT 181.900 43.100 182.200 43.400 ;
        RECT 184.600 43.100 185.000 43.500 ;
        RECT 179.500 41.100 180.100 43.100 ;
        RECT 181.800 41.100 182.200 43.100 ;
        RECT 184.000 42.800 185.000 43.100 ;
        RECT 184.000 41.100 184.400 42.800 ;
        RECT 186.200 41.100 186.600 45.300 ;
        RECT 187.000 45.500 189.800 45.600 ;
        RECT 187.000 45.400 189.900 45.500 ;
        RECT 187.000 45.300 191.900 45.400 ;
        RECT 187.000 41.100 187.400 45.300 ;
        RECT 189.500 45.100 191.900 45.300 ;
        RECT 188.600 44.500 191.300 44.800 ;
        RECT 188.600 44.400 189.000 44.500 ;
        RECT 190.900 44.400 191.300 44.500 ;
        RECT 191.600 44.500 191.900 45.100 ;
        RECT 192.600 45.200 192.900 46.800 ;
        RECT 193.400 46.400 193.800 46.500 ;
        RECT 193.400 46.100 195.300 46.400 ;
        RECT 194.900 46.000 195.300 46.100 ;
        RECT 194.100 45.700 194.500 45.800 ;
        RECT 195.800 45.700 196.200 47.400 ;
        RECT 199.100 47.200 199.400 48.200 ;
        RECT 202.200 48.100 202.600 48.200 ;
        RECT 205.400 48.100 205.800 49.900 ;
        RECT 207.000 48.900 207.400 49.900 ;
        RECT 206.200 48.100 206.600 48.600 ;
        RECT 207.100 48.100 207.400 48.900 ;
        RECT 210.300 48.200 210.700 48.600 ;
        RECT 210.200 48.100 210.600 48.200 ;
        RECT 202.200 47.800 204.200 48.100 ;
        RECT 205.400 47.800 206.600 48.100 ;
        RECT 207.000 47.800 210.600 48.100 ;
        RECT 211.000 47.800 211.400 49.900 ;
        RECT 203.800 47.700 204.300 47.800 ;
        RECT 205.400 47.700 205.800 47.800 ;
        RECT 203.800 47.400 205.800 47.700 ;
        RECT 197.000 47.100 197.800 47.200 ;
        RECT 199.000 47.100 199.400 47.200 ;
        RECT 201.900 47.100 202.300 47.200 ;
        RECT 197.000 46.800 202.500 47.100 ;
        RECT 198.500 46.700 198.900 46.800 ;
        RECT 197.700 46.200 198.100 46.300 ;
        RECT 197.700 45.900 200.200 46.200 ;
        RECT 199.800 45.800 200.200 45.900 ;
        RECT 194.100 45.400 196.200 45.700 ;
        RECT 192.600 44.900 193.800 45.200 ;
        RECT 192.300 44.500 192.700 44.600 ;
        RECT 191.600 44.200 192.700 44.500 ;
        RECT 193.500 44.400 193.800 44.900 ;
        RECT 193.500 44.000 194.200 44.400 ;
        RECT 190.300 43.700 190.700 43.800 ;
        RECT 191.700 43.700 192.100 43.800 ;
        RECT 188.600 43.100 189.000 43.500 ;
        RECT 190.300 43.400 192.100 43.700 ;
        RECT 191.400 43.100 191.700 43.400 ;
        RECT 193.400 43.100 193.800 43.500 ;
        RECT 188.600 42.800 189.600 43.100 ;
        RECT 189.200 41.100 189.600 42.800 ;
        RECT 191.400 41.100 191.800 43.100 ;
        RECT 193.500 41.100 194.100 43.100 ;
        RECT 195.800 41.100 196.200 45.400 ;
        RECT 196.600 45.500 199.400 45.600 ;
        RECT 196.600 45.400 199.500 45.500 ;
        RECT 196.600 45.300 201.500 45.400 ;
        RECT 196.600 41.100 197.000 45.300 ;
        RECT 199.100 45.100 201.500 45.300 ;
        RECT 198.200 44.500 200.900 44.800 ;
        RECT 198.200 44.400 198.600 44.500 ;
        RECT 200.500 44.400 200.900 44.500 ;
        RECT 201.200 44.500 201.500 45.100 ;
        RECT 202.200 45.200 202.500 46.800 ;
        RECT 203.000 46.400 203.400 46.500 ;
        RECT 203.000 46.100 204.900 46.400 ;
        RECT 204.500 46.000 204.900 46.100 ;
        RECT 203.700 45.700 204.100 45.800 ;
        RECT 205.400 45.700 205.800 47.400 ;
        RECT 207.100 47.200 207.400 47.800 ;
        RECT 207.000 46.800 207.400 47.200 ;
        RECT 203.700 45.400 205.800 45.700 ;
        RECT 202.200 44.900 203.400 45.200 ;
        RECT 201.900 44.500 202.300 44.600 ;
        RECT 201.200 44.200 202.300 44.500 ;
        RECT 203.100 44.400 203.400 44.900 ;
        RECT 203.100 44.000 203.800 44.400 ;
        RECT 199.900 43.700 200.300 43.800 ;
        RECT 201.300 43.700 201.700 43.800 ;
        RECT 198.200 43.100 198.600 43.500 ;
        RECT 199.900 43.400 201.700 43.700 ;
        RECT 201.000 43.100 201.300 43.400 ;
        RECT 203.000 43.100 203.400 43.500 ;
        RECT 198.200 42.800 199.200 43.100 ;
        RECT 198.800 41.100 199.200 42.800 ;
        RECT 201.000 41.100 201.400 43.100 ;
        RECT 203.100 41.100 203.700 43.100 ;
        RECT 205.400 41.100 205.800 45.400 ;
        RECT 207.100 45.100 207.400 46.800 ;
        RECT 207.800 45.400 208.200 46.200 ;
        RECT 210.200 46.100 210.600 46.200 ;
        RECT 211.100 46.100 211.400 47.800 ;
        RECT 213.400 48.500 213.800 49.500 ;
        RECT 215.500 49.200 215.900 49.500 ;
        RECT 218.500 49.200 218.900 49.900 ;
        RECT 215.500 48.800 216.200 49.200 ;
        RECT 218.200 48.800 218.900 49.200 ;
        RECT 213.400 47.400 213.700 48.500 ;
        RECT 215.500 48.000 215.900 48.800 ;
        RECT 218.500 48.200 218.900 48.800 ;
        RECT 220.600 48.500 221.000 49.500 ;
        RECT 222.700 49.200 223.100 49.500 ;
        RECT 222.700 48.800 223.400 49.200 ;
        RECT 215.500 47.700 216.300 48.000 ;
        RECT 218.500 47.900 219.400 48.200 ;
        RECT 215.900 47.500 216.300 47.700 ;
        RECT 211.800 46.400 212.200 47.200 ;
        RECT 213.400 47.100 215.500 47.400 ;
        RECT 215.000 46.900 215.500 47.100 ;
        RECT 216.000 47.200 216.300 47.500 ;
        RECT 212.600 46.100 213.000 46.200 ;
        RECT 210.200 45.800 211.400 46.100 ;
        RECT 212.200 45.800 213.000 46.100 ;
        RECT 213.400 45.800 213.800 46.600 ;
        RECT 214.200 45.800 214.600 46.600 ;
        RECT 215.000 46.500 215.700 46.900 ;
        RECT 216.000 46.800 217.000 47.200 ;
        RECT 210.300 45.100 210.600 45.800 ;
        RECT 212.200 45.600 212.600 45.800 ;
        RECT 215.000 45.500 215.300 46.500 ;
        RECT 213.400 45.200 215.300 45.500 ;
        RECT 207.000 44.700 207.900 45.100 ;
        RECT 207.500 41.100 207.900 44.700 ;
        RECT 210.200 41.100 210.600 45.100 ;
        RECT 211.000 44.800 213.000 45.100 ;
        RECT 211.000 41.100 211.400 44.800 ;
        RECT 212.600 41.100 213.000 44.800 ;
        RECT 213.400 43.500 213.700 45.200 ;
        RECT 216.000 44.900 216.300 46.800 ;
        RECT 216.600 45.400 217.000 46.200 ;
        RECT 217.400 46.100 217.800 46.200 ;
        RECT 217.400 45.800 218.500 46.100 ;
        RECT 215.500 44.600 216.300 44.900 ;
        RECT 218.200 45.200 218.500 45.800 ;
        RECT 213.400 41.500 213.800 43.500 ;
        RECT 215.500 41.100 215.900 44.600 ;
        RECT 218.200 44.400 218.600 45.200 ;
        RECT 219.000 41.100 219.400 47.900 ;
        RECT 219.800 46.800 220.200 47.600 ;
        RECT 220.600 47.400 220.900 48.500 ;
        RECT 222.700 48.000 223.100 48.800 ;
        RECT 225.400 48.500 225.800 49.500 ;
        RECT 227.500 49.200 227.900 49.500 ;
        RECT 227.000 48.800 227.900 49.200 ;
        RECT 222.700 47.700 223.500 48.000 ;
        RECT 223.100 47.500 223.500 47.700 ;
        RECT 220.600 47.100 222.700 47.400 ;
        RECT 222.200 46.900 222.700 47.100 ;
        RECT 223.200 47.200 223.500 47.500 ;
        RECT 225.400 47.400 225.700 48.500 ;
        RECT 227.500 48.000 227.900 48.800 ;
        RECT 230.200 48.000 230.600 49.900 ;
        RECT 231.800 48.000 232.200 49.900 ;
        RECT 227.500 47.700 228.300 48.000 ;
        RECT 230.200 47.900 232.200 48.000 ;
        RECT 232.600 47.900 233.000 49.900 ;
        RECT 233.700 48.200 234.100 49.900 ;
        RECT 237.100 49.200 237.500 49.900 ;
        RECT 237.100 48.800 237.800 49.200 ;
        RECT 237.100 48.200 237.500 48.800 ;
        RECT 233.700 47.900 234.600 48.200 ;
        RECT 230.300 47.700 232.100 47.900 ;
        RECT 227.900 47.500 228.300 47.700 ;
        RECT 220.600 45.800 221.000 46.600 ;
        RECT 221.400 45.800 221.800 46.600 ;
        RECT 222.200 46.500 222.900 46.900 ;
        RECT 223.200 46.800 224.200 47.200 ;
        RECT 225.400 47.100 227.500 47.400 ;
        RECT 227.000 46.900 227.500 47.100 ;
        RECT 228.000 47.200 228.300 47.500 ;
        RECT 230.600 47.200 231.000 47.400 ;
        RECT 232.600 47.200 232.900 47.900 ;
        RECT 222.200 45.500 222.500 46.500 ;
        RECT 220.600 45.200 222.500 45.500 ;
        RECT 220.600 43.500 220.900 45.200 ;
        RECT 223.200 44.900 223.500 46.800 ;
        RECT 223.800 45.400 224.200 46.200 ;
        RECT 225.400 45.800 225.800 46.600 ;
        RECT 226.200 45.800 226.600 46.600 ;
        RECT 227.000 46.500 227.700 46.900 ;
        RECT 228.000 46.800 229.000 47.200 ;
        RECT 230.200 46.900 231.000 47.200 ;
        RECT 231.700 47.100 233.000 47.200 ;
        RECT 233.400 47.100 233.800 47.200 ;
        RECT 230.200 46.800 230.600 46.900 ;
        RECT 231.700 46.800 233.800 47.100 ;
        RECT 227.000 45.500 227.300 46.500 ;
        RECT 222.700 44.600 223.500 44.900 ;
        RECT 225.400 45.200 227.300 45.500 ;
        RECT 220.600 41.500 221.000 43.500 ;
        RECT 222.700 41.100 223.100 44.600 ;
        RECT 225.400 43.500 225.700 45.200 ;
        RECT 228.000 44.900 228.300 46.800 ;
        RECT 228.600 45.400 229.000 46.200 ;
        RECT 231.000 45.800 231.400 46.600 ;
        RECT 231.700 45.100 232.000 46.800 ;
        RECT 234.200 46.100 234.600 47.900 ;
        RECT 236.600 47.900 237.500 48.200 ;
        RECT 235.000 46.800 235.400 47.600 ;
        RECT 235.800 46.800 236.200 47.600 ;
        RECT 232.600 45.800 234.600 46.100 ;
        RECT 232.600 45.200 232.900 45.800 ;
        RECT 232.600 45.100 233.000 45.200 ;
        RECT 227.500 44.600 228.300 44.900 ;
        RECT 231.500 44.800 232.000 45.100 ;
        RECT 232.300 44.800 233.000 45.100 ;
        RECT 225.400 41.500 225.800 43.500 ;
        RECT 227.500 41.100 227.900 44.600 ;
        RECT 231.500 41.100 231.900 44.800 ;
        RECT 232.300 44.200 232.600 44.800 ;
        RECT 233.400 44.400 233.800 45.200 ;
        RECT 232.200 43.800 232.600 44.200 ;
        RECT 234.200 41.100 234.600 45.800 ;
        RECT 236.600 41.100 237.000 47.900 ;
        RECT 238.200 47.700 238.600 49.900 ;
        RECT 240.300 49.200 240.900 49.900 ;
        RECT 240.300 48.900 241.000 49.200 ;
        RECT 242.600 48.900 243.000 49.900 ;
        RECT 244.800 49.200 245.200 49.900 ;
        RECT 244.800 48.900 245.800 49.200 ;
        RECT 240.600 48.500 241.000 48.900 ;
        RECT 242.700 48.600 243.000 48.900 ;
        RECT 242.700 48.300 244.100 48.600 ;
        RECT 243.700 48.200 244.100 48.300 ;
        RECT 244.600 48.200 245.000 48.600 ;
        RECT 245.400 48.500 245.800 48.900 ;
        RECT 239.700 47.700 240.100 47.800 ;
        RECT 238.200 47.400 240.100 47.700 ;
        RECT 238.200 45.700 238.600 47.400 ;
        RECT 241.700 47.100 242.100 47.200 ;
        RECT 244.600 47.100 244.900 48.200 ;
        RECT 247.000 47.500 247.400 49.900 ;
        RECT 248.600 48.800 249.000 49.900 ;
        RECT 248.600 47.200 248.900 48.800 ;
        RECT 249.400 47.800 249.800 48.600 ;
        RECT 250.200 47.500 250.600 49.900 ;
        RECT 252.400 49.200 252.800 49.900 ;
        RECT 251.800 48.900 252.800 49.200 ;
        RECT 254.600 48.900 255.000 49.900 ;
        RECT 256.700 49.200 257.300 49.900 ;
        RECT 256.600 48.900 257.300 49.200 ;
        RECT 251.800 48.500 252.200 48.900 ;
        RECT 254.600 48.600 254.900 48.900 ;
        RECT 252.600 47.800 253.000 48.600 ;
        RECT 253.500 48.300 254.900 48.600 ;
        RECT 256.600 48.500 257.000 48.900 ;
        RECT 253.500 48.200 253.900 48.300 ;
        RECT 246.200 47.100 247.000 47.200 ;
        RECT 241.500 46.800 247.000 47.100 ;
        RECT 248.600 46.800 249.000 47.200 ;
        RECT 250.600 47.100 251.400 47.200 ;
        RECT 252.700 47.100 253.000 47.800 ;
        RECT 257.500 47.700 257.900 47.800 ;
        RECT 259.000 47.700 259.400 49.900 ;
        RECT 261.100 48.200 261.500 49.900 ;
        RECT 257.500 47.400 259.400 47.700 ;
        RECT 260.600 47.900 261.500 48.200 ;
        RECT 262.200 48.000 262.600 49.900 ;
        RECT 263.800 48.000 264.200 49.900 ;
        RECT 262.200 47.900 264.200 48.000 ;
        RECT 264.600 47.900 265.000 49.900 ;
        RECT 255.500 47.100 255.900 47.200 ;
        RECT 250.600 46.800 256.100 47.100 ;
        RECT 240.600 46.400 241.000 46.500 ;
        RECT 239.100 46.100 241.000 46.400 ;
        RECT 241.500 46.200 241.800 46.800 ;
        RECT 245.100 46.700 245.500 46.800 ;
        RECT 245.900 46.200 246.300 46.300 ;
        RECT 239.100 46.000 239.500 46.100 ;
        RECT 241.400 45.800 241.800 46.200 ;
        RECT 243.800 45.900 246.300 46.200 ;
        RECT 243.800 45.800 244.200 45.900 ;
        RECT 239.900 45.700 240.300 45.800 ;
        RECT 238.200 45.400 240.300 45.700 ;
        RECT 237.400 44.400 237.800 45.200 ;
        RECT 238.200 41.100 238.600 45.400 ;
        RECT 241.500 45.200 241.800 45.800 ;
        RECT 244.600 45.500 247.400 45.600 ;
        RECT 244.500 45.400 247.400 45.500 ;
        RECT 247.800 45.400 248.200 46.200 ;
        RECT 240.600 44.900 241.800 45.200 ;
        RECT 242.500 45.300 247.400 45.400 ;
        RECT 242.500 45.100 244.900 45.300 ;
        RECT 240.600 44.400 240.900 44.900 ;
        RECT 240.200 44.000 240.900 44.400 ;
        RECT 241.700 44.500 242.100 44.600 ;
        RECT 242.500 44.500 242.800 45.100 ;
        RECT 241.700 44.200 242.800 44.500 ;
        RECT 243.100 44.500 245.800 44.800 ;
        RECT 243.100 44.400 243.500 44.500 ;
        RECT 245.400 44.400 245.800 44.500 ;
        RECT 242.300 43.700 242.700 43.800 ;
        RECT 243.700 43.700 244.100 43.800 ;
        RECT 240.600 43.100 241.000 43.500 ;
        RECT 242.300 43.400 244.100 43.700 ;
        RECT 242.700 43.100 243.000 43.400 ;
        RECT 245.400 43.100 245.800 43.500 ;
        RECT 240.300 41.100 240.900 43.100 ;
        RECT 242.600 41.100 243.000 43.100 ;
        RECT 244.800 42.800 245.800 43.100 ;
        RECT 244.800 41.100 245.200 42.800 ;
        RECT 247.000 41.100 247.400 45.300 ;
        RECT 248.600 45.100 248.900 46.800 ;
        RECT 252.100 46.700 252.500 46.800 ;
        RECT 251.300 46.200 251.700 46.300 ;
        RECT 252.600 46.200 253.000 46.300 ;
        RECT 251.300 45.900 253.800 46.200 ;
        RECT 253.400 45.800 253.800 45.900 ;
        RECT 250.200 45.500 253.000 45.600 ;
        RECT 250.200 45.400 253.100 45.500 ;
        RECT 250.200 45.300 255.100 45.400 ;
        RECT 248.100 44.700 249.000 45.100 ;
        RECT 248.100 41.100 248.500 44.700 ;
        RECT 250.200 41.100 250.600 45.300 ;
        RECT 252.700 45.100 255.100 45.300 ;
        RECT 251.800 44.500 254.500 44.800 ;
        RECT 251.800 44.400 252.200 44.500 ;
        RECT 254.100 44.400 254.500 44.500 ;
        RECT 254.800 44.500 255.100 45.100 ;
        RECT 255.800 45.200 256.100 46.800 ;
        RECT 256.600 46.400 257.000 46.500 ;
        RECT 256.600 46.100 258.500 46.400 ;
        RECT 258.100 46.000 258.500 46.100 ;
        RECT 257.300 45.700 257.700 45.800 ;
        RECT 259.000 45.700 259.400 47.400 ;
        RECT 259.800 46.800 260.200 47.600 ;
        RECT 257.300 45.400 259.400 45.700 ;
        RECT 255.800 44.900 257.000 45.200 ;
        RECT 255.500 44.500 255.900 44.600 ;
        RECT 254.800 44.200 255.900 44.500 ;
        RECT 256.700 44.400 257.000 44.900 ;
        RECT 256.700 44.000 257.400 44.400 ;
        RECT 253.500 43.700 253.900 43.800 ;
        RECT 254.900 43.700 255.300 43.800 ;
        RECT 251.800 43.100 252.200 43.500 ;
        RECT 253.500 43.400 255.300 43.700 ;
        RECT 254.600 43.100 254.900 43.400 ;
        RECT 256.600 43.100 257.000 43.500 ;
        RECT 251.800 42.800 252.800 43.100 ;
        RECT 252.400 41.100 252.800 42.800 ;
        RECT 254.600 41.100 255.000 43.100 ;
        RECT 256.700 41.100 257.300 43.100 ;
        RECT 259.000 41.100 259.400 45.400 ;
        RECT 259.800 44.100 260.200 44.200 ;
        RECT 260.600 44.100 261.000 47.900 ;
        RECT 262.300 47.700 264.100 47.900 ;
        RECT 262.600 47.200 263.000 47.400 ;
        RECT 264.600 47.200 264.900 47.900 ;
        RECT 261.400 47.100 261.800 47.200 ;
        RECT 262.200 47.100 263.000 47.200 ;
        RECT 261.400 46.900 263.000 47.100 ;
        RECT 261.400 46.800 262.600 46.900 ;
        RECT 263.700 46.800 265.000 47.200 ;
        RECT 263.000 46.100 263.400 46.600 ;
        RECT 261.400 45.800 263.400 46.100 ;
        RECT 261.400 45.200 261.700 45.800 ;
        RECT 261.400 44.400 261.800 45.200 ;
        RECT 263.700 45.100 264.000 46.800 ;
        RECT 264.600 45.100 265.000 45.200 ;
        RECT 263.500 44.800 264.000 45.100 ;
        RECT 264.300 44.800 265.000 45.100 ;
        RECT 259.800 43.800 261.000 44.100 ;
        RECT 260.600 41.100 261.000 43.800 ;
        RECT 263.500 42.200 263.900 44.800 ;
        RECT 264.300 44.200 264.600 44.800 ;
        RECT 264.200 43.800 264.600 44.200 ;
        RECT 263.000 41.800 263.900 42.200 ;
        RECT 263.500 41.100 263.900 41.800 ;
        RECT 0.600 36.200 1.000 39.900 ;
        RECT 2.200 36.200 2.600 39.900 ;
        RECT 0.600 35.900 2.600 36.200 ;
        RECT 3.000 35.900 3.400 39.900 ;
        RECT 4.100 36.300 4.500 39.900 ;
        RECT 6.200 37.500 6.600 39.500 ;
        RECT 8.300 39.200 8.700 39.900 ;
        RECT 8.300 38.800 9.000 39.200 ;
        RECT 4.100 35.900 5.000 36.300 ;
        RECT 1.000 35.200 1.400 35.400 ;
        RECT 3.000 35.200 3.300 35.900 ;
        RECT 0.600 34.900 1.400 35.200 ;
        RECT 2.200 34.900 3.400 35.200 ;
        RECT 0.600 34.800 1.000 34.900 ;
        RECT 1.400 33.800 1.800 34.600 ;
        RECT 2.200 34.100 2.500 34.900 ;
        RECT 3.000 34.800 3.400 34.900 ;
        RECT 3.800 34.800 4.200 35.600 ;
        RECT 4.600 34.200 4.900 35.900 ;
        RECT 6.200 35.800 6.500 37.500 ;
        RECT 8.300 36.400 8.700 38.800 ;
        RECT 8.300 36.100 9.100 36.400 ;
        RECT 6.200 35.500 8.100 35.800 ;
        RECT 6.200 34.400 6.600 35.200 ;
        RECT 7.000 34.400 7.400 35.200 ;
        RECT 7.800 34.500 8.100 35.500 ;
        RECT 3.000 34.100 3.400 34.200 ;
        RECT 2.200 33.800 3.400 34.100 ;
        RECT 4.600 33.800 5.000 34.200 ;
        RECT 7.800 34.100 8.500 34.500 ;
        RECT 8.800 34.200 9.100 36.100 ;
        RECT 9.400 35.100 9.800 35.600 ;
        RECT 11.000 35.100 11.400 35.200 ;
        RECT 9.400 34.800 11.400 35.100 ;
        RECT 7.800 33.900 8.300 34.100 ;
        RECT 2.200 33.100 2.500 33.800 ;
        RECT 3.000 33.100 3.400 33.200 ;
        RECT 4.600 33.100 4.900 33.800 ;
        RECT 6.200 33.600 8.300 33.900 ;
        RECT 8.800 33.800 9.800 34.200 ;
        RECT 2.200 31.100 2.600 33.100 ;
        RECT 3.000 32.800 4.900 33.100 ;
        RECT 2.900 32.400 3.300 32.800 ;
        RECT 4.600 32.100 4.900 32.800 ;
        RECT 5.400 32.400 5.800 33.200 ;
        RECT 6.200 32.500 6.500 33.600 ;
        RECT 8.800 33.500 9.100 33.800 ;
        RECT 8.700 33.300 9.100 33.500 ;
        RECT 8.300 33.000 9.100 33.300 ;
        RECT 4.600 31.100 5.000 32.100 ;
        RECT 6.200 31.500 6.600 32.500 ;
        RECT 8.300 31.500 8.700 33.000 ;
        RECT 11.000 32.400 11.400 33.200 ;
        RECT 11.800 31.100 12.200 39.900 ;
        RECT 12.600 35.600 13.000 39.900 ;
        RECT 14.700 37.900 15.300 39.900 ;
        RECT 17.000 37.900 17.400 39.900 ;
        RECT 19.200 38.200 19.600 39.900 ;
        RECT 19.200 37.900 20.200 38.200 ;
        RECT 15.000 37.500 15.400 37.900 ;
        RECT 17.100 37.600 17.400 37.900 ;
        RECT 16.700 37.300 18.500 37.600 ;
        RECT 19.800 37.500 20.200 37.900 ;
        RECT 16.700 37.200 17.100 37.300 ;
        RECT 18.100 37.200 18.500 37.300 ;
        RECT 14.600 36.600 15.300 37.000 ;
        RECT 15.000 36.100 15.300 36.600 ;
        RECT 16.100 36.500 17.200 36.800 ;
        RECT 16.100 36.400 16.500 36.500 ;
        RECT 15.000 35.800 16.200 36.100 ;
        RECT 12.600 35.300 14.700 35.600 ;
        RECT 12.600 33.600 13.000 35.300 ;
        RECT 14.300 35.200 14.700 35.300 ;
        RECT 13.500 34.900 13.900 35.000 ;
        RECT 13.500 34.600 15.400 34.900 ;
        RECT 15.000 34.500 15.400 34.600 ;
        RECT 15.900 34.200 16.200 35.800 ;
        RECT 16.900 35.900 17.200 36.500 ;
        RECT 17.500 36.500 17.900 36.600 ;
        RECT 19.800 36.500 20.200 36.600 ;
        RECT 17.500 36.200 20.200 36.500 ;
        RECT 16.900 35.700 19.300 35.900 ;
        RECT 21.400 35.700 21.800 39.900 ;
        RECT 24.100 36.400 24.500 39.900 ;
        RECT 26.200 37.500 26.600 39.500 ;
        RECT 16.900 35.600 21.800 35.700 ;
        RECT 23.700 36.100 24.500 36.400 ;
        RECT 18.900 35.500 21.800 35.600 ;
        RECT 19.000 35.400 21.800 35.500 ;
        RECT 18.200 35.100 18.600 35.200 ;
        RECT 18.200 34.800 20.700 35.100 ;
        RECT 23.000 34.800 23.400 35.600 ;
        RECT 19.000 34.700 19.400 34.800 ;
        RECT 20.300 34.700 20.700 34.800 ;
        RECT 19.500 34.200 19.900 34.300 ;
        RECT 23.700 34.200 24.000 36.100 ;
        RECT 26.300 35.800 26.600 37.500 ;
        RECT 28.300 36.200 28.700 39.900 ;
        RECT 29.000 36.800 29.400 37.200 ;
        RECT 29.100 36.200 29.400 36.800 ;
        RECT 28.300 35.900 28.800 36.200 ;
        RECT 29.100 35.900 29.800 36.200 ;
        RECT 24.700 35.500 26.600 35.800 ;
        RECT 24.700 34.500 25.000 35.500 ;
        RECT 15.900 33.900 21.400 34.200 ;
        RECT 16.100 33.800 16.500 33.900 ;
        RECT 12.600 33.300 14.500 33.600 ;
        RECT 12.600 31.100 13.000 33.300 ;
        RECT 14.100 33.200 14.500 33.300 ;
        RECT 19.000 32.800 19.300 33.900 ;
        RECT 20.600 33.800 21.400 33.900 ;
        RECT 22.200 34.100 22.600 34.200 ;
        RECT 23.000 34.100 24.000 34.200 ;
        RECT 24.300 34.100 25.000 34.500 ;
        RECT 25.400 34.400 25.800 35.200 ;
        RECT 26.200 35.100 26.600 35.200 ;
        RECT 27.000 35.100 27.400 35.200 ;
        RECT 26.200 34.800 27.400 35.100 ;
        RECT 26.200 34.400 26.600 34.800 ;
        RECT 27.800 34.400 28.200 35.200 ;
        RECT 28.500 34.200 28.800 35.900 ;
        RECT 29.400 35.800 29.800 35.900 ;
        RECT 30.200 35.800 30.600 36.600 ;
        RECT 29.400 35.100 29.700 35.800 ;
        RECT 31.000 35.100 31.400 39.900 ;
        RECT 33.900 36.200 34.300 39.900 ;
        RECT 34.600 36.800 35.000 37.200 ;
        RECT 34.700 36.200 35.000 36.800 ;
        RECT 33.900 35.900 34.400 36.200 ;
        RECT 34.700 35.900 35.400 36.200 ;
        RECT 29.400 34.800 31.400 35.100 ;
        RECT 22.200 33.800 24.000 34.100 ;
        RECT 23.700 33.500 24.000 33.800 ;
        RECT 24.500 33.900 25.000 34.100 ;
        RECT 27.000 34.100 27.400 34.200 ;
        RECT 24.500 33.600 26.600 33.900 ;
        RECT 27.000 33.800 27.800 34.100 ;
        RECT 28.500 33.800 29.800 34.200 ;
        RECT 27.400 33.600 27.800 33.800 ;
        RECT 18.100 32.700 18.500 32.800 ;
        RECT 15.000 32.100 15.400 32.500 ;
        RECT 17.100 32.400 18.500 32.700 ;
        RECT 19.000 32.400 19.400 32.800 ;
        RECT 17.100 32.100 17.400 32.400 ;
        RECT 19.800 32.100 20.200 32.500 ;
        RECT 14.700 31.800 15.400 32.100 ;
        RECT 14.700 31.100 15.300 31.800 ;
        RECT 17.000 31.100 17.400 32.100 ;
        RECT 19.200 31.800 20.200 32.100 ;
        RECT 19.200 31.100 19.600 31.800 ;
        RECT 21.400 31.100 21.800 33.500 ;
        RECT 23.700 33.300 24.100 33.500 ;
        RECT 23.700 33.000 24.500 33.300 ;
        RECT 24.100 31.500 24.500 33.000 ;
        RECT 26.300 32.500 26.600 33.600 ;
        RECT 27.100 33.100 28.900 33.300 ;
        RECT 29.400 33.100 29.700 33.800 ;
        RECT 31.000 33.100 31.400 34.800 ;
        RECT 33.400 34.400 33.800 35.200 ;
        RECT 34.100 34.200 34.400 35.900 ;
        RECT 35.000 35.800 35.400 35.900 ;
        RECT 35.800 35.800 36.200 36.600 ;
        RECT 35.000 35.100 35.300 35.800 ;
        RECT 36.600 35.100 37.000 39.900 ;
        RECT 38.200 37.500 38.600 39.500 ;
        RECT 40.300 39.200 40.700 39.900 ;
        RECT 40.300 38.800 41.000 39.200 ;
        RECT 38.200 35.800 38.500 37.500 ;
        RECT 40.300 36.400 40.700 38.800 ;
        RECT 40.300 36.100 41.100 36.400 ;
        RECT 38.200 35.500 40.100 35.800 ;
        RECT 35.000 34.800 37.000 35.100 ;
        RECT 31.800 33.400 32.200 34.200 ;
        RECT 32.600 34.100 33.000 34.200 ;
        RECT 32.600 33.800 33.400 34.100 ;
        RECT 34.100 33.800 35.400 34.200 ;
        RECT 33.000 33.600 33.400 33.800 ;
        RECT 32.700 33.100 34.500 33.300 ;
        RECT 35.000 33.100 35.300 33.800 ;
        RECT 36.600 33.100 37.000 34.800 ;
        RECT 38.200 34.400 38.600 35.200 ;
        RECT 39.000 34.400 39.400 35.200 ;
        RECT 39.800 34.500 40.100 35.500 ;
        RECT 37.400 33.400 37.800 34.200 ;
        RECT 39.800 34.100 40.500 34.500 ;
        RECT 40.800 34.200 41.100 36.100 ;
        RECT 43.300 36.300 43.700 39.900 ;
        RECT 43.300 35.900 44.200 36.300 ;
        RECT 41.400 34.800 41.800 35.600 ;
        RECT 42.200 35.100 42.600 35.200 ;
        RECT 43.000 35.100 43.400 35.600 ;
        RECT 42.200 34.800 43.400 35.100 ;
        RECT 43.800 34.200 44.100 35.900 ;
        RECT 45.400 35.700 45.800 39.900 ;
        RECT 47.600 38.200 48.000 39.900 ;
        RECT 47.000 37.900 48.000 38.200 ;
        RECT 49.800 37.900 50.200 39.900 ;
        RECT 51.900 37.900 52.500 39.900 ;
        RECT 47.000 37.500 47.400 37.900 ;
        RECT 49.800 37.600 50.100 37.900 ;
        RECT 48.700 37.300 50.500 37.600 ;
        RECT 51.800 37.500 52.200 37.900 ;
        RECT 48.700 37.200 49.100 37.300 ;
        RECT 50.100 37.200 50.500 37.300 ;
        RECT 47.000 36.500 47.400 36.600 ;
        RECT 49.300 36.500 49.700 36.600 ;
        RECT 47.000 36.200 49.700 36.500 ;
        RECT 50.000 36.500 51.100 36.800 ;
        RECT 50.000 35.900 50.300 36.500 ;
        RECT 50.700 36.400 51.100 36.500 ;
        RECT 51.900 36.600 52.600 37.000 ;
        RECT 51.900 36.100 52.200 36.600 ;
        RECT 47.900 35.700 50.300 35.900 ;
        RECT 45.400 35.600 50.300 35.700 ;
        RECT 51.000 35.800 52.200 36.100 ;
        RECT 45.400 35.500 48.300 35.600 ;
        RECT 45.400 35.400 48.200 35.500 ;
        RECT 48.600 35.100 49.000 35.200 ;
        RECT 46.500 34.800 49.000 35.100 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 51.000 35.100 51.300 35.800 ;
        RECT 54.200 35.600 54.600 39.900 ;
        RECT 58.500 36.400 58.900 39.900 ;
        RECT 60.600 37.500 61.000 39.500 ;
        RECT 58.100 36.100 58.900 36.400 ;
        RECT 52.500 35.300 54.600 35.600 ;
        RECT 52.500 35.200 52.900 35.300 ;
        RECT 50.200 34.800 51.300 35.100 ;
        RECT 54.200 35.100 54.600 35.300 ;
        RECT 57.400 35.100 57.800 35.600 ;
        RECT 53.300 34.900 53.700 35.000 ;
        RECT 46.500 34.700 46.900 34.800 ;
        RECT 47.800 34.700 48.200 34.800 ;
        RECT 47.300 34.200 47.700 34.300 ;
        RECT 51.000 34.200 51.300 34.800 ;
        RECT 51.800 34.600 53.700 34.900 ;
        RECT 54.200 34.800 57.800 35.100 ;
        RECT 51.800 34.500 52.200 34.600 ;
        RECT 39.800 33.900 40.300 34.100 ;
        RECT 38.200 33.600 40.300 33.900 ;
        RECT 40.800 33.800 41.800 34.200 ;
        RECT 43.800 33.800 44.200 34.200 ;
        RECT 45.800 33.900 51.300 34.200 ;
        RECT 45.800 33.800 46.600 33.900 ;
        RECT 26.200 31.500 26.600 32.500 ;
        RECT 27.000 33.000 29.000 33.100 ;
        RECT 27.000 31.100 27.400 33.000 ;
        RECT 28.600 31.100 29.000 33.000 ;
        RECT 29.400 31.100 29.800 33.100 ;
        RECT 30.500 32.800 31.400 33.100 ;
        RECT 32.600 33.000 34.600 33.100 ;
        RECT 30.500 31.100 30.900 32.800 ;
        RECT 32.600 31.100 33.000 33.000 ;
        RECT 34.200 31.100 34.600 33.000 ;
        RECT 35.000 31.100 35.400 33.100 ;
        RECT 36.100 32.800 37.000 33.100 ;
        RECT 36.100 31.100 36.500 32.800 ;
        RECT 38.200 32.500 38.500 33.600 ;
        RECT 40.800 33.500 41.100 33.800 ;
        RECT 40.700 33.300 41.100 33.500 ;
        RECT 40.300 33.000 41.100 33.300 ;
        RECT 38.200 31.500 38.600 32.500 ;
        RECT 40.300 31.500 40.700 33.000 ;
        RECT 43.800 32.200 44.100 33.800 ;
        RECT 44.600 32.400 45.000 33.200 ;
        RECT 43.800 31.100 44.200 32.200 ;
        RECT 45.400 31.100 45.800 33.500 ;
        RECT 47.900 32.800 48.200 33.900 ;
        RECT 50.700 33.800 51.100 33.900 ;
        RECT 54.200 33.600 54.600 34.800 ;
        RECT 58.100 34.200 58.400 36.100 ;
        RECT 60.700 35.800 61.000 37.500 ;
        RECT 59.100 35.500 61.000 35.800 ;
        RECT 59.100 34.500 59.400 35.500 ;
        RECT 57.400 33.800 58.400 34.200 ;
        RECT 58.700 34.100 59.400 34.500 ;
        RECT 59.800 34.400 60.200 35.200 ;
        RECT 60.600 34.400 61.000 35.200 ;
        RECT 52.700 33.300 54.600 33.600 ;
        RECT 52.700 33.200 53.100 33.300 ;
        RECT 47.000 32.100 47.400 32.500 ;
        RECT 47.800 32.400 48.200 32.800 ;
        RECT 48.700 32.700 49.100 32.800 ;
        RECT 48.700 32.400 50.100 32.700 ;
        RECT 49.800 32.100 50.100 32.400 ;
        RECT 51.800 32.100 52.200 32.500 ;
        RECT 47.000 31.800 48.000 32.100 ;
        RECT 47.600 31.100 48.000 31.800 ;
        RECT 49.800 31.100 50.200 32.100 ;
        RECT 51.800 31.800 52.500 32.100 ;
        RECT 51.900 31.100 52.500 31.800 ;
        RECT 54.200 31.100 54.600 33.300 ;
        RECT 58.100 33.500 58.400 33.800 ;
        RECT 58.900 33.900 59.400 34.100 ;
        RECT 58.900 33.600 61.000 33.900 ;
        RECT 58.100 33.300 58.500 33.500 ;
        RECT 58.100 33.000 58.900 33.300 ;
        RECT 58.500 32.200 58.900 33.000 ;
        RECT 60.700 32.500 61.000 33.600 ;
        RECT 61.400 33.400 61.800 34.200 ;
        RECT 62.200 33.100 62.600 39.900 ;
        RECT 63.800 37.500 64.200 39.500 ;
        RECT 65.900 39.200 66.300 39.900 ;
        RECT 65.900 38.800 66.600 39.200 ;
        RECT 63.000 35.800 63.400 36.600 ;
        RECT 63.800 35.800 64.100 37.500 ;
        RECT 65.900 36.400 66.300 38.800 ;
        RECT 65.900 36.100 66.700 36.400 ;
        RECT 63.800 35.500 65.700 35.800 ;
        RECT 63.800 34.400 64.200 35.200 ;
        RECT 64.600 34.400 65.000 35.200 ;
        RECT 65.400 34.500 65.700 35.500 ;
        RECT 65.400 34.100 66.100 34.500 ;
        RECT 66.400 34.200 66.700 36.100 ;
        RECT 69.900 36.200 70.300 39.900 ;
        RECT 70.600 36.800 71.000 37.200 ;
        RECT 70.700 36.200 71.000 36.800 ;
        RECT 69.900 35.900 70.400 36.200 ;
        RECT 70.700 35.900 71.400 36.200 ;
        RECT 67.000 34.800 67.400 35.600 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 69.400 35.100 69.800 35.200 ;
        RECT 67.800 34.800 69.800 35.100 ;
        RECT 69.400 34.400 69.800 34.800 ;
        RECT 70.100 34.200 70.400 35.900 ;
        RECT 71.000 35.800 71.400 35.900 ;
        RECT 71.800 35.800 72.200 36.600 ;
        RECT 71.000 35.100 71.300 35.800 ;
        RECT 72.600 35.100 73.000 39.900 ;
        RECT 74.200 35.700 74.600 39.900 ;
        RECT 76.400 38.200 76.800 39.900 ;
        RECT 75.800 37.900 76.800 38.200 ;
        RECT 78.600 37.900 79.000 39.900 ;
        RECT 80.700 37.900 81.300 39.900 ;
        RECT 75.800 37.500 76.200 37.900 ;
        RECT 78.600 37.600 78.900 37.900 ;
        RECT 77.500 37.300 79.300 37.600 ;
        RECT 80.600 37.500 81.000 37.900 ;
        RECT 77.500 37.200 77.900 37.300 ;
        RECT 78.900 37.200 79.300 37.300 ;
        RECT 75.800 36.500 76.200 36.600 ;
        RECT 78.100 36.500 78.500 36.600 ;
        RECT 75.800 36.200 78.500 36.500 ;
        RECT 78.800 36.500 79.900 36.800 ;
        RECT 78.800 35.900 79.100 36.500 ;
        RECT 79.500 36.400 79.900 36.500 ;
        RECT 80.700 36.600 81.400 37.000 ;
        RECT 80.700 36.100 81.000 36.600 ;
        RECT 76.700 35.700 79.100 35.900 ;
        RECT 74.200 35.600 79.100 35.700 ;
        RECT 79.800 35.800 81.000 36.100 ;
        RECT 74.200 35.500 77.100 35.600 ;
        RECT 74.200 35.400 77.000 35.500 ;
        RECT 79.800 35.200 80.100 35.800 ;
        RECT 83.000 35.600 83.400 39.900 ;
        RECT 81.300 35.300 83.400 35.600 ;
        RECT 83.800 37.500 84.200 39.500 ;
        RECT 85.900 39.200 86.300 39.900 ;
        RECT 90.500 39.200 90.900 39.900 ;
        RECT 85.900 38.800 86.600 39.200 ;
        RECT 90.500 38.800 91.400 39.200 ;
        RECT 83.800 35.800 84.100 37.500 ;
        RECT 85.900 36.400 86.300 38.800 ;
        RECT 90.500 36.400 90.900 38.800 ;
        RECT 92.600 37.500 93.000 39.500 ;
        RECT 85.900 36.100 86.700 36.400 ;
        RECT 83.800 35.500 85.700 35.800 ;
        RECT 81.300 35.200 81.700 35.300 ;
        RECT 77.400 35.100 77.800 35.200 ;
        RECT 71.000 34.800 73.000 35.100 ;
        RECT 65.400 33.900 65.900 34.100 ;
        RECT 63.800 33.600 65.900 33.900 ;
        RECT 66.400 33.800 67.400 34.200 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 70.100 34.100 71.400 34.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 68.600 33.800 69.400 34.100 ;
        RECT 70.100 33.800 72.200 34.100 ;
        RECT 62.200 32.800 63.100 33.100 ;
        RECT 58.500 31.800 59.400 32.200 ;
        RECT 58.500 31.500 58.900 31.800 ;
        RECT 60.600 31.500 61.000 32.500 ;
        RECT 62.700 32.200 63.100 32.800 ;
        RECT 63.800 32.500 64.100 33.600 ;
        RECT 66.400 33.500 66.700 33.800 ;
        RECT 69.000 33.600 69.400 33.800 ;
        RECT 66.300 33.300 66.700 33.500 ;
        RECT 65.900 33.000 66.700 33.300 ;
        RECT 68.700 33.100 70.500 33.300 ;
        RECT 71.000 33.100 71.300 33.800 ;
        RECT 72.600 33.100 73.000 34.800 ;
        RECT 75.300 34.800 77.800 35.100 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 82.100 34.900 82.500 35.000 ;
        RECT 75.300 34.700 75.700 34.800 ;
        RECT 76.600 34.700 77.000 34.800 ;
        RECT 76.100 34.200 76.500 34.300 ;
        RECT 79.800 34.200 80.100 34.800 ;
        RECT 80.600 34.600 82.500 34.900 ;
        RECT 80.600 34.500 81.000 34.600 ;
        RECT 73.400 33.400 73.800 34.200 ;
        RECT 74.600 33.900 80.100 34.200 ;
        RECT 74.600 33.800 75.400 33.900 ;
        RECT 68.600 33.000 70.600 33.100 ;
        RECT 62.700 31.800 63.400 32.200 ;
        RECT 62.700 31.100 63.100 31.800 ;
        RECT 63.800 31.500 64.200 32.500 ;
        RECT 65.900 31.500 66.300 33.000 ;
        RECT 68.600 31.100 69.000 33.000 ;
        RECT 70.200 31.100 70.600 33.000 ;
        RECT 71.000 31.100 71.400 33.100 ;
        RECT 72.100 32.800 73.000 33.100 ;
        RECT 72.100 31.100 72.500 32.800 ;
        RECT 74.200 31.100 74.600 33.500 ;
        RECT 76.700 32.800 77.000 33.900 ;
        RECT 78.200 33.800 78.600 33.900 ;
        RECT 79.500 33.800 79.900 33.900 ;
        RECT 83.000 33.600 83.400 35.300 ;
        RECT 83.800 34.400 84.200 35.200 ;
        RECT 84.600 34.400 85.000 35.200 ;
        RECT 85.400 34.500 85.700 35.500 ;
        RECT 85.400 34.100 86.100 34.500 ;
        RECT 86.400 34.200 86.700 36.100 ;
        RECT 90.100 36.100 90.900 36.400 ;
        RECT 87.000 34.800 87.400 35.600 ;
        RECT 88.600 35.100 89.000 35.200 ;
        RECT 89.400 35.100 89.800 35.600 ;
        RECT 88.600 34.800 89.800 35.100 ;
        RECT 90.100 34.200 90.400 36.100 ;
        RECT 92.700 35.800 93.000 37.500 ;
        RECT 91.100 35.500 93.000 35.800 ;
        RECT 93.400 35.700 93.800 39.900 ;
        RECT 95.600 38.200 96.000 39.900 ;
        RECT 95.000 37.900 96.000 38.200 ;
        RECT 97.800 37.900 98.200 39.900 ;
        RECT 99.900 37.900 100.500 39.900 ;
        RECT 95.000 37.500 95.400 37.900 ;
        RECT 97.800 37.600 98.100 37.900 ;
        RECT 96.700 37.300 98.500 37.600 ;
        RECT 99.800 37.500 100.200 37.900 ;
        RECT 96.700 37.200 97.100 37.300 ;
        RECT 98.100 37.200 98.500 37.300 ;
        RECT 95.000 36.500 95.400 36.600 ;
        RECT 97.300 36.500 97.700 36.600 ;
        RECT 95.000 36.200 97.700 36.500 ;
        RECT 98.000 36.500 99.100 36.800 ;
        RECT 98.000 35.900 98.300 36.500 ;
        RECT 98.700 36.400 99.100 36.500 ;
        RECT 99.900 36.600 100.600 37.000 ;
        RECT 99.900 36.100 100.200 36.600 ;
        RECT 95.900 35.700 98.300 35.900 ;
        RECT 93.400 35.600 98.300 35.700 ;
        RECT 99.000 35.800 100.200 36.100 ;
        RECT 93.400 35.500 96.300 35.600 ;
        RECT 91.100 34.500 91.400 35.500 ;
        RECT 93.400 35.400 96.200 35.500 ;
        RECT 85.400 33.900 85.900 34.100 ;
        RECT 81.500 33.300 83.400 33.600 ;
        RECT 81.500 33.200 81.900 33.300 ;
        RECT 75.800 32.100 76.200 32.500 ;
        RECT 76.600 32.400 77.000 32.800 ;
        RECT 77.500 32.700 77.900 32.800 ;
        RECT 77.500 32.400 78.900 32.700 ;
        RECT 78.600 32.100 78.900 32.400 ;
        RECT 80.600 32.100 81.000 32.500 ;
        RECT 75.800 31.800 76.800 32.100 ;
        RECT 76.400 31.100 76.800 31.800 ;
        RECT 78.600 31.100 79.000 32.100 ;
        RECT 80.600 31.800 81.300 32.100 ;
        RECT 80.700 31.100 81.300 31.800 ;
        RECT 83.000 31.100 83.400 33.300 ;
        RECT 83.800 33.600 85.900 33.900 ;
        RECT 86.400 33.800 87.400 34.200 ;
        RECT 89.400 33.800 90.400 34.200 ;
        RECT 90.700 34.100 91.400 34.500 ;
        RECT 91.800 34.400 92.200 35.200 ;
        RECT 92.600 34.400 93.000 35.200 ;
        RECT 96.600 35.100 97.000 35.200 ;
        RECT 97.400 35.100 97.800 35.200 ;
        RECT 94.500 34.800 97.800 35.100 ;
        RECT 94.500 34.700 94.900 34.800 ;
        RECT 95.300 34.200 95.700 34.300 ;
        RECT 99.000 34.200 99.300 35.800 ;
        RECT 102.200 35.600 102.600 39.900 ;
        RECT 100.500 35.300 102.600 35.600 ;
        RECT 100.500 35.200 100.900 35.300 ;
        RECT 101.300 34.900 101.700 35.000 ;
        RECT 99.800 34.600 101.700 34.900 ;
        RECT 99.800 34.500 100.200 34.600 ;
        RECT 83.800 32.500 84.100 33.600 ;
        RECT 86.400 33.500 86.700 33.800 ;
        RECT 86.300 33.300 86.700 33.500 ;
        RECT 85.900 33.000 86.700 33.300 ;
        RECT 90.100 33.500 90.400 33.800 ;
        RECT 90.900 33.900 91.400 34.100 ;
        RECT 93.800 33.900 99.300 34.200 ;
        RECT 90.900 33.600 93.000 33.900 ;
        RECT 93.800 33.800 94.600 33.900 ;
        RECT 90.100 33.300 90.500 33.500 ;
        RECT 90.100 33.000 90.900 33.300 ;
        RECT 83.800 31.500 84.200 32.500 ;
        RECT 85.900 31.500 86.300 33.000 ;
        RECT 90.500 31.500 90.900 33.000 ;
        RECT 92.700 32.500 93.000 33.600 ;
        RECT 92.600 31.500 93.000 32.500 ;
        RECT 93.400 31.100 93.800 33.500 ;
        RECT 95.900 32.800 96.200 33.900 ;
        RECT 96.600 33.800 97.000 33.900 ;
        RECT 98.700 33.800 99.100 33.900 ;
        RECT 102.200 33.600 102.600 35.300 ;
        RECT 103.800 35.100 104.200 39.900 ;
        RECT 108.100 36.400 108.500 39.900 ;
        RECT 110.200 37.500 110.600 39.500 ;
        RECT 107.700 36.100 108.500 36.400 ;
        RECT 107.000 35.100 107.400 35.600 ;
        RECT 103.800 34.800 107.400 35.100 ;
        RECT 100.700 33.300 102.600 33.600 ;
        RECT 100.700 33.200 101.100 33.300 ;
        RECT 102.200 33.100 102.600 33.300 ;
        RECT 103.000 33.800 103.400 34.200 ;
        RECT 103.000 33.200 103.300 33.800 ;
        RECT 103.000 33.100 103.400 33.200 ;
        RECT 102.200 32.800 103.400 33.100 ;
        RECT 95.000 32.100 95.400 32.500 ;
        RECT 95.800 32.400 96.200 32.800 ;
        RECT 96.700 32.700 97.100 32.800 ;
        RECT 96.700 32.400 98.100 32.700 ;
        RECT 97.800 32.100 98.100 32.400 ;
        RECT 99.800 32.100 100.200 32.500 ;
        RECT 95.000 31.800 96.000 32.100 ;
        RECT 95.600 31.100 96.000 31.800 ;
        RECT 97.800 31.100 98.200 32.100 ;
        RECT 99.800 31.800 100.500 32.100 ;
        RECT 99.900 31.100 100.500 31.800 ;
        RECT 102.200 31.100 102.600 32.800 ;
        RECT 103.000 32.400 103.400 32.800 ;
        RECT 103.800 31.100 104.200 34.800 ;
        RECT 107.700 34.200 108.000 36.100 ;
        RECT 110.300 35.800 110.600 37.500 ;
        RECT 108.700 35.500 110.600 35.800 ;
        RECT 111.800 35.600 112.200 39.900 ;
        RECT 113.400 35.600 113.800 39.900 ;
        RECT 115.000 35.600 115.400 39.900 ;
        RECT 116.600 35.600 117.000 39.900 ;
        RECT 119.000 35.600 119.400 39.900 ;
        RECT 120.600 35.600 121.000 39.900 ;
        RECT 122.200 35.600 122.600 39.900 ;
        RECT 123.800 35.600 124.200 39.900 ;
        RECT 108.700 34.500 109.000 35.500 ;
        RECT 111.000 35.200 112.200 35.600 ;
        RECT 112.700 35.200 113.800 35.600 ;
        RECT 114.300 35.200 115.400 35.600 ;
        RECT 116.100 35.200 117.000 35.600 ;
        RECT 118.200 35.200 119.400 35.600 ;
        RECT 119.900 35.200 121.000 35.600 ;
        RECT 121.500 35.200 122.600 35.600 ;
        RECT 123.300 35.200 124.200 35.600 ;
        RECT 125.400 37.500 125.800 39.500 ;
        RECT 127.500 39.200 127.900 39.900 ;
        RECT 127.500 38.800 128.200 39.200 ;
        RECT 125.400 35.800 125.700 37.500 ;
        RECT 127.500 36.400 127.900 38.800 ;
        RECT 127.500 36.100 128.300 36.400 ;
        RECT 125.400 35.500 127.300 35.800 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 107.000 34.100 108.000 34.200 ;
        RECT 108.300 34.100 109.000 34.500 ;
        RECT 109.400 34.400 109.800 35.200 ;
        RECT 110.200 34.400 110.600 35.200 ;
        RECT 105.400 33.800 108.000 34.100 ;
        RECT 107.700 33.500 108.000 33.800 ;
        RECT 108.500 33.900 109.000 34.100 ;
        RECT 108.500 33.600 110.600 33.900 ;
        RECT 107.700 33.300 108.100 33.500 ;
        RECT 107.700 33.000 108.500 33.300 ;
        RECT 108.100 31.500 108.500 33.000 ;
        RECT 110.300 32.500 110.600 33.600 ;
        RECT 111.000 33.800 111.400 35.200 ;
        RECT 112.700 34.500 113.100 35.200 ;
        RECT 114.300 34.500 114.700 35.200 ;
        RECT 116.100 34.500 116.500 35.200 ;
        RECT 111.800 34.100 113.100 34.500 ;
        RECT 113.500 34.100 114.700 34.500 ;
        RECT 115.200 34.100 116.500 34.500 ;
        RECT 116.900 34.100 117.800 34.500 ;
        RECT 112.700 33.800 113.100 34.100 ;
        RECT 114.300 33.800 114.700 34.100 ;
        RECT 116.100 33.800 116.500 34.100 ;
        RECT 117.400 33.800 117.800 34.100 ;
        RECT 118.200 33.800 118.600 35.200 ;
        RECT 119.900 34.500 120.300 35.200 ;
        RECT 121.500 34.500 121.900 35.200 ;
        RECT 123.300 34.500 123.700 35.200 ;
        RECT 119.000 34.100 120.300 34.500 ;
        RECT 120.700 34.100 121.900 34.500 ;
        RECT 122.400 34.100 123.700 34.500 ;
        RECT 124.100 34.100 125.000 34.500 ;
        RECT 125.400 34.400 125.800 35.200 ;
        RECT 126.200 34.400 126.600 35.200 ;
        RECT 127.000 34.500 127.300 35.500 ;
        RECT 119.900 33.800 120.300 34.100 ;
        RECT 121.500 33.800 121.900 34.100 ;
        RECT 123.300 33.800 123.700 34.100 ;
        RECT 124.600 33.800 125.000 34.100 ;
        RECT 127.000 34.100 127.700 34.500 ;
        RECT 128.000 34.200 128.300 36.100 ;
        RECT 130.200 36.200 130.600 39.900 ;
        RECT 131.800 36.400 132.200 39.900 ;
        RECT 133.400 37.500 133.800 39.500 ;
        RECT 135.500 39.200 135.900 39.900 ;
        RECT 135.500 38.800 136.200 39.200 ;
        RECT 130.200 35.900 131.500 36.200 ;
        RECT 131.800 35.900 132.300 36.400 ;
        RECT 128.600 34.800 129.000 35.600 ;
        RECT 130.200 34.800 130.700 35.200 ;
        RECT 130.300 34.400 130.700 34.800 ;
        RECT 131.200 34.900 131.500 35.900 ;
        RECT 131.200 34.500 131.700 34.900 ;
        RECT 127.000 33.900 127.500 34.100 ;
        RECT 111.000 33.400 112.200 33.800 ;
        RECT 112.700 33.400 113.800 33.800 ;
        RECT 114.300 33.400 115.400 33.800 ;
        RECT 116.100 33.400 117.000 33.800 ;
        RECT 118.200 33.400 119.400 33.800 ;
        RECT 119.900 33.400 121.000 33.800 ;
        RECT 121.500 33.400 122.600 33.800 ;
        RECT 123.300 33.400 124.200 33.800 ;
        RECT 110.200 31.500 110.600 32.500 ;
        RECT 111.800 31.100 112.200 33.400 ;
        RECT 113.400 31.100 113.800 33.400 ;
        RECT 115.000 31.100 115.400 33.400 ;
        RECT 116.600 31.100 117.000 33.400 ;
        RECT 119.000 31.100 119.400 33.400 ;
        RECT 120.600 31.100 121.000 33.400 ;
        RECT 122.200 31.100 122.600 33.400 ;
        RECT 123.800 31.100 124.200 33.400 ;
        RECT 125.400 33.600 127.500 33.900 ;
        RECT 128.000 33.800 129.000 34.200 ;
        RECT 125.400 32.500 125.700 33.600 ;
        RECT 128.000 33.500 128.300 33.800 ;
        RECT 131.200 33.700 131.500 34.500 ;
        RECT 132.000 34.200 132.300 35.900 ;
        RECT 133.400 35.800 133.700 37.500 ;
        RECT 135.500 36.400 135.900 38.800 ;
        RECT 135.500 36.100 136.300 36.400 ;
        RECT 139.500 36.300 139.900 39.900 ;
        RECT 133.400 35.500 135.300 35.800 ;
        RECT 133.400 34.400 133.800 35.200 ;
        RECT 134.200 34.400 134.600 35.200 ;
        RECT 135.000 34.500 135.300 35.500 ;
        RECT 131.800 33.800 132.300 34.200 ;
        RECT 135.000 34.100 135.700 34.500 ;
        RECT 136.000 34.200 136.300 36.100 ;
        RECT 139.000 35.900 139.900 36.300 ;
        RECT 140.600 35.900 141.000 39.900 ;
        RECT 141.400 36.200 141.800 39.900 ;
        RECT 143.000 36.200 143.400 39.900 ;
        RECT 141.400 35.900 143.400 36.200 ;
        RECT 136.600 35.100 137.000 35.600 ;
        RECT 138.200 35.100 138.600 35.200 ;
        RECT 136.600 34.800 138.600 35.100 ;
        RECT 139.100 34.200 139.400 35.900 ;
        RECT 139.800 34.800 140.200 35.600 ;
        RECT 140.700 35.200 141.000 35.900 ;
        RECT 143.800 35.700 144.200 39.900 ;
        RECT 146.000 38.200 146.400 39.900 ;
        RECT 145.400 37.900 146.400 38.200 ;
        RECT 148.200 37.900 148.600 39.900 ;
        RECT 150.300 37.900 150.900 39.900 ;
        RECT 145.400 37.500 145.800 37.900 ;
        RECT 148.200 37.600 148.500 37.900 ;
        RECT 147.100 37.300 148.900 37.600 ;
        RECT 150.200 37.500 150.600 37.900 ;
        RECT 147.100 37.200 147.500 37.300 ;
        RECT 148.500 37.200 148.900 37.300 ;
        RECT 145.400 36.500 145.800 36.600 ;
        RECT 147.700 36.500 148.100 36.600 ;
        RECT 145.400 36.200 148.100 36.500 ;
        RECT 148.400 36.500 149.500 36.800 ;
        RECT 148.400 35.900 148.700 36.500 ;
        RECT 149.100 36.400 149.500 36.500 ;
        RECT 150.300 36.600 151.000 37.000 ;
        RECT 150.300 36.100 150.600 36.600 ;
        RECT 146.300 35.700 148.700 35.900 ;
        RECT 143.800 35.600 148.700 35.700 ;
        RECT 149.400 35.800 150.600 36.100 ;
        RECT 143.800 35.500 146.700 35.600 ;
        RECT 143.800 35.400 146.600 35.500 ;
        RECT 142.600 35.200 143.000 35.400 ;
        RECT 149.400 35.200 149.700 35.800 ;
        RECT 152.600 35.600 153.000 39.900 ;
        RECT 150.900 35.300 153.000 35.600 ;
        RECT 153.400 35.600 153.800 39.900 ;
        RECT 155.500 39.200 155.900 39.900 ;
        RECT 155.500 38.800 156.200 39.200 ;
        RECT 155.500 36.200 155.900 38.800 ;
        RECT 155.500 35.900 156.200 36.200 ;
        RECT 153.400 35.400 155.400 35.600 ;
        RECT 153.400 35.300 155.500 35.400 ;
        RECT 150.900 35.200 151.300 35.300 ;
        RECT 140.600 34.900 141.800 35.200 ;
        RECT 142.600 34.900 143.400 35.200 ;
        RECT 147.000 35.100 147.400 35.200 ;
        RECT 140.600 34.800 141.000 34.900 ;
        RECT 135.000 33.900 135.500 34.100 ;
        RECT 127.900 33.300 128.300 33.500 ;
        RECT 127.500 33.000 128.300 33.300 ;
        RECT 130.200 33.400 131.500 33.700 ;
        RECT 125.400 31.500 125.800 32.500 ;
        RECT 127.500 31.500 127.900 33.000 ;
        RECT 130.200 31.100 130.600 33.400 ;
        RECT 132.000 33.100 132.300 33.800 ;
        RECT 131.800 32.800 132.300 33.100 ;
        RECT 133.400 33.600 135.500 33.900 ;
        RECT 136.000 33.800 137.000 34.200 ;
        RECT 139.000 33.800 139.400 34.200 ;
        RECT 131.800 31.100 132.200 32.800 ;
        RECT 133.400 32.500 133.700 33.600 ;
        RECT 136.000 33.500 136.300 33.800 ;
        RECT 135.900 33.300 136.300 33.500 ;
        RECT 135.500 33.000 136.300 33.300 ;
        RECT 133.400 31.500 133.800 32.500 ;
        RECT 135.500 31.500 135.900 33.000 ;
        RECT 138.200 32.400 138.600 33.200 ;
        RECT 139.100 33.100 139.400 33.800 ;
        RECT 140.600 33.100 141.000 33.200 ;
        RECT 141.500 33.100 141.800 34.900 ;
        RECT 143.000 34.800 143.400 34.900 ;
        RECT 144.900 34.800 147.400 35.100 ;
        RECT 149.400 34.800 149.800 35.200 ;
        RECT 151.700 34.900 152.100 35.000 ;
        RECT 144.900 34.700 145.300 34.800 ;
        RECT 142.200 33.800 142.600 34.600 ;
        RECT 145.700 34.200 146.100 34.300 ;
        RECT 149.400 34.200 149.700 34.800 ;
        RECT 150.200 34.600 152.100 34.900 ;
        RECT 150.200 34.500 150.600 34.600 ;
        RECT 144.200 33.900 149.700 34.200 ;
        RECT 144.200 33.800 145.000 33.900 ;
        RECT 139.000 32.800 141.000 33.100 ;
        RECT 139.100 32.100 139.400 32.800 ;
        RECT 140.700 32.400 141.100 32.800 ;
        RECT 139.000 31.100 139.400 32.100 ;
        RECT 141.400 31.100 141.800 33.100 ;
        RECT 143.800 31.100 144.200 33.500 ;
        RECT 146.300 32.800 146.600 33.900 ;
        RECT 149.100 33.800 149.500 33.900 ;
        RECT 152.600 33.600 153.000 35.300 ;
        RECT 155.100 35.000 155.500 35.300 ;
        RECT 155.900 35.200 156.200 35.900 ;
        RECT 158.200 35.700 158.600 39.900 ;
        RECT 160.400 38.200 160.800 39.900 ;
        RECT 159.800 37.900 160.800 38.200 ;
        RECT 162.600 37.900 163.000 39.900 ;
        RECT 164.700 37.900 165.300 39.900 ;
        RECT 159.800 37.500 160.200 37.900 ;
        RECT 162.600 37.600 162.900 37.900 ;
        RECT 161.500 37.300 163.300 37.600 ;
        RECT 164.600 37.500 165.000 37.900 ;
        RECT 161.500 37.200 161.900 37.300 ;
        RECT 162.900 37.200 163.300 37.300 ;
        RECT 159.800 36.500 160.200 36.600 ;
        RECT 162.100 36.500 162.500 36.600 ;
        RECT 159.800 36.200 162.500 36.500 ;
        RECT 162.800 36.500 163.900 36.800 ;
        RECT 162.800 35.900 163.100 36.500 ;
        RECT 163.500 36.400 163.900 36.500 ;
        RECT 164.700 36.600 165.400 37.000 ;
        RECT 164.700 36.100 165.000 36.600 ;
        RECT 160.700 35.700 163.100 35.900 ;
        RECT 158.200 35.600 163.100 35.700 ;
        RECT 163.800 35.800 165.000 36.100 ;
        RECT 158.200 35.500 161.100 35.600 ;
        RECT 158.200 35.400 161.000 35.500 ;
        RECT 154.400 34.200 154.800 34.600 ;
        RECT 154.200 33.800 154.700 34.200 ;
        RECT 151.100 33.300 153.000 33.600 ;
        RECT 155.200 33.500 155.500 35.000 ;
        RECT 155.800 34.800 156.200 35.200 ;
        RECT 161.400 35.100 161.800 35.200 ;
        RECT 151.100 33.200 151.500 33.300 ;
        RECT 145.400 32.100 145.800 32.500 ;
        RECT 146.200 32.400 146.600 32.800 ;
        RECT 147.100 32.700 147.500 32.800 ;
        RECT 147.100 32.400 148.500 32.700 ;
        RECT 148.200 32.100 148.500 32.400 ;
        RECT 150.200 32.100 150.600 32.500 ;
        RECT 145.400 31.800 146.400 32.100 ;
        RECT 146.000 31.100 146.400 31.800 ;
        RECT 148.200 31.100 148.600 32.100 ;
        RECT 150.200 31.800 150.900 32.100 ;
        RECT 150.300 31.100 150.900 31.800 ;
        RECT 152.600 31.100 153.000 33.300 ;
        RECT 154.300 33.200 155.500 33.500 ;
        RECT 153.400 32.400 153.800 33.200 ;
        RECT 154.300 32.100 154.600 33.200 ;
        RECT 155.900 33.100 156.200 34.800 ;
        RECT 159.300 34.800 161.800 35.100 ;
        RECT 159.300 34.700 159.700 34.800 ;
        RECT 160.100 34.200 160.500 34.300 ;
        RECT 163.800 34.200 164.100 35.800 ;
        RECT 167.000 35.600 167.400 39.900 ;
        RECT 165.300 35.300 167.400 35.600 ;
        RECT 167.800 37.500 168.200 39.500 ;
        RECT 169.900 39.200 170.300 39.900 ;
        RECT 169.900 38.800 170.600 39.200 ;
        RECT 167.800 35.800 168.100 37.500 ;
        RECT 169.900 36.400 170.300 38.800 ;
        RECT 169.900 36.100 170.700 36.400 ;
        RECT 173.900 36.300 174.300 39.900 ;
        RECT 167.800 35.500 169.700 35.800 ;
        RECT 165.300 35.200 165.700 35.300 ;
        RECT 166.100 34.900 166.500 35.000 ;
        RECT 164.600 34.600 166.500 34.900 ;
        RECT 164.600 34.500 165.000 34.600 ;
        RECT 158.600 33.900 164.100 34.200 ;
        RECT 158.600 33.800 159.400 33.900 ;
        RECT 154.200 31.100 154.600 32.100 ;
        RECT 155.800 31.100 156.200 33.100 ;
        RECT 158.200 31.100 158.600 33.500 ;
        RECT 160.700 32.800 161.000 33.900 ;
        RECT 163.500 33.800 163.900 33.900 ;
        RECT 167.000 33.600 167.400 35.300 ;
        RECT 167.800 34.400 168.200 35.200 ;
        RECT 168.600 34.400 169.000 35.200 ;
        RECT 169.400 34.500 169.700 35.500 ;
        RECT 169.400 34.100 170.100 34.500 ;
        RECT 170.400 34.200 170.700 36.100 ;
        RECT 173.400 35.900 174.300 36.300 ;
        RECT 175.000 35.900 175.400 39.900 ;
        RECT 175.800 36.200 176.200 39.900 ;
        RECT 177.400 36.200 177.800 39.900 ;
        RECT 175.800 35.900 177.800 36.200 ;
        RECT 171.000 35.100 171.400 35.600 ;
        RECT 171.800 35.100 172.200 35.200 ;
        RECT 171.000 34.800 172.200 35.100 ;
        RECT 173.500 34.200 173.800 35.900 ;
        RECT 174.200 34.800 174.600 35.600 ;
        RECT 175.100 35.200 175.400 35.900 ;
        RECT 178.200 35.700 178.600 39.900 ;
        RECT 180.400 38.200 180.800 39.900 ;
        RECT 179.800 37.900 180.800 38.200 ;
        RECT 182.600 37.900 183.000 39.900 ;
        RECT 184.700 37.900 185.300 39.900 ;
        RECT 179.800 37.500 180.200 37.900 ;
        RECT 182.600 37.600 182.900 37.900 ;
        RECT 181.500 37.300 183.300 37.600 ;
        RECT 184.600 37.500 185.000 37.900 ;
        RECT 181.500 37.200 181.900 37.300 ;
        RECT 182.900 37.200 183.300 37.300 ;
        RECT 185.100 37.000 185.800 37.200 ;
        RECT 184.700 36.800 185.800 37.000 ;
        RECT 179.800 36.500 180.200 36.600 ;
        RECT 182.100 36.500 182.500 36.600 ;
        RECT 179.800 36.200 182.500 36.500 ;
        RECT 182.800 36.500 183.900 36.800 ;
        RECT 182.800 35.900 183.100 36.500 ;
        RECT 183.500 36.400 183.900 36.500 ;
        RECT 184.700 36.600 185.400 36.800 ;
        RECT 184.700 36.100 185.000 36.600 ;
        RECT 180.700 35.700 183.100 35.900 ;
        RECT 178.200 35.600 183.100 35.700 ;
        RECT 183.800 35.800 185.000 36.100 ;
        RECT 178.200 35.500 181.100 35.600 ;
        RECT 178.200 35.400 181.000 35.500 ;
        RECT 177.000 35.200 177.400 35.400 ;
        RECT 175.000 34.900 176.200 35.200 ;
        RECT 177.000 34.900 177.800 35.200 ;
        RECT 181.400 35.100 181.800 35.200 ;
        RECT 175.000 34.800 175.400 34.900 ;
        RECT 169.400 33.900 169.900 34.100 ;
        RECT 165.500 33.300 167.400 33.600 ;
        RECT 165.500 33.200 165.900 33.300 ;
        RECT 159.800 32.100 160.200 32.500 ;
        RECT 160.600 32.400 161.000 32.800 ;
        RECT 161.500 32.700 161.900 32.800 ;
        RECT 161.500 32.400 162.900 32.700 ;
        RECT 162.600 32.100 162.900 32.400 ;
        RECT 164.600 32.100 165.000 32.500 ;
        RECT 159.800 31.800 160.800 32.100 ;
        RECT 160.400 31.100 160.800 31.800 ;
        RECT 162.600 31.100 163.000 32.100 ;
        RECT 164.600 31.800 165.300 32.100 ;
        RECT 164.700 31.100 165.300 31.800 ;
        RECT 167.000 31.100 167.400 33.300 ;
        RECT 167.800 33.600 169.900 33.900 ;
        RECT 170.400 33.800 171.400 34.200 ;
        RECT 173.400 33.800 173.800 34.200 ;
        RECT 167.800 32.500 168.100 33.600 ;
        RECT 170.400 33.500 170.700 33.800 ;
        RECT 170.300 33.300 170.700 33.500 ;
        RECT 169.900 33.000 170.700 33.300 ;
        RECT 167.800 31.500 168.200 32.500 ;
        RECT 169.900 31.500 170.300 33.000 ;
        RECT 172.600 32.400 173.000 33.200 ;
        RECT 173.500 33.100 173.800 33.800 ;
        RECT 175.900 33.200 176.200 34.900 ;
        RECT 177.400 34.800 177.800 34.900 ;
        RECT 179.300 34.800 181.800 35.100 ;
        RECT 179.300 34.700 179.700 34.800 ;
        RECT 176.600 33.800 177.000 34.600 ;
        RECT 180.100 34.200 180.500 34.300 ;
        RECT 183.800 34.200 184.100 35.800 ;
        RECT 187.000 35.600 187.400 39.900 ;
        RECT 185.300 35.300 187.400 35.600 ;
        RECT 187.800 37.500 188.200 39.500 ;
        RECT 187.800 35.800 188.100 37.500 ;
        RECT 189.900 36.400 190.300 39.900 ;
        RECT 189.900 36.100 190.700 36.400 ;
        RECT 187.800 35.500 189.700 35.800 ;
        RECT 185.300 35.200 185.700 35.300 ;
        RECT 186.100 34.900 186.500 35.000 ;
        RECT 184.600 34.600 186.500 34.900 ;
        RECT 184.600 34.500 185.000 34.600 ;
        RECT 178.600 33.900 184.100 34.200 ;
        RECT 178.600 33.800 179.400 33.900 ;
        RECT 175.000 33.100 175.400 33.200 ;
        RECT 173.400 32.800 175.400 33.100 ;
        RECT 173.500 32.100 173.800 32.800 ;
        RECT 175.100 32.400 175.500 32.800 ;
        RECT 173.400 31.100 173.800 32.100 ;
        RECT 175.800 31.100 176.200 33.200 ;
        RECT 178.200 31.100 178.600 33.500 ;
        RECT 180.700 32.800 181.000 33.900 ;
        RECT 183.500 33.800 183.900 33.900 ;
        RECT 187.000 33.600 187.400 35.300 ;
        RECT 187.800 34.400 188.200 35.200 ;
        RECT 188.600 34.400 189.000 35.200 ;
        RECT 189.400 34.500 189.700 35.500 ;
        RECT 189.400 34.100 190.100 34.500 ;
        RECT 190.400 34.200 190.700 36.100 ;
        RECT 191.000 35.100 191.400 35.600 ;
        RECT 192.600 35.100 193.000 39.900 ;
        RECT 194.200 37.500 194.600 39.500 ;
        RECT 196.300 39.200 196.700 39.900 ;
        RECT 200.900 39.200 201.300 39.900 ;
        RECT 196.300 38.800 197.000 39.200 ;
        RECT 200.900 38.800 201.800 39.200 ;
        RECT 194.200 35.800 194.500 37.500 ;
        RECT 196.300 36.400 196.700 38.800 ;
        RECT 200.900 36.400 201.300 38.800 ;
        RECT 203.000 37.500 203.400 39.500 ;
        RECT 196.300 36.100 197.100 36.400 ;
        RECT 194.200 35.500 196.100 35.800 ;
        RECT 191.000 34.800 193.000 35.100 ;
        RECT 189.400 33.900 189.900 34.100 ;
        RECT 185.500 33.300 187.400 33.600 ;
        RECT 185.500 33.200 185.900 33.300 ;
        RECT 179.800 32.100 180.200 32.500 ;
        RECT 180.600 32.400 181.000 32.800 ;
        RECT 181.500 32.700 181.900 32.800 ;
        RECT 181.500 32.400 182.900 32.700 ;
        RECT 182.600 32.100 182.900 32.400 ;
        RECT 184.600 32.100 185.000 32.500 ;
        RECT 179.800 31.800 180.800 32.100 ;
        RECT 180.400 31.100 180.800 31.800 ;
        RECT 182.600 31.100 183.000 32.100 ;
        RECT 184.600 31.800 185.300 32.100 ;
        RECT 184.700 31.100 185.300 31.800 ;
        RECT 187.000 31.100 187.400 33.300 ;
        RECT 187.800 33.600 189.900 33.900 ;
        RECT 190.400 33.800 191.400 34.200 ;
        RECT 187.800 32.500 188.100 33.600 ;
        RECT 190.400 33.500 190.700 33.800 ;
        RECT 190.300 33.300 190.700 33.500 ;
        RECT 189.900 33.000 190.700 33.300 ;
        RECT 189.900 32.800 190.600 33.000 ;
        RECT 187.800 31.500 188.200 32.500 ;
        RECT 189.900 31.500 190.300 32.800 ;
        RECT 192.600 31.100 193.000 34.800 ;
        RECT 194.200 34.400 194.600 35.200 ;
        RECT 195.000 34.400 195.400 35.200 ;
        RECT 195.800 34.500 196.100 35.500 ;
        RECT 193.400 33.800 193.800 34.200 ;
        RECT 195.800 34.100 196.500 34.500 ;
        RECT 196.800 34.200 197.100 36.100 ;
        RECT 200.500 36.100 201.300 36.400 ;
        RECT 197.400 34.800 197.800 35.600 ;
        RECT 199.000 35.100 199.400 35.200 ;
        RECT 199.800 35.100 200.200 35.600 ;
        RECT 199.000 34.800 200.200 35.100 ;
        RECT 200.500 34.200 200.800 36.100 ;
        RECT 203.100 35.800 203.400 37.500 ;
        RECT 203.800 36.200 204.200 39.900 ;
        RECT 205.400 36.200 205.800 39.900 ;
        RECT 203.800 35.900 205.800 36.200 ;
        RECT 206.200 35.900 206.600 39.900 ;
        RECT 207.300 36.300 207.700 39.900 ;
        RECT 212.900 39.200 213.300 39.900 ;
        RECT 212.900 38.800 213.800 39.200 ;
        RECT 212.900 36.400 213.300 38.800 ;
        RECT 215.000 37.500 215.400 39.500 ;
        RECT 207.300 35.900 208.200 36.300 ;
        RECT 212.500 36.100 213.300 36.400 ;
        RECT 201.500 35.500 203.400 35.800 ;
        RECT 201.500 34.500 201.800 35.500 ;
        RECT 204.200 35.200 204.600 35.400 ;
        RECT 206.200 35.200 206.500 35.900 ;
        RECT 195.800 33.900 196.300 34.100 ;
        RECT 193.400 33.200 193.700 33.800 ;
        RECT 194.200 33.600 196.300 33.900 ;
        RECT 196.800 33.800 197.800 34.200 ;
        RECT 199.800 33.800 200.800 34.200 ;
        RECT 201.100 34.100 201.800 34.500 ;
        RECT 202.200 34.400 202.600 35.200 ;
        RECT 203.000 34.400 203.400 35.200 ;
        RECT 203.800 34.900 204.600 35.200 ;
        RECT 205.400 34.900 206.600 35.200 ;
        RECT 203.800 34.800 204.200 34.900 ;
        RECT 193.400 32.400 193.800 33.200 ;
        RECT 194.200 32.500 194.500 33.600 ;
        RECT 196.800 33.500 197.100 33.800 ;
        RECT 196.700 33.300 197.100 33.500 ;
        RECT 196.300 33.000 197.100 33.300 ;
        RECT 200.500 33.500 200.800 33.800 ;
        RECT 201.300 33.900 201.800 34.100 ;
        RECT 201.300 33.600 203.400 33.900 ;
        RECT 204.600 33.800 205.000 34.600 ;
        RECT 200.500 33.300 200.900 33.500 ;
        RECT 200.500 33.000 201.300 33.300 ;
        RECT 194.200 31.500 194.600 32.500 ;
        RECT 196.300 31.500 196.700 33.000 ;
        RECT 200.900 31.500 201.300 33.000 ;
        RECT 203.100 32.500 203.400 33.600 ;
        RECT 203.000 31.500 203.400 32.500 ;
        RECT 205.400 33.100 205.700 34.900 ;
        RECT 206.200 34.800 206.600 34.900 ;
        RECT 207.000 34.800 207.400 35.600 ;
        RECT 207.800 34.200 208.100 35.900 ;
        RECT 211.800 34.800 212.200 35.600 ;
        RECT 212.500 34.200 212.800 36.100 ;
        RECT 215.100 35.800 215.400 37.500 ;
        RECT 217.700 39.200 218.100 39.900 ;
        RECT 217.700 38.800 218.600 39.200 ;
        RECT 217.700 36.400 218.100 38.800 ;
        RECT 219.800 37.500 220.200 39.500 ;
        RECT 213.500 35.500 215.400 35.800 ;
        RECT 217.300 36.100 218.100 36.400 ;
        RECT 213.500 34.500 213.800 35.500 ;
        RECT 207.800 33.800 208.200 34.200 ;
        RECT 211.800 33.800 212.800 34.200 ;
        RECT 213.100 34.100 213.800 34.500 ;
        RECT 214.200 34.400 214.600 35.200 ;
        RECT 215.000 34.400 215.400 35.200 ;
        RECT 215.800 35.100 216.200 35.200 ;
        RECT 216.600 35.100 217.000 35.600 ;
        RECT 215.800 34.800 217.000 35.100 ;
        RECT 217.300 34.200 217.600 36.100 ;
        RECT 219.900 35.800 220.200 37.500 ;
        RECT 220.600 36.200 221.000 39.900 ;
        RECT 222.200 36.200 222.600 39.900 ;
        RECT 220.600 35.900 222.600 36.200 ;
        RECT 223.000 35.900 223.400 39.900 ;
        RECT 225.100 36.300 225.500 39.900 ;
        RECT 224.600 35.900 225.500 36.300 ;
        RECT 226.200 37.500 226.600 39.500 ;
        RECT 228.300 39.200 228.700 39.900 ;
        RECT 227.800 38.800 228.700 39.200 ;
        RECT 218.300 35.500 220.200 35.800 ;
        RECT 218.300 34.500 218.600 35.500 ;
        RECT 221.000 35.200 221.400 35.400 ;
        RECT 223.000 35.200 223.300 35.900 ;
        RECT 206.200 33.100 206.600 33.200 ;
        RECT 207.800 33.100 208.100 33.800 ;
        RECT 212.500 33.500 212.800 33.800 ;
        RECT 213.300 33.900 213.800 34.100 ;
        RECT 213.300 33.600 215.400 33.900 ;
        RECT 216.600 33.800 217.600 34.200 ;
        RECT 217.900 34.100 218.600 34.500 ;
        RECT 219.000 34.400 219.400 35.200 ;
        RECT 219.800 34.400 220.200 35.200 ;
        RECT 220.600 34.900 221.400 35.200 ;
        RECT 222.200 34.900 223.400 35.200 ;
        RECT 220.600 34.800 221.000 34.900 ;
        RECT 212.500 33.300 212.900 33.500 ;
        RECT 205.400 31.100 205.800 33.100 ;
        RECT 206.200 32.800 208.100 33.100 ;
        RECT 206.100 32.400 206.500 32.800 ;
        RECT 207.800 32.100 208.100 32.800 ;
        RECT 208.600 33.100 209.000 33.200 ;
        RECT 209.400 33.100 209.800 33.200 ;
        RECT 208.600 32.800 209.800 33.100 ;
        RECT 212.500 33.000 213.300 33.300 ;
        RECT 208.600 32.400 209.000 32.800 ;
        RECT 207.800 31.100 208.200 32.100 ;
        RECT 212.900 31.500 213.300 33.000 ;
        RECT 215.100 32.500 215.400 33.600 ;
        RECT 217.300 33.500 217.600 33.800 ;
        RECT 218.100 33.900 218.600 34.100 ;
        RECT 218.100 33.600 220.200 33.900 ;
        RECT 221.400 33.800 221.800 34.600 ;
        RECT 217.300 33.300 217.700 33.500 ;
        RECT 217.300 33.000 218.100 33.300 ;
        RECT 215.000 31.500 215.400 32.500 ;
        RECT 217.700 31.500 218.100 33.000 ;
        RECT 219.900 32.500 220.200 33.600 ;
        RECT 219.800 31.500 220.200 32.500 ;
        RECT 222.200 33.100 222.500 34.900 ;
        RECT 223.000 34.800 223.400 34.900 ;
        RECT 224.700 34.200 225.000 35.900 ;
        RECT 226.200 35.800 226.500 37.500 ;
        RECT 228.300 36.400 228.700 38.800 ;
        RECT 228.300 36.100 229.100 36.400 ;
        RECT 225.400 34.800 225.800 35.600 ;
        RECT 226.200 35.500 228.100 35.800 ;
        RECT 226.200 34.400 226.600 35.200 ;
        RECT 227.000 34.400 227.400 35.200 ;
        RECT 227.800 34.500 228.100 35.500 ;
        RECT 224.600 34.100 225.000 34.200 ;
        RECT 223.000 33.800 225.000 34.100 ;
        RECT 227.800 34.100 228.500 34.500 ;
        RECT 228.800 34.200 229.100 36.100 ;
        RECT 229.400 35.100 229.800 35.600 ;
        RECT 231.800 35.100 232.200 39.900 ;
        RECT 234.500 37.200 234.900 39.900 ;
        RECT 233.800 36.800 234.200 37.200 ;
        RECT 234.500 36.800 235.400 37.200 ;
        RECT 232.600 35.800 233.000 36.600 ;
        RECT 233.800 36.200 234.100 36.800 ;
        RECT 234.500 36.200 234.900 36.800 ;
        RECT 233.400 35.900 234.100 36.200 ;
        RECT 234.400 35.900 234.900 36.200 ;
        RECT 233.400 35.800 233.800 35.900 ;
        RECT 233.400 35.100 233.700 35.800 ;
        RECT 229.400 34.800 230.500 35.100 ;
        RECT 227.800 33.900 228.300 34.100 ;
        RECT 223.000 33.200 223.300 33.800 ;
        RECT 222.200 31.100 222.600 33.100 ;
        RECT 223.000 32.800 223.400 33.200 ;
        RECT 222.900 32.400 223.300 32.800 ;
        RECT 223.800 32.400 224.200 33.200 ;
        RECT 224.700 32.100 225.000 33.800 ;
        RECT 224.600 31.100 225.000 32.100 ;
        RECT 226.200 33.600 228.300 33.900 ;
        RECT 228.800 33.800 229.800 34.200 ;
        RECT 230.200 34.100 230.500 34.800 ;
        RECT 231.800 34.800 233.700 35.100 ;
        RECT 231.000 34.100 231.400 34.200 ;
        RECT 230.200 33.800 231.400 34.100 ;
        RECT 226.200 32.500 226.500 33.600 ;
        RECT 228.800 33.500 229.100 33.800 ;
        RECT 228.700 33.300 229.100 33.500 ;
        RECT 231.000 33.400 231.400 33.800 ;
        RECT 228.300 33.000 229.100 33.300 ;
        RECT 231.800 33.100 232.200 34.800 ;
        RECT 234.400 34.200 234.700 35.900 ;
        RECT 236.600 35.600 237.000 39.900 ;
        RECT 238.700 37.900 239.300 39.900 ;
        RECT 241.000 37.900 241.400 39.900 ;
        RECT 243.200 38.200 243.600 39.900 ;
        RECT 243.200 37.900 244.200 38.200 ;
        RECT 239.000 37.500 239.400 37.900 ;
        RECT 241.100 37.600 241.400 37.900 ;
        RECT 240.700 37.300 242.500 37.600 ;
        RECT 243.800 37.500 244.200 37.900 ;
        RECT 240.700 37.200 241.100 37.300 ;
        RECT 242.100 37.200 242.500 37.300 ;
        RECT 238.600 36.600 239.300 37.000 ;
        RECT 239.000 36.100 239.300 36.600 ;
        RECT 240.100 36.500 241.200 36.800 ;
        RECT 240.100 36.400 240.500 36.500 ;
        RECT 239.000 35.800 240.200 36.100 ;
        RECT 236.600 35.300 238.700 35.600 ;
        RECT 235.000 34.400 235.400 35.200 ;
        RECT 233.400 33.800 234.700 34.200 ;
        RECT 235.800 34.100 236.200 34.200 ;
        RECT 235.400 33.800 236.200 34.100 ;
        RECT 233.500 33.100 233.800 33.800 ;
        RECT 235.400 33.600 235.800 33.800 ;
        RECT 236.600 33.600 237.000 35.300 ;
        RECT 238.300 35.200 238.700 35.300 ;
        RECT 237.500 34.900 237.900 35.000 ;
        RECT 237.500 34.600 239.400 34.900 ;
        RECT 239.000 34.500 239.400 34.600 ;
        RECT 239.900 34.200 240.200 35.800 ;
        RECT 240.900 35.900 241.200 36.500 ;
        RECT 241.500 36.500 241.900 36.600 ;
        RECT 243.800 36.500 244.200 36.600 ;
        RECT 241.500 36.200 244.200 36.500 ;
        RECT 240.900 35.700 243.300 35.900 ;
        RECT 245.400 35.700 245.800 39.900 ;
        RECT 247.500 36.200 247.900 39.900 ;
        RECT 248.200 36.800 248.600 37.200 ;
        RECT 248.300 36.200 248.600 36.800 ;
        RECT 247.500 35.900 248.000 36.200 ;
        RECT 248.300 35.900 249.000 36.200 ;
        RECT 240.900 35.600 245.800 35.700 ;
        RECT 242.900 35.500 245.800 35.600 ;
        RECT 243.000 35.400 245.800 35.500 ;
        RECT 241.400 35.100 241.800 35.200 ;
        RECT 242.200 35.100 242.600 35.200 ;
        RECT 241.400 34.800 244.700 35.100 ;
        RECT 244.300 34.700 244.700 34.800 ;
        RECT 247.000 34.400 247.400 35.200 ;
        RECT 243.500 34.200 243.900 34.300 ;
        RECT 247.700 34.200 248.000 35.900 ;
        RECT 248.600 35.800 249.000 35.900 ;
        RECT 249.400 35.800 249.800 36.600 ;
        RECT 248.600 35.100 248.900 35.800 ;
        RECT 250.200 35.100 250.600 39.900 ;
        RECT 251.000 37.100 251.400 37.200 ;
        RECT 251.800 37.100 252.200 39.900 ;
        RECT 253.900 37.900 254.500 39.900 ;
        RECT 256.200 37.900 256.600 39.900 ;
        RECT 258.400 38.200 258.800 39.900 ;
        RECT 258.400 37.900 259.400 38.200 ;
        RECT 254.200 37.500 254.600 37.900 ;
        RECT 256.300 37.600 256.600 37.900 ;
        RECT 255.900 37.300 257.700 37.600 ;
        RECT 259.000 37.500 259.400 37.900 ;
        RECT 255.900 37.200 256.300 37.300 ;
        RECT 257.300 37.200 257.700 37.300 ;
        RECT 251.000 36.800 252.200 37.100 ;
        RECT 248.600 34.800 250.600 35.100 ;
        RECT 239.800 33.900 245.400 34.200 ;
        RECT 239.800 33.800 240.500 33.900 ;
        RECT 236.600 33.300 238.500 33.600 ;
        RECT 234.300 33.100 236.100 33.300 ;
        RECT 226.200 31.500 226.600 32.500 ;
        RECT 228.300 31.500 228.700 33.000 ;
        RECT 231.800 32.800 232.700 33.100 ;
        RECT 232.300 31.100 232.700 32.800 ;
        RECT 233.400 31.100 233.800 33.100 ;
        RECT 234.200 33.000 236.200 33.100 ;
        RECT 234.200 31.100 234.600 33.000 ;
        RECT 235.800 31.100 236.200 33.000 ;
        RECT 236.600 31.100 237.000 33.300 ;
        RECT 238.100 33.200 238.500 33.300 ;
        RECT 243.000 32.800 243.300 33.900 ;
        RECT 244.600 33.800 245.400 33.900 ;
        RECT 246.200 34.100 246.600 34.200 ;
        RECT 247.700 34.100 249.000 34.200 ;
        RECT 249.400 34.100 249.800 34.200 ;
        RECT 246.200 33.800 247.000 34.100 ;
        RECT 247.700 33.800 249.800 34.100 ;
        RECT 246.600 33.600 247.000 33.800 ;
        RECT 242.100 32.700 242.500 32.800 ;
        RECT 239.000 32.100 239.400 32.500 ;
        RECT 241.100 32.400 242.500 32.700 ;
        RECT 243.000 32.400 243.400 32.800 ;
        RECT 241.100 32.100 241.400 32.400 ;
        RECT 243.800 32.100 244.200 32.500 ;
        RECT 238.700 31.800 239.400 32.100 ;
        RECT 238.700 31.100 239.300 31.800 ;
        RECT 241.000 31.100 241.400 32.100 ;
        RECT 243.200 31.800 244.200 32.100 ;
        RECT 243.200 31.100 243.600 31.800 ;
        RECT 245.400 31.100 245.800 33.500 ;
        RECT 246.300 33.100 248.100 33.300 ;
        RECT 248.600 33.100 248.900 33.800 ;
        RECT 250.200 33.100 250.600 34.800 ;
        RECT 251.800 35.600 252.200 36.800 ;
        RECT 253.800 36.600 254.500 37.000 ;
        RECT 254.200 36.100 254.500 36.600 ;
        RECT 255.300 36.500 256.400 36.800 ;
        RECT 255.300 36.400 255.700 36.500 ;
        RECT 254.200 35.800 255.400 36.100 ;
        RECT 251.800 35.300 253.900 35.600 ;
        RECT 251.000 33.400 251.400 34.200 ;
        RECT 251.800 33.600 252.200 35.300 ;
        RECT 253.500 35.200 253.900 35.300 ;
        RECT 252.700 34.900 253.100 35.000 ;
        RECT 252.700 34.600 254.600 34.900 ;
        RECT 254.200 34.500 254.600 34.600 ;
        RECT 255.100 34.200 255.400 35.800 ;
        RECT 256.100 35.900 256.400 36.500 ;
        RECT 256.700 36.500 257.100 36.600 ;
        RECT 259.000 36.500 259.400 36.600 ;
        RECT 256.700 36.200 259.400 36.500 ;
        RECT 256.100 35.700 258.500 35.900 ;
        RECT 260.600 35.700 261.000 39.900 ;
        RECT 262.700 36.200 263.100 39.900 ;
        RECT 263.400 36.800 263.800 37.200 ;
        RECT 263.500 36.200 263.800 36.800 ;
        RECT 262.700 35.900 263.200 36.200 ;
        RECT 263.500 35.900 264.200 36.200 ;
        RECT 256.100 35.600 261.000 35.700 ;
        RECT 258.100 35.500 261.000 35.600 ;
        RECT 258.200 35.400 261.000 35.500 ;
        RECT 257.400 35.100 257.800 35.200 ;
        RECT 261.400 35.100 261.800 35.200 ;
        RECT 262.200 35.100 262.600 35.200 ;
        RECT 257.400 34.800 259.900 35.100 ;
        RECT 261.400 34.800 262.600 35.100 ;
        RECT 259.500 34.700 259.900 34.800 ;
        RECT 262.200 34.400 262.600 34.800 ;
        RECT 258.700 34.200 259.100 34.300 ;
        RECT 262.900 34.200 263.200 35.900 ;
        RECT 263.800 35.800 264.200 35.900 ;
        RECT 255.100 33.900 260.600 34.200 ;
        RECT 255.300 33.800 255.700 33.900 ;
        RECT 256.600 33.800 257.000 33.900 ;
        RECT 246.200 33.000 248.200 33.100 ;
        RECT 246.200 31.100 246.600 33.000 ;
        RECT 247.800 31.100 248.200 33.000 ;
        RECT 248.600 31.100 249.000 33.100 ;
        RECT 249.700 32.800 250.600 33.100 ;
        RECT 251.800 33.300 253.700 33.600 ;
        RECT 249.700 31.100 250.100 32.800 ;
        RECT 251.800 31.100 252.200 33.300 ;
        RECT 253.300 33.200 253.700 33.300 ;
        RECT 258.200 32.800 258.500 33.900 ;
        RECT 259.800 33.800 260.600 33.900 ;
        RECT 261.400 34.100 261.800 34.200 ;
        RECT 261.400 33.800 262.200 34.100 ;
        RECT 262.900 33.800 264.200 34.200 ;
        RECT 261.800 33.600 262.200 33.800 ;
        RECT 257.300 32.700 257.700 32.800 ;
        RECT 254.200 32.100 254.600 32.500 ;
        RECT 256.300 32.400 257.700 32.700 ;
        RECT 258.200 32.400 258.600 32.800 ;
        RECT 256.300 32.100 256.600 32.400 ;
        RECT 259.000 32.100 259.400 32.500 ;
        RECT 253.900 31.800 254.600 32.100 ;
        RECT 253.900 31.100 254.500 31.800 ;
        RECT 256.200 31.100 256.600 32.100 ;
        RECT 258.400 31.800 259.400 32.100 ;
        RECT 258.400 31.100 258.800 31.800 ;
        RECT 260.600 31.100 261.000 33.500 ;
        RECT 261.500 33.100 263.300 33.300 ;
        RECT 263.800 33.100 264.100 33.800 ;
        RECT 261.400 33.000 263.400 33.100 ;
        RECT 261.400 31.100 261.800 33.000 ;
        RECT 263.000 31.100 263.400 33.000 ;
        RECT 263.800 31.100 264.200 33.100 ;
        RECT 0.600 27.500 1.000 29.900 ;
        RECT 2.800 29.200 3.200 29.900 ;
        RECT 2.200 28.900 3.200 29.200 ;
        RECT 5.000 28.900 5.400 29.900 ;
        RECT 7.100 29.200 7.700 29.900 ;
        RECT 7.000 28.900 7.700 29.200 ;
        RECT 2.200 28.500 2.600 28.900 ;
        RECT 5.000 28.600 5.300 28.900 ;
        RECT 3.000 28.200 3.400 28.600 ;
        RECT 3.900 28.300 5.300 28.600 ;
        RECT 7.000 28.500 7.400 28.900 ;
        RECT 3.900 28.200 4.300 28.300 ;
        RECT 1.000 27.100 1.800 27.200 ;
        RECT 3.100 27.100 3.400 28.200 ;
        RECT 7.900 27.700 8.300 27.800 ;
        RECT 9.400 27.700 9.800 29.900 ;
        RECT 7.900 27.400 9.800 27.700 ;
        RECT 5.900 27.100 6.300 27.200 ;
        RECT 1.000 26.800 6.500 27.100 ;
        RECT 2.500 26.700 2.900 26.800 ;
        RECT 1.700 26.200 2.100 26.300 ;
        RECT 3.000 26.200 3.400 26.300 ;
        RECT 6.200 26.200 6.500 26.800 ;
        RECT 7.000 26.400 7.400 26.500 ;
        RECT 1.700 25.900 4.200 26.200 ;
        RECT 3.800 25.800 4.200 25.900 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 7.000 26.100 8.900 26.400 ;
        RECT 8.500 26.000 8.900 26.100 ;
        RECT 0.600 25.500 3.400 25.600 ;
        RECT 0.600 25.400 3.500 25.500 ;
        RECT 0.600 25.300 5.500 25.400 ;
        RECT 0.600 21.100 1.000 25.300 ;
        RECT 3.100 25.100 5.500 25.300 ;
        RECT 2.200 24.500 4.900 24.800 ;
        RECT 2.200 24.400 2.600 24.500 ;
        RECT 4.500 24.400 4.900 24.500 ;
        RECT 5.200 24.500 5.500 25.100 ;
        RECT 6.200 25.200 6.500 25.800 ;
        RECT 7.700 25.700 8.100 25.800 ;
        RECT 9.400 25.700 9.800 27.400 ;
        RECT 11.000 27.600 11.400 29.900 ;
        RECT 12.600 27.600 13.000 29.900 ;
        RECT 14.200 27.600 14.600 29.900 ;
        RECT 15.800 27.600 16.200 29.900 ;
        RECT 17.400 28.500 17.800 29.500 ;
        RECT 11.000 27.200 11.900 27.600 ;
        RECT 12.600 27.200 13.700 27.600 ;
        RECT 14.200 27.200 15.300 27.600 ;
        RECT 15.800 27.200 17.000 27.600 ;
        RECT 10.200 26.900 10.600 27.200 ;
        RECT 11.500 26.900 11.900 27.200 ;
        RECT 13.300 26.900 13.700 27.200 ;
        RECT 14.900 26.900 15.300 27.200 ;
        RECT 10.200 26.500 11.100 26.900 ;
        RECT 11.500 26.500 12.800 26.900 ;
        RECT 13.300 26.500 14.500 26.900 ;
        RECT 14.900 26.500 16.200 26.900 ;
        RECT 11.500 25.800 11.900 26.500 ;
        RECT 13.300 25.800 13.700 26.500 ;
        RECT 14.900 25.800 15.300 26.500 ;
        RECT 16.600 25.800 17.000 27.200 ;
        RECT 17.400 27.400 17.700 28.500 ;
        RECT 19.500 28.000 19.900 29.500 ;
        RECT 24.100 29.200 24.500 29.500 ;
        RECT 24.100 28.800 25.000 29.200 ;
        RECT 24.100 28.000 24.500 28.800 ;
        RECT 26.200 28.500 26.600 29.500 ;
        RECT 19.500 27.700 20.300 28.000 ;
        RECT 19.900 27.500 20.300 27.700 ;
        RECT 17.400 27.100 19.500 27.400 ;
        RECT 19.000 26.900 19.500 27.100 ;
        RECT 20.000 27.200 20.300 27.500 ;
        RECT 23.700 27.700 24.500 28.000 ;
        RECT 23.700 27.500 24.100 27.700 ;
        RECT 23.700 27.200 24.000 27.500 ;
        RECT 26.300 27.400 26.600 28.500 ;
        RECT 27.000 27.500 27.400 29.900 ;
        RECT 29.200 29.200 29.600 29.900 ;
        RECT 28.600 28.900 29.600 29.200 ;
        RECT 31.400 28.900 31.800 29.900 ;
        RECT 33.500 29.200 34.100 29.900 ;
        RECT 33.400 28.900 34.100 29.200 ;
        RECT 28.600 28.500 29.000 28.900 ;
        RECT 31.400 28.600 31.700 28.900 ;
        RECT 29.400 28.200 29.800 28.600 ;
        RECT 30.300 28.300 31.700 28.600 ;
        RECT 33.400 28.500 33.800 28.900 ;
        RECT 30.300 28.200 30.700 28.300 ;
        RECT 20.000 27.100 21.000 27.200 ;
        RECT 17.400 25.800 17.800 26.600 ;
        RECT 18.200 25.800 18.600 26.600 ;
        RECT 19.000 26.500 19.700 26.900 ;
        RECT 20.000 26.800 22.500 27.100 ;
        RECT 23.000 26.800 24.000 27.200 ;
        RECT 24.500 27.100 26.600 27.400 ;
        RECT 29.500 27.200 29.800 28.200 ;
        RECT 34.300 27.700 34.700 27.800 ;
        RECT 35.800 27.700 36.200 29.900 ;
        RECT 34.300 27.400 36.200 27.700 ;
        RECT 36.600 27.500 37.000 29.900 ;
        RECT 38.800 29.200 39.200 29.900 ;
        RECT 38.200 28.900 39.200 29.200 ;
        RECT 41.000 28.900 41.400 29.900 ;
        RECT 43.100 29.200 43.700 29.900 ;
        RECT 43.000 28.900 43.700 29.200 ;
        RECT 38.200 28.500 38.600 28.900 ;
        RECT 41.000 28.600 41.300 28.900 ;
        RECT 39.000 28.200 39.400 28.600 ;
        RECT 39.900 28.300 41.300 28.600 ;
        RECT 43.000 28.500 43.400 28.900 ;
        RECT 39.900 28.200 40.300 28.300 ;
        RECT 27.400 27.100 28.200 27.200 ;
        RECT 29.400 27.100 29.800 27.200 ;
        RECT 32.300 27.100 32.700 27.200 ;
        RECT 24.500 26.900 25.000 27.100 ;
        RECT 7.700 25.400 9.800 25.700 ;
        RECT 6.200 24.900 7.400 25.200 ;
        RECT 5.900 24.500 6.300 24.600 ;
        RECT 5.200 24.200 6.300 24.500 ;
        RECT 7.100 24.400 7.400 24.900 ;
        RECT 7.100 24.000 7.800 24.400 ;
        RECT 3.900 23.700 4.300 23.800 ;
        RECT 5.300 23.700 5.700 23.800 ;
        RECT 2.200 23.100 2.600 23.500 ;
        RECT 3.900 23.400 5.700 23.700 ;
        RECT 5.000 23.100 5.300 23.400 ;
        RECT 7.000 23.100 7.400 23.500 ;
        RECT 2.200 22.800 3.200 23.100 ;
        RECT 2.800 21.100 3.200 22.800 ;
        RECT 5.000 21.100 5.400 23.100 ;
        RECT 7.100 21.100 7.700 23.100 ;
        RECT 9.400 21.100 9.800 25.400 ;
        RECT 11.000 25.400 11.900 25.800 ;
        RECT 12.600 25.400 13.700 25.800 ;
        RECT 14.200 25.400 15.300 25.800 ;
        RECT 15.800 25.400 17.000 25.800 ;
        RECT 19.000 25.500 19.300 26.500 ;
        RECT 11.000 21.100 11.400 25.400 ;
        RECT 12.600 21.100 13.000 25.400 ;
        RECT 14.200 21.100 14.600 25.400 ;
        RECT 15.800 21.100 16.200 25.400 ;
        RECT 17.400 25.200 19.300 25.500 ;
        RECT 17.400 23.500 17.700 25.200 ;
        RECT 20.000 24.900 20.300 26.800 ;
        RECT 20.600 25.400 21.000 26.200 ;
        RECT 22.200 26.100 22.500 26.800 ;
        RECT 23.000 26.100 23.400 26.200 ;
        RECT 22.200 25.800 23.400 26.100 ;
        RECT 23.000 25.400 23.400 25.800 ;
        RECT 19.500 24.600 20.300 24.900 ;
        RECT 23.700 24.900 24.000 26.800 ;
        RECT 24.300 26.500 25.000 26.900 ;
        RECT 27.400 26.800 32.900 27.100 ;
        RECT 28.900 26.700 29.300 26.800 ;
        RECT 24.700 25.500 25.000 26.500 ;
        RECT 25.400 25.800 25.800 26.600 ;
        RECT 26.200 25.800 26.600 26.600 ;
        RECT 28.100 26.200 28.500 26.300 ;
        RECT 28.100 25.900 30.600 26.200 ;
        RECT 30.200 25.800 30.600 25.900 ;
        RECT 27.000 25.500 29.800 25.600 ;
        RECT 24.700 25.200 26.600 25.500 ;
        RECT 23.700 24.600 24.500 24.900 ;
        RECT 17.400 21.500 17.800 23.500 ;
        RECT 19.500 21.100 19.900 24.600 ;
        RECT 24.100 21.100 24.500 24.600 ;
        RECT 26.300 23.500 26.600 25.200 ;
        RECT 26.200 21.500 26.600 23.500 ;
        RECT 27.000 25.400 29.900 25.500 ;
        RECT 27.000 25.300 31.900 25.400 ;
        RECT 27.000 21.100 27.400 25.300 ;
        RECT 29.500 25.100 31.900 25.300 ;
        RECT 28.600 24.500 31.300 24.800 ;
        RECT 28.600 24.400 29.000 24.500 ;
        RECT 30.900 24.400 31.300 24.500 ;
        RECT 31.600 24.500 31.900 25.100 ;
        RECT 32.600 25.200 32.900 26.800 ;
        RECT 33.400 26.400 33.800 26.500 ;
        RECT 33.400 26.100 35.300 26.400 ;
        RECT 34.900 26.000 35.300 26.100 ;
        RECT 34.100 25.700 34.500 25.800 ;
        RECT 35.800 25.700 36.200 27.400 ;
        RECT 37.000 27.100 37.800 27.200 ;
        RECT 39.100 27.100 39.400 28.200 ;
        RECT 43.900 27.700 44.300 27.800 ;
        RECT 45.400 27.700 45.800 29.900 ;
        RECT 46.300 28.200 46.700 28.600 ;
        RECT 46.200 27.800 46.600 28.200 ;
        RECT 47.000 27.900 47.400 29.900 ;
        RECT 43.900 27.400 45.800 27.700 ;
        RECT 41.900 27.100 42.300 27.200 ;
        RECT 37.000 26.800 42.500 27.100 ;
        RECT 38.500 26.700 38.900 26.800 ;
        RECT 37.700 26.200 38.100 26.300 ;
        RECT 39.000 26.200 39.400 26.300 ;
        RECT 42.200 26.200 42.500 26.800 ;
        RECT 43.000 26.400 43.400 26.500 ;
        RECT 37.700 25.900 40.200 26.200 ;
        RECT 39.800 25.800 40.200 25.900 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 43.000 26.100 44.900 26.400 ;
        RECT 44.500 26.000 44.900 26.100 ;
        RECT 34.100 25.400 36.200 25.700 ;
        RECT 32.600 24.900 33.800 25.200 ;
        RECT 32.300 24.500 32.700 24.600 ;
        RECT 31.600 24.200 32.700 24.500 ;
        RECT 33.500 24.400 33.800 24.900 ;
        RECT 33.500 24.000 34.200 24.400 ;
        RECT 30.300 23.700 30.700 23.800 ;
        RECT 31.700 23.700 32.100 23.800 ;
        RECT 28.600 23.100 29.000 23.500 ;
        RECT 30.300 23.400 32.100 23.700 ;
        RECT 31.400 23.100 31.700 23.400 ;
        RECT 33.400 23.100 33.800 23.500 ;
        RECT 28.600 22.800 29.600 23.100 ;
        RECT 29.200 21.100 29.600 22.800 ;
        RECT 31.400 21.100 31.800 23.100 ;
        RECT 33.500 21.100 34.100 23.100 ;
        RECT 35.800 21.100 36.200 25.400 ;
        RECT 36.600 25.500 39.400 25.600 ;
        RECT 36.600 25.400 39.500 25.500 ;
        RECT 36.600 25.300 41.500 25.400 ;
        RECT 36.600 21.100 37.000 25.300 ;
        RECT 39.100 25.100 41.500 25.300 ;
        RECT 38.200 24.500 40.900 24.800 ;
        RECT 38.200 24.400 38.600 24.500 ;
        RECT 40.500 24.400 40.900 24.500 ;
        RECT 41.200 24.500 41.500 25.100 ;
        RECT 42.200 25.200 42.500 25.800 ;
        RECT 43.700 25.700 44.100 25.800 ;
        RECT 45.400 25.700 45.800 27.400 ;
        RECT 46.200 26.100 46.600 26.200 ;
        RECT 47.100 26.100 47.400 27.900 ;
        RECT 49.400 27.500 49.800 29.900 ;
        RECT 51.600 29.200 52.000 29.900 ;
        RECT 51.000 28.900 52.000 29.200 ;
        RECT 53.800 28.900 54.200 29.900 ;
        RECT 55.900 29.200 56.500 29.900 ;
        RECT 55.800 28.900 56.500 29.200 ;
        RECT 58.200 29.100 58.600 29.900 ;
        RECT 59.800 29.100 60.200 29.200 ;
        RECT 51.000 28.500 51.400 28.900 ;
        RECT 53.800 28.600 54.100 28.900 ;
        RECT 51.800 28.200 52.200 28.600 ;
        RECT 52.700 28.300 54.100 28.600 ;
        RECT 55.800 28.500 56.200 28.900 ;
        RECT 58.200 28.800 60.200 29.100 ;
        RECT 52.700 28.200 53.100 28.300 ;
        RECT 47.800 27.100 48.200 27.200 ;
        RECT 48.600 27.100 49.000 27.200 ;
        RECT 47.800 26.800 49.000 27.100 ;
        RECT 49.800 27.100 50.600 27.200 ;
        RECT 51.900 27.100 52.200 28.200 ;
        RECT 56.700 27.700 57.100 27.800 ;
        RECT 58.200 27.700 58.600 28.800 ;
        RECT 60.600 28.000 61.000 29.900 ;
        RECT 62.200 28.000 62.600 29.900 ;
        RECT 60.600 27.900 62.600 28.000 ;
        RECT 63.000 27.900 63.400 29.900 ;
        RECT 60.700 27.700 62.500 27.900 ;
        RECT 56.700 27.400 58.600 27.700 ;
        RECT 54.700 27.100 55.100 27.200 ;
        RECT 49.800 26.800 55.300 27.100 ;
        RECT 47.800 26.400 48.200 26.800 ;
        RECT 51.300 26.700 51.700 26.800 ;
        RECT 50.500 26.200 50.900 26.300 ;
        RECT 48.600 26.100 49.000 26.200 ;
        RECT 46.200 25.800 47.400 26.100 ;
        RECT 48.200 25.800 49.000 26.100 ;
        RECT 50.500 25.900 53.000 26.200 ;
        RECT 52.600 25.800 53.000 25.900 ;
        RECT 43.700 25.400 45.800 25.700 ;
        RECT 42.200 24.900 43.400 25.200 ;
        RECT 41.900 24.500 42.300 24.600 ;
        RECT 41.200 24.200 42.300 24.500 ;
        RECT 43.100 24.400 43.400 24.900 ;
        RECT 43.100 24.000 43.800 24.400 ;
        RECT 39.900 23.700 40.300 23.800 ;
        RECT 41.300 23.700 41.700 23.800 ;
        RECT 38.200 23.100 38.600 23.500 ;
        RECT 39.900 23.400 41.700 23.700 ;
        RECT 41.000 23.100 41.300 23.400 ;
        RECT 43.000 23.100 43.400 23.500 ;
        RECT 38.200 22.800 39.200 23.100 ;
        RECT 38.800 21.100 39.200 22.800 ;
        RECT 41.000 21.100 41.400 23.100 ;
        RECT 43.100 21.100 43.700 23.100 ;
        RECT 45.400 21.100 45.800 25.400 ;
        RECT 46.300 25.100 46.600 25.800 ;
        RECT 48.200 25.600 48.600 25.800 ;
        RECT 49.400 25.500 52.200 25.600 ;
        RECT 49.400 25.400 52.300 25.500 ;
        RECT 49.400 25.300 54.300 25.400 ;
        RECT 46.200 21.100 46.600 25.100 ;
        RECT 47.000 24.800 49.000 25.100 ;
        RECT 47.000 21.100 47.400 24.800 ;
        RECT 48.600 21.100 49.000 24.800 ;
        RECT 49.400 21.100 49.800 25.300 ;
        RECT 51.900 25.100 54.300 25.300 ;
        RECT 51.000 24.500 53.700 24.800 ;
        RECT 51.000 24.400 51.400 24.500 ;
        RECT 53.300 24.400 53.700 24.500 ;
        RECT 54.000 24.500 54.300 25.100 ;
        RECT 55.000 25.200 55.300 26.800 ;
        RECT 55.800 26.400 56.200 26.500 ;
        RECT 55.800 26.100 57.700 26.400 ;
        RECT 57.300 26.000 57.700 26.100 ;
        RECT 56.500 25.700 56.900 25.800 ;
        RECT 58.200 25.700 58.600 27.400 ;
        RECT 61.000 27.200 61.400 27.400 ;
        RECT 63.000 27.200 63.300 27.900 ;
        RECT 63.800 27.600 64.200 29.900 ;
        RECT 65.400 28.200 65.800 29.900 ;
        RECT 65.400 27.900 65.900 28.200 ;
        RECT 67.000 28.000 67.400 29.900 ;
        RECT 68.600 28.000 69.000 29.900 ;
        RECT 67.000 27.900 69.000 28.000 ;
        RECT 69.400 27.900 69.800 29.900 ;
        RECT 70.500 28.200 70.900 29.900 ;
        RECT 70.500 27.900 71.400 28.200 ;
        RECT 63.800 27.300 65.100 27.600 ;
        RECT 60.600 26.900 61.400 27.200 ;
        RECT 60.600 26.800 61.000 26.900 ;
        RECT 62.100 26.800 63.400 27.200 ;
        RECT 61.400 25.800 61.800 26.600 ;
        RECT 56.500 25.400 58.600 25.700 ;
        RECT 55.000 24.900 56.200 25.200 ;
        RECT 54.700 24.500 55.100 24.600 ;
        RECT 54.000 24.200 55.100 24.500 ;
        RECT 55.900 24.400 56.200 24.900 ;
        RECT 55.900 24.000 56.600 24.400 ;
        RECT 52.700 23.700 53.100 23.800 ;
        RECT 54.100 23.700 54.500 23.800 ;
        RECT 51.000 23.100 51.400 23.500 ;
        RECT 52.700 23.400 54.500 23.700 ;
        RECT 53.800 23.100 54.100 23.400 ;
        RECT 55.800 23.100 56.200 23.500 ;
        RECT 51.000 22.800 52.000 23.100 ;
        RECT 51.600 21.100 52.000 22.800 ;
        RECT 53.800 21.100 54.200 23.100 ;
        RECT 55.900 21.100 56.500 23.100 ;
        RECT 58.200 21.100 58.600 25.400 ;
        RECT 62.100 25.200 62.400 26.800 ;
        RECT 63.900 26.200 64.300 26.600 ;
        RECT 63.800 25.800 64.300 26.200 ;
        RECT 64.800 26.500 65.100 27.300 ;
        RECT 65.600 27.200 65.900 27.900 ;
        RECT 67.100 27.700 68.900 27.900 ;
        RECT 67.400 27.200 67.800 27.400 ;
        RECT 69.400 27.200 69.700 27.900 ;
        RECT 65.400 27.100 65.900 27.200 ;
        RECT 67.000 27.100 67.800 27.200 ;
        RECT 65.400 26.900 67.800 27.100 ;
        RECT 65.400 26.800 67.400 26.900 ;
        RECT 68.500 26.800 69.800 27.200 ;
        RECT 64.800 26.100 65.300 26.500 ;
        RECT 61.400 24.800 62.400 25.200 ;
        RECT 63.000 25.100 63.400 25.200 ;
        RECT 64.800 25.100 65.100 26.100 ;
        RECT 65.600 25.100 65.900 26.800 ;
        RECT 67.800 25.800 68.200 26.600 ;
        RECT 68.500 25.100 68.800 26.800 ;
        RECT 71.000 26.100 71.400 27.900 ;
        RECT 72.600 27.700 73.000 29.900 ;
        RECT 74.700 29.200 75.300 29.900 ;
        RECT 74.700 28.900 75.400 29.200 ;
        RECT 77.000 28.900 77.400 29.900 ;
        RECT 79.200 29.200 79.600 29.900 ;
        RECT 79.200 28.900 80.200 29.200 ;
        RECT 75.000 28.500 75.400 28.900 ;
        RECT 77.100 28.600 77.400 28.900 ;
        RECT 77.100 28.300 78.500 28.600 ;
        RECT 78.100 28.200 78.500 28.300 ;
        RECT 79.000 28.200 79.400 28.600 ;
        RECT 79.800 28.500 80.200 28.900 ;
        RECT 74.100 27.700 74.500 27.800 ;
        RECT 69.400 25.800 71.400 26.100 ;
        RECT 71.800 26.800 72.200 27.600 ;
        RECT 72.600 27.400 74.500 27.700 ;
        RECT 71.800 26.200 72.100 26.800 ;
        RECT 71.800 25.800 72.200 26.200 ;
        RECT 69.400 25.200 69.700 25.800 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 62.700 24.800 63.400 25.100 ;
        RECT 63.800 24.800 65.100 25.100 ;
        RECT 61.900 21.100 62.300 24.800 ;
        RECT 62.700 24.200 63.000 24.800 ;
        RECT 62.600 23.800 63.000 24.200 ;
        RECT 63.800 21.100 64.200 24.800 ;
        RECT 65.400 24.600 65.900 25.100 ;
        RECT 68.300 24.800 68.800 25.100 ;
        RECT 69.100 24.800 69.800 25.100 ;
        RECT 65.400 21.100 65.800 24.600 ;
        RECT 68.300 22.200 68.700 24.800 ;
        RECT 69.100 24.200 69.400 24.800 ;
        RECT 70.200 24.400 70.600 25.200 ;
        RECT 69.000 23.800 69.400 24.200 ;
        RECT 67.800 21.800 68.700 22.200 ;
        RECT 68.300 21.100 68.700 21.800 ;
        RECT 71.000 21.100 71.400 25.800 ;
        RECT 72.600 25.700 73.000 27.400 ;
        RECT 76.100 27.100 76.500 27.200 ;
        RECT 78.200 27.100 78.600 27.200 ;
        RECT 79.000 27.100 79.300 28.200 ;
        RECT 81.400 27.500 81.800 29.900 ;
        RECT 84.100 29.200 84.500 29.500 ;
        RECT 83.800 28.800 84.500 29.200 ;
        RECT 84.100 28.000 84.500 28.800 ;
        RECT 86.200 28.500 86.600 29.500 ;
        RECT 83.700 27.700 84.500 28.000 ;
        RECT 83.700 27.500 84.100 27.700 ;
        RECT 83.700 27.200 84.000 27.500 ;
        RECT 86.300 27.400 86.600 28.500 ;
        RECT 80.600 27.100 81.400 27.200 ;
        RECT 75.900 26.800 81.400 27.100 ;
        RECT 83.000 26.800 84.000 27.200 ;
        RECT 84.500 27.100 86.600 27.400 ;
        RECT 87.000 27.800 87.400 28.600 ;
        RECT 87.000 27.200 87.300 27.800 ;
        RECT 84.500 26.900 85.000 27.100 ;
        RECT 75.000 26.400 75.400 26.500 ;
        RECT 73.500 26.100 75.400 26.400 ;
        RECT 73.500 26.000 73.900 26.100 ;
        RECT 74.300 25.700 74.700 25.800 ;
        RECT 72.600 25.400 74.700 25.700 ;
        RECT 72.600 21.100 73.000 25.400 ;
        RECT 75.900 25.200 76.200 26.800 ;
        RECT 79.500 26.700 79.900 26.800 ;
        RECT 79.000 26.200 79.400 26.300 ;
        RECT 80.300 26.200 80.700 26.300 ;
        RECT 78.200 25.900 80.700 26.200 ;
        RECT 78.200 25.800 78.600 25.900 ;
        RECT 79.000 25.500 81.800 25.600 ;
        RECT 78.900 25.400 81.800 25.500 ;
        RECT 83.000 25.400 83.400 26.200 ;
        RECT 75.000 24.900 76.200 25.200 ;
        RECT 76.900 25.300 81.800 25.400 ;
        RECT 76.900 25.100 79.300 25.300 ;
        RECT 75.000 24.400 75.300 24.900 ;
        RECT 74.600 24.000 75.300 24.400 ;
        RECT 76.100 24.500 76.500 24.600 ;
        RECT 76.900 24.500 77.200 25.100 ;
        RECT 76.100 24.200 77.200 24.500 ;
        RECT 77.500 24.500 80.200 24.800 ;
        RECT 77.500 24.400 77.900 24.500 ;
        RECT 79.800 24.400 80.200 24.500 ;
        RECT 76.700 23.700 77.100 23.800 ;
        RECT 78.100 23.700 78.500 23.800 ;
        RECT 75.000 23.100 75.400 23.500 ;
        RECT 76.700 23.400 78.500 23.700 ;
        RECT 77.100 23.100 77.400 23.400 ;
        RECT 79.800 23.100 80.200 23.500 ;
        RECT 74.700 21.100 75.300 23.100 ;
        RECT 77.000 21.100 77.400 23.100 ;
        RECT 79.200 22.800 80.200 23.100 ;
        RECT 79.200 21.100 79.600 22.800 ;
        RECT 81.400 21.100 81.800 25.300 ;
        RECT 83.700 24.900 84.000 26.800 ;
        RECT 84.300 26.500 85.000 26.900 ;
        RECT 87.000 26.800 87.400 27.200 ;
        RECT 84.700 25.500 85.000 26.500 ;
        RECT 85.400 25.800 85.800 26.600 ;
        RECT 86.200 25.800 86.600 26.600 ;
        RECT 87.800 26.100 88.200 29.900 ;
        RECT 90.500 28.000 90.900 29.500 ;
        RECT 92.600 28.500 93.000 29.500 ;
        RECT 90.100 27.700 90.900 28.000 ;
        RECT 90.100 27.500 90.500 27.700 ;
        RECT 90.100 27.200 90.400 27.500 ;
        RECT 92.700 27.400 93.000 28.500 ;
        RECT 88.600 27.100 89.000 27.200 ;
        RECT 89.400 27.100 90.400 27.200 ;
        RECT 88.600 26.800 90.400 27.100 ;
        RECT 90.900 27.100 93.000 27.400 ;
        RECT 93.400 28.500 93.800 29.500 ;
        RECT 95.500 29.200 95.900 29.500 ;
        RECT 95.000 28.800 95.900 29.200 ;
        RECT 93.400 27.400 93.700 28.500 ;
        RECT 95.500 28.000 95.900 28.800 ;
        RECT 99.000 28.200 99.400 29.900 ;
        RECT 95.500 27.700 96.300 28.000 ;
        RECT 95.900 27.500 96.300 27.700 ;
        RECT 93.400 27.100 95.500 27.400 ;
        RECT 90.900 26.900 91.400 27.100 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 87.800 25.800 89.800 26.100 ;
        RECT 84.700 25.200 86.600 25.500 ;
        RECT 83.700 24.600 84.500 24.900 ;
        RECT 84.100 21.100 84.500 24.600 ;
        RECT 86.300 23.500 86.600 25.200 ;
        RECT 86.200 21.500 86.600 23.500 ;
        RECT 87.800 21.100 88.200 25.800 ;
        RECT 89.400 25.400 89.800 25.800 ;
        RECT 90.100 24.900 90.400 26.800 ;
        RECT 90.700 26.500 91.400 26.900 ;
        RECT 95.000 26.900 95.500 27.100 ;
        RECT 96.000 27.200 96.300 27.500 ;
        RECT 98.900 27.900 99.400 28.200 ;
        RECT 98.900 27.200 99.200 27.900 ;
        RECT 100.600 27.600 101.000 29.900 ;
        RECT 101.400 28.000 101.800 29.900 ;
        RECT 103.000 28.000 103.400 29.900 ;
        RECT 101.400 27.900 103.400 28.000 ;
        RECT 103.800 27.900 104.200 29.900 ;
        RECT 104.900 28.200 105.300 29.900 ;
        RECT 107.800 29.100 108.200 29.200 ;
        RECT 108.600 29.100 109.000 29.900 ;
        RECT 107.800 28.800 109.000 29.100 ;
        RECT 110.700 29.200 111.300 29.900 ;
        RECT 110.700 28.900 111.400 29.200 ;
        RECT 113.000 28.900 113.400 29.900 ;
        RECT 115.200 29.200 115.600 29.900 ;
        RECT 115.200 28.900 116.200 29.200 ;
        RECT 104.900 27.900 105.800 28.200 ;
        RECT 101.500 27.700 103.300 27.900 ;
        RECT 99.700 27.300 101.000 27.600 ;
        RECT 91.100 25.500 91.400 26.500 ;
        RECT 91.800 25.800 92.200 26.600 ;
        RECT 92.600 25.800 93.000 26.600 ;
        RECT 93.400 25.800 93.800 26.600 ;
        RECT 94.200 25.800 94.600 26.600 ;
        RECT 95.000 26.500 95.700 26.900 ;
        RECT 96.000 26.800 97.000 27.200 ;
        RECT 98.900 26.800 99.400 27.200 ;
        RECT 95.000 25.500 95.300 26.500 ;
        RECT 91.100 25.200 93.000 25.500 ;
        RECT 90.100 24.600 90.900 24.900 ;
        RECT 90.500 21.100 90.900 24.600 ;
        RECT 92.700 23.500 93.000 25.200 ;
        RECT 92.600 21.500 93.000 23.500 ;
        RECT 93.400 25.200 95.300 25.500 ;
        RECT 93.400 23.500 93.700 25.200 ;
        RECT 96.000 24.900 96.300 26.800 ;
        RECT 96.600 26.100 97.000 26.200 ;
        RECT 98.200 26.100 98.600 26.200 ;
        RECT 96.600 25.800 98.600 26.100 ;
        RECT 96.600 25.400 97.000 25.800 ;
        RECT 95.500 24.600 96.300 24.900 ;
        RECT 98.900 25.100 99.200 26.800 ;
        RECT 99.700 26.500 100.000 27.300 ;
        RECT 101.800 27.200 102.200 27.400 ;
        RECT 103.800 27.200 104.100 27.900 ;
        RECT 101.400 26.900 102.200 27.200 ;
        RECT 102.900 27.100 104.200 27.200 ;
        RECT 104.600 27.100 105.000 27.200 ;
        RECT 101.400 26.800 101.800 26.900 ;
        RECT 102.900 26.800 105.000 27.100 ;
        RECT 99.500 26.100 100.000 26.500 ;
        RECT 99.700 25.100 100.000 26.100 ;
        RECT 100.500 26.200 100.900 26.600 ;
        RECT 100.500 25.800 101.000 26.200 ;
        RECT 102.200 25.800 102.600 26.600 ;
        RECT 102.900 25.100 103.200 26.800 ;
        RECT 105.400 26.100 105.800 27.900 ;
        RECT 108.600 27.700 109.000 28.800 ;
        RECT 111.000 28.500 111.400 28.900 ;
        RECT 113.100 28.600 113.400 28.900 ;
        RECT 113.100 28.300 114.500 28.600 ;
        RECT 114.100 28.200 114.500 28.300 ;
        RECT 115.000 28.200 115.400 28.600 ;
        RECT 115.800 28.500 116.200 28.900 ;
        RECT 110.100 27.700 110.500 27.800 ;
        RECT 106.200 27.100 106.600 27.600 ;
        RECT 108.600 27.400 110.500 27.700 ;
        RECT 107.800 27.100 108.200 27.200 ;
        RECT 106.200 26.800 108.200 27.100 ;
        RECT 103.800 25.800 105.800 26.100 ;
        RECT 103.800 25.200 104.100 25.800 ;
        RECT 103.800 25.100 104.200 25.200 ;
        RECT 98.900 24.600 99.400 25.100 ;
        RECT 99.700 24.800 101.000 25.100 ;
        RECT 93.400 21.500 93.800 23.500 ;
        RECT 95.500 21.100 95.900 24.600 ;
        RECT 99.000 21.100 99.400 24.600 ;
        RECT 100.600 21.100 101.000 24.800 ;
        RECT 102.700 24.800 103.200 25.100 ;
        RECT 103.500 24.800 104.200 25.100 ;
        RECT 102.700 21.100 103.100 24.800 ;
        RECT 103.500 24.200 103.800 24.800 ;
        RECT 104.600 24.400 105.000 25.200 ;
        RECT 103.400 23.800 103.800 24.200 ;
        RECT 105.400 21.100 105.800 25.800 ;
        RECT 108.600 25.700 109.000 27.400 ;
        RECT 112.100 27.100 112.500 27.200 ;
        RECT 115.000 27.100 115.300 28.200 ;
        RECT 117.400 27.500 117.800 29.900 ;
        RECT 118.200 28.500 118.600 29.500 ;
        RECT 120.300 29.200 120.700 29.500 ;
        RECT 120.300 28.800 121.000 29.200 ;
        RECT 118.200 27.400 118.500 28.500 ;
        RECT 120.300 28.000 120.700 28.800 ;
        RECT 123.000 28.500 123.400 29.500 ;
        RECT 120.300 27.700 121.100 28.000 ;
        RECT 120.700 27.500 121.100 27.700 ;
        RECT 116.600 27.100 117.400 27.200 ;
        RECT 118.200 27.100 120.300 27.400 ;
        RECT 111.900 26.800 117.400 27.100 ;
        RECT 119.800 26.900 120.300 27.100 ;
        RECT 120.800 27.200 121.100 27.500 ;
        RECT 123.000 27.400 123.300 28.500 ;
        RECT 125.100 28.000 125.500 29.500 ;
        RECT 125.100 27.700 125.900 28.000 ;
        RECT 125.500 27.500 125.900 27.700 ;
        RECT 111.000 26.400 111.400 26.500 ;
        RECT 109.500 26.100 111.400 26.400 ;
        RECT 109.500 26.000 109.900 26.100 ;
        RECT 110.300 25.700 110.700 25.800 ;
        RECT 108.600 25.400 110.700 25.700 ;
        RECT 108.600 21.100 109.000 25.400 ;
        RECT 111.900 25.200 112.200 26.800 ;
        RECT 115.500 26.700 115.900 26.800 ;
        RECT 116.300 26.200 116.700 26.300 ;
        RECT 114.200 25.900 116.700 26.200 ;
        RECT 114.200 25.800 114.600 25.900 ;
        RECT 118.200 25.800 118.600 26.600 ;
        RECT 119.000 25.800 119.400 26.600 ;
        RECT 119.800 26.500 120.500 26.900 ;
        RECT 120.800 26.800 121.800 27.200 ;
        RECT 123.000 27.100 125.100 27.400 ;
        RECT 124.600 26.900 125.100 27.100 ;
        RECT 125.600 27.200 125.900 27.500 ;
        RECT 125.600 27.100 126.600 27.200 ;
        RECT 127.000 27.100 127.400 27.200 ;
        RECT 115.000 25.500 117.800 25.600 ;
        RECT 119.800 25.500 120.100 26.500 ;
        RECT 114.900 25.400 117.800 25.500 ;
        RECT 111.000 24.900 112.200 25.200 ;
        RECT 112.900 25.300 117.800 25.400 ;
        RECT 112.900 25.100 115.300 25.300 ;
        RECT 111.000 24.400 111.300 24.900 ;
        RECT 110.600 24.000 111.300 24.400 ;
        RECT 112.100 24.500 112.500 24.600 ;
        RECT 112.900 24.500 113.200 25.100 ;
        RECT 112.100 24.200 113.200 24.500 ;
        RECT 113.500 24.500 116.200 24.800 ;
        RECT 113.500 24.400 113.900 24.500 ;
        RECT 115.800 24.400 116.200 24.500 ;
        RECT 112.700 23.700 113.100 23.800 ;
        RECT 114.100 23.700 114.500 23.800 ;
        RECT 111.000 23.100 111.400 23.500 ;
        RECT 112.700 23.400 114.500 23.700 ;
        RECT 113.100 23.100 113.400 23.400 ;
        RECT 115.800 23.100 116.200 23.500 ;
        RECT 110.700 21.100 111.300 23.100 ;
        RECT 113.000 21.100 113.400 23.100 ;
        RECT 115.200 22.800 116.200 23.100 ;
        RECT 115.200 21.100 115.600 22.800 ;
        RECT 117.400 21.100 117.800 25.300 ;
        RECT 118.200 25.200 120.100 25.500 ;
        RECT 118.200 23.500 118.500 25.200 ;
        RECT 120.800 24.900 121.100 26.800 ;
        RECT 121.400 25.400 121.800 26.200 ;
        RECT 123.000 25.800 123.400 26.600 ;
        RECT 123.800 25.800 124.200 26.600 ;
        RECT 124.600 26.500 125.300 26.900 ;
        RECT 125.600 26.800 127.400 27.100 ;
        RECT 124.600 25.500 124.900 26.500 ;
        RECT 120.300 24.600 121.100 24.900 ;
        RECT 123.000 25.200 124.900 25.500 ;
        RECT 118.200 21.500 118.600 23.500 ;
        RECT 120.300 21.100 120.700 24.600 ;
        RECT 123.000 23.500 123.300 25.200 ;
        RECT 125.600 24.900 125.900 26.800 ;
        RECT 126.200 26.100 126.600 26.200 ;
        RECT 127.800 26.100 128.200 29.900 ;
        RECT 128.600 28.100 129.000 28.600 ;
        RECT 129.400 28.100 129.800 29.900 ;
        RECT 131.500 29.200 132.100 29.900 ;
        RECT 131.500 28.900 132.200 29.200 ;
        RECT 133.800 28.900 134.200 29.900 ;
        RECT 136.000 29.200 136.400 29.900 ;
        RECT 136.000 28.900 137.000 29.200 ;
        RECT 131.800 28.500 132.200 28.900 ;
        RECT 133.900 28.600 134.200 28.900 ;
        RECT 133.900 28.300 135.300 28.600 ;
        RECT 134.900 28.200 135.300 28.300 ;
        RECT 135.800 28.200 136.200 28.600 ;
        RECT 136.600 28.500 137.000 28.900 ;
        RECT 128.600 27.800 129.800 28.100 ;
        RECT 126.200 25.800 128.200 26.100 ;
        RECT 126.200 25.400 126.600 25.800 ;
        RECT 125.100 24.600 125.900 24.900 ;
        RECT 123.000 21.500 123.400 23.500 ;
        RECT 125.100 21.100 125.500 24.600 ;
        RECT 127.800 21.100 128.200 25.800 ;
        RECT 129.400 27.700 129.800 27.800 ;
        RECT 130.900 27.700 131.300 27.800 ;
        RECT 129.400 27.400 131.300 27.700 ;
        RECT 129.400 25.700 129.800 27.400 ;
        RECT 132.900 27.100 133.300 27.200 ;
        RECT 135.800 27.100 136.100 28.200 ;
        RECT 138.200 27.500 138.600 29.900 ;
        RECT 139.000 27.700 139.400 29.900 ;
        RECT 141.100 29.200 141.700 29.900 ;
        RECT 141.100 28.900 141.800 29.200 ;
        RECT 143.400 28.900 143.800 29.900 ;
        RECT 145.600 29.200 146.000 29.900 ;
        RECT 145.600 28.900 146.600 29.200 ;
        RECT 141.400 28.500 141.800 28.900 ;
        RECT 143.500 28.600 143.800 28.900 ;
        RECT 143.500 28.300 144.900 28.600 ;
        RECT 144.500 28.200 144.900 28.300 ;
        RECT 145.400 28.200 145.800 28.600 ;
        RECT 146.200 28.500 146.600 28.900 ;
        RECT 140.500 27.700 140.900 27.800 ;
        RECT 139.000 27.400 140.900 27.700 ;
        RECT 137.400 27.100 138.200 27.200 ;
        RECT 132.700 26.800 138.200 27.100 ;
        RECT 131.800 26.400 132.200 26.500 ;
        RECT 130.300 26.100 132.200 26.400 ;
        RECT 130.300 26.000 130.700 26.100 ;
        RECT 131.100 25.700 131.500 25.800 ;
        RECT 129.400 25.400 131.500 25.700 ;
        RECT 129.400 21.100 129.800 25.400 ;
        RECT 132.700 25.200 133.000 26.800 ;
        RECT 136.300 26.700 136.700 26.800 ;
        RECT 137.100 26.200 137.500 26.300 ;
        RECT 135.000 25.900 137.500 26.200 ;
        RECT 135.000 25.800 135.400 25.900 ;
        RECT 139.000 25.700 139.400 27.400 ;
        RECT 142.500 27.100 142.900 27.200 ;
        RECT 145.400 27.100 145.700 28.200 ;
        RECT 147.800 27.500 148.200 29.900 ;
        RECT 148.600 28.000 149.000 29.900 ;
        RECT 150.200 28.000 150.600 29.900 ;
        RECT 148.600 27.900 150.600 28.000 ;
        RECT 151.000 27.900 151.400 29.900 ;
        RECT 152.100 28.200 152.500 29.900 ;
        RECT 152.100 27.900 153.000 28.200 ;
        RECT 148.700 27.700 150.500 27.900 ;
        RECT 149.000 27.200 149.400 27.400 ;
        RECT 151.000 27.200 151.300 27.900 ;
        RECT 147.000 27.100 147.800 27.200 ;
        RECT 142.300 26.800 147.800 27.100 ;
        RECT 148.600 26.900 149.400 27.200 ;
        RECT 148.600 26.800 149.000 26.900 ;
        RECT 150.100 26.800 151.400 27.200 ;
        RECT 141.400 26.400 141.800 26.500 ;
        RECT 139.900 26.100 141.800 26.400 ;
        RECT 142.300 26.200 142.600 26.800 ;
        RECT 145.900 26.700 146.300 26.800 ;
        RECT 146.700 26.200 147.100 26.300 ;
        RECT 139.900 26.000 140.300 26.100 ;
        RECT 142.200 25.800 142.600 26.200 ;
        RECT 144.600 25.900 147.100 26.200 ;
        RECT 144.600 25.800 145.000 25.900 ;
        RECT 149.400 25.800 149.800 26.600 ;
        RECT 140.700 25.700 141.100 25.800 ;
        RECT 135.800 25.500 138.600 25.600 ;
        RECT 135.700 25.400 138.600 25.500 ;
        RECT 131.800 24.900 133.000 25.200 ;
        RECT 133.700 25.300 138.600 25.400 ;
        RECT 133.700 25.100 136.100 25.300 ;
        RECT 131.800 24.400 132.100 24.900 ;
        RECT 131.400 24.000 132.100 24.400 ;
        RECT 132.900 24.500 133.300 24.600 ;
        RECT 133.700 24.500 134.000 25.100 ;
        RECT 132.900 24.200 134.000 24.500 ;
        RECT 134.300 24.500 137.000 24.800 ;
        RECT 134.300 24.400 134.700 24.500 ;
        RECT 136.600 24.400 137.000 24.500 ;
        RECT 133.500 23.700 133.900 23.800 ;
        RECT 134.900 23.700 135.300 23.800 ;
        RECT 131.800 23.100 132.200 23.500 ;
        RECT 133.500 23.400 135.300 23.700 ;
        RECT 133.900 23.100 134.200 23.400 ;
        RECT 136.600 23.100 137.000 23.500 ;
        RECT 131.500 21.100 132.100 23.100 ;
        RECT 133.800 21.100 134.200 23.100 ;
        RECT 136.000 22.800 137.000 23.100 ;
        RECT 136.000 21.100 136.400 22.800 ;
        RECT 138.200 21.100 138.600 25.300 ;
        RECT 139.000 25.400 141.100 25.700 ;
        RECT 139.000 21.100 139.400 25.400 ;
        RECT 142.300 25.200 142.600 25.800 ;
        RECT 145.400 25.500 148.200 25.600 ;
        RECT 145.300 25.400 148.200 25.500 ;
        RECT 141.400 24.900 142.600 25.200 ;
        RECT 143.300 25.300 148.200 25.400 ;
        RECT 143.300 25.100 145.700 25.300 ;
        RECT 141.400 24.400 141.700 24.900 ;
        RECT 141.000 24.200 141.700 24.400 ;
        RECT 142.500 24.500 142.900 24.600 ;
        RECT 143.300 24.500 143.600 25.100 ;
        RECT 142.500 24.200 143.600 24.500 ;
        RECT 143.900 24.500 146.600 24.800 ;
        RECT 143.900 24.400 144.300 24.500 ;
        RECT 146.200 24.400 146.600 24.500 ;
        RECT 140.600 24.000 141.700 24.200 ;
        RECT 140.600 23.800 141.300 24.000 ;
        RECT 143.100 23.700 143.500 23.800 ;
        RECT 144.500 23.700 144.900 23.800 ;
        RECT 141.400 23.100 141.800 23.500 ;
        RECT 143.100 23.400 144.900 23.700 ;
        RECT 143.500 23.100 143.800 23.400 ;
        RECT 146.200 23.100 146.600 23.500 ;
        RECT 141.100 21.100 141.700 23.100 ;
        RECT 143.400 21.100 143.800 23.100 ;
        RECT 145.600 22.800 146.600 23.100 ;
        RECT 145.600 21.100 146.000 22.800 ;
        RECT 147.800 21.100 148.200 25.300 ;
        RECT 150.100 25.100 150.400 26.800 ;
        RECT 152.600 26.100 153.000 27.900 ;
        RECT 153.400 27.100 153.800 27.600 ;
        RECT 155.800 27.500 156.200 29.900 ;
        RECT 158.000 29.200 158.400 29.900 ;
        RECT 157.400 28.900 158.400 29.200 ;
        RECT 160.200 28.900 160.600 29.900 ;
        RECT 162.300 29.200 162.900 29.900 ;
        RECT 162.200 28.900 162.900 29.200 ;
        RECT 157.400 28.500 157.800 28.900 ;
        RECT 160.200 28.600 160.500 28.900 ;
        RECT 158.200 28.200 158.600 28.600 ;
        RECT 159.100 28.300 160.500 28.600 ;
        RECT 162.200 28.500 162.600 28.900 ;
        RECT 159.100 28.200 159.500 28.300 ;
        RECT 155.000 27.100 155.400 27.200 ;
        RECT 153.400 26.800 155.400 27.100 ;
        RECT 156.200 27.100 157.000 27.200 ;
        RECT 158.300 27.100 158.600 28.200 ;
        RECT 163.100 27.700 163.500 27.800 ;
        RECT 164.600 27.700 165.000 29.900 ;
        RECT 165.400 28.000 165.800 29.900 ;
        RECT 167.000 28.000 167.400 29.900 ;
        RECT 165.400 27.900 167.400 28.000 ;
        RECT 167.800 27.900 168.200 29.900 ;
        RECT 168.900 28.200 169.300 29.900 ;
        RECT 168.900 27.900 169.800 28.200 ;
        RECT 165.500 27.700 167.300 27.900 ;
        RECT 163.100 27.400 165.000 27.700 ;
        RECT 161.100 27.100 161.500 27.200 ;
        RECT 156.200 26.800 161.700 27.100 ;
        RECT 157.700 26.700 158.100 26.800 ;
        RECT 151.000 25.800 153.000 26.100 ;
        RECT 156.900 26.200 157.300 26.300 ;
        RECT 158.200 26.200 158.600 26.300 ;
        RECT 156.900 25.900 159.400 26.200 ;
        RECT 159.000 25.800 159.400 25.900 ;
        RECT 151.000 25.200 151.300 25.800 ;
        RECT 151.000 25.100 151.400 25.200 ;
        RECT 149.900 24.800 150.400 25.100 ;
        RECT 150.700 24.800 151.400 25.100 ;
        RECT 149.900 21.100 150.300 24.800 ;
        RECT 150.700 24.200 151.000 24.800 ;
        RECT 151.800 24.400 152.200 25.200 ;
        RECT 150.600 23.800 151.000 24.200 ;
        RECT 152.600 21.100 153.000 25.800 ;
        RECT 155.800 25.500 158.600 25.600 ;
        RECT 155.800 25.400 158.700 25.500 ;
        RECT 155.800 25.300 160.700 25.400 ;
        RECT 155.800 21.100 156.200 25.300 ;
        RECT 158.300 25.100 160.700 25.300 ;
        RECT 157.400 24.500 160.100 24.800 ;
        RECT 157.400 24.400 157.800 24.500 ;
        RECT 159.700 24.400 160.100 24.500 ;
        RECT 160.400 24.500 160.700 25.100 ;
        RECT 161.400 25.200 161.700 26.800 ;
        RECT 162.200 26.400 162.600 26.500 ;
        RECT 162.200 26.100 164.100 26.400 ;
        RECT 163.700 26.000 164.100 26.100 ;
        RECT 162.900 25.700 163.300 25.800 ;
        RECT 164.600 25.700 165.000 27.400 ;
        RECT 165.800 27.200 166.200 27.400 ;
        RECT 167.800 27.200 168.100 27.900 ;
        RECT 165.400 26.900 166.200 27.200 ;
        RECT 165.400 26.800 165.800 26.900 ;
        RECT 166.900 26.800 168.200 27.200 ;
        RECT 166.200 25.800 166.600 26.600 ;
        RECT 162.900 25.400 165.000 25.700 ;
        RECT 161.400 24.900 162.600 25.200 ;
        RECT 161.100 24.500 161.500 24.600 ;
        RECT 160.400 24.200 161.500 24.500 ;
        RECT 162.300 24.400 162.600 24.900 ;
        RECT 162.300 24.000 163.000 24.400 ;
        RECT 159.100 23.700 159.500 23.800 ;
        RECT 160.500 23.700 160.900 23.800 ;
        RECT 157.400 23.100 157.800 23.500 ;
        RECT 159.100 23.400 160.900 23.700 ;
        RECT 160.200 23.100 160.500 23.400 ;
        RECT 162.200 23.100 162.600 23.500 ;
        RECT 157.400 22.800 158.400 23.100 ;
        RECT 158.000 21.100 158.400 22.800 ;
        RECT 160.200 21.100 160.600 23.100 ;
        RECT 162.300 21.100 162.900 23.100 ;
        RECT 164.600 21.100 165.000 25.400 ;
        RECT 166.900 25.100 167.200 26.800 ;
        RECT 169.400 26.100 169.800 27.900 ;
        RECT 171.000 27.700 171.400 29.900 ;
        RECT 173.100 29.200 173.700 29.900 ;
        RECT 173.100 28.900 173.800 29.200 ;
        RECT 175.400 28.900 175.800 29.900 ;
        RECT 177.600 29.200 178.000 29.900 ;
        RECT 177.600 28.900 178.600 29.200 ;
        RECT 173.400 28.500 173.800 28.900 ;
        RECT 175.500 28.600 175.800 28.900 ;
        RECT 175.500 28.300 176.900 28.600 ;
        RECT 176.500 28.200 176.900 28.300 ;
        RECT 177.400 28.200 177.800 28.600 ;
        RECT 178.200 28.500 178.600 28.900 ;
        RECT 172.500 27.700 172.900 27.800 ;
        RECT 170.200 27.100 170.600 27.600 ;
        RECT 171.000 27.400 172.900 27.700 ;
        RECT 171.000 27.100 171.400 27.400 ;
        RECT 174.500 27.100 174.900 27.200 ;
        RECT 177.400 27.100 177.700 28.200 ;
        RECT 179.800 27.500 180.200 29.900 ;
        RECT 181.400 28.200 181.800 29.900 ;
        RECT 181.300 27.900 181.800 28.200 ;
        RECT 181.300 27.200 181.600 27.900 ;
        RECT 183.000 27.600 183.400 29.900 ;
        RECT 182.100 27.300 183.400 27.600 ;
        RECT 183.800 28.500 184.200 29.500 ;
        RECT 183.800 27.400 184.100 28.500 ;
        RECT 185.900 28.000 186.300 29.500 ;
        RECT 185.900 27.700 186.700 28.000 ;
        RECT 186.300 27.500 186.700 27.700 ;
        RECT 179.000 27.100 179.800 27.200 ;
        RECT 170.200 26.800 171.400 27.100 ;
        RECT 167.800 25.800 169.800 26.100 ;
        RECT 167.800 25.200 168.100 25.800 ;
        RECT 167.800 25.100 168.200 25.200 ;
        RECT 166.700 24.800 167.200 25.100 ;
        RECT 167.500 24.800 168.200 25.100 ;
        RECT 166.700 24.200 167.100 24.800 ;
        RECT 167.500 24.200 167.800 24.800 ;
        RECT 168.600 24.400 169.000 25.200 ;
        RECT 166.200 23.800 167.100 24.200 ;
        RECT 167.400 23.800 167.800 24.200 ;
        RECT 166.700 21.100 167.100 23.800 ;
        RECT 169.400 21.100 169.800 25.800 ;
        RECT 171.000 25.700 171.400 26.800 ;
        RECT 174.300 26.800 179.800 27.100 ;
        RECT 181.300 26.800 181.800 27.200 ;
        RECT 173.400 26.400 173.800 26.500 ;
        RECT 171.900 26.100 173.800 26.400 ;
        RECT 171.900 26.000 172.300 26.100 ;
        RECT 172.700 25.700 173.100 25.800 ;
        RECT 171.000 25.400 173.100 25.700 ;
        RECT 171.000 21.100 171.400 25.400 ;
        RECT 174.300 25.200 174.600 26.800 ;
        RECT 177.900 26.700 178.300 26.800 ;
        RECT 178.700 26.200 179.100 26.300 ;
        RECT 175.800 26.100 176.200 26.200 ;
        RECT 176.600 26.100 179.100 26.200 ;
        RECT 175.800 25.900 179.100 26.100 ;
        RECT 175.800 25.800 177.000 25.900 ;
        RECT 177.400 25.500 180.200 25.600 ;
        RECT 177.300 25.400 180.200 25.500 ;
        RECT 173.400 24.900 174.600 25.200 ;
        RECT 175.300 25.300 180.200 25.400 ;
        RECT 175.300 25.100 177.700 25.300 ;
        RECT 173.400 24.400 173.700 24.900 ;
        RECT 173.000 24.000 173.700 24.400 ;
        RECT 174.500 24.500 174.900 24.600 ;
        RECT 175.300 24.500 175.600 25.100 ;
        RECT 174.500 24.200 175.600 24.500 ;
        RECT 175.900 24.500 178.600 24.800 ;
        RECT 175.900 24.400 176.300 24.500 ;
        RECT 178.200 24.400 178.600 24.500 ;
        RECT 175.100 23.700 175.500 23.800 ;
        RECT 176.500 23.700 176.900 23.800 ;
        RECT 173.400 23.100 173.800 23.500 ;
        RECT 175.100 23.400 176.900 23.700 ;
        RECT 175.500 23.100 175.800 23.400 ;
        RECT 178.200 23.100 178.600 23.500 ;
        RECT 173.100 21.100 173.700 23.100 ;
        RECT 175.400 21.100 175.800 23.100 ;
        RECT 177.600 22.800 178.600 23.100 ;
        RECT 177.600 21.100 178.000 22.800 ;
        RECT 179.800 21.100 180.200 25.300 ;
        RECT 181.300 25.100 181.600 26.800 ;
        RECT 182.100 26.500 182.400 27.300 ;
        RECT 183.800 27.100 185.900 27.400 ;
        RECT 185.400 26.900 185.900 27.100 ;
        RECT 186.400 27.200 186.700 27.500 ;
        RECT 181.900 26.100 182.400 26.500 ;
        RECT 182.100 25.100 182.400 26.100 ;
        RECT 182.900 26.200 183.300 26.600 ;
        RECT 182.900 25.800 183.400 26.200 ;
        RECT 183.800 25.800 184.200 26.600 ;
        RECT 184.600 25.800 185.000 26.600 ;
        RECT 185.400 26.500 186.100 26.900 ;
        RECT 186.400 26.800 187.400 27.200 ;
        RECT 185.400 25.500 185.700 26.500 ;
        RECT 183.800 25.200 185.700 25.500 ;
        RECT 181.300 24.600 181.800 25.100 ;
        RECT 182.100 24.800 183.400 25.100 ;
        RECT 181.400 21.100 181.800 24.600 ;
        RECT 183.000 21.100 183.400 24.800 ;
        RECT 183.800 23.500 184.100 25.200 ;
        RECT 186.400 24.900 186.700 26.800 ;
        RECT 187.000 26.100 187.400 26.200 ;
        RECT 188.600 26.100 189.000 29.900 ;
        RECT 189.400 27.800 189.800 28.600 ;
        RECT 187.000 25.800 189.000 26.100 ;
        RECT 187.000 25.400 187.400 25.800 ;
        RECT 185.900 24.600 186.700 24.900 ;
        RECT 183.800 21.500 184.200 23.500 ;
        RECT 185.900 22.200 186.300 24.600 ;
        RECT 185.900 21.800 186.600 22.200 ;
        RECT 185.900 21.100 186.300 21.800 ;
        RECT 188.600 21.100 189.000 25.800 ;
        RECT 190.200 27.700 190.600 29.900 ;
        RECT 192.300 29.200 192.900 29.900 ;
        RECT 192.300 28.900 193.000 29.200 ;
        RECT 194.600 28.900 195.000 29.900 ;
        RECT 196.800 29.200 197.200 29.900 ;
        RECT 196.800 28.900 197.800 29.200 ;
        RECT 192.600 28.500 193.000 28.900 ;
        RECT 194.700 28.600 195.000 28.900 ;
        RECT 194.700 28.300 196.100 28.600 ;
        RECT 195.700 28.200 196.100 28.300 ;
        RECT 196.600 28.200 197.000 28.600 ;
        RECT 197.400 28.500 197.800 28.900 ;
        RECT 191.700 27.700 192.100 27.800 ;
        RECT 190.200 27.400 192.100 27.700 ;
        RECT 190.200 25.700 190.600 27.400 ;
        RECT 196.600 27.200 196.900 28.200 ;
        RECT 199.000 27.500 199.400 29.900 ;
        RECT 199.800 28.000 200.200 29.900 ;
        RECT 201.400 28.000 201.800 29.900 ;
        RECT 199.800 27.900 201.800 28.000 ;
        RECT 202.200 27.900 202.600 29.900 ;
        RECT 203.000 27.900 203.400 29.900 ;
        RECT 203.800 28.000 204.200 29.900 ;
        RECT 205.400 28.000 205.800 29.900 ;
        RECT 203.800 27.900 205.800 28.000 ;
        RECT 199.900 27.700 201.700 27.900 ;
        RECT 200.200 27.200 200.600 27.400 ;
        RECT 202.200 27.200 202.500 27.900 ;
        RECT 203.100 27.200 203.400 27.900 ;
        RECT 203.900 27.700 205.700 27.900 ;
        RECT 207.800 27.500 208.200 29.900 ;
        RECT 210.000 29.200 210.400 29.900 ;
        RECT 209.400 28.900 210.400 29.200 ;
        RECT 212.200 28.900 212.600 29.900 ;
        RECT 214.300 29.200 214.900 29.900 ;
        RECT 214.200 28.900 214.900 29.200 ;
        RECT 209.400 28.500 209.800 28.900 ;
        RECT 212.200 28.600 212.500 28.900 ;
        RECT 210.200 28.200 210.600 28.600 ;
        RECT 211.100 28.300 212.500 28.600 ;
        RECT 214.200 28.500 214.600 28.900 ;
        RECT 211.100 28.200 211.500 28.300 ;
        RECT 205.000 27.200 205.400 27.400 ;
        RECT 193.700 27.100 194.100 27.200 ;
        RECT 196.600 27.100 197.000 27.200 ;
        RECT 198.200 27.100 199.000 27.200 ;
        RECT 193.500 26.800 199.000 27.100 ;
        RECT 199.800 26.900 200.600 27.200 ;
        RECT 199.800 26.800 200.200 26.900 ;
        RECT 201.300 26.800 202.600 27.200 ;
        RECT 203.000 26.800 204.300 27.200 ;
        RECT 205.000 26.900 205.800 27.200 ;
        RECT 205.400 26.800 205.800 26.900 ;
        RECT 208.200 27.100 209.000 27.200 ;
        RECT 210.300 27.100 210.600 28.200 ;
        RECT 215.100 27.700 215.500 27.800 ;
        RECT 216.600 27.700 217.000 29.900 ;
        RECT 215.100 27.400 217.000 27.700 ;
        RECT 213.100 27.100 213.500 27.200 ;
        RECT 208.200 26.800 213.700 27.100 ;
        RECT 192.600 26.400 193.000 26.500 ;
        RECT 191.100 26.100 193.000 26.400 ;
        RECT 191.100 26.000 191.500 26.100 ;
        RECT 191.900 25.700 192.300 25.800 ;
        RECT 190.200 25.400 192.300 25.700 ;
        RECT 190.200 21.100 190.600 25.400 ;
        RECT 193.500 25.200 193.800 26.800 ;
        RECT 197.100 26.700 197.500 26.800 ;
        RECT 197.900 26.200 198.300 26.300 ;
        RECT 195.800 25.900 198.300 26.200 ;
        RECT 195.800 25.800 196.200 25.900 ;
        RECT 200.600 25.800 201.000 26.600 ;
        RECT 196.600 25.500 199.400 25.600 ;
        RECT 196.500 25.400 199.400 25.500 ;
        RECT 192.600 24.900 193.800 25.200 ;
        RECT 194.500 25.300 199.400 25.400 ;
        RECT 194.500 25.100 196.900 25.300 ;
        RECT 192.600 24.400 192.900 24.900 ;
        RECT 192.200 24.000 192.900 24.400 ;
        RECT 193.700 24.500 194.100 24.600 ;
        RECT 194.500 24.500 194.800 25.100 ;
        RECT 193.700 24.200 194.800 24.500 ;
        RECT 195.100 24.500 197.800 24.800 ;
        RECT 195.100 24.400 195.500 24.500 ;
        RECT 197.400 24.400 197.800 24.500 ;
        RECT 194.300 23.700 194.700 23.800 ;
        RECT 195.700 23.700 196.100 23.800 ;
        RECT 192.600 23.100 193.000 23.500 ;
        RECT 194.300 23.400 196.100 23.700 ;
        RECT 194.700 23.100 195.000 23.400 ;
        RECT 197.400 23.100 197.800 23.500 ;
        RECT 192.300 21.100 192.900 23.100 ;
        RECT 194.600 21.100 195.000 23.100 ;
        RECT 196.800 22.800 197.800 23.100 ;
        RECT 196.800 21.100 197.200 22.800 ;
        RECT 199.000 21.100 199.400 25.300 ;
        RECT 201.300 25.100 201.600 26.800 ;
        RECT 204.000 26.100 204.300 26.800 ;
        RECT 209.700 26.700 210.100 26.800 ;
        RECT 202.200 25.800 204.300 26.100 ;
        RECT 204.600 25.800 205.000 26.600 ;
        RECT 208.900 26.200 209.300 26.300 ;
        RECT 210.200 26.200 210.600 26.300 ;
        RECT 213.400 26.200 213.700 26.800 ;
        RECT 214.200 26.400 214.600 26.500 ;
        RECT 208.900 25.900 211.400 26.200 ;
        RECT 211.000 25.800 211.400 25.900 ;
        RECT 213.400 25.800 213.800 26.200 ;
        RECT 214.200 26.100 216.100 26.400 ;
        RECT 215.700 26.000 216.100 26.100 ;
        RECT 202.200 25.200 202.500 25.800 ;
        RECT 202.200 25.100 202.600 25.200 ;
        RECT 201.100 24.800 201.600 25.100 ;
        RECT 201.900 24.800 202.600 25.100 ;
        RECT 203.000 25.100 203.400 25.200 ;
        RECT 204.000 25.100 204.300 25.800 ;
        RECT 207.800 25.500 210.600 25.600 ;
        RECT 207.800 25.400 210.700 25.500 ;
        RECT 207.800 25.300 212.700 25.400 ;
        RECT 203.000 24.800 203.700 25.100 ;
        RECT 204.000 24.800 204.500 25.100 ;
        RECT 201.100 21.100 201.500 24.800 ;
        RECT 201.900 24.200 202.200 24.800 ;
        RECT 201.800 23.800 202.200 24.200 ;
        RECT 203.400 24.200 203.700 24.800 ;
        RECT 203.400 23.800 203.800 24.200 ;
        RECT 204.100 21.100 204.500 24.800 ;
        RECT 207.800 21.100 208.200 25.300 ;
        RECT 210.300 25.100 212.700 25.300 ;
        RECT 209.400 24.500 212.100 24.800 ;
        RECT 209.400 24.400 209.800 24.500 ;
        RECT 211.700 24.400 212.100 24.500 ;
        RECT 212.400 24.500 212.700 25.100 ;
        RECT 213.400 25.200 213.700 25.800 ;
        RECT 214.900 25.700 215.300 25.800 ;
        RECT 216.600 25.700 217.000 27.400 ;
        RECT 217.400 28.500 217.800 29.500 ;
        RECT 219.500 29.200 219.900 29.500 ;
        RECT 219.000 28.800 219.900 29.200 ;
        RECT 217.400 27.400 217.700 28.500 ;
        RECT 219.500 28.000 219.900 28.800 ;
        RECT 219.500 27.700 220.300 28.000 ;
        RECT 219.900 27.500 220.300 27.700 ;
        RECT 217.400 27.100 219.500 27.400 ;
        RECT 219.000 26.900 219.500 27.100 ;
        RECT 220.000 27.200 220.300 27.500 ;
        RECT 222.200 27.700 222.600 29.900 ;
        RECT 224.300 29.200 224.900 29.900 ;
        RECT 224.300 28.900 225.000 29.200 ;
        RECT 226.600 28.900 227.000 29.900 ;
        RECT 228.800 29.200 229.200 29.900 ;
        RECT 228.800 28.900 229.800 29.200 ;
        RECT 224.600 28.500 225.000 28.900 ;
        RECT 226.700 28.600 227.000 28.900 ;
        RECT 226.700 28.300 228.100 28.600 ;
        RECT 227.700 28.200 228.100 28.300 ;
        RECT 228.600 28.200 229.000 28.600 ;
        RECT 229.400 28.500 229.800 28.900 ;
        RECT 223.700 27.700 224.100 27.800 ;
        RECT 222.200 27.400 224.100 27.700 ;
        RECT 217.400 25.800 217.800 26.600 ;
        RECT 218.200 25.800 218.600 26.600 ;
        RECT 219.000 26.500 219.700 26.900 ;
        RECT 220.000 26.800 221.000 27.200 ;
        RECT 214.900 25.400 217.000 25.700 ;
        RECT 219.000 25.500 219.300 26.500 ;
        RECT 213.400 24.900 214.600 25.200 ;
        RECT 213.100 24.500 213.500 24.600 ;
        RECT 212.400 24.200 213.500 24.500 ;
        RECT 214.300 24.400 214.600 24.900 ;
        RECT 214.300 24.000 215.000 24.400 ;
        RECT 211.100 23.700 211.500 23.800 ;
        RECT 212.500 23.700 212.900 23.800 ;
        RECT 209.400 23.100 209.800 23.500 ;
        RECT 211.100 23.400 212.900 23.700 ;
        RECT 212.200 23.100 212.500 23.400 ;
        RECT 214.200 23.100 214.600 23.500 ;
        RECT 209.400 22.800 210.400 23.100 ;
        RECT 210.000 21.100 210.400 22.800 ;
        RECT 212.200 21.100 212.600 23.100 ;
        RECT 214.300 21.100 214.900 23.100 ;
        RECT 216.600 21.100 217.000 25.400 ;
        RECT 217.400 25.200 219.300 25.500 ;
        RECT 217.400 23.500 217.700 25.200 ;
        RECT 220.000 24.900 220.300 26.800 ;
        RECT 220.600 25.400 221.000 26.200 ;
        RECT 222.200 25.700 222.600 27.400 ;
        RECT 225.700 27.100 226.100 27.200 ;
        RECT 228.600 27.100 228.900 28.200 ;
        RECT 231.000 27.500 231.400 29.900 ;
        RECT 230.200 27.100 231.000 27.200 ;
        RECT 225.500 26.800 231.000 27.100 ;
        RECT 224.600 26.400 225.000 26.500 ;
        RECT 223.100 26.100 225.000 26.400 ;
        RECT 223.100 26.000 223.500 26.100 ;
        RECT 223.900 25.700 224.300 25.800 ;
        RECT 222.200 25.400 224.300 25.700 ;
        RECT 219.500 24.600 220.300 24.900 ;
        RECT 217.400 21.500 217.800 23.500 ;
        RECT 219.500 21.100 219.900 24.600 ;
        RECT 222.200 21.100 222.600 25.400 ;
        RECT 225.500 25.200 225.800 26.800 ;
        RECT 229.100 26.700 229.500 26.800 ;
        RECT 229.900 26.200 230.300 26.300 ;
        RECT 226.200 26.100 226.600 26.200 ;
        RECT 227.800 26.100 230.300 26.200 ;
        RECT 226.200 25.900 230.300 26.100 ;
        RECT 226.200 25.800 228.200 25.900 ;
        RECT 228.600 25.500 231.400 25.600 ;
        RECT 228.500 25.400 231.400 25.500 ;
        RECT 224.600 24.900 225.800 25.200 ;
        RECT 226.500 25.300 231.400 25.400 ;
        RECT 226.500 25.100 228.900 25.300 ;
        RECT 224.600 24.400 224.900 24.900 ;
        RECT 224.200 24.000 224.900 24.400 ;
        RECT 225.700 24.500 226.100 24.600 ;
        RECT 226.500 24.500 226.800 25.100 ;
        RECT 225.700 24.200 226.800 24.500 ;
        RECT 227.100 24.500 229.800 24.800 ;
        RECT 227.100 24.400 227.500 24.500 ;
        RECT 229.400 24.400 229.800 24.500 ;
        RECT 226.300 23.700 226.700 23.800 ;
        RECT 227.700 23.700 228.100 23.800 ;
        RECT 224.600 23.100 225.000 23.500 ;
        RECT 226.300 23.400 228.100 23.700 ;
        RECT 226.700 23.100 227.000 23.400 ;
        RECT 229.400 23.100 229.800 23.500 ;
        RECT 224.300 21.100 224.900 23.100 ;
        RECT 226.600 21.100 227.000 23.100 ;
        RECT 228.800 22.800 229.800 23.100 ;
        RECT 228.800 21.100 229.200 22.800 ;
        RECT 231.000 21.100 231.400 25.300 ;
        RECT 231.800 21.100 232.200 29.900 ;
        RECT 232.600 27.800 233.000 28.600 ;
        RECT 233.400 27.700 233.800 29.900 ;
        RECT 235.500 29.200 236.100 29.900 ;
        RECT 235.500 28.900 236.200 29.200 ;
        RECT 237.800 28.900 238.200 29.900 ;
        RECT 240.000 29.200 240.400 29.900 ;
        RECT 240.000 28.900 241.000 29.200 ;
        RECT 235.800 28.500 236.200 28.900 ;
        RECT 237.900 28.600 238.200 28.900 ;
        RECT 237.900 28.300 239.300 28.600 ;
        RECT 238.900 28.200 239.300 28.300 ;
        RECT 239.800 28.200 240.200 28.600 ;
        RECT 240.600 28.500 241.000 28.900 ;
        RECT 234.900 27.700 235.300 27.800 ;
        RECT 233.400 27.400 235.300 27.700 ;
        RECT 233.400 25.700 233.800 27.400 ;
        RECT 236.900 27.100 237.300 27.200 ;
        RECT 238.200 27.100 238.600 27.200 ;
        RECT 239.800 27.100 240.100 28.200 ;
        RECT 242.200 27.500 242.600 29.900 ;
        RECT 244.300 28.200 244.700 29.900 ;
        RECT 243.800 27.900 244.700 28.200 ;
        RECT 245.400 27.900 245.800 29.900 ;
        RECT 246.200 28.000 246.600 29.900 ;
        RECT 247.800 28.000 248.200 29.900 ;
        RECT 246.200 27.900 248.200 28.000 ;
        RECT 248.600 28.500 249.000 29.500 ;
        RECT 250.700 29.200 251.100 29.500 ;
        RECT 250.200 28.800 251.100 29.200 ;
        RECT 241.400 27.100 242.200 27.200 ;
        RECT 236.700 26.800 242.200 27.100 ;
        RECT 243.000 26.800 243.400 27.600 ;
        RECT 235.800 26.400 236.200 26.500 ;
        RECT 234.300 26.100 236.200 26.400 ;
        RECT 234.300 26.000 234.700 26.100 ;
        RECT 235.100 25.700 235.500 25.800 ;
        RECT 233.400 25.400 235.500 25.700 ;
        RECT 233.400 21.100 233.800 25.400 ;
        RECT 236.700 25.200 237.000 26.800 ;
        RECT 240.300 26.700 240.700 26.800 ;
        RECT 239.800 26.200 240.200 26.300 ;
        RECT 241.100 26.200 241.500 26.300 ;
        RECT 239.000 25.900 241.500 26.200 ;
        RECT 243.800 26.100 244.200 27.900 ;
        RECT 245.500 27.200 245.800 27.900 ;
        RECT 246.300 27.700 248.100 27.900 ;
        RECT 248.600 27.400 248.900 28.500 ;
        RECT 250.700 28.000 251.100 28.800 ;
        RECT 250.700 27.700 251.500 28.000 ;
        RECT 251.100 27.500 251.500 27.700 ;
        RECT 247.400 27.200 247.800 27.400 ;
        RECT 244.600 27.100 245.000 27.200 ;
        RECT 245.400 27.100 246.700 27.200 ;
        RECT 244.600 26.800 246.700 27.100 ;
        RECT 247.400 26.900 248.200 27.200 ;
        RECT 248.600 27.100 250.700 27.400 ;
        RECT 247.800 26.800 248.200 26.900 ;
        RECT 250.200 26.900 250.700 27.100 ;
        RECT 251.200 27.200 251.500 27.500 ;
        RECT 253.400 27.700 253.800 29.900 ;
        RECT 255.500 29.200 256.100 29.900 ;
        RECT 255.500 28.900 256.200 29.200 ;
        RECT 257.800 28.900 258.200 29.900 ;
        RECT 260.000 29.200 260.400 29.900 ;
        RECT 260.000 28.900 261.000 29.200 ;
        RECT 255.800 28.500 256.200 28.900 ;
        RECT 257.900 28.600 258.200 28.900 ;
        RECT 257.900 28.300 259.300 28.600 ;
        RECT 258.900 28.200 259.300 28.300 ;
        RECT 259.800 28.200 260.200 28.600 ;
        RECT 260.600 28.500 261.000 28.900 ;
        RECT 254.900 27.700 255.300 27.800 ;
        RECT 253.400 27.400 255.300 27.700 ;
        RECT 239.000 25.800 239.400 25.900 ;
        RECT 243.800 25.800 245.700 26.100 ;
        RECT 239.800 25.500 242.600 25.600 ;
        RECT 239.700 25.400 242.600 25.500 ;
        RECT 235.800 24.900 237.000 25.200 ;
        RECT 237.700 25.300 242.600 25.400 ;
        RECT 237.700 25.100 240.100 25.300 ;
        RECT 235.800 24.400 236.100 24.900 ;
        RECT 235.400 24.000 236.100 24.400 ;
        RECT 236.900 24.500 237.300 24.600 ;
        RECT 237.700 24.500 238.000 25.100 ;
        RECT 236.900 24.200 238.000 24.500 ;
        RECT 238.300 24.500 241.000 24.800 ;
        RECT 238.300 24.400 238.700 24.500 ;
        RECT 240.600 24.400 241.000 24.500 ;
        RECT 237.500 23.700 237.900 23.800 ;
        RECT 238.900 23.700 239.300 23.800 ;
        RECT 235.800 23.100 236.200 23.500 ;
        RECT 237.500 23.400 239.300 23.700 ;
        RECT 237.900 23.100 238.200 23.400 ;
        RECT 240.600 23.100 241.000 23.500 ;
        RECT 235.500 21.100 236.100 23.100 ;
        RECT 237.800 21.100 238.200 23.100 ;
        RECT 240.000 22.800 241.000 23.100 ;
        RECT 240.000 21.100 240.400 22.800 ;
        RECT 242.200 21.100 242.600 25.300 ;
        RECT 243.800 21.100 244.200 25.800 ;
        RECT 245.400 25.200 245.700 25.800 ;
        RECT 244.600 24.400 245.000 25.200 ;
        RECT 245.400 25.100 245.800 25.200 ;
        RECT 246.400 25.100 246.700 26.800 ;
        RECT 247.000 25.800 247.400 26.600 ;
        RECT 248.600 25.800 249.000 26.600 ;
        RECT 249.400 25.800 249.800 26.600 ;
        RECT 250.200 26.500 250.900 26.900 ;
        RECT 251.200 26.800 252.200 27.200 ;
        RECT 250.200 25.500 250.500 26.500 ;
        RECT 248.600 25.200 250.500 25.500 ;
        RECT 245.400 24.800 246.100 25.100 ;
        RECT 246.400 24.800 246.900 25.100 ;
        RECT 245.800 24.200 246.100 24.800 ;
        RECT 245.800 23.800 246.200 24.200 ;
        RECT 246.500 21.100 246.900 24.800 ;
        RECT 248.600 23.500 248.900 25.200 ;
        RECT 251.200 24.900 251.500 26.800 ;
        RECT 251.800 26.100 252.200 26.200 ;
        RECT 252.600 26.100 253.000 26.200 ;
        RECT 251.800 25.800 253.000 26.100 ;
        RECT 251.800 25.400 252.200 25.800 ;
        RECT 253.400 25.700 253.800 27.400 ;
        RECT 256.900 27.100 257.300 27.200 ;
        RECT 259.800 27.100 260.100 28.200 ;
        RECT 262.200 27.500 262.600 29.900 ;
        RECT 261.400 27.100 262.200 27.200 ;
        RECT 256.700 26.800 262.200 27.100 ;
        RECT 255.800 26.400 256.200 26.500 ;
        RECT 254.300 26.100 256.200 26.400 ;
        RECT 254.300 26.000 254.700 26.100 ;
        RECT 255.100 25.700 255.500 25.800 ;
        RECT 253.400 25.400 255.500 25.700 ;
        RECT 250.700 24.600 251.500 24.900 ;
        RECT 248.600 21.500 249.000 23.500 ;
        RECT 250.700 21.100 251.100 24.600 ;
        RECT 253.400 21.100 253.800 25.400 ;
        RECT 256.700 25.200 257.000 26.800 ;
        RECT 260.300 26.700 260.700 26.800 ;
        RECT 259.800 26.200 260.200 26.300 ;
        RECT 261.100 26.200 261.500 26.300 ;
        RECT 259.000 25.900 261.500 26.200 ;
        RECT 259.000 25.800 259.400 25.900 ;
        RECT 259.800 25.500 262.600 25.600 ;
        RECT 259.700 25.400 262.600 25.500 ;
        RECT 255.800 24.900 257.000 25.200 ;
        RECT 257.700 25.300 262.600 25.400 ;
        RECT 257.700 25.100 260.100 25.300 ;
        RECT 255.800 24.400 256.100 24.900 ;
        RECT 255.400 24.000 256.100 24.400 ;
        RECT 256.900 24.500 257.300 24.600 ;
        RECT 257.700 24.500 258.000 25.100 ;
        RECT 256.900 24.200 258.000 24.500 ;
        RECT 258.300 24.500 261.000 24.800 ;
        RECT 258.300 24.400 258.700 24.500 ;
        RECT 260.600 24.400 261.000 24.500 ;
        RECT 257.500 23.700 257.900 23.800 ;
        RECT 258.900 23.700 259.300 23.800 ;
        RECT 255.800 23.100 256.200 23.500 ;
        RECT 257.500 23.400 259.300 23.700 ;
        RECT 257.900 23.100 258.200 23.400 ;
        RECT 260.600 23.100 261.000 23.500 ;
        RECT 255.500 21.100 256.100 23.100 ;
        RECT 257.800 21.100 258.200 23.100 ;
        RECT 260.000 22.800 261.000 23.100 ;
        RECT 260.000 21.100 260.400 22.800 ;
        RECT 262.200 21.100 262.600 25.300 ;
        RECT 0.600 15.600 1.000 19.900 ;
        RECT 2.700 17.900 3.300 19.900 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.200 18.200 7.600 19.900 ;
        RECT 7.200 17.900 8.200 18.200 ;
        RECT 3.000 17.500 3.400 17.900 ;
        RECT 5.100 17.600 5.400 17.900 ;
        RECT 4.700 17.300 6.500 17.600 ;
        RECT 7.800 17.500 8.200 17.900 ;
        RECT 4.700 17.200 5.100 17.300 ;
        RECT 6.100 17.200 6.500 17.300 ;
        RECT 2.600 16.600 3.300 17.000 ;
        RECT 3.000 16.100 3.300 16.600 ;
        RECT 4.100 16.500 5.200 16.800 ;
        RECT 4.100 16.400 4.500 16.500 ;
        RECT 3.000 15.800 4.200 16.100 ;
        RECT 0.600 15.300 2.700 15.600 ;
        RECT 0.600 13.600 1.000 15.300 ;
        RECT 2.300 15.200 2.700 15.300 ;
        RECT 1.500 14.900 1.900 15.000 ;
        RECT 1.500 14.600 3.400 14.900 ;
        RECT 3.000 14.500 3.400 14.600 ;
        RECT 3.900 14.200 4.200 15.800 ;
        RECT 4.900 15.900 5.200 16.500 ;
        RECT 5.500 16.500 5.900 16.600 ;
        RECT 7.800 16.500 8.200 16.600 ;
        RECT 5.500 16.200 8.200 16.500 ;
        RECT 4.900 15.700 7.300 15.900 ;
        RECT 9.400 15.700 9.800 19.900 ;
        RECT 10.600 16.800 11.000 17.200 ;
        RECT 10.600 16.200 10.900 16.800 ;
        RECT 11.300 16.200 11.700 19.900 ;
        RECT 10.200 15.900 10.900 16.200 ;
        RECT 11.200 15.900 11.700 16.200 ;
        RECT 14.700 16.200 15.100 19.900 ;
        RECT 15.400 16.800 15.800 17.200 ;
        RECT 15.500 16.200 15.800 16.800 ;
        RECT 14.700 15.900 15.200 16.200 ;
        RECT 15.500 15.900 16.200 16.200 ;
        RECT 10.200 15.800 10.600 15.900 ;
        RECT 4.900 15.600 9.800 15.700 ;
        RECT 6.900 15.500 9.800 15.600 ;
        RECT 7.000 15.400 9.800 15.500 ;
        RECT 11.200 15.200 11.500 15.900 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 6.200 14.800 8.700 15.100 ;
        RECT 11.000 14.800 11.500 15.200 ;
        RECT 7.000 14.700 7.400 14.800 ;
        RECT 8.300 14.700 8.700 14.800 ;
        RECT 7.500 14.200 7.900 14.300 ;
        RECT 11.200 14.200 11.500 14.800 ;
        RECT 11.800 14.400 12.200 15.200 ;
        RECT 14.200 14.400 14.600 15.200 ;
        RECT 14.900 14.200 15.200 15.900 ;
        RECT 15.800 15.800 16.200 15.900 ;
        RECT 16.600 15.800 17.000 16.600 ;
        RECT 15.800 15.100 16.100 15.800 ;
        RECT 17.400 15.100 17.800 19.900 ;
        RECT 19.000 17.500 19.400 19.500 ;
        RECT 21.100 19.200 21.500 19.900 ;
        RECT 21.100 18.800 21.800 19.200 ;
        RECT 19.000 15.800 19.300 17.500 ;
        RECT 21.100 16.400 21.500 18.800 ;
        RECT 21.100 16.100 21.900 16.400 ;
        RECT 19.000 15.500 20.900 15.800 ;
        RECT 15.800 14.800 17.800 15.100 ;
        RECT 3.900 13.900 9.400 14.200 ;
        RECT 4.100 13.800 4.500 13.900 ;
        RECT 0.600 13.300 2.500 13.600 ;
        RECT 0.600 11.100 1.000 13.300 ;
        RECT 2.100 13.200 2.500 13.300 ;
        RECT 7.000 13.200 7.300 13.900 ;
        RECT 8.600 13.800 9.400 13.900 ;
        RECT 10.200 13.800 11.500 14.200 ;
        RECT 12.600 14.100 13.000 14.200 ;
        RECT 13.400 14.100 13.800 14.200 ;
        RECT 12.200 13.800 14.200 14.100 ;
        RECT 14.900 13.800 16.200 14.200 ;
        RECT 6.100 12.700 6.500 12.800 ;
        RECT 3.000 12.100 3.400 12.500 ;
        RECT 5.100 12.400 6.500 12.700 ;
        RECT 7.000 12.400 7.400 13.200 ;
        RECT 5.100 12.100 5.400 12.400 ;
        RECT 7.800 12.100 8.200 12.500 ;
        RECT 2.700 11.800 3.400 12.100 ;
        RECT 2.700 11.100 3.300 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.200 11.800 8.200 12.100 ;
        RECT 7.200 11.100 7.600 11.800 ;
        RECT 9.400 11.100 9.800 13.500 ;
        RECT 10.300 13.100 10.600 13.800 ;
        RECT 12.200 13.600 12.600 13.800 ;
        RECT 13.800 13.600 14.200 13.800 ;
        RECT 11.100 13.100 12.900 13.300 ;
        RECT 13.500 13.100 15.300 13.300 ;
        RECT 15.800 13.100 16.100 13.800 ;
        RECT 17.400 13.100 17.800 14.800 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 18.200 14.200 18.500 14.800 ;
        RECT 19.000 14.400 19.400 15.200 ;
        RECT 19.800 14.400 20.200 15.200 ;
        RECT 20.600 14.500 20.900 15.500 ;
        RECT 18.200 13.400 18.600 14.200 ;
        RECT 20.600 14.100 21.300 14.500 ;
        RECT 21.600 14.200 21.900 16.100 ;
        RECT 23.800 15.600 24.200 19.900 ;
        RECT 25.900 17.900 26.500 19.900 ;
        RECT 28.200 17.900 28.600 19.900 ;
        RECT 30.400 18.200 30.800 19.900 ;
        RECT 30.400 17.900 31.400 18.200 ;
        RECT 26.200 17.500 26.600 17.900 ;
        RECT 28.300 17.600 28.600 17.900 ;
        RECT 27.900 17.300 29.700 17.600 ;
        RECT 31.000 17.500 31.400 17.900 ;
        RECT 27.900 17.200 28.300 17.300 ;
        RECT 29.300 17.200 29.700 17.300 ;
        RECT 25.800 16.600 26.500 17.000 ;
        RECT 26.200 16.100 26.500 16.600 ;
        RECT 27.300 16.500 28.400 16.800 ;
        RECT 27.300 16.400 27.700 16.500 ;
        RECT 26.200 15.800 27.400 16.100 ;
        RECT 22.200 15.100 22.600 15.600 ;
        RECT 23.800 15.300 25.900 15.600 ;
        RECT 23.800 15.100 24.200 15.300 ;
        RECT 25.500 15.200 25.900 15.300 ;
        RECT 22.200 14.800 24.200 15.100 ;
        RECT 20.600 13.900 21.100 14.100 ;
        RECT 19.000 13.600 21.100 13.900 ;
        RECT 21.600 13.800 22.600 14.200 ;
        RECT 10.200 11.100 10.600 13.100 ;
        RECT 11.000 13.000 13.000 13.100 ;
        RECT 11.000 11.100 11.400 13.000 ;
        RECT 12.600 11.100 13.000 13.000 ;
        RECT 13.400 13.000 15.400 13.100 ;
        RECT 13.400 11.100 13.800 13.000 ;
        RECT 15.000 11.100 15.400 13.000 ;
        RECT 15.800 11.100 16.200 13.100 ;
        RECT 16.900 12.800 17.800 13.100 ;
        RECT 16.900 11.100 17.300 12.800 ;
        RECT 19.000 12.500 19.300 13.600 ;
        RECT 21.600 13.500 21.900 13.800 ;
        RECT 21.500 13.300 21.900 13.500 ;
        RECT 21.100 13.000 21.900 13.300 ;
        RECT 23.800 13.600 24.200 14.800 ;
        RECT 24.700 14.900 25.100 15.000 ;
        RECT 24.700 14.600 26.600 14.900 ;
        RECT 26.200 14.500 26.600 14.600 ;
        RECT 27.100 14.200 27.400 15.800 ;
        RECT 28.100 15.900 28.400 16.500 ;
        RECT 28.700 16.500 29.100 16.600 ;
        RECT 31.000 16.500 31.400 16.600 ;
        RECT 28.700 16.200 31.400 16.500 ;
        RECT 28.100 15.700 30.500 15.900 ;
        RECT 32.600 15.700 33.000 19.900 ;
        RECT 34.700 16.300 35.100 19.900 ;
        RECT 34.200 15.900 35.100 16.300 ;
        RECT 35.800 15.900 36.200 19.900 ;
        RECT 36.600 16.200 37.000 19.900 ;
        RECT 38.200 16.200 38.600 19.900 ;
        RECT 39.800 16.400 40.200 19.900 ;
        RECT 36.600 15.900 38.600 16.200 ;
        RECT 39.700 15.900 40.200 16.400 ;
        RECT 41.400 16.200 41.800 19.900 ;
        RECT 40.500 15.900 41.800 16.200 ;
        RECT 28.100 15.600 33.000 15.700 ;
        RECT 30.100 15.500 33.000 15.600 ;
        RECT 30.200 15.400 33.000 15.500 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 29.400 14.800 31.900 15.100 ;
        RECT 30.200 14.700 30.600 14.800 ;
        RECT 31.500 14.700 31.900 14.800 ;
        RECT 30.700 14.200 31.100 14.300 ;
        RECT 34.300 14.200 34.600 15.900 ;
        RECT 35.000 14.800 35.400 15.600 ;
        RECT 35.900 15.200 36.200 15.900 ;
        RECT 37.800 15.200 38.200 15.400 ;
        RECT 35.800 14.900 37.000 15.200 ;
        RECT 37.800 14.900 38.600 15.200 ;
        RECT 35.800 14.800 36.200 14.900 ;
        RECT 27.100 13.900 32.600 14.200 ;
        RECT 27.300 13.800 27.700 13.900 ;
        RECT 29.400 13.800 29.800 13.900 ;
        RECT 23.800 13.300 25.700 13.600 ;
        RECT 19.000 11.500 19.400 12.500 ;
        RECT 21.100 11.500 21.500 13.000 ;
        RECT 23.800 11.100 24.200 13.300 ;
        RECT 25.300 13.200 25.700 13.300 ;
        RECT 30.200 12.800 30.500 13.900 ;
        RECT 31.800 13.800 32.600 13.900 ;
        RECT 34.200 13.800 34.600 14.200 ;
        RECT 29.300 12.700 29.700 12.800 ;
        RECT 26.200 12.100 26.600 12.500 ;
        RECT 28.300 12.400 29.700 12.700 ;
        RECT 30.200 12.400 30.600 12.800 ;
        RECT 28.300 12.100 28.600 12.400 ;
        RECT 31.000 12.100 31.400 12.500 ;
        RECT 25.900 11.800 26.600 12.100 ;
        RECT 25.900 11.100 26.500 11.800 ;
        RECT 28.200 11.100 28.600 12.100 ;
        RECT 30.400 11.800 31.400 12.100 ;
        RECT 30.400 11.100 30.800 11.800 ;
        RECT 32.600 11.100 33.000 13.500 ;
        RECT 33.400 12.400 33.800 13.200 ;
        RECT 34.300 13.100 34.600 13.800 ;
        RECT 35.800 13.100 36.200 13.200 ;
        RECT 36.700 13.100 37.000 14.900 ;
        RECT 38.200 14.800 38.600 14.900 ;
        RECT 37.400 13.800 37.800 14.600 ;
        RECT 39.700 14.200 40.000 15.900 ;
        RECT 40.500 14.900 40.800 15.900 ;
        RECT 43.000 15.600 43.400 19.900 ;
        RECT 44.600 15.600 45.000 19.900 ;
        RECT 46.200 15.600 46.600 19.900 ;
        RECT 47.800 15.600 48.200 19.900 ;
        RECT 50.200 15.600 50.600 19.900 ;
        RECT 51.800 15.600 52.200 19.900 ;
        RECT 55.800 16.400 56.200 19.900 ;
        RECT 43.000 15.200 43.900 15.600 ;
        RECT 44.600 15.200 45.700 15.600 ;
        RECT 46.200 15.200 47.300 15.600 ;
        RECT 47.800 15.200 49.000 15.600 ;
        RECT 40.300 14.500 40.800 14.900 ;
        RECT 39.700 13.800 40.200 14.200 ;
        RECT 34.200 12.800 36.200 13.100 ;
        RECT 34.300 12.100 34.600 12.800 ;
        RECT 35.900 12.400 36.300 12.800 ;
        RECT 34.200 11.100 34.600 12.100 ;
        RECT 36.600 11.100 37.000 13.100 ;
        RECT 39.700 13.200 40.000 13.800 ;
        RECT 40.500 13.700 40.800 14.500 ;
        RECT 41.300 14.800 41.800 15.200 ;
        RECT 41.300 14.400 41.700 14.800 ;
        RECT 43.500 14.500 43.900 15.200 ;
        RECT 45.300 14.500 45.700 15.200 ;
        RECT 46.900 14.500 47.300 15.200 ;
        RECT 42.200 14.100 43.100 14.500 ;
        RECT 43.500 14.100 44.800 14.500 ;
        RECT 45.300 14.100 46.500 14.500 ;
        RECT 46.900 14.100 48.200 14.500 ;
        RECT 42.200 13.800 42.600 14.100 ;
        RECT 43.500 13.800 43.900 14.100 ;
        RECT 45.300 13.800 45.700 14.100 ;
        RECT 46.900 13.800 47.300 14.100 ;
        RECT 48.600 13.800 49.000 15.200 ;
        RECT 40.500 13.400 41.800 13.700 ;
        RECT 39.700 12.800 40.200 13.200 ;
        RECT 39.800 11.100 40.200 12.800 ;
        RECT 41.400 11.100 41.800 13.400 ;
        RECT 43.000 13.400 43.900 13.800 ;
        RECT 44.600 13.400 45.700 13.800 ;
        RECT 46.200 13.400 47.300 13.800 ;
        RECT 47.800 13.400 49.000 13.800 ;
        RECT 50.200 15.200 52.200 15.600 ;
        RECT 55.700 15.900 56.200 16.400 ;
        RECT 57.400 16.200 57.800 19.900 ;
        RECT 56.500 15.900 57.800 16.200 ;
        RECT 59.500 16.200 59.900 19.900 ;
        RECT 60.200 16.800 60.600 17.200 ;
        RECT 60.300 16.200 60.600 16.800 ;
        RECT 59.500 15.900 60.000 16.200 ;
        RECT 60.300 15.900 61.000 16.200 ;
        RECT 50.200 13.800 50.600 15.200 ;
        RECT 55.700 14.200 56.000 15.900 ;
        RECT 56.500 14.900 56.800 15.900 ;
        RECT 56.300 14.500 56.800 14.900 ;
        RECT 55.700 13.800 56.200 14.200 ;
        RECT 50.200 13.400 52.200 13.800 ;
        RECT 43.000 11.100 43.400 13.400 ;
        RECT 44.600 11.100 45.000 13.400 ;
        RECT 46.200 11.100 46.600 13.400 ;
        RECT 47.800 11.100 48.200 13.400 ;
        RECT 50.200 11.100 50.600 13.400 ;
        RECT 51.800 11.100 52.200 13.400 ;
        RECT 55.700 13.100 56.000 13.800 ;
        RECT 56.500 13.700 56.800 14.500 ;
        RECT 57.300 14.800 57.800 15.200 ;
        RECT 57.300 14.400 57.700 14.800 ;
        RECT 59.000 14.400 59.400 15.200 ;
        RECT 59.700 14.200 60.000 15.900 ;
        RECT 60.600 15.800 61.000 15.900 ;
        RECT 61.400 15.800 61.800 16.600 ;
        RECT 60.600 15.100 60.900 15.800 ;
        RECT 62.200 15.100 62.600 19.900 ;
        RECT 63.800 15.700 64.200 19.900 ;
        RECT 66.000 18.200 66.400 19.900 ;
        RECT 65.400 17.900 66.400 18.200 ;
        RECT 68.200 17.900 68.600 19.900 ;
        RECT 70.300 17.900 70.900 19.900 ;
        RECT 65.400 17.500 65.800 17.900 ;
        RECT 68.200 17.600 68.500 17.900 ;
        RECT 67.100 17.300 68.900 17.600 ;
        RECT 70.200 17.500 70.600 17.900 ;
        RECT 67.100 17.200 67.500 17.300 ;
        RECT 68.500 17.200 68.900 17.300 ;
        RECT 65.400 16.500 65.800 16.600 ;
        RECT 67.700 16.500 68.100 16.600 ;
        RECT 65.400 16.200 68.100 16.500 ;
        RECT 68.400 16.500 69.500 16.800 ;
        RECT 68.400 15.900 68.700 16.500 ;
        RECT 69.100 16.400 69.500 16.500 ;
        RECT 70.300 16.600 71.000 17.000 ;
        RECT 70.300 16.100 70.600 16.600 ;
        RECT 66.300 15.700 68.700 15.900 ;
        RECT 63.800 15.600 68.700 15.700 ;
        RECT 69.400 15.800 70.600 16.100 ;
        RECT 63.800 15.500 66.700 15.600 ;
        RECT 63.800 15.400 66.600 15.500 ;
        RECT 67.000 15.100 67.400 15.200 ;
        RECT 60.600 14.800 62.600 15.100 ;
        RECT 58.200 14.100 58.600 14.200 ;
        RECT 59.700 14.100 61.000 14.200 ;
        RECT 61.400 14.100 61.800 14.200 ;
        RECT 58.200 13.800 59.000 14.100 ;
        RECT 59.700 13.800 61.800 14.100 ;
        RECT 56.500 13.400 57.800 13.700 ;
        RECT 58.600 13.600 59.000 13.800 ;
        RECT 55.700 12.800 56.200 13.100 ;
        RECT 55.800 11.100 56.200 12.800 ;
        RECT 57.400 11.100 57.800 13.400 ;
        RECT 58.300 13.100 60.100 13.300 ;
        RECT 60.600 13.100 60.900 13.800 ;
        RECT 62.200 13.100 62.600 14.800 ;
        RECT 64.900 14.800 67.400 15.100 ;
        RECT 64.900 14.700 65.300 14.800 ;
        RECT 66.200 14.700 66.600 14.800 ;
        RECT 65.700 14.200 66.100 14.300 ;
        RECT 69.400 14.200 69.700 15.800 ;
        RECT 72.600 15.600 73.000 19.900 ;
        RECT 70.900 15.300 73.000 15.600 ;
        RECT 73.400 17.500 73.800 19.500 ;
        RECT 75.500 19.200 75.900 19.900 ;
        RECT 75.000 18.800 75.900 19.200 ;
        RECT 73.400 15.800 73.700 17.500 ;
        RECT 75.500 16.400 75.900 18.800 ;
        RECT 75.500 16.100 76.300 16.400 ;
        RECT 73.400 15.500 75.300 15.800 ;
        RECT 70.900 15.200 71.300 15.300 ;
        RECT 71.700 14.900 72.100 15.000 ;
        RECT 70.200 14.600 72.100 14.900 ;
        RECT 70.200 14.500 70.600 14.600 ;
        RECT 63.000 13.400 63.400 14.200 ;
        RECT 64.200 13.900 69.700 14.200 ;
        RECT 64.200 13.800 65.000 13.900 ;
        RECT 58.200 13.000 60.200 13.100 ;
        RECT 58.200 11.100 58.600 13.000 ;
        RECT 59.800 11.100 60.200 13.000 ;
        RECT 60.600 11.100 61.000 13.100 ;
        RECT 61.700 12.800 62.600 13.100 ;
        RECT 61.700 11.100 62.100 12.800 ;
        RECT 63.800 11.100 64.200 13.500 ;
        RECT 66.300 12.800 66.600 13.900 ;
        RECT 69.100 13.800 69.500 13.900 ;
        RECT 72.600 13.600 73.000 15.300 ;
        RECT 73.400 14.400 73.800 15.200 ;
        RECT 74.200 14.400 74.600 15.200 ;
        RECT 75.000 14.500 75.300 15.500 ;
        RECT 75.000 14.100 75.700 14.500 ;
        RECT 76.000 14.200 76.300 16.100 ;
        RECT 78.200 15.700 78.600 19.900 ;
        RECT 80.400 18.200 80.800 19.900 ;
        RECT 79.800 17.900 80.800 18.200 ;
        RECT 82.600 17.900 83.000 19.900 ;
        RECT 84.700 17.900 85.300 19.900 ;
        RECT 79.800 17.500 80.200 17.900 ;
        RECT 82.600 17.600 82.900 17.900 ;
        RECT 81.500 17.300 83.300 17.600 ;
        RECT 84.600 17.500 85.000 17.900 ;
        RECT 81.500 17.200 81.900 17.300 ;
        RECT 82.900 17.200 83.300 17.300 ;
        RECT 79.800 16.500 80.200 16.600 ;
        RECT 82.100 16.500 82.500 16.600 ;
        RECT 79.800 16.200 82.500 16.500 ;
        RECT 82.800 16.500 83.900 16.800 ;
        RECT 82.800 15.900 83.100 16.500 ;
        RECT 83.500 16.400 83.900 16.500 ;
        RECT 84.700 16.600 85.400 17.000 ;
        RECT 84.700 16.100 85.000 16.600 ;
        RECT 80.700 15.700 83.100 15.900 ;
        RECT 78.200 15.600 83.100 15.700 ;
        RECT 83.800 15.800 85.000 16.100 ;
        RECT 76.600 14.800 77.000 15.600 ;
        RECT 78.200 15.500 81.100 15.600 ;
        RECT 78.200 15.400 81.000 15.500 ;
        RECT 83.800 15.200 84.100 15.800 ;
        RECT 87.000 15.600 87.400 19.900 ;
        RECT 85.300 15.300 87.400 15.600 ;
        RECT 85.300 15.200 85.700 15.300 ;
        RECT 81.400 15.100 81.800 15.200 ;
        RECT 79.300 14.800 81.800 15.100 ;
        RECT 83.800 14.800 84.200 15.200 ;
        RECT 86.100 14.900 86.500 15.000 ;
        RECT 79.300 14.700 79.700 14.800 ;
        RECT 80.600 14.700 81.000 14.800 ;
        RECT 80.100 14.200 80.500 14.300 ;
        RECT 83.800 14.200 84.100 14.800 ;
        RECT 84.600 14.600 86.500 14.900 ;
        RECT 84.600 14.500 85.000 14.600 ;
        RECT 75.000 13.900 75.500 14.100 ;
        RECT 71.100 13.300 73.000 13.600 ;
        RECT 71.100 13.200 71.500 13.300 ;
        RECT 65.400 12.100 65.800 12.500 ;
        RECT 66.200 12.400 66.600 12.800 ;
        RECT 67.100 12.700 67.500 12.800 ;
        RECT 67.100 12.400 68.500 12.700 ;
        RECT 68.200 12.100 68.500 12.400 ;
        RECT 70.200 12.100 70.600 12.500 ;
        RECT 65.400 11.800 66.400 12.100 ;
        RECT 66.000 11.100 66.400 11.800 ;
        RECT 68.200 11.100 68.600 12.100 ;
        RECT 70.200 11.800 70.900 12.100 ;
        RECT 70.300 11.100 70.900 11.800 ;
        RECT 72.600 11.100 73.000 13.300 ;
        RECT 73.400 13.600 75.500 13.900 ;
        RECT 76.000 13.800 77.000 14.200 ;
        RECT 78.600 13.900 84.100 14.200 ;
        RECT 78.600 13.800 79.400 13.900 ;
        RECT 73.400 12.500 73.700 13.600 ;
        RECT 76.000 13.500 76.300 13.800 ;
        RECT 75.900 13.300 76.300 13.500 ;
        RECT 75.500 13.000 76.300 13.300 ;
        RECT 73.400 11.500 73.800 12.500 ;
        RECT 75.500 11.500 75.900 13.000 ;
        RECT 78.200 11.100 78.600 13.500 ;
        RECT 80.700 12.800 81.000 13.900 ;
        RECT 83.500 13.800 83.900 13.900 ;
        RECT 87.000 13.600 87.400 15.300 ;
        RECT 85.500 13.300 87.400 13.600 ;
        RECT 85.500 13.200 85.900 13.300 ;
        RECT 79.800 12.100 80.200 12.500 ;
        RECT 80.600 12.400 81.000 12.800 ;
        RECT 81.500 12.700 81.900 12.800 ;
        RECT 81.500 12.400 82.900 12.700 ;
        RECT 82.600 12.100 82.900 12.400 ;
        RECT 84.600 12.100 85.000 12.500 ;
        RECT 79.800 11.800 80.800 12.100 ;
        RECT 80.400 11.100 80.800 11.800 ;
        RECT 82.600 11.100 83.000 12.100 ;
        RECT 84.600 11.800 85.300 12.100 ;
        RECT 84.700 11.100 85.300 11.800 ;
        RECT 87.000 11.100 87.400 13.300 ;
        RECT 88.600 15.100 89.000 19.900 ;
        RECT 91.300 16.400 91.700 19.900 ;
        RECT 93.400 17.500 93.800 19.500 ;
        RECT 90.900 16.100 91.700 16.400 ;
        RECT 90.900 15.800 91.400 16.100 ;
        RECT 93.500 15.800 93.800 17.500 ;
        RECT 90.200 15.100 90.600 15.600 ;
        RECT 88.600 14.800 90.600 15.100 ;
        RECT 87.800 12.400 88.200 13.200 ;
        RECT 88.600 11.100 89.000 14.800 ;
        RECT 90.900 14.200 91.200 15.800 ;
        RECT 91.900 15.500 93.800 15.800 ;
        RECT 94.200 15.600 94.600 19.900 ;
        RECT 96.300 17.900 96.900 19.900 ;
        RECT 98.600 17.900 99.000 19.900 ;
        RECT 100.800 18.200 101.200 19.900 ;
        RECT 100.800 17.900 101.800 18.200 ;
        RECT 96.600 17.500 97.000 17.900 ;
        RECT 98.700 17.600 99.000 17.900 ;
        RECT 98.300 17.300 100.100 17.600 ;
        RECT 101.400 17.500 101.800 17.900 ;
        RECT 98.300 17.200 98.700 17.300 ;
        RECT 99.700 17.200 100.100 17.300 ;
        RECT 96.200 16.600 96.900 17.000 ;
        RECT 96.600 16.100 96.900 16.600 ;
        RECT 97.700 16.500 98.800 16.800 ;
        RECT 97.700 16.400 98.100 16.500 ;
        RECT 96.600 15.800 97.800 16.100 ;
        RECT 91.900 14.500 92.200 15.500 ;
        RECT 94.200 15.300 96.300 15.600 ;
        RECT 90.200 13.800 91.200 14.200 ;
        RECT 91.500 14.100 92.200 14.500 ;
        RECT 92.600 14.400 93.000 15.200 ;
        RECT 93.400 14.400 93.800 15.200 ;
        RECT 90.900 13.500 91.200 13.800 ;
        RECT 91.700 13.900 92.200 14.100 ;
        RECT 91.700 13.600 93.800 13.900 ;
        RECT 90.900 13.300 91.300 13.500 ;
        RECT 90.900 13.000 91.700 13.300 ;
        RECT 91.300 11.500 91.700 13.000 ;
        RECT 93.500 12.500 93.800 13.600 ;
        RECT 93.400 11.500 93.800 12.500 ;
        RECT 94.200 13.600 94.600 15.300 ;
        RECT 95.900 15.200 96.300 15.300 ;
        RECT 97.500 15.200 97.800 15.800 ;
        RECT 98.500 15.900 98.800 16.500 ;
        RECT 99.100 16.500 99.500 16.600 ;
        RECT 101.400 16.500 101.800 16.600 ;
        RECT 99.100 16.200 101.800 16.500 ;
        RECT 98.500 15.700 100.900 15.900 ;
        RECT 103.000 15.700 103.400 19.900 ;
        RECT 104.600 16.400 105.000 19.900 ;
        RECT 98.500 15.600 103.400 15.700 ;
        RECT 100.500 15.500 103.400 15.600 ;
        RECT 100.600 15.400 103.400 15.500 ;
        RECT 104.500 15.900 105.000 16.400 ;
        RECT 106.200 16.200 106.600 19.900 ;
        RECT 105.300 15.900 106.600 16.200 ;
        RECT 108.600 16.200 109.000 19.900 ;
        RECT 110.200 16.200 110.600 19.900 ;
        RECT 108.600 15.900 110.600 16.200 ;
        RECT 111.000 15.900 111.400 19.900 ;
        RECT 112.100 16.300 112.500 19.900 ;
        RECT 116.100 19.200 116.500 19.900 ;
        RECT 116.100 18.800 117.000 19.200 ;
        RECT 116.100 16.400 116.500 18.800 ;
        RECT 118.200 17.500 118.600 19.500 ;
        RECT 112.100 15.900 113.000 16.300 ;
        RECT 115.700 16.100 116.500 16.400 ;
        RECT 95.100 14.900 95.500 15.000 ;
        RECT 95.100 14.600 97.000 14.900 ;
        RECT 97.400 14.800 97.800 15.200 ;
        RECT 99.800 15.100 100.200 15.200 ;
        RECT 99.800 14.800 102.300 15.100 ;
        RECT 96.600 14.500 97.000 14.600 ;
        RECT 97.500 14.200 97.800 14.800 ;
        RECT 101.900 14.700 102.300 14.800 ;
        RECT 101.100 14.200 101.500 14.300 ;
        RECT 104.500 14.200 104.800 15.900 ;
        RECT 105.300 14.900 105.600 15.900 ;
        RECT 109.000 15.200 109.400 15.400 ;
        RECT 111.000 15.200 111.300 15.900 ;
        RECT 105.100 14.500 105.600 14.900 ;
        RECT 97.500 13.900 103.000 14.200 ;
        RECT 97.700 13.800 98.100 13.900 ;
        RECT 94.200 13.300 96.100 13.600 ;
        RECT 94.200 11.100 94.600 13.300 ;
        RECT 95.700 13.200 96.100 13.300 ;
        RECT 100.600 12.800 100.900 13.900 ;
        RECT 102.200 13.800 103.000 13.900 ;
        RECT 104.500 13.800 105.000 14.200 ;
        RECT 99.700 12.700 100.100 12.800 ;
        RECT 96.600 12.100 97.000 12.500 ;
        RECT 98.700 12.400 100.100 12.700 ;
        RECT 100.600 12.400 101.000 12.800 ;
        RECT 98.700 12.100 99.000 12.400 ;
        RECT 101.400 12.100 101.800 12.500 ;
        RECT 96.300 11.800 97.000 12.100 ;
        RECT 96.300 11.100 96.900 11.800 ;
        RECT 98.600 11.100 99.000 12.100 ;
        RECT 100.800 11.800 101.800 12.100 ;
        RECT 100.800 11.100 101.200 11.800 ;
        RECT 103.000 11.100 103.400 13.500 ;
        RECT 104.500 13.100 104.800 13.800 ;
        RECT 105.300 13.700 105.600 14.500 ;
        RECT 106.100 14.800 106.600 15.200 ;
        RECT 108.600 14.900 109.400 15.200 ;
        RECT 110.200 14.900 111.400 15.200 ;
        RECT 108.600 14.800 109.000 14.900 ;
        RECT 106.100 14.400 106.500 14.800 ;
        RECT 109.400 13.800 109.800 14.600 ;
        RECT 105.300 13.400 106.600 13.700 ;
        RECT 104.500 12.800 105.000 13.100 ;
        RECT 104.600 11.100 105.000 12.800 ;
        RECT 106.200 11.100 106.600 13.400 ;
        RECT 110.200 13.100 110.500 14.900 ;
        RECT 111.000 14.800 111.400 14.900 ;
        RECT 111.800 14.800 112.200 15.600 ;
        RECT 111.000 14.200 111.300 14.800 ;
        RECT 112.600 14.200 112.900 15.900 ;
        RECT 113.400 15.100 113.800 15.200 ;
        RECT 115.000 15.100 115.400 15.600 ;
        RECT 113.400 14.800 115.400 15.100 ;
        RECT 115.700 14.200 116.000 16.100 ;
        RECT 118.300 15.800 118.600 17.500 ;
        RECT 120.900 19.200 121.300 19.900 ;
        RECT 120.900 18.800 121.800 19.200 ;
        RECT 120.900 16.400 121.300 18.800 ;
        RECT 123.000 17.500 123.400 19.500 ;
        RECT 116.700 15.500 118.600 15.800 ;
        RECT 120.500 16.100 121.300 16.400 ;
        RECT 116.700 14.500 117.000 15.500 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 112.600 13.800 113.000 14.200 ;
        RECT 115.000 13.800 116.000 14.200 ;
        RECT 116.300 14.100 117.000 14.500 ;
        RECT 117.400 14.400 117.800 15.200 ;
        RECT 118.200 14.400 118.600 15.200 ;
        RECT 119.800 14.800 120.200 15.600 ;
        RECT 120.500 14.200 120.800 16.100 ;
        RECT 123.100 15.800 123.400 17.500 ;
        RECT 121.500 15.500 123.400 15.800 ;
        RECT 123.800 15.600 124.200 19.900 ;
        RECT 125.900 17.900 126.500 19.900 ;
        RECT 128.200 17.900 128.600 19.900 ;
        RECT 130.400 18.200 130.800 19.900 ;
        RECT 130.400 17.900 131.400 18.200 ;
        RECT 126.200 17.500 126.600 17.900 ;
        RECT 128.300 17.600 128.600 17.900 ;
        RECT 127.900 17.300 129.700 17.600 ;
        RECT 131.000 17.500 131.400 17.900 ;
        RECT 127.900 17.200 128.300 17.300 ;
        RECT 129.300 17.200 129.700 17.300 ;
        RECT 125.800 16.600 126.500 17.000 ;
        RECT 126.200 16.100 126.500 16.600 ;
        RECT 127.300 16.500 128.400 16.800 ;
        RECT 127.300 16.400 127.700 16.500 ;
        RECT 126.200 15.800 127.400 16.100 ;
        RECT 121.500 14.500 121.800 15.500 ;
        RECT 123.800 15.300 125.900 15.600 ;
        RECT 111.000 13.100 111.400 13.200 ;
        RECT 112.600 13.100 112.900 13.800 ;
        RECT 115.700 13.500 116.000 13.800 ;
        RECT 116.500 13.900 117.000 14.100 ;
        RECT 116.500 13.600 118.600 13.900 ;
        RECT 119.800 13.800 120.800 14.200 ;
        RECT 121.100 14.100 121.800 14.500 ;
        RECT 122.200 14.400 122.600 15.200 ;
        RECT 123.000 14.400 123.400 15.200 ;
        RECT 115.700 13.300 116.100 13.500 ;
        RECT 110.200 11.100 110.600 13.100 ;
        RECT 111.000 12.800 112.900 13.100 ;
        RECT 110.900 12.400 111.300 12.800 ;
        RECT 112.600 12.100 112.900 12.800 ;
        RECT 113.400 12.400 113.800 13.200 ;
        RECT 115.700 13.000 116.500 13.300 ;
        RECT 112.600 11.100 113.000 12.100 ;
        RECT 116.100 11.500 116.500 13.000 ;
        RECT 118.300 12.500 118.600 13.600 ;
        RECT 120.500 13.500 120.800 13.800 ;
        RECT 121.300 13.900 121.800 14.100 ;
        RECT 121.300 13.600 123.400 13.900 ;
        RECT 120.500 13.300 120.900 13.500 ;
        RECT 120.500 13.000 121.300 13.300 ;
        RECT 118.200 11.500 118.600 12.500 ;
        RECT 120.900 11.500 121.300 13.000 ;
        RECT 123.100 12.500 123.400 13.600 ;
        RECT 123.000 11.500 123.400 12.500 ;
        RECT 123.800 13.600 124.200 15.300 ;
        RECT 125.500 15.200 125.900 15.300 ;
        RECT 124.700 14.900 125.100 15.000 ;
        RECT 124.700 14.600 126.600 14.900 ;
        RECT 126.200 14.500 126.600 14.600 ;
        RECT 127.100 14.200 127.400 15.800 ;
        RECT 128.100 15.900 128.400 16.500 ;
        RECT 128.700 16.500 129.100 16.600 ;
        RECT 131.000 16.500 131.400 16.600 ;
        RECT 128.700 16.200 131.400 16.500 ;
        RECT 128.100 15.700 130.500 15.900 ;
        RECT 132.600 15.700 133.000 19.900 ;
        RECT 128.100 15.600 133.000 15.700 ;
        RECT 130.100 15.500 133.000 15.600 ;
        RECT 130.200 15.400 133.000 15.500 ;
        RECT 134.200 15.600 134.600 19.900 ;
        RECT 135.800 15.600 136.200 19.900 ;
        RECT 137.400 15.600 137.800 19.900 ;
        RECT 139.000 15.600 139.400 19.900 ;
        RECT 141.400 15.600 141.800 19.900 ;
        RECT 143.000 15.600 143.400 19.900 ;
        RECT 144.600 15.600 145.000 19.900 ;
        RECT 146.200 15.600 146.600 19.900 ;
        RECT 134.200 15.200 135.100 15.600 ;
        RECT 135.800 15.200 136.900 15.600 ;
        RECT 137.400 15.200 138.500 15.600 ;
        RECT 139.000 15.200 140.200 15.600 ;
        RECT 129.400 15.100 129.800 15.200 ;
        RECT 129.400 14.800 131.900 15.100 ;
        RECT 131.500 14.700 131.900 14.800 ;
        RECT 134.700 14.500 135.100 15.200 ;
        RECT 136.500 14.500 136.900 15.200 ;
        RECT 138.100 14.500 138.500 15.200 ;
        RECT 130.700 14.200 131.100 14.300 ;
        RECT 127.100 13.900 132.600 14.200 ;
        RECT 127.300 13.800 127.700 13.900 ;
        RECT 123.800 13.300 125.700 13.600 ;
        RECT 123.800 11.100 124.200 13.300 ;
        RECT 125.300 13.200 125.700 13.300 ;
        RECT 130.200 12.800 130.500 13.900 ;
        RECT 131.800 13.800 132.600 13.900 ;
        RECT 133.400 14.100 134.300 14.500 ;
        RECT 134.700 14.100 136.000 14.500 ;
        RECT 136.500 14.100 137.700 14.500 ;
        RECT 138.100 14.100 139.400 14.500 ;
        RECT 133.400 13.800 133.800 14.100 ;
        RECT 134.700 13.800 135.100 14.100 ;
        RECT 136.500 13.800 136.900 14.100 ;
        RECT 138.100 13.800 138.500 14.100 ;
        RECT 139.800 13.800 140.200 15.200 ;
        RECT 129.300 12.700 129.700 12.800 ;
        RECT 126.200 12.100 126.600 12.500 ;
        RECT 128.300 12.400 129.700 12.700 ;
        RECT 130.200 12.400 130.600 12.800 ;
        RECT 128.300 12.100 128.600 12.400 ;
        RECT 131.000 12.100 131.400 12.500 ;
        RECT 125.900 11.800 126.600 12.100 ;
        RECT 125.900 11.100 126.500 11.800 ;
        RECT 128.200 11.100 128.600 12.100 ;
        RECT 130.400 11.800 131.400 12.100 ;
        RECT 130.400 11.100 130.800 11.800 ;
        RECT 132.600 11.100 133.000 13.500 ;
        RECT 134.200 13.400 135.100 13.800 ;
        RECT 135.800 13.400 136.900 13.800 ;
        RECT 137.400 13.400 138.500 13.800 ;
        RECT 139.000 13.400 140.200 13.800 ;
        RECT 140.600 15.200 141.800 15.600 ;
        RECT 142.300 15.200 143.400 15.600 ;
        RECT 143.900 15.200 145.000 15.600 ;
        RECT 145.700 15.200 146.600 15.600 ;
        RECT 147.800 15.700 148.200 19.900 ;
        RECT 150.000 18.200 150.400 19.900 ;
        RECT 149.400 17.900 150.400 18.200 ;
        RECT 152.200 17.900 152.600 19.900 ;
        RECT 154.300 17.900 154.900 19.900 ;
        RECT 149.400 17.500 149.800 17.900 ;
        RECT 152.200 17.600 152.500 17.900 ;
        RECT 151.100 17.300 152.900 17.600 ;
        RECT 154.200 17.500 154.600 17.900 ;
        RECT 151.100 17.200 151.500 17.300 ;
        RECT 152.500 17.200 152.900 17.300 ;
        RECT 149.400 16.500 149.800 16.600 ;
        RECT 151.700 16.500 152.100 16.600 ;
        RECT 149.400 16.200 152.100 16.500 ;
        RECT 152.400 16.500 153.500 16.800 ;
        RECT 152.400 15.900 152.700 16.500 ;
        RECT 153.100 16.400 153.500 16.500 ;
        RECT 154.300 16.600 155.000 17.000 ;
        RECT 154.300 16.100 154.600 16.600 ;
        RECT 150.300 15.700 152.700 15.900 ;
        RECT 147.800 15.600 152.700 15.700 ;
        RECT 153.400 15.800 154.600 16.100 ;
        RECT 147.800 15.500 150.700 15.600 ;
        RECT 147.800 15.400 150.600 15.500 ;
        RECT 140.600 13.800 141.000 15.200 ;
        RECT 142.300 14.500 142.700 15.200 ;
        RECT 143.900 14.500 144.300 15.200 ;
        RECT 145.700 14.500 146.100 15.200 ;
        RECT 151.000 15.100 151.400 15.200 ;
        RECT 148.900 14.800 151.400 15.100 ;
        RECT 148.900 14.700 149.300 14.800 ;
        RECT 141.400 14.100 142.700 14.500 ;
        RECT 143.100 14.100 144.300 14.500 ;
        RECT 144.800 14.100 146.100 14.500 ;
        RECT 149.700 14.200 150.100 14.300 ;
        RECT 153.400 14.200 153.700 15.800 ;
        RECT 156.600 15.600 157.000 19.900 ;
        RECT 154.900 15.300 157.000 15.600 ;
        RECT 159.000 17.500 159.400 19.500 ;
        RECT 159.000 15.800 159.300 17.500 ;
        RECT 161.100 16.400 161.500 19.900 ;
        RECT 161.100 16.100 161.900 16.400 ;
        RECT 159.000 15.500 160.900 15.800 ;
        RECT 154.900 15.200 155.300 15.300 ;
        RECT 155.700 14.900 156.100 15.000 ;
        RECT 154.200 14.600 156.100 14.900 ;
        RECT 154.200 14.500 154.600 14.600 ;
        RECT 142.300 13.800 142.700 14.100 ;
        RECT 143.900 13.800 144.300 14.100 ;
        RECT 145.700 13.800 146.100 14.100 ;
        RECT 148.200 13.900 153.700 14.200 ;
        RECT 148.200 13.800 149.000 13.900 ;
        RECT 140.600 13.400 141.800 13.800 ;
        RECT 142.300 13.400 143.400 13.800 ;
        RECT 143.900 13.400 145.000 13.800 ;
        RECT 145.700 13.400 146.600 13.800 ;
        RECT 134.200 11.100 134.600 13.400 ;
        RECT 135.800 11.100 136.200 13.400 ;
        RECT 137.400 11.100 137.800 13.400 ;
        RECT 139.000 11.100 139.400 13.400 ;
        RECT 141.400 11.100 141.800 13.400 ;
        RECT 143.000 11.100 143.400 13.400 ;
        RECT 144.600 11.100 145.000 13.400 ;
        RECT 146.200 11.100 146.600 13.400 ;
        RECT 147.800 11.100 148.200 13.500 ;
        RECT 150.300 12.800 150.600 13.900 ;
        RECT 153.100 13.800 153.500 13.900 ;
        RECT 156.600 13.600 157.000 15.300 ;
        RECT 159.000 14.400 159.400 15.200 ;
        RECT 159.800 14.400 160.200 15.200 ;
        RECT 160.600 14.500 160.900 15.500 ;
        RECT 160.600 14.100 161.300 14.500 ;
        RECT 161.600 14.200 161.900 16.100 ;
        RECT 162.200 15.100 162.600 15.600 ;
        RECT 163.800 15.100 164.200 19.900 ;
        RECT 165.400 17.500 165.800 19.500 ;
        RECT 167.500 19.200 167.900 19.900 ;
        RECT 167.500 18.800 168.200 19.200 ;
        RECT 165.400 15.800 165.700 17.500 ;
        RECT 167.500 16.400 167.900 18.800 ;
        RECT 167.500 16.100 168.300 16.400 ;
        RECT 165.400 15.500 167.300 15.800 ;
        RECT 162.200 14.800 164.200 15.100 ;
        RECT 160.600 13.900 161.100 14.100 ;
        RECT 155.100 13.300 157.000 13.600 ;
        RECT 155.100 13.200 155.500 13.300 ;
        RECT 149.400 12.100 149.800 12.500 ;
        RECT 150.200 12.400 150.600 12.800 ;
        RECT 151.100 12.700 151.500 12.800 ;
        RECT 151.100 12.400 152.500 12.700 ;
        RECT 152.200 12.100 152.500 12.400 ;
        RECT 154.200 12.100 154.600 12.500 ;
        RECT 149.400 11.800 150.400 12.100 ;
        RECT 150.000 11.100 150.400 11.800 ;
        RECT 152.200 11.100 152.600 12.100 ;
        RECT 154.200 11.800 154.900 12.100 ;
        RECT 154.300 11.100 154.900 11.800 ;
        RECT 156.600 11.100 157.000 13.300 ;
        RECT 159.000 13.600 161.100 13.900 ;
        RECT 161.600 13.800 162.600 14.200 ;
        RECT 159.000 12.500 159.300 13.600 ;
        RECT 161.600 13.500 161.900 13.800 ;
        RECT 161.500 13.300 161.900 13.500 ;
        RECT 161.100 13.200 161.900 13.300 ;
        RECT 160.600 13.000 161.900 13.200 ;
        RECT 160.600 12.800 161.500 13.000 ;
        RECT 159.000 11.500 159.400 12.500 ;
        RECT 161.100 11.500 161.500 12.800 ;
        RECT 163.800 11.100 164.200 14.800 ;
        RECT 165.400 14.400 165.800 15.200 ;
        RECT 166.200 14.400 166.600 15.200 ;
        RECT 167.000 14.500 167.300 15.500 ;
        RECT 167.000 14.100 167.700 14.500 ;
        RECT 168.000 14.200 168.300 16.100 ;
        RECT 171.000 15.600 171.400 19.900 ;
        RECT 172.600 15.600 173.000 19.900 ;
        RECT 175.500 16.200 175.900 19.900 ;
        RECT 176.200 16.800 176.600 17.200 ;
        RECT 176.300 16.200 176.600 16.800 ;
        RECT 175.500 15.900 176.000 16.200 ;
        RECT 176.300 15.900 177.000 16.200 ;
        RECT 168.600 14.800 169.000 15.600 ;
        RECT 171.000 15.200 173.000 15.600 ;
        RECT 167.000 13.900 167.500 14.100 ;
        RECT 165.400 13.600 167.500 13.900 ;
        RECT 168.000 13.800 169.000 14.200 ;
        RECT 172.600 13.800 173.000 15.200 ;
        RECT 175.000 14.400 175.400 15.200 ;
        RECT 175.700 14.200 176.000 15.900 ;
        RECT 176.600 15.800 177.000 15.900 ;
        RECT 177.400 15.800 177.800 16.600 ;
        RECT 176.600 15.100 176.900 15.800 ;
        RECT 178.200 15.100 178.600 19.900 ;
        RECT 181.700 19.200 182.100 19.900 ;
        RECT 181.400 18.800 182.100 19.200 ;
        RECT 181.700 16.400 182.100 18.800 ;
        RECT 183.800 17.500 184.200 19.500 ;
        RECT 181.300 16.100 182.100 16.400 ;
        RECT 180.600 15.100 181.000 15.600 ;
        RECT 176.600 14.800 178.600 15.100 ;
        RECT 174.200 14.100 174.600 14.200 ;
        RECT 175.700 14.100 177.000 14.200 ;
        RECT 177.400 14.100 177.800 14.200 ;
        RECT 174.200 13.800 175.000 14.100 ;
        RECT 175.700 13.800 177.800 14.100 ;
        RECT 164.600 12.400 165.000 13.200 ;
        RECT 165.400 12.500 165.700 13.600 ;
        RECT 168.000 13.500 168.300 13.800 ;
        RECT 167.900 13.300 168.300 13.500 ;
        RECT 167.500 13.000 168.300 13.300 ;
        RECT 171.000 13.400 173.000 13.800 ;
        RECT 174.600 13.600 175.000 13.800 ;
        RECT 165.400 11.500 165.800 12.500 ;
        RECT 167.500 11.500 167.900 13.000 ;
        RECT 171.000 11.100 171.400 13.400 ;
        RECT 172.600 11.100 173.000 13.400 ;
        RECT 174.300 13.100 176.100 13.300 ;
        RECT 176.600 13.100 176.900 13.800 ;
        RECT 178.200 13.100 178.600 14.800 ;
        RECT 179.800 14.800 181.000 15.100 ;
        RECT 179.800 14.200 180.100 14.800 ;
        RECT 181.300 14.200 181.600 16.100 ;
        RECT 183.900 15.800 184.200 17.500 ;
        RECT 182.300 15.500 184.200 15.800 ;
        RECT 184.600 15.700 185.000 19.900 ;
        RECT 186.800 18.200 187.200 19.900 ;
        RECT 186.200 17.900 187.200 18.200 ;
        RECT 189.000 17.900 189.400 19.900 ;
        RECT 191.100 17.900 191.700 19.900 ;
        RECT 186.200 17.500 186.600 17.900 ;
        RECT 189.000 17.600 189.300 17.900 ;
        RECT 187.900 17.300 189.700 17.600 ;
        RECT 191.000 17.500 191.400 17.900 ;
        RECT 187.900 17.200 188.300 17.300 ;
        RECT 189.300 17.200 189.700 17.300 ;
        RECT 186.200 16.500 186.600 16.600 ;
        RECT 188.500 16.500 188.900 16.600 ;
        RECT 186.200 16.200 188.900 16.500 ;
        RECT 189.200 16.500 190.300 16.800 ;
        RECT 189.200 15.900 189.500 16.500 ;
        RECT 189.900 16.400 190.300 16.500 ;
        RECT 191.100 16.600 191.800 17.000 ;
        RECT 191.100 16.100 191.400 16.600 ;
        RECT 187.100 15.700 189.500 15.900 ;
        RECT 184.600 15.600 189.500 15.700 ;
        RECT 190.200 15.800 191.400 16.100 ;
        RECT 184.600 15.500 187.500 15.600 ;
        RECT 182.300 14.500 182.600 15.500 ;
        RECT 184.600 15.400 187.400 15.500 ;
        RECT 179.000 14.100 179.400 14.200 ;
        RECT 179.800 14.100 180.200 14.200 ;
        RECT 179.000 13.800 180.200 14.100 ;
        RECT 180.600 13.800 181.600 14.200 ;
        RECT 181.900 14.100 182.600 14.500 ;
        RECT 183.000 14.400 183.400 15.200 ;
        RECT 183.800 14.400 184.200 15.200 ;
        RECT 187.800 15.100 188.200 15.200 ;
        RECT 185.700 14.800 188.200 15.100 ;
        RECT 185.700 14.700 186.100 14.800 ;
        RECT 187.000 14.700 187.400 14.800 ;
        RECT 186.500 14.200 186.900 14.300 ;
        RECT 190.200 14.200 190.500 15.800 ;
        RECT 193.400 15.600 193.800 19.900 ;
        RECT 194.200 16.200 194.600 19.900 ;
        RECT 195.800 16.400 196.200 19.900 ;
        RECT 194.200 15.900 195.500 16.200 ;
        RECT 195.800 15.900 196.300 16.400 ;
        RECT 191.700 15.300 193.800 15.600 ;
        RECT 191.700 15.200 192.100 15.300 ;
        RECT 192.500 14.900 192.900 15.000 ;
        RECT 191.000 14.600 192.900 14.900 ;
        RECT 191.000 14.500 191.400 14.600 ;
        RECT 179.000 13.400 179.400 13.800 ;
        RECT 181.300 13.500 181.600 13.800 ;
        RECT 182.100 13.900 182.600 14.100 ;
        RECT 185.000 13.900 190.500 14.200 ;
        RECT 182.100 13.600 184.200 13.900 ;
        RECT 185.000 13.800 185.800 13.900 ;
        RECT 174.200 13.000 176.200 13.100 ;
        RECT 174.200 11.100 174.600 13.000 ;
        RECT 175.800 11.100 176.200 13.000 ;
        RECT 176.600 11.100 177.000 13.100 ;
        RECT 177.700 12.800 178.600 13.100 ;
        RECT 181.300 13.300 181.700 13.500 ;
        RECT 181.300 13.000 182.100 13.300 ;
        RECT 177.700 11.100 178.100 12.800 ;
        RECT 181.700 11.500 182.100 13.000 ;
        RECT 183.900 12.500 184.200 13.600 ;
        RECT 183.800 11.500 184.200 12.500 ;
        RECT 184.600 11.100 185.000 13.500 ;
        RECT 187.100 12.800 187.400 13.900 ;
        RECT 189.900 13.800 190.300 13.900 ;
        RECT 193.400 13.600 193.800 15.300 ;
        RECT 194.200 14.800 194.700 15.200 ;
        RECT 194.300 14.400 194.700 14.800 ;
        RECT 195.200 14.900 195.500 15.900 ;
        RECT 195.200 14.500 195.700 14.900 ;
        RECT 195.200 13.700 195.500 14.500 ;
        RECT 196.000 14.200 196.300 15.900 ;
        RECT 198.200 15.600 198.600 19.900 ;
        RECT 199.800 15.600 200.200 19.900 ;
        RECT 201.400 15.600 201.800 19.900 ;
        RECT 203.000 15.600 203.400 19.900 ;
        RECT 205.900 16.200 206.300 19.900 ;
        RECT 206.600 16.800 207.400 17.200 ;
        RECT 209.800 16.800 210.200 17.200 ;
        RECT 206.700 16.200 207.000 16.800 ;
        RECT 209.800 16.200 210.100 16.800 ;
        RECT 210.500 16.200 210.900 19.900 ;
        RECT 205.900 15.900 206.400 16.200 ;
        RECT 206.700 15.900 207.400 16.200 ;
        RECT 197.400 15.200 198.600 15.600 ;
        RECT 199.100 15.200 200.200 15.600 ;
        RECT 200.700 15.200 201.800 15.600 ;
        RECT 202.500 15.200 203.400 15.600 ;
        RECT 195.800 14.100 196.300 14.200 ;
        RECT 196.600 14.100 197.000 14.200 ;
        RECT 195.800 13.800 197.000 14.100 ;
        RECT 197.400 13.800 197.800 15.200 ;
        RECT 199.100 14.500 199.500 15.200 ;
        RECT 200.700 14.500 201.100 15.200 ;
        RECT 202.500 14.500 202.900 15.200 ;
        RECT 204.600 15.100 205.000 15.200 ;
        RECT 205.400 15.100 205.800 15.200 ;
        RECT 204.600 14.800 205.800 15.100 ;
        RECT 198.200 14.100 199.500 14.500 ;
        RECT 199.900 14.100 201.100 14.500 ;
        RECT 201.600 14.100 202.900 14.500 ;
        RECT 203.300 14.100 204.200 14.500 ;
        RECT 205.400 14.400 205.800 14.800 ;
        RECT 206.100 15.100 206.400 15.900 ;
        RECT 207.000 15.800 207.400 15.900 ;
        RECT 209.400 15.900 210.100 16.200 ;
        RECT 209.400 15.800 209.800 15.900 ;
        RECT 210.400 15.800 211.400 16.200 ;
        RECT 209.400 15.100 209.700 15.800 ;
        RECT 206.100 14.800 209.700 15.100 ;
        RECT 206.100 14.200 206.400 14.800 ;
        RECT 210.400 14.200 210.700 15.800 ;
        RECT 212.600 15.600 213.000 19.900 ;
        RECT 214.700 17.900 215.300 19.900 ;
        RECT 217.000 17.900 217.400 19.900 ;
        RECT 219.200 18.200 219.600 19.900 ;
        RECT 219.200 17.900 220.200 18.200 ;
        RECT 215.000 17.500 215.400 17.900 ;
        RECT 217.100 17.600 217.400 17.900 ;
        RECT 216.700 17.300 218.500 17.600 ;
        RECT 219.800 17.500 220.200 17.900 ;
        RECT 216.700 17.200 217.100 17.300 ;
        RECT 218.100 17.200 218.500 17.300 ;
        RECT 214.600 16.600 215.300 17.000 ;
        RECT 215.000 16.100 215.300 16.600 ;
        RECT 216.100 16.500 217.200 16.800 ;
        RECT 216.100 16.400 216.500 16.500 ;
        RECT 215.000 15.800 216.200 16.100 ;
        RECT 212.600 15.300 214.700 15.600 ;
        RECT 211.000 14.400 211.400 15.200 ;
        RECT 199.100 13.800 199.500 14.100 ;
        RECT 200.700 13.800 201.100 14.100 ;
        RECT 202.500 13.800 202.900 14.100 ;
        RECT 203.800 13.800 204.200 14.100 ;
        RECT 204.600 14.100 205.000 14.200 ;
        RECT 204.600 13.800 205.400 14.100 ;
        RECT 206.100 13.800 207.400 14.200 ;
        RECT 209.400 13.800 210.700 14.200 ;
        RECT 211.800 14.100 212.200 14.200 ;
        RECT 211.400 13.800 212.200 14.100 ;
        RECT 191.900 13.300 193.800 13.600 ;
        RECT 191.900 13.200 192.300 13.300 ;
        RECT 186.200 12.100 186.600 12.500 ;
        RECT 187.000 12.400 187.400 12.800 ;
        RECT 187.900 12.700 188.300 12.800 ;
        RECT 187.900 12.400 189.300 12.700 ;
        RECT 189.000 12.100 189.300 12.400 ;
        RECT 191.000 12.100 191.400 12.500 ;
        RECT 186.200 11.800 187.200 12.100 ;
        RECT 186.800 11.100 187.200 11.800 ;
        RECT 189.000 11.100 189.400 12.100 ;
        RECT 191.000 11.800 191.700 12.100 ;
        RECT 191.100 11.100 191.700 11.800 ;
        RECT 193.400 11.100 193.800 13.300 ;
        RECT 194.200 13.400 195.500 13.700 ;
        RECT 194.200 11.100 194.600 13.400 ;
        RECT 196.000 13.100 196.300 13.800 ;
        RECT 197.400 13.400 198.600 13.800 ;
        RECT 199.100 13.400 200.200 13.800 ;
        RECT 200.700 13.400 201.800 13.800 ;
        RECT 202.500 13.400 203.400 13.800 ;
        RECT 205.000 13.600 205.400 13.800 ;
        RECT 195.800 12.800 196.300 13.100 ;
        RECT 195.800 11.100 196.200 12.800 ;
        RECT 198.200 11.100 198.600 13.400 ;
        RECT 199.800 11.100 200.200 13.400 ;
        RECT 201.400 11.100 201.800 13.400 ;
        RECT 203.000 11.100 203.400 13.400 ;
        RECT 204.700 13.100 206.500 13.300 ;
        RECT 207.000 13.100 207.300 13.800 ;
        RECT 209.500 13.100 209.800 13.800 ;
        RECT 211.400 13.600 211.800 13.800 ;
        RECT 212.600 13.600 213.000 15.300 ;
        RECT 214.300 15.200 214.700 15.300 ;
        RECT 213.500 14.900 213.900 15.000 ;
        RECT 213.500 14.600 215.400 14.900 ;
        RECT 215.000 14.500 215.400 14.600 ;
        RECT 215.900 14.200 216.200 15.800 ;
        RECT 216.900 15.900 217.200 16.500 ;
        RECT 217.500 16.500 217.900 16.600 ;
        RECT 219.800 16.500 220.200 16.600 ;
        RECT 217.500 16.200 220.200 16.500 ;
        RECT 216.900 15.700 219.300 15.900 ;
        RECT 221.400 15.700 221.800 19.900 ;
        RECT 222.200 16.200 222.600 19.900 ;
        RECT 223.800 16.400 224.200 19.900 ;
        RECT 222.200 15.900 223.500 16.200 ;
        RECT 223.800 15.900 224.300 16.400 ;
        RECT 216.900 15.600 221.800 15.700 ;
        RECT 218.900 15.500 221.800 15.600 ;
        RECT 219.000 15.400 221.800 15.500 ;
        RECT 218.200 15.100 218.600 15.200 ;
        RECT 218.200 14.800 220.700 15.100 ;
        RECT 222.200 14.800 222.700 15.200 ;
        RECT 220.300 14.700 220.700 14.800 ;
        RECT 222.300 14.400 222.700 14.800 ;
        RECT 223.200 14.900 223.500 15.900 ;
        RECT 223.200 14.500 223.700 14.900 ;
        RECT 219.500 14.200 219.900 14.300 ;
        RECT 215.900 13.900 221.400 14.200 ;
        RECT 216.100 13.800 216.500 13.900 ;
        RECT 212.600 13.300 214.500 13.600 ;
        RECT 210.300 13.100 212.100 13.300 ;
        RECT 204.600 13.000 206.600 13.100 ;
        RECT 204.600 11.100 205.000 13.000 ;
        RECT 206.200 11.100 206.600 13.000 ;
        RECT 207.000 11.100 207.400 13.100 ;
        RECT 209.400 11.100 209.800 13.100 ;
        RECT 210.200 13.000 212.200 13.100 ;
        RECT 210.200 11.100 210.600 13.000 ;
        RECT 211.800 11.100 212.200 13.000 ;
        RECT 212.600 11.100 213.000 13.300 ;
        RECT 214.100 13.200 214.500 13.300 ;
        RECT 219.000 13.200 219.300 13.900 ;
        RECT 220.600 13.800 221.400 13.900 ;
        RECT 223.200 13.700 223.500 14.500 ;
        RECT 224.000 14.200 224.300 15.900 ;
        RECT 223.800 14.100 224.300 14.200 ;
        RECT 224.600 14.800 225.000 15.200 ;
        RECT 224.600 14.100 224.900 14.800 ;
        RECT 223.800 13.800 224.900 14.100 ;
        RECT 218.100 12.700 218.500 12.800 ;
        RECT 215.000 12.100 215.400 12.500 ;
        RECT 217.100 12.400 218.500 12.700 ;
        RECT 219.000 12.400 219.400 13.200 ;
        RECT 217.100 12.100 217.400 12.400 ;
        RECT 219.800 12.100 220.200 12.500 ;
        RECT 214.700 11.800 215.400 12.100 ;
        RECT 214.700 11.100 215.300 11.800 ;
        RECT 217.000 11.100 217.400 12.100 ;
        RECT 219.200 11.800 220.200 12.100 ;
        RECT 219.200 11.100 219.600 11.800 ;
        RECT 221.400 11.100 221.800 13.500 ;
        RECT 222.200 13.400 223.500 13.700 ;
        RECT 222.200 11.100 222.600 13.400 ;
        RECT 224.000 13.100 224.300 13.800 ;
        RECT 225.400 13.400 225.800 14.200 ;
        RECT 223.800 12.800 224.300 13.100 ;
        RECT 226.200 13.100 226.600 19.900 ;
        RECT 227.800 17.500 228.200 19.500 ;
        RECT 227.000 15.800 227.400 16.600 ;
        RECT 227.800 15.800 228.100 17.500 ;
        RECT 229.900 16.400 230.300 19.900 ;
        RECT 229.900 16.100 230.700 16.400 ;
        RECT 227.800 15.500 229.700 15.800 ;
        RECT 227.800 14.400 228.200 15.200 ;
        RECT 228.600 14.400 229.000 15.200 ;
        RECT 229.400 14.500 229.700 15.500 ;
        RECT 229.400 14.100 230.100 14.500 ;
        RECT 230.400 14.200 230.700 16.100 ;
        RECT 232.600 15.600 233.000 19.900 ;
        RECT 234.700 17.900 235.300 19.900 ;
        RECT 237.000 17.900 237.400 19.900 ;
        RECT 239.200 18.200 239.600 19.900 ;
        RECT 239.200 17.900 240.200 18.200 ;
        RECT 235.000 17.500 235.400 17.900 ;
        RECT 237.100 17.600 237.400 17.900 ;
        RECT 236.700 17.300 238.500 17.600 ;
        RECT 239.800 17.500 240.200 17.900 ;
        RECT 236.700 17.200 237.100 17.300 ;
        RECT 238.100 17.200 238.500 17.300 ;
        RECT 234.600 16.600 235.300 17.000 ;
        RECT 235.000 16.100 235.300 16.600 ;
        RECT 236.100 16.500 237.200 16.800 ;
        RECT 236.100 16.400 236.500 16.500 ;
        RECT 235.000 15.800 236.200 16.100 ;
        RECT 231.000 15.100 231.400 15.600 ;
        RECT 232.600 15.300 234.700 15.600 ;
        RECT 231.800 15.100 232.200 15.200 ;
        RECT 231.000 14.800 232.200 15.100 ;
        RECT 229.400 13.900 229.900 14.100 ;
        RECT 227.800 13.600 229.900 13.900 ;
        RECT 230.400 13.800 231.400 14.200 ;
        RECT 226.200 12.800 227.100 13.100 ;
        RECT 223.800 11.100 224.200 12.800 ;
        RECT 226.700 12.200 227.100 12.800 ;
        RECT 226.200 11.800 227.100 12.200 ;
        RECT 226.700 11.100 227.100 11.800 ;
        RECT 227.800 12.500 228.100 13.600 ;
        RECT 230.400 13.500 230.700 13.800 ;
        RECT 230.300 13.300 230.700 13.500 ;
        RECT 229.900 13.000 230.700 13.300 ;
        RECT 232.600 13.600 233.000 15.300 ;
        RECT 234.300 15.200 234.700 15.300 ;
        RECT 233.500 14.900 233.900 15.000 ;
        RECT 233.500 14.600 235.400 14.900 ;
        RECT 235.000 14.500 235.400 14.600 ;
        RECT 235.900 14.200 236.200 15.800 ;
        RECT 236.900 15.900 237.200 16.500 ;
        RECT 237.500 16.500 237.900 16.600 ;
        RECT 239.800 16.500 240.200 16.600 ;
        RECT 237.500 16.200 240.200 16.500 ;
        RECT 236.900 15.700 239.300 15.900 ;
        RECT 241.400 15.700 241.800 19.900 ;
        RECT 236.900 15.600 241.800 15.700 ;
        RECT 238.900 15.500 241.800 15.600 ;
        RECT 239.000 15.400 241.800 15.500 ;
        RECT 243.000 15.600 243.400 19.900 ;
        RECT 244.600 15.600 245.000 19.900 ;
        RECT 246.200 15.600 246.600 19.900 ;
        RECT 247.800 15.600 248.200 19.900 ;
        RECT 250.700 16.200 251.100 19.900 ;
        RECT 251.400 16.800 251.800 17.200 ;
        RECT 251.500 16.200 251.800 16.800 ;
        RECT 250.700 15.900 251.200 16.200 ;
        RECT 251.500 15.900 252.200 16.200 ;
        RECT 243.000 15.200 243.900 15.600 ;
        RECT 244.600 15.200 245.700 15.600 ;
        RECT 246.200 15.200 247.300 15.600 ;
        RECT 247.800 15.200 249.000 15.600 ;
        RECT 238.200 15.100 238.600 15.200 ;
        RECT 238.200 14.800 240.700 15.100 ;
        RECT 240.300 14.700 240.700 14.800 ;
        RECT 243.500 14.500 243.900 15.200 ;
        RECT 245.300 14.500 245.700 15.200 ;
        RECT 246.900 14.500 247.300 15.200 ;
        RECT 239.500 14.200 239.900 14.300 ;
        RECT 235.900 13.900 241.400 14.200 ;
        RECT 236.100 13.800 236.500 13.900 ;
        RECT 239.000 13.800 239.400 13.900 ;
        RECT 240.600 13.800 241.400 13.900 ;
        RECT 242.200 14.100 243.100 14.500 ;
        RECT 243.500 14.100 244.800 14.500 ;
        RECT 245.300 14.100 246.500 14.500 ;
        RECT 246.900 14.100 248.200 14.500 ;
        RECT 242.200 13.800 242.600 14.100 ;
        RECT 243.500 13.800 243.900 14.100 ;
        RECT 245.300 13.800 245.700 14.100 ;
        RECT 246.900 13.800 247.300 14.100 ;
        RECT 248.600 13.800 249.000 15.200 ;
        RECT 250.200 14.400 250.600 15.200 ;
        RECT 250.900 15.100 251.200 15.900 ;
        RECT 251.800 15.800 252.200 15.900 ;
        RECT 251.800 15.100 252.200 15.200 ;
        RECT 250.900 14.800 252.200 15.100 ;
        RECT 250.900 14.200 251.200 14.800 ;
        RECT 249.400 14.100 249.800 14.200 ;
        RECT 249.400 13.800 250.200 14.100 ;
        RECT 250.900 13.800 252.200 14.200 ;
        RECT 232.600 13.300 234.500 13.600 ;
        RECT 227.800 11.500 228.200 12.500 ;
        RECT 229.900 11.500 230.300 13.000 ;
        RECT 232.600 11.100 233.000 13.300 ;
        RECT 234.100 13.200 234.500 13.300 ;
        RECT 239.000 12.800 239.300 13.800 ;
        RECT 238.100 12.700 238.500 12.800 ;
        RECT 235.000 12.100 235.400 12.500 ;
        RECT 237.100 12.400 238.500 12.700 ;
        RECT 239.000 12.400 239.400 12.800 ;
        RECT 237.100 12.100 237.400 12.400 ;
        RECT 239.800 12.100 240.200 12.500 ;
        RECT 234.700 11.800 235.400 12.100 ;
        RECT 234.700 11.100 235.300 11.800 ;
        RECT 237.000 11.100 237.400 12.100 ;
        RECT 239.200 11.800 240.200 12.100 ;
        RECT 239.200 11.100 239.600 11.800 ;
        RECT 241.400 11.100 241.800 13.500 ;
        RECT 243.000 13.400 243.900 13.800 ;
        RECT 244.600 13.400 245.700 13.800 ;
        RECT 246.200 13.400 247.300 13.800 ;
        RECT 247.800 13.400 249.000 13.800 ;
        RECT 249.800 13.600 250.200 13.800 ;
        RECT 243.000 11.100 243.400 13.400 ;
        RECT 244.600 11.100 245.000 13.400 ;
        RECT 246.200 11.100 246.600 13.400 ;
        RECT 247.800 11.100 248.200 13.400 ;
        RECT 249.500 13.100 251.300 13.300 ;
        RECT 251.800 13.100 252.100 13.800 ;
        RECT 252.600 13.400 253.000 14.200 ;
        RECT 253.400 13.100 253.800 19.900 ;
        RECT 254.200 15.800 254.600 16.600 ;
        RECT 255.000 15.600 255.400 19.900 ;
        RECT 257.100 17.900 257.700 19.900 ;
        RECT 259.400 17.900 259.800 19.900 ;
        RECT 261.600 18.200 262.000 19.900 ;
        RECT 261.600 17.900 262.600 18.200 ;
        RECT 257.400 17.500 257.800 17.900 ;
        RECT 259.500 17.600 259.800 17.900 ;
        RECT 259.100 17.300 260.900 17.600 ;
        RECT 262.200 17.500 262.600 17.900 ;
        RECT 259.100 17.200 259.500 17.300 ;
        RECT 260.500 17.200 260.900 17.300 ;
        RECT 256.600 17.000 257.300 17.200 ;
        RECT 256.600 16.800 257.700 17.000 ;
        RECT 257.000 16.600 257.700 16.800 ;
        RECT 257.400 16.100 257.700 16.600 ;
        RECT 258.500 16.500 259.600 16.800 ;
        RECT 258.500 16.400 258.900 16.500 ;
        RECT 257.400 15.800 258.600 16.100 ;
        RECT 255.000 15.300 257.100 15.600 ;
        RECT 255.000 13.600 255.400 15.300 ;
        RECT 256.700 15.200 257.100 15.300 ;
        RECT 255.900 14.900 256.300 15.000 ;
        RECT 255.900 14.600 257.800 14.900 ;
        RECT 257.400 14.500 257.800 14.600 ;
        RECT 258.300 14.200 258.600 15.800 ;
        RECT 259.300 15.900 259.600 16.500 ;
        RECT 259.900 16.500 260.300 16.600 ;
        RECT 262.200 16.500 262.600 16.600 ;
        RECT 259.900 16.200 262.600 16.500 ;
        RECT 259.300 15.700 261.700 15.900 ;
        RECT 263.800 15.700 264.200 19.900 ;
        RECT 259.300 15.600 264.200 15.700 ;
        RECT 261.300 15.500 264.200 15.600 ;
        RECT 261.400 15.400 264.200 15.500 ;
        RECT 260.600 15.100 261.000 15.200 ;
        RECT 260.600 14.800 263.100 15.100 ;
        RECT 262.700 14.700 263.100 14.800 ;
        RECT 261.900 14.200 262.300 14.300 ;
        RECT 258.300 13.900 263.800 14.200 ;
        RECT 258.500 13.800 258.900 13.900 ;
        RECT 255.000 13.300 256.900 13.600 ;
        RECT 249.400 13.000 251.400 13.100 ;
        RECT 249.400 11.100 249.800 13.000 ;
        RECT 251.000 11.100 251.400 13.000 ;
        RECT 251.800 11.100 252.200 13.100 ;
        RECT 253.400 12.800 254.300 13.100 ;
        RECT 253.900 11.100 254.300 12.800 ;
        RECT 255.000 11.100 255.400 13.300 ;
        RECT 256.500 13.200 256.900 13.300 ;
        RECT 261.400 13.200 261.700 13.900 ;
        RECT 263.000 13.800 263.800 13.900 ;
        RECT 260.500 12.700 260.900 12.800 ;
        RECT 257.400 12.100 257.800 12.500 ;
        RECT 259.500 12.400 260.900 12.700 ;
        RECT 261.400 12.400 261.800 13.200 ;
        RECT 259.500 12.100 259.800 12.400 ;
        RECT 262.200 12.100 262.600 12.500 ;
        RECT 257.100 11.800 257.800 12.100 ;
        RECT 257.100 11.100 257.700 11.800 ;
        RECT 259.400 11.100 259.800 12.100 ;
        RECT 261.600 11.800 262.600 12.100 ;
        RECT 261.600 11.100 262.000 11.800 ;
        RECT 263.800 11.100 264.200 13.500 ;
        RECT 1.400 7.600 1.800 9.900 ;
        RECT 3.000 7.600 3.400 9.900 ;
        RECT 4.600 7.600 5.000 9.900 ;
        RECT 6.200 7.600 6.600 9.900 ;
        RECT 9.100 9.200 9.500 9.900 ;
        RECT 8.600 8.800 9.500 9.200 ;
        RECT 9.100 8.200 9.500 8.800 ;
        RECT 8.600 7.900 9.500 8.200 ;
        RECT 1.400 7.200 2.300 7.600 ;
        RECT 3.000 7.200 4.100 7.600 ;
        RECT 4.600 7.200 5.700 7.600 ;
        RECT 6.200 7.200 7.400 7.600 ;
        RECT 1.900 6.900 2.300 7.200 ;
        RECT 3.700 6.900 4.100 7.200 ;
        RECT 5.300 6.900 5.700 7.200 ;
        RECT 1.900 6.500 3.200 6.900 ;
        RECT 3.700 6.500 4.900 6.900 ;
        RECT 5.300 6.500 6.600 6.900 ;
        RECT 1.900 5.800 2.300 6.500 ;
        RECT 3.700 5.800 4.100 6.500 ;
        RECT 5.300 5.800 5.700 6.500 ;
        RECT 7.000 5.800 7.400 7.200 ;
        RECT 7.800 6.800 8.200 7.600 ;
        RECT 1.400 5.400 2.300 5.800 ;
        RECT 3.000 5.400 4.100 5.800 ;
        RECT 4.600 5.400 5.700 5.800 ;
        RECT 6.200 5.400 7.400 5.800 ;
        RECT 1.400 1.100 1.800 5.400 ;
        RECT 3.000 1.100 3.400 5.400 ;
        RECT 4.600 1.100 5.000 5.400 ;
        RECT 6.200 1.100 6.600 5.400 ;
        RECT 8.600 1.100 9.000 7.900 ;
        RECT 10.200 7.500 10.600 9.900 ;
        RECT 12.400 9.200 12.800 9.900 ;
        RECT 11.800 8.900 12.800 9.200 ;
        RECT 14.600 8.900 15.000 9.900 ;
        RECT 16.700 9.200 17.300 9.900 ;
        RECT 16.600 8.900 17.300 9.200 ;
        RECT 11.800 8.500 12.200 8.900 ;
        RECT 14.600 8.600 14.900 8.900 ;
        RECT 12.600 7.800 13.000 8.600 ;
        RECT 13.500 8.300 14.900 8.600 ;
        RECT 16.600 8.500 17.000 8.900 ;
        RECT 13.500 8.200 13.900 8.300 ;
        RECT 10.600 7.100 11.400 7.200 ;
        RECT 12.700 7.100 13.000 7.800 ;
        RECT 17.500 7.700 17.900 7.800 ;
        RECT 19.000 7.700 19.400 9.900 ;
        RECT 17.500 7.400 19.400 7.700 ;
        RECT 15.500 7.100 15.900 7.200 ;
        RECT 10.600 6.800 16.100 7.100 ;
        RECT 12.100 6.700 12.500 6.800 ;
        RECT 11.300 6.200 11.700 6.300 ;
        RECT 11.300 6.100 13.800 6.200 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 11.300 5.900 15.400 6.100 ;
        RECT 13.400 5.800 15.400 5.900 ;
        RECT 10.200 5.500 13.000 5.600 ;
        RECT 10.200 5.400 13.100 5.500 ;
        RECT 10.200 5.300 15.100 5.400 ;
        RECT 9.400 4.400 9.800 5.200 ;
        RECT 10.200 1.100 10.600 5.300 ;
        RECT 12.700 5.100 15.100 5.300 ;
        RECT 11.800 4.500 14.500 4.800 ;
        RECT 11.800 4.400 12.200 4.500 ;
        RECT 14.100 4.400 14.500 4.500 ;
        RECT 14.800 4.500 15.100 5.100 ;
        RECT 15.800 5.200 16.100 6.800 ;
        RECT 16.600 6.400 17.000 6.500 ;
        RECT 16.600 6.100 18.500 6.400 ;
        RECT 18.100 6.000 18.500 6.100 ;
        RECT 17.300 5.700 17.700 5.800 ;
        RECT 19.000 5.700 19.400 7.400 ;
        RECT 17.300 5.400 19.400 5.700 ;
        RECT 15.800 4.900 17.000 5.200 ;
        RECT 15.500 4.500 15.900 4.600 ;
        RECT 14.800 4.200 15.900 4.500 ;
        RECT 16.700 4.400 17.000 4.900 ;
        RECT 16.700 4.000 17.400 4.400 ;
        RECT 13.500 3.700 13.900 3.800 ;
        RECT 14.900 3.700 15.300 3.800 ;
        RECT 11.800 3.100 12.200 3.500 ;
        RECT 13.500 3.400 15.300 3.700 ;
        RECT 14.600 3.100 14.900 3.400 ;
        RECT 16.600 3.100 17.000 3.500 ;
        RECT 11.800 2.800 12.800 3.100 ;
        RECT 12.400 1.100 12.800 2.800 ;
        RECT 14.600 1.100 15.000 3.100 ;
        RECT 16.700 1.100 17.300 3.100 ;
        RECT 19.000 1.100 19.400 5.400 ;
        RECT 19.800 7.700 20.200 9.900 ;
        RECT 21.900 9.200 22.500 9.900 ;
        RECT 21.900 8.900 22.600 9.200 ;
        RECT 24.200 8.900 24.600 9.900 ;
        RECT 26.400 9.200 26.800 9.900 ;
        RECT 26.400 8.900 27.400 9.200 ;
        RECT 22.200 8.500 22.600 8.900 ;
        RECT 24.300 8.600 24.600 8.900 ;
        RECT 24.300 8.300 25.700 8.600 ;
        RECT 25.300 8.200 25.700 8.300 ;
        RECT 26.200 8.200 26.600 8.600 ;
        RECT 27.000 8.500 27.400 8.900 ;
        RECT 21.300 7.700 21.700 7.800 ;
        RECT 19.800 7.400 21.700 7.700 ;
        RECT 19.800 5.700 20.200 7.400 ;
        RECT 23.300 7.100 23.700 7.200 ;
        RECT 26.200 7.100 26.500 8.200 ;
        RECT 28.600 7.500 29.000 9.900 ;
        RECT 30.700 8.200 31.100 9.900 ;
        RECT 30.200 7.900 31.100 8.200 ;
        RECT 31.800 7.900 32.200 9.900 ;
        RECT 32.600 8.000 33.000 9.900 ;
        RECT 34.200 8.000 34.600 9.900 ;
        RECT 32.600 7.900 34.600 8.000 ;
        RECT 27.800 7.100 28.600 7.200 ;
        RECT 23.100 6.800 28.600 7.100 ;
        RECT 29.400 6.800 29.800 7.600 ;
        RECT 22.200 6.400 22.600 6.500 ;
        RECT 20.700 6.100 22.600 6.400 ;
        RECT 20.700 6.000 21.100 6.100 ;
        RECT 21.500 5.700 21.900 5.800 ;
        RECT 19.800 5.400 21.900 5.700 ;
        RECT 19.800 1.100 20.200 5.400 ;
        RECT 23.100 5.200 23.400 6.800 ;
        RECT 26.700 6.700 27.100 6.800 ;
        RECT 27.500 6.200 27.900 6.300 ;
        RECT 25.400 5.900 27.900 6.200 ;
        RECT 30.200 6.100 30.600 7.900 ;
        RECT 31.900 7.200 32.200 7.900 ;
        RECT 32.700 7.700 34.500 7.900 ;
        RECT 35.800 7.600 36.200 9.900 ;
        RECT 37.400 7.600 37.800 9.900 ;
        RECT 39.000 7.600 39.400 9.900 ;
        RECT 40.600 7.600 41.000 9.900 ;
        RECT 33.800 7.200 34.200 7.400 ;
        RECT 35.000 7.200 36.200 7.600 ;
        RECT 36.700 7.200 37.800 7.600 ;
        RECT 38.300 7.200 39.400 7.600 ;
        RECT 40.100 7.200 41.000 7.600 ;
        RECT 43.000 7.600 43.400 9.900 ;
        RECT 44.600 7.600 45.000 9.900 ;
        RECT 46.200 7.600 46.600 9.900 ;
        RECT 47.800 7.600 48.200 9.900 ;
        RECT 50.200 7.600 50.600 9.900 ;
        RECT 51.800 7.600 52.200 9.900 ;
        RECT 53.400 7.600 53.800 9.900 ;
        RECT 55.000 7.600 55.400 9.900 ;
        RECT 43.000 7.200 43.900 7.600 ;
        RECT 44.600 7.200 45.700 7.600 ;
        RECT 46.200 7.200 47.300 7.600 ;
        RECT 47.800 7.200 49.000 7.600 ;
        RECT 31.000 7.100 31.400 7.200 ;
        RECT 31.800 7.100 33.100 7.200 ;
        RECT 31.000 6.800 33.100 7.100 ;
        RECT 33.800 6.900 34.600 7.200 ;
        RECT 34.200 6.800 34.600 6.900 ;
        RECT 25.400 5.800 25.800 5.900 ;
        RECT 30.200 5.800 32.100 6.100 ;
        RECT 26.200 5.500 29.000 5.600 ;
        RECT 26.100 5.400 29.000 5.500 ;
        RECT 22.200 4.900 23.400 5.200 ;
        RECT 24.100 5.300 29.000 5.400 ;
        RECT 24.100 5.100 26.500 5.300 ;
        RECT 22.200 4.400 22.500 4.900 ;
        RECT 21.800 4.000 22.500 4.400 ;
        RECT 23.300 4.500 23.700 4.600 ;
        RECT 24.100 4.500 24.400 5.100 ;
        RECT 23.300 4.200 24.400 4.500 ;
        RECT 24.700 4.500 27.400 4.800 ;
        RECT 24.700 4.400 25.100 4.500 ;
        RECT 27.000 4.400 27.400 4.500 ;
        RECT 23.900 3.700 24.300 3.800 ;
        RECT 25.300 3.700 25.700 3.800 ;
        RECT 22.200 3.100 22.600 3.500 ;
        RECT 23.900 3.400 25.700 3.700 ;
        RECT 24.300 3.100 24.600 3.400 ;
        RECT 27.000 3.100 27.400 3.500 ;
        RECT 21.900 1.100 22.500 3.100 ;
        RECT 24.200 1.100 24.600 3.100 ;
        RECT 26.400 2.800 27.400 3.100 ;
        RECT 26.400 1.100 26.800 2.800 ;
        RECT 28.600 1.100 29.000 5.300 ;
        RECT 30.200 1.100 30.600 5.800 ;
        RECT 31.800 5.200 32.100 5.800 ;
        RECT 31.000 4.400 31.400 5.200 ;
        RECT 31.800 5.100 32.200 5.200 ;
        RECT 32.800 5.100 33.100 6.800 ;
        RECT 33.400 5.800 33.800 6.600 ;
        RECT 35.000 5.800 35.400 7.200 ;
        RECT 36.700 6.900 37.100 7.200 ;
        RECT 38.300 6.900 38.700 7.200 ;
        RECT 40.100 6.900 40.500 7.200 ;
        RECT 41.400 6.900 41.800 7.200 ;
        RECT 35.800 6.500 37.100 6.900 ;
        RECT 37.500 6.500 38.700 6.900 ;
        RECT 39.200 6.500 40.500 6.900 ;
        RECT 40.900 6.500 41.800 6.900 ;
        RECT 43.500 6.900 43.900 7.200 ;
        RECT 45.300 6.900 45.700 7.200 ;
        RECT 46.900 6.900 47.300 7.200 ;
        RECT 43.500 6.500 44.800 6.900 ;
        RECT 45.300 6.500 46.500 6.900 ;
        RECT 46.900 6.500 48.200 6.900 ;
        RECT 36.700 5.800 37.100 6.500 ;
        RECT 38.300 5.800 38.700 6.500 ;
        RECT 40.100 5.800 40.500 6.500 ;
        RECT 43.500 5.800 43.900 6.500 ;
        RECT 45.300 5.800 45.700 6.500 ;
        RECT 46.900 5.800 47.300 6.500 ;
        RECT 48.600 5.800 49.000 7.200 ;
        RECT 35.000 5.400 36.200 5.800 ;
        RECT 36.700 5.400 37.800 5.800 ;
        RECT 38.300 5.400 39.400 5.800 ;
        RECT 40.100 5.400 41.000 5.800 ;
        RECT 31.800 4.800 32.500 5.100 ;
        RECT 32.800 4.800 33.300 5.100 ;
        RECT 32.200 4.200 32.500 4.800 ;
        RECT 32.200 3.800 32.600 4.200 ;
        RECT 32.900 1.100 33.300 4.800 ;
        RECT 35.800 1.100 36.200 5.400 ;
        RECT 37.400 1.100 37.800 5.400 ;
        RECT 39.000 1.100 39.400 5.400 ;
        RECT 40.600 1.100 41.000 5.400 ;
        RECT 43.000 5.400 43.900 5.800 ;
        RECT 44.600 5.400 45.700 5.800 ;
        RECT 46.200 5.400 47.300 5.800 ;
        RECT 47.800 5.400 49.000 5.800 ;
        RECT 49.400 7.200 50.600 7.600 ;
        RECT 51.100 7.200 52.200 7.600 ;
        RECT 52.700 7.200 53.800 7.600 ;
        RECT 54.500 7.200 55.400 7.600 ;
        RECT 59.000 7.600 59.400 9.900 ;
        RECT 60.600 7.600 61.000 9.900 ;
        RECT 62.200 7.600 62.600 9.900 ;
        RECT 63.800 7.600 64.200 9.900 ;
        RECT 65.400 8.500 65.800 9.500 ;
        RECT 59.000 7.200 59.900 7.600 ;
        RECT 60.600 7.200 61.700 7.600 ;
        RECT 62.200 7.200 63.300 7.600 ;
        RECT 63.800 7.200 65.000 7.600 ;
        RECT 49.400 5.800 49.800 7.200 ;
        RECT 51.100 6.900 51.500 7.200 ;
        RECT 52.700 6.900 53.100 7.200 ;
        RECT 54.500 6.900 54.900 7.200 ;
        RECT 55.800 7.100 56.200 7.200 ;
        RECT 58.200 7.100 58.600 7.200 ;
        RECT 55.800 6.900 58.600 7.100 ;
        RECT 59.500 6.900 59.900 7.200 ;
        RECT 61.300 6.900 61.700 7.200 ;
        RECT 62.900 6.900 63.300 7.200 ;
        RECT 50.200 6.500 51.500 6.900 ;
        RECT 51.900 6.500 53.100 6.900 ;
        RECT 53.600 6.500 54.900 6.900 ;
        RECT 55.300 6.800 59.100 6.900 ;
        RECT 55.300 6.500 56.200 6.800 ;
        RECT 58.200 6.500 59.100 6.800 ;
        RECT 59.500 6.500 60.800 6.900 ;
        RECT 61.300 6.500 62.500 6.900 ;
        RECT 62.900 6.500 64.200 6.900 ;
        RECT 51.100 5.800 51.500 6.500 ;
        RECT 52.700 5.800 53.100 6.500 ;
        RECT 54.500 5.800 54.900 6.500 ;
        RECT 55.800 6.200 56.100 6.500 ;
        RECT 55.800 5.800 56.200 6.200 ;
        RECT 59.500 5.800 59.900 6.500 ;
        RECT 61.300 5.800 61.700 6.500 ;
        RECT 62.900 5.800 63.300 6.500 ;
        RECT 64.600 5.800 65.000 7.200 ;
        RECT 65.400 7.400 65.700 8.500 ;
        RECT 67.500 8.000 67.900 9.500 ;
        RECT 67.500 7.700 68.300 8.000 ;
        RECT 67.900 7.500 68.300 7.700 ;
        RECT 65.400 7.100 67.500 7.400 ;
        RECT 67.000 6.900 67.500 7.100 ;
        RECT 68.000 7.200 68.300 7.500 ;
        RECT 68.000 7.100 69.000 7.200 ;
        RECT 69.400 7.100 69.800 7.200 ;
        RECT 65.400 5.800 65.800 6.600 ;
        RECT 66.200 5.800 66.600 6.600 ;
        RECT 67.000 6.500 67.700 6.900 ;
        RECT 68.000 6.800 69.800 7.100 ;
        RECT 49.400 5.400 50.600 5.800 ;
        RECT 51.100 5.400 52.200 5.800 ;
        RECT 52.700 5.400 53.800 5.800 ;
        RECT 54.500 5.400 55.400 5.800 ;
        RECT 43.000 1.100 43.400 5.400 ;
        RECT 44.600 1.100 45.000 5.400 ;
        RECT 46.200 1.100 46.600 5.400 ;
        RECT 47.800 1.100 48.200 5.400 ;
        RECT 50.200 1.100 50.600 5.400 ;
        RECT 51.800 1.100 52.200 5.400 ;
        RECT 53.400 1.100 53.800 5.400 ;
        RECT 55.000 1.100 55.400 5.400 ;
        RECT 59.000 5.400 59.900 5.800 ;
        RECT 60.600 5.400 61.700 5.800 ;
        RECT 62.200 5.400 63.300 5.800 ;
        RECT 63.800 5.400 65.000 5.800 ;
        RECT 67.000 5.500 67.300 6.500 ;
        RECT 59.000 1.100 59.400 5.400 ;
        RECT 60.600 1.100 61.000 5.400 ;
        RECT 62.200 1.100 62.600 5.400 ;
        RECT 63.800 1.100 64.200 5.400 ;
        RECT 65.400 5.200 67.300 5.500 ;
        RECT 65.400 3.500 65.700 5.200 ;
        RECT 68.000 4.900 68.300 6.800 ;
        RECT 68.600 6.100 69.000 6.200 ;
        RECT 70.200 6.100 70.600 9.900 ;
        RECT 71.000 7.800 71.400 8.600 ;
        RECT 71.800 7.500 72.200 9.900 ;
        RECT 74.000 9.200 74.400 9.900 ;
        RECT 73.400 8.900 74.400 9.200 ;
        RECT 76.200 8.900 76.600 9.900 ;
        RECT 78.300 9.200 78.900 9.900 ;
        RECT 78.200 8.900 78.900 9.200 ;
        RECT 73.400 8.500 73.800 8.900 ;
        RECT 76.200 8.600 76.500 8.900 ;
        RECT 74.200 8.200 74.600 8.600 ;
        RECT 75.100 8.300 76.500 8.600 ;
        RECT 78.200 8.500 78.600 8.900 ;
        RECT 75.100 8.200 75.500 8.300 ;
        RECT 72.200 7.100 73.000 7.200 ;
        RECT 74.300 7.100 74.600 8.200 ;
        RECT 79.100 7.700 79.500 7.800 ;
        RECT 80.600 7.700 81.000 9.900 ;
        RECT 79.100 7.400 81.000 7.700 ;
        RECT 77.100 7.100 77.500 7.200 ;
        RECT 72.200 6.800 77.700 7.100 ;
        RECT 73.700 6.700 74.100 6.800 ;
        RECT 68.600 5.800 70.600 6.100 ;
        RECT 72.900 6.200 73.300 6.300 ;
        RECT 74.200 6.200 74.600 6.300 ;
        RECT 72.900 5.900 75.400 6.200 ;
        RECT 75.000 5.800 75.400 5.900 ;
        RECT 68.600 5.400 69.000 5.800 ;
        RECT 67.500 4.600 68.300 4.900 ;
        RECT 65.400 1.500 65.800 3.500 ;
        RECT 67.500 1.100 67.900 4.600 ;
        RECT 70.200 1.100 70.600 5.800 ;
        RECT 71.800 5.500 74.600 5.600 ;
        RECT 71.800 5.400 74.700 5.500 ;
        RECT 71.800 5.300 76.700 5.400 ;
        RECT 71.800 1.100 72.200 5.300 ;
        RECT 74.300 5.100 76.700 5.300 ;
        RECT 73.400 4.500 76.100 4.800 ;
        RECT 73.400 4.400 73.800 4.500 ;
        RECT 75.700 4.400 76.100 4.500 ;
        RECT 76.400 4.500 76.700 5.100 ;
        RECT 77.400 5.200 77.700 6.800 ;
        RECT 78.200 6.400 78.600 6.500 ;
        RECT 78.200 6.100 80.100 6.400 ;
        RECT 79.700 6.000 80.100 6.100 ;
        RECT 78.900 5.700 79.300 5.800 ;
        RECT 80.600 5.700 81.000 7.400 ;
        RECT 78.900 5.400 81.000 5.700 ;
        RECT 77.400 4.900 78.600 5.200 ;
        RECT 77.100 4.500 77.500 4.600 ;
        RECT 76.400 4.200 77.500 4.500 ;
        RECT 78.300 4.400 78.600 4.900 ;
        RECT 78.300 4.000 79.000 4.400 ;
        RECT 75.100 3.700 75.500 3.800 ;
        RECT 76.500 3.700 76.900 3.800 ;
        RECT 73.400 3.100 73.800 3.500 ;
        RECT 75.100 3.400 76.900 3.700 ;
        RECT 76.200 3.100 76.500 3.400 ;
        RECT 78.200 3.100 78.600 3.500 ;
        RECT 73.400 2.800 74.400 3.100 ;
        RECT 74.000 1.100 74.400 2.800 ;
        RECT 76.200 1.100 76.600 3.100 ;
        RECT 78.300 1.100 78.900 3.100 ;
        RECT 80.600 1.100 81.000 5.400 ;
        RECT 81.400 7.700 81.800 9.900 ;
        RECT 83.500 9.200 84.100 9.900 ;
        RECT 83.500 8.900 84.200 9.200 ;
        RECT 85.800 8.900 86.200 9.900 ;
        RECT 88.000 9.200 88.400 9.900 ;
        RECT 88.000 8.900 89.000 9.200 ;
        RECT 83.800 8.500 84.200 8.900 ;
        RECT 85.900 8.600 86.200 8.900 ;
        RECT 85.900 8.300 87.300 8.600 ;
        RECT 86.900 8.200 87.300 8.300 ;
        RECT 87.800 8.200 88.200 8.600 ;
        RECT 88.600 8.500 89.000 8.900 ;
        RECT 82.900 7.700 83.300 7.800 ;
        RECT 81.400 7.400 83.300 7.700 ;
        RECT 81.400 5.700 81.800 7.400 ;
        RECT 84.900 7.100 85.300 7.200 ;
        RECT 87.000 7.100 87.400 7.200 ;
        RECT 87.800 7.100 88.100 8.200 ;
        RECT 90.200 7.500 90.600 9.900 ;
        RECT 92.300 8.200 92.700 9.900 ;
        RECT 91.800 7.900 92.700 8.200 ;
        RECT 93.400 7.900 93.800 9.900 ;
        RECT 94.200 8.000 94.600 9.900 ;
        RECT 95.800 8.000 96.200 9.900 ;
        RECT 94.200 7.900 96.200 8.000 ;
        RECT 89.400 7.100 90.200 7.200 ;
        RECT 84.700 6.800 90.200 7.100 ;
        RECT 91.000 6.800 91.400 7.600 ;
        RECT 83.800 6.400 84.200 6.500 ;
        RECT 82.300 6.100 84.200 6.400 ;
        RECT 82.300 6.000 82.700 6.100 ;
        RECT 83.100 5.700 83.500 5.800 ;
        RECT 81.400 5.400 83.500 5.700 ;
        RECT 81.400 1.100 81.800 5.400 ;
        RECT 84.700 5.200 85.000 6.800 ;
        RECT 88.300 6.700 88.700 6.800 ;
        RECT 87.800 6.200 88.200 6.300 ;
        RECT 89.100 6.200 89.500 6.300 ;
        RECT 87.000 5.900 89.500 6.200 ;
        RECT 91.800 6.100 92.200 7.900 ;
        RECT 93.500 7.200 93.800 7.900 ;
        RECT 94.300 7.700 96.100 7.900 ;
        RECT 96.600 7.500 97.000 9.900 ;
        RECT 98.800 9.200 99.200 9.900 ;
        RECT 98.200 8.900 99.200 9.200 ;
        RECT 101.000 8.900 101.400 9.900 ;
        RECT 103.100 9.200 103.700 9.900 ;
        RECT 103.000 8.900 103.700 9.200 ;
        RECT 105.400 9.100 105.800 9.900 ;
        RECT 98.200 8.500 98.600 8.900 ;
        RECT 101.000 8.600 101.300 8.900 ;
        RECT 99.000 8.200 99.400 8.600 ;
        RECT 99.900 8.300 101.300 8.600 ;
        RECT 103.000 8.500 103.400 8.900 ;
        RECT 105.400 8.800 106.500 9.100 ;
        RECT 99.900 8.200 100.300 8.300 ;
        RECT 95.400 7.200 95.800 7.400 ;
        RECT 92.600 7.100 93.000 7.200 ;
        RECT 93.400 7.100 94.700 7.200 ;
        RECT 92.600 6.800 94.700 7.100 ;
        RECT 95.400 6.900 96.200 7.200 ;
        RECT 95.800 6.800 96.200 6.900 ;
        RECT 97.000 7.100 97.800 7.200 ;
        RECT 99.100 7.100 99.400 8.200 ;
        RECT 103.900 7.700 104.300 7.800 ;
        RECT 105.400 7.700 105.800 8.800 ;
        RECT 106.200 8.100 106.500 8.800 ;
        RECT 107.800 8.100 108.200 8.600 ;
        RECT 106.200 7.800 108.200 8.100 ;
        RECT 103.900 7.400 105.800 7.700 ;
        RECT 101.900 7.100 102.300 7.200 ;
        RECT 97.000 6.800 102.500 7.100 ;
        RECT 87.000 5.800 87.400 5.900 ;
        RECT 91.800 5.800 93.700 6.100 ;
        RECT 87.800 5.500 90.600 5.600 ;
        RECT 87.700 5.400 90.600 5.500 ;
        RECT 83.800 4.900 85.000 5.200 ;
        RECT 85.700 5.300 90.600 5.400 ;
        RECT 85.700 5.100 88.100 5.300 ;
        RECT 83.800 4.400 84.100 4.900 ;
        RECT 83.400 4.000 84.100 4.400 ;
        RECT 84.900 4.500 85.300 4.600 ;
        RECT 85.700 4.500 86.000 5.100 ;
        RECT 84.900 4.200 86.000 4.500 ;
        RECT 86.300 4.500 89.000 4.800 ;
        RECT 86.300 4.400 86.700 4.500 ;
        RECT 88.600 4.400 89.000 4.500 ;
        RECT 85.500 3.700 85.900 3.800 ;
        RECT 86.900 3.700 87.300 3.800 ;
        RECT 83.800 3.100 84.200 3.500 ;
        RECT 85.500 3.400 87.300 3.700 ;
        RECT 85.900 3.100 86.200 3.400 ;
        RECT 88.600 3.100 89.000 3.500 ;
        RECT 83.500 1.100 84.100 3.100 ;
        RECT 85.800 1.100 86.200 3.100 ;
        RECT 88.000 2.800 89.000 3.100 ;
        RECT 88.000 1.100 88.400 2.800 ;
        RECT 90.200 1.100 90.600 5.300 ;
        RECT 91.800 1.100 92.200 5.800 ;
        RECT 93.400 5.200 93.700 5.800 ;
        RECT 92.600 4.400 93.000 5.200 ;
        RECT 93.400 5.100 93.800 5.200 ;
        RECT 94.400 5.100 94.700 6.800 ;
        RECT 98.500 6.700 98.900 6.800 ;
        RECT 95.000 5.800 95.400 6.600 ;
        RECT 97.700 6.200 98.100 6.300 ;
        RECT 97.700 6.100 100.200 6.200 ;
        RECT 101.400 6.100 101.800 6.200 ;
        RECT 97.700 5.900 101.800 6.100 ;
        RECT 99.800 5.800 101.800 5.900 ;
        RECT 96.600 5.500 99.400 5.600 ;
        RECT 96.600 5.400 99.500 5.500 ;
        RECT 96.600 5.300 101.500 5.400 ;
        RECT 93.400 4.800 94.100 5.100 ;
        RECT 94.400 4.800 94.900 5.100 ;
        RECT 93.800 4.200 94.100 4.800 ;
        RECT 93.800 3.800 94.200 4.200 ;
        RECT 94.500 1.100 94.900 4.800 ;
        RECT 96.600 1.100 97.000 5.300 ;
        RECT 99.100 5.100 101.500 5.300 ;
        RECT 98.200 4.500 100.900 4.800 ;
        RECT 98.200 4.400 98.600 4.500 ;
        RECT 100.500 4.400 100.900 4.500 ;
        RECT 101.200 4.500 101.500 5.100 ;
        RECT 102.200 5.200 102.500 6.800 ;
        RECT 103.000 6.400 103.400 6.500 ;
        RECT 103.000 6.100 104.900 6.400 ;
        RECT 104.500 6.000 104.900 6.100 ;
        RECT 103.700 5.700 104.100 5.800 ;
        RECT 105.400 5.700 105.800 7.400 ;
        RECT 103.700 5.400 105.800 5.700 ;
        RECT 102.200 4.900 103.400 5.200 ;
        RECT 101.900 4.500 102.300 4.600 ;
        RECT 101.200 4.200 102.300 4.500 ;
        RECT 103.100 4.400 103.400 4.900 ;
        RECT 103.100 4.000 103.800 4.400 ;
        RECT 99.900 3.700 100.300 3.800 ;
        RECT 101.300 3.700 101.700 3.800 ;
        RECT 98.200 3.100 98.600 3.500 ;
        RECT 99.900 3.400 101.700 3.700 ;
        RECT 101.000 3.100 101.300 3.400 ;
        RECT 103.000 3.100 103.400 3.500 ;
        RECT 98.200 2.800 99.200 3.100 ;
        RECT 98.800 1.100 99.200 2.800 ;
        RECT 101.000 1.100 101.400 3.100 ;
        RECT 103.100 1.100 103.700 3.100 ;
        RECT 105.400 1.100 105.800 5.400 ;
        RECT 108.600 6.100 109.000 9.900 ;
        RECT 111.300 8.000 111.700 9.500 ;
        RECT 113.400 8.500 113.800 9.500 ;
        RECT 110.900 7.700 111.700 8.000 ;
        RECT 110.900 7.500 111.300 7.700 ;
        RECT 110.900 7.200 111.200 7.500 ;
        RECT 113.500 7.400 113.800 8.500 ;
        RECT 114.200 8.000 114.600 9.900 ;
        RECT 115.800 8.000 116.200 9.900 ;
        RECT 114.200 7.900 116.200 8.000 ;
        RECT 116.600 7.900 117.000 9.900 ;
        RECT 117.700 8.200 118.100 9.900 ;
        RECT 117.700 7.900 118.600 8.200 ;
        RECT 114.300 7.700 116.100 7.900 ;
        RECT 110.200 6.800 111.200 7.200 ;
        RECT 111.700 7.100 113.800 7.400 ;
        RECT 114.600 7.200 115.000 7.400 ;
        RECT 116.600 7.200 116.900 7.900 ;
        RECT 111.700 6.900 112.200 7.100 ;
        RECT 110.200 6.100 110.600 6.200 ;
        RECT 108.600 5.800 110.600 6.100 ;
        RECT 108.600 1.100 109.000 5.800 ;
        RECT 110.200 5.400 110.600 5.800 ;
        RECT 110.900 4.900 111.200 6.800 ;
        RECT 111.500 6.500 112.200 6.900 ;
        RECT 114.200 6.900 115.000 7.200 ;
        RECT 115.700 7.100 117.000 7.200 ;
        RECT 117.400 7.100 117.800 7.200 ;
        RECT 114.200 6.800 114.600 6.900 ;
        RECT 115.700 6.800 117.800 7.100 ;
        RECT 111.900 5.500 112.200 6.500 ;
        RECT 112.600 5.800 113.000 6.600 ;
        RECT 113.400 5.800 113.800 6.600 ;
        RECT 115.000 5.800 115.400 6.600 ;
        RECT 111.900 5.200 113.800 5.500 ;
        RECT 110.900 4.600 111.700 4.900 ;
        RECT 111.300 1.100 111.700 4.600 ;
        RECT 113.500 3.500 113.800 5.200 ;
        RECT 115.700 5.100 116.000 6.800 ;
        RECT 118.200 6.100 118.600 7.900 ;
        RECT 119.800 7.700 120.200 9.900 ;
        RECT 121.900 9.200 122.500 9.900 ;
        RECT 121.900 8.900 122.600 9.200 ;
        RECT 124.200 8.900 124.600 9.900 ;
        RECT 126.400 9.200 126.800 9.900 ;
        RECT 126.400 8.900 127.400 9.200 ;
        RECT 122.200 8.500 122.600 8.900 ;
        RECT 124.300 8.600 124.600 8.900 ;
        RECT 124.300 8.300 125.700 8.600 ;
        RECT 125.300 8.200 125.700 8.300 ;
        RECT 126.200 8.200 126.600 8.600 ;
        RECT 127.000 8.500 127.400 8.900 ;
        RECT 121.300 7.700 121.700 7.800 ;
        RECT 119.000 7.100 119.400 7.600 ;
        RECT 119.800 7.400 121.700 7.700 ;
        RECT 119.800 7.100 120.200 7.400 ;
        RECT 123.300 7.100 123.700 7.200 ;
        RECT 126.200 7.100 126.500 8.200 ;
        RECT 128.600 7.500 129.000 9.900 ;
        RECT 130.700 8.200 131.100 9.900 ;
        RECT 130.200 7.900 131.100 8.200 ;
        RECT 131.800 7.900 132.200 9.900 ;
        RECT 132.600 8.000 133.000 9.900 ;
        RECT 134.200 8.000 134.600 9.900 ;
        RECT 132.600 7.900 134.600 8.000 ;
        RECT 127.800 7.100 128.600 7.200 ;
        RECT 119.000 6.800 120.200 7.100 ;
        RECT 116.600 5.800 118.600 6.100 ;
        RECT 116.600 5.200 116.900 5.800 ;
        RECT 116.600 5.100 117.000 5.200 ;
        RECT 113.400 1.500 113.800 3.500 ;
        RECT 115.500 4.800 116.000 5.100 ;
        RECT 116.300 4.800 117.000 5.100 ;
        RECT 115.500 1.100 115.900 4.800 ;
        RECT 116.300 4.200 116.600 4.800 ;
        RECT 117.400 4.400 117.800 5.200 ;
        RECT 116.200 3.800 116.600 4.200 ;
        RECT 118.200 1.100 118.600 5.800 ;
        RECT 119.800 5.700 120.200 6.800 ;
        RECT 123.100 6.800 128.600 7.100 ;
        RECT 129.400 6.800 129.800 7.600 ;
        RECT 122.200 6.400 122.600 6.500 ;
        RECT 120.700 6.100 122.600 6.400 ;
        RECT 120.700 6.000 121.100 6.100 ;
        RECT 121.500 5.700 121.900 5.800 ;
        RECT 119.800 5.400 121.900 5.700 ;
        RECT 119.800 1.100 120.200 5.400 ;
        RECT 123.100 5.200 123.400 6.800 ;
        RECT 126.700 6.700 127.100 6.800 ;
        RECT 127.500 6.200 127.900 6.300 ;
        RECT 125.400 5.900 127.900 6.200 ;
        RECT 130.200 6.100 130.600 7.900 ;
        RECT 131.900 7.200 132.200 7.900 ;
        RECT 132.700 7.700 134.500 7.900 ;
        RECT 135.000 7.700 135.400 9.900 ;
        RECT 137.100 9.200 137.700 9.900 ;
        RECT 137.100 8.900 137.800 9.200 ;
        RECT 139.400 8.900 139.800 9.900 ;
        RECT 141.600 9.200 142.000 9.900 ;
        RECT 141.600 8.900 142.600 9.200 ;
        RECT 137.400 8.500 137.800 8.900 ;
        RECT 139.500 8.600 139.800 8.900 ;
        RECT 139.500 8.300 140.900 8.600 ;
        RECT 140.500 8.200 140.900 8.300 ;
        RECT 141.400 8.200 141.800 8.600 ;
        RECT 142.200 8.500 142.600 8.900 ;
        RECT 136.500 7.700 136.900 7.800 ;
        RECT 135.000 7.400 136.900 7.700 ;
        RECT 133.800 7.200 134.200 7.400 ;
        RECT 131.800 6.800 133.100 7.200 ;
        RECT 133.800 6.900 134.600 7.200 ;
        RECT 134.200 6.800 134.600 6.900 ;
        RECT 132.800 6.200 133.100 6.800 ;
        RECT 125.400 5.800 125.800 5.900 ;
        RECT 130.200 5.800 132.100 6.100 ;
        RECT 132.600 5.800 133.100 6.200 ;
        RECT 133.400 5.800 133.800 6.600 ;
        RECT 126.200 5.500 129.000 5.600 ;
        RECT 126.100 5.400 129.000 5.500 ;
        RECT 122.200 4.900 123.400 5.200 ;
        RECT 124.100 5.300 129.000 5.400 ;
        RECT 124.100 5.100 126.500 5.300 ;
        RECT 122.200 4.400 122.500 4.900 ;
        RECT 121.800 4.000 122.500 4.400 ;
        RECT 123.300 4.500 123.700 4.600 ;
        RECT 124.100 4.500 124.400 5.100 ;
        RECT 123.300 4.200 124.400 4.500 ;
        RECT 124.700 4.500 127.400 4.800 ;
        RECT 124.700 4.400 125.100 4.500 ;
        RECT 127.000 4.400 127.400 4.500 ;
        RECT 123.900 3.700 124.300 3.800 ;
        RECT 125.300 3.700 125.700 3.800 ;
        RECT 122.200 3.100 122.600 3.500 ;
        RECT 123.900 3.400 125.700 3.700 ;
        RECT 124.300 3.100 124.600 3.400 ;
        RECT 127.000 3.100 127.400 3.500 ;
        RECT 121.900 1.100 122.500 3.100 ;
        RECT 124.200 1.100 124.600 3.100 ;
        RECT 126.400 2.800 127.400 3.100 ;
        RECT 126.400 1.100 126.800 2.800 ;
        RECT 128.600 1.100 129.000 5.300 ;
        RECT 130.200 1.100 130.600 5.800 ;
        RECT 131.800 5.200 132.100 5.800 ;
        RECT 131.000 4.400 131.400 5.200 ;
        RECT 131.800 5.100 132.200 5.200 ;
        RECT 132.800 5.100 133.100 5.800 ;
        RECT 135.000 5.700 135.400 7.400 ;
        RECT 138.500 7.100 138.900 7.200 ;
        RECT 141.400 7.100 141.700 8.200 ;
        RECT 143.800 7.500 144.200 9.900 ;
        RECT 145.400 7.600 145.800 9.900 ;
        RECT 147.000 7.600 147.400 9.900 ;
        RECT 148.600 7.600 149.000 9.900 ;
        RECT 150.200 7.600 150.600 9.900 ;
        RECT 152.600 8.200 153.000 9.900 ;
        RECT 152.500 7.900 153.000 8.200 ;
        RECT 145.400 7.200 146.300 7.600 ;
        RECT 147.000 7.200 148.100 7.600 ;
        RECT 148.600 7.200 149.700 7.600 ;
        RECT 150.200 7.200 151.400 7.600 ;
        RECT 143.000 7.100 143.800 7.200 ;
        RECT 138.300 6.800 143.800 7.100 ;
        RECT 144.600 6.900 145.000 7.200 ;
        RECT 145.900 6.900 146.300 7.200 ;
        RECT 147.700 6.900 148.100 7.200 ;
        RECT 149.300 6.900 149.700 7.200 ;
        RECT 137.400 6.400 137.800 6.500 ;
        RECT 135.900 6.100 137.800 6.400 ;
        RECT 135.900 6.000 136.300 6.100 ;
        RECT 136.700 5.700 137.100 5.800 ;
        RECT 135.000 5.400 137.100 5.700 ;
        RECT 131.800 4.800 132.500 5.100 ;
        RECT 132.800 4.800 133.300 5.100 ;
        RECT 132.200 4.200 132.500 4.800 ;
        RECT 132.200 3.800 132.600 4.200 ;
        RECT 132.900 1.100 133.300 4.800 ;
        RECT 135.000 1.100 135.400 5.400 ;
        RECT 138.300 5.200 138.600 6.800 ;
        RECT 141.900 6.700 142.300 6.800 ;
        RECT 144.600 6.500 145.500 6.900 ;
        RECT 145.900 6.500 147.200 6.900 ;
        RECT 147.700 6.500 148.900 6.900 ;
        RECT 149.300 6.500 150.600 6.900 ;
        RECT 142.700 6.200 143.100 6.300 ;
        RECT 139.000 6.100 139.400 6.200 ;
        RECT 140.600 6.100 143.100 6.200 ;
        RECT 139.000 5.900 143.100 6.100 ;
        RECT 139.000 5.800 141.000 5.900 ;
        RECT 145.900 5.800 146.300 6.500 ;
        RECT 147.700 5.800 148.100 6.500 ;
        RECT 149.300 5.800 149.700 6.500 ;
        RECT 151.000 5.800 151.400 7.200 ;
        RECT 141.400 5.500 144.200 5.600 ;
        RECT 141.300 5.400 144.200 5.500 ;
        RECT 137.400 4.900 138.600 5.200 ;
        RECT 139.300 5.300 144.200 5.400 ;
        RECT 139.300 5.100 141.700 5.300 ;
        RECT 137.400 4.400 137.700 4.900 ;
        RECT 137.000 4.000 137.700 4.400 ;
        RECT 138.500 4.500 138.900 4.600 ;
        RECT 139.300 4.500 139.600 5.100 ;
        RECT 138.500 4.200 139.600 4.500 ;
        RECT 139.900 4.500 142.600 4.800 ;
        RECT 139.900 4.400 140.300 4.500 ;
        RECT 142.200 4.400 142.600 4.500 ;
        RECT 139.100 3.700 139.500 3.800 ;
        RECT 140.500 3.700 140.900 3.800 ;
        RECT 137.400 3.100 137.800 3.500 ;
        RECT 139.100 3.400 140.900 3.700 ;
        RECT 139.500 3.100 139.800 3.400 ;
        RECT 142.200 3.100 142.600 3.500 ;
        RECT 137.100 1.100 137.700 3.100 ;
        RECT 139.400 1.100 139.800 3.100 ;
        RECT 141.600 2.800 142.600 3.100 ;
        RECT 141.600 1.100 142.000 2.800 ;
        RECT 143.800 1.100 144.200 5.300 ;
        RECT 145.400 5.400 146.300 5.800 ;
        RECT 147.000 5.400 148.100 5.800 ;
        RECT 148.600 5.400 149.700 5.800 ;
        RECT 150.200 5.400 151.400 5.800 ;
        RECT 152.500 7.200 152.800 7.900 ;
        RECT 154.200 7.600 154.600 9.900 ;
        RECT 153.300 7.300 154.600 7.600 ;
        RECT 156.600 7.500 157.000 9.900 ;
        RECT 158.800 9.200 159.200 9.900 ;
        RECT 158.200 8.900 159.200 9.200 ;
        RECT 161.000 8.900 161.400 9.900 ;
        RECT 163.100 9.200 163.700 9.900 ;
        RECT 163.000 8.900 163.700 9.200 ;
        RECT 158.200 8.500 158.600 8.900 ;
        RECT 161.000 8.600 161.300 8.900 ;
        RECT 159.000 8.200 159.400 8.600 ;
        RECT 159.900 8.300 161.300 8.600 ;
        RECT 163.000 8.500 163.400 8.900 ;
        RECT 159.900 8.200 160.300 8.300 ;
        RECT 152.500 6.800 153.000 7.200 ;
        RECT 145.400 1.100 145.800 5.400 ;
        RECT 147.000 1.100 147.400 5.400 ;
        RECT 148.600 1.100 149.000 5.400 ;
        RECT 150.200 1.100 150.600 5.400 ;
        RECT 152.500 5.100 152.800 6.800 ;
        RECT 153.300 6.500 153.600 7.300 ;
        RECT 157.000 7.100 157.800 7.200 ;
        RECT 159.100 7.100 159.400 8.200 ;
        RECT 165.400 8.100 165.800 9.900 ;
        RECT 166.200 8.100 166.600 8.600 ;
        RECT 165.400 7.800 166.600 8.100 ;
        RECT 163.900 7.700 164.300 7.800 ;
        RECT 165.400 7.700 165.800 7.800 ;
        RECT 163.900 7.400 165.800 7.700 ;
        RECT 161.900 7.100 162.300 7.200 ;
        RECT 157.000 6.800 162.500 7.100 ;
        RECT 158.500 6.700 158.900 6.800 ;
        RECT 153.100 6.100 153.600 6.500 ;
        RECT 153.300 5.100 153.600 6.100 ;
        RECT 154.100 6.200 154.500 6.600 ;
        RECT 157.700 6.200 158.100 6.300 ;
        RECT 154.100 5.800 154.600 6.200 ;
        RECT 157.700 6.100 160.200 6.200 ;
        RECT 161.400 6.100 161.800 6.200 ;
        RECT 157.700 5.900 161.800 6.100 ;
        RECT 159.800 5.800 161.800 5.900 ;
        RECT 156.600 5.500 159.400 5.600 ;
        RECT 156.600 5.400 159.500 5.500 ;
        RECT 156.600 5.300 161.500 5.400 ;
        RECT 152.500 4.600 153.000 5.100 ;
        RECT 153.300 4.800 154.600 5.100 ;
        RECT 152.600 1.100 153.000 4.600 ;
        RECT 154.200 1.100 154.600 4.800 ;
        RECT 156.600 1.100 157.000 5.300 ;
        RECT 159.100 5.100 161.500 5.300 ;
        RECT 158.200 4.500 160.900 4.800 ;
        RECT 158.200 4.400 158.600 4.500 ;
        RECT 160.500 4.400 160.900 4.500 ;
        RECT 161.200 4.500 161.500 5.100 ;
        RECT 162.200 5.200 162.500 6.800 ;
        RECT 163.000 6.400 163.400 6.500 ;
        RECT 163.000 6.100 164.900 6.400 ;
        RECT 164.500 6.000 164.900 6.100 ;
        RECT 163.700 5.700 164.100 5.800 ;
        RECT 165.400 5.700 165.800 7.400 ;
        RECT 163.700 5.400 165.800 5.700 ;
        RECT 162.200 4.900 163.400 5.200 ;
        RECT 161.900 4.500 162.300 4.600 ;
        RECT 161.200 4.200 162.300 4.500 ;
        RECT 163.100 4.400 163.400 4.900 ;
        RECT 163.100 4.000 163.800 4.400 ;
        RECT 159.900 3.700 160.300 3.800 ;
        RECT 161.300 3.700 161.700 3.800 ;
        RECT 158.200 3.100 158.600 3.500 ;
        RECT 159.900 3.400 161.700 3.700 ;
        RECT 161.000 3.100 161.300 3.400 ;
        RECT 163.000 3.100 163.400 3.500 ;
        RECT 158.200 2.800 159.200 3.100 ;
        RECT 158.800 1.100 159.200 2.800 ;
        RECT 161.000 1.100 161.400 3.100 ;
        RECT 163.100 1.100 163.700 3.100 ;
        RECT 165.400 1.100 165.800 5.400 ;
        RECT 167.000 6.100 167.400 9.900 ;
        RECT 169.700 8.000 170.100 9.500 ;
        RECT 171.800 8.500 172.200 9.500 ;
        RECT 169.300 7.700 170.100 8.000 ;
        RECT 169.300 7.500 169.700 7.700 ;
        RECT 169.300 7.200 169.600 7.500 ;
        RECT 171.900 7.400 172.200 8.500 ;
        RECT 168.600 6.800 169.600 7.200 ;
        RECT 170.100 7.100 172.200 7.400 ;
        RECT 173.400 7.600 173.800 9.900 ;
        RECT 175.000 7.600 175.400 9.900 ;
        RECT 173.400 7.200 175.400 7.600 ;
        RECT 176.600 8.500 177.000 9.500 ;
        RECT 176.600 7.400 176.900 8.500 ;
        RECT 178.700 8.000 179.100 9.500 ;
        RECT 178.700 7.700 179.500 8.000 ;
        RECT 179.100 7.500 179.500 7.700 ;
        RECT 170.100 6.900 170.600 7.100 ;
        RECT 168.600 6.100 169.000 6.200 ;
        RECT 167.000 5.800 169.000 6.100 ;
        RECT 167.000 1.100 167.400 5.800 ;
        RECT 168.600 5.400 169.000 5.800 ;
        RECT 169.300 4.900 169.600 6.800 ;
        RECT 169.900 6.500 170.600 6.900 ;
        RECT 170.300 5.500 170.600 6.500 ;
        RECT 171.000 5.800 171.400 6.600 ;
        RECT 171.800 5.800 172.200 6.600 ;
        RECT 172.600 6.100 173.000 6.200 ;
        RECT 173.400 6.100 173.800 7.200 ;
        RECT 176.600 7.100 178.700 7.400 ;
        RECT 178.200 6.900 178.700 7.100 ;
        RECT 179.200 7.200 179.500 7.500 ;
        RECT 179.200 7.100 180.200 7.200 ;
        RECT 180.600 7.100 181.000 7.200 ;
        RECT 172.600 5.800 173.800 6.100 ;
        RECT 176.600 5.800 177.000 6.600 ;
        RECT 177.400 5.800 177.800 6.600 ;
        RECT 178.200 6.500 178.900 6.900 ;
        RECT 179.200 6.800 181.000 7.100 ;
        RECT 170.300 5.200 172.200 5.500 ;
        RECT 169.300 4.600 170.100 4.900 ;
        RECT 169.700 1.100 170.100 4.600 ;
        RECT 171.900 3.500 172.200 5.200 ;
        RECT 171.800 1.500 172.200 3.500 ;
        RECT 173.400 5.400 175.400 5.800 ;
        RECT 178.200 5.500 178.500 6.500 ;
        RECT 173.400 1.100 173.800 5.400 ;
        RECT 175.000 1.100 175.400 5.400 ;
        RECT 176.600 5.200 178.500 5.500 ;
        RECT 176.600 3.500 176.900 5.200 ;
        RECT 179.200 4.900 179.500 6.800 ;
        RECT 179.800 6.100 180.200 6.200 ;
        RECT 181.400 6.100 181.800 9.900 ;
        RECT 182.200 8.100 182.600 8.600 ;
        RECT 183.000 8.100 183.400 9.900 ;
        RECT 185.100 9.200 185.700 9.900 ;
        RECT 185.100 8.900 185.800 9.200 ;
        RECT 187.400 8.900 187.800 9.900 ;
        RECT 189.600 9.200 190.000 9.900 ;
        RECT 189.600 8.900 190.600 9.200 ;
        RECT 185.400 8.500 185.800 8.900 ;
        RECT 187.500 8.600 187.800 8.900 ;
        RECT 187.500 8.300 188.900 8.600 ;
        RECT 188.500 8.200 188.900 8.300 ;
        RECT 189.400 8.200 189.800 8.600 ;
        RECT 190.200 8.500 190.600 8.900 ;
        RECT 182.200 7.800 183.400 8.100 ;
        RECT 179.800 5.800 181.800 6.100 ;
        RECT 179.800 5.400 180.200 5.800 ;
        RECT 178.700 4.600 179.500 4.900 ;
        RECT 176.600 1.500 177.000 3.500 ;
        RECT 178.700 1.100 179.100 4.600 ;
        RECT 181.400 1.100 181.800 5.800 ;
        RECT 183.000 7.700 183.400 7.800 ;
        RECT 184.500 7.700 184.900 7.800 ;
        RECT 183.000 7.400 184.900 7.700 ;
        RECT 183.000 5.700 183.400 7.400 ;
        RECT 186.500 7.100 186.900 7.200 ;
        RECT 189.400 7.100 189.700 8.200 ;
        RECT 191.800 7.500 192.200 9.900 ;
        RECT 192.600 7.500 193.000 9.900 ;
        RECT 194.800 9.200 195.200 9.900 ;
        RECT 194.200 8.900 195.200 9.200 ;
        RECT 197.000 8.900 197.400 9.900 ;
        RECT 199.100 9.200 199.700 9.900 ;
        RECT 199.000 8.900 199.700 9.200 ;
        RECT 194.200 8.500 194.600 8.900 ;
        RECT 197.000 8.600 197.300 8.900 ;
        RECT 195.000 8.200 195.400 8.600 ;
        RECT 195.900 8.300 197.300 8.600 ;
        RECT 199.000 8.500 199.400 8.900 ;
        RECT 195.900 8.200 196.300 8.300 ;
        RECT 191.000 7.100 191.800 7.200 ;
        RECT 186.300 6.800 191.800 7.100 ;
        RECT 193.000 7.100 193.800 7.200 ;
        RECT 195.100 7.100 195.400 8.200 ;
        RECT 199.900 7.700 200.300 7.800 ;
        RECT 201.400 7.700 201.800 9.900 ;
        RECT 199.900 7.400 201.800 7.700 ;
        RECT 202.200 7.500 202.600 9.900 ;
        RECT 204.400 9.200 204.800 9.900 ;
        RECT 203.800 8.900 204.800 9.200 ;
        RECT 206.600 8.900 207.000 9.900 ;
        RECT 208.700 9.200 209.300 9.900 ;
        RECT 208.600 8.900 209.300 9.200 ;
        RECT 203.800 8.500 204.200 8.900 ;
        RECT 206.600 8.600 206.900 8.900 ;
        RECT 204.600 8.200 205.000 8.600 ;
        RECT 205.500 8.300 206.900 8.600 ;
        RECT 208.600 8.500 209.000 8.900 ;
        RECT 205.500 8.200 205.900 8.300 ;
        RECT 197.900 7.100 198.600 7.200 ;
        RECT 193.000 6.800 198.600 7.100 ;
        RECT 185.400 6.400 185.800 6.500 ;
        RECT 183.900 6.100 185.800 6.400 ;
        RECT 183.900 6.000 184.300 6.100 ;
        RECT 184.700 5.700 185.100 5.800 ;
        RECT 183.000 5.400 185.100 5.700 ;
        RECT 183.000 1.100 183.400 5.400 ;
        RECT 186.300 5.200 186.600 6.800 ;
        RECT 189.900 6.700 190.300 6.800 ;
        RECT 194.500 6.700 194.900 6.800 ;
        RECT 190.700 6.200 191.100 6.300 ;
        RECT 188.600 5.900 191.100 6.200 ;
        RECT 193.700 6.200 194.100 6.300 ;
        RECT 193.700 5.900 196.200 6.200 ;
        RECT 188.600 5.800 189.000 5.900 ;
        RECT 195.800 5.800 196.200 5.900 ;
        RECT 189.400 5.500 192.200 5.600 ;
        RECT 189.300 5.400 192.200 5.500 ;
        RECT 185.400 4.900 186.600 5.200 ;
        RECT 187.300 5.300 192.200 5.400 ;
        RECT 187.300 5.100 189.700 5.300 ;
        RECT 185.400 4.400 185.700 4.900 ;
        RECT 185.000 4.000 185.700 4.400 ;
        RECT 186.500 4.500 186.900 4.600 ;
        RECT 187.300 4.500 187.600 5.100 ;
        RECT 186.500 4.200 187.600 4.500 ;
        RECT 187.900 4.500 190.600 4.800 ;
        RECT 187.900 4.400 188.300 4.500 ;
        RECT 190.200 4.400 190.600 4.500 ;
        RECT 187.100 3.700 187.500 3.800 ;
        RECT 188.500 3.700 188.900 3.800 ;
        RECT 185.400 3.100 185.800 3.500 ;
        RECT 187.100 3.400 188.900 3.700 ;
        RECT 187.500 3.100 187.800 3.400 ;
        RECT 190.200 3.100 190.600 3.500 ;
        RECT 185.100 1.100 185.700 3.100 ;
        RECT 187.400 1.100 187.800 3.100 ;
        RECT 189.600 2.800 190.600 3.100 ;
        RECT 189.600 1.100 190.000 2.800 ;
        RECT 191.800 1.100 192.200 5.300 ;
        RECT 192.600 5.500 195.400 5.600 ;
        RECT 192.600 5.400 195.500 5.500 ;
        RECT 192.600 5.300 197.500 5.400 ;
        RECT 192.600 1.100 193.000 5.300 ;
        RECT 195.100 5.100 197.500 5.300 ;
        RECT 194.200 4.500 196.900 4.800 ;
        RECT 194.200 4.400 194.600 4.500 ;
        RECT 196.500 4.400 196.900 4.500 ;
        RECT 197.200 4.500 197.500 5.100 ;
        RECT 198.200 5.200 198.500 6.800 ;
        RECT 199.000 6.400 199.400 6.500 ;
        RECT 199.000 6.100 200.900 6.400 ;
        RECT 200.500 6.000 200.900 6.100 ;
        RECT 199.700 5.700 200.100 5.800 ;
        RECT 201.400 5.700 201.800 7.400 ;
        RECT 202.600 7.100 203.400 7.200 ;
        RECT 204.700 7.100 205.000 8.200 ;
        RECT 209.500 7.700 209.900 7.800 ;
        RECT 211.000 7.700 211.400 9.900 ;
        RECT 213.400 8.000 213.800 9.900 ;
        RECT 215.000 8.000 215.400 9.900 ;
        RECT 213.400 7.900 215.400 8.000 ;
        RECT 215.800 7.900 216.200 9.900 ;
        RECT 216.900 8.200 217.300 9.900 ;
        RECT 216.900 7.900 217.800 8.200 ;
        RECT 213.500 7.700 215.300 7.900 ;
        RECT 209.500 7.400 211.400 7.700 ;
        RECT 206.200 7.100 206.600 7.200 ;
        RECT 207.500 7.100 207.900 7.200 ;
        RECT 202.600 6.800 208.100 7.100 ;
        RECT 204.100 6.700 204.500 6.800 ;
        RECT 203.300 6.200 203.700 6.300 ;
        RECT 203.300 5.900 205.800 6.200 ;
        RECT 205.400 5.800 205.800 5.900 ;
        RECT 199.700 5.400 201.800 5.700 ;
        RECT 198.200 4.900 199.400 5.200 ;
        RECT 197.900 4.500 198.300 4.600 ;
        RECT 197.200 4.200 198.300 4.500 ;
        RECT 199.100 4.400 199.400 4.900 ;
        RECT 199.100 4.000 199.800 4.400 ;
        RECT 195.900 3.700 196.300 3.800 ;
        RECT 197.300 3.700 197.700 3.800 ;
        RECT 194.200 3.100 194.600 3.500 ;
        RECT 195.900 3.400 197.700 3.700 ;
        RECT 197.000 3.100 197.300 3.400 ;
        RECT 199.000 3.100 199.400 3.500 ;
        RECT 194.200 2.800 195.200 3.100 ;
        RECT 194.800 1.100 195.200 2.800 ;
        RECT 197.000 1.100 197.400 3.100 ;
        RECT 199.100 1.100 199.700 3.100 ;
        RECT 201.400 1.100 201.800 5.400 ;
        RECT 202.200 5.500 205.000 5.600 ;
        RECT 202.200 5.400 205.100 5.500 ;
        RECT 202.200 5.300 207.100 5.400 ;
        RECT 202.200 1.100 202.600 5.300 ;
        RECT 204.700 5.100 207.100 5.300 ;
        RECT 203.800 4.500 206.500 4.800 ;
        RECT 203.800 4.400 204.200 4.500 ;
        RECT 206.100 4.400 206.500 4.500 ;
        RECT 206.800 4.500 207.100 5.100 ;
        RECT 207.800 5.200 208.100 6.800 ;
        RECT 208.600 6.400 209.000 6.500 ;
        RECT 208.600 6.100 210.500 6.400 ;
        RECT 210.100 6.000 210.500 6.100 ;
        RECT 209.300 5.700 209.700 5.800 ;
        RECT 211.000 5.700 211.400 7.400 ;
        RECT 213.800 7.200 214.200 7.400 ;
        RECT 215.800 7.200 216.100 7.900 ;
        RECT 213.400 6.900 214.200 7.200 ;
        RECT 213.400 6.800 213.800 6.900 ;
        RECT 214.900 6.800 216.200 7.200 ;
        RECT 214.200 5.800 214.600 6.600 ;
        RECT 214.900 6.200 215.200 6.800 ;
        RECT 214.900 5.800 215.400 6.200 ;
        RECT 217.400 6.100 217.800 7.900 ;
        RECT 219.800 7.600 220.200 9.900 ;
        RECT 221.400 7.600 221.800 9.900 ;
        RECT 223.000 7.600 223.400 9.900 ;
        RECT 224.600 7.600 225.000 9.900 ;
        RECT 226.200 7.900 226.600 9.900 ;
        RECT 227.000 8.000 227.400 9.900 ;
        RECT 228.600 8.000 229.000 9.900 ;
        RECT 227.000 7.900 229.000 8.000 ;
        RECT 218.200 6.800 218.600 7.600 ;
        RECT 219.000 7.200 220.200 7.600 ;
        RECT 220.700 7.200 221.800 7.600 ;
        RECT 222.300 7.200 223.400 7.600 ;
        RECT 224.100 7.200 225.000 7.600 ;
        RECT 226.300 7.200 226.600 7.900 ;
        RECT 227.100 7.700 228.900 7.900 ;
        RECT 229.400 7.700 229.800 9.900 ;
        RECT 231.500 9.200 232.100 9.900 ;
        RECT 231.500 8.900 232.200 9.200 ;
        RECT 233.800 8.900 234.200 9.900 ;
        RECT 236.000 9.200 236.400 9.900 ;
        RECT 236.000 8.900 237.000 9.200 ;
        RECT 231.800 8.500 232.200 8.900 ;
        RECT 233.900 8.600 234.200 8.900 ;
        RECT 233.900 8.300 235.300 8.600 ;
        RECT 234.900 8.200 235.300 8.300 ;
        RECT 235.800 8.200 236.200 8.600 ;
        RECT 236.600 8.500 237.000 8.900 ;
        RECT 230.900 7.700 231.300 7.800 ;
        RECT 229.400 7.400 231.300 7.700 ;
        RECT 228.200 7.200 228.600 7.400 ;
        RECT 215.800 5.800 217.800 6.100 ;
        RECT 209.300 5.400 211.400 5.700 ;
        RECT 207.800 4.900 209.000 5.200 ;
        RECT 207.500 4.500 207.900 4.600 ;
        RECT 206.800 4.200 207.900 4.500 ;
        RECT 208.700 4.400 209.000 4.900 ;
        RECT 208.700 4.000 209.400 4.400 ;
        RECT 205.500 3.700 205.900 3.800 ;
        RECT 206.900 3.700 207.300 3.800 ;
        RECT 203.800 3.100 204.200 3.500 ;
        RECT 205.500 3.400 207.300 3.700 ;
        RECT 206.600 3.100 206.900 3.400 ;
        RECT 208.600 3.100 209.000 3.500 ;
        RECT 203.800 2.800 204.800 3.100 ;
        RECT 204.400 1.100 204.800 2.800 ;
        RECT 206.600 1.100 207.000 3.100 ;
        RECT 208.700 1.100 209.300 3.100 ;
        RECT 211.000 1.100 211.400 5.400 ;
        RECT 214.900 5.100 215.200 5.800 ;
        RECT 215.800 5.200 216.100 5.800 ;
        RECT 215.800 5.100 216.200 5.200 ;
        RECT 214.700 4.800 215.200 5.100 ;
        RECT 215.500 4.800 216.200 5.100 ;
        RECT 214.700 1.100 215.100 4.800 ;
        RECT 215.500 4.200 215.800 4.800 ;
        RECT 216.600 4.400 217.000 5.200 ;
        RECT 215.400 3.800 215.800 4.200 ;
        RECT 217.400 1.100 217.800 5.800 ;
        RECT 219.000 5.800 219.400 7.200 ;
        RECT 220.700 6.900 221.100 7.200 ;
        RECT 222.300 6.900 222.700 7.200 ;
        RECT 224.100 6.900 224.500 7.200 ;
        RECT 225.400 6.900 225.800 7.200 ;
        RECT 219.800 6.500 221.100 6.900 ;
        RECT 221.500 6.500 222.700 6.900 ;
        RECT 223.200 6.500 224.500 6.900 ;
        RECT 224.900 6.500 225.800 6.900 ;
        RECT 226.200 6.800 227.500 7.200 ;
        RECT 228.200 6.900 229.000 7.200 ;
        RECT 228.600 6.800 229.000 6.900 ;
        RECT 220.700 5.800 221.100 6.500 ;
        RECT 222.300 5.800 222.700 6.500 ;
        RECT 224.100 5.800 224.500 6.500 ;
        RECT 227.200 6.200 227.500 6.800 ;
        RECT 227.000 5.800 227.500 6.200 ;
        RECT 227.800 5.800 228.200 6.600 ;
        RECT 219.000 5.400 220.200 5.800 ;
        RECT 220.700 5.400 221.800 5.800 ;
        RECT 222.300 5.400 223.400 5.800 ;
        RECT 224.100 5.400 225.000 5.800 ;
        RECT 219.800 1.100 220.200 5.400 ;
        RECT 221.400 1.100 221.800 5.400 ;
        RECT 223.000 1.100 223.400 5.400 ;
        RECT 224.600 1.100 225.000 5.400 ;
        RECT 226.200 5.100 226.600 5.200 ;
        RECT 227.200 5.100 227.500 5.800 ;
        RECT 229.400 5.700 229.800 7.400 ;
        RECT 232.900 7.100 233.300 7.200 ;
        RECT 235.800 7.100 236.100 8.200 ;
        RECT 238.200 7.500 238.600 9.900 ;
        RECT 239.800 7.600 240.200 9.900 ;
        RECT 241.400 7.600 241.800 9.900 ;
        RECT 243.000 7.600 243.400 9.900 ;
        RECT 244.600 7.600 245.000 9.900 ;
        RECT 247.000 7.600 247.400 9.900 ;
        RECT 248.600 7.600 249.000 9.900 ;
        RECT 250.200 7.600 250.600 9.900 ;
        RECT 251.800 7.600 252.200 9.900 ;
        RECT 253.400 7.700 253.800 9.900 ;
        RECT 255.500 9.200 256.100 9.900 ;
        RECT 255.500 8.900 256.200 9.200 ;
        RECT 257.800 8.900 258.200 9.900 ;
        RECT 260.000 9.200 260.400 9.900 ;
        RECT 260.000 8.900 261.000 9.200 ;
        RECT 255.800 8.500 256.200 8.900 ;
        RECT 257.900 8.600 258.200 8.900 ;
        RECT 257.900 8.300 259.300 8.600 ;
        RECT 258.900 8.200 259.300 8.300 ;
        RECT 259.800 8.200 260.200 8.600 ;
        RECT 260.600 8.500 261.000 8.900 ;
        RECT 254.900 7.700 255.300 7.800 ;
        RECT 239.800 7.200 240.700 7.600 ;
        RECT 241.400 7.200 242.500 7.600 ;
        RECT 243.000 7.200 244.100 7.600 ;
        RECT 244.600 7.200 245.800 7.600 ;
        RECT 247.000 7.200 247.900 7.600 ;
        RECT 248.600 7.200 249.700 7.600 ;
        RECT 250.200 7.200 251.300 7.600 ;
        RECT 251.800 7.200 253.000 7.600 ;
        RECT 237.400 7.100 238.200 7.200 ;
        RECT 232.700 6.800 238.200 7.100 ;
        RECT 240.300 6.900 240.700 7.200 ;
        RECT 242.100 6.900 242.500 7.200 ;
        RECT 243.700 6.900 244.100 7.200 ;
        RECT 231.800 6.400 232.200 6.500 ;
        RECT 230.300 6.100 232.200 6.400 ;
        RECT 230.300 6.000 230.700 6.100 ;
        RECT 231.100 5.700 231.500 5.800 ;
        RECT 229.400 5.400 231.500 5.700 ;
        RECT 226.200 4.800 226.900 5.100 ;
        RECT 227.200 4.800 227.700 5.100 ;
        RECT 226.600 4.200 226.900 4.800 ;
        RECT 226.600 3.800 227.000 4.200 ;
        RECT 227.300 1.100 227.700 4.800 ;
        RECT 229.400 1.100 229.800 5.400 ;
        RECT 232.700 5.200 233.000 6.800 ;
        RECT 236.300 6.700 236.700 6.800 ;
        RECT 240.300 6.500 241.600 6.900 ;
        RECT 242.100 6.500 243.300 6.900 ;
        RECT 243.700 6.500 245.000 6.900 ;
        RECT 237.100 6.200 237.500 6.300 ;
        RECT 235.000 5.900 237.500 6.200 ;
        RECT 235.000 5.800 235.400 5.900 ;
        RECT 240.300 5.800 240.700 6.500 ;
        RECT 242.100 5.800 242.500 6.500 ;
        RECT 243.700 5.800 244.100 6.500 ;
        RECT 245.400 5.800 245.800 7.200 ;
        RECT 246.200 6.900 246.600 7.200 ;
        RECT 247.500 6.900 247.900 7.200 ;
        RECT 249.300 6.900 249.700 7.200 ;
        RECT 250.900 6.900 251.300 7.200 ;
        RECT 246.200 6.500 247.100 6.900 ;
        RECT 247.500 6.500 248.800 6.900 ;
        RECT 249.300 6.500 250.500 6.900 ;
        RECT 250.900 6.500 252.200 6.900 ;
        RECT 247.500 5.800 247.900 6.500 ;
        RECT 249.300 5.800 249.700 6.500 ;
        RECT 250.900 5.800 251.300 6.500 ;
        RECT 252.600 5.800 253.000 7.200 ;
        RECT 235.800 5.500 238.600 5.600 ;
        RECT 235.700 5.400 238.600 5.500 ;
        RECT 231.800 4.900 233.000 5.200 ;
        RECT 233.700 5.300 238.600 5.400 ;
        RECT 233.700 5.100 236.100 5.300 ;
        RECT 231.800 4.400 232.100 4.900 ;
        RECT 231.400 4.000 232.100 4.400 ;
        RECT 232.900 4.500 233.300 4.600 ;
        RECT 233.700 4.500 234.000 5.100 ;
        RECT 232.900 4.200 234.000 4.500 ;
        RECT 234.300 4.500 237.000 4.800 ;
        RECT 234.300 4.400 234.700 4.500 ;
        RECT 236.600 4.400 237.000 4.500 ;
        RECT 233.500 3.700 233.900 3.800 ;
        RECT 234.900 3.700 235.300 3.800 ;
        RECT 231.800 3.100 232.200 3.500 ;
        RECT 233.500 3.400 235.300 3.700 ;
        RECT 233.900 3.100 234.200 3.400 ;
        RECT 236.600 3.100 237.000 3.500 ;
        RECT 231.500 1.100 232.100 3.100 ;
        RECT 233.800 1.100 234.200 3.100 ;
        RECT 236.000 2.800 237.000 3.100 ;
        RECT 236.000 1.100 236.400 2.800 ;
        RECT 238.200 1.100 238.600 5.300 ;
        RECT 239.800 5.400 240.700 5.800 ;
        RECT 241.400 5.400 242.500 5.800 ;
        RECT 243.000 5.400 244.100 5.800 ;
        RECT 244.600 5.400 245.800 5.800 ;
        RECT 247.000 5.400 247.900 5.800 ;
        RECT 248.600 5.400 249.700 5.800 ;
        RECT 250.200 5.400 251.300 5.800 ;
        RECT 251.800 5.400 253.000 5.800 ;
        RECT 253.400 7.400 255.300 7.700 ;
        RECT 253.400 5.700 253.800 7.400 ;
        RECT 256.900 7.100 257.300 7.200 ;
        RECT 259.800 7.100 260.100 8.200 ;
        RECT 262.200 7.500 262.600 9.900 ;
        RECT 261.400 7.100 262.200 7.200 ;
        RECT 256.700 6.800 262.200 7.100 ;
        RECT 255.800 6.400 256.200 6.500 ;
        RECT 254.300 6.100 256.200 6.400 ;
        RECT 256.700 6.200 257.000 6.800 ;
        RECT 260.300 6.700 260.700 6.800 ;
        RECT 259.800 6.200 260.200 6.300 ;
        RECT 261.100 6.200 261.500 6.300 ;
        RECT 254.300 6.000 254.700 6.100 ;
        RECT 256.600 5.800 257.000 6.200 ;
        RECT 259.000 5.900 261.500 6.200 ;
        RECT 259.000 5.800 259.400 5.900 ;
        RECT 255.100 5.700 255.500 5.800 ;
        RECT 253.400 5.400 255.500 5.700 ;
        RECT 239.800 1.100 240.200 5.400 ;
        RECT 241.400 1.100 241.800 5.400 ;
        RECT 243.000 1.100 243.400 5.400 ;
        RECT 244.600 1.100 245.000 5.400 ;
        RECT 247.000 1.100 247.400 5.400 ;
        RECT 248.600 1.100 249.000 5.400 ;
        RECT 250.200 1.100 250.600 5.400 ;
        RECT 251.800 1.100 252.200 5.400 ;
        RECT 253.400 1.100 253.800 5.400 ;
        RECT 256.700 5.200 257.000 5.800 ;
        RECT 259.800 5.500 262.600 5.600 ;
        RECT 259.700 5.400 262.600 5.500 ;
        RECT 255.800 4.900 257.000 5.200 ;
        RECT 257.700 5.300 262.600 5.400 ;
        RECT 257.700 5.100 260.100 5.300 ;
        RECT 255.800 4.400 256.100 4.900 ;
        RECT 255.400 4.000 256.100 4.400 ;
        RECT 256.900 4.500 257.300 4.600 ;
        RECT 257.700 4.500 258.000 5.100 ;
        RECT 256.900 4.200 258.000 4.500 ;
        RECT 258.300 4.500 261.000 4.800 ;
        RECT 258.300 4.400 258.700 4.500 ;
        RECT 260.600 4.400 261.000 4.500 ;
        RECT 257.500 3.700 257.900 3.800 ;
        RECT 258.900 3.700 259.300 3.800 ;
        RECT 255.800 3.100 256.200 3.500 ;
        RECT 257.500 3.400 259.300 3.700 ;
        RECT 257.900 3.100 258.200 3.400 ;
        RECT 260.600 3.100 261.000 3.500 ;
        RECT 255.500 1.100 256.100 3.100 ;
        RECT 257.800 1.100 258.200 3.100 ;
        RECT 260.000 2.800 261.000 3.100 ;
        RECT 260.000 1.100 260.400 2.800 ;
        RECT 262.200 1.100 262.600 5.300 ;
      LAYER via1 ;
        RECT 27.800 236.800 28.200 237.200 ;
        RECT 47.000 234.800 47.400 235.200 ;
        RECT 44.600 233.800 45.000 234.200 ;
        RECT 6.200 231.800 6.600 232.200 ;
        RECT 13.400 231.800 13.800 232.200 ;
        RECT 15.800 231.800 16.200 232.200 ;
        RECT 42.200 231.800 42.600 232.200 ;
        RECT 43.800 233.100 44.200 233.500 ;
        RECT 49.400 233.800 49.800 234.200 ;
        RECT 52.600 231.800 53.000 232.200 ;
        RECT 64.600 233.800 65.000 234.200 ;
        RECT 60.600 232.800 61.000 233.200 ;
        RECT 71.000 234.800 71.400 235.200 ;
        RECT 67.000 233.800 67.400 234.200 ;
        RECT 68.600 233.800 69.000 234.200 ;
        RECT 67.800 233.100 68.200 233.500 ;
        RECT 80.600 234.800 81.000 235.200 ;
        RECT 76.600 231.800 77.000 232.200 ;
        RECT 77.400 233.100 77.800 233.500 ;
        RECT 87.000 232.800 87.400 233.200 ;
        RECT 91.800 234.800 92.200 235.200 ;
        RECT 92.600 234.800 93.000 235.200 ;
        RECT 97.400 234.800 97.800 235.200 ;
        RECT 93.400 233.100 93.800 233.500 ;
        RECT 109.400 235.800 109.800 236.200 ;
        RECT 107.800 234.800 108.200 235.200 ;
        RECT 107.800 233.800 108.200 234.200 ;
        RECT 111.000 234.800 111.400 235.200 ;
        RECT 118.200 234.800 118.600 235.200 ;
        RECT 109.400 233.800 109.800 234.200 ;
        RECT 111.800 233.800 112.200 234.200 ;
        RECT 113.400 233.100 113.800 233.500 ;
        RECT 123.800 234.800 124.200 235.200 ;
        RECT 124.600 234.800 125.000 235.200 ;
        RECT 138.200 236.800 138.600 237.200 ;
        RECT 102.200 231.800 102.600 232.200 ;
        RECT 115.800 232.800 116.200 233.200 ;
        RECT 131.800 234.800 132.200 235.200 ;
        RECT 127.800 233.800 128.200 234.200 ;
        RECT 129.400 233.800 129.800 234.200 ;
        RECT 122.200 231.800 122.600 232.200 ;
        RECT 128.600 233.100 129.000 233.500 ;
        RECT 138.200 233.800 138.600 234.200 ;
        RECT 142.200 234.800 142.600 235.200 ;
        RECT 143.000 233.800 143.400 234.200 ;
        RECT 147.000 232.800 147.400 233.200 ;
        RECT 156.600 236.200 157.000 236.600 ;
        RECT 158.200 235.500 158.600 235.900 ;
        RECT 175.000 236.800 175.400 237.200 ;
        RECT 158.200 233.100 158.600 233.500 ;
        RECT 164.600 234.800 165.000 235.200 ;
        RECT 162.200 233.800 162.600 234.200 ;
        RECT 165.400 233.800 165.800 234.200 ;
        RECT 166.200 233.100 166.600 233.500 ;
        RECT 175.800 234.800 176.200 235.200 ;
        RECT 176.600 234.800 177.000 235.200 ;
        RECT 184.600 235.800 185.000 236.200 ;
        RECT 195.000 236.800 195.400 237.200 ;
        RECT 149.400 231.800 149.800 232.200 ;
        RECT 168.600 232.800 169.000 233.200 ;
        RECT 180.600 233.800 181.000 234.200 ;
        RECT 184.600 234.800 185.000 235.200 ;
        RECT 185.400 233.800 185.800 234.200 ;
        RECT 187.000 233.800 187.400 234.200 ;
        RECT 186.200 233.100 186.600 233.500 ;
        RECT 203.000 236.200 203.400 236.600 ;
        RECT 204.600 235.500 205.000 235.900 ;
        RECT 222.200 234.800 222.600 235.200 ;
        RECT 204.600 233.100 205.000 233.500 ;
        RECT 195.800 231.800 196.200 232.200 ;
        RECT 238.200 234.800 238.600 235.200 ;
        RECT 226.200 233.800 226.600 234.200 ;
        RECT 223.800 231.800 224.200 232.200 ;
        RECT 234.200 233.100 234.600 233.500 ;
        RECT 243.000 231.800 243.400 232.200 ;
        RECT 243.800 236.800 244.200 237.200 ;
        RECT 251.000 236.200 251.400 236.600 ;
        RECT 252.600 235.500 253.000 235.900 ;
        RECT 250.200 232.800 250.600 233.200 ;
        RECT 252.600 233.100 253.000 233.500 ;
        RECT 255.000 233.800 255.400 234.200 ;
        RECT 261.400 231.800 261.800 232.200 ;
        RECT 0.600 226.800 1.000 227.200 ;
        RECT 7.000 226.800 7.400 227.200 ;
        RECT 8.600 226.800 9.000 227.200 ;
        RECT 12.600 225.800 13.000 226.200 ;
        RECT 7.800 225.100 8.200 225.500 ;
        RECT 31.800 228.800 32.200 229.200 ;
        RECT 18.200 226.800 18.600 227.200 ;
        RECT 20.600 225.800 21.000 226.200 ;
        RECT 23.000 225.100 23.400 225.500 ;
        RECT 16.600 223.800 17.000 224.200 ;
        RECT 30.200 223.800 30.600 224.200 ;
        RECT 42.200 225.800 42.600 226.200 ;
        RECT 46.200 225.800 46.600 226.200 ;
        RECT 63.000 228.800 63.400 229.200 ;
        RECT 56.600 226.800 57.000 227.200 ;
        RECT 47.000 221.800 47.400 222.200 ;
        RECT 54.200 225.100 54.600 225.500 ;
        RECT 65.400 226.800 65.800 227.200 ;
        RECT 67.000 224.800 67.400 225.200 ;
        RECT 79.800 226.800 80.200 227.200 ;
        RECT 95.000 228.800 95.400 229.200 ;
        RECT 76.600 226.100 77.000 226.500 ;
        RECT 71.800 221.800 72.200 222.200 ;
        RECT 80.600 225.900 81.000 226.300 ;
        RECT 83.000 225.100 83.400 225.500 ;
        RECT 85.400 225.800 85.800 226.200 ;
        RECT 87.800 226.800 88.200 227.200 ;
        RECT 89.400 226.800 89.800 227.200 ;
        RECT 88.600 225.800 89.000 226.200 ;
        RECT 97.400 226.800 97.800 227.200 ;
        RECT 100.600 225.800 101.000 226.200 ;
        RECT 74.200 221.800 74.600 222.200 ;
        RECT 95.000 221.800 95.400 222.200 ;
        RECT 96.600 225.100 97.000 225.500 ;
        RECT 110.200 228.800 110.600 229.200 ;
        RECT 107.000 223.800 107.400 224.200 ;
        RECT 116.600 228.800 117.000 229.200 ;
        RECT 114.200 224.800 114.600 225.200 ;
        RECT 119.000 221.800 119.400 222.200 ;
        RECT 142.200 228.800 142.600 229.200 ;
        RECT 130.200 225.800 130.600 226.200 ;
        RECT 136.600 225.800 137.000 226.200 ;
        RECT 129.400 221.800 129.800 222.200 ;
        RECT 134.200 221.800 134.600 222.200 ;
        RECT 148.600 226.800 149.000 227.200 ;
        RECT 144.600 226.100 145.000 226.500 ;
        RECT 138.200 224.800 138.600 225.200 ;
        RECT 140.600 224.800 141.000 225.200 ;
        RECT 163.000 228.800 163.400 229.200 ;
        RECT 151.000 225.100 151.400 225.500 ;
        RECT 155.000 225.800 155.400 226.200 ;
        RECT 159.000 225.800 159.400 226.200 ;
        RECT 168.600 226.800 169.000 227.200 ;
        RECT 165.400 226.100 165.800 226.500 ;
        RECT 169.400 225.900 169.800 226.300 ;
        RECT 171.800 225.100 172.200 225.500 ;
        RECT 174.200 225.800 174.600 226.200 ;
        RECT 176.600 226.800 177.000 227.200 ;
        RECT 178.200 225.800 178.600 226.200 ;
        RECT 179.000 225.800 179.400 226.200 ;
        RECT 183.000 224.800 183.400 225.200 ;
        RECT 183.800 221.800 184.200 222.200 ;
        RECT 191.000 226.800 191.400 227.200 ;
        RECT 198.200 228.800 198.600 229.200 ;
        RECT 193.400 226.800 193.800 227.200 ;
        RECT 187.800 226.100 188.200 226.500 ;
        RECT 194.200 225.100 194.600 225.500 ;
        RECT 196.600 225.800 197.000 226.200 ;
        RECT 200.600 228.800 201.000 229.200 ;
        RECT 199.000 226.800 199.400 227.200 ;
        RECT 199.800 225.800 200.200 226.200 ;
        RECT 208.600 226.800 209.000 227.200 ;
        RECT 203.000 226.100 203.400 226.500 ;
        RECT 207.000 225.900 207.400 226.300 ;
        RECT 209.400 225.100 209.800 225.500 ;
        RECT 213.400 225.800 213.800 226.200 ;
        RECT 226.200 228.800 226.600 229.200 ;
        RECT 215.800 226.800 216.200 227.200 ;
        RECT 220.600 226.800 221.000 227.200 ;
        RECT 216.600 225.800 217.000 226.200 ;
        RECT 221.400 225.800 221.800 226.200 ;
        RECT 217.400 225.100 217.800 225.500 ;
        RECT 226.200 221.800 226.600 222.200 ;
        RECT 238.200 228.800 238.600 229.200 ;
        RECT 231.800 225.800 232.200 226.200 ;
        RECT 227.800 221.800 228.200 222.200 ;
        RECT 243.800 228.800 244.200 229.200 ;
        RECT 239.000 224.800 239.400 225.200 ;
        RECT 243.000 224.800 243.400 225.200 ;
        RECT 253.400 226.800 253.800 227.200 ;
        RECT 247.800 221.800 248.200 222.200 ;
        RECT 254.200 224.800 254.600 225.200 ;
        RECT 262.200 228.800 262.600 229.200 ;
        RECT 256.600 226.800 257.000 227.200 ;
        RECT 255.000 221.800 255.400 222.200 ;
        RECT 7.800 216.200 8.200 216.600 ;
        RECT 9.400 215.500 9.800 215.900 ;
        RECT 9.400 213.100 9.800 213.500 ;
        RECT 0.600 211.800 1.000 212.200 ;
        RECT 10.200 212.800 10.600 213.200 ;
        RECT 23.000 216.200 23.400 216.600 ;
        RECT 24.600 215.500 25.000 215.900 ;
        RECT 32.600 216.200 33.000 216.600 ;
        RECT 34.200 215.500 34.600 215.900 ;
        RECT 46.200 218.800 46.600 219.200 ;
        RECT 24.600 213.100 25.000 213.500 ;
        RECT 15.800 211.800 16.200 212.200 ;
        RECT 35.000 213.800 35.400 214.200 ;
        RECT 34.200 213.100 34.600 213.500 ;
        RECT 25.400 211.800 25.800 212.200 ;
        RECT 39.000 214.800 39.400 215.200 ;
        RECT 41.400 213.800 41.800 214.200 ;
        RECT 43.000 214.800 43.400 215.200 ;
        RECT 43.800 214.800 44.200 215.200 ;
        RECT 44.600 214.800 45.000 215.200 ;
        RECT 55.800 216.800 56.200 217.200 ;
        RECT 53.400 214.800 53.800 215.200 ;
        RECT 49.400 213.800 49.800 214.200 ;
        RECT 48.600 213.100 49.000 213.500 ;
        RECT 63.800 214.800 64.200 215.200 ;
        RECT 66.200 214.800 66.600 215.200 ;
        RECT 64.600 213.800 65.000 214.200 ;
        RECT 68.600 213.800 69.000 214.200 ;
        RECT 70.200 213.800 70.600 214.200 ;
        RECT 78.200 216.200 78.600 216.600 ;
        RECT 79.800 215.500 80.200 215.900 ;
        RECT 75.000 214.800 75.400 215.200 ;
        RECT 59.000 211.800 59.400 212.200 ;
        RECT 87.800 216.200 88.200 216.600 ;
        RECT 89.400 215.500 89.800 215.900 ;
        RECT 93.400 214.800 93.800 215.200 ;
        RECT 79.800 213.100 80.200 213.500 ;
        RECT 89.400 213.100 89.800 213.500 ;
        RECT 80.600 211.800 81.000 212.200 ;
        RECT 90.200 213.100 90.600 213.500 ;
        RECT 99.000 211.800 99.400 212.200 ;
        RECT 111.800 216.200 112.200 216.600 ;
        RECT 113.400 215.500 113.800 215.900 ;
        RECT 113.400 213.100 113.800 213.500 ;
        RECT 104.600 211.800 105.000 212.200 ;
        RECT 115.800 212.800 116.200 213.200 ;
        RECT 115.000 211.800 115.400 212.200 ;
        RECT 128.600 216.200 129.000 216.600 ;
        RECT 130.200 215.500 130.600 215.900 ;
        RECT 140.600 218.800 141.000 219.200 ;
        RECT 134.200 214.800 134.600 215.200 ;
        RECT 135.000 214.800 135.400 215.200 ;
        RECT 130.200 213.100 130.600 213.500 ;
        RECT 121.400 211.800 121.800 212.200 ;
        RECT 138.200 214.800 138.600 215.200 ;
        RECT 136.600 211.800 137.000 212.200 ;
        RECT 156.600 216.200 157.000 216.600 ;
        RECT 158.200 215.500 158.600 215.900 ;
        RECT 167.800 216.800 168.200 217.200 ;
        RECT 160.600 214.800 161.000 215.200 ;
        RECT 158.200 213.100 158.600 213.500 ;
        RECT 149.400 211.800 149.800 212.200 ;
        RECT 175.000 216.200 175.400 216.600 ;
        RECT 176.600 215.500 177.000 215.900 ;
        RECT 184.600 218.800 185.000 219.200 ;
        RECT 187.000 218.800 187.400 219.200 ;
        RECT 171.800 213.800 172.200 214.200 ;
        RECT 177.400 213.800 177.800 214.200 ;
        RECT 176.600 213.100 177.000 213.500 ;
        RECT 181.400 214.800 181.800 215.200 ;
        RECT 184.600 214.800 185.000 215.200 ;
        RECT 182.200 213.800 182.600 214.200 ;
        RECT 185.400 213.800 185.800 214.200 ;
        RECT 194.200 214.800 194.600 215.200 ;
        RECT 195.800 213.800 196.200 214.200 ;
        RECT 198.200 213.800 198.600 214.200 ;
        RECT 206.200 216.200 206.600 216.600 ;
        RECT 207.800 215.500 208.200 215.900 ;
        RECT 219.000 216.800 219.400 217.200 ;
        RECT 223.800 218.800 224.200 219.200 ;
        RECT 207.800 213.100 208.200 213.500 ;
        RECT 199.000 211.800 199.400 212.200 ;
        RECT 210.200 213.100 210.600 213.500 ;
        RECT 225.400 214.800 225.800 215.200 ;
        RECT 221.400 211.800 221.800 212.200 ;
        RECT 233.400 216.200 233.800 216.600 ;
        RECT 235.000 215.500 235.400 215.900 ;
        RECT 243.000 216.200 243.400 216.600 ;
        RECT 244.600 215.500 245.000 215.900 ;
        RECT 254.200 218.800 254.600 219.200 ;
        RECT 235.000 213.100 235.400 213.500 ;
        RECT 226.200 211.800 226.600 212.200 ;
        RECT 244.600 213.100 245.000 213.500 ;
        RECT 235.800 211.800 236.200 212.200 ;
        RECT 245.400 213.100 245.800 213.500 ;
        RECT 258.200 214.800 258.600 215.200 ;
        RECT 255.000 213.100 255.400 213.500 ;
        RECT 263.800 211.800 264.200 212.200 ;
        RECT 9.400 208.800 9.800 209.200 ;
        RECT 4.600 205.800 5.000 206.200 ;
        RECT 0.600 205.100 1.000 205.500 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 19.800 208.800 20.200 209.200 ;
        RECT 40.600 208.800 41.000 209.200 ;
        RECT 27.800 205.800 28.200 206.200 ;
        RECT 32.600 206.800 33.000 207.200 ;
        RECT 37.400 206.800 37.800 207.200 ;
        RECT 29.400 201.800 29.800 202.200 ;
        RECT 31.800 205.100 32.200 205.500 ;
        RECT 51.800 205.800 52.200 206.200 ;
        RECT 54.200 205.100 54.600 205.500 ;
        RECT 78.200 208.800 78.600 209.200 ;
        RECT 71.000 205.800 71.400 206.200 ;
        RECT 76.600 205.800 77.000 206.200 ;
        RECT 79.000 206.800 79.400 207.200 ;
        RECT 81.400 206.800 81.800 207.200 ;
        RECT 79.800 205.800 80.200 206.200 ;
        RECT 84.600 205.800 85.000 206.200 ;
        RECT 80.600 205.100 81.000 205.500 ;
        RECT 72.600 201.800 73.000 202.200 ;
        RECT 114.200 208.800 114.600 209.200 ;
        RECT 89.400 201.800 89.800 202.200 ;
        RECT 96.600 205.800 97.000 206.200 ;
        RECT 99.800 205.800 100.200 206.200 ;
        RECT 101.400 205.800 101.800 206.200 ;
        RECT 122.200 208.800 122.600 209.200 ;
        RECT 111.000 205.800 111.400 206.200 ;
        RECT 115.000 205.800 115.400 206.200 ;
        RECT 140.600 208.800 141.000 209.200 ;
        RECT 119.800 204.800 120.200 205.200 ;
        RECT 130.200 206.800 130.600 207.200 ;
        RECT 135.800 206.800 136.200 207.200 ;
        RECT 124.600 206.100 125.000 206.500 ;
        RECT 131.000 205.100 131.400 205.500 ;
        RECT 131.800 205.100 132.200 205.500 ;
        RECT 155.000 208.800 155.400 209.200 ;
        RECT 150.200 206.800 150.600 207.200 ;
        RECT 163.000 206.800 163.400 207.200 ;
        RECT 144.600 204.800 145.000 205.200 ;
        RECT 151.000 205.800 151.400 206.200 ;
        RECT 154.200 205.800 154.600 206.200 ;
        RECT 153.400 204.800 153.800 205.200 ;
        RECT 159.800 205.800 160.200 206.200 ;
        RECT 163.000 204.800 163.400 205.200 ;
        RECT 167.800 206.100 168.200 206.500 ;
        RECT 169.400 205.800 169.800 206.200 ;
        RECT 184.600 208.800 185.000 209.200 ;
        RECT 196.600 208.800 197.000 209.200 ;
        RECT 183.000 206.800 183.400 207.200 ;
        RECT 177.400 206.100 177.800 206.500 ;
        RECT 174.200 205.100 174.600 205.500 ;
        RECT 187.000 206.100 187.400 206.500 ;
        RECT 183.800 205.100 184.200 205.500 ;
        RECT 175.000 201.800 175.400 202.200 ;
        RECT 193.400 205.100 193.800 205.500 ;
        RECT 204.600 205.800 205.000 206.200 ;
        RECT 211.000 208.800 211.400 209.200 ;
        RECT 216.600 208.800 217.000 209.200 ;
        RECT 215.000 205.800 215.400 206.200 ;
        RECT 230.200 208.800 230.600 209.200 ;
        RECT 217.400 206.800 217.800 207.200 ;
        RECT 223.000 205.800 223.400 206.200 ;
        RECT 226.200 204.800 226.600 205.200 ;
        RECT 238.200 206.800 238.600 207.200 ;
        RECT 232.600 206.100 233.000 206.500 ;
        RECT 243.800 206.800 244.200 207.200 ;
        RECT 239.000 205.100 239.400 205.500 ;
        RECT 261.400 208.800 261.800 209.200 ;
        RECT 254.200 206.800 254.600 207.200 ;
        RECT 255.800 206.800 256.200 207.200 ;
        RECT 248.600 206.100 249.000 206.500 ;
        RECT 255.000 205.100 255.400 205.500 ;
        RECT 246.200 201.800 246.600 202.200 ;
        RECT 11.000 194.800 11.400 195.200 ;
        RECT 8.600 193.800 9.000 194.200 ;
        RECT 6.200 191.800 6.600 192.200 ;
        RECT 7.800 193.100 8.200 193.500 ;
        RECT 27.000 195.800 27.400 196.200 ;
        RECT 23.000 193.800 23.400 194.200 ;
        RECT 27.000 194.800 27.400 195.200 ;
        RECT 27.800 193.800 28.200 194.200 ;
        RECT 35.800 196.200 36.200 196.600 ;
        RECT 37.400 195.500 37.800 195.900 ;
        RECT 41.400 194.800 41.800 195.200 ;
        RECT 39.000 193.800 39.400 194.200 ;
        RECT 37.400 193.100 37.800 193.500 ;
        RECT 28.600 191.800 29.000 192.200 ;
        RECT 38.200 193.100 38.600 193.500 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 48.600 193.800 49.000 194.200 ;
        RECT 51.000 193.800 51.400 194.200 ;
        RECT 59.800 196.200 60.200 196.600 ;
        RECT 61.400 195.500 61.800 195.900 ;
        RECT 47.000 191.800 47.400 192.200 ;
        RECT 61.400 193.100 61.800 193.500 ;
        RECT 52.600 191.800 53.000 192.200 ;
        RECT 69.400 194.800 69.800 195.200 ;
        RECT 65.400 192.800 65.800 193.200 ;
        RECT 70.200 193.800 70.600 194.200 ;
        RECT 78.200 196.200 78.600 196.600 ;
        RECT 79.800 195.500 80.200 195.900 ;
        RECT 86.200 198.800 86.600 199.200 ;
        RECT 80.600 194.800 81.000 195.200 ;
        RECT 81.400 194.800 81.800 195.200 ;
        RECT 79.800 193.100 80.200 193.500 ;
        RECT 71.000 191.800 71.400 192.200 ;
        RECT 87.800 194.800 88.200 195.200 ;
        RECT 88.600 194.800 89.000 195.200 ;
        RECT 87.000 193.800 87.400 194.200 ;
        RECT 91.800 193.800 92.200 194.200 ;
        RECT 83.000 191.800 83.400 192.200 ;
        RECT 95.800 195.800 96.200 196.200 ;
        RECT 101.400 196.200 101.800 196.600 ;
        RECT 103.000 195.500 103.400 195.900 ;
        RECT 103.000 193.100 103.400 193.500 ;
        RECT 107.800 194.800 108.200 195.200 ;
        RECT 104.600 191.800 105.000 192.200 ;
        RECT 115.800 196.200 116.200 196.600 ;
        RECT 117.400 195.500 117.800 195.900 ;
        RECT 118.200 193.800 118.600 194.200 ;
        RECT 117.400 193.100 117.800 193.500 ;
        RECT 108.600 191.800 109.000 192.200 ;
        RECT 122.200 194.800 122.600 195.200 ;
        RECT 131.000 195.800 131.400 196.200 ;
        RECT 141.400 196.800 141.800 197.200 ;
        RECT 123.000 193.800 123.400 194.200 ;
        RECT 126.200 194.800 126.600 195.200 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 128.600 193.800 129.000 194.200 ;
        RECT 131.800 193.800 132.200 194.200 ;
        RECT 133.400 193.800 133.800 194.200 ;
        RECT 132.600 193.100 133.000 193.500 ;
        RECT 142.200 194.800 142.600 195.200 ;
        RECT 143.000 194.800 143.400 195.200 ;
        RECT 150.200 194.800 150.600 195.200 ;
        RECT 151.000 194.800 151.400 195.200 ;
        RECT 151.800 194.800 152.200 195.200 ;
        RECT 155.000 194.800 155.400 195.200 ;
        RECT 157.400 195.800 157.800 196.200 ;
        RECT 158.200 194.800 158.600 195.200 ;
        RECT 160.600 193.800 161.000 194.200 ;
        RECT 168.600 196.200 169.000 196.600 ;
        RECT 170.200 195.500 170.600 195.900 ;
        RECT 170.200 193.100 170.600 193.500 ;
        RECT 173.400 194.800 173.800 195.200 ;
        RECT 178.200 198.800 178.600 199.200 ;
        RECT 171.800 191.800 172.200 192.200 ;
        RECT 174.200 192.800 174.600 193.200 ;
        RECT 179.000 194.800 179.400 195.200 ;
        RECT 179.800 194.800 180.200 195.200 ;
        RECT 184.600 198.800 185.000 199.200 ;
        RECT 180.600 193.800 181.000 194.200 ;
        RECT 184.600 194.800 185.000 195.200 ;
        RECT 186.200 194.800 186.600 195.200 ;
        RECT 187.000 194.800 187.400 195.200 ;
        RECT 185.400 193.800 185.800 194.200 ;
        RECT 190.200 193.800 190.600 194.200 ;
        RECT 199.800 196.200 200.200 196.600 ;
        RECT 201.400 195.500 201.800 195.900 ;
        RECT 209.400 196.200 209.800 196.600 ;
        RECT 211.000 195.500 211.400 195.900 ;
        RECT 201.400 193.100 201.800 193.500 ;
        RECT 211.000 193.100 211.400 193.500 ;
        RECT 202.200 191.800 202.600 192.200 ;
        RECT 217.400 194.800 217.800 195.200 ;
        RECT 219.000 194.800 219.400 195.200 ;
        RECT 219.800 194.800 220.200 195.200 ;
        RECT 218.200 193.800 218.600 194.200 ;
        RECT 230.200 193.800 230.600 194.200 ;
        RECT 231.800 193.800 232.200 194.200 ;
        RECT 239.800 196.200 240.200 196.600 ;
        RECT 241.400 195.500 241.800 195.900 ;
        RECT 242.200 194.800 242.600 195.200 ;
        RECT 243.000 194.800 243.400 195.200 ;
        RECT 225.400 191.800 225.800 192.200 ;
        RECT 247.800 194.800 248.200 195.200 ;
        RECT 246.200 193.800 246.600 194.200 ;
        RECT 241.400 193.100 241.800 193.500 ;
        RECT 259.000 196.200 259.400 196.600 ;
        RECT 260.600 195.500 261.000 195.900 ;
        RECT 262.200 194.800 262.600 195.200 ;
        RECT 264.600 195.800 265.000 196.200 ;
        RECT 260.600 193.100 261.000 193.500 ;
        RECT 0.600 185.100 1.000 185.500 ;
        RECT 14.200 187.800 14.600 188.200 ;
        RECT 25.400 188.800 25.800 189.200 ;
        RECT 12.600 185.800 13.000 186.200 ;
        RECT 17.400 186.800 17.800 187.200 ;
        RECT 11.000 181.800 11.400 182.200 ;
        RECT 16.600 185.100 17.000 185.500 ;
        RECT 33.400 185.800 33.800 186.200 ;
        RECT 38.200 185.800 38.600 186.200 ;
        RECT 35.000 181.800 35.400 182.200 ;
        RECT 39.800 181.800 40.200 182.200 ;
        RECT 45.400 185.800 45.800 186.200 ;
        RECT 55.000 186.800 55.400 187.200 ;
        RECT 67.000 188.800 67.400 189.200 ;
        RECT 48.600 184.800 49.000 185.200 ;
        RECT 52.600 185.800 53.000 186.200 ;
        RECT 59.000 185.800 59.400 186.200 ;
        RECT 64.600 185.800 65.000 186.200 ;
        RECT 58.200 181.800 58.600 182.200 ;
        RECT 71.800 186.800 72.200 187.200 ;
        RECT 67.000 184.800 67.400 185.200 ;
        RECT 83.000 188.800 83.400 189.200 ;
        RECT 76.600 185.900 77.000 186.300 ;
        RECT 74.200 185.100 74.600 185.500 ;
        RECT 87.000 185.800 87.400 186.200 ;
        RECT 86.200 181.800 86.600 182.200 ;
        RECT 106.200 188.800 106.600 189.200 ;
        RECT 100.600 185.800 101.000 186.200 ;
        RECT 104.600 185.800 105.000 186.200 ;
        RECT 114.200 186.800 114.600 187.200 ;
        RECT 108.600 186.100 109.000 186.500 ;
        RECT 112.600 185.900 113.000 186.300 ;
        RECT 137.400 188.800 137.800 189.200 ;
        RECT 121.400 186.800 121.800 187.200 ;
        RECT 97.400 181.800 97.800 182.200 ;
        RECT 115.000 185.100 115.400 185.500 ;
        RECT 117.400 184.800 117.800 185.200 ;
        RECT 127.000 181.800 127.400 182.200 ;
        RECT 128.600 185.100 129.000 185.500 ;
        RECT 139.800 185.800 140.200 186.200 ;
        RECT 163.800 188.800 164.200 189.200 ;
        RECT 141.400 184.800 141.800 185.200 ;
        RECT 143.800 185.100 144.200 185.500 ;
        RECT 155.800 186.800 156.200 187.200 ;
        RECT 159.800 185.800 160.200 186.200 ;
        RECT 152.600 181.800 153.000 182.200 ;
        RECT 155.000 185.100 155.400 185.500 ;
        RECT 162.200 183.800 162.600 184.200 ;
        RECT 187.000 188.800 187.400 189.200 ;
        RECT 173.400 181.800 173.800 182.200 ;
        RECT 179.000 185.800 179.400 186.200 ;
        RECT 183.800 185.800 184.200 186.200 ;
        RECT 200.600 187.800 201.000 188.200 ;
        RECT 178.200 181.800 178.600 182.200 ;
        RECT 191.800 185.800 192.200 186.200 ;
        RECT 199.000 185.800 199.400 186.200 ;
        RECT 195.800 181.800 196.200 182.200 ;
        RECT 206.200 185.800 206.600 186.200 ;
        RECT 213.400 186.800 213.800 187.200 ;
        RECT 212.600 185.800 213.000 186.200 ;
        RECT 222.200 186.800 222.600 187.200 ;
        RECT 205.400 181.800 205.800 182.200 ;
        RECT 217.400 185.800 217.800 186.200 ;
        RECT 223.800 185.800 224.200 186.200 ;
        RECT 219.000 185.100 219.400 185.500 ;
        RECT 216.600 181.800 217.000 182.200 ;
        RECT 243.800 188.800 244.200 189.200 ;
        RECT 229.400 185.800 229.800 186.200 ;
        RECT 233.400 185.800 233.800 186.200 ;
        RECT 234.200 185.800 234.600 186.200 ;
        RECT 227.800 181.800 228.200 182.200 ;
        RECT 243.000 185.800 243.400 186.200 ;
        RECT 261.400 188.800 261.800 189.200 ;
        RECT 251.800 186.800 252.200 187.200 ;
        RECT 253.400 186.800 253.800 187.200 ;
        RECT 246.200 186.100 246.600 186.500 ;
        RECT 239.800 184.800 240.200 185.200 ;
        RECT 242.200 184.800 242.600 185.200 ;
        RECT 259.800 186.800 260.200 187.200 ;
        RECT 252.600 185.100 253.000 185.500 ;
        RECT 260.600 184.800 261.000 185.200 ;
        RECT 259.000 181.800 259.400 182.200 ;
        RECT 263.800 186.800 264.200 187.200 ;
        RECT 7.800 176.200 8.200 176.600 ;
        RECT 9.400 175.500 9.800 175.900 ;
        RECT 13.400 174.800 13.800 175.200 ;
        RECT 14.200 174.800 14.600 175.200 ;
        RECT 15.000 174.800 15.400 175.200 ;
        RECT 15.800 174.800 16.200 175.200 ;
        RECT 19.000 174.800 19.400 175.200 ;
        RECT 26.200 175.800 26.600 176.200 ;
        RECT 31.800 177.800 32.200 178.200 ;
        RECT 9.400 173.100 9.800 173.500 ;
        RECT 0.600 171.800 1.000 172.200 ;
        RECT 23.000 174.800 23.400 175.200 ;
        RECT 23.800 174.800 24.200 175.200 ;
        RECT 27.800 174.800 28.200 175.200 ;
        RECT 29.400 174.800 29.800 175.200 ;
        RECT 22.200 172.800 22.600 173.200 ;
        RECT 32.600 174.800 33.000 175.200 ;
        RECT 33.400 174.800 33.800 175.200 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 39.800 173.800 40.200 174.200 ;
        RECT 47.000 174.800 47.400 175.200 ;
        RECT 53.400 174.800 53.800 175.200 ;
        RECT 54.200 174.800 54.600 175.200 ;
        RECT 57.400 174.800 57.800 175.200 ;
        RECT 35.000 171.800 35.400 172.200 ;
        RECT 39.000 171.800 39.400 172.200 ;
        RECT 43.000 171.800 43.400 172.200 ;
        RECT 45.400 171.800 45.800 172.200 ;
        RECT 49.400 172.800 49.800 173.200 ;
        RECT 48.600 171.800 49.000 172.200 ;
        RECT 64.600 174.800 65.000 175.200 ;
        RECT 65.400 174.800 65.800 175.200 ;
        RECT 71.800 176.800 72.200 177.200 ;
        RECT 59.000 171.800 59.400 172.200 ;
        RECT 66.200 173.800 66.600 174.200 ;
        RECT 70.200 174.800 70.600 175.200 ;
        RECT 69.400 173.800 69.800 174.200 ;
        RECT 71.000 173.800 71.400 174.200 ;
        RECT 79.000 176.200 79.400 176.600 ;
        RECT 85.400 178.800 85.800 179.200 ;
        RECT 80.600 175.500 81.000 175.900 ;
        RECT 80.600 173.100 81.000 173.500 ;
        RECT 84.600 173.800 85.000 174.200 ;
        RECT 92.600 176.200 93.000 176.600 ;
        RECT 94.200 175.500 94.600 175.900 ;
        RECT 83.000 171.800 83.400 172.200 ;
        RECT 94.200 173.100 94.600 173.500 ;
        RECT 102.200 174.800 102.600 175.200 ;
        RECT 103.000 174.800 103.400 175.200 ;
        RECT 96.600 171.800 97.000 172.200 ;
        RECT 103.800 173.800 104.200 174.200 ;
        RECT 106.200 175.800 106.600 176.200 ;
        RECT 111.800 173.800 112.200 174.200 ;
        RECT 125.400 176.200 125.800 176.600 ;
        RECT 127.000 175.500 127.400 175.900 ;
        RECT 113.400 171.800 113.800 172.200 ;
        RECT 136.600 174.800 137.000 175.200 ;
        RECT 132.600 173.800 133.000 174.200 ;
        RECT 134.200 173.800 134.600 174.200 ;
        RECT 127.000 173.100 127.400 173.500 ;
        RECT 118.200 171.800 118.600 172.200 ;
        RECT 127.800 172.800 128.200 173.200 ;
        RECT 133.400 173.100 133.800 173.500 ;
        RECT 151.800 178.800 152.200 179.200 ;
        RECT 152.600 176.800 153.000 177.200 ;
        RECT 147.800 174.800 148.200 175.200 ;
        RECT 148.600 174.800 149.000 175.200 ;
        RECT 165.400 178.800 165.800 179.200 ;
        RECT 159.800 174.800 160.200 175.200 ;
        RECT 156.600 173.100 157.000 173.500 ;
        RECT 159.000 172.800 159.400 173.200 ;
        RECT 181.400 178.800 181.800 179.200 ;
        RECT 171.000 174.800 171.400 175.200 ;
        RECT 171.800 174.800 172.200 175.200 ;
        RECT 175.800 174.800 176.200 175.200 ;
        RECT 172.600 173.100 173.000 173.500 ;
        RECT 175.000 172.800 175.400 173.200 ;
        RECT 181.400 171.800 181.800 172.200 ;
        RECT 183.800 175.800 184.200 176.200 ;
        RECT 189.400 176.200 189.800 176.600 ;
        RECT 191.000 175.500 191.400 175.900 ;
        RECT 191.800 174.800 192.200 175.200 ;
        RECT 192.600 174.800 193.000 175.200 ;
        RECT 197.400 173.800 197.800 174.200 ;
        RECT 191.000 173.100 191.400 173.500 ;
        RECT 182.200 171.800 182.600 172.200 ;
        RECT 196.600 173.100 197.000 173.500 ;
        RECT 205.400 171.800 205.800 172.200 ;
        RECT 207.000 176.800 207.400 177.200 ;
        RECT 207.000 172.800 207.400 173.200 ;
        RECT 219.800 174.800 220.200 175.200 ;
        RECT 211.000 173.800 211.400 174.200 ;
        RECT 213.400 172.800 213.800 173.200 ;
        RECT 223.000 174.800 223.400 175.200 ;
        RECT 223.800 174.800 224.200 175.200 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 225.400 174.800 225.800 175.200 ;
        RECT 231.000 175.800 231.400 176.200 ;
        RECT 231.000 174.800 231.400 175.200 ;
        RECT 234.200 174.800 234.600 175.200 ;
        RECT 210.200 171.800 210.600 172.200 ;
        RECT 231.800 173.800 232.200 174.200 ;
        RECT 235.000 173.800 235.400 174.200 ;
        RECT 237.400 173.800 237.800 174.200 ;
        RECT 245.400 176.200 245.800 176.600 ;
        RECT 247.000 175.500 247.400 175.900 ;
        RECT 249.400 174.800 249.800 175.200 ;
        RECT 244.600 172.800 245.000 173.200 ;
        RECT 247.000 173.100 247.400 173.500 ;
        RECT 250.200 173.800 250.600 174.200 ;
        RECT 258.200 176.200 258.600 176.600 ;
        RECT 259.800 175.500 260.200 175.900 ;
        RECT 259.800 173.100 260.200 173.500 ;
        RECT 251.000 171.800 251.400 172.200 ;
        RECT 261.400 171.800 261.800 172.200 ;
        RECT 9.400 168.800 9.800 169.200 ;
        RECT 1.400 166.800 1.800 167.200 ;
        RECT 24.600 168.800 25.000 169.200 ;
        RECT 0.600 165.100 1.000 165.500 ;
        RECT 16.600 166.800 17.000 167.200 ;
        RECT 11.800 164.800 12.200 165.200 ;
        RECT 20.600 165.800 21.000 166.200 ;
        RECT 15.800 165.100 16.200 165.500 ;
        RECT 31.800 165.800 32.200 166.200 ;
        RECT 40.600 168.800 41.000 169.200 ;
        RECT 28.600 164.800 29.000 165.200 ;
        RECT 33.400 164.800 33.800 165.200 ;
        RECT 48.600 166.800 49.000 167.200 ;
        RECT 43.000 166.100 43.400 166.500 ;
        RECT 39.000 164.800 39.400 165.200 ;
        RECT 55.000 168.800 55.400 169.200 ;
        RECT 51.800 166.800 52.200 167.200 ;
        RECT 51.000 165.800 51.400 166.200 ;
        RECT 53.400 165.800 53.800 166.200 ;
        RECT 49.400 165.100 49.800 165.500 ;
        RECT 70.200 168.800 70.600 169.200 ;
        RECT 57.400 166.100 57.800 166.500 ;
        RECT 69.400 165.800 69.800 166.200 ;
        RECT 63.800 165.100 64.200 165.500 ;
        RECT 66.200 164.800 66.600 165.200 ;
        RECT 85.400 168.800 85.800 169.200 ;
        RECT 79.800 166.800 80.200 167.200 ;
        RECT 72.600 166.100 73.000 166.500 ;
        RECT 79.000 165.100 79.400 165.500 ;
        RECT 92.600 165.800 93.000 166.200 ;
        RECT 93.400 165.800 93.800 166.200 ;
        RECT 88.600 164.800 89.000 165.200 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 106.200 166.800 106.600 167.200 ;
        RECT 98.200 164.800 98.600 165.200 ;
        RECT 97.400 162.800 97.800 163.200 ;
        RECT 102.200 165.800 102.600 166.200 ;
        RECT 105.400 165.100 105.800 165.500 ;
        RECT 128.600 166.800 129.000 167.200 ;
        RECT 136.600 167.800 137.000 168.200 ;
        RECT 147.800 168.800 148.200 169.200 ;
        RECT 127.800 165.800 128.200 166.200 ;
        RECT 132.600 165.800 133.000 166.200 ;
        RECT 141.400 166.800 141.800 167.200 ;
        RECT 149.400 166.800 149.800 167.200 ;
        RECT 139.000 165.800 139.400 166.200 ;
        RECT 142.200 165.800 142.600 166.200 ;
        RECT 144.600 164.800 145.000 165.200 ;
        RECT 152.600 166.800 153.000 167.200 ;
        RECT 151.800 165.800 152.200 166.200 ;
        RECT 153.400 165.800 153.800 166.200 ;
        RECT 147.800 164.800 148.200 165.200 ;
        RECT 171.000 168.800 171.400 169.200 ;
        RECT 158.200 165.800 158.600 166.200 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 154.200 164.800 154.600 165.200 ;
        RECT 179.000 168.800 179.400 169.200 ;
        RECT 183.000 168.800 183.400 169.200 ;
        RECT 167.800 165.800 168.200 166.200 ;
        RECT 175.000 165.800 175.400 166.200 ;
        RECT 182.200 166.800 182.600 167.200 ;
        RECT 171.000 164.800 171.400 165.200 ;
        RECT 174.200 164.800 174.600 165.200 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 195.800 168.800 196.200 169.200 ;
        RECT 199.000 168.800 199.400 169.200 ;
        RECT 205.400 168.800 205.800 169.200 ;
        RECT 187.800 166.800 188.200 167.200 ;
        RECT 186.200 165.800 186.600 166.200 ;
        RECT 190.200 165.800 190.600 166.200 ;
        RECT 189.400 164.800 189.800 165.200 ;
        RECT 191.000 164.800 191.400 165.200 ;
        RECT 199.800 165.800 200.200 166.200 ;
        RECT 195.800 164.800 196.200 165.200 ;
        RECT 213.400 166.800 213.800 167.200 ;
        RECT 207.800 166.100 208.200 166.500 ;
        RECT 211.800 165.900 212.200 166.300 ;
        RECT 214.200 165.100 214.600 165.500 ;
        RECT 202.200 161.800 202.600 162.200 ;
        RECT 205.400 161.800 205.800 162.200 ;
        RECT 222.200 165.800 222.600 166.200 ;
        RECT 227.000 165.800 227.400 166.200 ;
        RECT 236.600 166.800 237.000 167.200 ;
        RECT 246.200 168.800 246.600 169.200 ;
        RECT 247.000 168.800 247.400 169.200 ;
        RECT 239.000 165.800 239.400 166.200 ;
        RECT 243.000 166.800 243.400 167.200 ;
        RECT 242.200 165.800 242.600 166.200 ;
        RECT 243.800 165.800 244.200 166.200 ;
        RECT 252.600 166.800 253.000 167.200 ;
        RECT 249.400 166.100 249.800 166.500 ;
        RECT 251.000 165.800 251.400 166.200 ;
        RECT 258.200 166.800 258.600 167.200 ;
        RECT 246.200 164.800 246.600 165.200 ;
        RECT 255.800 165.100 256.200 165.500 ;
        RECT 259.000 165.800 259.400 166.200 ;
        RECT 256.600 161.800 257.000 162.200 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 0.600 153.100 1.000 153.500 ;
        RECT 10.200 153.800 10.600 154.200 ;
        RECT 23.000 154.800 23.400 155.200 ;
        RECT 20.600 153.800 21.000 154.200 ;
        RECT 19.800 153.100 20.200 153.500 ;
        RECT 32.600 154.800 33.000 155.200 ;
        RECT 30.200 153.800 30.600 154.200 ;
        RECT 28.600 151.800 29.000 152.200 ;
        RECT 29.400 153.100 29.800 153.500 ;
        RECT 45.400 155.800 45.800 156.200 ;
        RECT 39.000 152.800 39.400 153.200 ;
        RECT 42.200 152.800 42.600 153.200 ;
        RECT 47.000 154.800 47.400 155.200 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 48.600 154.800 49.000 155.200 ;
        RECT 64.600 156.800 65.000 157.200 ;
        RECT 38.200 151.800 38.600 152.200 ;
        RECT 51.000 153.800 51.400 154.200 ;
        RECT 74.200 156.800 74.600 157.200 ;
        RECT 56.600 153.800 57.000 154.200 ;
        RECT 53.400 152.800 53.800 153.200 ;
        RECT 55.800 153.100 56.200 153.500 ;
        RECT 68.600 154.800 69.000 155.200 ;
        RECT 66.200 153.800 66.600 154.200 ;
        RECT 65.400 153.100 65.800 153.500 ;
        RECT 78.200 154.800 78.600 155.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 87.800 156.800 88.200 157.200 ;
        RECT 83.800 154.800 84.200 155.200 ;
        RECT 99.000 156.800 99.400 157.200 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 88.600 154.800 89.000 155.200 ;
        RECT 89.400 154.800 89.800 155.200 ;
        RECT 93.400 154.800 93.800 155.200 ;
        RECT 91.000 153.800 91.400 154.200 ;
        RECT 90.200 153.100 90.600 153.500 ;
        RECT 99.800 154.800 100.200 155.200 ;
        RECT 100.600 154.800 101.000 155.200 ;
        RECT 104.600 154.800 105.000 155.200 ;
        RECT 112.600 158.800 113.000 159.200 ;
        RECT 110.200 154.800 110.600 155.200 ;
        RECT 111.000 153.800 111.400 154.200 ;
        RECT 111.800 153.800 112.200 154.200 ;
        RECT 125.400 157.800 125.800 158.200 ;
        RECT 120.600 154.800 121.000 155.200 ;
        RECT 117.400 153.800 117.800 154.200 ;
        RECT 114.200 152.800 114.600 153.200 ;
        RECT 115.000 151.800 115.400 152.200 ;
        RECT 116.600 153.100 117.000 153.500 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 127.000 154.800 127.400 155.200 ;
        RECT 141.400 156.800 141.800 157.200 ;
        RECT 131.000 154.800 131.400 155.200 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 143.000 158.800 143.400 159.200 ;
        RECT 131.800 153.800 132.200 154.200 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 132.600 153.100 133.000 153.500 ;
        RECT 143.800 153.800 144.200 154.200 ;
        RECT 144.600 153.800 145.000 154.200 ;
        RECT 149.400 154.800 149.800 155.200 ;
        RECT 149.400 153.800 149.800 154.200 ;
        RECT 154.200 157.800 154.600 158.200 ;
        RECT 151.800 153.800 152.200 154.200 ;
        RECT 161.400 156.200 161.800 156.600 ;
        RECT 163.000 155.500 163.400 155.900 ;
        RECT 177.400 156.800 177.800 157.200 ;
        RECT 163.000 153.100 163.400 153.500 ;
        RECT 168.600 154.800 169.000 155.200 ;
        RECT 165.400 153.800 165.800 154.200 ;
        RECT 169.400 153.800 169.800 154.200 ;
        RECT 172.600 153.800 173.000 154.200 ;
        RECT 169.400 152.800 169.800 153.200 ;
        RECT 175.800 154.800 176.200 155.200 ;
        RECT 191.800 158.800 192.200 159.200 ;
        RECT 181.400 154.800 181.800 155.200 ;
        RECT 182.200 154.800 182.600 155.200 ;
        RECT 186.200 154.800 186.600 155.200 ;
        RECT 173.400 151.800 173.800 152.200 ;
        RECT 183.000 153.100 183.400 153.500 ;
        RECT 193.400 154.800 193.800 155.200 ;
        RECT 195.000 154.800 195.400 155.200 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 199.000 153.800 199.400 154.200 ;
        RECT 203.000 154.800 203.400 155.200 ;
        RECT 206.200 154.800 206.600 155.200 ;
        RECT 203.800 153.800 204.200 154.200 ;
        RECT 207.800 154.800 208.200 155.200 ;
        RECT 208.600 154.800 209.000 155.200 ;
        RECT 215.000 154.800 215.400 155.200 ;
        RECT 198.200 151.800 198.600 152.200 ;
        RECT 215.800 154.800 216.200 155.200 ;
        RECT 219.000 154.800 219.400 155.200 ;
        RECT 223.000 154.800 223.400 155.200 ;
        RECT 223.800 154.800 224.200 155.200 ;
        RECT 224.600 154.800 225.000 155.200 ;
        RECT 225.400 154.800 225.800 155.200 ;
        RECT 212.600 151.800 213.000 152.200 ;
        RECT 241.400 158.800 241.800 159.200 ;
        RECT 233.400 153.800 233.800 154.200 ;
        RECT 232.600 153.100 233.000 153.500 ;
        RECT 244.600 153.800 245.000 154.200 ;
        RECT 248.600 154.800 249.000 155.200 ;
        RECT 255.800 156.800 256.200 157.200 ;
        RECT 249.400 153.800 249.800 154.200 ;
        RECT 250.200 153.800 250.600 154.200 ;
        RECT 254.200 154.800 254.600 155.200 ;
        RECT 253.400 153.800 253.800 154.200 ;
        RECT 255.000 153.800 255.400 154.200 ;
        RECT 263.000 156.200 263.400 156.600 ;
        RECT 264.600 155.500 265.000 155.900 ;
        RECT 247.000 151.800 247.400 152.200 ;
        RECT 264.600 153.100 265.000 153.500 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 1.400 146.800 1.800 147.200 ;
        RECT 0.600 145.100 1.000 145.500 ;
        RECT 13.400 146.800 13.800 147.200 ;
        RECT 23.800 146.800 24.200 147.200 ;
        RECT 16.600 144.800 17.000 145.200 ;
        RECT 30.200 146.800 30.600 147.200 ;
        RECT 22.200 145.800 22.600 146.200 ;
        RECT 21.400 141.800 21.800 142.200 ;
        RECT 39.800 148.800 40.200 149.200 ;
        RECT 58.200 148.800 58.600 149.200 ;
        RECT 42.200 146.800 42.600 147.200 ;
        RECT 48.600 146.800 49.000 147.200 ;
        RECT 50.200 146.800 50.600 147.200 ;
        RECT 40.600 145.800 41.000 146.200 ;
        RECT 49.400 145.100 49.800 145.500 ;
        RECT 62.200 145.800 62.600 146.200 ;
        RECT 75.800 148.800 76.200 149.200 ;
        RECT 63.800 144.800 64.200 145.200 ;
        RECT 70.200 145.800 70.600 146.200 ;
        RECT 74.200 145.800 74.600 146.200 ;
        RECT 80.600 146.800 81.000 147.200 ;
        RECT 78.200 146.100 78.600 146.500 ;
        RECT 73.400 141.800 73.800 142.200 ;
        RECT 82.200 145.900 82.600 146.300 ;
        RECT 84.600 145.100 85.000 145.500 ;
        RECT 91.800 145.800 92.200 146.200 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 99.800 145.800 100.200 146.200 ;
        RECT 101.400 144.800 101.800 145.200 ;
        RECT 109.400 145.100 109.800 145.500 ;
        RECT 95.800 141.800 96.200 142.200 ;
        RECT 107.000 141.800 107.400 142.200 ;
        RECT 122.200 148.800 122.600 149.200 ;
        RECT 120.600 146.800 121.000 147.200 ;
        RECT 119.800 145.800 120.200 146.200 ;
        RECT 121.400 145.800 121.800 146.200 ;
        RECT 127.000 146.800 127.400 147.200 ;
        RECT 124.600 146.100 125.000 146.500 ;
        RECT 118.200 141.800 118.600 142.200 ;
        RECT 131.000 145.100 131.400 145.500 ;
        RECT 131.800 144.800 132.200 145.200 ;
        RECT 139.800 148.800 140.200 149.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 137.400 145.800 137.800 146.200 ;
        RECT 152.600 148.800 153.000 149.200 ;
        RECT 157.400 148.800 157.800 149.200 ;
        RECT 159.800 148.800 160.200 149.200 ;
        RECT 143.000 145.800 143.400 146.200 ;
        RECT 144.600 144.800 145.000 145.200 ;
        RECT 149.400 144.800 149.800 145.200 ;
        RECT 143.000 143.800 143.400 144.200 ;
        RECT 139.800 141.800 140.200 142.200 ;
        RECT 143.000 141.800 143.400 142.200 ;
        RECT 145.400 141.800 145.800 142.200 ;
        RECT 148.600 141.800 149.000 142.200 ;
        RECT 152.600 141.800 153.000 142.200 ;
        RECT 158.200 144.800 158.600 145.200 ;
        RECT 155.000 141.800 155.400 142.200 ;
        RECT 164.600 148.800 165.000 149.200 ;
        RECT 167.800 148.800 168.200 149.200 ;
        RECT 159.800 144.800 160.200 145.200 ;
        RECT 162.200 142.800 162.600 143.200 ;
        RECT 166.200 141.800 166.600 142.200 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 170.200 146.100 170.600 146.500 ;
        RECT 176.600 145.100 177.000 145.500 ;
        RECT 187.000 148.800 187.400 149.200 ;
        RECT 179.800 141.800 180.200 142.200 ;
        RECT 191.800 146.800 192.200 147.200 ;
        RECT 189.400 146.100 189.800 146.500 ;
        RECT 193.400 145.900 193.800 146.300 ;
        RECT 197.400 145.800 197.800 146.200 ;
        RECT 195.800 145.100 196.200 145.500 ;
        RECT 205.400 146.800 205.800 147.200 ;
        RECT 203.000 145.800 203.400 146.200 ;
        RECT 220.600 148.800 221.000 149.200 ;
        RECT 217.400 146.800 217.800 147.200 ;
        RECT 211.800 146.100 212.200 146.500 ;
        RECT 241.400 148.800 241.800 149.200 ;
        RECT 218.200 145.100 218.600 145.500 ;
        RECT 223.000 145.800 223.400 146.200 ;
        RECT 209.400 143.800 209.800 144.200 ;
        RECT 233.400 146.800 233.800 147.200 ;
        RECT 228.600 144.800 229.000 145.200 ;
        RECT 232.600 145.100 233.000 145.500 ;
        RECT 245.400 146.800 245.800 147.200 ;
        RECT 250.200 148.800 250.600 149.200 ;
        RECT 245.400 144.800 245.800 145.200 ;
        RECT 258.200 146.800 258.600 147.200 ;
        RECT 252.600 146.100 253.000 146.500 ;
        RECT 248.600 141.800 249.000 142.200 ;
        RECT 259.000 145.100 259.400 145.500 ;
        RECT 260.600 141.800 261.000 142.200 ;
        RECT 9.400 138.800 9.800 139.200 ;
        RECT 3.800 134.800 4.200 135.200 ;
        RECT 1.400 133.800 1.800 134.200 ;
        RECT 0.600 133.100 1.000 133.500 ;
        RECT 3.000 132.800 3.400 133.200 ;
        RECT 19.000 134.800 19.400 135.200 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 23.800 134.800 24.200 135.200 ;
        RECT 24.600 134.800 25.000 135.200 ;
        RECT 18.200 131.800 18.600 132.200 ;
        RECT 23.000 132.800 23.400 133.200 ;
        RECT 27.800 134.800 28.200 135.200 ;
        RECT 35.000 138.800 35.400 139.200 ;
        RECT 34.200 136.800 34.600 137.200 ;
        RECT 31.800 134.800 32.200 135.200 ;
        RECT 32.600 134.800 33.000 135.200 ;
        RECT 26.200 131.800 26.600 132.200 ;
        RECT 31.000 132.800 31.400 133.200 ;
        RECT 42.200 136.200 42.600 136.600 ;
        RECT 43.800 135.500 44.200 135.900 ;
        RECT 47.800 134.800 48.200 135.200 ;
        RECT 45.400 133.800 45.800 134.200 ;
        RECT 41.400 132.800 41.800 133.200 ;
        RECT 43.800 133.100 44.200 133.500 ;
        RECT 44.600 133.100 45.000 133.500 ;
        RECT 56.600 134.800 57.000 135.200 ;
        RECT 70.200 138.800 70.600 139.200 ;
        RECT 75.000 138.800 75.400 139.200 ;
        RECT 53.400 131.800 53.800 132.200 ;
        RECT 59.800 132.800 60.200 133.200 ;
        RECT 68.600 134.800 69.000 135.200 ;
        RECT 67.000 131.800 67.400 132.200 ;
        RECT 71.800 134.800 72.200 135.200 ;
        RECT 72.600 134.800 73.000 135.200 ;
        RECT 73.400 134.800 73.800 135.200 ;
        RECT 76.600 134.800 77.000 135.200 ;
        RECT 81.400 134.800 81.800 135.200 ;
        RECT 90.200 138.800 90.600 139.200 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 78.200 133.800 78.600 134.200 ;
        RECT 77.400 133.100 77.800 133.500 ;
        RECT 88.600 134.800 89.000 135.200 ;
        RECT 89.400 133.800 89.800 134.200 ;
        RECT 97.400 136.200 97.800 136.600 ;
        RECT 103.800 137.800 104.200 138.200 ;
        RECT 100.600 136.800 101.000 137.200 ;
        RECT 99.000 135.500 99.400 135.900 ;
        RECT 102.200 135.800 102.600 136.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 86.200 131.800 86.600 132.200 ;
        RECT 99.000 133.100 99.400 133.500 ;
        RECT 103.000 133.800 103.400 134.200 ;
        RECT 114.200 134.800 114.600 135.200 ;
        RECT 111.000 133.100 111.400 133.500 ;
        RECT 121.400 134.800 121.800 135.200 ;
        RECT 122.200 134.800 122.600 135.200 ;
        RECT 131.800 138.800 132.200 139.200 ;
        RECT 134.200 138.800 134.600 139.200 ;
        RECT 137.400 138.800 137.800 139.200 ;
        RECT 125.400 133.800 125.800 134.200 ;
        RECT 119.800 131.800 120.200 132.200 ;
        RECT 135.800 134.800 136.200 135.200 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 134.200 131.800 134.600 132.200 ;
        RECT 139.000 138.800 139.400 139.200 ;
        RECT 141.400 138.800 141.800 139.200 ;
        RECT 139.800 133.800 140.200 134.200 ;
        RECT 140.600 133.800 141.000 134.200 ;
        RECT 143.800 138.800 144.200 139.200 ;
        RECT 143.000 135.800 143.400 136.200 ;
        RECT 146.200 138.800 146.600 139.200 ;
        RECT 144.600 133.800 145.000 134.200 ;
        RECT 145.400 133.800 145.800 134.200 ;
        RECT 153.400 138.800 153.800 139.200 ;
        RECT 139.000 131.800 139.400 132.200 ;
        RECT 142.200 131.800 142.600 132.200 ;
        RECT 143.800 131.800 144.200 132.200 ;
        RECT 150.200 132.800 150.600 133.200 ;
        RECT 151.800 132.800 152.200 133.200 ;
        RECT 155.800 138.800 156.200 139.200 ;
        RECT 154.200 133.800 154.600 134.200 ;
        RECT 159.800 138.800 160.200 139.200 ;
        RECT 156.600 133.800 157.000 134.200 ;
        RECT 160.600 133.800 161.000 134.200 ;
        RECT 161.400 132.800 161.800 133.200 ;
        RECT 159.800 131.800 160.200 132.200 ;
        RECT 168.600 138.800 169.000 139.200 ;
        RECT 165.400 133.800 165.800 134.200 ;
        RECT 164.600 132.800 165.000 133.200 ;
        RECT 166.200 132.800 166.600 133.200 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 175.800 136.200 176.200 136.600 ;
        RECT 177.400 135.500 177.800 135.900 ;
        RECT 178.200 134.800 178.600 135.200 ;
        RECT 179.000 134.800 179.400 135.200 ;
        RECT 193.400 136.800 193.800 137.200 ;
        RECT 177.400 133.100 177.800 133.500 ;
        RECT 180.600 131.800 181.000 132.200 ;
        RECT 183.800 132.800 184.200 133.200 ;
        RECT 184.600 133.100 185.000 133.500 ;
        RECT 195.000 138.800 195.400 139.200 ;
        RECT 194.200 133.800 194.600 134.200 ;
        RECT 199.000 134.800 199.400 135.200 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 204.600 134.800 205.000 135.200 ;
        RECT 198.200 132.800 198.600 133.200 ;
        RECT 204.600 133.800 205.000 134.200 ;
        RECT 202.200 132.800 202.600 133.200 ;
        RECT 207.000 138.800 207.400 139.200 ;
        RECT 211.800 138.800 212.200 139.200 ;
        RECT 207.800 133.800 208.200 134.200 ;
        RECT 223.800 138.800 224.200 139.200 ;
        RECT 216.600 134.800 217.000 135.200 ;
        RECT 217.400 134.800 217.800 135.200 ;
        RECT 211.800 131.800 212.200 132.200 ;
        RECT 231.000 136.200 231.400 136.600 ;
        RECT 232.600 135.500 233.000 135.900 ;
        RECT 233.400 134.800 233.800 135.200 ;
        RECT 219.000 131.800 219.400 132.200 ;
        RECT 223.000 132.800 223.400 133.200 ;
        RECT 232.600 133.100 233.000 133.500 ;
        RECT 251.000 136.200 251.400 136.600 ;
        RECT 252.600 135.500 253.000 135.900 ;
        RECT 252.600 133.100 253.000 133.500 ;
        RECT 243.800 131.800 244.200 132.200 ;
        RECT 261.400 134.800 261.800 135.200 ;
        RECT 1.400 128.800 1.800 129.200 ;
        RECT 16.600 128.800 17.000 129.200 ;
        RECT 7.000 126.800 7.400 127.200 ;
        RECT 25.400 128.800 25.800 129.200 ;
        RECT 7.800 125.100 8.200 125.500 ;
        RECT 36.600 128.800 37.000 129.200 ;
        RECT 19.000 124.800 19.400 125.200 ;
        RECT 31.800 125.800 32.200 126.200 ;
        RECT 27.800 125.100 28.200 125.500 ;
        RECT 39.000 125.800 39.400 126.200 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 54.200 127.800 54.600 128.200 ;
        RECT 40.600 124.800 41.000 125.200 ;
        RECT 47.000 125.800 47.400 126.200 ;
        RECT 47.800 125.800 48.200 126.200 ;
        RECT 51.800 125.800 52.200 126.200 ;
        RECT 52.600 125.800 53.000 126.200 ;
        RECT 45.400 123.800 45.800 124.200 ;
        RECT 48.600 124.800 49.000 125.200 ;
        RECT 58.200 124.800 58.600 125.200 ;
        RECT 78.200 128.800 78.600 129.200 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 63.800 125.800 64.200 126.200 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 68.600 125.800 69.000 126.200 ;
        RECT 69.400 125.100 69.800 125.500 ;
        RECT 83.800 124.800 84.200 125.200 ;
        RECT 86.200 124.800 86.600 125.200 ;
        RECT 103.000 128.800 103.400 129.200 ;
        RECT 94.200 126.100 94.600 126.500 ;
        RECT 100.600 125.100 101.000 125.500 ;
        RECT 91.800 121.800 92.200 122.200 ;
        RECT 103.000 121.800 103.400 122.200 ;
        RECT 107.800 124.800 108.200 125.200 ;
        RECT 116.600 126.800 117.000 127.200 ;
        RECT 121.400 126.800 121.800 127.200 ;
        RECT 114.200 125.800 114.600 126.200 ;
        RECT 117.400 125.800 117.800 126.200 ;
        RECT 127.800 126.800 128.200 127.200 ;
        RECT 140.600 128.800 141.000 129.200 ;
        RECT 132.600 126.800 133.000 127.200 ;
        RECT 113.400 124.800 113.800 125.200 ;
        RECT 112.600 121.800 113.000 122.200 ;
        RECT 115.000 124.800 115.400 125.200 ;
        RECT 131.800 125.100 132.200 125.500 ;
        RECT 131.000 121.800 131.400 122.200 ;
        RECT 143.000 125.800 143.400 126.200 ;
        RECT 159.000 128.800 159.400 129.200 ;
        RECT 144.600 124.800 145.000 125.200 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 152.600 125.800 153.000 126.200 ;
        RECT 153.400 124.800 153.800 125.200 ;
        RECT 149.400 121.800 149.800 122.200 ;
        RECT 171.800 128.800 172.200 129.200 ;
        RECT 175.800 128.800 176.200 129.200 ;
        RECT 171.000 126.800 171.400 127.200 ;
        RECT 160.600 121.800 161.000 122.200 ;
        RECT 170.200 124.800 170.600 125.200 ;
        RECT 173.400 125.800 173.800 126.200 ;
        RECT 180.600 126.800 181.000 127.200 ;
        RECT 194.200 128.800 194.600 129.200 ;
        RECT 183.800 125.800 184.200 126.200 ;
        RECT 187.800 125.900 188.200 126.300 ;
        RECT 178.200 124.800 178.600 125.200 ;
        RECT 175.800 121.800 176.200 122.200 ;
        RECT 182.200 121.800 182.600 122.200 ;
        RECT 184.600 124.800 185.000 125.200 ;
        RECT 185.400 125.100 185.800 125.500 ;
        RECT 201.400 126.800 201.800 127.200 ;
        RECT 213.400 126.800 213.800 127.200 ;
        RECT 207.000 124.800 207.400 125.200 ;
        RECT 224.600 128.800 225.000 129.200 ;
        RECT 215.800 125.100 216.200 125.500 ;
        RECT 228.600 125.800 229.000 126.200 ;
        RECT 242.200 128.800 242.600 129.200 ;
        RECT 250.200 128.800 250.600 129.200 ;
        RECT 234.200 126.100 234.600 126.500 ;
        RECT 240.600 125.100 241.000 125.500 ;
        RECT 231.800 121.800 232.200 122.200 ;
        RECT 247.800 126.800 248.200 127.200 ;
        RECT 243.800 125.800 244.200 126.200 ;
        RECT 242.200 121.800 242.600 122.200 ;
        RECT 247.800 124.800 248.200 125.200 ;
        RECT 252.600 126.100 253.000 126.500 ;
        RECT 254.200 125.800 254.600 126.200 ;
        RECT 259.000 125.100 259.400 125.500 ;
        RECT 16.600 116.800 17.000 117.200 ;
        RECT 7.000 114.800 7.400 115.200 ;
        RECT 11.800 114.800 12.200 115.200 ;
        RECT 8.600 113.800 9.000 114.200 ;
        RECT 7.800 113.100 8.200 113.500 ;
        RECT 18.200 114.800 18.600 115.200 ;
        RECT 25.400 118.800 25.800 119.200 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 23.800 114.800 24.200 115.200 ;
        RECT 22.200 113.800 22.600 114.200 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 33.400 114.800 33.800 115.200 ;
        RECT 31.000 112.800 31.400 113.200 ;
        RECT 29.400 111.800 29.800 112.200 ;
        RECT 34.200 113.800 34.600 114.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 36.600 114.800 37.000 115.200 ;
        RECT 37.400 114.800 37.800 115.200 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 50.200 116.200 50.600 116.600 ;
        RECT 51.800 115.500 52.200 115.900 ;
        RECT 51.800 113.100 52.200 113.500 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 64.600 114.800 65.000 115.200 ;
        RECT 60.600 113.800 61.000 114.200 ;
        RECT 54.200 111.800 54.600 112.200 ;
        RECT 59.000 112.800 59.400 113.200 ;
        RECT 59.800 113.100 60.200 113.500 ;
        RECT 70.200 114.800 70.600 115.200 ;
        RECT 71.000 114.800 71.400 115.200 ;
        RECT 72.600 113.800 73.000 114.200 ;
        RECT 75.000 114.800 75.400 115.200 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 79.800 114.800 80.200 115.200 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 92.600 118.800 93.000 119.200 ;
        RECT 68.600 111.800 69.000 112.200 ;
        RECT 82.200 112.800 82.600 113.200 ;
        RECT 90.200 114.800 90.600 115.200 ;
        RECT 91.000 114.800 91.400 115.200 ;
        RECT 89.400 113.800 89.800 114.200 ;
        RECT 102.200 116.200 102.600 116.600 ;
        RECT 103.800 115.500 104.200 115.900 ;
        RECT 111.000 114.800 111.400 115.200 ;
        RECT 123.000 116.800 123.400 117.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 103.800 113.100 104.200 113.500 ;
        RECT 95.000 111.800 95.400 112.200 ;
        RECT 106.200 113.100 106.600 113.500 ;
        RECT 119.000 114.800 119.400 115.200 ;
        RECT 116.600 113.800 117.000 114.200 ;
        RECT 115.000 111.800 115.400 112.200 ;
        RECT 115.800 113.100 116.200 113.500 ;
        RECT 126.200 114.800 126.600 115.200 ;
        RECT 128.600 114.800 129.000 115.200 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 143.000 116.800 143.400 117.200 ;
        RECT 131.800 113.800 132.200 114.200 ;
        RECT 133.400 113.800 133.800 114.200 ;
        RECT 134.200 113.100 134.600 113.500 ;
        RECT 148.600 114.800 149.000 115.200 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 144.600 111.800 145.000 112.200 ;
        RECT 151.000 114.800 151.400 115.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 163.000 116.800 163.400 117.200 ;
        RECT 155.800 113.800 156.200 114.200 ;
        RECT 150.200 112.800 150.600 113.200 ;
        RECT 161.400 114.800 161.800 115.200 ;
        RECT 160.600 113.800 161.000 114.200 ;
        RECT 162.200 113.800 162.600 114.200 ;
        RECT 170.200 116.200 170.600 116.600 ;
        RECT 171.800 115.500 172.200 115.900 ;
        RECT 185.400 118.800 185.800 119.200 ;
        RECT 171.800 113.100 172.200 113.500 ;
        RECT 173.400 111.800 173.800 112.200 ;
        RECT 187.000 113.800 187.400 114.200 ;
        RECT 187.800 111.800 188.200 112.200 ;
        RECT 195.800 116.200 196.200 116.600 ;
        RECT 199.000 118.800 199.400 119.200 ;
        RECT 197.400 115.500 197.800 115.900 ;
        RECT 197.400 113.100 197.800 113.500 ;
        RECT 188.600 111.800 189.000 112.200 ;
        RECT 201.400 114.800 201.800 115.200 ;
        RECT 202.200 113.800 202.600 114.200 ;
        RECT 199.000 111.800 199.400 112.200 ;
        RECT 203.800 114.800 204.200 115.200 ;
        RECT 211.800 118.800 212.200 119.200 ;
        RECT 207.800 114.800 208.200 115.200 ;
        RECT 208.600 114.800 209.000 115.200 ;
        RECT 228.600 116.800 229.000 117.200 ;
        RECT 213.400 112.800 213.800 113.200 ;
        RECT 222.200 114.800 222.600 115.200 ;
        RECT 216.600 111.800 217.000 112.200 ;
        RECT 219.000 113.100 219.400 113.500 ;
        RECT 239.000 117.800 239.400 118.200 ;
        RECT 228.600 113.800 229.000 114.200 ;
        RECT 221.400 112.800 221.800 113.200 ;
        RECT 232.600 114.800 233.000 115.200 ;
        RECT 233.400 113.800 233.800 114.200 ;
        RECT 246.200 118.800 246.600 119.200 ;
        RECT 235.800 112.800 236.200 113.200 ;
        RECT 242.200 112.800 242.600 113.200 ;
        RECT 253.400 116.200 253.800 116.600 ;
        RECT 255.000 115.500 255.400 115.900 ;
        RECT 264.600 118.800 265.000 119.200 ;
        RECT 256.600 113.800 257.000 114.200 ;
        RECT 255.000 113.100 255.400 113.500 ;
        RECT 255.800 113.100 256.200 113.500 ;
        RECT 13.400 108.800 13.800 109.200 ;
        RECT 8.600 106.800 9.000 107.200 ;
        RECT 1.400 102.800 1.800 103.200 ;
        RECT 4.600 105.100 5.000 105.500 ;
        RECT 15.000 106.800 15.400 107.200 ;
        RECT 28.600 108.800 29.000 109.200 ;
        RECT 20.600 106.800 21.000 107.200 ;
        RECT 17.400 105.800 17.800 106.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 19.800 105.100 20.200 105.500 ;
        RECT 33.400 106.800 33.800 107.200 ;
        RECT 34.200 105.800 34.600 106.200 ;
        RECT 45.400 108.800 45.800 109.200 ;
        RECT 41.400 105.800 41.800 106.200 ;
        RECT 37.400 104.800 37.800 105.200 ;
        RECT 51.000 106.800 51.400 107.200 ;
        RECT 68.600 108.800 69.000 109.200 ;
        RECT 47.800 106.100 48.200 106.500 ;
        RECT 54.200 105.100 54.600 105.500 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 62.200 105.900 62.600 106.300 ;
        RECT 59.800 105.100 60.200 105.500 ;
        RECT 72.600 106.800 73.000 107.200 ;
        RECT 77.400 105.900 77.800 106.300 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 75.000 105.100 75.400 105.500 ;
        RECT 99.000 108.800 99.400 109.200 ;
        RECT 88.600 106.800 89.000 107.200 ;
        RECT 92.600 106.800 93.000 107.200 ;
        RECT 86.200 105.800 86.600 106.200 ;
        RECT 87.800 105.800 88.200 106.200 ;
        RECT 89.400 105.800 89.800 106.200 ;
        RECT 90.200 105.100 90.600 105.500 ;
        RECT 83.800 103.800 84.200 104.200 ;
        RECT 104.600 108.800 105.000 109.200 ;
        RECT 103.800 106.800 104.200 107.200 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 112.600 108.800 113.000 109.200 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 117.400 108.800 117.800 109.200 ;
        RECT 124.600 108.800 125.000 109.200 ;
        RECT 123.000 106.800 123.400 107.200 ;
        RECT 117.400 101.800 117.800 102.200 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 127.000 104.800 127.400 105.200 ;
        RECT 139.800 108.800 140.200 109.200 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 138.200 106.800 138.600 107.200 ;
        RECT 131.800 104.800 132.200 105.200 ;
        RECT 137.400 105.800 137.800 106.200 ;
        RECT 143.000 106.800 143.400 107.200 ;
        RECT 148.600 107.800 149.000 108.200 ;
        RECT 144.600 105.800 145.000 106.200 ;
        RECT 152.600 108.800 153.000 109.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 148.600 105.800 149.000 106.200 ;
        RECT 166.200 108.800 166.600 109.200 ;
        RECT 161.400 106.800 161.800 107.200 ;
        RECT 155.800 105.800 156.200 106.200 ;
        RECT 159.000 105.800 159.400 106.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 163.000 104.800 163.400 105.200 ;
        RECT 167.800 106.800 168.200 107.200 ;
        RECT 170.200 105.800 170.600 106.200 ;
        RECT 183.000 108.800 183.400 109.200 ;
        RECT 179.000 106.800 179.400 107.200 ;
        RECT 173.400 106.100 173.800 106.500 ;
        RECT 166.200 104.800 166.600 105.200 ;
        RECT 177.400 105.900 177.800 106.300 ;
        RECT 179.800 105.100 180.200 105.500 ;
        RECT 171.000 103.800 171.400 104.200 ;
        RECT 182.200 104.800 182.600 105.200 ;
        RECT 187.000 106.800 187.400 107.200 ;
        RECT 189.400 105.800 189.800 106.200 ;
        RECT 203.000 108.800 203.400 109.200 ;
        RECT 199.800 106.800 200.200 107.200 ;
        RECT 194.200 106.100 194.600 106.500 ;
        RECT 200.600 105.100 201.000 105.500 ;
        RECT 191.800 101.800 192.200 102.200 ;
        RECT 203.000 101.800 203.400 102.200 ;
        RECT 213.400 108.800 213.800 109.200 ;
        RECT 208.600 105.800 209.000 106.200 ;
        RECT 218.200 106.800 218.600 107.200 ;
        RECT 221.400 106.800 221.800 107.200 ;
        RECT 215.800 106.100 216.200 106.500 ;
        RECT 208.600 101.800 209.000 102.200 ;
        RECT 222.200 105.100 222.600 105.500 ;
        RECT 223.000 104.800 223.400 105.200 ;
        RECT 227.000 105.800 227.400 106.200 ;
        RECT 226.200 104.800 226.600 105.200 ;
        RECT 229.400 104.800 229.800 105.200 ;
        RECT 228.600 103.800 229.000 104.200 ;
        RECT 232.600 107.800 233.000 108.200 ;
        RECT 238.200 106.800 238.600 107.200 ;
        RECT 246.200 108.800 246.600 109.200 ;
        RECT 243.000 106.800 243.400 107.200 ;
        RECT 235.000 106.100 235.400 106.500 ;
        RECT 231.800 104.800 232.200 105.200 ;
        RECT 239.000 105.900 239.400 106.300 ;
        RECT 251.800 106.800 252.200 107.200 ;
        RECT 253.400 106.800 253.800 107.200 ;
        RECT 241.400 105.100 241.800 105.500 ;
        RECT 252.600 105.100 253.000 105.500 ;
        RECT 261.400 101.800 261.800 102.200 ;
        RECT 9.400 96.800 9.800 97.200 ;
        RECT 5.400 94.800 5.800 95.200 ;
        RECT 18.200 98.800 18.600 99.200 ;
        RECT 0.600 93.100 1.000 93.500 ;
        RECT 14.200 94.800 14.600 95.200 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 15.000 93.800 15.400 94.200 ;
        RECT 32.600 96.800 33.000 97.200 ;
        RECT 26.200 94.800 26.600 95.200 ;
        RECT 23.800 93.800 24.200 94.200 ;
        RECT 23.000 93.100 23.400 93.500 ;
        RECT 43.000 98.800 43.400 99.200 ;
        RECT 32.600 93.800 33.000 94.200 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 40.600 94.800 41.000 95.200 ;
        RECT 38.200 93.800 38.600 94.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 44.600 94.800 45.000 95.200 ;
        RECT 46.200 94.800 46.600 95.200 ;
        RECT 38.200 92.800 38.600 93.200 ;
        RECT 48.600 93.800 49.000 94.200 ;
        RECT 39.000 91.800 39.400 92.200 ;
        RECT 51.800 93.800 52.200 94.200 ;
        RECT 59.800 96.200 60.200 96.600 ;
        RECT 61.400 95.500 61.800 95.900 ;
        RECT 63.800 95.800 64.200 96.200 ;
        RECT 63.800 94.800 64.200 95.200 ;
        RECT 61.400 93.100 61.800 93.500 ;
        RECT 64.600 93.800 65.000 94.200 ;
        RECT 72.600 96.200 73.000 96.600 ;
        RECT 74.200 95.500 74.600 95.900 ;
        RECT 75.800 98.800 76.200 99.200 ;
        RECT 82.200 94.800 82.600 95.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 74.200 93.100 74.600 93.500 ;
        RECT 65.400 91.800 65.800 92.200 ;
        RECT 90.200 94.800 90.600 95.200 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 92.600 94.800 93.000 95.200 ;
        RECT 95.800 93.800 96.200 94.200 ;
        RECT 105.400 96.200 105.800 96.600 ;
        RECT 107.000 95.500 107.400 95.900 ;
        RECT 110.200 94.800 110.600 95.200 ;
        RECT 124.600 96.800 125.000 97.200 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 107.000 93.100 107.400 93.500 ;
        RECT 115.000 92.800 115.400 93.200 ;
        RECT 115.800 93.100 116.200 93.500 ;
        RECT 125.400 92.800 125.800 93.200 ;
        RECT 131.800 98.800 132.200 99.200 ;
        RECT 129.400 94.800 129.800 95.200 ;
        RECT 130.200 94.800 130.600 95.200 ;
        RECT 149.400 96.800 149.800 97.200 ;
        RECT 155.000 98.800 155.400 99.200 ;
        RECT 135.800 91.800 136.200 92.200 ;
        RECT 140.600 93.100 141.000 93.500 ;
        RECT 155.800 94.800 156.200 95.200 ;
        RECT 158.200 94.800 158.600 95.200 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 150.200 92.800 150.600 93.200 ;
        RECT 164.600 94.800 165.000 95.200 ;
        RECT 161.400 93.100 161.800 93.500 ;
        RECT 160.600 91.800 161.000 92.200 ;
        RECT 163.800 92.800 164.200 93.200 ;
        RECT 175.000 94.800 175.400 95.200 ;
        RECT 176.600 93.800 177.000 94.200 ;
        RECT 179.800 94.800 180.200 95.200 ;
        RECT 180.600 94.800 181.000 95.200 ;
        RECT 184.600 94.800 185.000 95.200 ;
        RECT 185.400 94.800 185.800 95.200 ;
        RECT 189.400 94.800 189.800 95.200 ;
        RECT 190.200 94.800 190.600 95.200 ;
        RECT 194.200 98.800 194.600 99.200 ;
        RECT 197.400 98.800 197.800 99.200 ;
        RECT 195.800 94.800 196.200 95.200 ;
        RECT 194.200 91.800 194.600 92.200 ;
        RECT 199.000 94.800 199.400 95.200 ;
        RECT 197.400 91.800 197.800 92.200 ;
        RECT 202.200 94.800 202.600 95.200 ;
        RECT 200.600 91.800 201.000 92.200 ;
        RECT 215.000 96.200 215.400 96.600 ;
        RECT 216.600 95.500 217.000 95.900 ;
        RECT 204.600 91.800 205.000 92.200 ;
        RECT 216.600 93.100 217.000 93.500 ;
        RECT 207.800 91.800 208.200 92.200 ;
        RECT 219.000 96.800 219.400 97.200 ;
        RECT 228.600 96.800 229.000 97.200 ;
        RECT 223.000 94.800 223.400 95.200 ;
        RECT 230.200 98.800 230.600 99.200 ;
        RECT 219.800 93.100 220.200 93.500 ;
        RECT 222.200 92.800 222.600 93.200 ;
        RECT 231.800 94.800 232.200 95.200 ;
        RECT 238.200 94.800 238.600 95.200 ;
        RECT 233.400 91.800 233.800 92.200 ;
        RECT 239.800 98.800 240.200 99.200 ;
        RECT 247.000 96.200 247.400 96.600 ;
        RECT 248.600 95.500 249.000 95.900 ;
        RECT 249.400 93.800 249.800 94.200 ;
        RECT 248.600 93.100 249.000 93.500 ;
        RECT 255.000 94.800 255.400 95.200 ;
        RECT 253.400 92.800 253.800 93.200 ;
        RECT 251.000 91.800 251.400 92.200 ;
        RECT 259.000 92.800 259.400 93.200 ;
        RECT 261.400 96.800 261.800 97.200 ;
        RECT 262.200 94.800 262.600 95.200 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 0.600 85.100 1.000 85.500 ;
        RECT 16.600 88.800 17.000 89.200 ;
        RECT 24.600 86.800 25.000 87.200 ;
        RECT 31.800 86.800 32.200 87.200 ;
        RECT 19.000 86.100 19.400 86.500 ;
        RECT 25.400 85.100 25.800 85.500 ;
        RECT 33.400 85.800 33.800 86.200 ;
        RECT 29.400 85.100 29.800 85.500 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 49.400 88.800 49.800 89.200 ;
        RECT 41.400 85.800 41.800 86.200 ;
        RECT 59.800 88.800 60.200 89.200 ;
        RECT 60.600 88.800 61.000 89.200 ;
        RECT 38.200 83.800 38.600 84.200 ;
        RECT 43.800 84.800 44.200 85.200 ;
        RECT 52.600 85.800 53.000 86.200 ;
        RECT 56.600 85.800 57.000 86.200 ;
        RECT 82.200 88.800 82.600 89.200 ;
        RECT 63.000 86.100 63.400 86.500 ;
        RECT 67.000 85.900 67.400 86.300 ;
        RECT 59.800 84.800 60.200 85.200 ;
        RECT 69.400 85.100 69.800 85.500 ;
        RECT 70.200 84.800 70.600 85.200 ;
        RECT 78.200 86.800 78.600 87.200 ;
        RECT 90.200 88.800 90.600 89.200 ;
        RECT 75.800 85.800 76.200 86.200 ;
        RECT 79.000 85.800 79.400 86.200 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 93.400 88.800 93.800 89.200 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 95.800 86.100 96.200 86.500 ;
        RECT 99.800 85.900 100.200 86.300 ;
        RECT 110.200 86.800 110.600 87.200 ;
        RECT 119.000 87.800 119.400 88.200 ;
        RECT 102.200 85.100 102.600 85.500 ;
        RECT 106.200 85.800 106.600 86.200 ;
        RECT 109.400 85.100 109.800 85.500 ;
        RECT 125.400 85.100 125.800 85.500 ;
        RECT 148.600 88.800 149.000 89.200 ;
        RECT 141.400 85.800 141.800 86.200 ;
        RECT 142.200 85.800 142.600 86.200 ;
        RECT 146.200 86.800 146.600 87.200 ;
        RECT 150.200 81.800 150.600 82.200 ;
        RECT 151.000 88.800 151.400 89.200 ;
        RECT 167.800 88.800 168.200 89.200 ;
        RECT 159.000 86.800 159.400 87.200 ;
        RECT 179.000 88.800 179.400 89.200 ;
        RECT 153.400 86.100 153.800 86.500 ;
        RECT 157.400 85.900 157.800 86.300 ;
        RECT 159.800 85.100 160.200 85.500 ;
        RECT 173.400 86.800 173.800 87.200 ;
        RECT 175.000 85.800 175.400 86.200 ;
        RECT 170.200 85.100 170.600 85.500 ;
        RECT 189.400 88.800 189.800 89.200 ;
        RECT 182.200 85.800 182.600 86.200 ;
        RECT 207.000 88.800 207.400 89.200 ;
        RECT 215.000 88.800 215.400 89.200 ;
        RECT 219.800 88.800 220.200 89.200 ;
        RECT 197.400 86.800 197.800 87.200 ;
        RECT 199.000 86.800 199.400 87.200 ;
        RECT 191.800 86.100 192.200 86.500 ;
        RECT 181.400 83.800 181.800 84.200 ;
        RECT 188.600 84.800 189.000 85.200 ;
        RECT 205.400 86.800 205.800 87.200 ;
        RECT 219.000 86.800 219.400 87.200 ;
        RECT 198.200 85.100 198.600 85.500 ;
        RECT 239.800 88.800 240.200 89.200 ;
        RECT 213.400 83.800 213.800 84.200 ;
        RECT 231.800 86.800 232.200 87.200 ;
        RECT 241.400 88.800 241.800 89.200 ;
        RECT 227.000 85.800 227.400 86.200 ;
        RECT 229.400 85.800 229.800 86.200 ;
        RECT 233.400 85.900 233.800 86.300 ;
        RECT 223.000 81.800 223.400 82.200 ;
        RECT 225.400 81.800 225.800 82.200 ;
        RECT 230.200 84.800 230.600 85.200 ;
        RECT 231.000 85.100 231.400 85.500 ;
        RECT 255.800 88.800 256.200 89.200 ;
        RECT 247.000 86.800 247.400 87.200 ;
        RECT 263.800 88.800 264.200 89.200 ;
        RECT 256.600 86.800 257.000 87.200 ;
        RECT 258.200 86.800 258.600 87.200 ;
        RECT 238.200 83.800 238.600 84.200 ;
        RECT 257.400 85.800 257.800 86.200 ;
        RECT 253.400 81.800 253.800 82.200 ;
        RECT 263.800 81.800 264.200 82.200 ;
        RECT 10.200 76.800 10.600 77.200 ;
        RECT 3.800 74.800 4.200 75.200 ;
        RECT 1.400 73.800 1.800 74.200 ;
        RECT 0.600 73.100 1.000 73.500 ;
        RECT 10.200 73.800 10.600 74.200 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 15.800 73.100 16.200 73.500 ;
        RECT 18.200 72.800 18.600 73.200 ;
        RECT 24.600 71.800 25.000 72.200 ;
        RECT 35.800 74.800 36.200 75.200 ;
        RECT 27.000 72.800 27.400 73.200 ;
        RECT 28.600 72.800 29.000 73.200 ;
        RECT 31.000 73.100 31.400 73.500 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 41.400 74.800 41.800 75.200 ;
        RECT 33.400 72.800 33.800 73.200 ;
        RECT 39.800 71.800 40.200 72.200 ;
        RECT 44.600 73.800 45.000 74.200 ;
        RECT 54.200 76.200 54.600 76.600 ;
        RECT 55.800 75.500 56.200 75.900 ;
        RECT 57.400 73.800 57.800 74.200 ;
        RECT 65.400 76.200 65.800 76.600 ;
        RECT 67.000 75.500 67.400 75.900 ;
        RECT 55.800 73.100 56.200 73.500 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 67.000 73.100 67.400 73.500 ;
        RECT 58.200 71.800 58.600 72.200 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 72.600 73.800 73.000 74.200 ;
        RECT 77.400 73.800 77.800 74.200 ;
        RECT 70.200 72.800 70.600 73.200 ;
        RECT 79.800 78.800 80.200 79.200 ;
        RECT 87.000 76.200 87.400 76.600 ;
        RECT 88.600 75.500 89.000 75.900 ;
        RECT 91.800 78.800 92.200 79.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 88.600 73.100 89.000 73.500 ;
        RECT 98.200 78.800 98.600 79.200 ;
        RECT 94.200 74.800 94.600 75.200 ;
        RECT 95.000 73.800 95.400 74.200 ;
        RECT 100.600 74.800 101.000 75.200 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 121.400 78.800 121.800 79.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 106.200 73.800 106.600 74.200 ;
        RECT 110.200 73.800 110.600 74.200 ;
        RECT 111.800 73.800 112.200 74.200 ;
        RECT 102.200 71.800 102.600 72.200 ;
        RECT 111.000 73.100 111.400 73.500 ;
        RECT 119.800 71.800 120.200 72.200 ;
        RECT 139.000 78.800 139.400 79.200 ;
        RECT 133.400 74.800 133.800 75.200 ;
        RECT 144.600 78.800 145.000 79.200 ;
        RECT 130.200 73.100 130.600 73.500 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 151.000 74.800 151.400 75.200 ;
        RECT 132.600 72.800 133.000 73.200 ;
        RECT 140.600 71.800 141.000 72.200 ;
        RECT 147.800 73.800 148.200 74.200 ;
        RECT 147.000 73.100 147.400 73.500 ;
        RECT 159.000 78.800 159.400 79.200 ;
        RECT 158.200 73.800 158.600 74.200 ;
        RECT 163.000 78.800 163.400 79.200 ;
        RECT 165.400 78.800 165.800 79.200 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 166.200 73.800 166.600 74.200 ;
        RECT 170.200 74.800 170.600 75.200 ;
        RECT 171.000 74.800 171.400 75.200 ;
        RECT 171.800 74.800 172.200 75.200 ;
        RECT 172.600 74.800 173.000 75.200 ;
        RECT 155.800 71.800 156.200 72.200 ;
        RECT 183.800 76.200 184.200 76.600 ;
        RECT 185.400 75.500 185.800 75.900 ;
        RECT 178.200 73.800 178.600 74.200 ;
        RECT 198.200 78.800 198.600 79.200 ;
        RECT 200.600 78.800 201.000 79.200 ;
        RECT 195.000 74.800 195.400 75.200 ;
        RECT 195.800 74.800 196.200 75.200 ;
        RECT 210.200 77.800 210.600 78.200 ;
        RECT 220.600 78.800 221.000 79.200 ;
        RECT 198.200 74.800 198.600 75.200 ;
        RECT 185.400 73.100 185.800 73.500 ;
        RECT 186.200 72.800 186.600 73.200 ;
        RECT 199.000 73.800 199.400 74.200 ;
        RECT 210.200 74.800 210.600 75.200 ;
        RECT 215.800 74.800 216.200 75.200 ;
        RECT 211.000 73.800 211.400 74.200 ;
        RECT 212.600 73.800 213.000 74.200 ;
        RECT 211.800 73.100 212.200 73.500 ;
        RECT 223.000 74.800 223.400 75.200 ;
        RECT 233.400 77.800 233.800 78.200 ;
        RECT 231.800 76.800 232.200 77.200 ;
        RECT 227.000 74.800 227.400 75.200 ;
        RECT 227.800 74.800 228.200 75.200 ;
        RECT 223.800 73.800 224.200 74.200 ;
        RECT 224.600 73.800 225.000 74.200 ;
        RECT 231.800 74.800 232.200 75.200 ;
        RECT 232.600 73.800 233.000 74.200 ;
        RECT 240.600 76.200 241.000 76.600 ;
        RECT 242.200 75.500 242.600 75.900 ;
        RECT 220.600 71.800 221.000 72.200 ;
        RECT 229.400 71.800 229.800 72.200 ;
        RECT 242.200 73.100 242.600 73.500 ;
        RECT 253.400 76.200 253.800 76.600 ;
        RECT 255.000 75.500 255.400 75.900 ;
        RECT 263.000 76.200 263.400 76.600 ;
        RECT 264.600 75.500 265.000 75.900 ;
        RECT 255.000 73.100 255.400 73.500 ;
        RECT 246.200 71.800 246.600 72.200 ;
        RECT 264.600 73.100 265.000 73.500 ;
        RECT 255.800 71.800 256.200 72.200 ;
        RECT 1.400 68.800 1.800 69.200 ;
        RECT 23.800 68.800 24.200 69.200 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 19.800 65.800 20.200 66.200 ;
        RECT 15.000 65.100 15.400 65.500 ;
        RECT 26.200 68.800 26.600 69.200 ;
        RECT 25.400 66.800 25.800 67.200 ;
        RECT 37.400 68.800 37.800 69.200 ;
        RECT 27.800 65.800 28.200 66.200 ;
        RECT 32.600 62.800 33.000 63.200 ;
        RECT 53.400 68.800 53.800 69.200 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 47.000 65.800 47.400 66.200 ;
        RECT 43.800 63.800 44.200 64.200 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 48.600 63.800 49.000 64.200 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 88.600 68.800 89.000 69.200 ;
        RECT 70.200 66.800 70.600 67.200 ;
        RECT 69.400 65.800 69.800 66.200 ;
        RECT 76.600 66.800 77.000 67.200 ;
        RECT 80.600 66.800 81.000 67.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 79.800 65.100 80.200 65.500 ;
        RECT 78.200 62.800 78.600 63.200 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 95.800 65.800 96.200 66.200 ;
        RECT 100.600 65.800 101.000 66.200 ;
        RECT 111.000 66.800 111.400 67.200 ;
        RECT 110.200 65.800 110.600 66.200 ;
        RECT 111.000 64.800 111.400 65.200 ;
        RECT 124.600 68.800 125.000 69.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 111.800 61.800 112.200 62.200 ;
        RECT 116.600 65.800 117.000 66.200 ;
        RECT 122.200 66.800 122.600 67.200 ;
        RECT 121.400 65.800 121.800 66.200 ;
        RECT 127.800 66.800 128.200 67.200 ;
        RECT 131.800 66.800 132.200 67.200 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 142.200 68.800 142.600 69.200 ;
        RECT 125.400 65.800 125.800 66.200 ;
        RECT 128.600 65.800 129.000 66.200 ;
        RECT 129.400 65.800 129.800 66.200 ;
        RECT 134.200 65.800 134.600 66.200 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 126.200 63.800 126.600 64.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 151.000 68.800 151.400 69.200 ;
        RECT 168.600 68.800 169.000 69.200 ;
        RECT 171.000 68.800 171.400 69.200 ;
        RECT 152.600 65.800 153.000 66.200 ;
        RECT 151.000 64.800 151.400 65.200 ;
        RECT 158.200 64.800 158.600 65.200 ;
        RECT 160.600 66.800 161.000 67.200 ;
        RECT 163.000 66.800 163.400 67.200 ;
        RECT 163.800 65.800 164.200 66.200 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 187.000 68.800 187.400 69.200 ;
        RECT 173.400 66.100 173.800 66.500 ;
        RECT 177.400 65.900 177.800 66.300 ;
        RECT 166.200 64.800 166.600 65.200 ;
        RECT 179.800 65.100 180.200 65.500 ;
        RECT 182.200 64.800 182.600 65.200 ;
        RECT 189.400 66.800 189.800 67.200 ;
        RECT 188.600 65.800 189.000 66.200 ;
        RECT 197.400 66.800 197.800 67.200 ;
        RECT 200.600 66.800 201.000 67.200 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 195.000 61.800 195.400 62.200 ;
        RECT 199.000 64.800 199.400 65.200 ;
        RECT 200.600 64.800 201.000 65.200 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 205.400 66.800 205.800 67.200 ;
        RECT 203.000 65.800 203.400 66.200 ;
        RECT 207.800 65.800 208.200 66.200 ;
        RECT 211.800 65.800 212.200 66.200 ;
        RECT 211.000 63.800 211.400 64.200 ;
        RECT 212.600 64.800 213.000 65.200 ;
        RECT 215.000 66.800 215.400 67.200 ;
        RECT 217.400 66.800 217.800 67.200 ;
        RECT 215.000 65.800 215.400 66.200 ;
        RECT 223.800 65.800 224.200 66.200 ;
        RECT 227.800 65.800 228.200 66.200 ;
        RECT 228.600 65.100 229.000 65.500 ;
        RECT 255.800 68.800 256.200 69.200 ;
        RECT 246.200 65.800 246.600 66.200 ;
        RECT 251.000 65.800 251.400 66.200 ;
        RECT 262.200 66.800 262.600 67.200 ;
        RECT 263.800 66.800 264.200 67.200 ;
        RECT 258.200 66.100 258.600 66.500 ;
        RECT 250.200 64.800 250.600 65.200 ;
        RECT 254.200 64.800 254.600 65.200 ;
        RECT 264.600 65.100 265.000 65.500 ;
        RECT 13.400 58.800 13.800 59.200 ;
        RECT 17.400 58.800 17.800 59.200 ;
        RECT 15.000 54.800 15.400 55.200 ;
        RECT 15.800 54.800 16.200 55.200 ;
        RECT 23.000 54.800 23.400 55.200 ;
        RECT 20.600 53.800 21.000 54.200 ;
        RECT 19.800 53.100 20.200 53.500 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 30.200 54.800 30.600 55.200 ;
        RECT 28.600 51.800 29.000 52.200 ;
        RECT 35.000 52.800 35.400 53.200 ;
        RECT 35.800 52.800 36.200 53.200 ;
        RECT 44.600 58.800 45.000 59.200 ;
        RECT 40.600 54.800 41.000 55.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 43.000 54.800 43.400 55.200 ;
        RECT 46.200 54.800 46.600 55.200 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 66.200 58.800 66.600 59.200 ;
        RECT 47.000 53.100 47.400 53.500 ;
        RECT 55.800 51.800 56.200 52.200 ;
        RECT 74.200 56.800 74.600 57.200 ;
        RECT 67.000 54.800 67.400 55.200 ;
        RECT 67.800 54.800 68.200 55.200 ;
        RECT 69.400 54.800 69.800 55.200 ;
        RECT 61.400 52.800 61.800 53.200 ;
        RECT 81.400 56.200 81.800 56.600 ;
        RECT 91.800 58.800 92.200 59.200 ;
        RECT 83.000 55.500 83.400 55.900 ;
        RECT 96.600 58.800 97.000 59.200 ;
        RECT 85.400 54.800 85.800 55.200 ;
        RECT 71.000 51.800 71.400 52.200 ;
        RECT 87.000 53.800 87.400 54.200 ;
        RECT 83.000 53.100 83.400 53.500 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 90.200 54.800 90.600 55.200 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 95.000 54.800 95.400 55.200 ;
        RECT 107.800 58.800 108.200 59.200 ;
        RECT 98.200 54.800 98.600 55.200 ;
        RECT 102.200 54.800 102.600 55.200 ;
        RECT 127.800 57.800 128.200 58.200 ;
        RECT 104.600 53.800 105.000 54.200 ;
        RECT 99.000 53.100 99.400 53.500 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 113.400 53.800 113.800 54.200 ;
        RECT 113.400 52.800 113.800 53.200 ;
        RECT 123.000 54.800 123.400 55.200 ;
        RECT 119.800 53.800 120.200 54.200 ;
        RECT 136.600 58.800 137.000 59.200 ;
        RECT 116.600 51.800 117.000 52.200 ;
        RECT 119.000 53.100 119.400 53.500 ;
        RECT 132.600 54.800 133.000 55.200 ;
        RECT 141.400 58.800 141.800 59.200 ;
        RECT 133.400 53.800 133.800 54.200 ;
        RECT 137.400 54.800 137.800 55.200 ;
        RECT 138.200 54.800 138.600 55.200 ;
        RECT 139.000 54.800 139.400 55.200 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 144.600 54.800 145.000 55.200 ;
        RECT 157.400 56.800 157.800 57.200 ;
        RECT 151.800 54.800 152.200 55.200 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 148.600 53.100 149.000 53.500 ;
        RECT 160.600 54.800 161.000 55.200 ;
        RECT 161.400 54.800 161.800 55.200 ;
        RECT 168.600 54.800 169.000 55.200 ;
        RECT 169.400 54.800 169.800 55.200 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 174.200 54.800 174.600 55.200 ;
        RECT 175.000 52.800 175.400 53.200 ;
        RECT 187.800 56.200 188.200 56.600 ;
        RECT 189.400 55.500 189.800 55.900 ;
        RECT 190.200 54.800 190.600 55.200 ;
        RECT 191.000 54.800 191.400 55.200 ;
        RECT 203.800 58.800 204.200 59.200 ;
        RECT 189.400 53.100 189.800 53.500 ;
        RECT 180.600 51.800 181.000 52.200 ;
        RECT 196.600 54.800 197.000 55.200 ;
        RECT 197.400 54.800 197.800 55.200 ;
        RECT 201.400 54.800 201.800 55.200 ;
        RECT 202.200 54.800 202.600 55.200 ;
        RECT 209.400 54.800 209.800 55.200 ;
        RECT 195.800 52.800 196.200 53.200 ;
        RECT 211.800 53.800 212.200 54.200 ;
        RECT 211.000 53.100 211.400 53.500 ;
        RECT 223.800 54.800 224.200 55.200 ;
        RECT 224.600 54.800 225.000 55.200 ;
        RECT 225.400 54.800 225.800 55.200 ;
        RECT 226.200 54.800 226.600 55.200 ;
        RECT 231.000 54.800 231.400 55.200 ;
        RECT 219.800 51.800 220.200 52.200 ;
        RECT 235.000 54.800 235.400 55.200 ;
        RECT 235.800 54.800 236.200 55.200 ;
        RECT 236.600 54.800 237.000 55.200 ;
        RECT 239.000 53.800 239.400 54.200 ;
        RECT 238.200 53.100 238.600 53.500 ;
        RECT 248.600 54.800 249.000 55.200 ;
        RECT 255.800 58.800 256.200 59.200 ;
        RECT 253.400 54.800 253.800 55.200 ;
        RECT 254.200 54.800 254.600 55.200 ;
        RECT 252.600 53.800 253.000 54.200 ;
        RECT 247.000 51.800 247.400 52.200 ;
        RECT 250.200 51.800 250.600 52.200 ;
        RECT 10.200 47.800 10.600 48.200 ;
        RECT 0.600 45.100 1.000 45.500 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 16.600 48.800 17.000 49.200 ;
        RECT 19.000 46.100 19.400 46.500 ;
        RECT 20.600 45.800 21.000 46.200 ;
        RECT 23.000 45.900 23.400 46.300 ;
        RECT 32.600 48.800 33.000 49.200 ;
        RECT 25.400 45.100 25.800 45.500 ;
        RECT 42.200 48.800 42.600 49.200 ;
        RECT 35.000 46.100 35.400 46.500 ;
        RECT 59.800 48.800 60.200 49.200 ;
        RECT 50.200 46.800 50.600 47.200 ;
        RECT 44.600 46.100 45.000 46.500 ;
        RECT 41.400 45.100 41.800 45.500 ;
        RECT 48.600 45.900 49.000 46.300 ;
        RECT 62.200 48.800 62.600 49.200 ;
        RECT 51.000 45.100 51.400 45.500 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 61.400 45.800 61.800 46.200 ;
        RECT 71.800 48.800 72.200 49.200 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 64.600 46.100 65.000 46.500 ;
        RECT 68.600 45.900 69.000 46.300 ;
        RECT 79.800 46.800 80.200 47.200 ;
        RECT 74.200 46.100 74.600 46.500 ;
        RECT 71.000 45.100 71.400 45.500 ;
        RECT 78.200 45.900 78.600 46.300 ;
        RECT 80.600 45.100 81.000 45.500 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 84.600 44.800 85.000 45.200 ;
        RECT 87.000 45.100 87.400 45.500 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 98.200 44.800 98.600 45.200 ;
        RECT 103.000 45.800 103.400 46.200 ;
        RECT 110.200 46.800 110.600 47.200 ;
        RECT 114.200 46.800 114.600 47.200 ;
        RECT 106.200 46.100 106.600 46.500 ;
        RECT 117.400 45.800 117.800 46.200 ;
        RECT 112.600 45.100 113.000 45.500 ;
        RECT 113.400 45.100 113.800 45.500 ;
        RECT 129.400 45.100 129.800 45.500 ;
        RECT 122.200 41.800 122.600 42.200 ;
        RECT 138.200 43.800 138.600 44.200 ;
        RECT 159.000 48.800 159.400 49.200 ;
        RECT 170.200 48.800 170.600 49.200 ;
        RECT 177.400 48.800 177.800 49.200 ;
        RECT 167.000 46.800 167.400 47.200 ;
        RECT 161.400 46.100 161.800 46.500 ;
        RECT 153.400 44.800 153.800 45.200 ;
        RECT 155.800 44.800 156.200 45.200 ;
        RECT 175.000 46.800 175.400 47.200 ;
        RECT 167.800 45.100 168.200 45.500 ;
        RECT 195.800 48.800 196.200 49.200 ;
        RECT 175.000 44.800 175.400 45.200 ;
        RECT 185.400 46.800 185.800 47.200 ;
        RECT 187.800 46.800 188.200 47.200 ;
        RECT 179.800 46.100 180.200 46.500 ;
        RECT 191.800 45.800 192.200 46.200 ;
        RECT 186.200 45.100 186.600 45.500 ;
        RECT 187.000 45.100 187.400 45.500 ;
        RECT 199.000 46.800 199.400 47.200 ;
        RECT 196.600 45.100 197.000 45.500 ;
        RECT 207.800 45.800 208.200 46.200 ;
        RECT 215.800 48.800 216.200 49.200 ;
        RECT 223.000 48.800 223.400 49.200 ;
        RECT 211.800 46.800 212.200 47.200 ;
        RECT 212.600 45.800 213.000 46.200 ;
        RECT 216.600 45.800 217.000 46.200 ;
        RECT 237.400 48.800 237.800 49.200 ;
        RECT 238.200 48.800 238.600 49.200 ;
        RECT 223.800 45.800 224.200 46.200 ;
        RECT 233.400 46.800 233.800 47.200 ;
        RECT 228.600 45.800 229.000 46.200 ;
        RECT 233.400 44.800 233.800 45.200 ;
        RECT 259.000 48.800 259.400 49.200 ;
        RECT 240.600 46.100 241.000 46.500 ;
        RECT 247.800 45.800 248.200 46.200 ;
        RECT 237.400 44.800 237.800 45.200 ;
        RECT 247.000 45.100 247.400 45.500 ;
        RECT 252.600 45.900 253.000 46.300 ;
        RECT 250.200 45.100 250.600 45.500 ;
        RECT 261.400 44.800 261.800 45.200 ;
        RECT 264.600 44.800 265.000 45.200 ;
        RECT 8.600 38.800 9.000 39.200 ;
        RECT 6.200 34.800 6.600 35.200 ;
        RECT 7.000 34.800 7.400 35.200 ;
        RECT 3.000 33.800 3.400 34.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 11.800 34.800 12.200 35.200 ;
        RECT 5.400 32.800 5.800 33.200 ;
        RECT 11.000 32.800 11.400 33.200 ;
        RECT 19.800 36.200 20.200 36.600 ;
        RECT 21.400 35.500 21.800 35.900 ;
        RECT 25.400 34.800 25.800 35.200 ;
        RECT 27.000 34.800 27.400 35.200 ;
        RECT 27.800 34.800 28.200 35.200 ;
        RECT 21.400 33.100 21.800 33.500 ;
        RECT 12.600 31.800 13.000 32.200 ;
        RECT 33.400 34.800 33.800 35.200 ;
        RECT 40.600 38.800 41.000 39.200 ;
        RECT 31.800 33.800 32.200 34.200 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 39.000 34.800 39.400 35.200 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 35.000 31.800 35.400 32.200 ;
        RECT 44.600 32.800 45.000 33.200 ;
        RECT 45.400 33.100 45.800 33.500 ;
        RECT 43.800 31.800 44.200 32.200 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 60.600 34.800 61.000 35.200 ;
        RECT 54.200 31.800 54.600 32.200 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 66.200 38.800 66.600 39.200 ;
        RECT 63.800 34.800 64.200 35.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 83.000 36.800 83.400 37.200 ;
        RECT 86.200 38.800 86.600 39.200 ;
        RECT 91.000 38.800 91.400 39.200 ;
        RECT 59.000 31.800 59.400 32.200 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 73.400 33.800 73.800 34.200 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 74.200 33.100 74.600 33.500 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 92.600 34.800 93.000 35.200 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 93.400 33.100 93.800 33.500 ;
        RECT 111.800 38.800 112.200 39.200 ;
        RECT 119.000 38.800 119.400 39.200 ;
        RECT 127.800 38.800 128.200 39.200 ;
        RECT 109.400 34.800 109.800 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 125.400 34.800 125.800 35.200 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 131.800 38.800 132.200 39.200 ;
        RECT 135.800 38.800 136.200 39.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 134.200 34.800 134.600 35.200 ;
        RECT 152.600 38.800 153.000 39.200 ;
        RECT 138.200 34.800 138.600 35.200 ;
        RECT 155.800 38.800 156.200 39.200 ;
        RECT 138.200 32.800 138.600 33.200 ;
        RECT 147.000 34.800 147.400 35.200 ;
        RECT 144.600 33.800 145.000 34.200 ;
        RECT 141.400 31.800 141.800 32.200 ;
        RECT 143.800 33.100 144.200 33.500 ;
        RECT 167.000 38.800 167.400 39.200 ;
        RECT 153.400 32.800 153.800 33.200 ;
        RECT 161.400 34.800 161.800 35.200 ;
        RECT 170.200 38.800 170.600 39.200 ;
        RECT 159.000 33.800 159.400 34.200 ;
        RECT 158.200 33.100 158.600 33.500 ;
        RECT 167.800 34.800 168.200 35.200 ;
        RECT 168.600 34.800 169.000 35.200 ;
        RECT 185.400 36.800 185.800 37.200 ;
        RECT 171.800 34.800 172.200 35.200 ;
        RECT 172.600 32.800 173.000 33.200 ;
        RECT 181.400 34.800 181.800 35.200 ;
        RECT 179.000 33.800 179.400 34.200 ;
        RECT 175.800 32.800 176.200 33.200 ;
        RECT 178.200 33.100 178.600 33.500 ;
        RECT 187.800 34.800 188.200 35.200 ;
        RECT 188.600 34.800 189.000 35.200 ;
        RECT 196.600 38.800 197.000 39.200 ;
        RECT 201.400 38.800 201.800 39.200 ;
        RECT 187.000 31.800 187.400 32.200 ;
        RECT 190.200 32.800 190.600 33.200 ;
        RECT 194.200 34.800 194.600 35.200 ;
        RECT 195.000 34.800 195.400 35.200 ;
        RECT 213.400 38.800 213.800 39.200 ;
        RECT 202.200 34.800 202.600 35.200 ;
        RECT 203.000 34.800 203.400 35.200 ;
        RECT 218.200 38.800 218.600 39.200 ;
        RECT 214.200 34.800 214.600 35.200 ;
        RECT 215.000 34.800 215.400 35.200 ;
        RECT 219.000 34.800 219.400 35.200 ;
        RECT 219.800 34.800 220.200 35.200 ;
        RECT 205.400 31.800 205.800 32.200 ;
        RECT 209.400 32.800 209.800 33.200 ;
        RECT 226.200 34.800 226.600 35.200 ;
        RECT 227.000 34.800 227.400 35.200 ;
        RECT 235.000 36.800 235.400 37.200 ;
        RECT 236.600 36.800 237.000 37.200 ;
        RECT 223.800 32.800 224.200 33.200 ;
        RECT 222.200 31.800 222.600 32.200 ;
        RECT 231.000 33.800 231.400 34.200 ;
        RECT 235.000 34.800 235.400 35.200 ;
        RECT 235.800 33.800 236.200 34.200 ;
        RECT 243.800 36.200 244.200 36.600 ;
        RECT 245.400 35.500 245.800 35.900 ;
        RECT 247.000 34.800 247.400 35.200 ;
        RECT 249.400 33.800 249.800 34.200 ;
        RECT 245.400 33.100 245.800 33.500 ;
        RECT 251.000 33.800 251.400 34.200 ;
        RECT 259.000 36.200 259.400 36.600 ;
        RECT 260.600 35.500 261.000 35.900 ;
        RECT 263.000 33.800 263.400 34.200 ;
        RECT 260.600 33.100 261.000 33.500 ;
        RECT 9.400 28.800 9.800 29.200 ;
        RECT 3.000 25.900 3.400 26.300 ;
        RECT 0.600 25.100 1.000 25.500 ;
        RECT 10.200 26.800 10.600 27.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 24.600 28.800 25.000 29.200 ;
        RECT 35.800 28.800 36.200 29.200 ;
        RECT 45.400 28.800 45.800 29.200 ;
        RECT 20.600 25.800 21.000 26.200 ;
        RECT 29.400 26.800 29.800 27.200 ;
        RECT 27.000 25.100 27.400 25.500 ;
        RECT 47.000 28.800 47.400 29.200 ;
        RECT 39.000 25.900 39.400 26.300 ;
        RECT 36.600 25.100 37.000 25.500 ;
        RECT 59.800 28.800 60.200 29.200 ;
        RECT 48.600 26.800 49.000 27.200 ;
        RECT 50.200 26.800 50.600 27.200 ;
        RECT 48.600 25.800 49.000 26.200 ;
        RECT 49.400 25.100 49.800 25.500 ;
        RECT 72.600 28.800 73.000 29.200 ;
        RECT 63.000 24.800 63.400 25.200 ;
        RECT 70.200 24.800 70.600 25.200 ;
        RECT 78.200 26.800 78.600 27.200 ;
        RECT 75.000 26.100 75.400 26.500 ;
        RECT 79.000 25.900 79.400 26.300 ;
        RECT 83.000 25.800 83.400 26.200 ;
        RECT 81.400 25.100 81.800 25.500 ;
        RECT 99.000 28.800 99.400 29.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 100.600 25.800 101.000 26.200 ;
        RECT 107.800 26.800 108.200 27.200 ;
        RECT 104.600 24.800 105.000 25.200 ;
        RECT 120.600 28.800 121.000 29.200 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 111.000 26.100 111.400 26.500 ;
        RECT 117.400 25.100 117.800 25.500 ;
        RECT 108.600 21.800 109.000 22.200 ;
        RECT 121.400 25.800 121.800 26.200 ;
        RECT 127.000 26.800 127.400 27.200 ;
        RECT 139.000 28.800 139.400 29.200 ;
        RECT 137.400 26.800 137.800 27.200 ;
        RECT 131.800 26.100 132.200 26.500 ;
        RECT 151.000 26.800 151.400 27.200 ;
        RECT 141.400 26.100 141.800 26.500 ;
        RECT 138.200 25.100 138.600 25.500 ;
        RECT 147.800 25.100 148.200 25.500 ;
        RECT 164.600 28.800 165.000 29.200 ;
        RECT 155.000 26.800 155.400 27.200 ;
        RECT 156.600 26.800 157.000 27.200 ;
        RECT 171.000 28.800 171.400 29.200 ;
        RECT 158.200 25.900 158.600 26.300 ;
        RECT 151.800 24.800 152.200 25.200 ;
        RECT 155.800 25.100 156.200 25.500 ;
        RECT 181.400 28.800 181.800 29.200 ;
        RECT 168.600 24.800 169.000 25.200 ;
        RECT 179.000 26.800 179.400 27.200 ;
        RECT 173.400 26.100 173.800 26.500 ;
        RECT 179.800 25.100 180.200 25.500 ;
        RECT 183.000 25.800 183.400 26.200 ;
        RECT 190.200 28.800 190.600 29.200 ;
        RECT 186.200 21.800 186.600 22.200 ;
        RECT 202.200 28.800 202.600 29.200 ;
        RECT 216.600 28.800 217.000 29.200 ;
        RECT 196.600 26.800 197.000 27.200 ;
        RECT 192.600 26.100 193.000 26.500 ;
        RECT 199.000 25.100 199.400 25.500 ;
        RECT 210.200 25.900 210.600 26.300 ;
        RECT 207.800 25.100 208.200 25.500 ;
        RECT 222.200 28.800 222.600 29.200 ;
        RECT 220.600 25.800 221.000 26.200 ;
        RECT 230.200 26.800 230.600 27.200 ;
        RECT 224.600 26.100 225.000 26.500 ;
        RECT 231.000 25.100 231.400 25.500 ;
        RECT 233.400 28.800 233.800 29.200 ;
        RECT 231.800 21.800 232.200 22.200 ;
        RECT 238.200 26.800 238.600 27.200 ;
        RECT 235.800 26.100 236.200 26.500 ;
        RECT 239.800 25.900 240.200 26.300 ;
        RECT 253.400 28.800 253.800 29.200 ;
        RECT 242.200 25.100 242.600 25.500 ;
        RECT 244.600 24.800 245.000 25.200 ;
        RECT 252.600 25.800 253.000 26.200 ;
        RECT 261.400 26.800 261.800 27.200 ;
        RECT 255.800 26.100 256.200 26.500 ;
        RECT 259.800 25.900 260.200 26.300 ;
        RECT 262.200 25.100 262.600 25.500 ;
        RECT 0.600 18.800 1.000 19.200 ;
        RECT 7.800 16.200 8.200 16.600 ;
        RECT 9.400 15.500 9.800 15.900 ;
        RECT 11.800 14.800 12.200 15.200 ;
        RECT 14.200 14.800 14.600 15.200 ;
        RECT 21.400 18.800 21.800 19.200 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 7.000 12.800 7.400 13.200 ;
        RECT 9.400 13.100 9.800 13.500 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 19.800 14.800 20.200 15.200 ;
        RECT 31.000 16.200 31.400 16.600 ;
        RECT 32.600 15.500 33.000 15.900 ;
        RECT 32.600 13.100 33.000 13.500 ;
        RECT 23.800 11.800 24.200 12.200 ;
        RECT 33.400 12.800 33.800 13.200 ;
        RECT 47.800 18.800 48.200 19.200 ;
        RECT 51.800 17.800 52.200 18.200 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 39.800 12.800 40.200 13.200 ;
        RECT 36.600 11.800 37.000 12.200 ;
        RECT 57.400 14.800 57.800 15.200 ;
        RECT 59.000 14.800 59.400 15.200 ;
        RECT 72.600 16.800 73.000 17.200 ;
        RECT 61.400 13.800 61.800 14.200 ;
        RECT 55.800 11.800 56.200 12.200 ;
        RECT 63.000 13.800 63.400 14.200 ;
        RECT 64.600 13.800 65.000 14.200 ;
        RECT 63.800 13.100 64.200 13.500 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 74.200 14.800 74.600 15.200 ;
        RECT 87.000 18.800 87.400 19.200 ;
        RECT 78.200 13.100 78.600 13.500 ;
        RECT 91.000 15.800 91.400 16.200 ;
        RECT 87.800 12.800 88.200 13.200 ;
        RECT 94.200 16.800 94.600 17.200 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 93.400 14.800 93.800 15.200 ;
        RECT 101.400 16.200 101.800 16.600 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 103.000 15.500 103.400 15.900 ;
        RECT 116.600 18.800 117.000 19.200 ;
        RECT 103.000 13.100 103.400 13.500 ;
        RECT 106.200 14.800 106.600 15.200 ;
        RECT 104.600 11.800 105.000 12.200 ;
        RECT 121.400 18.800 121.800 19.200 ;
        RECT 117.400 14.800 117.800 15.200 ;
        RECT 118.200 14.800 118.600 15.200 ;
        RECT 122.200 14.800 122.600 15.200 ;
        RECT 123.000 14.800 123.400 15.200 ;
        RECT 113.400 12.800 113.800 13.200 ;
        RECT 131.000 16.200 131.400 16.600 ;
        RECT 132.600 15.500 133.000 15.900 ;
        RECT 139.000 18.800 139.400 19.200 ;
        RECT 132.600 13.100 133.000 13.500 ;
        RECT 123.800 11.800 124.200 12.200 ;
        RECT 140.600 14.800 141.000 15.200 ;
        RECT 151.000 14.800 151.400 15.200 ;
        RECT 148.600 13.800 149.000 14.200 ;
        RECT 147.800 13.100 148.200 13.500 ;
        RECT 159.000 14.800 159.400 15.200 ;
        RECT 159.800 14.800 160.200 15.200 ;
        RECT 167.800 18.800 168.200 19.200 ;
        RECT 171.000 18.800 171.400 19.200 ;
        RECT 156.600 11.800 157.000 12.200 ;
        RECT 165.400 14.800 165.800 15.200 ;
        RECT 166.200 14.800 166.600 15.200 ;
        RECT 175.000 14.800 175.400 15.200 ;
        RECT 164.600 12.800 165.000 13.200 ;
        RECT 177.400 13.800 177.800 14.200 ;
        RECT 179.800 13.800 180.200 14.200 ;
        RECT 183.000 14.800 183.400 15.200 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 198.200 18.800 198.600 19.200 ;
        RECT 185.400 13.800 185.800 14.200 ;
        RECT 184.600 13.100 185.000 13.500 ;
        RECT 207.000 16.800 207.400 17.200 ;
        RECT 212.600 16.800 213.000 17.200 ;
        RECT 196.600 13.800 197.000 14.200 ;
        RECT 211.000 15.800 211.400 16.200 ;
        RECT 211.000 14.800 211.400 15.200 ;
        RECT 193.400 11.800 193.800 12.200 ;
        RECT 198.200 11.800 198.600 12.200 ;
        RECT 211.800 13.800 212.200 14.200 ;
        RECT 219.800 16.200 220.200 16.600 ;
        RECT 221.400 15.500 221.800 15.900 ;
        RECT 225.400 13.800 225.800 14.200 ;
        RECT 219.000 12.800 219.400 13.200 ;
        RECT 221.400 13.100 221.800 13.500 ;
        RECT 232.600 18.800 233.000 19.200 ;
        RECT 227.800 14.800 228.200 15.200 ;
        RECT 228.600 14.800 229.000 15.200 ;
        RECT 231.800 14.800 232.200 15.200 ;
        RECT 231.000 13.800 231.400 14.200 ;
        RECT 239.800 16.200 240.200 16.600 ;
        RECT 241.400 15.500 241.800 15.900 ;
        RECT 253.400 18.800 253.800 19.200 ;
        RECT 250.200 14.800 250.600 15.200 ;
        RECT 251.800 14.800 252.200 15.200 ;
        RECT 241.400 13.100 241.800 13.500 ;
        RECT 252.600 13.800 253.000 14.200 ;
        RECT 255.000 18.800 255.400 19.200 ;
        RECT 262.200 16.200 262.600 16.600 ;
        RECT 263.800 15.500 264.200 15.900 ;
        RECT 247.800 11.800 248.200 12.200 ;
        RECT 261.400 12.800 261.800 13.200 ;
        RECT 263.800 13.100 264.200 13.500 ;
        RECT 6.200 8.800 6.600 9.200 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 15.000 5.800 15.400 6.200 ;
        RECT 9.400 4.800 9.800 5.200 ;
        RECT 10.200 5.100 10.600 5.500 ;
        RECT 19.800 8.800 20.200 9.200 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 22.200 6.100 22.600 6.500 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 28.600 5.100 29.000 5.500 ;
        RECT 31.000 4.800 31.400 5.200 ;
        RECT 41.400 6.800 41.800 7.200 ;
        RECT 48.600 6.800 49.000 7.200 ;
        RECT 64.600 6.800 65.000 7.200 ;
        RECT 69.400 6.800 69.800 7.200 ;
        RECT 80.600 8.800 81.000 9.200 ;
        RECT 72.600 6.800 73.000 7.200 ;
        RECT 74.200 5.900 74.600 6.300 ;
        RECT 71.800 5.100 72.200 5.500 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 87.000 6.800 87.400 7.200 ;
        RECT 83.800 6.100 84.200 6.500 ;
        RECT 87.800 5.900 88.200 6.300 ;
        RECT 97.400 6.800 97.800 7.200 ;
        RECT 107.800 7.800 108.200 8.200 ;
        RECT 90.200 5.100 90.600 5.500 ;
        RECT 92.600 4.800 93.000 5.200 ;
        RECT 101.400 5.800 101.800 6.200 ;
        RECT 96.600 5.100 97.000 5.500 ;
        RECT 119.800 8.800 120.200 9.200 ;
        RECT 117.400 6.800 117.800 7.200 ;
        RECT 135.000 8.800 135.400 9.200 ;
        RECT 117.400 4.800 117.800 5.200 ;
        RECT 127.800 6.800 128.200 7.200 ;
        RECT 122.200 6.100 122.600 6.500 ;
        RECT 128.600 5.100 129.000 5.500 ;
        RECT 131.000 4.800 131.400 5.200 ;
        RECT 152.600 8.800 153.000 9.200 ;
        RECT 143.000 6.800 143.400 7.200 ;
        RECT 144.600 6.800 145.000 7.200 ;
        RECT 137.400 6.100 137.800 6.500 ;
        RECT 151.000 6.800 151.400 7.200 ;
        RECT 143.800 5.100 144.200 5.500 ;
        RECT 165.400 8.800 165.800 9.200 ;
        RECT 157.400 6.800 157.800 7.200 ;
        RECT 154.200 5.800 154.600 6.200 ;
        RECT 161.400 5.800 161.800 6.200 ;
        RECT 156.600 5.100 157.000 5.500 ;
        RECT 175.000 8.800 175.400 9.200 ;
        RECT 180.600 6.800 181.000 7.200 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 201.400 8.800 201.800 9.200 ;
        RECT 191.000 6.800 191.400 7.200 ;
        RECT 211.000 8.800 211.400 9.200 ;
        RECT 198.200 6.800 198.600 7.200 ;
        RECT 185.400 6.100 185.800 6.500 ;
        RECT 191.800 5.100 192.200 5.500 ;
        RECT 192.600 5.100 193.000 5.500 ;
        RECT 206.200 6.800 206.600 7.200 ;
        RECT 202.200 5.100 202.600 5.500 ;
        RECT 215.000 5.800 215.400 6.200 ;
        RECT 229.400 8.800 229.800 9.200 ;
        RECT 219.000 6.800 219.400 7.200 ;
        RECT 216.600 4.800 217.000 5.200 ;
        RECT 225.400 6.800 225.800 7.200 ;
        RECT 244.600 8.800 245.000 9.200 ;
        RECT 253.400 8.800 253.800 9.200 ;
        RECT 237.400 6.800 237.800 7.200 ;
        RECT 231.800 6.100 232.200 6.500 ;
        RECT 246.200 6.800 246.600 7.200 ;
        RECT 238.200 5.100 238.600 5.500 ;
        RECT 261.400 6.800 261.800 7.200 ;
        RECT 255.800 6.100 256.200 6.500 ;
        RECT 259.800 5.900 260.200 6.300 ;
        RECT 262.200 5.100 262.600 5.500 ;
      LAYER metal2 ;
        RECT 21.400 236.800 21.800 237.200 ;
        RECT 27.800 237.100 28.200 237.200 ;
        RECT 28.600 237.100 29.000 237.200 ;
        RECT 27.800 236.800 29.000 237.100 ;
        RECT 29.400 236.800 29.800 237.200 ;
        RECT 36.600 236.800 37.000 237.200 ;
        RECT 21.400 234.200 21.700 236.800 ;
        RECT 29.400 234.200 29.700 236.800 ;
        RECT 35.800 234.800 36.200 235.200 ;
        RECT 35.800 234.200 36.100 234.800 ;
        RECT 36.600 234.200 36.900 236.800 ;
        RECT 21.400 233.800 21.800 234.200 ;
        RECT 23.800 233.800 24.200 234.200 ;
        RECT 29.400 233.800 29.800 234.200 ;
        RECT 35.800 233.800 36.200 234.200 ;
        RECT 36.600 233.800 37.000 234.200 ;
        RECT 0.600 231.800 1.000 232.200 ;
        RECT 5.400 232.100 5.800 232.200 ;
        RECT 6.200 232.100 6.600 232.200 ;
        RECT 5.400 231.800 6.600 232.100 ;
        RECT 13.400 231.800 13.800 232.200 ;
        RECT 15.800 231.800 16.200 232.200 ;
        RECT 0.600 227.200 0.900 231.800 ;
        RECT 6.200 228.800 6.600 229.200 ;
        RECT 0.600 226.800 1.000 227.200 ;
        RECT 0.600 213.200 0.900 226.800 ;
        RECT 0.600 212.800 1.000 213.200 ;
        RECT 0.600 212.100 1.000 212.200 ;
        RECT 1.400 212.100 1.800 212.200 ;
        RECT 3.000 212.100 3.400 217.900 ;
        RECT 6.200 214.200 6.500 228.800 ;
        RECT 7.000 226.800 7.400 227.200 ;
        RECT 7.000 226.200 7.300 226.800 ;
        RECT 7.000 225.800 7.400 226.200 ;
        RECT 7.800 225.100 8.200 227.900 ;
        RECT 8.600 226.800 9.000 227.200 ;
        RECT 8.600 226.200 8.900 226.800 ;
        RECT 8.600 225.800 9.000 226.200 ;
        RECT 7.000 215.800 7.400 216.200 ;
        RECT 7.000 215.100 7.300 215.800 ;
        RECT 7.000 214.700 7.400 215.100 ;
        RECT 6.200 213.800 6.600 214.200 ;
        RECT 6.200 212.800 6.600 213.200 ;
        RECT 0.600 211.800 1.800 212.100 ;
        RECT 0.600 205.100 1.000 207.900 ;
        RECT 2.200 203.100 2.600 208.900 ;
        RECT 6.200 206.200 6.500 212.800 ;
        RECT 7.800 212.100 8.200 217.900 ;
        RECT 4.600 206.100 5.000 206.200 ;
        RECT 5.400 206.100 5.800 206.200 ;
        RECT 4.600 205.800 5.800 206.100 ;
        RECT 6.200 205.800 6.600 206.200 ;
        RECT 0.600 194.800 1.000 195.200 ;
        RECT 0.600 194.200 0.900 194.800 ;
        RECT 6.200 194.200 6.500 205.800 ;
        RECT 7.000 203.100 7.400 208.900 ;
        RECT 8.600 205.200 8.900 225.800 ;
        RECT 9.400 223.100 9.800 228.900 ;
        RECT 12.600 226.800 13.000 227.200 ;
        RECT 12.600 226.200 12.900 226.800 ;
        RECT 12.600 225.800 13.000 226.200 ;
        RECT 9.400 213.100 9.800 215.900 ;
        RECT 11.800 214.800 12.200 215.200 ;
        RECT 12.600 214.800 13.000 215.200 ;
        RECT 11.800 214.200 12.100 214.800 ;
        RECT 12.600 214.200 12.900 214.800 ;
        RECT 11.800 213.800 12.200 214.200 ;
        RECT 12.600 213.800 13.000 214.200 ;
        RECT 10.200 212.800 10.600 213.200 ;
        RECT 10.200 212.200 10.500 212.800 ;
        RECT 10.200 211.800 10.600 212.200 ;
        RECT 9.400 209.100 9.800 209.200 ;
        RECT 10.200 209.100 10.600 209.200 ;
        RECT 9.400 208.800 10.600 209.100 ;
        RECT 13.400 208.200 13.700 231.800 ;
        RECT 15.800 229.200 16.100 231.800 ;
        RECT 14.200 223.100 14.600 228.900 ;
        RECT 15.800 228.800 16.200 229.200 ;
        RECT 19.000 227.800 19.400 228.200 ;
        RECT 22.200 227.800 22.600 228.200 ;
        RECT 19.000 227.200 19.300 227.800 ;
        RECT 18.200 226.800 18.600 227.200 ;
        RECT 19.000 226.800 19.400 227.200 ;
        RECT 18.200 226.200 18.500 226.800 ;
        RECT 17.400 225.800 17.800 226.200 ;
        RECT 18.200 225.800 18.600 226.200 ;
        RECT 20.600 225.800 21.000 226.200 ;
        RECT 17.400 225.200 17.700 225.800 ;
        RECT 15.000 224.800 15.400 225.200 ;
        RECT 17.400 224.800 17.800 225.200 ;
        RECT 15.000 215.200 15.300 224.800 ;
        RECT 16.600 224.100 17.000 224.200 ;
        RECT 17.400 224.100 17.800 224.200 ;
        RECT 16.600 223.800 17.800 224.100 ;
        RECT 15.000 214.800 15.400 215.200 ;
        RECT 14.200 214.100 14.600 214.200 ;
        RECT 15.000 214.100 15.400 214.200 ;
        RECT 14.200 213.800 15.400 214.100 ;
        RECT 15.800 212.100 16.200 212.200 ;
        RECT 18.200 212.100 18.600 217.900 ;
        RECT 19.800 214.800 20.200 215.200 ;
        RECT 19.000 213.800 19.400 214.200 ;
        RECT 15.800 211.800 16.900 212.100 ;
        RECT 15.000 208.800 15.400 209.200 ;
        RECT 13.400 207.800 13.800 208.200 ;
        RECT 15.000 207.200 15.300 208.800 ;
        RECT 16.600 208.200 16.900 211.800 ;
        RECT 19.000 208.200 19.300 213.800 ;
        RECT 19.800 209.200 20.100 214.800 ;
        RECT 20.600 211.200 20.900 225.800 ;
        RECT 21.400 224.800 21.800 225.200 ;
        RECT 20.600 210.800 21.000 211.200 ;
        RECT 19.800 208.800 20.200 209.200 ;
        RECT 16.600 207.800 17.000 208.200 ;
        RECT 17.400 207.800 17.800 208.200 ;
        RECT 19.000 207.800 19.400 208.200 ;
        RECT 10.200 206.800 10.600 207.200 ;
        RECT 12.600 206.800 13.000 207.200 ;
        RECT 13.400 207.100 13.800 207.200 ;
        RECT 14.200 207.100 14.600 207.200 ;
        RECT 13.400 206.800 14.600 207.100 ;
        RECT 15.000 206.800 15.400 207.200 ;
        RECT 10.200 205.200 10.500 206.800 ;
        RECT 11.000 206.100 11.400 206.200 ;
        RECT 11.800 206.100 12.200 206.200 ;
        RECT 11.000 205.800 12.200 206.100 ;
        RECT 8.600 204.800 9.000 205.200 ;
        RECT 10.200 204.800 10.600 205.200 ;
        RECT 0.600 193.800 1.000 194.200 ;
        RECT 6.200 193.800 6.600 194.200 ;
        RECT 7.800 193.100 8.200 195.900 ;
        RECT 8.600 194.800 9.000 195.200 ;
        RECT 8.600 194.200 8.900 194.800 ;
        RECT 8.600 193.800 9.000 194.200 ;
        RECT 6.200 191.800 6.600 192.200 ;
        RECT 9.400 192.100 9.800 197.900 ;
        RECT 11.000 195.100 11.400 195.200 ;
        RECT 11.800 195.100 12.200 195.200 ;
        RECT 11.000 194.800 12.200 195.100 ;
        RECT 6.200 191.200 6.500 191.800 ;
        RECT 6.200 190.800 6.600 191.200 ;
        RECT 0.600 185.100 1.000 187.900 ;
        RECT 2.200 183.100 2.600 188.900 ;
        RECT 6.200 186.200 6.500 190.800 ;
        RECT 12.600 190.100 12.900 206.800 ;
        RECT 16.600 206.200 16.900 207.800 ;
        RECT 16.600 205.800 17.000 206.200 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 13.400 204.200 13.700 204.800 ;
        RECT 13.400 203.800 13.800 204.200 ;
        RECT 14.200 192.100 14.600 197.900 ;
        RECT 15.000 192.800 15.400 193.200 ;
        RECT 13.400 190.100 13.800 190.200 ;
        RECT 12.600 189.800 13.800 190.100 ;
        RECT 3.800 185.800 4.200 186.200 ;
        RECT 6.200 185.800 6.600 186.200 ;
        RECT 3.800 185.200 4.100 185.800 ;
        RECT 3.800 184.800 4.200 185.200 ;
        RECT 0.600 172.100 1.000 172.200 ;
        RECT 1.400 172.100 1.800 172.200 ;
        RECT 3.000 172.100 3.400 177.900 ;
        RECT 0.600 171.800 1.800 172.100 ;
        RECT 0.600 165.100 1.000 167.900 ;
        RECT 1.400 166.800 1.800 167.200 ;
        RECT 0.600 153.100 1.000 155.900 ;
        RECT 0.600 145.100 1.000 147.900 ;
        RECT 1.400 147.200 1.700 166.800 ;
        RECT 2.200 163.100 2.600 168.900 ;
        RECT 3.800 166.800 4.200 167.200 ;
        RECT 3.800 166.200 4.100 166.800 ;
        RECT 3.800 165.800 4.200 166.200 ;
        RECT 6.200 165.200 6.500 185.800 ;
        RECT 7.000 183.100 7.400 188.900 ;
        RECT 10.200 186.800 10.600 187.200 ;
        RECT 10.200 186.200 10.500 186.800 ;
        RECT 10.200 185.800 10.600 186.200 ;
        RECT 11.800 186.100 12.200 186.200 ;
        RECT 12.600 186.100 13.000 186.200 ;
        RECT 11.800 185.800 13.000 186.100 ;
        RECT 11.800 184.800 12.200 185.200 ;
        RECT 11.000 181.800 11.400 182.200 ;
        RECT 7.000 174.700 7.400 175.100 ;
        RECT 7.000 171.100 7.300 174.700 ;
        RECT 7.800 172.100 8.200 177.900 ;
        RECT 8.600 174.800 9.000 175.200 ;
        RECT 8.600 174.200 8.900 174.800 ;
        RECT 8.600 173.800 9.000 174.200 ;
        RECT 9.400 173.100 9.800 175.900 ;
        RECT 11.000 175.200 11.300 181.800 ;
        RECT 11.800 179.200 12.100 184.800 ;
        RECT 11.800 178.800 12.200 179.200 ;
        RECT 13.400 175.200 13.700 189.800 ;
        RECT 14.200 187.800 14.600 188.200 ;
        RECT 14.200 187.200 14.500 187.800 ;
        RECT 14.200 186.800 14.600 187.200 ;
        RECT 15.000 186.200 15.300 192.800 ;
        RECT 15.000 185.800 15.400 186.200 ;
        RECT 15.800 185.800 16.200 186.200 ;
        RECT 15.800 185.200 16.100 185.800 ;
        RECT 15.800 184.800 16.200 185.200 ;
        RECT 16.600 185.100 17.000 187.900 ;
        RECT 17.400 187.200 17.700 207.800 ;
        RECT 19.000 195.200 19.300 207.800 ;
        RECT 21.400 207.100 21.700 224.800 ;
        RECT 20.600 206.800 21.700 207.100 ;
        RECT 22.200 224.200 22.500 227.800 ;
        RECT 23.000 225.100 23.400 227.900 ;
        RECT 22.200 223.800 22.600 224.200 ;
        RECT 20.600 206.200 20.900 206.800 ;
        RECT 22.200 206.200 22.500 223.800 ;
        RECT 23.000 212.100 23.400 217.900 ;
        RECT 23.800 214.200 24.100 233.800 ;
        RECT 43.800 233.100 44.200 235.900 ;
        RECT 44.600 234.800 45.000 235.200 ;
        RECT 44.600 234.200 44.900 234.800 ;
        RECT 44.600 233.800 45.000 234.200 ;
        RECT 42.200 231.800 42.600 232.200 ;
        RECT 45.400 232.100 45.800 237.900 ;
        RECT 47.000 234.800 47.400 235.200 ;
        RECT 24.600 223.100 25.000 228.900 ;
        RECT 25.400 228.800 25.800 229.200 ;
        RECT 25.400 228.200 25.700 228.800 ;
        RECT 25.400 227.800 25.800 228.200 ;
        RECT 26.200 225.800 26.600 226.200 ;
        RECT 26.200 224.200 26.500 225.800 ;
        RECT 26.200 223.800 26.600 224.200 ;
        RECT 29.400 223.100 29.800 228.900 ;
        RECT 31.800 228.800 32.200 229.200 ;
        RECT 31.800 227.200 32.100 228.800 ;
        RECT 42.200 228.200 42.500 231.800 ;
        RECT 38.200 227.800 38.600 228.200 ;
        RECT 42.200 227.800 42.600 228.200 ;
        RECT 38.200 227.200 38.500 227.800 ;
        RECT 31.800 226.800 32.200 227.200 ;
        RECT 38.200 226.800 38.600 227.200 ;
        RECT 39.800 226.800 40.200 227.200 ;
        RECT 42.200 226.800 42.600 227.200 ;
        RECT 43.000 226.800 43.400 227.200 ;
        RECT 39.800 226.200 40.100 226.800 ;
        RECT 42.200 226.200 42.500 226.800 ;
        RECT 43.000 226.200 43.300 226.800 ;
        RECT 31.800 226.100 32.200 226.200 ;
        RECT 32.600 226.100 33.000 226.200 ;
        RECT 31.800 225.800 33.000 226.100 ;
        RECT 33.400 226.100 33.800 226.200 ;
        RECT 34.200 226.100 34.600 226.200 ;
        RECT 33.400 225.800 34.600 226.100 ;
        RECT 38.200 225.800 38.600 226.200 ;
        RECT 39.800 225.800 40.200 226.200 ;
        RECT 42.200 225.800 42.600 226.200 ;
        RECT 43.000 225.800 43.400 226.200 ;
        RECT 45.400 226.100 45.800 226.200 ;
        RECT 46.200 226.100 46.600 226.200 ;
        RECT 45.400 225.800 46.600 226.100 ;
        RECT 33.400 225.200 33.700 225.800 ;
        RECT 33.400 224.800 33.800 225.200 ;
        RECT 30.200 223.800 30.600 224.200 ;
        RECT 34.200 224.100 34.600 224.200 ;
        RECT 35.000 224.100 35.400 224.200 ;
        RECT 34.200 223.800 35.400 224.100 ;
        RECT 30.200 219.200 30.500 223.800 ;
        RECT 30.200 218.800 30.600 219.200 ;
        RECT 26.200 216.800 26.600 217.200 ;
        RECT 23.800 213.800 24.200 214.200 ;
        RECT 24.600 213.100 25.000 215.900 ;
        RECT 25.400 212.800 25.800 213.200 ;
        RECT 25.400 212.200 25.700 212.800 ;
        RECT 25.400 211.800 25.800 212.200 ;
        RECT 25.400 206.200 25.700 211.800 ;
        RECT 26.200 206.200 26.500 216.800 ;
        RECT 27.800 212.100 28.200 217.900 ;
        RECT 30.200 214.200 30.500 218.800 ;
        RECT 31.800 215.800 32.200 216.200 ;
        RECT 31.800 215.100 32.100 215.800 ;
        RECT 31.800 214.700 32.200 215.100 ;
        RECT 30.200 213.800 30.600 214.200 ;
        RECT 30.200 211.800 30.600 212.200 ;
        RECT 32.600 212.100 33.000 217.900 ;
        RECT 34.200 213.100 34.600 215.900 ;
        RECT 36.600 215.800 37.000 216.200 ;
        RECT 37.400 215.800 37.800 216.200 ;
        RECT 36.600 215.200 36.900 215.800 ;
        RECT 36.600 214.800 37.000 215.200 ;
        RECT 37.400 214.200 37.700 215.800 ;
        RECT 35.000 213.800 35.400 214.200 ;
        RECT 37.400 213.800 37.800 214.200 ;
        RECT 35.000 213.200 35.300 213.800 ;
        RECT 35.000 212.800 35.400 213.200 ;
        RECT 37.400 212.800 37.800 213.200 ;
        RECT 30.200 206.200 30.500 211.800 ;
        RECT 20.600 205.800 21.000 206.200 ;
        RECT 21.400 205.800 21.800 206.200 ;
        RECT 22.200 205.800 22.600 206.200 ;
        RECT 25.400 205.800 25.800 206.200 ;
        RECT 26.200 205.800 26.600 206.200 ;
        RECT 27.000 206.100 27.400 206.200 ;
        RECT 27.800 206.100 28.200 206.200 ;
        RECT 27.000 205.800 28.200 206.100 ;
        RECT 30.200 205.800 30.600 206.200 ;
        RECT 31.000 205.800 31.400 206.200 ;
        RECT 19.000 194.800 19.400 195.200 ;
        RECT 19.800 194.800 20.200 195.200 ;
        RECT 19.000 193.200 19.300 194.800 ;
        RECT 19.800 194.200 20.100 194.800 ;
        RECT 20.600 194.200 20.900 205.800 ;
        RECT 21.400 203.200 21.700 205.800 ;
        RECT 21.400 202.800 21.800 203.200 ;
        RECT 23.800 201.800 24.200 202.200 ;
        RECT 22.200 194.800 22.600 195.200 ;
        RECT 19.800 193.800 20.200 194.200 ;
        RECT 20.600 193.800 21.000 194.200 ;
        RECT 21.400 193.800 21.800 194.200 ;
        RECT 19.000 192.800 19.400 193.200 ;
        RECT 19.000 191.800 19.400 192.200 ;
        RECT 17.400 186.800 17.800 187.200 ;
        RECT 14.200 176.800 14.600 177.200 ;
        RECT 14.200 175.200 14.500 176.800 ;
        RECT 11.000 174.800 11.400 175.200 ;
        RECT 13.400 174.800 13.800 175.200 ;
        RECT 14.200 174.800 14.600 175.200 ;
        RECT 15.000 174.800 15.400 175.200 ;
        RECT 15.800 174.800 16.200 175.200 ;
        RECT 13.400 173.800 13.800 174.200 ;
        RECT 7.000 170.800 8.100 171.100 ;
        RECT 6.200 164.800 6.600 165.200 ;
        RECT 2.200 152.100 2.600 157.900 ;
        RECT 6.200 155.200 6.500 164.800 ;
        RECT 7.000 163.100 7.400 168.900 ;
        RECT 7.800 168.200 8.100 170.800 ;
        RECT 9.400 170.800 9.800 171.200 ;
        RECT 9.400 169.200 9.700 170.800 ;
        RECT 9.400 168.800 9.800 169.200 ;
        RECT 7.800 167.800 8.200 168.200 ;
        RECT 11.800 167.100 12.200 167.200 ;
        RECT 12.600 167.100 13.000 167.200 ;
        RECT 11.800 166.800 13.000 167.100 ;
        RECT 11.800 165.800 12.200 166.200 ;
        RECT 11.800 165.200 12.100 165.800 ;
        RECT 11.800 164.800 12.200 165.200 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 1.400 146.800 1.800 147.200 ;
        RECT 0.600 133.100 1.000 135.900 ;
        RECT 1.400 134.200 1.700 146.800 ;
        RECT 2.200 143.100 2.600 148.900 ;
        RECT 3.800 148.200 4.100 154.800 ;
        RECT 7.000 152.100 7.400 157.900 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 10.200 154.200 10.500 156.800 ;
        RECT 11.800 156.100 12.200 156.200 ;
        RECT 12.600 156.100 13.000 156.200 ;
        RECT 11.800 155.800 13.000 156.100 ;
        RECT 10.200 153.800 10.600 154.200 ;
        RECT 10.200 150.200 10.500 153.800 ;
        RECT 11.000 151.800 11.400 152.200 ;
        RECT 10.200 149.800 10.600 150.200 ;
        RECT 9.400 149.100 9.800 149.200 ;
        RECT 10.200 149.100 10.600 149.200 ;
        RECT 3.800 147.800 4.200 148.200 ;
        RECT 3.800 145.800 4.200 146.200 ;
        RECT 3.800 145.200 4.100 145.800 ;
        RECT 3.800 144.800 4.200 145.200 ;
        RECT 7.000 143.100 7.400 148.900 ;
        RECT 9.400 148.800 10.600 149.100 ;
        RECT 10.200 147.800 10.600 148.200 ;
        RECT 10.200 147.200 10.500 147.800 ;
        RECT 10.200 146.800 10.600 147.200 ;
        RECT 10.200 145.100 10.600 145.200 ;
        RECT 11.000 145.100 11.300 151.800 ;
        RECT 11.800 146.200 12.100 155.800 ;
        RECT 12.600 154.100 13.000 154.200 ;
        RECT 13.400 154.100 13.700 173.800 ;
        RECT 15.000 170.200 15.300 174.800 ;
        RECT 15.800 171.200 16.100 174.800 ;
        RECT 17.400 174.200 17.700 186.800 ;
        RECT 18.200 183.100 18.600 188.900 ;
        RECT 19.000 175.200 19.300 191.800 ;
        RECT 19.800 187.800 20.200 188.200 ;
        RECT 19.800 186.200 20.100 187.800 ;
        RECT 19.800 185.800 20.200 186.200 ;
        RECT 19.000 174.800 19.400 175.200 ;
        RECT 17.400 173.800 17.800 174.200 ;
        RECT 15.800 170.800 16.200 171.200 ;
        RECT 15.000 169.800 15.400 170.200 ;
        RECT 14.200 167.100 14.600 167.200 ;
        RECT 15.000 167.100 15.400 167.200 ;
        RECT 14.200 166.800 15.400 167.100 ;
        RECT 14.200 166.100 14.600 166.200 ;
        RECT 15.000 166.100 15.400 166.200 ;
        RECT 14.200 165.800 15.400 166.100 ;
        RECT 15.800 165.100 16.200 167.900 ;
        RECT 16.600 166.800 17.000 167.200 ;
        RECT 16.600 165.200 16.900 166.800 ;
        RECT 16.600 164.800 17.000 165.200 ;
        RECT 17.400 163.100 17.800 168.900 ;
        RECT 20.600 167.200 20.900 193.800 ;
        RECT 21.400 193.200 21.700 193.800 ;
        RECT 21.400 192.800 21.800 193.200 ;
        RECT 21.400 178.200 21.700 192.800 ;
        RECT 22.200 190.200 22.500 194.800 ;
        RECT 23.000 193.800 23.400 194.200 ;
        RECT 23.000 193.200 23.300 193.800 ;
        RECT 23.000 192.800 23.400 193.200 ;
        RECT 22.200 189.800 22.600 190.200 ;
        RECT 23.000 183.100 23.400 188.900 ;
        RECT 21.400 177.800 21.800 178.200 ;
        RECT 23.800 176.100 24.100 201.800 ;
        RECT 26.200 196.200 26.500 205.800 ;
        RECT 31.000 202.200 31.300 205.800 ;
        RECT 31.800 205.100 32.200 207.900 ;
        RECT 32.600 206.800 33.000 207.200 ;
        RECT 32.600 205.200 32.900 206.800 ;
        RECT 32.600 204.800 33.000 205.200 ;
        RECT 33.400 203.100 33.800 208.900 ;
        RECT 35.000 207.800 35.400 208.200 ;
        RECT 35.000 206.200 35.300 207.800 ;
        RECT 37.400 207.200 37.700 212.800 ;
        RECT 38.200 212.200 38.500 225.800 ;
        RECT 40.600 221.800 41.000 222.200 ;
        RECT 39.000 214.800 39.400 215.200 ;
        RECT 38.200 211.800 38.600 212.200 ;
        RECT 37.400 206.800 37.800 207.200 ;
        RECT 35.000 205.800 35.400 206.200 ;
        RECT 38.200 203.100 38.600 208.900 ;
        RECT 39.000 204.200 39.300 214.800 ;
        RECT 40.600 210.200 40.900 221.800 ;
        RECT 45.400 218.200 45.700 225.800 ;
        RECT 47.000 225.100 47.300 234.800 ;
        RECT 49.400 233.800 49.800 234.200 ;
        RECT 49.400 230.200 49.700 233.800 ;
        RECT 50.200 232.100 50.600 237.900 ;
        RECT 53.400 236.800 53.800 237.200 ;
        RECT 53.400 234.200 53.700 236.800 ;
        RECT 65.400 235.800 65.800 236.200 ;
        RECT 65.400 235.200 65.700 235.800 ;
        RECT 62.200 235.100 62.600 235.200 ;
        RECT 61.400 234.800 62.600 235.100 ;
        RECT 65.400 234.800 65.800 235.200 ;
        RECT 53.400 233.800 53.800 234.200 ;
        RECT 60.600 232.800 61.000 233.200 ;
        RECT 60.600 232.200 60.900 232.800 ;
        RECT 52.600 231.800 53.000 232.200 ;
        RECT 60.600 231.800 61.000 232.200 ;
        RECT 49.400 229.800 49.800 230.200 ;
        RECT 47.800 227.800 48.200 228.200 ;
        RECT 47.800 227.200 48.100 227.800 ;
        RECT 52.600 227.200 52.900 231.800 ;
        RECT 47.800 226.800 48.200 227.200 ;
        RECT 52.600 226.800 53.000 227.200 ;
        RECT 50.200 226.100 50.600 226.200 ;
        RECT 51.000 226.100 51.400 226.200 ;
        RECT 50.200 225.800 51.400 226.100 ;
        RECT 54.200 225.100 54.600 227.900 ;
        RECT 46.200 224.800 47.300 225.100 ;
        RECT 46.200 219.200 46.500 224.800 ;
        RECT 55.800 223.100 56.200 228.900 ;
        RECT 59.800 227.800 60.200 228.200 ;
        RECT 56.600 226.800 57.000 227.200 ;
        RECT 57.400 226.800 57.800 227.200 ;
        RECT 47.000 221.800 47.400 222.200 ;
        RECT 51.800 221.800 52.200 222.200 ;
        RECT 46.200 218.800 46.600 219.200 ;
        RECT 45.400 217.800 45.800 218.200 ;
        RECT 45.400 216.200 45.700 217.800 ;
        RECT 43.000 215.800 43.400 216.200 ;
        RECT 45.400 215.800 45.800 216.200 ;
        RECT 43.000 215.200 43.300 215.800 ;
        RECT 47.000 215.200 47.300 221.800 ;
        RECT 41.400 214.800 41.800 215.200 ;
        RECT 43.000 214.800 43.400 215.200 ;
        RECT 43.800 214.800 44.200 215.200 ;
        RECT 44.600 214.800 45.000 215.200 ;
        RECT 47.000 214.800 47.400 215.200 ;
        RECT 41.400 214.200 41.700 214.800 ;
        RECT 41.400 213.800 41.800 214.200 ;
        RECT 40.600 209.800 41.000 210.200 ;
        RECT 40.600 209.100 41.000 209.200 ;
        RECT 41.400 209.100 41.800 209.200 ;
        RECT 40.600 208.800 41.800 209.100 ;
        RECT 42.200 208.100 42.600 208.200 ;
        RECT 43.000 208.100 43.400 208.200 ;
        RECT 42.200 207.800 43.400 208.100 ;
        RECT 43.800 206.200 44.100 214.800 ;
        RECT 44.600 214.200 44.900 214.800 ;
        RECT 44.600 213.800 45.000 214.200 ;
        RECT 48.600 213.100 49.000 215.900 ;
        RECT 49.400 213.800 49.800 214.200 ;
        RECT 49.400 213.200 49.700 213.800 ;
        RECT 49.400 212.800 49.800 213.200 ;
        RECT 50.200 212.100 50.600 217.900 ;
        RECT 51.000 213.800 51.400 214.200 ;
        RECT 51.000 213.200 51.300 213.800 ;
        RECT 51.000 212.800 51.400 213.200 ;
        RECT 45.400 208.800 45.800 209.200 ;
        RECT 47.000 208.800 47.400 209.200 ;
        RECT 40.600 206.100 41.000 206.200 ;
        RECT 41.400 206.100 41.800 206.200 ;
        RECT 40.600 205.800 41.800 206.100 ;
        RECT 42.200 205.800 42.600 206.200 ;
        RECT 43.800 205.800 44.200 206.200 ;
        RECT 39.000 203.800 39.400 204.200 ;
        RECT 29.400 201.800 29.800 202.200 ;
        RECT 31.000 201.800 31.400 202.200 ;
        RECT 27.000 196.800 27.400 197.200 ;
        RECT 27.000 196.200 27.300 196.800 ;
        RECT 24.600 195.800 25.000 196.200 ;
        RECT 26.200 195.800 26.600 196.200 ;
        RECT 27.000 195.800 27.400 196.200 ;
        RECT 24.600 192.200 24.900 195.800 ;
        RECT 27.000 194.800 27.400 195.200 ;
        RECT 27.800 194.800 28.200 195.200 ;
        RECT 27.000 192.200 27.300 194.800 ;
        RECT 27.800 194.200 28.100 194.800 ;
        RECT 27.800 193.800 28.200 194.200 ;
        RECT 28.600 192.800 29.000 193.200 ;
        RECT 28.600 192.200 28.900 192.800 ;
        RECT 24.600 191.800 25.000 192.200 ;
        RECT 27.000 191.800 27.400 192.200 ;
        RECT 28.600 191.800 29.000 192.200 ;
        RECT 27.000 189.800 27.400 190.200 ;
        RECT 25.400 189.100 25.800 189.200 ;
        RECT 26.200 189.100 26.600 189.200 ;
        RECT 25.400 188.800 26.600 189.100 ;
        RECT 27.000 186.200 27.300 189.800 ;
        RECT 27.800 188.100 28.200 188.200 ;
        RECT 28.600 188.100 29.000 188.200 ;
        RECT 27.800 187.800 29.000 188.100 ;
        RECT 29.400 186.200 29.700 201.800 ;
        RECT 31.000 192.100 31.400 197.900 ;
        RECT 32.600 197.800 33.000 198.200 ;
        RECT 31.800 188.800 32.200 189.200 ;
        RECT 31.800 188.200 32.100 188.800 ;
        RECT 31.800 187.800 32.200 188.200 ;
        RECT 26.200 185.800 26.600 186.200 ;
        RECT 27.000 185.800 27.400 186.200 ;
        RECT 29.400 185.800 29.800 186.200 ;
        RECT 26.200 185.100 26.500 185.800 ;
        RECT 27.000 185.100 27.400 185.200 ;
        RECT 26.200 184.800 27.400 185.100 ;
        RECT 23.000 175.800 24.100 176.100 ;
        RECT 26.200 176.800 26.600 177.200 ;
        RECT 26.200 176.200 26.500 176.800 ;
        RECT 26.200 175.800 26.600 176.200 ;
        RECT 23.000 175.200 23.300 175.800 ;
        RECT 23.000 174.800 23.400 175.200 ;
        RECT 23.800 174.800 24.200 175.200 ;
        RECT 25.400 174.800 25.800 175.200 ;
        RECT 23.800 174.200 24.100 174.800 ;
        RECT 23.800 173.800 24.200 174.200 ;
        RECT 21.400 173.100 21.800 173.200 ;
        RECT 22.200 173.100 22.600 173.200 ;
        RECT 21.400 172.800 22.600 173.100 ;
        RECT 25.400 171.200 25.700 174.800 ;
        RECT 25.400 170.800 25.800 171.200 ;
        RECT 24.600 169.100 25.000 169.200 ;
        RECT 25.400 169.100 25.800 169.200 ;
        RECT 20.600 166.800 21.000 167.200 ;
        RECT 20.600 165.800 21.000 166.200 ;
        RECT 20.600 165.200 20.900 165.800 ;
        RECT 20.600 164.800 21.000 165.200 ;
        RECT 22.200 163.100 22.600 168.900 ;
        RECT 24.600 168.800 25.800 169.100 ;
        RECT 12.600 153.800 13.700 154.100 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 19.000 154.200 19.300 154.800 ;
        RECT 19.000 153.800 19.400 154.200 ;
        RECT 13.400 148.200 13.700 153.800 ;
        RECT 19.800 153.100 20.200 155.900 ;
        RECT 20.600 154.800 21.000 155.200 ;
        RECT 20.600 154.200 20.900 154.800 ;
        RECT 20.600 153.800 21.000 154.200 ;
        RECT 21.400 152.100 21.800 157.900 ;
        RECT 25.400 157.800 25.800 158.200 ;
        RECT 25.400 155.200 25.700 157.800 ;
        RECT 23.000 154.800 23.400 155.200 ;
        RECT 25.400 154.800 25.800 155.200 ;
        RECT 23.000 153.200 23.300 154.800 ;
        RECT 23.000 152.800 23.400 153.200 ;
        RECT 26.200 152.100 26.600 157.900 ;
        RECT 15.800 149.800 16.200 150.200 ;
        RECT 13.400 147.800 13.800 148.200 ;
        RECT 13.400 147.100 13.800 147.200 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 13.400 146.800 14.600 147.100 ;
        RECT 15.000 146.800 15.400 147.200 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 13.400 146.100 13.800 146.200 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 13.400 145.800 14.600 146.100 ;
        RECT 10.200 144.800 11.300 145.100 ;
        RECT 14.200 144.800 14.600 145.200 ;
        RECT 14.200 144.200 14.500 144.800 ;
        RECT 14.200 143.800 14.600 144.200 ;
        RECT 9.400 140.800 9.800 141.200 ;
        RECT 9.400 139.200 9.700 140.800 ;
        RECT 9.400 138.800 9.800 139.200 ;
        RECT 1.400 133.800 1.800 134.200 ;
        RECT 1.400 129.200 1.700 133.800 ;
        RECT 2.200 132.100 2.600 137.900 ;
        RECT 3.800 135.100 4.200 135.200 ;
        RECT 4.600 135.100 5.000 135.200 ;
        RECT 3.800 134.800 5.000 135.100 ;
        RECT 3.000 132.800 3.400 133.200 ;
        RECT 1.400 128.800 1.800 129.200 ;
        RECT 3.000 107.200 3.300 132.800 ;
        RECT 7.000 132.100 7.400 137.900 ;
        RECT 11.800 135.800 12.200 136.200 ;
        RECT 14.200 135.800 14.600 136.200 ;
        RECT 11.800 135.200 12.100 135.800 ;
        RECT 11.800 134.800 12.200 135.200 ;
        RECT 12.600 134.800 13.000 135.200 ;
        RECT 12.600 134.200 12.900 134.800 ;
        RECT 14.200 134.200 14.500 135.800 ;
        RECT 15.000 135.200 15.300 146.800 ;
        RECT 15.800 135.200 16.100 149.800 ;
        RECT 18.200 148.800 18.600 149.200 ;
        RECT 18.200 147.200 18.500 148.800 ;
        RECT 23.800 147.800 24.200 148.200 ;
        RECT 23.800 147.200 24.100 147.800 ;
        RECT 18.200 147.100 18.600 147.200 ;
        RECT 19.000 147.100 19.400 147.200 ;
        RECT 18.200 146.800 19.400 147.100 ;
        RECT 19.800 146.800 20.200 147.200 ;
        RECT 23.800 146.800 24.200 147.200 ;
        RECT 19.800 146.200 20.100 146.800 ;
        RECT 16.600 145.800 17.000 146.200 ;
        RECT 18.200 146.100 18.600 146.200 ;
        RECT 19.000 146.100 19.400 146.200 ;
        RECT 18.200 145.800 19.400 146.100 ;
        RECT 19.800 145.800 20.200 146.200 ;
        RECT 22.200 145.800 22.600 146.200 ;
        RECT 16.600 145.200 16.900 145.800 ;
        RECT 16.600 144.800 17.000 145.200 ;
        RECT 16.600 144.200 16.900 144.800 ;
        RECT 16.600 143.800 17.000 144.200 ;
        RECT 21.400 141.800 21.800 142.200 ;
        RECT 19.800 137.800 20.200 138.200 ;
        RECT 19.800 135.200 20.100 137.800 ;
        RECT 21.400 135.200 21.700 141.800 ;
        RECT 22.200 141.200 22.500 145.800 ;
        RECT 27.000 142.200 27.300 184.800 ;
        RECT 31.000 178.100 31.400 178.200 ;
        RECT 31.800 178.100 32.200 178.200 ;
        RECT 31.000 177.800 32.200 178.100 ;
        RECT 29.400 176.800 29.800 177.200 ;
        RECT 29.400 175.200 29.700 176.800 ;
        RECT 30.200 175.800 30.600 176.200 ;
        RECT 30.200 175.200 30.500 175.800 ;
        RECT 32.600 175.200 32.900 197.800 ;
        RECT 34.200 195.800 34.600 196.200 ;
        RECT 34.200 195.200 34.500 195.800 ;
        RECT 34.200 194.800 34.600 195.200 ;
        RECT 34.200 191.800 34.600 192.200 ;
        RECT 35.800 192.100 36.200 197.900 ;
        RECT 39.000 197.200 39.300 203.800 ;
        RECT 39.000 196.800 39.400 197.200 ;
        RECT 36.600 194.800 37.000 195.200 ;
        RECT 36.600 194.200 36.900 194.800 ;
        RECT 36.600 193.800 37.000 194.200 ;
        RECT 37.400 193.100 37.800 195.900 ;
        RECT 38.200 193.100 38.600 195.900 ;
        RECT 39.000 193.800 39.400 194.200 ;
        RECT 33.400 185.800 33.800 186.200 ;
        RECT 33.400 185.200 33.700 185.800 ;
        RECT 33.400 184.800 33.800 185.200 ;
        RECT 34.200 176.200 34.500 191.800 ;
        RECT 39.000 191.200 39.300 193.800 ;
        RECT 39.800 192.100 40.200 197.900 ;
        RECT 41.400 194.800 41.800 195.200 ;
        RECT 41.400 194.200 41.700 194.800 ;
        RECT 41.400 193.800 41.800 194.200 ;
        RECT 39.000 190.800 39.400 191.200 ;
        RECT 42.200 190.200 42.500 205.800 ;
        RECT 43.800 199.200 44.100 205.800 ;
        RECT 43.800 198.800 44.200 199.200 ;
        RECT 44.600 192.100 45.000 197.900 ;
        RECT 42.200 189.800 42.600 190.200 ;
        RECT 43.000 188.800 43.400 189.200 ;
        RECT 38.200 186.800 38.600 187.200 ;
        RECT 40.600 186.800 41.000 187.200 ;
        RECT 38.200 186.200 38.500 186.800 ;
        RECT 40.600 186.200 40.900 186.800 ;
        RECT 43.000 186.200 43.300 188.800 ;
        RECT 43.800 187.800 44.200 188.200 ;
        RECT 43.800 187.200 44.100 187.800 ;
        RECT 43.800 186.800 44.200 187.200 ;
        RECT 45.400 186.200 45.700 208.800 ;
        RECT 47.000 208.200 47.300 208.800 ;
        RECT 47.000 207.800 47.400 208.200 ;
        RECT 47.800 205.800 48.200 206.200 ;
        RECT 48.600 206.100 49.000 206.200 ;
        RECT 49.400 206.100 49.800 206.200 ;
        RECT 48.600 205.800 49.800 206.100 ;
        RECT 47.800 205.200 48.100 205.800 ;
        RECT 47.800 204.800 48.200 205.200 ;
        RECT 49.400 201.800 49.800 202.200 ;
        RECT 49.400 198.200 49.700 201.800 ;
        RECT 49.400 197.800 49.800 198.200 ;
        RECT 47.800 195.800 48.200 196.200 ;
        RECT 47.000 191.800 47.400 192.200 ;
        RECT 47.000 187.200 47.300 191.800 ;
        RECT 47.800 189.200 48.100 195.800 ;
        RECT 51.000 194.200 51.300 212.800 ;
        RECT 51.800 206.200 52.100 221.800 ;
        RECT 56.600 219.100 56.900 226.800 ;
        RECT 57.400 226.200 57.700 226.800 ;
        RECT 57.400 225.800 57.800 226.200 ;
        RECT 55.800 218.800 56.900 219.100 ;
        RECT 59.800 223.200 60.100 227.800 ;
        RECT 59.800 222.800 60.200 223.200 ;
        RECT 60.600 223.100 61.000 228.900 ;
        RECT 53.400 214.800 53.800 215.200 ;
        RECT 53.400 214.200 53.700 214.800 ;
        RECT 53.400 213.800 53.800 214.200 ;
        RECT 55.000 212.100 55.400 217.900 ;
        RECT 55.800 217.200 56.100 218.800 ;
        RECT 55.800 216.800 56.200 217.200 ;
        RECT 55.800 210.200 56.100 216.800 ;
        RECT 59.000 211.800 59.400 212.200 ;
        RECT 55.800 209.800 56.200 210.200 ;
        RECT 58.200 209.800 58.600 210.200 ;
        RECT 52.600 206.800 53.000 207.200 ;
        RECT 51.800 205.800 52.200 206.200 ;
        RECT 52.600 195.200 52.900 206.800 ;
        RECT 54.200 205.100 54.600 207.900 ;
        RECT 55.800 203.100 56.200 208.900 ;
        RECT 56.600 206.100 57.000 206.200 ;
        RECT 57.400 206.100 57.800 206.200 ;
        RECT 56.600 205.800 57.800 206.100 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 52.600 194.800 53.000 195.200 ;
        RECT 48.600 194.100 49.000 194.200 ;
        RECT 49.400 194.100 49.800 194.200 ;
        RECT 48.600 193.800 49.800 194.100 ;
        RECT 51.000 193.800 51.400 194.200 ;
        RECT 47.800 188.800 48.200 189.200 ;
        RECT 47.000 186.800 47.400 187.200 ;
        RECT 50.200 186.800 50.600 187.200 ;
        RECT 47.000 186.200 47.300 186.800 ;
        RECT 50.200 186.200 50.500 186.800 ;
        RECT 35.000 186.100 35.400 186.200 ;
        RECT 35.800 186.100 36.200 186.200 ;
        RECT 35.000 185.800 36.200 186.100 ;
        RECT 36.600 185.800 37.000 186.200 ;
        RECT 38.200 185.800 38.600 186.200 ;
        RECT 40.600 185.800 41.000 186.200 ;
        RECT 41.400 185.800 41.800 186.200 ;
        RECT 42.200 185.800 42.600 186.200 ;
        RECT 43.000 185.800 43.400 186.200 ;
        RECT 45.400 185.800 45.800 186.200 ;
        RECT 47.000 185.800 47.400 186.200 ;
        RECT 49.400 185.800 49.800 186.200 ;
        RECT 50.200 185.800 50.600 186.200 ;
        RECT 36.600 184.200 36.900 185.800 ;
        RECT 41.400 184.200 41.700 185.800 ;
        RECT 42.200 185.200 42.500 185.800 ;
        RECT 42.200 184.800 42.600 185.200 ;
        RECT 48.600 184.800 49.000 185.200 ;
        RECT 48.600 184.200 48.900 184.800 ;
        RECT 36.600 183.800 37.000 184.200 ;
        RECT 41.400 183.800 41.800 184.200 ;
        RECT 48.600 183.800 49.000 184.200 ;
        RECT 49.400 182.200 49.700 185.800 ;
        RECT 51.800 184.200 52.100 194.800 ;
        RECT 52.600 192.100 53.000 192.200 ;
        RECT 53.400 192.100 53.800 192.200 ;
        RECT 55.000 192.100 55.400 197.900 ;
        RECT 57.400 195.800 57.800 196.200 ;
        RECT 57.400 195.200 57.700 195.800 ;
        RECT 57.400 194.800 57.800 195.200 ;
        RECT 58.200 194.200 58.500 209.800 ;
        RECT 58.200 193.800 58.600 194.200 ;
        RECT 52.600 191.800 53.800 192.100 ;
        RECT 52.600 186.200 52.900 191.800 ;
        RECT 53.400 190.800 53.800 191.200 ;
        RECT 52.600 185.800 53.000 186.200 ;
        RECT 51.800 183.800 52.200 184.200 ;
        RECT 35.000 181.800 35.400 182.200 ;
        RECT 39.800 181.800 40.200 182.200 ;
        RECT 49.400 181.800 49.800 182.200 ;
        RECT 33.400 176.100 33.800 176.200 ;
        RECT 34.200 176.100 34.600 176.200 ;
        RECT 33.400 175.800 34.600 176.100 ;
        RECT 27.800 175.100 28.200 175.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 27.800 174.800 29.000 175.100 ;
        RECT 29.400 174.800 29.800 175.200 ;
        RECT 30.200 174.800 30.600 175.200 ;
        RECT 31.800 174.800 32.200 175.200 ;
        RECT 32.600 174.800 33.000 175.200 ;
        RECT 33.400 174.800 33.800 175.200 ;
        RECT 35.000 175.100 35.300 181.800 ;
        RECT 38.200 175.800 38.600 176.200 ;
        RECT 39.800 176.100 40.100 181.800 ;
        RECT 43.000 177.800 43.400 178.200 ;
        RECT 39.800 175.800 40.900 176.100 ;
        RECT 35.800 175.100 36.200 175.200 ;
        RECT 35.000 174.800 36.200 175.100 ;
        RECT 27.800 172.200 28.100 174.800 ;
        RECT 27.800 171.800 28.200 172.200 ;
        RECT 31.800 167.200 32.100 174.800 ;
        RECT 33.400 174.200 33.700 174.800 ;
        RECT 33.400 173.800 33.800 174.200 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 37.400 173.800 37.800 174.200 ;
        RECT 35.000 171.800 35.400 172.200 ;
        RECT 34.200 167.800 34.600 168.200 ;
        RECT 34.200 167.200 34.500 167.800 ;
        RECT 30.200 166.800 30.600 167.200 ;
        RECT 31.800 166.800 32.200 167.200 ;
        RECT 34.200 166.800 34.600 167.200 ;
        RECT 30.200 166.200 30.500 166.800 ;
        RECT 35.000 166.200 35.300 171.800 ;
        RECT 36.600 171.200 36.900 173.800 ;
        RECT 37.400 173.200 37.700 173.800 ;
        RECT 37.400 172.800 37.800 173.200 ;
        RECT 36.600 170.800 37.000 171.200 ;
        RECT 36.600 167.800 37.000 168.200 ;
        RECT 36.600 167.200 36.900 167.800 ;
        RECT 36.600 166.800 37.000 167.200 ;
        RECT 30.200 165.800 30.600 166.200 ;
        RECT 31.800 165.800 32.200 166.200 ;
        RECT 33.400 165.800 33.800 166.200 ;
        RECT 35.000 165.800 35.400 166.200 ;
        RECT 35.800 165.800 36.200 166.200 ;
        RECT 37.400 165.800 37.800 166.200 ;
        RECT 38.200 166.100 38.500 175.800 ;
        RECT 40.600 175.200 40.900 175.800 ;
        RECT 39.000 175.100 39.400 175.200 ;
        RECT 39.800 175.100 40.200 175.200 ;
        RECT 39.000 174.800 40.200 175.100 ;
        RECT 40.600 174.800 41.000 175.200 ;
        RECT 43.000 174.200 43.300 177.800 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 52.600 175.200 52.900 176.800 ;
        RECT 53.400 175.200 53.700 190.800 ;
        RECT 59.000 189.200 59.300 211.800 ;
        RECT 59.800 206.200 60.100 222.800 ;
        RECT 61.400 216.200 61.700 234.800 ;
        RECT 62.200 233.800 62.600 234.200 ;
        RECT 64.600 234.100 65.000 234.200 ;
        RECT 65.400 234.100 65.800 234.200 ;
        RECT 64.600 233.800 65.800 234.100 ;
        RECT 67.000 233.800 67.400 234.200 ;
        RECT 62.200 224.200 62.500 233.800 ;
        RECT 67.000 232.200 67.300 233.800 ;
        RECT 67.800 233.100 68.200 235.900 ;
        RECT 68.600 233.800 69.000 234.200 ;
        RECT 68.600 233.200 68.900 233.800 ;
        RECT 68.600 232.800 69.000 233.200 ;
        RECT 67.000 231.800 67.400 232.200 ;
        RECT 69.400 232.100 69.800 237.900 ;
        RECT 71.000 234.800 71.400 235.200 ;
        RECT 71.000 234.200 71.300 234.800 ;
        RECT 71.000 233.800 71.400 234.200 ;
        RECT 72.600 231.800 73.000 232.200 ;
        RECT 74.200 232.100 74.600 237.900 ;
        RECT 77.400 233.100 77.800 235.900 ;
        RECT 75.800 232.100 76.200 232.200 ;
        RECT 76.600 232.100 77.000 232.200 ;
        RECT 79.000 232.100 79.400 237.900 ;
        RECT 80.600 235.100 81.000 235.200 ;
        RECT 81.400 235.100 81.800 235.200 ;
        RECT 80.600 234.800 81.800 235.100 ;
        RECT 83.000 234.800 83.400 235.200 ;
        RECT 79.800 232.800 80.200 233.200 ;
        RECT 75.800 231.800 77.000 232.100 ;
        RECT 63.000 229.100 63.400 229.200 ;
        RECT 63.800 229.100 64.200 229.200 ;
        RECT 63.000 228.800 64.200 229.100 ;
        RECT 68.600 228.800 69.000 229.200 ;
        RECT 68.600 227.200 68.900 228.800 ;
        RECT 63.800 226.800 64.200 227.200 ;
        RECT 65.400 227.100 65.800 227.200 ;
        RECT 66.200 227.100 66.600 227.200 ;
        RECT 65.400 226.800 66.600 227.100 ;
        RECT 68.600 226.800 69.000 227.200 ;
        RECT 63.800 224.200 64.100 226.800 ;
        RECT 72.600 226.200 72.900 231.800 ;
        RECT 75.000 229.800 75.400 230.200 ;
        RECT 75.000 228.200 75.300 229.800 ;
        RECT 75.000 227.800 75.400 228.200 ;
        RECT 64.600 225.800 65.000 226.200 ;
        RECT 72.600 225.800 73.000 226.200 ;
        RECT 73.400 225.800 73.800 226.200 ;
        RECT 64.600 225.200 64.900 225.800 ;
        RECT 73.400 225.200 73.700 225.800 ;
        RECT 64.600 224.800 65.000 225.200 ;
        RECT 67.000 224.800 67.400 225.200 ;
        RECT 73.400 224.800 73.800 225.200 ;
        RECT 62.200 223.800 62.600 224.200 ;
        RECT 63.800 223.800 64.200 224.200 ;
        RECT 67.000 216.200 67.300 224.800 ;
        RECT 71.800 221.800 72.200 222.200 ;
        RECT 73.400 222.100 73.800 222.200 ;
        RECT 74.200 222.100 74.600 222.200 ;
        RECT 73.400 221.800 74.600 222.100 ;
        RECT 70.200 216.800 70.600 217.200 ;
        RECT 61.400 215.800 61.800 216.200 ;
        RECT 66.200 215.800 66.600 216.200 ;
        RECT 67.000 215.800 67.400 216.200 ;
        RECT 67.800 216.100 68.200 216.200 ;
        RECT 68.600 216.100 69.000 216.200 ;
        RECT 67.800 215.800 69.000 216.100 ;
        RECT 61.400 215.200 61.700 215.800 ;
        RECT 66.200 215.200 66.500 215.800 ;
        RECT 61.400 214.800 61.800 215.200 ;
        RECT 63.800 214.800 64.200 215.200 ;
        RECT 66.200 214.800 66.600 215.200 ;
        RECT 68.600 214.800 69.000 215.200 ;
        RECT 63.800 214.200 64.100 214.800 ;
        RECT 61.400 214.100 61.800 214.200 ;
        RECT 62.200 214.100 62.600 214.200 ;
        RECT 61.400 213.800 62.600 214.100 ;
        RECT 63.800 213.800 64.200 214.200 ;
        RECT 64.600 213.800 65.000 214.200 ;
        RECT 64.600 213.200 64.900 213.800 ;
        RECT 64.600 212.800 65.000 213.200 ;
        RECT 59.800 205.800 60.200 206.200 ;
        RECT 60.600 203.100 61.000 208.900 ;
        RECT 63.800 207.800 64.200 208.200 ;
        RECT 63.800 207.200 64.100 207.800 ;
        RECT 63.800 206.800 64.200 207.200 ;
        RECT 65.400 206.800 65.800 207.200 ;
        RECT 65.400 206.200 65.700 206.800 ;
        RECT 65.400 205.800 65.800 206.200 ;
        RECT 59.800 192.100 60.200 197.900 ;
        RECT 65.400 197.800 65.800 198.200 ;
        RECT 61.400 193.100 61.800 195.900 ;
        RECT 62.200 194.800 62.600 195.200 ;
        RECT 63.800 195.100 64.200 195.200 ;
        RECT 64.600 195.100 65.000 195.200 ;
        RECT 63.800 194.800 65.000 195.100 ;
        RECT 62.200 194.200 62.500 194.800 ;
        RECT 62.200 193.800 62.600 194.200 ;
        RECT 63.000 193.800 63.400 194.200 ;
        RECT 65.400 194.100 65.700 197.800 ;
        RECT 64.600 193.800 65.700 194.100 ;
        RECT 63.000 193.200 63.300 193.800 ;
        RECT 63.000 192.800 63.400 193.200 ;
        RECT 59.000 188.800 59.400 189.200 ;
        RECT 61.400 188.800 61.800 189.200 ;
        RECT 55.000 186.800 55.400 187.200 ;
        RECT 55.800 186.800 56.200 187.200 ;
        RECT 60.600 186.800 61.000 187.200 ;
        RECT 55.000 185.200 55.300 186.800 ;
        RECT 55.800 186.200 56.100 186.800 ;
        RECT 60.600 186.200 60.900 186.800 ;
        RECT 61.400 186.200 61.700 188.800 ;
        RECT 64.600 186.200 64.900 193.800 ;
        RECT 65.400 192.800 65.800 193.200 ;
        RECT 65.400 192.200 65.700 192.800 ;
        RECT 66.200 192.200 66.500 214.800 ;
        RECT 68.600 214.200 68.900 214.800 ;
        RECT 70.200 214.200 70.500 216.800 ;
        RECT 68.600 213.800 69.000 214.200 ;
        RECT 70.200 213.800 70.600 214.200 ;
        RECT 67.800 206.100 68.200 206.200 ;
        RECT 68.600 206.100 69.000 206.200 ;
        RECT 67.800 205.800 69.000 206.100 ;
        RECT 69.400 205.800 69.800 206.200 ;
        RECT 69.400 203.200 69.700 205.800 ;
        RECT 69.400 202.800 69.800 203.200 ;
        RECT 67.000 199.800 67.400 200.200 ;
        RECT 67.000 195.200 67.300 199.800 ;
        RECT 70.200 198.200 70.500 213.800 ;
        RECT 71.000 207.800 71.400 208.200 ;
        RECT 71.000 206.200 71.300 207.800 ;
        RECT 71.000 205.800 71.400 206.200 ;
        RECT 71.800 198.200 72.100 221.800 ;
        RECT 74.200 220.800 74.600 221.200 ;
        RECT 73.400 212.100 73.800 217.900 ;
        RECT 74.200 217.200 74.500 220.800 ;
        RECT 74.200 216.800 74.600 217.200 ;
        RECT 73.400 207.800 73.800 208.200 ;
        RECT 73.400 206.200 73.700 207.800 ;
        RECT 74.200 206.200 74.500 216.800 ;
        RECT 75.000 215.200 75.300 227.800 ;
        RECT 76.600 223.100 77.000 228.900 ;
        RECT 79.800 227.200 80.100 232.800 ;
        RECT 83.000 231.200 83.300 234.800 ;
        RECT 83.800 232.100 84.200 237.900 ;
        RECT 92.600 235.800 93.000 236.200 ;
        RECT 92.600 235.200 92.900 235.800 ;
        RECT 88.600 234.800 89.000 235.200 ;
        RECT 91.800 234.800 92.200 235.200 ;
        RECT 92.600 234.800 93.000 235.200 ;
        RECT 88.600 234.200 88.900 234.800 ;
        RECT 88.600 233.800 89.000 234.200 ;
        RECT 91.800 234.100 92.100 234.800 ;
        RECT 91.800 233.800 92.900 234.100 ;
        RECT 87.000 232.800 87.400 233.200 ;
        RECT 83.000 230.800 83.400 231.200 ;
        RECT 87.000 230.200 87.300 232.800 ;
        RECT 87.000 229.800 87.400 230.200 ;
        RECT 79.800 226.800 80.200 227.200 ;
        RECT 80.600 226.800 81.000 227.200 ;
        RECT 77.400 215.800 77.800 216.200 ;
        RECT 75.000 214.800 75.400 215.200 ;
        RECT 75.800 215.100 76.200 215.200 ;
        RECT 76.600 215.100 77.000 215.200 ;
        RECT 75.800 214.800 77.000 215.100 ;
        RECT 75.000 209.800 75.400 210.200 ;
        RECT 75.000 208.200 75.300 209.800 ;
        RECT 75.000 207.800 75.400 208.200 ;
        RECT 75.000 207.200 75.300 207.800 ;
        RECT 75.000 206.800 75.400 207.200 ;
        RECT 76.600 206.800 77.000 207.200 ;
        RECT 76.600 206.200 76.900 206.800 ;
        RECT 73.400 205.800 73.800 206.200 ;
        RECT 74.200 206.100 74.600 206.200 ;
        RECT 74.200 205.800 75.300 206.100 ;
        RECT 76.600 205.800 77.000 206.200 ;
        RECT 72.600 201.800 73.000 202.200 ;
        RECT 70.200 197.800 70.600 198.200 ;
        RECT 71.800 197.800 72.200 198.200 ;
        RECT 69.400 196.800 69.800 197.200 ;
        RECT 67.800 195.800 68.200 196.200 ;
        RECT 68.600 195.800 69.000 196.200 ;
        RECT 67.000 194.800 67.400 195.200 ;
        RECT 67.000 193.200 67.300 194.800 ;
        RECT 67.000 192.800 67.400 193.200 ;
        RECT 65.400 191.800 65.800 192.200 ;
        RECT 66.200 191.800 66.600 192.200 ;
        RECT 67.800 192.100 68.100 195.800 ;
        RECT 68.600 195.200 68.900 195.800 ;
        RECT 69.400 195.200 69.700 196.800 ;
        RECT 68.600 194.800 69.000 195.200 ;
        RECT 69.400 194.800 69.800 195.200 ;
        RECT 67.000 191.800 68.100 192.100 ;
        RECT 65.400 190.800 65.800 191.200 ;
        RECT 65.400 187.200 65.700 190.800 ;
        RECT 67.000 189.200 67.300 191.800 ;
        RECT 67.000 188.800 67.400 189.200 ;
        RECT 69.400 188.200 69.700 194.800 ;
        RECT 70.200 193.800 70.600 194.200 ;
        RECT 67.000 187.800 67.400 188.200 ;
        RECT 69.400 187.800 69.800 188.200 ;
        RECT 65.400 186.800 65.800 187.200 ;
        RECT 55.800 185.800 56.200 186.200 ;
        RECT 56.600 185.800 57.000 186.200 ;
        RECT 59.000 186.100 59.400 186.200 ;
        RECT 59.800 186.100 60.200 186.200 ;
        RECT 59.000 185.800 60.200 186.100 ;
        RECT 60.600 185.800 61.000 186.200 ;
        RECT 61.400 185.800 61.800 186.200 ;
        RECT 63.000 186.100 63.400 186.200 ;
        RECT 63.800 186.100 64.200 186.200 ;
        RECT 63.000 185.800 64.200 186.100 ;
        RECT 64.600 185.800 65.000 186.200 ;
        RECT 56.600 185.200 56.900 185.800 ;
        RECT 67.000 185.200 67.300 187.800 ;
        RECT 70.200 186.200 70.500 193.800 ;
        RECT 71.000 191.800 71.400 192.200 ;
        RECT 71.000 191.200 71.300 191.800 ;
        RECT 71.000 190.800 71.400 191.200 ;
        RECT 71.800 186.800 72.200 187.200 ;
        RECT 71.800 186.200 72.100 186.800 ;
        RECT 67.800 185.800 68.200 186.200 ;
        RECT 68.600 185.800 69.000 186.200 ;
        RECT 70.200 185.800 70.600 186.200 ;
        RECT 71.800 185.800 72.200 186.200 ;
        RECT 55.000 184.800 55.400 185.200 ;
        RECT 56.600 184.800 57.000 185.200 ;
        RECT 66.200 185.100 66.600 185.200 ;
        RECT 67.000 185.100 67.400 185.200 ;
        RECT 66.200 184.800 67.400 185.100 ;
        RECT 61.400 183.800 61.800 184.200 ;
        RECT 58.200 181.800 58.600 182.200 ;
        RECT 58.200 178.200 58.500 181.800 ;
        RECT 58.200 177.800 58.600 178.200 ;
        RECT 55.800 176.800 56.200 177.200 ;
        RECT 55.800 175.200 56.100 176.800 ;
        RECT 43.800 175.100 44.200 175.200 ;
        RECT 44.600 175.100 45.000 175.200 ;
        RECT 43.800 174.800 45.000 175.100 ;
        RECT 47.000 174.800 47.400 175.200 ;
        RECT 47.800 175.100 48.200 175.200 ;
        RECT 48.600 175.100 49.000 175.200 ;
        RECT 47.800 174.800 49.000 175.100 ;
        RECT 49.400 174.800 49.800 175.200 ;
        RECT 52.600 174.800 53.000 175.200 ;
        RECT 53.400 174.800 53.800 175.200 ;
        RECT 54.200 174.800 54.600 175.200 ;
        RECT 55.800 174.800 56.200 175.200 ;
        RECT 56.600 175.100 57.000 175.200 ;
        RECT 57.400 175.100 57.800 175.200 ;
        RECT 56.600 174.800 57.800 175.100 ;
        RECT 47.000 174.200 47.300 174.800 ;
        RECT 39.800 174.100 40.200 174.200 ;
        RECT 40.600 174.100 41.000 174.200 ;
        RECT 39.800 173.800 41.000 174.100 ;
        RECT 41.400 173.800 41.800 174.200 ;
        RECT 43.000 173.800 43.400 174.200 ;
        RECT 47.000 173.800 47.400 174.200 ;
        RECT 41.400 173.200 41.700 173.800 ;
        RECT 41.400 172.800 41.800 173.200 ;
        RECT 39.000 171.800 39.400 172.200 ;
        RECT 42.200 172.100 42.600 172.200 ;
        RECT 43.000 172.100 43.400 172.200 ;
        RECT 42.200 171.800 43.400 172.100 ;
        RECT 45.400 171.800 45.800 172.200 ;
        RECT 39.000 168.200 39.300 171.800 ;
        RECT 45.400 171.200 45.700 171.800 ;
        RECT 40.600 170.800 41.000 171.200 ;
        RECT 45.400 170.800 45.800 171.200 ;
        RECT 40.600 169.200 40.900 170.800 ;
        RECT 40.600 168.800 41.000 169.200 ;
        RECT 39.000 167.800 39.400 168.200 ;
        RECT 39.000 167.100 39.400 167.200 ;
        RECT 39.800 167.100 40.200 167.200 ;
        RECT 39.000 166.800 40.200 167.100 ;
        RECT 39.000 166.100 39.400 166.200 ;
        RECT 38.200 165.800 39.400 166.100 ;
        RECT 39.800 165.800 40.200 166.200 ;
        RECT 27.800 165.100 28.200 165.200 ;
        RECT 28.600 165.100 29.000 165.200 ;
        RECT 27.800 164.800 29.000 165.100 ;
        RECT 29.400 153.100 29.800 155.900 ;
        RECT 30.200 153.800 30.600 154.200 ;
        RECT 28.600 152.100 29.000 152.200 ;
        RECT 29.400 152.100 29.800 152.200 ;
        RECT 28.600 151.800 29.800 152.100 ;
        RECT 30.200 147.200 30.500 153.800 ;
        RECT 31.000 152.100 31.400 157.900 ;
        RECT 31.800 154.200 32.100 165.800 ;
        RECT 33.400 165.200 33.700 165.800 ;
        RECT 35.800 165.200 36.100 165.800 ;
        RECT 37.400 165.200 37.700 165.800 ;
        RECT 33.400 165.100 33.800 165.200 ;
        RECT 34.200 165.100 34.600 165.200 ;
        RECT 33.400 164.800 34.600 165.100 ;
        RECT 35.800 164.800 36.200 165.200 ;
        RECT 37.400 164.800 37.800 165.200 ;
        RECT 32.600 154.800 33.000 155.200 ;
        RECT 31.800 153.800 32.200 154.200 ;
        RECT 32.600 149.200 32.900 154.800 ;
        RECT 35.800 152.100 36.200 157.900 ;
        RECT 38.200 156.200 38.500 165.800 ;
        RECT 39.000 165.100 39.400 165.200 ;
        RECT 39.800 165.100 40.100 165.800 ;
        RECT 39.000 164.800 40.100 165.100 ;
        RECT 43.000 163.100 43.400 168.900 ;
        RECT 45.400 166.100 45.800 166.200 ;
        RECT 46.200 166.100 46.600 166.200 ;
        RECT 45.400 165.800 46.600 166.100 ;
        RECT 45.400 156.800 45.800 157.200 ;
        RECT 45.400 156.200 45.700 156.800 ;
        RECT 38.200 155.800 38.600 156.200 ;
        RECT 45.400 155.800 45.800 156.200 ;
        RECT 47.000 155.200 47.300 173.800 ;
        RECT 49.400 173.200 49.700 174.800 ;
        RECT 54.200 174.200 54.500 174.800 ;
        RECT 54.200 173.800 54.600 174.200 ;
        RECT 49.400 172.800 49.800 173.200 ;
        RECT 49.400 172.200 49.700 172.800 ;
        RECT 48.600 171.800 49.000 172.200 ;
        RECT 49.400 171.800 49.800 172.200 ;
        RECT 55.000 171.800 55.400 172.200 ;
        RECT 58.200 172.100 58.600 172.200 ;
        RECT 59.000 172.100 59.400 172.200 ;
        RECT 58.200 171.800 59.400 172.100 ;
        RECT 48.600 169.200 48.900 171.800 ;
        RECT 53.400 170.800 53.800 171.200 ;
        RECT 47.800 163.100 48.200 168.900 ;
        RECT 48.600 168.800 49.000 169.200 ;
        RECT 50.200 168.800 50.600 169.200 ;
        RECT 50.200 168.200 50.500 168.800 ;
        RECT 48.600 166.800 49.000 167.200 ;
        RECT 48.600 159.200 48.900 166.800 ;
        RECT 49.400 165.100 49.800 167.900 ;
        RECT 50.200 167.800 50.600 168.200 ;
        RECT 51.800 167.100 52.200 167.200 ;
        RECT 52.600 167.100 53.000 167.200 ;
        RECT 51.800 166.800 53.000 167.100 ;
        RECT 53.400 166.200 53.700 170.800 ;
        RECT 55.000 169.200 55.300 171.800 ;
        RECT 60.600 169.800 61.000 170.200 ;
        RECT 55.000 168.800 55.400 169.200 ;
        RECT 51.000 166.100 51.400 166.200 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 51.000 165.800 52.200 166.100 ;
        RECT 53.400 165.800 53.800 166.200 ;
        RECT 57.400 163.100 57.800 168.900 ;
        RECT 58.200 165.800 58.600 166.200 ;
        RECT 59.000 166.100 59.400 166.200 ;
        RECT 59.800 166.100 60.200 166.200 ;
        RECT 59.000 165.800 60.200 166.100 ;
        RECT 58.200 162.200 58.500 165.800 ;
        RECT 58.200 161.800 58.600 162.200 ;
        RECT 48.600 158.800 49.000 159.200 ;
        RECT 58.200 158.200 58.500 161.800 ;
        RECT 59.000 158.800 59.400 159.200 ;
        RECT 56.600 157.800 57.000 158.200 ;
        RECT 48.600 155.800 49.000 156.200 ;
        RECT 48.600 155.200 48.900 155.800 ;
        RECT 40.600 155.100 41.000 155.200 ;
        RECT 41.400 155.100 41.800 155.200 ;
        RECT 40.600 154.800 41.800 155.100 ;
        RECT 43.000 154.800 43.400 155.200 ;
        RECT 47.000 154.800 47.400 155.200 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 48.600 154.800 49.000 155.200 ;
        RECT 53.400 154.800 53.800 155.200 ;
        RECT 43.000 154.200 43.300 154.800 ;
        RECT 47.800 154.200 48.100 154.800 ;
        RECT 43.000 153.800 43.400 154.200 ;
        RECT 47.800 153.800 48.200 154.200 ;
        RECT 51.000 154.100 51.400 154.200 ;
        RECT 51.800 154.100 52.200 154.200 ;
        RECT 51.000 153.800 52.200 154.100 ;
        RECT 39.000 152.800 39.400 153.200 ;
        RECT 42.200 152.800 42.600 153.200 ;
        RECT 39.000 152.200 39.300 152.800 ;
        RECT 42.200 152.200 42.500 152.800 ;
        RECT 38.200 151.800 38.600 152.200 ;
        RECT 39.000 151.800 39.400 152.200 ;
        RECT 42.200 151.800 42.600 152.200 ;
        RECT 32.600 148.800 33.000 149.200 ;
        RECT 36.600 147.800 37.000 148.200 ;
        RECT 30.200 146.800 30.600 147.200 ;
        RECT 27.000 141.800 27.400 142.200 ;
        RECT 22.200 140.800 22.600 141.200 ;
        RECT 27.800 136.800 28.200 137.200 ;
        RECT 29.400 136.800 29.800 137.200 ;
        RECT 27.800 135.200 28.100 136.800 ;
        RECT 29.400 135.200 29.700 136.800 ;
        RECT 15.000 134.800 15.400 135.200 ;
        RECT 15.800 134.800 16.200 135.200 ;
        RECT 19.000 134.800 19.400 135.200 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 20.600 134.800 21.000 135.200 ;
        RECT 21.400 134.800 21.800 135.200 ;
        RECT 23.000 135.100 23.400 135.200 ;
        RECT 23.800 135.100 24.200 135.200 ;
        RECT 23.000 134.800 24.200 135.100 ;
        RECT 24.600 135.100 25.000 135.200 ;
        RECT 25.400 135.100 25.800 135.200 ;
        RECT 24.600 134.800 25.800 135.100 ;
        RECT 27.800 134.800 28.200 135.200 ;
        RECT 29.400 134.800 29.800 135.200 ;
        RECT 12.600 133.800 13.000 134.200 ;
        RECT 14.200 133.800 14.600 134.200 ;
        RECT 7.000 126.800 7.400 127.200 ;
        RECT 7.000 115.200 7.300 126.800 ;
        RECT 7.800 125.100 8.200 127.900 ;
        RECT 9.400 123.100 9.800 128.900 ;
        RECT 11.000 126.100 11.400 126.200 ;
        RECT 11.800 126.100 12.200 126.200 ;
        RECT 11.000 125.800 12.200 126.100 ;
        RECT 14.200 123.100 14.600 128.900 ;
        RECT 15.000 128.200 15.300 134.800 ;
        RECT 18.200 131.800 18.600 132.200 ;
        RECT 16.600 129.100 17.000 129.200 ;
        RECT 17.400 129.100 17.800 129.200 ;
        RECT 16.600 128.800 17.800 129.100 ;
        RECT 15.000 127.800 15.400 128.200 ;
        RECT 17.400 127.800 17.800 128.200 ;
        RECT 7.000 114.800 7.400 115.200 ;
        RECT 3.000 106.800 3.400 107.200 ;
        RECT 1.400 103.100 1.800 103.200 ;
        RECT 2.200 103.100 2.600 103.200 ;
        RECT 1.400 102.800 2.600 103.100 ;
        RECT 0.600 93.100 1.000 95.900 ;
        RECT 2.200 92.100 2.600 97.900 ;
        RECT 3.000 94.200 3.300 106.800 ;
        RECT 4.600 105.100 5.000 107.900 ;
        RECT 6.200 103.100 6.600 108.900 ;
        RECT 7.000 108.200 7.300 114.800 ;
        RECT 7.800 113.100 8.200 115.900 ;
        RECT 8.600 113.800 9.000 114.200 ;
        RECT 7.000 107.800 7.400 108.200 ;
        RECT 8.600 107.200 8.900 113.800 ;
        RECT 9.400 112.100 9.800 117.900 ;
        RECT 11.800 116.800 12.200 117.200 ;
        RECT 11.800 115.200 12.100 116.800 ;
        RECT 11.800 114.800 12.200 115.200 ;
        RECT 14.200 112.100 14.600 117.900 ;
        RECT 16.600 116.800 17.000 117.200 ;
        RECT 16.600 115.200 16.900 116.800 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 17.400 114.200 17.700 127.800 ;
        RECT 18.200 127.200 18.500 131.800 ;
        RECT 19.000 129.200 19.300 134.800 ;
        RECT 19.000 128.800 19.400 129.200 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 19.000 126.800 19.400 127.200 ;
        RECT 19.000 126.200 19.300 126.800 ;
        RECT 19.000 125.800 19.400 126.200 ;
        RECT 19.000 125.100 19.400 125.200 ;
        RECT 19.800 125.100 20.200 125.200 ;
        RECT 19.000 124.800 20.200 125.100 ;
        RECT 20.600 124.100 20.900 134.800 ;
        RECT 30.200 134.100 30.500 146.800 ;
        RECT 36.600 146.200 36.900 147.800 ;
        RECT 38.200 146.200 38.500 151.800 ;
        RECT 39.000 150.200 39.300 151.800 ;
        RECT 39.000 149.800 39.400 150.200 ;
        RECT 39.000 149.100 39.400 149.200 ;
        RECT 39.800 149.100 40.200 149.200 ;
        RECT 39.000 148.800 40.200 149.100 ;
        RECT 41.400 147.100 41.800 147.200 ;
        RECT 42.200 147.100 42.600 147.200 ;
        RECT 41.400 146.800 42.600 147.100 ;
        RECT 31.000 145.800 31.400 146.200 ;
        RECT 31.800 145.800 32.200 146.200 ;
        RECT 36.600 145.800 37.000 146.200 ;
        RECT 37.400 145.800 37.800 146.200 ;
        RECT 38.200 146.100 38.600 146.200 ;
        RECT 39.000 146.100 39.400 146.200 ;
        RECT 38.200 145.800 39.400 146.100 ;
        RECT 40.600 145.800 41.000 146.200 ;
        RECT 31.000 142.200 31.300 145.800 ;
        RECT 31.000 141.800 31.400 142.200 ;
        RECT 31.800 135.200 32.100 145.800 ;
        RECT 35.000 144.800 35.400 145.200 ;
        RECT 35.000 139.200 35.300 144.800 ;
        RECT 37.400 143.200 37.700 145.800 ;
        RECT 40.600 145.200 40.900 145.800 ;
        RECT 40.600 144.800 41.000 145.200 ;
        RECT 37.400 142.800 37.800 143.200 ;
        RECT 35.000 138.800 35.400 139.200 ;
        RECT 33.400 137.100 33.800 137.200 ;
        RECT 34.200 137.100 34.600 137.200 ;
        RECT 33.400 136.800 34.600 137.100 ;
        RECT 31.800 134.800 32.200 135.200 ;
        RECT 32.600 134.800 33.000 135.200 ;
        RECT 31.800 134.200 32.100 134.800 ;
        RECT 31.000 134.100 31.400 134.200 ;
        RECT 30.200 133.800 31.400 134.100 ;
        RECT 31.800 133.800 32.200 134.200 ;
        RECT 22.200 133.100 22.600 133.200 ;
        RECT 23.000 133.100 23.400 133.200 ;
        RECT 22.200 132.800 23.400 133.100 ;
        RECT 30.200 133.100 30.600 133.200 ;
        RECT 31.000 133.100 31.400 133.200 ;
        RECT 30.200 132.800 31.400 133.100 ;
        RECT 26.200 131.800 26.600 132.200 ;
        RECT 21.400 129.800 21.800 130.200 ;
        RECT 21.400 126.200 21.700 129.800 ;
        RECT 24.600 129.100 25.000 129.200 ;
        RECT 25.400 129.100 25.800 129.200 ;
        RECT 24.600 128.800 25.800 129.100 ;
        RECT 26.200 128.200 26.500 131.800 ;
        RECT 32.600 131.200 32.900 134.800 ;
        RECT 37.400 132.100 37.800 137.900 ;
        RECT 40.600 134.800 41.000 135.200 ;
        RECT 38.200 133.800 38.600 134.200 ;
        RECT 32.600 130.800 33.000 131.200 ;
        RECT 22.200 127.800 22.600 128.200 ;
        RECT 26.200 127.800 26.600 128.200 ;
        RECT 22.200 127.200 22.500 127.800 ;
        RECT 22.200 126.800 22.600 127.200 ;
        RECT 23.000 126.800 23.400 127.200 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 23.000 126.200 23.300 126.800 ;
        RECT 27.000 126.200 27.300 126.800 ;
        RECT 21.400 125.800 21.800 126.200 ;
        RECT 23.000 125.800 23.400 126.200 ;
        RECT 26.200 126.100 26.600 126.200 ;
        RECT 25.400 125.800 26.600 126.100 ;
        RECT 27.000 125.800 27.400 126.200 ;
        RECT 21.400 125.200 21.700 125.800 ;
        RECT 21.400 124.800 21.800 125.200 ;
        RECT 19.800 123.800 20.900 124.100 ;
        RECT 18.200 117.100 18.600 117.200 ;
        RECT 19.000 117.100 19.400 117.200 ;
        RECT 18.200 116.800 19.400 117.100 ;
        RECT 18.200 115.800 18.600 116.200 ;
        RECT 18.200 115.200 18.500 115.800 ;
        RECT 18.200 114.800 18.600 115.200 ;
        RECT 17.400 113.800 17.800 114.200 ;
        RECT 19.800 113.200 20.100 123.800 ;
        RECT 25.400 119.200 25.700 125.800 ;
        RECT 27.800 125.100 28.200 127.900 ;
        RECT 29.400 123.100 29.800 128.900 ;
        RECT 30.200 128.800 30.600 129.200 ;
        RECT 30.200 128.200 30.500 128.800 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 31.800 126.100 32.200 126.200 ;
        RECT 32.600 126.100 33.000 126.200 ;
        RECT 31.800 125.800 33.000 126.100 ;
        RECT 32.600 124.800 33.000 125.200 ;
        RECT 25.400 118.800 25.800 119.200 ;
        RECT 20.600 116.100 21.000 116.200 ;
        RECT 21.400 116.100 21.800 116.200 ;
        RECT 20.600 115.800 21.800 116.100 ;
        RECT 22.200 114.800 22.600 115.200 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 23.800 115.100 24.200 115.200 ;
        RECT 24.600 115.100 25.000 115.200 ;
        RECT 23.800 114.800 25.000 115.100 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 27.800 114.800 28.200 115.200 ;
        RECT 22.200 114.200 22.500 114.800 ;
        RECT 22.200 113.800 22.600 114.200 ;
        RECT 23.000 113.200 23.300 114.800 ;
        RECT 27.000 113.200 27.300 114.800 ;
        RECT 27.800 114.200 28.100 114.800 ;
        RECT 27.800 113.800 28.200 114.200 ;
        RECT 28.600 114.100 29.000 114.200 ;
        RECT 29.400 114.100 29.800 114.200 ;
        RECT 28.600 113.800 29.800 114.100 ;
        RECT 18.200 112.800 18.600 113.200 ;
        RECT 19.800 112.800 20.200 113.200 ;
        RECT 23.000 112.800 23.400 113.200 ;
        RECT 27.000 112.800 27.400 113.200 ;
        RECT 28.600 112.800 29.000 113.200 ;
        RECT 30.200 113.100 30.600 113.200 ;
        RECT 31.000 113.100 31.400 113.200 ;
        RECT 30.200 112.800 31.400 113.100 ;
        RECT 13.400 109.100 13.800 109.200 ;
        RECT 14.200 109.100 14.600 109.200 ;
        RECT 8.600 106.800 9.000 107.200 ;
        RECT 7.800 106.100 8.200 106.200 ;
        RECT 8.600 106.100 9.000 106.200 ;
        RECT 7.800 105.800 9.000 106.100 ;
        RECT 11.000 103.100 11.400 108.900 ;
        RECT 13.400 108.800 14.600 109.100 ;
        RECT 15.000 107.800 15.400 108.200 ;
        RECT 17.400 107.800 17.800 108.200 ;
        RECT 15.000 107.200 15.300 107.800 ;
        RECT 15.000 106.800 15.400 107.200 ;
        RECT 17.400 106.200 17.700 107.800 ;
        RECT 14.200 106.100 14.600 106.200 ;
        RECT 15.800 106.100 16.200 106.200 ;
        RECT 16.600 106.100 17.000 106.200 ;
        RECT 14.200 105.800 15.300 106.100 ;
        RECT 15.800 105.800 17.000 106.100 ;
        RECT 17.400 105.800 17.800 106.200 ;
        RECT 11.800 99.800 12.200 100.200 ;
        RECT 14.200 99.800 14.600 100.200 ;
        RECT 5.400 94.800 5.800 95.200 ;
        RECT 6.200 94.800 6.600 95.200 ;
        RECT 5.400 94.200 5.700 94.800 ;
        RECT 3.000 93.800 3.400 94.200 ;
        RECT 5.400 93.800 5.800 94.200 ;
        RECT 0.600 85.100 1.000 87.900 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 0.600 73.100 1.000 75.900 ;
        RECT 1.400 74.200 1.700 86.800 ;
        RECT 2.200 83.100 2.600 88.900 ;
        RECT 3.800 86.100 4.200 86.200 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 3.800 85.800 5.000 86.100 ;
        RECT 1.400 73.800 1.800 74.200 ;
        RECT 1.400 69.200 1.700 73.800 ;
        RECT 2.200 72.100 2.600 77.900 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 3.800 74.800 5.000 75.100 ;
        RECT 1.400 68.800 1.800 69.200 ;
        RECT 0.600 66.800 1.000 67.200 ;
        RECT 0.600 66.200 0.900 66.800 ;
        RECT 0.600 65.800 1.000 66.200 ;
        RECT 0.600 54.200 0.900 65.800 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 0.600 45.100 1.000 47.900 ;
        RECT 2.200 43.100 2.600 48.900 ;
        RECT 3.800 46.100 4.200 46.200 ;
        RECT 4.600 46.100 5.000 46.200 ;
        RECT 3.800 45.800 5.000 46.100 ;
        RECT 5.400 45.800 5.800 46.200 ;
        RECT 0.600 38.800 1.000 39.200 ;
        RECT 0.600 35.200 0.900 38.800 ;
        RECT 1.400 36.800 1.800 37.200 ;
        RECT 3.800 36.800 4.200 37.200 ;
        RECT 0.600 34.800 1.000 35.200 ;
        RECT 1.400 34.200 1.700 36.800 ;
        RECT 3.800 35.200 4.100 36.800 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 1.400 33.800 1.800 34.200 ;
        RECT 3.000 33.800 3.400 34.200 ;
        RECT 5.400 34.100 5.700 45.800 ;
        RECT 6.200 35.200 6.500 94.800 ;
        RECT 7.000 92.100 7.400 97.900 ;
        RECT 9.400 97.100 9.800 97.200 ;
        RECT 10.200 97.100 10.600 97.200 ;
        RECT 9.400 96.800 10.600 97.100 ;
        RECT 11.800 96.200 12.100 99.800 ;
        RECT 11.800 95.800 12.200 96.200 ;
        RECT 14.200 95.200 14.500 99.800 ;
        RECT 14.200 94.800 14.600 95.200 ;
        RECT 15.000 94.200 15.300 105.800 ;
        RECT 18.200 99.200 18.500 112.800 ;
        RECT 24.600 111.800 25.000 112.200 ;
        RECT 19.000 108.800 19.400 109.200 ;
        RECT 19.000 108.200 19.300 108.800 ;
        RECT 19.000 107.800 19.400 108.200 ;
        RECT 19.800 105.100 20.200 107.900 ;
        RECT 20.600 106.800 21.000 107.200 ;
        RECT 20.600 106.200 20.900 106.800 ;
        RECT 20.600 105.800 21.000 106.200 ;
        RECT 21.400 103.100 21.800 108.900 ;
        RECT 24.600 106.200 24.900 111.800 ;
        RECT 28.600 109.200 28.900 112.800 ;
        RECT 29.400 111.800 29.800 112.200 ;
        RECT 29.400 111.200 29.700 111.800 ;
        RECT 29.400 110.800 29.800 111.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 26.200 103.100 26.600 108.900 ;
        RECT 28.600 108.800 29.000 109.200 ;
        RECT 30.200 108.800 30.600 109.200 ;
        RECT 30.200 106.200 30.500 108.800 ;
        RECT 29.400 105.800 29.800 106.200 ;
        RECT 30.200 105.800 30.600 106.200 ;
        RECT 29.400 99.200 29.700 105.800 ;
        RECT 18.200 98.800 18.600 99.200 ;
        RECT 29.400 98.800 29.800 99.200 ;
        RECT 16.600 96.800 17.000 97.200 ;
        RECT 15.800 95.800 16.200 96.200 ;
        RECT 15.800 95.200 16.100 95.800 ;
        RECT 16.600 95.200 16.900 96.800 ;
        RECT 22.200 95.800 22.600 96.200 ;
        RECT 22.200 95.200 22.500 95.800 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 11.800 94.100 12.200 94.200 ;
        RECT 12.600 94.100 13.000 94.200 ;
        RECT 11.800 93.800 13.000 94.100 ;
        RECT 15.000 94.100 15.400 94.200 ;
        RECT 15.800 94.100 16.200 94.200 ;
        RECT 15.000 93.800 16.200 94.100 ;
        RECT 19.800 93.800 20.200 94.200 ;
        RECT 10.200 91.800 10.600 92.200 ;
        RECT 7.000 83.100 7.400 88.900 ;
        RECT 10.200 88.200 10.500 91.800 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 11.800 86.800 12.200 87.200 ;
        RECT 11.800 86.200 12.100 86.800 ;
        RECT 15.000 86.200 15.300 93.800 ;
        RECT 19.800 89.200 20.100 93.800 ;
        RECT 23.000 93.100 23.400 95.900 ;
        RECT 23.800 93.800 24.200 94.200 ;
        RECT 23.800 93.200 24.100 93.800 ;
        RECT 23.800 92.800 24.200 93.200 ;
        RECT 21.400 91.800 21.800 92.200 ;
        RECT 24.600 92.100 25.000 97.900 ;
        RECT 26.200 95.800 26.600 96.200 ;
        RECT 26.200 95.200 26.500 95.800 ;
        RECT 26.200 94.800 26.600 95.200 ;
        RECT 27.800 94.800 28.200 95.200 ;
        RECT 16.600 89.100 17.000 89.200 ;
        RECT 17.400 89.100 17.800 89.200 ;
        RECT 16.600 88.800 17.800 89.100 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 15.000 85.800 15.400 86.200 ;
        RECT 15.800 86.100 16.200 86.200 ;
        RECT 16.600 86.100 17.000 86.200 ;
        RECT 15.800 85.800 17.000 86.100 ;
        RECT 19.000 83.100 19.400 88.900 ;
        RECT 19.800 88.800 20.200 89.200 ;
        RECT 21.400 85.200 21.700 91.800 ;
        RECT 22.200 86.800 22.600 87.200 ;
        RECT 22.200 86.200 22.500 86.800 ;
        RECT 22.200 85.800 22.600 86.200 ;
        RECT 21.400 84.800 21.800 85.200 ;
        RECT 23.800 83.100 24.200 88.900 ;
        RECT 24.600 86.800 25.000 87.200 ;
        RECT 24.600 81.200 24.900 86.800 ;
        RECT 25.400 85.100 25.800 87.900 ;
        RECT 26.200 87.100 26.600 87.200 ;
        RECT 27.000 87.100 27.400 87.200 ;
        RECT 26.200 86.800 27.400 87.100 ;
        RECT 27.800 86.200 28.100 94.800 ;
        RECT 28.600 93.800 29.000 94.200 ;
        RECT 28.600 87.200 28.900 93.800 ;
        RECT 29.400 92.100 29.800 97.900 ;
        RECT 32.600 97.200 32.900 124.800 ;
        RECT 34.200 123.100 34.600 128.900 ;
        RECT 36.600 128.800 37.000 129.200 ;
        RECT 36.600 128.200 36.900 128.800 ;
        RECT 36.600 127.800 37.000 128.200 ;
        RECT 38.200 128.100 38.500 133.800 ;
        RECT 40.600 133.200 40.900 134.800 ;
        RECT 40.600 132.800 41.000 133.200 ;
        RECT 41.400 132.800 41.800 133.200 ;
        RECT 41.400 131.200 41.700 132.800 ;
        RECT 42.200 132.100 42.600 137.900 ;
        RECT 43.000 136.200 43.300 153.800 ;
        RECT 53.400 153.200 53.700 154.800 ;
        RECT 53.400 152.800 53.800 153.200 ;
        RECT 55.800 153.100 56.200 155.900 ;
        RECT 56.600 154.200 56.900 157.800 ;
        RECT 56.600 153.800 57.000 154.200 ;
        RECT 57.400 152.100 57.800 157.900 ;
        RECT 58.200 157.800 58.600 158.200 ;
        RECT 58.200 154.700 58.600 155.100 ;
        RECT 58.200 154.200 58.500 154.700 ;
        RECT 58.200 153.800 58.600 154.200 ;
        RECT 45.400 150.800 45.800 151.200 ;
        RECT 43.000 135.800 43.400 136.200 ;
        RECT 41.400 130.800 41.800 131.200 ;
        RECT 37.400 127.800 38.500 128.100 ;
        RECT 42.200 127.800 42.600 128.200 ;
        RECT 37.400 127.200 37.700 127.800 ;
        RECT 42.200 127.200 42.500 127.800 ;
        RECT 37.400 126.800 37.800 127.200 ;
        RECT 38.200 126.800 38.600 127.200 ;
        RECT 40.600 126.800 41.000 127.200 ;
        RECT 42.200 126.800 42.600 127.200 ;
        RECT 35.800 116.800 36.200 117.200 ;
        RECT 35.800 115.200 36.100 116.800 ;
        RECT 37.400 116.100 37.700 126.800 ;
        RECT 38.200 126.200 38.500 126.800 ;
        RECT 38.200 125.800 38.600 126.200 ;
        RECT 39.000 126.100 39.400 126.200 ;
        RECT 39.800 126.100 40.200 126.200 ;
        RECT 39.000 125.800 40.200 126.100 ;
        RECT 40.600 125.200 40.900 126.800 ;
        RECT 42.200 125.800 42.600 126.200 ;
        RECT 40.600 124.800 41.000 125.200 ;
        RECT 37.400 115.800 38.500 116.100 ;
        RECT 33.400 114.800 33.800 115.200 ;
        RECT 34.200 114.800 34.600 115.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 36.600 114.800 37.000 115.200 ;
        RECT 37.400 114.800 37.800 115.200 ;
        RECT 33.400 114.200 33.700 114.800 ;
        RECT 34.200 114.200 34.500 114.800 ;
        RECT 33.400 113.800 33.800 114.200 ;
        RECT 34.200 113.800 34.600 114.200 ;
        RECT 33.400 111.200 33.700 113.800 ;
        RECT 36.600 113.200 36.900 114.800 ;
        RECT 37.400 114.200 37.700 114.800 ;
        RECT 37.400 113.800 37.800 114.200 ;
        RECT 36.600 112.800 37.000 113.200 ;
        RECT 33.400 110.800 33.800 111.200 ;
        RECT 34.200 108.800 34.600 109.200 ;
        RECT 34.200 108.200 34.500 108.800 ;
        RECT 34.200 107.800 34.600 108.200 ;
        RECT 33.400 106.800 33.800 107.200 ;
        RECT 33.400 106.200 33.700 106.800 ;
        RECT 34.200 106.200 34.500 107.800 ;
        RECT 33.400 105.800 33.800 106.200 ;
        RECT 34.200 105.800 34.600 106.200 ;
        RECT 37.400 105.800 37.800 106.200 ;
        RECT 37.400 105.200 37.700 105.800 ;
        RECT 37.400 104.800 37.800 105.200 ;
        RECT 34.200 97.800 34.600 98.200 ;
        RECT 36.600 97.800 37.000 98.200 ;
        RECT 32.600 96.800 33.000 97.200 ;
        RECT 32.600 94.200 32.900 96.800 ;
        RECT 34.200 96.200 34.500 97.800 ;
        RECT 34.200 95.800 34.600 96.200 ;
        RECT 35.000 95.800 35.400 96.200 ;
        RECT 35.000 94.200 35.300 95.800 ;
        RECT 36.600 95.200 36.900 97.800 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 38.200 94.200 38.500 115.800 ;
        RECT 40.600 114.800 41.000 115.200 ;
        RECT 40.600 114.200 40.900 114.800 ;
        RECT 39.000 113.800 39.400 114.200 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 39.000 106.200 39.300 113.800 ;
        RECT 39.800 111.800 40.200 112.200 ;
        RECT 39.800 106.200 40.100 111.800 ;
        RECT 42.200 109.200 42.500 125.800 ;
        RECT 43.000 117.200 43.300 135.800 ;
        RECT 43.800 133.100 44.200 135.900 ;
        RECT 44.600 133.100 45.000 135.900 ;
        RECT 45.400 134.200 45.700 150.800 ;
        RECT 48.600 146.800 49.000 147.200 ;
        RECT 48.600 146.200 48.900 146.800 ;
        RECT 48.600 145.800 49.000 146.200 ;
        RECT 45.400 133.800 45.800 134.200 ;
        RECT 45.400 132.200 45.700 133.800 ;
        RECT 45.400 131.800 45.800 132.200 ;
        RECT 46.200 132.100 46.600 137.900 ;
        RECT 47.800 135.800 48.200 136.200 ;
        RECT 47.800 135.200 48.100 135.800 ;
        RECT 47.800 134.800 48.200 135.200 ;
        RECT 44.600 129.800 45.000 130.200 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 43.800 126.200 44.100 126.800 ;
        RECT 43.800 125.800 44.200 126.200 ;
        RECT 43.000 116.800 43.400 117.200 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 42.200 108.800 42.600 109.200 ;
        RECT 41.400 106.800 41.800 107.200 ;
        RECT 41.400 106.200 41.700 106.800 ;
        RECT 39.000 105.800 39.400 106.200 ;
        RECT 39.800 105.800 40.200 106.200 ;
        RECT 41.400 105.800 41.800 106.200 ;
        RECT 39.000 94.200 39.300 105.800 ;
        RECT 43.000 104.200 43.300 111.800 ;
        RECT 44.600 106.200 44.900 129.800 ;
        RECT 45.400 127.800 45.800 128.200 ;
        RECT 45.400 127.200 45.700 127.800 ;
        RECT 45.400 126.800 45.800 127.200 ;
        RECT 47.000 125.800 47.400 126.200 ;
        RECT 47.800 125.800 48.200 126.200 ;
        RECT 48.600 126.100 48.900 145.800 ;
        RECT 49.400 145.100 49.800 147.900 ;
        RECT 50.200 146.800 50.600 147.200 ;
        RECT 50.200 146.200 50.500 146.800 ;
        RECT 50.200 145.800 50.600 146.200 ;
        RECT 51.000 143.100 51.400 148.900 ;
        RECT 51.800 147.800 52.200 148.200 ;
        RECT 51.000 132.100 51.400 137.900 ;
        RECT 50.200 126.800 50.600 127.200 ;
        RECT 50.200 126.200 50.500 126.800 ;
        RECT 51.800 126.200 52.100 147.800 ;
        RECT 52.600 146.100 53.000 146.200 ;
        RECT 53.400 146.100 53.800 146.200 ;
        RECT 52.600 145.800 53.800 146.100 ;
        RECT 55.800 143.100 56.200 148.900 ;
        RECT 58.200 148.800 58.600 149.200 ;
        RECT 58.200 147.200 58.500 148.800 ;
        RECT 58.200 146.800 58.600 147.200 ;
        RECT 56.600 136.800 57.000 137.200 ;
        RECT 56.600 136.200 56.900 136.800 ;
        RECT 56.600 135.800 57.000 136.200 ;
        RECT 58.200 135.800 58.600 136.200 ;
        RECT 56.600 134.800 57.000 135.200 ;
        RECT 55.000 134.100 55.400 134.200 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 55.000 133.800 56.200 134.100 ;
        RECT 53.400 131.800 53.800 132.200 ;
        RECT 48.600 125.800 49.700 126.100 ;
        RECT 50.200 125.800 50.600 126.200 ;
        RECT 51.800 125.800 52.200 126.200 ;
        RECT 52.600 125.800 53.000 126.200 ;
        RECT 45.400 123.800 45.800 124.200 ;
        RECT 45.400 123.200 45.700 123.800 ;
        RECT 45.400 122.800 45.800 123.200 ;
        RECT 46.200 122.800 46.600 123.200 ;
        RECT 45.400 112.100 45.800 117.900 ;
        RECT 46.200 116.200 46.500 122.800 ;
        RECT 47.000 122.200 47.300 125.800 ;
        RECT 47.800 125.200 48.100 125.800 ;
        RECT 47.800 124.800 48.200 125.200 ;
        RECT 48.600 124.800 49.000 125.200 ;
        RECT 48.600 124.200 48.900 124.800 ;
        RECT 48.600 123.800 49.000 124.200 ;
        RECT 47.000 121.800 47.400 122.200 ;
        RECT 47.000 117.800 47.400 118.200 ;
        RECT 46.200 115.800 46.600 116.200 ;
        RECT 45.400 109.800 45.800 110.200 ;
        RECT 45.400 109.200 45.700 109.800 ;
        RECT 45.400 108.800 45.800 109.200 ;
        RECT 43.800 105.800 44.200 106.200 ;
        RECT 44.600 105.800 45.000 106.200 ;
        RECT 41.400 103.800 41.800 104.200 ;
        RECT 43.000 103.800 43.400 104.200 ;
        RECT 40.600 95.800 41.000 96.200 ;
        RECT 40.600 95.200 40.900 95.800 ;
        RECT 41.400 95.200 41.700 103.800 ;
        RECT 43.800 103.100 44.100 105.800 ;
        RECT 43.000 102.800 44.100 103.100 ;
        RECT 43.000 99.200 43.300 102.800 ;
        RECT 43.000 98.800 43.400 99.200 ;
        RECT 46.200 96.200 46.500 115.800 ;
        RECT 46.200 95.800 46.600 96.200 ;
        RECT 46.200 95.200 46.500 95.800 ;
        RECT 40.600 94.800 41.000 95.200 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 44.600 94.800 45.000 95.200 ;
        RECT 46.200 94.800 46.600 95.200 ;
        RECT 32.600 93.800 33.000 94.200 ;
        RECT 35.000 93.800 35.400 94.200 ;
        RECT 38.200 93.800 38.600 94.200 ;
        RECT 39.000 93.800 39.400 94.200 ;
        RECT 38.200 92.800 38.600 93.200 ;
        RECT 28.600 86.800 29.000 87.200 ;
        RECT 26.200 85.800 26.600 86.200 ;
        RECT 27.800 85.800 28.200 86.200 ;
        RECT 26.200 85.200 26.500 85.800 ;
        RECT 26.200 84.800 26.600 85.200 ;
        RECT 29.400 85.100 29.800 87.900 ;
        RECT 25.400 82.800 25.800 83.200 ;
        RECT 31.000 83.100 31.400 88.900 ;
        RECT 31.800 86.800 32.200 87.200 ;
        RECT 24.600 80.800 25.000 81.200 ;
        RECT 7.000 72.100 7.400 77.900 ;
        RECT 10.200 76.800 10.600 77.200 ;
        RECT 10.200 74.200 10.500 76.800 ;
        RECT 11.800 76.100 12.200 76.200 ;
        RECT 12.600 76.100 13.000 76.200 ;
        RECT 11.800 75.800 13.000 76.100 ;
        RECT 14.200 75.800 14.600 76.200 ;
        RECT 14.200 75.200 14.500 75.800 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 11.800 74.200 12.100 74.800 ;
        RECT 10.200 73.800 10.600 74.200 ;
        RECT 11.800 73.800 12.200 74.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 15.000 72.100 15.300 73.800 ;
        RECT 15.800 73.100 16.200 75.900 ;
        RECT 17.400 72.100 17.800 77.900 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 19.000 73.200 19.300 74.800 ;
        RECT 18.200 72.800 18.600 73.200 ;
        RECT 19.000 72.800 19.400 73.200 ;
        RECT 15.000 71.800 16.100 72.100 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 13.400 66.800 13.800 67.200 ;
        RECT 7.800 66.200 8.100 66.800 ;
        RECT 7.800 65.800 8.200 66.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 7.000 54.200 7.300 54.800 ;
        RECT 7.000 53.800 7.400 54.200 ;
        RECT 7.800 53.800 8.200 54.200 ;
        RECT 7.000 43.100 7.400 48.900 ;
        RECT 7.800 44.200 8.100 53.800 ;
        RECT 7.800 43.800 8.200 44.200 ;
        RECT 8.600 39.200 8.900 65.800 ;
        RECT 13.400 59.200 13.700 66.800 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 13.400 58.800 13.800 59.200 ;
        RECT 10.200 52.800 10.600 53.200 ;
        RECT 10.200 48.200 10.500 52.800 ;
        RECT 14.200 48.200 14.500 65.800 ;
        RECT 15.000 65.100 15.400 67.900 ;
        RECT 15.800 65.200 16.100 71.800 ;
        RECT 18.200 71.200 18.500 72.800 ;
        RECT 22.200 72.100 22.600 77.900 ;
        RECT 25.400 75.200 25.700 82.800 ;
        RECT 27.800 76.800 28.200 77.200 ;
        RECT 25.400 74.800 25.800 75.200 ;
        RECT 27.000 72.800 27.400 73.200 ;
        RECT 27.000 72.200 27.300 72.800 ;
        RECT 24.600 72.100 25.000 72.200 ;
        RECT 25.400 72.100 25.800 72.200 ;
        RECT 24.600 71.800 25.800 72.100 ;
        RECT 27.000 71.800 27.400 72.200 ;
        RECT 18.200 70.800 18.600 71.200 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 16.600 63.100 17.000 68.900 ;
        RECT 18.200 67.200 18.500 70.800 ;
        RECT 27.000 70.200 27.300 71.800 ;
        RECT 27.000 69.800 27.400 70.200 ;
        RECT 19.800 68.800 20.200 69.200 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 19.800 66.200 20.100 68.800 ;
        RECT 19.800 65.800 20.200 66.200 ;
        RECT 20.600 65.800 21.000 66.200 ;
        RECT 17.400 63.800 17.800 64.200 ;
        RECT 17.400 59.200 17.700 63.800 ;
        RECT 17.400 58.800 17.800 59.200 ;
        RECT 15.000 55.800 15.400 56.200 ;
        RECT 15.000 55.200 15.300 55.800 ;
        RECT 15.000 54.800 15.400 55.200 ;
        RECT 15.800 54.800 16.200 55.200 ;
        RECT 18.200 54.800 18.600 55.200 ;
        RECT 15.800 53.200 16.100 54.800 ;
        RECT 15.800 52.800 16.200 53.200 ;
        RECT 15.000 51.800 15.400 52.200 ;
        RECT 10.200 47.800 10.600 48.200 ;
        RECT 14.200 47.800 14.600 48.200 ;
        RECT 11.800 46.800 12.200 47.200 ;
        RECT 11.800 46.200 12.100 46.800 ;
        RECT 15.000 46.200 15.300 51.800 ;
        RECT 18.200 49.200 18.500 54.800 ;
        RECT 19.800 53.100 20.200 55.900 ;
        RECT 20.600 55.200 20.900 65.800 ;
        RECT 21.400 63.100 21.800 68.900 ;
        RECT 23.800 68.800 24.200 69.200 ;
        RECT 25.400 69.100 25.800 69.200 ;
        RECT 26.200 69.100 26.600 69.200 ;
        RECT 25.400 68.800 26.600 69.100 ;
        RECT 23.800 68.200 24.100 68.800 ;
        RECT 23.800 67.800 24.200 68.200 ;
        RECT 27.800 67.200 28.100 76.800 ;
        RECT 29.400 74.800 29.800 75.200 ;
        RECT 30.200 74.800 30.600 75.200 ;
        RECT 29.400 74.200 29.700 74.800 ;
        RECT 29.400 73.800 29.800 74.200 ;
        RECT 28.600 72.800 29.000 73.200 ;
        RECT 28.600 72.200 28.900 72.800 ;
        RECT 28.600 71.800 29.000 72.200 ;
        RECT 29.400 68.800 29.800 69.200 ;
        RECT 29.400 68.200 29.700 68.800 ;
        RECT 29.400 67.800 29.800 68.200 ;
        RECT 25.400 67.100 25.800 67.200 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 25.400 66.800 26.600 67.100 ;
        RECT 27.800 66.800 28.200 67.200 ;
        RECT 27.800 66.200 28.100 66.800 ;
        RECT 24.600 65.800 25.000 66.200 ;
        RECT 27.800 65.800 28.200 66.200 ;
        RECT 28.600 66.100 29.000 66.200 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 28.600 65.800 29.800 66.100 ;
        RECT 24.600 65.200 24.900 65.800 ;
        RECT 24.600 64.800 25.000 65.200 ;
        RECT 20.600 54.800 21.000 55.200 ;
        RECT 20.600 54.200 20.900 54.800 ;
        RECT 20.600 53.800 21.000 54.200 ;
        RECT 21.400 52.100 21.800 57.900 ;
        RECT 23.000 55.100 23.400 55.200 ;
        RECT 23.800 55.100 24.200 55.200 ;
        RECT 23.000 54.800 24.200 55.100 ;
        RECT 24.600 52.200 24.900 64.800 ;
        RECT 25.400 58.800 25.800 59.200 ;
        RECT 24.600 51.800 25.000 52.200 ;
        RECT 25.400 51.100 25.700 58.800 ;
        RECT 30.200 58.200 30.500 74.800 ;
        RECT 31.000 73.100 31.400 75.900 ;
        RECT 26.200 52.100 26.600 57.900 ;
        RECT 30.200 57.800 30.600 58.200 ;
        RECT 27.000 56.800 27.400 57.200 ;
        RECT 24.600 50.800 25.700 51.100 ;
        RECT 16.600 49.100 17.000 49.200 ;
        RECT 17.400 49.100 17.800 49.200 ;
        RECT 16.600 48.800 17.800 49.100 ;
        RECT 18.200 48.800 18.600 49.200 ;
        RECT 11.800 45.800 12.200 46.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.800 46.100 16.200 46.200 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 15.800 45.800 17.000 46.100 ;
        RECT 15.000 39.200 15.300 45.800 ;
        RECT 19.000 43.100 19.400 48.900 ;
        RECT 22.200 46.200 22.600 46.300 ;
        RECT 23.000 46.200 23.400 46.300 ;
        RECT 20.600 45.800 21.000 46.200 ;
        RECT 22.200 45.900 23.400 46.200 ;
        RECT 8.600 38.800 9.000 39.200 ;
        RECT 13.400 38.800 13.800 39.200 ;
        RECT 15.000 38.800 15.400 39.200 ;
        RECT 11.800 35.800 12.200 36.200 ;
        RECT 11.800 35.200 12.100 35.800 ;
        RECT 6.200 34.800 6.600 35.200 ;
        RECT 7.000 34.800 7.400 35.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 11.800 34.800 12.200 35.200 ;
        RECT 5.400 33.800 6.500 34.100 ;
        RECT 0.600 25.100 1.000 27.900 ;
        RECT 2.200 23.100 2.600 28.900 ;
        RECT 3.000 26.300 3.300 33.800 ;
        RECT 4.600 33.100 5.000 33.200 ;
        RECT 5.400 33.100 5.800 33.200 ;
        RECT 4.600 32.800 5.800 33.100 ;
        RECT 6.200 27.200 6.500 33.800 ;
        RECT 7.000 33.200 7.300 34.800 ;
        RECT 11.000 33.200 11.300 34.800 ;
        RECT 7.000 32.800 7.400 33.200 ;
        RECT 9.400 32.800 9.800 33.200 ;
        RECT 11.000 32.800 11.400 33.200 ;
        RECT 12.600 32.800 13.000 33.200 ;
        RECT 9.400 29.200 9.700 32.800 ;
        RECT 12.600 32.200 12.900 32.800 ;
        RECT 12.600 31.800 13.000 32.200 ;
        RECT 6.200 26.800 6.600 27.200 ;
        RECT 3.000 25.900 3.400 26.300 ;
        RECT 6.200 26.200 6.500 26.800 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 0.600 19.100 1.000 19.200 ;
        RECT 1.400 19.100 1.800 19.200 ;
        RECT 0.600 18.800 1.800 19.100 ;
        RECT 3.000 12.100 3.400 17.900 ;
        RECT 6.200 9.200 6.500 25.800 ;
        RECT 7.000 23.100 7.400 28.900 ;
        RECT 9.400 28.800 9.800 29.200 ;
        RECT 10.200 26.800 10.600 27.200 ;
        RECT 10.200 26.200 10.500 26.800 ;
        RECT 10.200 25.800 10.600 26.200 ;
        RECT 12.600 25.800 13.000 26.200 ;
        RECT 7.000 14.700 7.400 15.100 ;
        RECT 7.000 14.200 7.300 14.700 ;
        RECT 7.000 13.800 7.400 14.200 ;
        RECT 7.000 12.800 7.400 13.200 ;
        RECT 7.000 12.200 7.300 12.800 ;
        RECT 7.000 11.800 7.400 12.200 ;
        RECT 7.800 12.100 8.200 17.900 ;
        RECT 8.600 15.800 9.000 16.200 ;
        RECT 10.200 16.100 10.600 16.200 ;
        RECT 11.000 16.100 11.400 16.200 ;
        RECT 8.600 9.200 8.900 15.800 ;
        RECT 9.400 13.100 9.800 15.900 ;
        RECT 10.200 15.800 11.400 16.100 ;
        RECT 11.800 15.800 12.200 16.200 ;
        RECT 11.800 15.200 12.100 15.800 ;
        RECT 10.200 15.100 10.600 15.200 ;
        RECT 11.000 15.100 11.400 15.200 ;
        RECT 10.200 14.800 11.400 15.100 ;
        RECT 11.800 14.800 12.200 15.200 ;
        RECT 12.600 13.200 12.900 25.800 ;
        RECT 13.400 14.200 13.700 38.800 ;
        RECT 15.000 32.100 15.400 37.900 ;
        RECT 19.000 34.700 19.400 35.100 ;
        RECT 17.400 33.800 17.800 34.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 16.600 26.200 16.900 26.800 ;
        RECT 17.400 26.200 17.700 33.800 ;
        RECT 19.000 33.200 19.300 34.700 ;
        RECT 19.000 32.800 19.400 33.200 ;
        RECT 19.800 32.100 20.200 37.900 ;
        RECT 20.600 34.200 20.900 45.800 ;
        RECT 23.800 43.100 24.200 48.900 ;
        RECT 20.600 33.800 21.000 34.200 ;
        RECT 20.600 29.200 20.900 33.800 ;
        RECT 21.400 33.100 21.800 35.900 ;
        RECT 22.200 35.100 22.600 35.200 ;
        RECT 23.000 35.100 23.400 35.200 ;
        RECT 22.200 34.800 23.400 35.100 ;
        RECT 22.200 33.800 22.600 34.200 ;
        RECT 22.200 33.200 22.500 33.800 ;
        RECT 22.200 32.800 22.600 33.200 ;
        RECT 24.600 29.200 24.900 50.800 ;
        RECT 26.200 48.800 26.600 49.200 ;
        RECT 26.200 48.200 26.500 48.800 ;
        RECT 25.400 45.100 25.800 47.900 ;
        RECT 26.200 47.800 26.600 48.200 ;
        RECT 26.200 46.800 26.600 47.200 ;
        RECT 26.200 46.200 26.500 46.800 ;
        RECT 26.200 45.800 26.600 46.200 ;
        RECT 27.000 35.200 27.300 56.800 ;
        RECT 29.400 55.800 29.800 56.200 ;
        RECT 29.400 55.200 29.700 55.800 ;
        RECT 30.200 55.200 30.500 57.800 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 30.200 54.800 30.600 55.200 ;
        RECT 31.000 54.800 31.400 55.200 ;
        RECT 31.000 53.200 31.300 54.800 ;
        RECT 31.000 52.800 31.400 53.200 ;
        RECT 28.600 52.100 29.000 52.200 ;
        RECT 29.400 52.100 29.800 52.200 ;
        RECT 28.600 51.800 29.800 52.100 ;
        RECT 31.800 47.200 32.100 86.800 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 34.200 86.100 34.600 86.200 ;
        RECT 33.400 85.800 34.600 86.100 ;
        RECT 35.800 83.100 36.200 88.900 ;
        RECT 38.200 84.200 38.500 92.800 ;
        RECT 39.000 91.800 39.400 92.200 ;
        RECT 39.000 88.200 39.300 91.800 ;
        RECT 39.000 87.800 39.400 88.200 ;
        RECT 40.600 87.200 40.900 94.800 ;
        RECT 43.800 92.200 44.100 94.800 ;
        RECT 43.800 91.800 44.200 92.200 ;
        RECT 41.400 90.800 41.800 91.200 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 39.000 86.100 39.400 86.200 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 39.000 85.800 40.200 86.100 ;
        RECT 38.200 84.100 38.600 84.200 ;
        RECT 39.000 84.100 39.400 84.200 ;
        RECT 38.200 83.800 39.400 84.100 ;
        RECT 32.600 72.100 33.000 77.900 ;
        RECT 35.800 74.800 36.200 75.200 ;
        RECT 33.400 72.800 33.800 73.200 ;
        RECT 33.400 71.200 33.700 72.800 ;
        RECT 33.400 70.800 33.800 71.200 ;
        RECT 34.200 70.800 34.600 71.200 ;
        RECT 34.200 66.200 34.500 70.800 ;
        RECT 35.800 68.200 36.100 74.800 ;
        RECT 37.400 72.100 37.800 77.900 ;
        RECT 40.600 77.200 40.900 86.800 ;
        RECT 41.400 86.200 41.700 90.800 ;
        RECT 41.400 85.800 41.800 86.200 ;
        RECT 42.200 85.800 42.600 86.200 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 42.200 84.200 42.500 85.800 ;
        RECT 43.800 85.200 44.100 85.800 ;
        RECT 43.800 84.800 44.200 85.200 ;
        RECT 44.600 85.100 44.900 94.800 ;
        RECT 45.400 93.800 45.800 94.200 ;
        RECT 45.400 91.200 45.700 93.800 ;
        RECT 45.400 90.800 45.800 91.200 ;
        RECT 45.400 86.800 45.800 87.200 ;
        RECT 45.400 86.200 45.700 86.800 ;
        RECT 47.000 86.200 47.300 117.800 ;
        RECT 47.800 115.100 48.200 115.200 ;
        RECT 48.600 115.100 49.000 115.200 ;
        RECT 47.800 114.800 49.000 115.100 ;
        RECT 49.400 114.200 49.700 125.800 ;
        RECT 51.800 118.200 52.100 125.800 ;
        RECT 52.600 125.200 52.900 125.800 ;
        RECT 53.400 125.200 53.700 131.800 ;
        RECT 55.800 128.800 56.200 129.200 ;
        RECT 54.200 127.800 54.600 128.200 ;
        RECT 55.000 127.800 55.400 128.200 ;
        RECT 54.200 127.200 54.500 127.800 ;
        RECT 54.200 126.800 54.600 127.200 ;
        RECT 55.000 126.200 55.300 127.800 ;
        RECT 55.800 126.200 56.100 128.800 ;
        RECT 55.000 125.800 55.400 126.200 ;
        RECT 55.800 125.800 56.200 126.200 ;
        RECT 56.600 125.200 56.900 134.800 ;
        RECT 58.200 129.200 58.500 135.800 ;
        RECT 59.000 133.200 59.300 158.800 ;
        RECT 59.800 155.800 60.200 156.200 ;
        RECT 59.800 152.200 60.100 155.800 ;
        RECT 59.800 151.800 60.200 152.200 ;
        RECT 59.800 147.200 60.100 151.800 ;
        RECT 59.800 146.800 60.200 147.200 ;
        RECT 60.600 137.200 60.900 169.800 ;
        RECT 61.400 146.200 61.700 183.800 ;
        RECT 67.800 183.200 68.100 185.800 ;
        RECT 68.600 185.200 68.900 185.800 ;
        RECT 68.600 184.800 69.000 185.200 ;
        RECT 67.800 182.800 68.200 183.200 ;
        RECT 67.000 176.800 67.400 177.200 ;
        RECT 71.000 177.100 71.400 177.200 ;
        RECT 71.800 177.100 72.200 177.200 ;
        RECT 71.000 176.800 72.200 177.100 ;
        RECT 62.200 174.800 62.600 175.200 ;
        RECT 64.600 174.800 65.000 175.200 ;
        RECT 65.400 175.100 65.800 175.200 ;
        RECT 66.200 175.100 66.600 175.200 ;
        RECT 65.400 174.800 66.600 175.100 ;
        RECT 62.200 174.200 62.500 174.800 ;
        RECT 62.200 173.800 62.600 174.200 ;
        RECT 64.600 169.200 64.900 174.800 ;
        RECT 67.000 174.200 67.300 176.800 ;
        RECT 67.800 176.100 68.200 176.200 ;
        RECT 68.600 176.100 69.000 176.200 ;
        RECT 67.800 175.800 69.000 176.100 ;
        RECT 70.200 175.800 70.600 176.200 ;
        RECT 70.200 175.200 70.500 175.800 ;
        RECT 70.200 174.800 70.600 175.200 ;
        RECT 66.200 174.100 66.600 174.200 ;
        RECT 67.000 174.100 67.400 174.200 ;
        RECT 66.200 173.800 67.400 174.100 ;
        RECT 68.600 174.100 69.000 174.200 ;
        RECT 69.400 174.100 69.800 174.200 ;
        RECT 68.600 173.800 69.800 174.100 ;
        RECT 71.000 173.800 71.400 174.200 ;
        RECT 71.000 171.200 71.300 173.800 ;
        RECT 69.400 170.800 69.800 171.200 ;
        RECT 71.000 170.800 71.400 171.200 ;
        RECT 62.200 163.100 62.600 168.900 ;
        RECT 64.600 168.800 65.000 169.200 ;
        RECT 63.800 165.100 64.200 167.900 ;
        RECT 64.600 167.200 64.900 168.800 ;
        RECT 69.400 167.200 69.700 170.800 ;
        RECT 72.600 170.200 72.900 201.800 ;
        RECT 73.400 192.100 73.800 197.900 ;
        RECT 73.400 188.800 73.800 189.200 ;
        RECT 73.400 188.200 73.700 188.800 ;
        RECT 73.400 187.800 73.800 188.200 ;
        RECT 74.200 185.100 74.600 187.900 ;
        RECT 74.200 172.100 74.600 177.900 ;
        RECT 75.000 175.200 75.300 205.800 ;
        RECT 75.800 195.100 76.200 195.200 ;
        RECT 76.600 195.100 77.000 195.200 ;
        RECT 75.800 194.800 77.000 195.100 ;
        RECT 77.400 194.200 77.700 215.800 ;
        RECT 78.200 212.100 78.600 217.900 ;
        RECT 79.800 217.200 80.100 226.800 ;
        RECT 80.600 226.300 80.900 226.800 ;
        RECT 80.600 225.900 81.000 226.300 ;
        RECT 80.600 225.800 80.900 225.900 ;
        RECT 81.400 223.100 81.800 228.900 ;
        RECT 88.600 228.800 89.000 229.200 ;
        RECT 83.000 225.100 83.400 227.900 ;
        RECT 83.800 227.800 84.200 228.200 ;
        RECT 83.800 222.200 84.100 227.800 ;
        RECT 86.200 227.100 86.600 227.200 ;
        RECT 87.000 227.100 87.400 227.200 ;
        RECT 86.200 226.800 87.400 227.100 ;
        RECT 87.800 226.800 88.200 227.200 ;
        RECT 87.800 226.200 88.100 226.800 ;
        RECT 88.600 226.200 88.900 228.800 ;
        RECT 89.400 227.100 89.800 227.200 ;
        RECT 90.200 227.100 90.600 227.200 ;
        RECT 89.400 226.800 90.600 227.100 ;
        RECT 84.600 226.100 85.000 226.200 ;
        RECT 85.400 226.100 85.800 226.200 ;
        RECT 84.600 225.800 85.800 226.100 ;
        RECT 87.800 225.800 88.200 226.200 ;
        RECT 88.600 225.800 89.000 226.200 ;
        RECT 88.600 224.200 88.900 225.800 ;
        RECT 88.600 223.800 89.000 224.200 ;
        RECT 83.800 221.800 84.200 222.200 ;
        RECT 81.400 218.800 81.800 219.200 ;
        RECT 79.800 216.800 80.200 217.200 ;
        RECT 79.000 214.800 79.400 215.200 ;
        RECT 78.200 210.800 78.600 211.200 ;
        RECT 78.200 209.200 78.500 210.800 ;
        RECT 78.200 208.800 78.600 209.200 ;
        RECT 79.000 207.200 79.300 214.800 ;
        RECT 79.800 213.100 80.200 215.900 ;
        RECT 80.600 211.800 81.000 212.200 ;
        RECT 80.600 210.200 80.900 211.800 ;
        RECT 80.600 209.800 81.000 210.200 ;
        RECT 78.200 207.100 78.600 207.200 ;
        RECT 79.000 207.100 79.400 207.200 ;
        RECT 78.200 206.800 79.400 207.100 ;
        RECT 79.000 206.100 79.400 206.200 ;
        RECT 79.800 206.100 80.200 206.200 ;
        RECT 79.000 205.800 80.200 206.100 ;
        RECT 80.600 205.100 81.000 207.900 ;
        RECT 81.400 207.200 81.700 218.800 ;
        RECT 83.000 212.100 83.400 217.900 ;
        RECT 83.800 216.800 84.200 217.200 ;
        RECT 83.800 215.200 84.100 216.800 ;
        RECT 83.800 214.800 84.200 215.200 ;
        RECT 86.200 214.800 86.600 215.200 ;
        RECT 86.200 211.200 86.500 214.800 ;
        RECT 87.800 212.100 88.200 217.900 ;
        RECT 89.400 213.100 89.800 215.900 ;
        RECT 90.200 213.100 90.600 215.900 ;
        RECT 91.800 212.100 92.200 217.900 ;
        RECT 86.200 210.800 86.600 211.200 ;
        RECT 81.400 206.800 81.800 207.200 ;
        RECT 82.200 203.100 82.600 208.900 ;
        RECT 84.600 206.100 85.000 206.200 ;
        RECT 85.400 206.100 85.800 206.200 ;
        RECT 84.600 205.800 85.800 206.100 ;
        RECT 86.200 203.800 86.600 204.200 ;
        RECT 86.200 199.200 86.500 203.800 ;
        RECT 87.000 203.100 87.400 208.900 ;
        RECT 92.600 207.200 92.900 233.800 ;
        RECT 93.400 233.100 93.800 235.900 ;
        RECT 95.000 232.100 95.400 237.900 ;
        RECT 97.400 235.100 97.800 235.200 ;
        RECT 98.200 235.100 98.600 235.200 ;
        RECT 97.400 234.800 98.600 235.100 ;
        RECT 97.400 233.800 97.800 234.200 ;
        RECT 95.000 230.800 95.400 231.200 ;
        RECT 94.200 229.800 94.600 230.200 ;
        RECT 93.400 214.800 93.800 215.200 ;
        RECT 93.400 214.200 93.700 214.800 ;
        RECT 93.400 213.800 93.800 214.200 ;
        RECT 90.200 206.800 90.600 207.200 ;
        RECT 92.600 206.800 93.000 207.200 ;
        RECT 90.200 206.200 90.500 206.800 ;
        RECT 92.600 206.200 92.900 206.800 ;
        RECT 94.200 206.200 94.500 229.800 ;
        RECT 95.000 229.200 95.300 230.800 ;
        RECT 95.000 228.800 95.400 229.200 ;
        RECT 96.600 225.100 97.000 227.900 ;
        RECT 97.400 227.200 97.700 233.800 ;
        RECT 99.800 232.100 100.200 237.900 ;
        RECT 103.000 236.100 103.400 236.200 ;
        RECT 103.800 236.100 104.200 236.200 ;
        RECT 103.000 235.800 104.200 236.100 ;
        RECT 107.800 235.800 108.200 236.200 ;
        RECT 108.600 236.100 109.000 236.200 ;
        RECT 109.400 236.100 109.800 236.200 ;
        RECT 108.600 235.800 109.800 236.100 ;
        RECT 112.600 235.800 113.000 236.200 ;
        RECT 107.800 235.200 108.100 235.800 ;
        RECT 102.200 235.100 102.600 235.200 ;
        RECT 103.000 235.100 103.400 235.200 ;
        RECT 102.200 234.800 103.400 235.100 ;
        RECT 107.800 234.800 108.200 235.200 ;
        RECT 111.000 234.800 111.400 235.200 ;
        RECT 111.000 234.200 111.300 234.800 ;
        RECT 107.800 233.800 108.200 234.200 ;
        RECT 109.400 234.100 109.800 234.200 ;
        RECT 108.600 233.800 109.800 234.100 ;
        RECT 110.200 233.800 110.600 234.200 ;
        RECT 111.000 233.800 111.400 234.200 ;
        RECT 111.800 233.800 112.200 234.200 ;
        RECT 100.600 232.800 101.000 233.200 ;
        RECT 97.400 226.800 97.800 227.200 ;
        RECT 97.400 223.200 97.700 226.800 ;
        RECT 97.400 222.800 97.800 223.200 ;
        RECT 98.200 223.100 98.600 228.900 ;
        RECT 100.600 226.200 100.900 232.800 ;
        RECT 102.200 232.100 102.600 232.200 ;
        RECT 103.000 232.100 103.400 232.200 ;
        RECT 102.200 231.800 103.400 232.100 ;
        RECT 107.800 230.200 108.100 233.800 ;
        RECT 108.600 232.200 108.900 233.800 ;
        RECT 108.600 231.800 109.000 232.200 ;
        RECT 107.800 229.800 108.200 230.200 ;
        RECT 102.200 228.800 102.600 229.200 ;
        RECT 100.600 225.800 101.000 226.200 ;
        RECT 95.000 221.800 95.400 222.200 ;
        RECT 95.000 216.200 95.300 221.800 ;
        RECT 95.000 215.800 95.400 216.200 ;
        RECT 96.600 212.100 97.000 217.900 ;
        RECT 102.200 215.200 102.500 228.800 ;
        RECT 103.000 223.100 103.400 228.900 ;
        RECT 108.600 226.200 108.900 231.800 ;
        RECT 110.200 230.200 110.500 233.800 ;
        RECT 111.800 233.200 112.100 233.800 ;
        RECT 111.800 232.800 112.200 233.200 ;
        RECT 112.600 232.100 112.900 235.800 ;
        RECT 113.400 233.100 113.800 235.900 ;
        RECT 114.200 235.800 114.600 236.200 ;
        RECT 114.200 234.200 114.500 235.800 ;
        RECT 114.200 233.800 114.600 234.200 ;
        RECT 112.600 231.800 113.700 232.100 ;
        RECT 110.200 229.800 110.600 230.200 ;
        RECT 113.400 229.200 113.700 231.800 ;
        RECT 109.400 229.100 109.800 229.200 ;
        RECT 110.200 229.100 110.600 229.200 ;
        RECT 109.400 228.800 110.600 229.100 ;
        RECT 113.400 228.800 113.800 229.200 ;
        RECT 110.200 226.800 110.600 227.200 ;
        RECT 107.000 225.800 107.400 226.200 ;
        RECT 107.800 225.800 108.200 226.200 ;
        RECT 108.600 225.800 109.000 226.200 ;
        RECT 107.000 224.200 107.300 225.800 ;
        RECT 107.800 225.200 108.100 225.800 ;
        RECT 107.800 224.800 108.200 225.200 ;
        RECT 107.000 223.800 107.400 224.200 ;
        RECT 107.800 221.200 108.100 224.800 ;
        RECT 107.800 220.800 108.200 221.200 ;
        RECT 108.600 218.800 109.000 219.200 ;
        RECT 102.200 214.800 102.600 215.200 ;
        RECT 99.800 214.100 100.200 214.200 ;
        RECT 100.600 214.100 101.000 214.200 ;
        RECT 99.800 213.800 101.000 214.100 ;
        RECT 101.400 213.800 101.800 214.200 ;
        RECT 99.800 212.800 100.200 213.200 ;
        RECT 99.000 212.100 99.400 212.200 ;
        RECT 98.200 211.800 99.400 212.100 ;
        RECT 98.200 208.200 98.500 211.800 ;
        RECT 99.800 211.100 100.100 212.800 ;
        RECT 99.000 210.800 100.100 211.100 ;
        RECT 99.000 209.200 99.300 210.800 ;
        RECT 101.400 210.200 101.700 213.800 ;
        RECT 99.800 209.800 100.200 210.200 ;
        RECT 101.400 209.800 101.800 210.200 ;
        RECT 99.000 208.800 99.400 209.200 ;
        RECT 98.200 207.800 98.600 208.200 ;
        RECT 99.800 206.200 100.100 209.800 ;
        RECT 102.200 208.200 102.500 214.800 ;
        RECT 104.600 212.100 105.000 212.200 ;
        RECT 105.400 212.100 105.800 212.200 ;
        RECT 107.000 212.100 107.400 217.900 ;
        RECT 107.800 215.800 108.200 216.200 ;
        RECT 107.800 215.200 108.100 215.800 ;
        RECT 107.800 214.800 108.200 215.200 ;
        RECT 104.600 211.800 105.800 212.100 ;
        RECT 107.800 211.800 108.200 212.200 ;
        RECT 103.800 208.800 104.200 209.200 ;
        RECT 101.400 207.800 101.800 208.200 ;
        RECT 102.200 207.800 102.600 208.200 ;
        RECT 101.400 206.200 101.700 207.800 ;
        RECT 103.800 206.200 104.100 208.800 ;
        RECT 107.000 206.800 107.400 207.200 ;
        RECT 107.000 206.200 107.300 206.800 ;
        RECT 107.800 206.200 108.100 211.800 ;
        RECT 90.200 205.800 90.600 206.200 ;
        RECT 91.800 205.800 92.200 206.200 ;
        RECT 92.600 205.800 93.000 206.200 ;
        RECT 93.400 205.800 93.800 206.200 ;
        RECT 94.200 205.800 94.600 206.200 ;
        RECT 96.600 205.800 97.000 206.200 ;
        RECT 99.800 205.800 100.200 206.200 ;
        RECT 101.400 205.800 101.800 206.200 ;
        RECT 103.800 205.800 104.200 206.200 ;
        RECT 104.600 205.800 105.000 206.200 ;
        RECT 107.000 205.800 107.400 206.200 ;
        RECT 107.800 205.800 108.200 206.200 ;
        RECT 90.200 204.800 90.600 205.200 ;
        RECT 90.200 204.200 90.500 204.800 ;
        RECT 90.200 203.800 90.600 204.200 ;
        RECT 89.400 201.800 89.800 202.200 ;
        RECT 89.400 201.200 89.700 201.800 ;
        RECT 87.000 200.800 87.400 201.200 ;
        RECT 89.400 200.800 89.800 201.200 ;
        RECT 86.200 198.800 86.600 199.200 ;
        RECT 77.400 193.800 77.800 194.200 ;
        RECT 75.800 183.100 76.200 188.900 ;
        RECT 76.600 185.900 77.000 186.300 ;
        RECT 76.600 185.200 76.900 185.900 ;
        RECT 76.600 184.800 77.000 185.200 ;
        RECT 75.000 174.800 75.400 175.200 ;
        RECT 76.600 174.800 77.000 175.200 ;
        RECT 76.600 174.200 76.900 174.800 ;
        RECT 76.600 173.800 77.000 174.200 ;
        RECT 70.200 169.800 70.600 170.200 ;
        RECT 71.000 169.800 71.400 170.200 ;
        RECT 72.600 169.800 73.000 170.200 ;
        RECT 77.400 170.100 77.700 193.800 ;
        RECT 78.200 192.100 78.600 197.900 ;
        RECT 83.800 196.800 84.200 197.200 ;
        RECT 79.800 193.100 80.200 195.900 ;
        RECT 83.800 195.200 84.100 196.800 ;
        RECT 84.600 196.100 85.000 196.200 ;
        RECT 85.400 196.100 85.800 196.200 ;
        RECT 84.600 195.800 85.800 196.100 ;
        RECT 80.600 194.800 81.000 195.200 ;
        RECT 81.400 195.100 81.800 195.200 ;
        RECT 82.200 195.100 82.600 195.200 ;
        RECT 81.400 194.800 82.600 195.100 ;
        RECT 83.800 194.800 84.200 195.200 ;
        RECT 80.600 193.200 80.900 194.800 ;
        RECT 87.000 194.200 87.300 200.800 ;
        RECT 87.800 198.800 88.200 199.200 ;
        RECT 87.800 195.200 88.100 198.800 ;
        RECT 91.800 196.200 92.100 205.800 ;
        RECT 93.400 205.200 93.700 205.800 ;
        RECT 93.400 204.800 93.800 205.200 ;
        RECT 96.600 205.100 96.900 205.800 ;
        RECT 95.800 204.800 96.900 205.100 ;
        RECT 93.400 196.200 93.700 204.800 ;
        RECT 95.000 201.800 95.400 202.200 ;
        RECT 95.000 199.200 95.300 201.800 ;
        RECT 95.000 198.800 95.400 199.200 ;
        RECT 95.000 197.800 95.400 198.200 ;
        RECT 91.800 195.800 92.200 196.200 ;
        RECT 93.400 195.800 93.800 196.200 ;
        RECT 87.800 194.800 88.200 195.200 ;
        RECT 88.600 194.800 89.000 195.200 ;
        RECT 91.800 194.800 92.200 195.200 ;
        RECT 88.600 194.200 88.900 194.800 ;
        RECT 91.800 194.200 92.100 194.800 ;
        RECT 87.000 193.800 87.400 194.200 ;
        RECT 88.600 193.800 89.000 194.200 ;
        RECT 91.800 193.800 92.200 194.200 ;
        RECT 80.600 192.800 81.000 193.200 ;
        RECT 83.000 191.800 83.400 192.200 ;
        RECT 83.000 191.200 83.300 191.800 ;
        RECT 83.000 190.800 83.400 191.200 ;
        RECT 82.200 189.100 82.600 189.200 ;
        RECT 83.000 189.100 83.400 189.200 ;
        RECT 79.800 185.800 80.200 186.200 ;
        RECT 79.000 172.100 79.400 177.900 ;
        RECT 79.800 175.200 80.100 185.800 ;
        RECT 80.600 183.100 81.000 188.900 ;
        RECT 82.200 188.800 83.400 189.100 ;
        RECT 84.600 188.800 85.000 189.200 ;
        RECT 84.600 186.200 84.900 188.800 ;
        RECT 87.000 186.200 87.300 193.800 ;
        RECT 88.600 187.800 89.000 188.200 ;
        RECT 93.400 187.800 93.800 188.200 ;
        RECT 83.800 185.800 84.200 186.200 ;
        RECT 84.600 185.800 85.000 186.200 ;
        RECT 87.000 185.800 87.400 186.200 ;
        RECT 83.800 185.200 84.100 185.800 ;
        RECT 83.800 184.800 84.200 185.200 ;
        RECT 86.200 181.800 86.600 182.200 ;
        RECT 85.400 179.800 85.800 180.200 ;
        RECT 85.400 179.200 85.700 179.800 ;
        RECT 85.400 178.800 85.800 179.200 ;
        RECT 79.800 174.800 80.200 175.200 ;
        RECT 79.800 174.200 80.100 174.800 ;
        RECT 79.800 173.800 80.200 174.200 ;
        RECT 80.600 173.100 81.000 175.900 ;
        RECT 81.400 175.100 81.800 175.200 ;
        RECT 82.200 175.100 82.600 175.200 ;
        RECT 81.400 174.800 82.600 175.100 ;
        RECT 83.800 175.100 84.200 175.200 ;
        RECT 84.600 175.100 85.000 175.200 ;
        RECT 83.800 174.800 85.000 175.100 ;
        RECT 82.200 173.800 82.600 174.200 ;
        RECT 84.600 173.800 85.000 174.200 ;
        RECT 85.400 173.800 85.800 174.200 ;
        RECT 82.200 172.200 82.500 173.800 ;
        RECT 84.600 173.200 84.900 173.800 ;
        RECT 84.600 172.800 85.000 173.200 ;
        RECT 82.200 171.800 82.600 172.200 ;
        RECT 83.000 172.100 83.400 172.200 ;
        RECT 83.800 172.100 84.200 172.200 ;
        RECT 83.000 171.800 84.200 172.100 ;
        RECT 76.600 169.800 77.700 170.100 ;
        RECT 80.600 170.800 81.000 171.200 ;
        RECT 70.200 169.200 70.500 169.800 ;
        RECT 70.200 168.800 70.600 169.200 ;
        RECT 64.600 166.800 65.000 167.200 ;
        RECT 69.400 166.800 69.800 167.200 ;
        RECT 67.800 166.100 68.200 166.200 ;
        RECT 68.600 166.100 69.000 166.200 ;
        RECT 67.800 165.800 69.000 166.100 ;
        RECT 69.400 165.800 69.800 166.200 ;
        RECT 69.400 165.200 69.700 165.800 ;
        RECT 66.200 165.100 66.600 165.200 ;
        RECT 67.000 165.100 67.400 165.200 ;
        RECT 66.200 164.800 67.400 165.100 ;
        RECT 69.400 164.800 69.800 165.200 ;
        RECT 69.400 160.200 69.700 164.800 ;
        RECT 69.400 159.800 69.800 160.200 ;
        RECT 62.200 152.100 62.600 157.900 ;
        RECT 64.600 156.800 65.000 157.200 ;
        RECT 64.600 155.200 64.900 156.800 ;
        RECT 64.600 154.800 65.000 155.200 ;
        RECT 65.400 153.100 65.800 155.900 ;
        RECT 66.200 153.800 66.600 154.200 ;
        RECT 66.200 151.200 66.500 153.800 ;
        RECT 67.000 152.100 67.400 157.900 ;
        RECT 68.600 155.800 69.000 156.200 ;
        RECT 68.600 155.200 68.900 155.800 ;
        RECT 68.600 154.800 69.000 155.200 ;
        RECT 66.200 150.800 66.600 151.200 ;
        RECT 67.000 148.800 67.400 149.200 ;
        RECT 65.400 146.800 65.800 147.200 ;
        RECT 65.400 146.200 65.700 146.800 ;
        RECT 67.000 146.200 67.300 148.800 ;
        RECT 71.000 147.100 71.300 169.800 ;
        RECT 72.600 163.100 73.000 168.900 ;
        RECT 76.600 168.200 76.900 169.800 ;
        RECT 76.600 167.800 77.000 168.200 ;
        RECT 75.000 166.100 75.400 166.200 ;
        RECT 75.800 166.100 76.200 166.200 ;
        RECT 75.000 165.800 76.200 166.100 ;
        RECT 76.600 165.200 76.900 167.800 ;
        RECT 76.600 164.800 77.000 165.200 ;
        RECT 76.600 162.800 77.000 163.200 ;
        RECT 77.400 163.100 77.800 168.900 ;
        RECT 79.000 165.100 79.400 167.900 ;
        RECT 79.800 167.100 80.200 167.200 ;
        RECT 80.600 167.100 80.900 170.800 ;
        RECT 79.800 166.800 80.900 167.100 ;
        RECT 76.600 159.200 76.900 162.800 ;
        RECT 76.600 158.800 77.000 159.200 ;
        RECT 71.800 152.100 72.200 157.900 ;
        RECT 74.200 157.100 74.600 157.200 ;
        RECT 75.000 157.100 75.400 157.200 ;
        RECT 74.200 156.800 75.400 157.100 ;
        RECT 79.800 156.800 80.200 157.200 ;
        RECT 79.800 155.200 80.100 156.800 ;
        RECT 75.000 154.800 75.400 155.200 ;
        RECT 78.200 154.800 78.600 155.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 79.800 154.800 80.200 155.200 ;
        RECT 75.000 154.200 75.300 154.800 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 78.200 150.200 78.500 154.800 ;
        RECT 79.000 154.200 79.300 154.800 ;
        RECT 79.800 154.200 80.100 154.800 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 79.800 153.800 80.200 154.200 ;
        RECT 80.600 153.200 80.900 166.800 ;
        RECT 84.600 161.200 84.900 172.800 ;
        RECT 85.400 169.200 85.700 173.800 ;
        RECT 85.400 168.800 85.800 169.200 ;
        RECT 86.200 168.200 86.500 181.800 ;
        RECT 88.600 180.200 88.900 187.800 ;
        RECT 93.400 186.200 93.700 187.800 ;
        RECT 95.000 186.200 95.300 197.800 ;
        RECT 95.800 196.200 96.100 204.800 ;
        RECT 99.800 200.200 100.100 205.800 ;
        RECT 104.600 202.200 104.900 205.800 ;
        RECT 108.600 203.100 108.900 218.800 ;
        RECT 107.800 202.800 108.900 203.100 ;
        RECT 102.200 201.800 102.600 202.200 ;
        RECT 104.600 201.800 105.000 202.200 ;
        RECT 99.800 199.800 100.200 200.200 ;
        RECT 95.800 195.800 96.200 196.200 ;
        RECT 96.600 192.100 97.000 197.900 ;
        RECT 99.000 195.100 99.400 195.200 ;
        RECT 99.800 195.100 100.200 195.200 ;
        RECT 99.000 194.800 100.200 195.100 ;
        RECT 100.600 194.800 101.000 195.200 ;
        RECT 100.600 194.200 100.900 194.800 ;
        RECT 100.600 193.800 101.000 194.200 ;
        RECT 101.400 192.100 101.800 197.900 ;
        RECT 100.600 188.800 101.000 189.200 ;
        RECT 98.200 186.800 98.600 187.200 ;
        RECT 98.200 186.200 98.500 186.800 ;
        RECT 100.600 186.200 100.900 188.800 ;
        RECT 102.200 186.200 102.500 201.800 ;
        RECT 107.800 198.200 108.100 202.800 ;
        RECT 108.600 201.800 109.000 202.200 ;
        RECT 107.800 197.800 108.200 198.200 ;
        RECT 103.000 193.100 103.400 195.900 ;
        RECT 107.800 195.200 108.100 197.800 ;
        RECT 108.600 197.200 108.900 201.800 ;
        RECT 110.200 197.200 110.500 226.800 ;
        RECT 111.000 226.100 111.400 226.200 ;
        RECT 111.800 226.100 112.200 226.200 ;
        RECT 111.000 225.800 112.200 226.100 ;
        RECT 114.200 225.200 114.500 233.800 ;
        RECT 115.000 232.100 115.400 237.900 ;
        RECT 118.200 236.800 118.600 237.200 ;
        RECT 118.200 235.200 118.500 236.800 ;
        RECT 118.200 234.800 118.600 235.200 ;
        RECT 115.800 233.800 116.200 234.200 ;
        RECT 115.800 233.200 116.100 233.800 ;
        RECT 115.800 232.800 116.200 233.200 ;
        RECT 115.800 227.200 116.100 232.800 ;
        RECT 119.800 232.100 120.200 237.900 ;
        RECT 124.600 236.800 125.000 237.200 ;
        RECT 126.200 236.800 126.600 237.200 ;
        RECT 124.600 235.200 124.900 236.800 ;
        RECT 126.200 236.200 126.500 236.800 ;
        RECT 126.200 235.800 126.600 236.200 ;
        RECT 126.200 235.200 126.500 235.800 ;
        RECT 123.800 234.800 124.200 235.200 ;
        RECT 124.600 234.800 125.000 235.200 ;
        RECT 126.200 234.800 126.600 235.200 ;
        RECT 123.000 233.800 123.400 234.200 ;
        RECT 123.000 232.200 123.300 233.800 ;
        RECT 120.600 231.800 121.000 232.200 ;
        RECT 122.200 231.800 122.600 232.200 ;
        RECT 123.000 231.800 123.400 232.200 ;
        RECT 116.600 229.800 117.000 230.200 ;
        RECT 116.600 229.200 116.900 229.800 ;
        RECT 116.600 228.800 117.000 229.200 ;
        RECT 115.800 226.800 116.200 227.200 ;
        RECT 115.000 225.800 115.400 226.200 ;
        RECT 114.200 224.800 114.600 225.200 ;
        RECT 111.000 214.700 111.400 215.100 ;
        RECT 111.000 214.200 111.300 214.700 ;
        RECT 111.000 213.800 111.400 214.200 ;
        RECT 111.000 212.800 111.400 213.200 ;
        RECT 111.000 206.200 111.300 212.800 ;
        RECT 111.800 212.100 112.200 217.900 ;
        RECT 112.600 216.800 113.000 217.200 ;
        RECT 112.600 206.200 112.900 216.800 ;
        RECT 114.200 216.200 114.500 224.800 ;
        RECT 115.000 219.200 115.300 225.800 ;
        RECT 119.000 222.100 119.400 222.200 ;
        RECT 119.800 222.100 120.200 222.200 ;
        RECT 119.000 221.800 120.200 222.100 ;
        RECT 115.000 218.800 115.400 219.200 ;
        RECT 120.600 217.200 120.900 231.800 ;
        RECT 122.200 231.200 122.500 231.800 ;
        RECT 122.200 230.800 122.600 231.200 ;
        RECT 123.800 231.100 124.100 234.800 ;
        RECT 123.000 230.800 124.100 231.100 ;
        RECT 127.800 233.800 128.200 234.200 ;
        RECT 127.800 231.200 128.100 233.800 ;
        RECT 128.600 233.100 129.000 235.900 ;
        RECT 129.400 233.800 129.800 234.200 ;
        RECT 129.400 233.200 129.700 233.800 ;
        RECT 129.400 232.800 129.800 233.200 ;
        RECT 130.200 232.100 130.600 237.900 ;
        RECT 131.800 235.100 132.200 235.200 ;
        RECT 132.600 235.100 133.000 235.200 ;
        RECT 131.800 234.800 133.000 235.100 ;
        RECT 135.000 232.100 135.400 237.900 ;
        RECT 138.200 236.800 138.600 237.200 ;
        RECT 138.200 234.200 138.500 236.800 ;
        RECT 139.000 236.100 139.400 236.200 ;
        RECT 139.800 236.100 140.200 236.200 ;
        RECT 139.000 235.800 140.200 236.100 ;
        RECT 142.200 235.800 142.600 236.200 ;
        RECT 146.200 236.100 146.600 236.200 ;
        RECT 147.000 236.100 147.400 236.200 ;
        RECT 146.200 235.800 147.400 236.100 ;
        RECT 142.200 235.200 142.500 235.800 ;
        RECT 139.800 234.800 140.200 235.200 ;
        RECT 142.200 234.800 142.600 235.200 ;
        RECT 148.600 234.800 149.000 235.200 ;
        RECT 139.800 234.200 140.100 234.800 ;
        RECT 138.200 233.800 138.600 234.200 ;
        RECT 139.800 233.800 140.200 234.200 ;
        RECT 143.000 233.800 143.400 234.200 ;
        RECT 144.600 233.800 145.000 234.200 ;
        RECT 136.600 232.800 137.000 233.200 ;
        RECT 127.800 230.800 128.200 231.200 ;
        RECT 122.200 228.800 122.600 229.200 ;
        RECT 122.200 226.200 122.500 228.800 ;
        RECT 122.200 225.800 122.600 226.200 ;
        RECT 120.600 216.800 121.000 217.200 ;
        RECT 113.400 213.100 113.800 215.900 ;
        RECT 114.200 215.800 114.600 216.200 ;
        RECT 120.600 215.200 120.900 216.800 ;
        RECT 116.600 215.100 117.000 215.200 ;
        RECT 117.400 215.100 117.800 215.200 ;
        RECT 116.600 214.800 117.800 215.100 ;
        RECT 119.800 214.800 120.200 215.200 ;
        RECT 120.600 214.800 121.000 215.200 ;
        RECT 119.800 214.200 120.100 214.800 ;
        RECT 114.200 213.800 114.600 214.200 ;
        RECT 117.400 214.100 117.800 214.200 ;
        RECT 118.200 214.100 118.600 214.200 ;
        RECT 117.400 213.800 118.600 214.100 ;
        RECT 119.800 213.800 120.200 214.200 ;
        RECT 114.200 213.200 114.500 213.800 ;
        RECT 114.200 212.800 114.600 213.200 ;
        RECT 115.800 212.800 116.200 213.200 ;
        RECT 121.400 212.800 121.800 213.200 ;
        RECT 115.800 212.200 116.100 212.800 ;
        RECT 121.400 212.200 121.700 212.800 ;
        RECT 115.000 211.800 115.400 212.200 ;
        RECT 115.800 211.800 116.200 212.200 ;
        RECT 121.400 211.800 121.800 212.200 ;
        RECT 114.200 210.800 114.600 211.200 ;
        RECT 114.200 209.200 114.500 210.800 ;
        RECT 114.200 208.800 114.600 209.200 ;
        RECT 115.000 206.200 115.300 211.800 ;
        RECT 122.200 209.800 122.600 210.200 ;
        RECT 122.200 209.200 122.500 209.800 ;
        RECT 119.000 208.800 119.400 209.200 ;
        RECT 122.200 208.800 122.600 209.200 ;
        RECT 119.000 208.200 119.300 208.800 ;
        RECT 116.600 207.800 117.000 208.200 ;
        RECT 119.000 207.800 119.400 208.200 ;
        RECT 116.600 207.200 116.900 207.800 ;
        RECT 116.600 206.800 117.000 207.200 ;
        RECT 111.000 205.800 111.400 206.200 ;
        RECT 111.800 205.800 112.200 206.200 ;
        RECT 112.600 205.800 113.000 206.200 ;
        RECT 115.000 205.800 115.400 206.200 ;
        RECT 116.600 206.100 117.000 206.200 ;
        RECT 117.400 206.100 117.800 206.200 ;
        RECT 116.600 205.800 117.800 206.100 ;
        RECT 111.800 203.200 112.100 205.800 ;
        RECT 119.000 205.100 119.400 205.200 ;
        RECT 119.800 205.100 120.200 205.200 ;
        RECT 119.000 204.800 120.200 205.100 ;
        RECT 111.800 202.800 112.200 203.200 ;
        RECT 108.600 196.800 109.000 197.200 ;
        RECT 110.200 196.800 110.600 197.200 ;
        RECT 107.800 194.800 108.200 195.200 ;
        RECT 103.000 191.800 103.400 192.200 ;
        RECT 104.600 191.800 105.000 192.200 ;
        RECT 107.800 192.100 108.200 192.200 ;
        RECT 108.600 192.100 109.000 192.200 ;
        RECT 111.000 192.100 111.400 197.900 ;
        RECT 107.800 191.800 109.000 192.100 ;
        RECT 103.000 186.200 103.300 191.800 ;
        RECT 104.600 190.200 104.900 191.800 ;
        RECT 104.600 189.800 105.000 190.200 ;
        RECT 106.200 189.100 106.600 189.200 ;
        RECT 107.000 189.100 107.400 189.200 ;
        RECT 106.200 188.800 107.400 189.100 ;
        RECT 91.000 185.800 91.400 186.200 ;
        RECT 93.400 185.800 93.800 186.200 ;
        RECT 94.200 185.800 94.600 186.200 ;
        RECT 95.000 185.800 95.400 186.200 ;
        RECT 98.200 185.800 98.600 186.200 ;
        RECT 99.000 185.800 99.400 186.200 ;
        RECT 100.600 185.800 101.000 186.200 ;
        RECT 102.200 185.800 102.600 186.200 ;
        RECT 103.000 185.800 103.400 186.200 ;
        RECT 104.600 185.800 105.000 186.200 ;
        RECT 88.600 179.800 89.000 180.200 ;
        RECT 90.200 179.800 90.600 180.200 ;
        RECT 87.800 172.100 88.200 177.900 ;
        RECT 88.600 174.800 89.000 175.200 ;
        RECT 88.600 171.200 88.900 174.800 ;
        RECT 88.600 170.800 89.000 171.200 ;
        RECT 86.200 167.800 86.600 168.200 ;
        RECT 87.000 166.800 87.400 167.200 ;
        RECT 87.000 166.200 87.300 166.800 ;
        RECT 90.200 166.200 90.500 179.800 ;
        RECT 91.000 166.200 91.300 185.800 ;
        RECT 94.200 185.200 94.500 185.800 ;
        RECT 94.200 184.800 94.600 185.200 ;
        RECT 93.400 183.800 93.800 184.200 ;
        RECT 91.800 181.800 92.200 182.200 ;
        RECT 91.800 175.100 92.100 181.800 ;
        RECT 91.800 174.700 92.200 175.100 ;
        RECT 92.600 172.100 93.000 177.900 ;
        RECT 93.400 174.200 93.700 183.800 ;
        RECT 97.400 181.800 97.800 182.200 ;
        RECT 95.800 177.800 96.200 178.200 ;
        RECT 93.400 173.800 93.800 174.200 ;
        RECT 94.200 173.100 94.600 175.900 ;
        RECT 95.000 174.800 95.400 175.200 ;
        RECT 95.000 174.200 95.300 174.800 ;
        RECT 95.800 174.200 96.100 177.800 ;
        RECT 97.400 177.200 97.700 181.800 ;
        RECT 99.000 179.200 99.300 185.800 ;
        RECT 101.400 181.800 101.800 182.200 ;
        RECT 99.000 178.800 99.400 179.200 ;
        RECT 97.400 176.800 97.800 177.200 ;
        RECT 101.400 176.200 101.700 181.800 ;
        RECT 104.600 181.200 104.900 185.800 ;
        RECT 108.600 183.100 109.000 188.900 ;
        RECT 109.400 185.800 109.800 186.200 ;
        RECT 109.400 184.200 109.700 185.800 ;
        RECT 111.800 185.100 112.100 202.800 ;
        RECT 115.000 195.800 115.400 196.200 ;
        RECT 115.000 195.100 115.300 195.800 ;
        RECT 115.000 194.700 115.400 195.100 ;
        RECT 114.200 193.800 114.600 194.200 ;
        RECT 112.600 186.800 113.000 187.200 ;
        RECT 112.600 186.300 112.900 186.800 ;
        RECT 112.600 185.900 113.000 186.300 ;
        RECT 111.800 184.800 112.900 185.100 ;
        RECT 109.400 183.800 109.800 184.200 ;
        RECT 104.600 180.800 105.000 181.200 ;
        RECT 105.400 176.800 105.800 177.200 ;
        RECT 99.800 175.800 100.200 176.200 ;
        RECT 101.400 175.800 101.800 176.200 ;
        RECT 99.800 175.200 100.100 175.800 ;
        RECT 97.400 174.800 97.800 175.200 ;
        RECT 99.800 174.800 100.200 175.200 ;
        RECT 102.200 175.100 102.600 175.200 ;
        RECT 101.400 174.800 102.600 175.100 ;
        RECT 103.000 174.800 103.400 175.200 ;
        RECT 97.400 174.200 97.700 174.800 ;
        RECT 95.000 173.800 95.400 174.200 ;
        RECT 95.800 173.800 96.200 174.200 ;
        RECT 97.400 173.800 97.800 174.200 ;
        RECT 96.600 171.800 97.000 172.200 ;
        RECT 96.600 168.200 96.900 171.800 ;
        RECT 92.600 167.800 93.000 168.200 ;
        RECT 96.600 167.800 97.000 168.200 ;
        RECT 98.200 167.800 98.600 168.200 ;
        RECT 92.600 166.200 92.900 167.800 ;
        RECT 95.800 167.100 96.200 167.200 ;
        RECT 96.600 167.100 97.000 167.200 ;
        RECT 95.800 166.800 97.000 167.100 ;
        RECT 87.000 165.800 87.400 166.200 ;
        RECT 88.600 165.800 89.000 166.200 ;
        RECT 90.200 165.800 90.600 166.200 ;
        RECT 91.000 165.800 91.400 166.200 ;
        RECT 92.600 165.800 93.000 166.200 ;
        RECT 93.400 166.100 93.800 166.200 ;
        RECT 94.200 166.100 94.600 166.200 ;
        RECT 93.400 165.800 94.600 166.100 ;
        RECT 95.000 165.800 95.400 166.200 ;
        RECT 95.800 166.100 96.200 166.200 ;
        RECT 96.600 166.100 97.000 166.200 ;
        RECT 95.800 165.800 97.000 166.100 ;
        RECT 88.600 165.200 88.900 165.800 ;
        RECT 88.600 164.800 89.000 165.200 ;
        RECT 84.600 160.800 85.000 161.200 ;
        RECT 91.000 158.200 91.300 165.800 ;
        RECT 95.000 163.200 95.300 165.800 ;
        RECT 98.200 165.200 98.500 167.800 ;
        RECT 99.000 165.800 99.400 166.200 ;
        RECT 99.800 165.800 100.200 166.200 ;
        RECT 99.000 165.200 99.300 165.800 ;
        RECT 98.200 164.800 98.600 165.200 ;
        RECT 99.000 164.800 99.400 165.200 ;
        RECT 99.800 164.200 100.100 165.800 ;
        RECT 97.400 163.800 97.800 164.200 ;
        RECT 99.800 163.800 100.200 164.200 ;
        RECT 97.400 163.200 97.700 163.800 ;
        RECT 95.000 162.800 95.400 163.200 ;
        RECT 97.400 162.800 97.800 163.200 ;
        RECT 98.200 159.800 98.600 160.200 ;
        RECT 91.000 157.800 91.400 158.200 ;
        RECT 87.000 157.100 87.400 157.200 ;
        RECT 87.800 157.100 88.200 157.200 ;
        RECT 87.000 156.800 88.200 157.100 ;
        RECT 81.400 155.800 81.800 156.200 ;
        RECT 82.200 155.800 82.600 156.200 ;
        RECT 81.400 155.200 81.700 155.800 ;
        RECT 81.400 154.800 81.800 155.200 ;
        RECT 82.200 154.200 82.500 155.800 ;
        RECT 83.800 154.800 84.200 155.200 ;
        RECT 86.200 154.800 86.600 155.200 ;
        RECT 88.600 154.800 89.000 155.200 ;
        RECT 89.400 154.800 89.800 155.200 ;
        RECT 82.200 153.800 82.600 154.200 ;
        RECT 80.600 152.800 81.000 153.200 ;
        RECT 74.200 149.800 74.600 150.200 ;
        RECT 75.800 149.800 76.200 150.200 ;
        RECT 78.200 149.800 78.600 150.200 ;
        RECT 70.200 146.800 71.300 147.100 ;
        RECT 71.800 146.800 72.200 147.200 ;
        RECT 70.200 146.200 70.500 146.800 ;
        RECT 71.800 146.200 72.100 146.800 ;
        RECT 74.200 146.200 74.500 149.800 ;
        RECT 75.800 149.200 76.100 149.800 ;
        RECT 75.800 148.800 76.200 149.200 ;
        RECT 61.400 145.800 61.800 146.200 ;
        RECT 62.200 146.100 62.600 146.200 ;
        RECT 63.000 146.100 63.400 146.200 ;
        RECT 62.200 145.800 63.400 146.100 ;
        RECT 65.400 145.800 65.800 146.200 ;
        RECT 66.200 145.800 66.600 146.200 ;
        RECT 67.000 145.800 67.400 146.200 ;
        RECT 70.200 145.800 70.600 146.200 ;
        RECT 71.000 145.800 71.400 146.200 ;
        RECT 71.800 145.800 72.200 146.200 ;
        RECT 74.200 145.800 74.600 146.200 ;
        RECT 61.400 145.200 61.700 145.800 ;
        RECT 66.200 145.200 66.500 145.800 ;
        RECT 71.000 145.200 71.300 145.800 ;
        RECT 61.400 144.800 61.800 145.200 ;
        RECT 63.800 144.800 64.200 145.200 ;
        RECT 66.200 144.800 66.600 145.200 ;
        RECT 70.200 144.800 70.600 145.200 ;
        RECT 71.000 144.800 71.400 145.200 ;
        RECT 75.000 144.800 75.400 145.200 ;
        RECT 60.600 136.800 61.000 137.200 ;
        RECT 59.000 133.100 59.400 133.200 ;
        RECT 59.800 133.100 60.200 133.200 ;
        RECT 59.000 132.800 60.200 133.100 ;
        RECT 58.200 128.800 58.600 129.200 ;
        RECT 59.800 126.800 60.200 127.200 ;
        RECT 59.800 125.200 60.100 126.800 ;
        RECT 60.600 126.200 60.900 136.800 ;
        RECT 63.800 132.100 64.100 144.800 ;
        RECT 67.800 141.800 68.200 142.200 ;
        RECT 65.400 134.100 65.800 134.200 ;
        RECT 66.200 134.100 66.600 134.200 ;
        RECT 65.400 133.800 66.600 134.100 ;
        RECT 63.800 131.800 64.900 132.100 ;
        RECT 62.200 128.100 62.600 128.200 ;
        RECT 63.000 128.100 63.400 128.200 ;
        RECT 62.200 127.800 63.400 128.100 ;
        RECT 60.600 125.800 61.000 126.200 ;
        RECT 61.400 125.800 61.800 126.200 ;
        RECT 63.800 125.800 64.200 126.200 ;
        RECT 61.400 125.200 61.700 125.800 ;
        RECT 52.600 124.800 53.000 125.200 ;
        RECT 53.400 124.800 53.800 125.200 ;
        RECT 56.600 124.800 57.000 125.200 ;
        RECT 58.200 124.800 58.600 125.200 ;
        RECT 59.800 124.800 60.200 125.200 ;
        RECT 61.400 124.800 61.800 125.200 ;
        RECT 58.200 123.200 58.500 124.800 ;
        RECT 58.200 122.800 58.600 123.200 ;
        RECT 63.800 118.200 64.100 125.800 ;
        RECT 64.600 124.200 64.900 131.800 ;
        RECT 67.000 131.800 67.400 132.200 ;
        RECT 67.000 129.200 67.300 131.800 ;
        RECT 67.000 128.800 67.400 129.200 ;
        RECT 67.000 127.800 67.400 128.200 ;
        RECT 67.800 128.100 68.100 141.800 ;
        RECT 70.200 139.200 70.500 144.800 ;
        RECT 73.400 141.800 73.800 142.200 ;
        RECT 70.200 138.800 70.600 139.200 ;
        RECT 73.400 135.200 73.700 141.800 ;
        RECT 75.000 139.200 75.300 144.800 ;
        RECT 78.200 143.100 78.600 148.900 ;
        RECT 80.600 147.200 80.900 152.800 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 80.600 147.100 81.000 147.200 ;
        RECT 79.800 146.800 81.000 147.100 ;
        RECT 82.200 146.800 82.600 147.200 ;
        RECT 82.200 146.300 82.500 146.800 ;
        RECT 82.200 145.900 82.600 146.300 ;
        RECT 83.000 143.100 83.400 148.900 ;
        RECT 83.800 142.200 84.100 154.800 ;
        RECT 86.200 154.200 86.500 154.800 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 86.200 153.800 86.600 154.200 ;
        RECT 84.600 151.200 84.900 153.800 ;
        RECT 84.600 150.800 85.000 151.200 ;
        RECT 88.600 150.200 88.900 154.800 ;
        RECT 89.400 154.200 89.700 154.800 ;
        RECT 89.400 153.800 89.800 154.200 ;
        RECT 90.200 153.100 90.600 155.900 ;
        RECT 91.000 153.800 91.400 154.200 ;
        RECT 91.000 153.200 91.300 153.800 ;
        RECT 91.000 152.800 91.400 153.200 ;
        RECT 90.200 151.800 90.600 152.200 ;
        RECT 91.800 152.100 92.200 157.900 ;
        RECT 93.400 154.800 93.800 155.200 ;
        RECT 93.400 154.200 93.700 154.800 ;
        RECT 93.400 153.800 93.800 154.200 ;
        RECT 96.600 152.100 97.000 157.900 ;
        RECT 85.400 149.800 85.800 150.200 ;
        RECT 88.600 149.800 89.000 150.200 ;
        RECT 85.400 148.200 85.700 149.800 ;
        RECT 84.600 145.100 85.000 147.900 ;
        RECT 85.400 147.800 85.800 148.200 ;
        RECT 87.000 146.800 87.400 147.200 ;
        RECT 87.000 146.200 87.300 146.800 ;
        RECT 87.000 145.800 87.400 146.200 ;
        RECT 83.800 141.800 84.200 142.200 ;
        RECT 88.600 139.200 88.900 149.800 ;
        RECT 90.200 146.200 90.500 151.800 ;
        RECT 96.600 150.800 97.000 151.200 ;
        RECT 91.800 149.800 92.200 150.200 ;
        RECT 91.800 148.200 92.100 149.800 ;
        RECT 91.800 147.800 92.200 148.200 ;
        RECT 96.600 147.200 96.900 150.800 ;
        RECT 98.200 149.200 98.500 159.800 ;
        RECT 101.400 159.200 101.700 174.800 ;
        RECT 102.200 165.800 102.600 166.200 ;
        RECT 101.400 158.800 101.800 159.200 ;
        RECT 99.800 157.800 100.200 158.200 ;
        RECT 99.000 156.800 99.400 157.200 ;
        RECT 99.000 155.200 99.300 156.800 ;
        RECT 99.800 155.200 100.100 157.800 ;
        RECT 102.200 157.200 102.500 165.800 ;
        RECT 103.000 160.200 103.300 174.800 ;
        RECT 105.400 174.200 105.700 176.800 ;
        RECT 106.200 176.100 106.600 176.200 ;
        RECT 107.000 176.100 107.400 176.200 ;
        RECT 106.200 175.800 107.400 176.100 ;
        RECT 108.600 176.100 109.000 176.200 ;
        RECT 109.400 176.100 109.800 176.200 ;
        RECT 108.600 175.800 109.800 176.100 ;
        RECT 107.800 174.800 108.200 175.200 ;
        RECT 110.200 174.800 110.600 175.200 ;
        RECT 111.000 175.100 111.400 175.200 ;
        RECT 111.800 175.100 112.200 175.200 ;
        RECT 111.000 174.800 112.200 175.100 ;
        RECT 107.800 174.200 108.100 174.800 ;
        RECT 110.200 174.200 110.500 174.800 ;
        RECT 103.800 173.800 104.200 174.200 ;
        RECT 105.400 173.800 105.800 174.200 ;
        RECT 107.800 173.800 108.200 174.200 ;
        RECT 110.200 173.800 110.600 174.200 ;
        RECT 111.800 173.800 112.200 174.200 ;
        RECT 103.800 173.200 104.100 173.800 ;
        RECT 103.800 172.800 104.200 173.200 ;
        RECT 104.600 171.800 105.000 172.200 ;
        RECT 104.600 171.200 104.900 171.800 ;
        RECT 104.600 170.800 105.000 171.200 ;
        RECT 104.600 167.800 105.000 168.200 ;
        RECT 104.600 167.200 104.900 167.800 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 105.400 165.100 105.800 167.900 ;
        RECT 106.200 166.800 106.600 167.200 ;
        RECT 106.200 162.200 106.500 166.800 ;
        RECT 107.000 163.100 107.400 168.900 ;
        RECT 106.200 161.800 106.600 162.200 ;
        RECT 103.000 159.800 103.400 160.200 ;
        RECT 102.200 156.800 102.600 157.200 ;
        RECT 106.200 155.800 106.600 156.200 ;
        RECT 106.200 155.200 106.500 155.800 ;
        RECT 99.000 154.800 99.400 155.200 ;
        RECT 99.800 154.800 100.200 155.200 ;
        RECT 100.600 155.100 101.000 155.200 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 100.600 154.800 101.800 155.100 ;
        RECT 103.800 154.800 104.200 155.200 ;
        RECT 104.600 154.800 105.000 155.200 ;
        RECT 106.200 154.800 106.600 155.200 ;
        RECT 98.200 148.800 98.600 149.200 ;
        RECT 99.800 148.200 100.100 154.800 ;
        RECT 103.800 154.200 104.100 154.800 ;
        RECT 103.800 153.800 104.200 154.200 ;
        RECT 104.600 153.200 104.900 154.800 ;
        RECT 106.200 154.100 106.600 154.200 ;
        RECT 107.000 154.100 107.400 154.200 ;
        RECT 106.200 153.800 107.400 154.100 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 99.800 147.800 100.200 148.200 ;
        RECT 96.600 146.800 97.000 147.200 ;
        RECT 96.600 146.200 96.900 146.800 ;
        RECT 90.200 145.800 90.600 146.200 ;
        RECT 91.800 146.100 92.200 146.200 ;
        RECT 92.600 146.100 93.000 146.200 ;
        RECT 91.800 145.800 93.000 146.100 ;
        RECT 96.600 145.800 97.000 146.200 ;
        RECT 97.400 146.100 97.800 146.200 ;
        RECT 98.200 146.100 98.600 146.200 ;
        RECT 97.400 145.800 98.600 146.100 ;
        RECT 99.800 146.100 100.200 146.200 ;
        RECT 100.600 146.100 101.000 146.200 ;
        RECT 99.800 145.800 101.000 146.100 ;
        RECT 102.200 145.800 102.600 146.200 ;
        RECT 107.000 145.800 107.400 146.200 ;
        RECT 102.200 145.200 102.500 145.800 ;
        RECT 107.000 145.200 107.300 145.800 ;
        RECT 101.400 144.800 101.800 145.200 ;
        RECT 102.200 144.800 102.600 145.200 ;
        RECT 106.200 144.800 106.600 145.200 ;
        RECT 107.000 144.800 107.400 145.200 ;
        RECT 99.000 144.100 99.400 144.200 ;
        RECT 99.800 144.100 100.200 144.200 ;
        RECT 99.000 143.800 100.200 144.100 ;
        RECT 95.800 141.800 96.200 142.200 ;
        RECT 75.000 138.800 75.400 139.200 ;
        RECT 88.600 138.800 89.000 139.200 ;
        RECT 90.200 139.100 90.600 139.200 ;
        RECT 91.000 139.100 91.400 139.200 ;
        RECT 90.200 138.800 91.400 139.100 ;
        RECT 68.600 134.800 69.000 135.200 ;
        RECT 71.800 134.800 72.200 135.200 ;
        RECT 72.600 134.800 73.000 135.200 ;
        RECT 73.400 134.800 73.800 135.200 ;
        RECT 76.600 134.800 77.000 135.200 ;
        RECT 68.600 129.200 68.900 134.800 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 70.200 130.200 70.500 131.800 ;
        RECT 70.200 129.800 70.600 130.200 ;
        RECT 71.800 129.200 72.100 134.800 ;
        RECT 72.600 130.200 72.900 134.800 ;
        RECT 72.600 129.800 73.000 130.200 ;
        RECT 68.600 128.800 69.000 129.200 ;
        RECT 67.800 127.800 68.900 128.100 ;
        RECT 67.000 127.200 67.300 127.800 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 65.400 126.800 66.600 127.100 ;
        RECT 67.000 126.800 67.400 127.200 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 67.800 126.200 68.100 126.800 ;
        RECT 68.600 126.200 68.900 127.800 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 67.800 125.800 68.200 126.200 ;
        RECT 68.600 125.800 69.000 126.200 ;
        RECT 65.400 125.200 65.700 125.800 ;
        RECT 65.400 124.800 65.800 125.200 ;
        RECT 64.600 123.800 65.000 124.200 ;
        RECT 65.400 122.200 65.700 124.800 ;
        RECT 65.400 121.800 65.800 122.200 ;
        RECT 49.400 113.800 49.800 114.200 ;
        RECT 50.200 112.100 50.600 117.900 ;
        RECT 51.800 117.800 52.200 118.200 ;
        RECT 59.000 117.800 59.400 118.200 ;
        RECT 51.000 113.800 51.400 114.200 ;
        RECT 47.800 103.100 48.200 108.900 ;
        RECT 51.000 107.200 51.300 113.800 ;
        RECT 51.800 113.100 52.200 115.900 ;
        RECT 52.600 115.100 53.000 115.200 ;
        RECT 53.400 115.100 53.800 115.200 ;
        RECT 52.600 114.800 53.800 115.100 ;
        RECT 55.000 114.800 55.400 115.200 ;
        RECT 57.400 114.800 57.800 115.200 ;
        RECT 53.400 113.800 53.800 114.200 ;
        RECT 53.400 111.200 53.700 113.800 ;
        RECT 54.200 111.800 54.600 112.200 ;
        RECT 54.200 111.200 54.500 111.800 ;
        RECT 53.400 110.800 53.800 111.200 ;
        RECT 54.200 110.800 54.600 111.200 ;
        RECT 53.400 110.200 53.700 110.800 ;
        RECT 53.400 109.800 53.800 110.200 ;
        RECT 51.000 106.800 51.400 107.200 ;
        RECT 51.000 105.800 51.400 106.200 ;
        RECT 51.000 105.200 51.300 105.800 ;
        RECT 51.000 104.800 51.400 105.200 ;
        RECT 52.600 103.100 53.000 108.900 ;
        RECT 54.200 105.100 54.600 107.900 ;
        RECT 55.000 107.200 55.300 114.800 ;
        RECT 57.400 110.200 57.700 114.800 ;
        RECT 59.000 113.200 59.300 117.800 ;
        RECT 59.000 112.800 59.400 113.200 ;
        RECT 59.800 113.100 60.200 115.900 ;
        RECT 60.600 113.800 61.000 114.200 ;
        RECT 60.600 113.200 60.900 113.800 ;
        RECT 60.600 112.800 61.000 113.200 ;
        RECT 61.400 112.100 61.800 117.900 ;
        RECT 63.800 117.800 64.200 118.200 ;
        RECT 62.200 110.800 62.600 111.200 ;
        RECT 57.400 109.800 57.800 110.200 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 59.000 104.200 59.300 105.800 ;
        RECT 59.800 105.100 60.200 107.900 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 59.000 103.800 59.400 104.200 ;
        RECT 56.600 98.800 57.000 99.200 ;
        RECT 47.800 96.100 48.200 96.200 ;
        RECT 48.600 96.100 49.000 96.200 ;
        RECT 47.800 95.800 49.000 96.100 ;
        RECT 47.800 94.100 48.200 94.200 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 47.800 93.800 49.000 94.100 ;
        RECT 51.800 93.800 52.200 94.200 ;
        RECT 51.800 92.200 52.100 93.800 ;
        RECT 51.800 91.800 52.200 92.200 ;
        RECT 55.000 92.100 55.400 97.900 ;
        RECT 48.600 89.100 49.000 89.200 ;
        RECT 49.400 89.100 49.800 89.200 ;
        RECT 48.600 88.800 49.800 89.100 ;
        RECT 51.800 86.200 52.100 91.800 ;
        RECT 52.600 87.800 53.000 88.200 ;
        RECT 52.600 86.200 52.900 87.800 ;
        RECT 55.000 86.800 55.400 87.200 ;
        RECT 55.000 86.200 55.300 86.800 ;
        RECT 56.600 86.200 56.900 98.800 ;
        RECT 58.200 94.800 58.600 95.200 ;
        RECT 58.200 94.200 58.500 94.800 ;
        RECT 58.200 93.800 58.600 94.200 ;
        RECT 59.000 92.800 59.400 93.200 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 57.400 86.200 57.700 86.800 ;
        RECT 45.400 85.800 45.800 86.200 ;
        RECT 46.200 85.800 46.600 86.200 ;
        RECT 47.000 85.800 47.400 86.200 ;
        RECT 47.800 85.800 48.200 86.200 ;
        RECT 51.800 85.800 52.200 86.200 ;
        RECT 52.600 85.800 53.000 86.200 ;
        RECT 55.000 85.800 55.400 86.200 ;
        RECT 56.600 85.800 57.000 86.200 ;
        RECT 57.400 85.800 57.800 86.200 ;
        RECT 46.200 85.100 46.500 85.800 ;
        RECT 44.600 84.800 46.500 85.100 ;
        RECT 42.200 83.800 42.600 84.200 ;
        RECT 40.600 76.800 41.000 77.200 ;
        RECT 40.600 75.800 41.000 76.200 ;
        RECT 40.600 75.200 40.900 75.800 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 41.400 74.800 41.800 75.200 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 39.000 73.800 39.400 74.200 ;
        RECT 37.400 68.800 37.800 69.200 ;
        RECT 37.400 68.200 37.700 68.800 ;
        RECT 35.800 67.800 36.200 68.200 ;
        RECT 37.400 67.800 37.800 68.200 ;
        RECT 35.000 66.800 35.400 67.200 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 39.000 66.200 39.300 73.800 ;
        RECT 39.800 71.800 40.200 72.200 ;
        RECT 39.800 68.200 40.100 71.800 ;
        RECT 39.800 68.100 40.200 68.200 ;
        RECT 40.600 68.100 41.000 68.200 ;
        RECT 39.800 67.800 41.000 68.100 ;
        RECT 33.400 65.800 33.800 66.200 ;
        RECT 34.200 65.800 34.600 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 35.800 65.800 36.200 66.200 ;
        RECT 39.000 65.800 39.400 66.200 ;
        RECT 33.400 64.200 33.700 65.800 ;
        RECT 35.800 65.200 36.100 65.800 ;
        RECT 35.800 64.800 36.200 65.200 ;
        RECT 33.400 63.800 33.800 64.200 ;
        RECT 35.800 63.800 36.200 64.200 ;
        RECT 32.600 63.100 33.000 63.200 ;
        RECT 33.400 63.100 33.800 63.200 ;
        RECT 32.600 62.800 33.800 63.100 ;
        RECT 35.000 53.800 35.400 54.200 ;
        RECT 35.000 53.200 35.300 53.800 ;
        RECT 35.800 53.200 36.100 63.800 ;
        RECT 41.400 58.200 41.700 74.800 ;
        RECT 44.600 74.200 44.900 74.800 ;
        RECT 44.600 73.800 45.000 74.200 ;
        RECT 44.600 69.800 45.000 70.200 ;
        RECT 44.600 66.200 44.900 69.800 ;
        RECT 45.400 66.200 45.700 84.800 ;
        RECT 46.200 72.800 46.600 73.200 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 45.400 65.800 45.800 66.200 ;
        RECT 42.200 64.200 42.500 65.800 ;
        RECT 42.200 63.800 42.600 64.200 ;
        RECT 43.000 64.100 43.400 64.200 ;
        RECT 43.800 64.100 44.200 64.200 ;
        RECT 43.000 63.800 44.200 64.100 ;
        RECT 45.400 62.200 45.700 65.800 ;
        RECT 45.400 61.800 45.800 62.200 ;
        RECT 44.600 60.800 45.000 61.200 ;
        RECT 44.600 59.200 44.900 60.800 ;
        RECT 44.600 58.800 45.000 59.200 ;
        RECT 40.600 57.800 41.000 58.200 ;
        RECT 41.400 57.800 41.800 58.200 ;
        RECT 40.600 55.200 40.900 57.800 ;
        RECT 41.400 56.800 41.800 57.200 ;
        RECT 41.400 55.200 41.700 56.800 ;
        RECT 42.200 55.800 42.600 56.200 ;
        RECT 42.200 55.200 42.500 55.800 ;
        RECT 46.200 55.200 46.500 72.800 ;
        RECT 47.000 72.200 47.300 85.800 ;
        RECT 47.800 85.200 48.100 85.800 ;
        RECT 47.800 84.800 48.200 85.200 ;
        RECT 59.000 85.100 59.300 92.800 ;
        RECT 59.800 92.100 60.200 97.900 ;
        RECT 60.600 94.200 60.900 106.800 ;
        RECT 61.400 103.100 61.800 108.900 ;
        RECT 62.200 106.300 62.500 110.800 ;
        RECT 63.800 109.200 64.100 117.800 ;
        RECT 64.600 115.100 65.000 115.200 ;
        RECT 65.400 115.100 65.800 115.200 ;
        RECT 64.600 114.800 65.800 115.100 ;
        RECT 66.200 112.100 66.600 117.900 ;
        RECT 67.800 111.200 68.100 125.800 ;
        RECT 69.400 125.100 69.800 127.900 ;
        RECT 71.000 123.100 71.400 128.900 ;
        RECT 71.800 128.800 72.200 129.200 ;
        RECT 71.800 128.100 72.200 128.200 ;
        RECT 72.600 128.100 73.000 128.200 ;
        RECT 71.800 127.800 73.000 128.100 ;
        RECT 72.600 125.800 73.000 126.200 ;
        RECT 72.600 122.200 72.900 125.800 ;
        RECT 74.200 124.800 74.600 125.200 ;
        RECT 72.600 121.800 73.000 122.200 ;
        RECT 74.200 116.200 74.500 124.800 ;
        RECT 75.800 123.100 76.200 128.900 ;
        RECT 76.600 119.200 76.900 134.800 ;
        RECT 77.400 133.100 77.800 135.900 ;
        RECT 78.200 133.800 78.600 134.200 ;
        RECT 78.200 133.200 78.500 133.800 ;
        RECT 78.200 132.800 78.600 133.200 ;
        RECT 79.000 132.100 79.400 137.900 ;
        RECT 81.400 135.100 81.800 135.200 ;
        RECT 82.200 135.100 82.600 135.200 ;
        RECT 81.400 134.800 82.600 135.100 ;
        RECT 83.800 132.100 84.200 137.900 ;
        RECT 85.400 135.800 85.800 136.200 ;
        RECT 86.200 136.100 86.600 136.200 ;
        RECT 87.000 136.100 87.400 136.200 ;
        RECT 86.200 135.800 87.400 136.100 ;
        RECT 88.600 135.800 89.000 136.200 ;
        RECT 85.400 129.200 85.700 135.800 ;
        RECT 88.600 135.200 88.900 135.800 ;
        RECT 86.200 135.100 86.600 135.200 ;
        RECT 87.000 135.100 87.400 135.200 ;
        RECT 86.200 134.800 87.400 135.100 ;
        RECT 88.600 134.800 89.000 135.200 ;
        RECT 86.200 131.800 86.600 132.200 ;
        RECT 78.200 128.800 78.600 129.200 ;
        RECT 85.400 128.800 85.800 129.200 ;
        RECT 78.200 128.200 78.500 128.800 ;
        RECT 86.200 128.200 86.500 131.800 ;
        RECT 78.200 127.800 78.600 128.200 ;
        RECT 80.600 127.800 81.000 128.200 ;
        RECT 82.200 127.800 82.600 128.200 ;
        RECT 84.600 127.800 85.000 128.200 ;
        RECT 86.200 127.800 86.600 128.200 ;
        RECT 87.800 127.800 88.200 128.200 ;
        RECT 79.000 126.800 79.400 127.200 ;
        RECT 79.000 126.200 79.300 126.800 ;
        RECT 79.000 125.800 79.400 126.200 ;
        RECT 79.800 125.800 80.200 126.200 ;
        RECT 79.800 124.200 80.100 125.800 ;
        RECT 79.800 123.800 80.200 124.200 ;
        RECT 79.000 122.100 79.400 122.200 ;
        RECT 79.800 122.100 80.200 122.200 ;
        RECT 79.000 121.800 80.200 122.100 ;
        RECT 79.800 120.800 80.200 121.200 ;
        RECT 76.600 118.800 77.000 119.200 ;
        RECT 70.200 115.800 70.600 116.200 ;
        RECT 74.200 115.800 74.600 116.200 ;
        RECT 70.200 115.200 70.500 115.800 ;
        RECT 79.800 115.200 80.100 120.800 ;
        RECT 80.600 115.200 80.900 127.800 ;
        RECT 82.200 127.200 82.500 127.800 ;
        RECT 84.600 127.200 84.900 127.800 ;
        RECT 82.200 126.800 82.600 127.200 ;
        RECT 84.600 126.800 85.000 127.200 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 84.600 125.800 85.000 126.200 ;
        RECT 83.800 124.800 84.200 125.200 ;
        RECT 83.800 124.200 84.100 124.800 ;
        RECT 83.800 123.800 84.200 124.200 ;
        RECT 84.600 122.200 84.900 125.800 ;
        RECT 86.200 125.200 86.500 126.800 ;
        RECT 87.800 126.200 88.100 127.800 ;
        RECT 88.600 127.200 88.900 134.800 ;
        RECT 89.400 133.800 89.800 134.200 ;
        RECT 88.600 126.800 89.000 127.200 ;
        RECT 87.000 125.800 87.400 126.200 ;
        RECT 87.800 125.800 88.200 126.200 ;
        RECT 87.000 125.200 87.300 125.800 ;
        RECT 86.200 124.800 86.600 125.200 ;
        RECT 87.000 124.800 87.400 125.200 ;
        RECT 89.400 122.200 89.700 133.800 ;
        RECT 92.600 132.100 93.000 137.900 ;
        RECT 95.800 135.200 96.100 141.800 ;
        RECT 95.800 134.800 96.200 135.200 ;
        RECT 97.400 132.100 97.800 137.900 ;
        RECT 99.800 136.800 100.200 137.200 ;
        RECT 100.600 136.800 101.000 137.200 ;
        RECT 99.800 136.200 100.100 136.800 ;
        RECT 100.600 136.200 100.900 136.800 ;
        RECT 98.200 133.800 98.600 134.200 ;
        RECT 98.200 132.200 98.500 133.800 ;
        RECT 99.000 133.100 99.400 135.900 ;
        RECT 99.800 135.800 100.200 136.200 ;
        RECT 100.600 135.800 101.000 136.200 ;
        RECT 101.400 136.100 101.700 144.800 ;
        RECT 102.200 143.800 102.600 144.200 ;
        RECT 103.000 144.100 103.400 144.200 ;
        RECT 103.800 144.100 104.200 144.200 ;
        RECT 103.000 143.800 104.200 144.100 ;
        RECT 102.200 143.200 102.500 143.800 ;
        RECT 102.200 142.800 102.600 143.200 ;
        RECT 103.800 138.800 104.200 139.200 ;
        RECT 103.800 138.200 104.100 138.800 ;
        RECT 103.800 137.800 104.200 138.200 ;
        RECT 104.600 136.800 105.000 137.200 ;
        RECT 104.600 136.200 104.900 136.800 ;
        RECT 102.200 136.100 102.600 136.200 ;
        RECT 101.400 135.800 102.600 136.100 ;
        RECT 104.600 135.800 105.000 136.200 ;
        RECT 102.200 135.200 102.500 135.800 ;
        RECT 106.200 135.200 106.500 144.800 ;
        RECT 107.800 144.200 108.100 173.800 ;
        RECT 110.200 173.200 110.500 173.800 ;
        RECT 110.200 172.800 110.600 173.200 ;
        RECT 111.800 172.200 112.100 173.800 ;
        RECT 111.800 171.800 112.200 172.200 ;
        RECT 108.600 166.800 109.000 167.200 ;
        RECT 108.600 166.200 108.900 166.800 ;
        RECT 108.600 165.800 109.000 166.200 ;
        RECT 111.800 163.100 112.200 168.900 ;
        RECT 112.600 159.200 112.900 184.800 ;
        RECT 113.400 183.100 113.800 188.900 ;
        RECT 114.200 187.200 114.500 193.800 ;
        RECT 115.800 192.100 116.200 197.900 ;
        RECT 117.400 193.100 117.800 195.900 ;
        RECT 119.800 195.800 120.200 196.200 ;
        RECT 121.400 195.800 121.800 196.200 ;
        RECT 119.800 195.200 120.100 195.800 ;
        RECT 121.400 195.200 121.700 195.800 ;
        RECT 119.800 194.800 120.200 195.200 ;
        RECT 121.400 194.800 121.800 195.200 ;
        RECT 122.200 195.100 122.600 195.200 ;
        RECT 123.000 195.100 123.300 230.800 ;
        RECT 125.400 226.800 125.800 227.200 ;
        RECT 125.400 226.200 125.700 226.800 ;
        RECT 127.800 226.200 128.100 230.800 ;
        RECT 135.800 228.800 136.200 229.200 ;
        RECT 135.800 227.200 136.100 228.800 ;
        RECT 130.200 226.800 130.600 227.200 ;
        RECT 135.800 226.800 136.200 227.200 ;
        RECT 130.200 226.200 130.500 226.800 ;
        RECT 135.800 226.200 136.100 226.800 ;
        RECT 136.600 226.200 136.900 232.800 ;
        RECT 138.200 227.200 138.500 233.800 ;
        RECT 143.000 232.200 143.300 233.800 ;
        RECT 143.000 231.800 143.400 232.200 ;
        RECT 141.400 229.100 141.800 229.200 ;
        RECT 142.200 229.100 142.600 229.200 ;
        RECT 141.400 228.800 142.600 229.100 ;
        RECT 138.200 226.800 138.600 227.200 ;
        RECT 141.400 226.800 141.800 227.200 ;
        RECT 141.400 226.200 141.700 226.800 ;
        RECT 125.400 225.800 125.800 226.200 ;
        RECT 126.200 225.800 126.600 226.200 ;
        RECT 127.000 225.800 127.400 226.200 ;
        RECT 127.800 225.800 128.200 226.200 ;
        RECT 130.200 225.800 130.600 226.200 ;
        RECT 131.000 226.100 131.400 226.200 ;
        RECT 131.800 226.100 132.200 226.200 ;
        RECT 131.000 225.800 132.200 226.100 ;
        RECT 132.600 226.100 133.000 226.200 ;
        RECT 133.400 226.100 133.800 226.200 ;
        RECT 132.600 225.800 133.800 226.100 ;
        RECT 135.800 225.800 136.200 226.200 ;
        RECT 136.600 225.800 137.000 226.200 ;
        RECT 138.200 225.800 138.600 226.200 ;
        RECT 139.800 226.100 140.200 226.200 ;
        RECT 140.600 226.100 141.000 226.200 ;
        RECT 139.800 225.800 141.000 226.100 ;
        RECT 141.400 225.800 141.800 226.200 ;
        RECT 142.200 225.800 142.600 226.200 ;
        RECT 126.200 225.200 126.500 225.800 ;
        RECT 126.200 224.800 126.600 225.200 ;
        RECT 127.000 224.200 127.300 225.800 ;
        RECT 138.200 225.200 138.500 225.800 ;
        RECT 138.200 224.800 138.600 225.200 ;
        RECT 140.600 225.100 141.000 225.200 ;
        RECT 142.200 225.100 142.500 225.800 ;
        RECT 140.600 224.800 142.500 225.100 ;
        RECT 138.200 224.200 138.500 224.800 ;
        RECT 127.000 223.800 127.400 224.200 ;
        RECT 138.200 223.800 138.600 224.200 ;
        RECT 123.800 221.800 124.200 222.200 ;
        RECT 123.800 221.200 124.100 221.800 ;
        RECT 127.000 221.200 127.300 223.800 ;
        RECT 143.000 223.200 143.300 231.800 ;
        RECT 144.600 230.200 144.900 233.800 ;
        RECT 146.200 233.100 146.600 233.200 ;
        RECT 147.000 233.100 147.400 233.200 ;
        RECT 146.200 232.800 147.400 233.100 ;
        RECT 148.600 230.200 148.900 234.800 ;
        RECT 149.400 232.800 149.800 233.200 ;
        RECT 149.400 232.200 149.700 232.800 ;
        RECT 149.400 231.800 149.800 232.200 ;
        RECT 151.800 232.100 152.200 237.900 ;
        RECT 153.400 235.800 153.800 236.200 ;
        RECT 153.400 235.200 153.700 235.800 ;
        RECT 152.600 234.800 153.000 235.200 ;
        RECT 153.400 234.800 153.800 235.200 ;
        RECT 144.600 229.800 145.000 230.200 ;
        RECT 148.600 229.800 149.000 230.200 ;
        RECT 152.600 229.200 152.900 234.800 ;
        RECT 156.600 232.100 157.000 237.900 ;
        RECT 160.600 236.800 161.000 237.200 ;
        RECT 162.200 236.800 162.600 237.200 ;
        RECT 160.600 236.200 160.900 236.800 ;
        RECT 158.200 233.100 158.600 235.900 ;
        RECT 160.600 235.800 161.000 236.200 ;
        RECT 160.600 234.200 160.900 235.800 ;
        RECT 162.200 234.200 162.500 236.800 ;
        RECT 163.800 235.800 164.200 236.200 ;
        RECT 163.800 235.200 164.100 235.800 ;
        RECT 163.800 234.800 164.200 235.200 ;
        RECT 164.600 234.800 165.000 235.200 ;
        RECT 164.600 234.200 164.900 234.800 ;
        RECT 160.600 233.800 161.000 234.200 ;
        RECT 162.200 233.800 162.600 234.200 ;
        RECT 164.600 233.800 165.000 234.200 ;
        RECT 165.400 233.800 165.800 234.200 ;
        RECT 165.400 233.200 165.700 233.800 ;
        RECT 165.400 232.800 165.800 233.200 ;
        RECT 166.200 233.100 166.600 235.900 ;
        RECT 167.800 232.100 168.200 237.900 ;
        RECT 168.600 235.800 169.000 236.200 ;
        RECT 168.600 235.100 168.900 235.800 ;
        RECT 168.600 234.700 169.000 235.100 ;
        RECT 168.600 232.800 169.000 233.200 ;
        RECT 140.600 222.800 141.000 223.200 ;
        RECT 143.000 222.800 143.400 223.200 ;
        RECT 144.600 223.100 145.000 228.900 ;
        RECT 148.600 228.800 149.000 229.200 ;
        RECT 148.600 227.200 148.900 228.800 ;
        RECT 148.600 226.800 149.000 227.200 ;
        RECT 147.000 226.100 147.400 226.200 ;
        RECT 147.800 226.100 148.200 226.200 ;
        RECT 147.000 225.800 148.200 226.100 ;
        RECT 129.400 221.800 129.800 222.200 ;
        RECT 134.200 221.800 134.600 222.200 ;
        RECT 138.200 221.800 138.600 222.200 ;
        RECT 123.800 220.800 124.200 221.200 ;
        RECT 127.000 220.800 127.400 221.200 ;
        RECT 123.800 212.100 124.200 217.900 ;
        RECT 126.200 217.800 126.600 218.200 ;
        RECT 124.600 203.100 125.000 208.900 ;
        RECT 122.200 194.800 123.300 195.100 ;
        RECT 126.200 195.200 126.500 217.800 ;
        RECT 127.000 214.800 127.400 215.200 ;
        RECT 127.000 211.200 127.300 214.800 ;
        RECT 128.600 212.100 129.000 217.900 ;
        RECT 129.400 215.200 129.700 221.800 ;
        RECT 129.400 214.800 129.800 215.200 ;
        RECT 129.400 213.800 129.800 214.200 ;
        RECT 129.400 213.200 129.700 213.800 ;
        RECT 129.400 212.800 129.800 213.200 ;
        RECT 130.200 213.100 130.600 215.900 ;
        RECT 134.200 215.200 134.500 221.800 ;
        RECT 138.200 215.200 138.500 221.800 ;
        RECT 140.600 219.200 140.900 222.800 ;
        RECT 140.600 218.800 141.000 219.200 ;
        RECT 148.600 215.200 148.900 226.800 ;
        RECT 149.400 223.100 149.800 228.900 ;
        RECT 152.600 228.800 153.000 229.200 ;
        RECT 155.000 228.800 155.400 229.200 ;
        RECT 163.000 228.800 163.400 229.200 ;
        RECT 151.000 225.100 151.400 227.900 ;
        RECT 155.000 226.200 155.300 228.800 ;
        RECT 163.000 227.200 163.300 228.800 ;
        RECT 155.800 226.800 156.200 227.200 ;
        RECT 159.000 226.800 159.400 227.200 ;
        RECT 163.000 226.800 163.400 227.200 ;
        RECT 155.800 226.200 156.100 226.800 ;
        RECT 159.000 226.200 159.300 226.800 ;
        RECT 151.800 225.800 152.200 226.200 ;
        RECT 152.600 226.100 153.000 226.200 ;
        RECT 153.400 226.100 153.800 226.200 ;
        RECT 152.600 225.800 153.800 226.100 ;
        RECT 155.000 225.800 155.400 226.200 ;
        RECT 155.800 225.800 156.200 226.200 ;
        RECT 159.000 225.800 159.400 226.200 ;
        RECT 161.400 225.800 161.800 226.200 ;
        RECT 162.200 225.800 162.600 226.200 ;
        RECT 151.800 225.200 152.100 225.800 ;
        RECT 151.800 224.800 152.200 225.200 ;
        RECT 153.400 221.800 153.800 222.200 ;
        RECT 153.400 220.200 153.700 221.800 ;
        RECT 153.400 219.800 153.800 220.200 ;
        RECT 131.000 215.100 131.400 215.200 ;
        RECT 131.800 215.100 132.200 215.200 ;
        RECT 131.000 214.800 132.200 215.100 ;
        RECT 134.200 214.800 134.600 215.200 ;
        RECT 135.000 214.800 135.400 215.200 ;
        RECT 138.200 214.800 138.600 215.200 ;
        RECT 148.600 214.800 149.000 215.200 ;
        RECT 135.000 214.200 135.300 214.800 ;
        RECT 148.600 214.200 148.900 214.800 ;
        RECT 135.000 213.800 135.400 214.200 ;
        RECT 142.200 213.800 142.600 214.200 ;
        RECT 148.600 213.800 149.000 214.200 ;
        RECT 142.200 213.200 142.500 213.800 ;
        RECT 142.200 212.800 142.600 213.200 ;
        RECT 132.600 212.100 133.000 212.200 ;
        RECT 133.400 212.100 133.800 212.200 ;
        RECT 132.600 211.800 133.800 212.100 ;
        RECT 136.600 211.800 137.000 212.200 ;
        RECT 149.400 212.100 149.800 212.200 ;
        RECT 150.200 212.100 150.600 212.200 ;
        RECT 149.400 211.800 150.600 212.100 ;
        RECT 151.000 211.800 151.400 212.200 ;
        RECT 151.800 212.100 152.200 217.900 ;
        RECT 152.600 215.800 153.000 216.200 ;
        RECT 152.600 215.200 152.900 215.800 ;
        RECT 152.600 214.800 153.000 215.200 ;
        RECT 155.000 214.800 155.400 215.200 ;
        RECT 127.000 210.800 127.400 211.200 ;
        RECT 127.800 207.800 128.200 208.200 ;
        RECT 127.800 206.200 128.100 207.800 ;
        RECT 127.800 205.800 128.200 206.200 ;
        RECT 129.400 203.100 129.800 208.900 ;
        RECT 130.200 206.800 130.600 207.200 ;
        RECT 128.600 196.800 129.000 197.200 ;
        RECT 127.000 195.800 127.400 196.200 ;
        RECT 127.000 195.200 127.300 195.800 ;
        RECT 126.200 194.800 126.600 195.200 ;
        RECT 127.000 194.800 127.400 195.200 ;
        RECT 118.200 193.800 118.600 194.200 ;
        RECT 118.200 192.200 118.500 193.800 ;
        RECT 118.200 191.800 118.600 192.200 ;
        RECT 115.800 188.800 116.200 189.200 ;
        RECT 114.200 186.800 114.600 187.200 ;
        RECT 114.200 186.200 114.500 186.800 ;
        RECT 114.200 185.800 114.600 186.200 ;
        RECT 115.000 185.100 115.400 187.900 ;
        RECT 115.800 187.200 116.100 188.800 ;
        RECT 120.600 187.800 121.000 188.200 ;
        RECT 120.600 187.200 120.900 187.800 ;
        RECT 115.800 186.800 116.200 187.200 ;
        RECT 117.400 187.100 117.800 187.200 ;
        RECT 118.200 187.100 118.600 187.200 ;
        RECT 117.400 186.800 118.600 187.100 ;
        RECT 120.600 186.800 121.000 187.200 ;
        RECT 121.400 186.800 121.800 187.200 ;
        RECT 121.400 186.200 121.700 186.800 ;
        RECT 119.800 185.800 120.200 186.200 ;
        RECT 121.400 185.800 121.800 186.200 ;
        RECT 119.800 185.200 120.100 185.800 ;
        RECT 122.200 185.200 122.500 194.800 ;
        RECT 123.000 193.800 123.400 194.200 ;
        RECT 123.000 187.200 123.300 193.800 ;
        RECT 126.200 190.200 126.500 194.800 ;
        RECT 128.600 194.200 128.900 196.800 ;
        RECT 128.600 193.800 129.000 194.200 ;
        RECT 130.200 193.200 130.500 206.800 ;
        RECT 131.000 205.100 131.400 207.900 ;
        RECT 131.800 205.100 132.200 207.900 ;
        RECT 133.400 203.100 133.800 208.900 ;
        RECT 136.600 208.200 136.900 211.800 ;
        RECT 140.600 209.100 141.000 209.200 ;
        RECT 141.400 209.100 141.800 209.200 ;
        RECT 136.600 207.800 137.000 208.200 ;
        RECT 135.800 206.800 136.200 207.200 ;
        RECT 135.000 205.800 135.400 206.200 ;
        RECT 135.000 204.200 135.300 205.800 ;
        RECT 135.000 203.800 135.400 204.200 ;
        RECT 131.000 196.100 131.400 196.200 ;
        RECT 131.800 196.100 132.200 196.200 ;
        RECT 131.000 195.800 132.200 196.100 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 131.800 194.800 132.200 195.200 ;
        RECT 131.000 194.200 131.300 194.800 ;
        RECT 131.800 194.200 132.100 194.800 ;
        RECT 131.000 193.800 131.400 194.200 ;
        RECT 131.800 193.800 132.200 194.200 ;
        RECT 130.200 192.800 130.600 193.200 ;
        RECT 132.600 193.100 133.000 195.900 ;
        RECT 133.400 193.800 133.800 194.200 ;
        RECT 126.200 189.800 126.600 190.200 ;
        RECT 123.000 186.800 123.400 187.200 ;
        RECT 117.400 185.100 117.800 185.200 ;
        RECT 118.200 185.100 118.600 185.200 ;
        RECT 117.400 184.800 118.600 185.100 ;
        RECT 119.800 184.800 120.200 185.200 ;
        RECT 122.200 184.800 122.600 185.200 ;
        RECT 128.600 185.100 129.000 187.900 ;
        RECT 115.000 176.800 115.400 177.200 ;
        RECT 115.000 176.200 115.300 176.800 ;
        RECT 113.400 176.100 113.800 176.200 ;
        RECT 114.200 176.100 114.600 176.200 ;
        RECT 113.400 175.800 114.600 176.100 ;
        RECT 115.000 175.800 115.400 176.200 ;
        RECT 113.400 174.800 113.800 175.200 ;
        RECT 117.400 175.100 117.800 175.200 ;
        RECT 118.200 175.100 118.600 175.200 ;
        RECT 117.400 174.800 118.600 175.100 ;
        RECT 113.400 174.200 113.700 174.800 ;
        RECT 113.400 173.800 113.800 174.200 ;
        RECT 114.200 173.800 114.600 174.200 ;
        RECT 116.600 173.800 117.000 174.200 ;
        RECT 113.400 171.800 113.800 172.200 ;
        RECT 113.400 170.200 113.700 171.800 ;
        RECT 113.400 169.800 113.800 170.200 ;
        RECT 114.200 166.200 114.500 173.800 ;
        RECT 116.600 173.200 116.900 173.800 ;
        RECT 116.600 172.800 117.000 173.200 ;
        RECT 118.200 172.800 118.600 173.200 ;
        RECT 118.200 172.200 118.500 172.800 ;
        RECT 118.200 171.800 118.600 172.200 ;
        RECT 119.800 169.200 120.100 184.800 ;
        RECT 130.200 183.100 130.600 188.900 ;
        RECT 131.000 188.800 131.400 189.200 ;
        RECT 131.000 188.200 131.300 188.800 ;
        RECT 131.000 187.800 131.400 188.200 ;
        RECT 131.800 186.100 132.200 186.200 ;
        RECT 132.600 186.100 133.000 186.200 ;
        RECT 131.800 185.800 133.000 186.100 ;
        RECT 127.000 181.800 127.400 182.200 ;
        RECT 127.000 178.200 127.300 181.800 ;
        RECT 133.400 178.200 133.700 193.800 ;
        RECT 134.200 192.100 134.600 197.900 ;
        RECT 135.000 195.800 135.400 196.200 ;
        RECT 135.000 195.100 135.300 195.800 ;
        RECT 135.000 194.700 135.400 195.100 ;
        RECT 135.800 194.200 136.100 206.800 ;
        RECT 136.600 194.200 136.900 207.800 ;
        RECT 138.200 203.100 138.600 208.900 ;
        RECT 140.600 208.800 141.800 209.100 ;
        RECT 141.400 207.800 141.800 208.200 ;
        RECT 146.200 207.800 146.600 208.200 ;
        RECT 147.800 207.800 148.200 208.200 ;
        RECT 141.400 207.200 141.700 207.800 ;
        RECT 146.200 207.200 146.500 207.800 ;
        RECT 141.400 206.800 141.800 207.200 ;
        RECT 146.200 206.800 146.600 207.200 ;
        RECT 147.800 206.200 148.100 207.800 ;
        RECT 150.200 206.800 150.600 207.200 ;
        RECT 142.200 205.800 142.600 206.200 ;
        RECT 146.200 206.100 146.600 206.200 ;
        RECT 147.000 206.100 147.400 206.200 ;
        RECT 146.200 205.800 147.400 206.100 ;
        RECT 147.800 205.800 148.200 206.200 ;
        RECT 142.200 205.200 142.500 205.800 ;
        RECT 142.200 204.800 142.600 205.200 ;
        RECT 144.600 204.800 145.000 205.200 ;
        RECT 144.600 204.200 144.900 204.800 ;
        RECT 142.200 203.800 142.600 204.200 ;
        RECT 144.600 203.800 145.000 204.200 ;
        RECT 142.200 203.200 142.500 203.800 ;
        RECT 142.200 202.800 142.600 203.200 ;
        RECT 142.200 201.800 142.600 202.200 ;
        RECT 135.800 193.800 136.200 194.200 ;
        RECT 136.600 193.800 137.000 194.200 ;
        RECT 139.000 192.100 139.400 197.900 ;
        RECT 140.600 197.100 141.000 197.200 ;
        RECT 141.400 197.100 141.800 197.200 ;
        RECT 140.600 196.800 141.800 197.100 ;
        RECT 142.200 195.200 142.500 201.800 ;
        RECT 145.400 196.800 145.800 197.200 ;
        RECT 145.400 195.200 145.700 196.800 ;
        RECT 150.200 195.200 150.500 206.800 ;
        RECT 151.000 206.200 151.300 211.800 ;
        RECT 155.000 209.200 155.300 214.800 ;
        RECT 156.600 212.100 157.000 217.900 ;
        RECT 161.400 217.200 161.700 225.800 ;
        RECT 161.400 216.800 161.800 217.200 ;
        RECT 158.200 213.100 158.600 215.900 ;
        RECT 159.800 215.100 160.200 215.200 ;
        RECT 160.600 215.100 161.000 215.200 ;
        RECT 159.800 214.800 161.000 215.100 ;
        RECT 155.000 208.800 155.400 209.200 ;
        RECT 154.200 207.800 154.600 208.200 ;
        RECT 154.200 207.200 154.500 207.800 ;
        RECT 162.200 207.200 162.500 225.800 ;
        RECT 165.400 223.100 165.800 228.900 ;
        RECT 166.200 227.800 166.600 228.200 ;
        RECT 166.200 226.200 166.500 227.800 ;
        RECT 168.600 227.200 168.900 232.800 ;
        RECT 172.600 232.100 173.000 237.900 ;
        RECT 175.000 237.100 175.400 237.200 ;
        RECT 175.800 237.100 176.200 237.200 ;
        RECT 175.000 236.800 176.200 237.100 ;
        RECT 176.600 236.800 177.000 237.200 ;
        RECT 180.600 236.800 181.000 237.200 ;
        RECT 176.600 235.200 176.900 236.800 ;
        RECT 175.800 234.800 176.200 235.200 ;
        RECT 176.600 234.800 177.000 235.200 ;
        RECT 175.800 234.200 176.100 234.800 ;
        RECT 180.600 234.200 180.900 236.800 ;
        RECT 182.200 235.800 182.600 236.200 ;
        RECT 184.600 236.100 185.000 236.200 ;
        RECT 185.400 236.100 185.800 236.200 ;
        RECT 184.600 235.800 185.800 236.100 ;
        RECT 182.200 235.200 182.500 235.800 ;
        RECT 182.200 234.800 182.600 235.200 ;
        RECT 183.800 235.100 184.200 235.200 ;
        RECT 184.600 235.100 185.000 235.200 ;
        RECT 183.800 234.800 185.000 235.100 ;
        RECT 175.800 233.800 176.200 234.200 ;
        RECT 180.600 233.800 181.000 234.200 ;
        RECT 182.200 233.800 182.600 234.200 ;
        RECT 185.400 233.800 185.800 234.200 ;
        RECT 177.400 231.800 177.800 232.200 ;
        RECT 174.200 229.800 174.600 230.200 ;
        RECT 176.600 229.800 177.000 230.200 ;
        RECT 168.600 226.800 169.000 227.200 ;
        RECT 166.200 225.800 166.600 226.200 ;
        RECT 168.600 226.100 169.000 226.200 ;
        RECT 169.400 226.100 169.800 226.300 ;
        RECT 168.600 225.900 169.800 226.100 ;
        RECT 168.600 225.800 169.700 225.900 ;
        RECT 170.200 223.100 170.600 228.900 ;
        RECT 171.800 225.100 172.200 227.900 ;
        RECT 172.600 227.800 173.000 228.200 ;
        RECT 172.600 227.200 172.900 227.800 ;
        RECT 172.600 226.800 173.000 227.200 ;
        RECT 174.200 226.200 174.500 229.800 ;
        RECT 176.600 227.200 176.900 229.800 ;
        RECT 177.400 229.200 177.700 231.800 ;
        RECT 177.400 228.800 177.800 229.200 ;
        RECT 179.000 227.800 179.400 228.200 ;
        RECT 176.600 226.800 177.000 227.200 ;
        RECT 177.400 227.100 177.800 227.200 ;
        RECT 178.200 227.100 178.600 227.200 ;
        RECT 177.400 226.800 178.600 227.100 ;
        RECT 179.000 226.200 179.300 227.800 ;
        RECT 181.400 226.800 181.800 227.200 ;
        RECT 181.400 226.200 181.700 226.800 ;
        RECT 182.200 226.200 182.500 233.800 ;
        RECT 185.400 233.200 185.700 233.800 ;
        RECT 185.400 232.800 185.800 233.200 ;
        RECT 186.200 233.100 186.600 235.900 ;
        RECT 187.000 233.800 187.400 234.200 ;
        RECT 184.600 226.800 185.000 227.200 ;
        RECT 184.600 226.200 184.900 226.800 ;
        RECT 185.400 226.200 185.700 232.800 ;
        RECT 174.200 225.800 174.600 226.200 ;
        RECT 175.000 226.100 175.400 226.200 ;
        RECT 175.800 226.100 176.200 226.200 ;
        RECT 175.000 225.800 176.200 226.100 ;
        RECT 178.200 225.800 178.600 226.200 ;
        RECT 179.000 225.800 179.400 226.200 ;
        RECT 181.400 225.800 181.800 226.200 ;
        RECT 182.200 225.800 182.600 226.200 ;
        RECT 184.600 225.800 185.000 226.200 ;
        RECT 185.400 225.800 185.800 226.200 ;
        RECT 167.800 217.100 168.200 217.200 ;
        RECT 168.600 217.100 169.000 217.200 ;
        RECT 167.800 216.800 169.000 217.100 ;
        RECT 170.200 212.100 170.600 217.900 ;
        RECT 174.200 215.800 174.600 216.200 ;
        RECT 174.200 215.100 174.500 215.800 ;
        RECT 174.200 214.700 174.600 215.100 ;
        RECT 171.800 213.800 172.200 214.200 ;
        RECT 154.200 206.800 154.600 207.200 ;
        RECT 157.400 206.800 157.800 207.200 ;
        RECT 159.800 206.800 160.200 207.200 ;
        RECT 162.200 206.800 162.600 207.200 ;
        RECT 163.000 207.100 163.400 207.200 ;
        RECT 163.800 207.100 164.200 207.200 ;
        RECT 163.000 206.800 164.200 207.100 ;
        RECT 164.600 206.800 165.000 207.200 ;
        RECT 151.000 205.800 151.400 206.200 ;
        RECT 154.200 205.800 154.600 206.200 ;
        RECT 153.400 204.800 153.800 205.200 ;
        RECT 153.400 204.200 153.700 204.800 ;
        RECT 153.400 203.800 153.800 204.200 ;
        RECT 154.200 203.200 154.500 205.800 ;
        RECT 155.000 204.800 155.400 205.200 ;
        RECT 155.000 204.200 155.300 204.800 ;
        RECT 155.000 203.800 155.400 204.200 ;
        RECT 154.200 202.800 154.600 203.200 ;
        RECT 157.400 202.200 157.700 206.800 ;
        RECT 159.800 206.200 160.100 206.800 ;
        RECT 159.800 205.800 160.200 206.200 ;
        RECT 160.600 205.800 161.000 206.200 ;
        RECT 157.400 201.800 157.800 202.200 ;
        RECT 157.400 195.800 157.800 196.200 ;
        RECT 158.200 195.800 158.600 196.200 ;
        RECT 159.000 195.800 159.400 196.200 ;
        RECT 142.200 194.800 142.600 195.200 ;
        RECT 143.000 194.800 143.400 195.200 ;
        RECT 145.400 194.800 145.800 195.200 ;
        RECT 150.200 194.800 150.600 195.200 ;
        RECT 151.000 194.800 151.400 195.200 ;
        RECT 151.800 194.800 152.200 195.200 ;
        RECT 155.000 195.100 155.400 195.200 ;
        RECT 155.800 195.100 156.200 195.200 ;
        RECT 155.000 194.800 156.200 195.100 ;
        RECT 135.000 183.100 135.400 188.900 ;
        RECT 137.400 188.800 137.800 189.200 ;
        RECT 137.400 188.200 137.700 188.800 ;
        RECT 137.400 187.800 137.800 188.200 ;
        RECT 138.200 186.800 138.600 187.200 ;
        RECT 139.800 186.800 140.200 187.200 ;
        RECT 120.600 172.100 121.000 177.900 ;
        RECT 123.000 174.800 123.400 175.200 ;
        RECT 117.400 168.800 117.800 169.200 ;
        RECT 119.800 168.800 120.200 169.200 ;
        RECT 115.000 166.800 115.400 167.200 ;
        RECT 115.800 167.100 116.200 167.200 ;
        RECT 116.600 167.100 117.000 167.200 ;
        RECT 115.800 166.800 117.000 167.100 ;
        RECT 115.000 166.200 115.300 166.800 ;
        RECT 114.200 165.800 114.600 166.200 ;
        RECT 115.000 165.800 115.400 166.200 ;
        RECT 112.600 158.800 113.000 159.200 ;
        RECT 113.400 155.800 113.800 156.200 ;
        RECT 110.200 155.100 110.600 155.200 ;
        RECT 111.000 155.100 111.400 155.200 ;
        RECT 110.200 154.800 111.400 155.100 ;
        RECT 110.200 154.100 110.600 154.200 ;
        RECT 111.000 154.100 111.400 154.200 ;
        RECT 110.200 153.800 111.400 154.100 ;
        RECT 111.800 153.800 112.200 154.200 ;
        RECT 111.000 151.200 111.300 153.800 ;
        RECT 111.000 150.800 111.400 151.200 ;
        RECT 110.200 148.800 110.600 149.200 ;
        RECT 109.400 145.100 109.800 147.900 ;
        RECT 110.200 147.200 110.500 148.800 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 107.800 143.800 108.200 144.200 ;
        RECT 107.000 141.800 107.400 142.200 ;
        RECT 107.000 140.200 107.300 141.800 ;
        RECT 107.000 139.800 107.400 140.200 ;
        RECT 107.800 136.200 108.100 143.800 ;
        RECT 111.000 143.100 111.400 148.900 ;
        RECT 111.800 148.200 112.100 153.800 ;
        RECT 113.400 153.200 113.700 155.800 ;
        RECT 115.800 154.800 116.200 155.200 ;
        RECT 115.800 154.200 116.100 154.800 ;
        RECT 114.200 153.800 114.600 154.200 ;
        RECT 115.800 153.800 116.200 154.200 ;
        RECT 114.200 153.200 114.500 153.800 ;
        RECT 113.400 152.800 113.800 153.200 ;
        RECT 114.200 152.800 114.600 153.200 ;
        RECT 116.600 153.100 117.000 155.900 ;
        RECT 117.400 154.200 117.700 168.800 ;
        RECT 123.000 168.200 123.300 174.800 ;
        RECT 124.600 174.700 125.000 175.100 ;
        RECT 124.600 174.200 124.900 174.700 ;
        RECT 124.600 173.800 125.000 174.200 ;
        RECT 125.400 172.100 125.800 177.900 ;
        RECT 127.000 177.800 127.400 178.200 ;
        RECT 133.400 177.800 133.800 178.200 ;
        RECT 134.200 177.800 134.600 178.200 ;
        RECT 127.000 177.100 127.300 177.800 ;
        RECT 126.200 176.800 127.300 177.100 ;
        RECT 126.200 174.200 126.500 176.800 ;
        RECT 126.200 173.800 126.600 174.200 ;
        RECT 127.000 173.100 127.400 175.900 ;
        RECT 129.400 174.800 129.800 175.200 ;
        RECT 131.800 175.100 132.200 175.200 ;
        RECT 132.600 175.100 133.000 175.200 ;
        RECT 131.800 174.800 133.000 175.100 ;
        RECT 129.400 173.200 129.700 174.800 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 131.000 174.100 131.400 174.200 ;
        RECT 130.200 173.800 131.400 174.100 ;
        RECT 132.600 173.800 133.000 174.200 ;
        RECT 132.600 173.200 132.900 173.800 ;
        RECT 127.800 172.800 128.200 173.200 ;
        RECT 129.400 172.800 129.800 173.200 ;
        RECT 132.600 172.800 133.000 173.200 ;
        RECT 133.400 173.100 133.800 175.900 ;
        RECT 134.200 174.200 134.500 177.800 ;
        RECT 134.200 173.800 134.600 174.200 ;
        RECT 124.600 170.800 125.000 171.200 ;
        RECT 121.400 167.800 121.800 168.200 ;
        RECT 123.000 167.800 123.400 168.200 ;
        RECT 119.800 166.800 120.200 167.200 ;
        RECT 119.800 166.200 120.100 166.800 ;
        RECT 121.400 166.200 121.700 167.800 ;
        RECT 123.000 167.200 123.300 167.800 ;
        RECT 123.000 166.800 123.400 167.200 ;
        RECT 124.600 166.200 124.900 170.800 ;
        RECT 127.800 166.200 128.100 172.800 ;
        RECT 135.000 172.100 135.400 177.900 ;
        RECT 138.200 175.200 138.500 186.800 ;
        RECT 139.800 186.200 140.100 186.800 ;
        RECT 139.000 185.800 139.400 186.200 ;
        RECT 139.800 185.800 140.200 186.200 ;
        RECT 139.000 183.200 139.300 185.800 ;
        RECT 142.200 185.200 142.500 194.800 ;
        RECT 143.000 188.200 143.300 194.800 ;
        RECT 148.600 191.800 149.000 192.200 ;
        RECT 143.000 187.800 143.400 188.200 ;
        RECT 143.000 187.200 143.300 187.800 ;
        RECT 143.000 186.800 143.400 187.200 ;
        RECT 141.400 184.800 141.800 185.200 ;
        RECT 142.200 184.800 142.600 185.200 ;
        RECT 143.800 185.100 144.200 187.900 ;
        RECT 141.400 183.200 141.700 184.800 ;
        RECT 139.000 182.800 139.400 183.200 ;
        RECT 141.400 182.800 141.800 183.200 ;
        RECT 145.400 183.100 145.800 188.900 ;
        RECT 146.200 188.800 146.600 189.200 ;
        RECT 146.200 188.200 146.500 188.800 ;
        RECT 146.200 187.800 146.600 188.200 ;
        RECT 147.000 186.100 147.400 186.200 ;
        RECT 147.800 186.100 148.200 186.200 ;
        RECT 147.000 185.800 148.200 186.100 ;
        RECT 136.600 174.800 137.000 175.200 ;
        RECT 138.200 174.800 138.600 175.200 ;
        RECT 136.600 174.200 136.900 174.800 ;
        RECT 136.600 173.800 137.000 174.200 ;
        RECT 139.000 172.800 139.400 173.200 ;
        RECT 135.800 168.100 136.200 168.200 ;
        RECT 136.600 168.100 137.000 168.200 ;
        RECT 135.800 167.800 137.000 168.100 ;
        RECT 139.000 167.200 139.300 172.800 ;
        RECT 139.800 172.100 140.200 177.900 ;
        RECT 148.600 177.200 148.900 191.800 ;
        RECT 150.200 183.100 150.600 188.900 ;
        RECT 151.000 183.200 151.300 194.800 ;
        RECT 151.800 187.200 152.100 194.800 ;
        RECT 157.400 194.200 157.700 195.800 ;
        RECT 158.200 195.200 158.500 195.800 ;
        RECT 159.000 195.200 159.300 195.800 ;
        RECT 158.200 194.800 158.600 195.200 ;
        RECT 159.000 194.800 159.400 195.200 ;
        RECT 159.800 194.200 160.100 205.800 ;
        RECT 160.600 205.200 160.900 205.800 ;
        RECT 160.600 204.800 161.000 205.200 ;
        RECT 160.600 196.800 161.000 197.200 ;
        RECT 160.600 194.200 160.900 196.800 ;
        RECT 153.400 194.100 153.800 194.200 ;
        RECT 154.200 194.100 154.600 194.200 ;
        RECT 153.400 193.800 154.600 194.100 ;
        RECT 157.400 193.800 157.800 194.200 ;
        RECT 159.800 193.800 160.200 194.200 ;
        RECT 160.600 193.800 161.000 194.200 ;
        RECT 155.800 192.800 156.200 193.200 ;
        RECT 151.800 186.800 152.200 187.200 ;
        RECT 151.800 185.800 152.200 186.200 ;
        RECT 151.000 182.800 151.400 183.200 ;
        RECT 151.800 179.200 152.100 185.800 ;
        RECT 155.000 185.100 155.400 187.900 ;
        RECT 155.800 187.200 156.100 192.800 ;
        RECT 155.800 186.800 156.200 187.200 ;
        RECT 156.600 183.100 157.000 188.900 ;
        RECT 159.800 186.800 160.200 187.200 ;
        RECT 159.800 186.200 160.100 186.800 ;
        RECT 159.800 185.800 160.200 186.200 ;
        RECT 152.600 181.800 153.000 182.200 ;
        RECT 151.800 178.800 152.200 179.200 ;
        RECT 152.600 177.200 152.900 181.800 ;
        RECT 142.200 176.800 142.600 177.200 ;
        RECT 148.600 176.800 149.000 177.200 ;
        RECT 152.600 176.800 153.000 177.200 ;
        RECT 139.800 167.800 140.200 168.200 ;
        RECT 140.600 167.800 141.000 168.200 ;
        RECT 139.800 167.200 140.100 167.800 ;
        RECT 140.600 167.200 140.900 167.800 ;
        RECT 128.600 166.800 129.000 167.200 ;
        RECT 132.600 166.800 133.000 167.200 ;
        RECT 139.000 166.800 139.400 167.200 ;
        RECT 139.800 166.800 140.200 167.200 ;
        RECT 140.600 166.800 141.000 167.200 ;
        RECT 141.400 166.800 141.800 167.200 ;
        RECT 128.600 166.200 128.900 166.800 ;
        RECT 132.600 166.200 132.900 166.800 ;
        RECT 119.800 165.800 120.200 166.200 ;
        RECT 120.600 165.800 121.000 166.200 ;
        RECT 121.400 165.800 121.800 166.200 ;
        RECT 124.600 165.800 125.000 166.200 ;
        RECT 125.400 165.800 125.800 166.200 ;
        RECT 127.800 165.800 128.200 166.200 ;
        RECT 128.600 165.800 129.000 166.200 ;
        RECT 129.400 165.800 129.800 166.200 ;
        RECT 130.200 165.800 130.600 166.200 ;
        RECT 132.600 165.800 133.000 166.200 ;
        RECT 136.600 166.100 137.000 166.200 ;
        RECT 137.400 166.100 137.800 166.200 ;
        RECT 136.600 165.800 137.800 166.100 ;
        RECT 138.200 165.800 138.600 166.200 ;
        RECT 139.000 166.100 139.400 166.200 ;
        RECT 139.800 166.100 140.200 166.200 ;
        RECT 139.000 165.800 140.200 166.100 ;
        RECT 120.600 165.200 120.900 165.800 ;
        RECT 120.600 164.800 121.000 165.200 ;
        RECT 124.600 158.200 124.900 165.800 ;
        RECT 125.400 165.200 125.700 165.800 ;
        RECT 125.400 164.800 125.800 165.200 ;
        RECT 129.400 164.200 129.700 165.800 ;
        RECT 129.400 163.800 129.800 164.200 ;
        RECT 117.400 153.800 117.800 154.200 ;
        RECT 112.600 152.100 113.000 152.200 ;
        RECT 113.400 152.100 113.800 152.200 ;
        RECT 112.600 151.800 113.800 152.100 ;
        RECT 114.200 150.200 114.500 152.800 ;
        RECT 115.000 151.800 115.400 152.200 ;
        RECT 118.200 152.100 118.600 157.900 ;
        RECT 120.600 156.800 121.000 157.200 ;
        RECT 120.600 155.200 120.900 156.800 ;
        RECT 120.600 154.800 121.000 155.200 ;
        RECT 120.600 153.800 121.000 154.200 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 114.200 149.800 114.600 150.200 ;
        RECT 115.000 148.200 115.300 151.800 ;
        RECT 111.800 147.800 112.200 148.200 ;
        RECT 115.000 147.800 115.400 148.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 113.400 146.100 113.800 146.200 ;
        RECT 112.600 145.800 113.800 146.100 ;
        RECT 115.800 143.100 116.200 148.900 ;
        RECT 118.200 148.100 118.600 148.200 ;
        RECT 119.000 148.100 119.400 148.200 ;
        RECT 118.200 147.800 119.400 148.100 ;
        RECT 120.600 147.200 120.900 153.800 ;
        RECT 122.200 153.200 122.500 153.800 ;
        RECT 122.200 152.800 122.600 153.200 ;
        RECT 123.000 152.100 123.400 157.900 ;
        RECT 124.600 157.800 125.000 158.200 ;
        RECT 125.400 158.100 125.800 158.200 ;
        RECT 126.200 158.100 126.600 158.200 ;
        RECT 125.400 157.800 126.600 158.100 ;
        RECT 129.400 158.100 129.800 158.200 ;
        RECT 130.200 158.100 130.500 165.800 ;
        RECT 129.400 157.800 130.500 158.100 ;
        RECT 129.400 157.200 129.700 157.800 ;
        RECT 127.000 157.100 127.400 157.200 ;
        RECT 127.800 157.100 128.200 157.200 ;
        RECT 127.000 156.800 128.200 157.100 ;
        RECT 129.400 156.800 129.800 157.200 ;
        RECT 127.000 155.800 127.400 156.200 ;
        RECT 127.000 155.200 127.300 155.800 ;
        RECT 127.000 154.800 127.400 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 131.000 154.800 131.400 155.200 ;
        RECT 126.200 153.800 126.600 154.200 ;
        RECT 126.200 151.200 126.500 153.800 ;
        RECT 121.400 150.800 121.800 151.200 ;
        RECT 126.200 150.800 126.600 151.200 ;
        RECT 120.600 146.800 121.000 147.200 ;
        RECT 119.000 146.100 119.400 146.200 ;
        RECT 119.800 146.100 120.200 146.200 ;
        RECT 119.000 145.800 120.200 146.100 ;
        RECT 120.600 144.200 120.900 146.800 ;
        RECT 121.400 146.200 121.700 150.800 ;
        RECT 122.200 149.800 122.600 150.200 ;
        RECT 122.200 149.200 122.500 149.800 ;
        RECT 122.200 148.800 122.600 149.200 ;
        RECT 121.400 145.800 121.800 146.200 ;
        RECT 120.600 143.800 121.000 144.200 ;
        RECT 124.600 143.100 125.000 148.900 ;
        RECT 127.000 147.800 127.400 148.200 ;
        RECT 127.000 147.200 127.300 147.800 ;
        RECT 127.000 146.800 127.400 147.200 ;
        RECT 126.200 146.100 126.600 146.200 ;
        RECT 127.000 146.100 127.400 146.200 ;
        RECT 126.200 145.800 127.400 146.100 ;
        RECT 129.400 143.100 129.800 148.900 ;
        RECT 118.200 141.800 118.600 142.200 ;
        RECT 118.200 141.200 118.500 141.800 ;
        RECT 118.200 140.800 118.600 141.200 ;
        RECT 107.000 135.800 107.400 136.200 ;
        RECT 107.800 135.800 108.200 136.200 ;
        RECT 107.000 135.200 107.300 135.800 ;
        RECT 100.600 135.100 101.000 135.200 ;
        RECT 101.400 135.100 101.800 135.200 ;
        RECT 100.600 134.800 101.800 135.100 ;
        RECT 102.200 134.800 102.600 135.200 ;
        RECT 106.200 134.800 106.600 135.200 ;
        RECT 107.000 134.800 107.400 135.200 ;
        RECT 109.400 135.100 109.800 135.200 ;
        RECT 110.200 135.100 110.600 135.200 ;
        RECT 109.400 134.800 110.600 135.100 ;
        RECT 103.000 133.800 103.400 134.200 ;
        RECT 107.800 133.800 108.200 134.200 ;
        RECT 109.400 133.800 109.800 134.200 ;
        RECT 103.000 133.200 103.300 133.800 ;
        RECT 107.800 133.200 108.100 133.800 ;
        RECT 109.400 133.200 109.700 133.800 ;
        RECT 103.000 132.800 103.400 133.200 ;
        RECT 107.800 132.800 108.200 133.200 ;
        RECT 109.400 132.800 109.800 133.200 ;
        RECT 111.000 133.100 111.400 135.900 ;
        RECT 98.200 131.800 98.600 132.200 ;
        RECT 103.800 131.800 104.200 132.200 ;
        RECT 107.800 131.800 108.200 132.200 ;
        RECT 112.600 132.100 113.000 137.900 ;
        RECT 114.200 135.100 114.600 135.200 ;
        RECT 115.000 135.100 115.400 135.200 ;
        RECT 114.200 134.800 115.400 135.100 ;
        RECT 115.000 134.100 115.400 134.200 ;
        RECT 115.800 134.100 116.200 134.200 ;
        RECT 115.000 133.800 116.200 134.100 ;
        RECT 116.600 132.800 117.000 133.200 ;
        RECT 98.200 131.200 98.500 131.800 ;
        RECT 98.200 130.800 98.600 131.200 ;
        RECT 90.200 129.800 90.600 130.200 ;
        RECT 84.600 121.800 85.000 122.200 ;
        RECT 88.600 121.800 89.000 122.200 ;
        RECT 89.400 121.800 89.800 122.200 ;
        RECT 70.200 114.800 70.600 115.200 ;
        RECT 71.000 114.800 71.400 115.200 ;
        RECT 74.200 114.800 74.600 115.200 ;
        RECT 75.000 114.800 75.400 115.200 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 77.400 115.100 77.800 115.200 ;
        RECT 78.200 115.100 78.600 115.200 ;
        RECT 77.400 114.800 78.600 115.100 ;
        RECT 79.800 114.800 80.200 115.200 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 83.000 114.800 83.400 115.200 ;
        RECT 71.000 114.200 71.300 114.800 ;
        RECT 68.600 114.100 69.000 114.200 ;
        RECT 69.400 114.100 69.800 114.200 ;
        RECT 68.600 113.800 69.800 114.100 ;
        RECT 71.000 113.800 71.400 114.200 ;
        RECT 72.600 114.100 73.000 114.200 ;
        RECT 73.400 114.100 73.800 114.200 ;
        RECT 72.600 113.800 73.800 114.100 ;
        RECT 68.600 112.800 69.000 113.200 ;
        RECT 68.600 112.200 68.900 112.800 ;
        RECT 68.600 111.800 69.000 112.200 ;
        RECT 67.800 110.800 68.200 111.200 ;
        RECT 63.800 108.800 64.200 109.200 ;
        RECT 67.800 109.100 68.200 109.200 ;
        RECT 68.600 109.100 69.000 109.200 ;
        RECT 62.200 105.900 62.600 106.300 ;
        RECT 62.200 105.800 62.500 105.900 ;
        RECT 65.400 105.800 65.800 106.200 ;
        RECT 65.400 105.200 65.700 105.800 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 66.200 103.100 66.600 108.900 ;
        RECT 67.800 108.800 69.000 109.100 ;
        RECT 69.400 107.200 69.700 113.800 ;
        RECT 72.600 113.200 72.900 113.800 ;
        RECT 72.600 112.800 73.000 113.200 ;
        RECT 74.200 107.200 74.500 114.800 ;
        RECT 75.000 113.200 75.300 114.800 ;
        RECT 75.800 114.200 76.100 114.800 ;
        RECT 75.800 113.800 76.200 114.200 ;
        RECT 75.000 112.800 75.400 113.200 ;
        RECT 78.200 110.800 78.600 111.200 ;
        RECT 69.400 106.800 69.800 107.200 ;
        RECT 71.800 107.100 72.200 107.200 ;
        RECT 72.600 107.100 73.000 107.200 ;
        RECT 71.800 106.800 73.000 107.100 ;
        RECT 74.200 106.800 74.600 107.200 ;
        RECT 67.000 105.800 67.400 106.200 ;
        RECT 70.200 106.100 70.600 106.200 ;
        RECT 71.000 106.100 71.400 106.200 ;
        RECT 70.200 105.800 71.400 106.100 ;
        RECT 72.600 105.800 73.000 106.200 ;
        RECT 67.000 97.200 67.300 105.800 ;
        RECT 67.000 96.800 67.400 97.200 ;
        RECT 60.600 93.800 61.000 94.200 ;
        RECT 61.400 93.100 61.800 95.900 ;
        RECT 62.200 95.800 62.600 96.200 ;
        RECT 63.800 96.100 64.200 96.200 ;
        RECT 64.600 96.100 65.000 96.200 ;
        RECT 63.800 95.800 65.000 96.100 ;
        RECT 62.200 90.200 62.500 95.800 ;
        RECT 63.800 94.800 64.200 95.200 ;
        RECT 63.800 93.200 64.100 94.800 ;
        RECT 64.600 93.800 65.000 94.200 ;
        RECT 64.600 93.200 64.900 93.800 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 64.600 92.800 65.000 93.200 ;
        RECT 64.600 91.200 64.900 92.800 ;
        RECT 65.400 91.800 65.800 92.200 ;
        RECT 67.800 92.100 68.200 97.900 ;
        RECT 70.200 95.200 70.500 105.800 ;
        RECT 72.600 105.200 72.900 105.800 ;
        RECT 74.200 105.200 74.500 106.800 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 74.200 104.800 74.600 105.200 ;
        RECT 75.000 105.100 75.400 107.900 ;
        RECT 76.600 103.100 77.000 108.900 ;
        RECT 77.400 106.800 77.800 107.200 ;
        RECT 77.400 106.300 77.700 106.800 ;
        RECT 77.400 105.900 77.800 106.300 ;
        RECT 75.800 101.800 76.200 102.200 ;
        RECT 75.800 99.200 76.100 101.800 ;
        RECT 75.800 98.800 76.200 99.200 ;
        RECT 71.000 95.800 71.400 96.200 ;
        RECT 71.000 95.200 71.300 95.800 ;
        RECT 70.200 94.800 70.600 95.200 ;
        RECT 71.000 94.800 71.400 95.200 ;
        RECT 70.200 93.800 70.600 94.200 ;
        RECT 64.600 90.800 65.000 91.200 ;
        RECT 59.800 89.800 60.200 90.200 ;
        RECT 62.200 89.800 62.600 90.200 ;
        RECT 59.800 89.200 60.100 89.800 ;
        RECT 59.800 88.800 60.200 89.200 ;
        RECT 60.600 88.800 61.000 89.200 ;
        RECT 60.600 88.200 60.900 88.800 ;
        RECT 60.600 87.800 61.000 88.200 ;
        RECT 59.800 85.100 60.200 85.200 ;
        RECT 59.000 84.800 60.200 85.100 ;
        RECT 57.400 79.800 57.800 80.200 ;
        RECT 47.000 71.800 47.400 72.200 ;
        RECT 49.400 72.100 49.800 77.900 ;
        RECT 51.800 75.100 52.200 75.200 ;
        RECT 52.600 75.100 53.000 75.200 ;
        RECT 51.800 74.800 53.000 75.100 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 47.000 68.800 47.400 69.200 ;
        RECT 47.000 66.200 47.300 68.800 ;
        RECT 51.800 67.800 52.200 68.200 ;
        RECT 51.800 67.200 52.100 67.800 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 50.200 66.200 50.500 66.800 ;
        RECT 47.000 65.800 47.400 66.200 ;
        RECT 48.600 66.100 49.000 66.200 ;
        RECT 49.400 66.100 49.800 66.200 ;
        RECT 48.600 65.800 49.800 66.100 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 47.800 64.100 48.200 64.200 ;
        RECT 48.600 64.100 49.000 64.200 ;
        RECT 47.800 63.800 49.000 64.100 ;
        RECT 51.000 63.200 51.300 65.800 ;
        RECT 51.000 62.800 51.400 63.200 ;
        RECT 51.800 62.800 52.200 63.200 ;
        RECT 40.600 54.800 41.000 55.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 42.200 54.800 42.600 55.200 ;
        RECT 43.000 54.800 43.400 55.200 ;
        RECT 46.200 54.800 46.600 55.200 ;
        RECT 43.000 54.200 43.300 54.800 ;
        RECT 38.200 53.800 38.600 54.200 ;
        RECT 43.000 53.800 43.400 54.200 ;
        RECT 35.000 52.800 35.400 53.200 ;
        RECT 35.800 52.800 36.200 53.200 ;
        RECT 35.000 52.200 35.300 52.800 ;
        RECT 35.000 51.800 35.400 52.200 ;
        RECT 35.800 49.200 36.100 52.800 ;
        RECT 32.600 49.100 33.000 49.200 ;
        RECT 33.400 49.100 33.800 49.200 ;
        RECT 32.600 48.800 33.800 49.100 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 27.800 46.200 28.100 46.800 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 31.000 45.800 31.400 46.200 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 31.800 45.800 33.000 46.100 ;
        RECT 31.000 45.200 31.300 45.800 ;
        RECT 31.000 44.800 31.400 45.200 ;
        RECT 27.800 35.800 28.200 36.200 ;
        RECT 29.400 36.100 29.800 36.200 ;
        RECT 30.200 36.100 30.600 36.200 ;
        RECT 29.400 35.800 30.600 36.100 ;
        RECT 27.800 35.200 28.100 35.800 ;
        RECT 25.400 34.800 25.800 35.200 ;
        RECT 27.000 34.800 27.400 35.200 ;
        RECT 27.800 34.800 28.200 35.200 ;
        RECT 25.400 32.200 25.700 34.800 ;
        RECT 27.000 33.800 27.400 34.200 ;
        RECT 27.000 33.200 27.300 33.800 ;
        RECT 27.000 32.800 27.400 33.200 ;
        RECT 31.000 32.200 31.300 44.800 ;
        RECT 35.000 43.100 35.400 48.900 ;
        RECT 35.800 48.800 36.200 49.200 ;
        RECT 38.200 46.200 38.500 53.800 ;
        RECT 47.000 53.100 47.400 55.900 ;
        RECT 40.600 51.800 41.000 52.200 ;
        RECT 48.600 52.100 49.000 57.900 ;
        RECT 51.000 55.800 51.400 56.200 ;
        RECT 51.000 55.200 51.300 55.800 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 50.200 53.800 50.600 54.200 ;
        RECT 39.000 48.800 39.400 49.200 ;
        RECT 39.000 48.200 39.300 48.800 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 35.800 45.800 36.200 46.200 ;
        RECT 38.200 45.800 38.600 46.200 ;
        RECT 35.800 36.200 36.100 45.800 ;
        RECT 39.800 43.100 40.200 48.900 ;
        RECT 38.200 41.800 38.600 42.200 ;
        RECT 35.800 35.800 36.200 36.200 ;
        RECT 35.800 35.200 36.100 35.800 ;
        RECT 38.200 35.200 38.500 41.800 ;
        RECT 40.600 39.200 40.900 51.800 ;
        RECT 42.200 49.100 42.600 49.200 ;
        RECT 43.000 49.100 43.400 49.200 ;
        RECT 42.200 48.800 43.400 49.100 ;
        RECT 41.400 45.100 41.800 47.900 ;
        RECT 44.600 43.100 45.000 48.900 ;
        RECT 48.600 46.800 49.000 47.200 ;
        RECT 48.600 46.300 48.900 46.800 ;
        RECT 48.600 45.900 49.000 46.300 ;
        RECT 49.400 43.100 49.800 48.900 ;
        RECT 50.200 47.200 50.500 53.800 ;
        RECT 51.800 49.200 52.100 62.800 ;
        RECT 51.800 48.800 52.200 49.200 ;
        RECT 50.200 46.800 50.600 47.200 ;
        RECT 40.600 38.800 41.000 39.200 ;
        RECT 33.400 35.100 33.800 35.200 ;
        RECT 34.200 35.100 34.600 35.200 ;
        RECT 33.400 34.800 34.600 35.100 ;
        RECT 35.800 34.800 36.200 35.200 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 39.000 34.800 39.400 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 41.400 35.100 41.800 35.200 ;
        RECT 40.600 34.800 41.800 35.100 ;
        RECT 42.200 34.800 42.600 35.200 ;
        RECT 37.400 34.200 37.700 34.800 ;
        RECT 38.200 34.200 38.500 34.800 ;
        RECT 31.800 33.800 32.200 34.200 ;
        RECT 32.600 33.800 33.000 34.200 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 38.200 33.800 38.600 34.200 ;
        RECT 25.400 31.800 25.800 32.200 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 31.000 31.800 31.400 32.200 ;
        RECT 26.200 30.800 26.600 31.200 ;
        RECT 20.600 28.800 21.000 29.200 ;
        RECT 24.600 28.800 25.000 29.200 ;
        RECT 26.200 26.200 26.500 30.800 ;
        RECT 27.800 28.800 28.200 29.200 ;
        RECT 29.400 29.100 29.700 31.800 ;
        RECT 31.800 29.200 32.100 33.800 ;
        RECT 32.600 33.200 32.900 33.800 ;
        RECT 32.600 32.800 33.000 33.200 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 17.400 25.800 17.800 26.200 ;
        RECT 18.200 25.800 18.600 26.200 ;
        RECT 20.600 25.800 21.000 26.200 ;
        RECT 21.400 25.800 21.800 26.200 ;
        RECT 24.600 26.100 25.000 26.200 ;
        RECT 25.400 26.100 25.800 26.200 ;
        RECT 24.600 25.800 25.800 26.100 ;
        RECT 26.200 25.800 26.600 26.200 ;
        RECT 18.200 19.200 18.500 25.800 ;
        RECT 18.200 18.800 18.600 19.200 ;
        RECT 19.000 16.800 19.400 17.200 ;
        RECT 14.200 15.800 14.600 16.200 ;
        RECT 16.600 16.100 17.000 16.200 ;
        RECT 17.400 16.100 17.800 16.200 ;
        RECT 16.600 15.800 17.800 16.100 ;
        RECT 14.200 15.200 14.500 15.800 ;
        RECT 19.000 15.200 19.300 16.800 ;
        RECT 14.200 14.800 14.600 15.200 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 19.800 14.800 20.200 15.200 ;
        RECT 18.200 14.200 18.500 14.800 ;
        RECT 19.800 14.200 20.100 14.800 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 18.200 13.800 18.600 14.200 ;
        RECT 19.000 13.800 19.400 14.200 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 13.400 13.200 13.700 13.800 ;
        RECT 12.600 12.800 13.000 13.200 ;
        RECT 13.400 12.800 13.800 13.200 ;
        RECT 6.200 8.800 6.600 9.200 ;
        RECT 8.600 8.800 9.000 9.200 ;
        RECT 7.800 7.100 8.200 7.200 ;
        RECT 8.600 7.100 9.000 7.200 ;
        RECT 7.800 6.800 9.000 7.100 ;
        RECT 9.400 5.800 9.800 6.200 ;
        RECT 9.400 5.200 9.700 5.800 ;
        RECT 9.400 4.800 9.800 5.200 ;
        RECT 10.200 5.100 10.600 7.900 ;
        RECT 11.800 3.100 12.200 8.900 ;
        RECT 12.600 8.200 12.900 12.800 ;
        RECT 12.600 7.800 13.000 8.200 ;
        RECT 15.000 6.200 15.300 13.800 ;
        RECT 19.000 9.200 19.300 13.800 ;
        RECT 20.600 9.200 20.900 25.800 ;
        RECT 21.400 19.200 21.700 25.800 ;
        RECT 27.000 25.100 27.400 27.900 ;
        RECT 21.400 18.800 21.800 19.200 ;
        RECT 23.800 13.800 24.200 14.200 ;
        RECT 23.800 12.200 24.100 13.800 ;
        RECT 23.800 11.800 24.200 12.200 ;
        RECT 26.200 12.100 26.600 17.900 ;
        RECT 15.000 5.800 15.400 6.200 ;
        RECT 16.600 3.100 17.000 8.900 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 19.800 9.100 20.200 9.200 ;
        RECT 20.600 9.100 21.000 9.200 ;
        RECT 19.800 8.800 21.000 9.100 ;
        RECT 22.200 3.100 22.600 8.900 ;
        RECT 25.400 6.800 25.800 7.200 ;
        RECT 25.400 6.200 25.700 6.800 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 27.000 3.100 27.400 8.900 ;
        RECT 27.800 7.200 28.100 28.800 ;
        RECT 28.600 23.100 29.000 28.900 ;
        RECT 29.400 28.800 30.500 29.100 ;
        RECT 31.800 28.800 32.200 29.200 ;
        RECT 29.400 27.800 29.800 28.200 ;
        RECT 29.400 27.200 29.700 27.800 ;
        RECT 29.400 26.800 29.800 27.200 ;
        RECT 29.400 14.200 29.700 26.800 ;
        RECT 30.200 26.200 30.500 28.800 ;
        RECT 32.600 28.200 32.900 32.800 ;
        RECT 34.200 31.800 34.600 32.200 ;
        RECT 35.000 31.800 35.400 32.200 ;
        RECT 32.600 27.800 33.000 28.200 ;
        RECT 30.200 25.800 30.600 26.200 ;
        RECT 33.400 23.100 33.800 28.900 ;
        RECT 30.200 14.700 30.600 15.100 ;
        RECT 29.400 13.800 29.800 14.200 ;
        RECT 30.200 12.200 30.500 14.700 ;
        RECT 30.200 11.800 30.600 12.200 ;
        RECT 31.000 12.100 31.400 17.900 ;
        RECT 32.600 13.100 33.000 15.900 ;
        RECT 33.400 13.800 33.800 14.200 ;
        RECT 33.400 13.200 33.700 13.800 ;
        RECT 33.400 12.800 33.800 13.200 ;
        RECT 29.400 8.800 29.800 9.200 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 27.800 5.200 28.100 6.800 ;
        RECT 27.800 4.800 28.200 5.200 ;
        RECT 28.600 5.100 29.000 7.900 ;
        RECT 29.400 7.200 29.700 8.800 ;
        RECT 34.200 7.200 34.500 31.800 ;
        RECT 35.000 26.200 35.300 31.800 ;
        RECT 39.000 30.200 39.300 34.800 ;
        RECT 41.400 30.200 41.700 34.800 ;
        RECT 35.800 29.800 36.200 30.200 ;
        RECT 39.000 29.800 39.400 30.200 ;
        RECT 41.400 29.800 41.800 30.200 ;
        RECT 35.800 29.200 36.100 29.800 ;
        RECT 42.200 29.200 42.500 34.800 ;
        RECT 44.600 32.800 45.000 33.200 ;
        RECT 45.400 33.100 45.800 35.900 ;
        RECT 44.600 32.200 44.900 32.800 ;
        RECT 43.800 31.800 44.200 32.200 ;
        RECT 44.600 31.800 45.000 32.200 ;
        RECT 47.000 32.100 47.400 37.900 ;
        RECT 50.200 35.200 50.500 46.800 ;
        RECT 51.000 45.100 51.400 47.900 ;
        RECT 51.800 47.200 52.100 48.800 ;
        RECT 52.600 48.200 52.900 73.800 ;
        RECT 54.200 72.100 54.600 77.900 ;
        RECT 55.800 73.100 56.200 75.900 ;
        RECT 57.400 74.200 57.700 79.800 ;
        RECT 59.800 77.200 60.100 84.800 ;
        RECT 63.000 83.100 63.400 88.900 ;
        RECT 65.400 86.200 65.700 91.800 ;
        RECT 63.800 85.800 64.200 86.200 ;
        RECT 65.400 85.800 65.800 86.200 ;
        RECT 67.000 85.900 67.400 86.300 ;
        RECT 63.800 80.200 64.100 85.800 ;
        RECT 67.000 85.200 67.300 85.900 ;
        RECT 67.000 84.800 67.400 85.200 ;
        RECT 67.800 83.100 68.200 88.900 ;
        RECT 69.400 85.100 69.800 87.900 ;
        RECT 70.200 85.200 70.500 93.800 ;
        RECT 72.600 92.100 73.000 97.900 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 73.400 94.200 73.700 94.800 ;
        RECT 73.400 93.800 73.800 94.200 ;
        RECT 74.200 93.100 74.600 95.900 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 75.000 94.200 75.300 94.800 ;
        RECT 75.000 93.800 75.400 94.200 ;
        RECT 75.000 92.800 75.400 93.200 ;
        RECT 75.000 91.200 75.300 92.800 ;
        RECT 78.200 92.200 78.500 110.800 ;
        RECT 79.800 100.200 80.100 114.800 ;
        RECT 82.200 113.800 82.600 114.200 ;
        RECT 82.200 113.200 82.500 113.800 ;
        RECT 82.200 112.800 82.600 113.200 ;
        RECT 83.000 111.200 83.300 114.800 ;
        RECT 84.600 114.200 84.900 121.800 ;
        RECT 85.400 119.800 85.800 120.200 ;
        RECT 85.400 119.200 85.700 119.800 ;
        RECT 85.400 118.800 85.800 119.200 ;
        RECT 86.200 116.800 86.600 117.200 ;
        RECT 87.800 116.800 88.200 117.200 ;
        RECT 85.400 115.800 85.800 116.200 ;
        RECT 85.400 115.200 85.700 115.800 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 84.600 114.100 85.000 114.200 ;
        RECT 83.800 113.800 85.000 114.100 ;
        RECT 83.000 110.800 83.400 111.200 ;
        RECT 80.600 105.800 81.000 106.200 ;
        RECT 79.800 99.800 80.200 100.200 ;
        RECT 78.200 91.800 78.600 92.200 ;
        RECT 75.000 90.800 75.400 91.200 ;
        RECT 71.800 87.800 72.200 88.200 ;
        RECT 71.800 87.200 72.100 87.800 ;
        RECT 75.000 87.200 75.300 90.800 ;
        RECT 76.600 88.800 77.000 89.200 ;
        RECT 76.600 87.200 76.900 88.800 ;
        RECT 78.200 87.200 78.500 91.800 ;
        RECT 79.000 89.800 79.400 90.200 ;
        RECT 71.800 86.800 72.200 87.200 ;
        RECT 72.600 86.800 73.000 87.200 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 76.600 86.800 77.000 87.200 ;
        RECT 78.200 86.800 78.600 87.200 ;
        RECT 72.600 86.200 72.900 86.800 ;
        RECT 72.600 85.800 73.000 86.200 ;
        RECT 74.200 85.800 74.600 86.200 ;
        RECT 74.200 85.200 74.500 85.800 ;
        RECT 70.200 84.800 70.600 85.200 ;
        RECT 74.200 84.800 74.600 85.200 ;
        RECT 63.800 79.800 64.200 80.200 ;
        RECT 63.800 78.200 64.100 79.800 ;
        RECT 59.800 76.800 60.200 77.200 ;
        RECT 57.400 73.800 57.800 74.200 ;
        RECT 56.600 71.800 57.000 72.200 ;
        RECT 58.200 72.100 58.600 72.200 ;
        RECT 59.000 72.100 59.400 72.200 ;
        RECT 60.600 72.100 61.000 77.900 ;
        RECT 63.800 77.800 64.200 78.200 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 63.800 73.200 64.100 74.800 ;
        RECT 63.800 72.800 64.200 73.200 ;
        RECT 65.400 72.100 65.800 77.900 ;
        RECT 69.400 76.800 69.800 77.200 ;
        RECT 71.800 76.800 72.200 77.200 ;
        RECT 69.400 76.200 69.700 76.800 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 66.200 74.200 66.500 74.800 ;
        RECT 66.200 73.800 66.600 74.200 ;
        RECT 67.000 73.100 67.400 75.900 ;
        RECT 69.400 75.800 69.800 76.200 ;
        RECT 71.800 75.200 72.100 76.800 ;
        RECT 73.400 75.800 73.800 76.200 ;
        RECT 73.400 75.200 73.700 75.800 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 74.200 75.100 74.600 75.200 ;
        RECT 75.000 75.100 75.300 86.800 ;
        RECT 79.000 86.200 79.300 89.800 ;
        RECT 80.600 89.200 80.900 105.800 ;
        RECT 81.400 103.100 81.800 108.900 ;
        RECT 83.800 107.200 84.100 113.800 ;
        RECT 84.600 110.800 85.000 111.200 ;
        RECT 84.600 108.200 84.900 110.800 ;
        RECT 84.600 107.800 85.000 108.200 ;
        RECT 83.800 106.800 84.200 107.200 ;
        RECT 85.400 106.200 85.700 114.800 ;
        RECT 86.200 106.200 86.500 116.800 ;
        RECT 87.800 116.200 88.100 116.800 ;
        RECT 87.800 115.800 88.200 116.200 ;
        RECT 88.600 115.200 88.900 121.800 ;
        RECT 89.400 120.800 89.800 121.200 ;
        RECT 88.600 114.800 89.000 115.200 ;
        RECT 89.400 114.200 89.700 120.800 ;
        RECT 90.200 116.200 90.500 129.800 ;
        RECT 92.600 127.800 93.000 128.200 ;
        RECT 91.800 121.800 92.200 122.200 ;
        RECT 91.800 121.200 92.100 121.800 ;
        RECT 91.800 120.800 92.200 121.200 ;
        RECT 92.600 119.200 92.900 127.800 ;
        RECT 94.200 123.100 94.600 128.900 ;
        RECT 98.200 128.200 98.500 130.800 ;
        RECT 103.800 130.200 104.100 131.800 ;
        RECT 103.800 129.800 104.200 130.200 ;
        RECT 98.200 127.800 98.600 128.200 ;
        RECT 97.400 125.800 97.800 126.200 ;
        RECT 97.400 120.200 97.700 125.800 ;
        RECT 99.000 123.100 99.400 128.900 ;
        RECT 101.400 128.800 101.800 129.200 ;
        RECT 103.000 129.100 103.400 129.200 ;
        RECT 103.800 129.100 104.200 129.200 ;
        RECT 103.000 128.800 104.200 129.100 ;
        RECT 100.600 125.100 101.000 127.900 ;
        RECT 101.400 126.200 101.700 128.800 ;
        RECT 103.800 127.100 104.200 127.200 ;
        RECT 104.600 127.100 105.000 127.200 ;
        RECT 103.800 126.800 105.000 127.100 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 107.800 125.200 108.100 131.800 ;
        RECT 110.200 130.800 110.600 131.200 ;
        RECT 109.400 129.800 109.800 130.200 ;
        RECT 109.400 126.200 109.700 129.800 ;
        RECT 109.400 125.800 109.800 126.200 ;
        RECT 104.600 125.100 105.000 125.200 ;
        RECT 105.400 125.100 105.800 125.200 ;
        RECT 104.600 124.800 105.800 125.100 ;
        RECT 107.800 124.800 108.200 125.200 ;
        RECT 108.600 125.100 109.000 125.200 ;
        RECT 109.400 125.100 109.800 125.200 ;
        RECT 108.600 124.800 109.800 125.100 ;
        RECT 110.200 124.200 110.500 130.800 ;
        RECT 115.000 127.800 115.400 128.200 ;
        RECT 115.000 127.200 115.300 127.800 ;
        RECT 116.600 127.200 116.900 132.800 ;
        RECT 117.400 132.100 117.800 137.900 ;
        RECT 121.400 135.800 121.800 136.200 ;
        RECT 123.800 136.100 124.200 136.200 ;
        RECT 124.600 136.100 125.000 136.200 ;
        RECT 123.800 135.800 125.000 136.100 ;
        RECT 121.400 135.200 121.700 135.800 ;
        RECT 121.400 134.800 121.800 135.200 ;
        RECT 122.200 135.100 122.600 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 122.200 134.800 123.400 135.100 ;
        RECT 125.400 134.800 125.800 135.200 ;
        RECT 125.400 134.200 125.700 134.800 ;
        RECT 120.600 133.800 121.000 134.200 ;
        RECT 121.400 133.800 121.800 134.200 ;
        RECT 125.400 133.800 125.800 134.200 ;
        RECT 126.200 133.800 126.600 134.200 ;
        RECT 128.600 133.800 129.000 134.200 ;
        RECT 119.800 132.800 120.200 133.200 ;
        RECT 119.800 132.200 120.100 132.800 ;
        RECT 119.800 131.800 120.200 132.200 ;
        RECT 120.600 131.200 120.900 133.800 ;
        RECT 120.600 130.800 121.000 131.200 ;
        RECT 119.800 129.800 120.200 130.200 ;
        RECT 119.800 127.200 120.100 129.800 ;
        RECT 121.400 127.200 121.700 133.800 ;
        RECT 125.400 133.200 125.700 133.800 ;
        RECT 126.200 133.200 126.500 133.800 ;
        RECT 125.400 132.800 125.800 133.200 ;
        RECT 126.200 132.800 126.600 133.200 ;
        RECT 127.800 131.800 128.200 132.200 ;
        RECT 125.400 130.800 125.800 131.200 ;
        RECT 111.000 127.100 111.400 127.200 ;
        RECT 111.800 127.100 112.200 127.200 ;
        RECT 111.000 126.800 112.200 127.100 ;
        RECT 115.000 126.800 115.400 127.200 ;
        RECT 116.600 127.100 117.000 127.200 ;
        RECT 117.400 127.100 117.800 127.200 ;
        RECT 116.600 126.800 117.800 127.100 ;
        RECT 119.800 126.800 120.200 127.200 ;
        RECT 121.400 126.800 121.800 127.200 ;
        RECT 119.800 126.200 120.100 126.800 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 114.200 125.800 114.600 126.200 ;
        RECT 117.400 126.100 117.800 126.200 ;
        RECT 118.200 126.100 118.600 126.200 ;
        RECT 117.400 125.800 118.600 126.100 ;
        RECT 119.800 125.800 120.200 126.200 ;
        RECT 113.400 125.200 113.700 125.800 ;
        RECT 113.400 124.800 113.800 125.200 ;
        RECT 109.400 123.800 109.800 124.200 ;
        RECT 110.200 123.800 110.600 124.200 ;
        RECT 109.400 123.200 109.700 123.800 ;
        RECT 109.400 122.800 109.800 123.200 ;
        RECT 103.000 121.800 103.400 122.200 ;
        RECT 97.400 119.800 97.800 120.200 ;
        RECT 92.600 118.800 93.000 119.200 ;
        RECT 90.200 115.800 90.600 116.200 ;
        RECT 90.200 115.200 90.500 115.800 ;
        RECT 90.200 114.800 90.600 115.200 ;
        RECT 91.000 114.800 91.400 115.200 ;
        RECT 92.600 115.100 93.000 115.200 ;
        RECT 93.400 115.100 93.800 115.200 ;
        RECT 92.600 114.800 93.800 115.100 ;
        RECT 91.000 114.200 91.300 114.800 ;
        RECT 89.400 113.800 89.800 114.200 ;
        RECT 91.000 113.800 91.400 114.200 ;
        RECT 91.000 112.800 91.400 113.200 ;
        RECT 88.600 106.800 89.000 107.200 ;
        RECT 89.400 106.800 89.800 107.200 ;
        RECT 85.400 105.800 85.800 106.200 ;
        RECT 86.200 105.800 86.600 106.200 ;
        RECT 87.000 106.100 87.400 106.200 ;
        RECT 87.800 106.100 88.200 106.200 ;
        RECT 87.000 105.800 88.200 106.100 ;
        RECT 86.200 105.200 86.500 105.800 ;
        RECT 88.600 105.200 88.900 106.800 ;
        RECT 89.400 106.200 89.700 106.800 ;
        RECT 89.400 105.800 89.800 106.200 ;
        RECT 83.800 104.800 84.200 105.200 ;
        RECT 86.200 104.800 86.600 105.200 ;
        RECT 88.600 104.800 89.000 105.200 ;
        RECT 90.200 105.100 90.600 107.900 ;
        RECT 83.800 104.200 84.100 104.800 ;
        RECT 83.800 103.800 84.200 104.200 ;
        RECT 82.200 96.800 82.600 97.200 ;
        RECT 82.200 95.200 82.500 96.800 ;
        RECT 82.200 94.800 82.600 95.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 87.800 94.800 88.200 95.200 ;
        RECT 81.400 94.100 81.800 94.200 ;
        RECT 82.200 94.100 82.600 94.200 ;
        RECT 81.400 93.800 82.600 94.100 ;
        RECT 80.600 88.800 81.000 89.200 ;
        RECT 75.800 86.100 76.200 86.200 ;
        RECT 76.600 86.100 77.000 86.200 ;
        RECT 75.800 85.800 77.000 86.100 ;
        RECT 79.000 85.800 79.400 86.200 ;
        RECT 79.800 85.800 80.200 86.200 ;
        RECT 76.600 83.200 76.900 85.800 ;
        RECT 76.600 82.800 77.000 83.200 ;
        RECT 79.000 82.800 79.400 83.200 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 76.600 80.200 76.900 81.800 ;
        RECT 76.600 79.800 77.000 80.200 ;
        RECT 74.200 74.800 75.300 75.100 ;
        RECT 77.400 74.800 77.800 75.200 ;
        RECT 77.400 74.200 77.700 74.800 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 72.600 73.800 73.000 74.200 ;
        RECT 77.400 73.800 77.800 74.200 ;
        RECT 67.800 72.200 68.100 73.800 ;
        RECT 70.200 73.100 70.600 73.200 ;
        RECT 71.000 73.100 71.400 73.200 ;
        RECT 70.200 72.800 71.400 73.100 ;
        RECT 58.200 71.800 59.400 72.100 ;
        RECT 67.800 71.800 68.200 72.200 ;
        RECT 53.400 69.800 53.800 70.200 ;
        RECT 53.400 69.200 53.700 69.800 ;
        RECT 53.400 68.800 53.800 69.200 ;
        RECT 54.200 68.800 54.600 69.200 ;
        RECT 54.200 67.200 54.500 68.800 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 56.600 66.200 56.900 71.800 ;
        RECT 58.200 69.100 58.600 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 58.200 68.800 59.400 69.100 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 69.400 67.100 69.800 67.200 ;
        RECT 70.200 67.100 70.600 67.200 ;
        RECT 69.400 66.800 70.600 67.100 ;
        RECT 64.600 66.200 64.900 66.800 ;
        RECT 65.400 66.200 65.700 66.800 ;
        RECT 66.200 66.200 66.500 66.800 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 57.400 66.100 57.800 66.200 ;
        RECT 58.200 66.100 58.600 66.200 ;
        RECT 57.400 65.800 58.600 66.100 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 67.000 65.800 67.400 66.200 ;
        RECT 69.400 65.800 69.800 66.200 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 71.800 65.800 72.200 66.200 ;
        RECT 54.200 65.200 54.500 65.800 ;
        RECT 54.200 64.800 54.600 65.200 ;
        RECT 62.200 63.200 62.500 65.800 ;
        RECT 67.000 65.100 67.300 65.800 ;
        RECT 66.200 64.800 67.300 65.100 ;
        RECT 62.200 62.800 62.600 63.200 ;
        RECT 66.200 59.200 66.500 64.800 ;
        RECT 66.200 58.800 66.600 59.200 ;
        RECT 69.400 58.200 69.700 65.800 ;
        RECT 71.800 64.200 72.100 65.800 ;
        RECT 71.800 63.800 72.200 64.200 ;
        RECT 53.400 52.100 53.800 57.900 ;
        RECT 57.400 57.800 57.800 58.200 ;
        RECT 69.400 57.800 69.800 58.200 ;
        RECT 57.400 55.200 57.700 57.800 ;
        RECT 69.400 56.800 69.800 57.200 ;
        RECT 59.800 56.100 60.200 56.200 ;
        RECT 60.600 56.100 61.000 56.200 ;
        RECT 59.800 55.800 61.000 56.100 ;
        RECT 67.800 55.800 68.200 56.200 ;
        RECT 67.800 55.200 68.100 55.800 ;
        RECT 69.400 55.200 69.700 56.800 ;
        RECT 57.400 54.800 57.800 55.200 ;
        RECT 63.000 54.800 63.400 55.200 ;
        RECT 63.800 54.800 64.200 55.200 ;
        RECT 67.000 54.800 67.400 55.200 ;
        RECT 67.800 54.800 68.200 55.200 ;
        RECT 69.400 54.800 69.800 55.200 ;
        RECT 71.800 54.800 72.200 55.200 ;
        RECT 55.800 52.800 56.200 53.200 ;
        RECT 55.800 52.200 56.100 52.800 ;
        RECT 55.800 51.800 56.200 52.200 ;
        RECT 57.400 51.200 57.700 54.800 ;
        RECT 63.000 54.200 63.300 54.800 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 58.200 53.800 59.400 54.100 ;
        RECT 63.000 53.800 63.400 54.200 ;
        RECT 63.800 53.200 64.100 54.800 ;
        RECT 67.000 54.200 67.300 54.800 ;
        RECT 71.800 54.200 72.100 54.800 ;
        RECT 67.000 53.800 67.400 54.200 ;
        RECT 68.600 53.800 69.000 54.200 ;
        RECT 71.800 53.800 72.200 54.200 ;
        RECT 61.400 53.100 61.800 53.200 ;
        RECT 62.200 53.100 62.600 53.200 ;
        RECT 61.400 52.800 62.600 53.100 ;
        RECT 63.800 52.800 64.200 53.200 ;
        RECT 57.400 50.800 57.800 51.200 ;
        RECT 59.800 50.800 60.200 51.200 ;
        RECT 59.800 49.200 60.100 50.800 ;
        RECT 67.000 49.200 67.300 53.800 ;
        RECT 68.600 51.200 68.900 53.800 ;
        RECT 71.000 51.800 71.400 52.200 ;
        RECT 68.600 50.800 69.000 51.200 ;
        RECT 71.000 49.200 71.300 51.800 ;
        RECT 71.800 49.800 72.200 50.200 ;
        RECT 71.800 49.200 72.100 49.800 ;
        RECT 59.800 48.800 60.200 49.200 ;
        RECT 62.200 49.100 62.600 49.200 ;
        RECT 63.000 49.100 63.400 49.200 ;
        RECT 62.200 48.800 63.400 49.100 ;
        RECT 52.600 47.800 53.000 48.200 ;
        RECT 51.800 46.800 52.200 47.200 ;
        RECT 53.400 47.100 53.800 47.200 ;
        RECT 54.200 47.100 54.600 47.200 ;
        RECT 53.400 46.800 54.600 47.100 ;
        RECT 57.400 46.800 57.800 47.200 ;
        RECT 58.200 46.800 58.600 47.200 ;
        RECT 57.400 46.200 57.700 46.800 ;
        RECT 53.400 45.800 53.800 46.200 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 53.400 45.200 53.700 45.800 ;
        RECT 58.200 45.200 58.500 46.800 ;
        RECT 61.400 45.800 61.800 46.200 ;
        RECT 61.400 45.200 61.700 45.800 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 58.200 44.800 58.600 45.200 ;
        RECT 61.400 44.800 61.800 45.200 ;
        RECT 64.600 43.100 65.000 48.900 ;
        RECT 67.000 48.800 67.400 49.200 ;
        RECT 68.600 48.800 69.000 49.200 ;
        RECT 68.600 46.300 68.900 48.800 ;
        RECT 68.600 45.900 69.000 46.300 ;
        RECT 69.400 43.100 69.800 48.900 ;
        RECT 71.000 48.800 71.400 49.200 ;
        RECT 71.800 48.800 72.200 49.200 ;
        RECT 70.200 46.800 70.600 47.200 ;
        RECT 66.200 38.800 66.600 39.200 ;
        RECT 66.200 38.200 66.500 38.800 ;
        RECT 47.800 34.700 48.200 35.100 ;
        RECT 50.200 34.800 50.600 35.200 ;
        RECT 43.800 29.200 44.100 31.800 ;
        RECT 47.800 31.100 48.100 34.700 ;
        RECT 47.000 30.800 48.100 31.100 ;
        RECT 45.400 29.800 45.800 30.200 ;
        RECT 45.400 29.200 45.700 29.800 ;
        RECT 47.000 29.200 47.300 30.800 ;
        RECT 35.800 28.800 36.200 29.200 ;
        RECT 37.400 28.800 37.800 29.200 ;
        RECT 35.000 25.800 35.400 26.200 ;
        RECT 36.600 25.100 37.000 27.900 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 35.000 14.200 35.300 14.800 ;
        RECT 37.400 14.200 37.700 28.800 ;
        RECT 38.200 23.100 38.600 28.900 ;
        RECT 42.200 28.800 42.600 29.200 ;
        RECT 42.200 27.200 42.500 28.800 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 42.200 26.800 42.600 27.200 ;
        RECT 39.000 26.300 39.300 26.800 ;
        RECT 39.000 25.900 39.400 26.300 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 42.200 23.200 42.500 25.800 ;
        RECT 42.200 22.800 42.600 23.200 ;
        RECT 43.000 23.100 43.400 28.900 ;
        RECT 43.800 28.800 44.200 29.200 ;
        RECT 45.400 28.800 45.800 29.200 ;
        RECT 46.200 28.800 46.600 29.200 ;
        RECT 47.000 28.800 47.400 29.200 ;
        RECT 46.200 28.200 46.500 28.800 ;
        RECT 46.200 27.800 46.600 28.200 ;
        RECT 47.800 27.800 48.200 28.200 ;
        RECT 48.600 27.800 49.000 28.200 ;
        RECT 47.800 26.200 48.100 27.800 ;
        RECT 48.600 27.200 48.900 27.800 ;
        RECT 48.600 26.800 49.000 27.200 ;
        RECT 47.800 26.100 48.200 26.200 ;
        RECT 48.600 26.100 49.000 26.200 ;
        RECT 47.800 25.800 49.000 26.100 ;
        RECT 47.800 24.800 48.200 25.200 ;
        RECT 49.400 25.100 49.800 27.900 ;
        RECT 50.200 27.200 50.500 34.800 ;
        RECT 51.800 32.100 52.200 37.900 ;
        RECT 66.200 37.800 66.600 38.200 ;
        RECT 69.400 37.800 69.800 38.200 ;
        RECT 62.200 35.800 62.600 36.200 ;
        RECT 63.000 36.100 63.400 36.200 ;
        RECT 63.800 36.100 64.200 36.200 ;
        RECT 63.000 35.800 64.200 36.100 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 61.400 35.100 61.800 35.200 ;
        RECT 60.600 34.800 61.800 35.100 ;
        RECT 59.800 33.200 60.100 34.800 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 61.400 33.200 61.700 33.800 ;
        RECT 59.800 32.800 60.200 33.200 ;
        RECT 61.400 32.800 61.800 33.200 ;
        RECT 53.400 32.100 53.800 32.200 ;
        RECT 54.200 32.100 54.600 32.200 ;
        RECT 53.400 31.800 54.600 32.100 ;
        RECT 58.200 32.100 58.600 32.200 ;
        RECT 59.000 32.100 59.400 32.200 ;
        RECT 58.200 31.800 59.400 32.100 ;
        RECT 59.800 29.200 60.100 32.800 ;
        RECT 50.200 26.800 50.600 27.200 ;
        RECT 50.200 25.200 50.500 26.800 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 47.800 19.200 48.100 24.800 ;
        RECT 50.200 22.800 50.600 23.200 ;
        RECT 51.000 23.100 51.400 28.900 ;
        RECT 52.600 25.800 53.000 26.200 ;
        RECT 52.600 25.200 52.900 25.800 ;
        RECT 52.600 24.800 53.000 25.200 ;
        RECT 55.800 23.100 56.200 28.900 ;
        RECT 59.800 28.800 60.200 29.200 ;
        RECT 60.600 27.100 61.000 27.200 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 60.600 26.800 61.800 27.100 ;
        RECT 60.600 26.200 60.900 26.800 ;
        RECT 60.600 25.800 61.000 26.200 ;
        RECT 61.400 26.100 61.800 26.200 ;
        RECT 62.200 26.100 62.500 35.800 ;
        RECT 69.400 35.200 69.700 37.800 ;
        RECT 63.000 35.100 63.400 35.200 ;
        RECT 63.800 35.100 64.200 35.200 ;
        RECT 63.000 34.800 64.200 35.100 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 67.800 34.800 68.200 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 63.800 33.800 64.200 34.200 ;
        RECT 61.400 25.800 62.500 26.100 ;
        RECT 47.800 18.800 48.200 19.200 ;
        RECT 41.400 17.800 41.800 18.200 ;
        RECT 41.400 15.200 41.700 17.800 ;
        RECT 38.200 14.800 38.600 15.200 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 35.000 13.800 35.400 14.200 ;
        RECT 37.400 13.800 37.800 14.200 ;
        RECT 36.600 12.100 37.000 12.200 ;
        RECT 37.400 12.100 37.800 12.200 ;
        RECT 36.600 11.800 37.800 12.100 ;
        RECT 38.200 9.200 38.500 14.800 ;
        RECT 39.800 13.800 40.200 14.200 ;
        RECT 42.200 14.100 42.600 14.200 ;
        RECT 41.400 13.800 42.600 14.100 ;
        RECT 39.800 13.200 40.100 13.800 ;
        RECT 39.800 12.800 40.200 13.200 ;
        RECT 38.200 8.800 38.600 9.200 ;
        RECT 38.200 7.200 38.500 8.800 ;
        RECT 41.400 7.200 41.700 13.800 ;
        RECT 50.200 12.200 50.500 22.800 ;
        RECT 51.800 18.100 52.200 18.200 ;
        RECT 52.600 18.100 53.000 18.200 ;
        RECT 51.800 17.800 53.000 18.100 ;
        RECT 57.400 17.800 57.800 18.200 ;
        RECT 57.400 15.200 57.700 17.800 ;
        RECT 57.400 14.800 57.800 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 59.000 15.100 59.400 15.200 ;
        RECT 58.200 14.800 59.400 15.100 ;
        RECT 60.600 14.200 60.900 25.800 ;
        RECT 61.400 24.800 61.800 25.200 ;
        RECT 61.400 24.200 61.700 24.800 ;
        RECT 61.400 23.800 61.800 24.200 ;
        RECT 62.200 16.200 62.500 25.800 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 63.000 25.200 63.300 31.800 ;
        RECT 63.800 26.200 64.100 33.800 ;
        RECT 64.600 32.200 64.900 34.800 ;
        RECT 64.600 31.800 65.000 32.200 ;
        RECT 65.400 27.100 65.800 27.200 ;
        RECT 66.200 27.100 66.600 27.200 ;
        RECT 65.400 26.800 66.600 27.100 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 63.000 24.800 63.400 25.200 ;
        RECT 63.800 21.200 64.100 25.800 ;
        RECT 67.000 22.200 67.300 34.800 ;
        RECT 67.800 26.200 68.100 34.800 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 69.400 34.100 69.800 34.200 ;
        RECT 68.600 33.800 69.800 34.100 ;
        RECT 70.200 32.200 70.500 46.800 ;
        RECT 71.000 45.100 71.400 47.900 ;
        RECT 72.600 47.200 72.900 73.800 ;
        RECT 76.600 72.800 77.000 73.200 ;
        RECT 76.600 68.200 76.900 72.800 ;
        RECT 76.600 67.800 77.000 68.200 ;
        RECT 76.600 67.200 76.900 67.800 ;
        RECT 76.600 66.800 77.000 67.200 ;
        RECT 77.400 67.100 77.800 67.200 ;
        RECT 78.200 67.100 78.600 67.200 ;
        RECT 77.400 66.800 78.600 67.100 ;
        RECT 79.000 66.200 79.300 82.800 ;
        RECT 79.800 79.200 80.100 85.800 ;
        RECT 79.800 78.800 80.200 79.200 ;
        RECT 80.600 77.800 81.000 78.200 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 73.400 65.800 74.600 66.100 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 79.000 65.200 79.300 65.800 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 79.800 65.100 80.200 67.900 ;
        RECT 80.600 67.200 80.900 77.800 ;
        RECT 81.400 74.200 81.700 93.800 ;
        RECT 83.000 93.100 83.300 94.800 ;
        RECT 82.200 92.800 83.300 93.100 ;
        RECT 87.800 93.200 88.100 94.800 ;
        RECT 87.800 92.800 88.200 93.200 ;
        RECT 82.200 89.200 82.500 92.800 ;
        RECT 83.800 91.800 84.200 92.200 ;
        RECT 83.800 90.200 84.100 91.800 ;
        RECT 83.800 89.800 84.200 90.200 ;
        RECT 82.200 88.800 82.600 89.200 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 83.000 86.200 83.300 88.800 ;
        RECT 83.800 86.800 84.200 87.200 ;
        RECT 83.800 86.200 84.100 86.800 ;
        RECT 83.000 85.800 83.400 86.200 ;
        RECT 83.800 85.800 84.200 86.200 ;
        RECT 88.600 84.200 88.900 104.800 ;
        RECT 91.000 103.200 91.300 112.800 ;
        RECT 95.000 111.800 95.400 112.200 ;
        RECT 97.400 112.100 97.800 117.900 ;
        RECT 101.400 114.700 101.800 115.100 ;
        RECT 101.400 114.200 101.700 114.700 ;
        RECT 101.400 113.800 101.800 114.200 ;
        RECT 102.200 112.100 102.600 117.900 ;
        RECT 103.000 116.200 103.300 121.800 ;
        RECT 108.600 120.800 109.000 121.200 ;
        RECT 103.000 115.800 103.400 116.200 ;
        RECT 103.800 113.100 104.200 115.900 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 95.000 109.200 95.300 111.800 ;
        RECT 99.000 110.800 99.400 111.200 ;
        RECT 99.000 109.200 99.300 110.800 ;
        RECT 104.600 109.200 104.900 114.800 ;
        RECT 106.200 113.100 106.600 115.900 ;
        RECT 107.800 112.100 108.200 117.900 ;
        RECT 91.000 102.800 91.400 103.200 ;
        RECT 91.800 103.100 92.200 108.900 ;
        RECT 95.000 108.800 95.400 109.200 ;
        RECT 92.600 106.800 93.000 107.200 ;
        RECT 90.200 97.800 90.600 98.200 ;
        RECT 90.200 95.200 90.500 97.800 ;
        RECT 91.000 95.200 91.300 102.800 ;
        RECT 92.600 102.200 92.900 106.800 ;
        RECT 93.400 105.800 93.800 106.200 ;
        RECT 93.400 105.200 93.700 105.800 ;
        RECT 93.400 104.800 93.800 105.200 ;
        RECT 92.600 101.800 93.000 102.200 ;
        RECT 95.000 98.200 95.300 108.800 ;
        RECT 96.600 103.100 97.000 108.900 ;
        RECT 99.000 108.800 99.400 109.200 ;
        RECT 104.600 108.800 105.000 109.200 ;
        RECT 106.200 108.800 106.600 109.200 ;
        RECT 106.200 108.200 106.500 108.800 ;
        RECT 103.800 107.800 104.200 108.200 ;
        RECT 106.200 107.800 106.600 108.200 ;
        RECT 103.800 107.200 104.100 107.800 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 103.800 106.800 104.200 107.200 ;
        RECT 99.800 106.200 100.100 106.800 ;
        RECT 99.800 105.800 100.200 106.200 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 103.000 105.800 103.400 106.200 ;
        RECT 102.200 105.200 102.500 105.800 ;
        RECT 102.200 104.800 102.600 105.200 ;
        RECT 99.000 99.800 99.400 100.200 ;
        RECT 95.000 97.800 95.400 98.200 ;
        RECT 91.800 95.800 92.200 96.200 ;
        RECT 91.800 95.200 92.100 95.800 ;
        RECT 90.200 94.800 90.600 95.200 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 92.600 94.800 93.000 95.200 ;
        RECT 95.800 94.800 96.200 95.200 ;
        RECT 90.200 93.800 90.600 94.200 ;
        RECT 90.200 89.200 90.500 93.800 ;
        RECT 92.600 91.200 92.900 94.800 ;
        RECT 95.800 94.200 96.100 94.800 ;
        RECT 95.800 93.800 96.200 94.200 ;
        RECT 97.400 93.800 97.800 94.200 ;
        RECT 97.400 93.200 97.700 93.800 ;
        RECT 97.400 92.800 97.800 93.200 ;
        RECT 92.600 90.800 93.000 91.200 ;
        RECT 98.200 90.800 98.600 91.200 ;
        RECT 90.200 88.800 90.600 89.200 ;
        RECT 91.800 88.800 92.200 89.200 ;
        RECT 92.600 89.100 93.000 89.200 ;
        RECT 93.400 89.100 93.800 89.200 ;
        RECT 92.600 88.800 93.800 89.100 ;
        RECT 91.800 88.200 92.100 88.800 ;
        RECT 91.800 87.800 92.200 88.200 ;
        RECT 91.800 85.100 92.200 85.200 ;
        RECT 92.600 85.100 93.000 85.200 ;
        RECT 91.800 84.800 93.000 85.100 ;
        RECT 88.600 83.800 89.000 84.200 ;
        RECT 91.800 83.800 92.200 84.200 ;
        RECT 91.800 79.200 92.100 83.800 ;
        RECT 95.800 83.100 96.200 88.900 ;
        RECT 98.200 79.200 98.500 90.800 ;
        RECT 99.000 87.200 99.300 99.800 ;
        RECT 100.600 92.100 101.000 97.900 ;
        RECT 101.400 93.800 101.800 94.200 ;
        RECT 99.800 87.800 100.200 88.200 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 99.800 86.300 100.100 87.800 ;
        RECT 99.800 85.900 100.200 86.300 ;
        RECT 100.600 83.100 101.000 88.900 ;
        RECT 91.800 78.800 92.200 79.200 ;
        RECT 98.200 78.800 98.600 79.200 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 82.200 72.100 82.600 77.900 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 85.400 75.100 85.800 75.200 ;
        RECT 84.600 74.800 85.800 75.100 ;
        RECT 87.000 72.100 87.400 77.900 ;
        RECT 94.200 77.800 94.600 78.200 ;
        RECT 89.400 76.800 89.800 77.200 ;
        RECT 93.400 76.800 93.800 77.200 ;
        RECT 89.400 76.200 89.700 76.800 ;
        RECT 87.800 74.800 88.200 75.200 ;
        RECT 87.800 74.200 88.100 74.800 ;
        RECT 87.800 73.800 88.200 74.200 ;
        RECT 88.600 73.100 89.000 75.900 ;
        RECT 89.400 75.800 89.800 76.200 ;
        RECT 91.000 76.100 91.400 76.200 ;
        RECT 91.800 76.100 92.200 76.200 ;
        RECT 91.000 75.800 92.200 76.100 ;
        RECT 93.400 75.200 93.700 76.800 ;
        RECT 94.200 76.200 94.500 77.800 ;
        RECT 94.200 75.800 94.600 76.200 ;
        RECT 95.000 76.100 95.400 76.200 ;
        RECT 95.800 76.100 96.200 76.200 ;
        RECT 95.000 75.800 96.200 76.100 ;
        RECT 96.600 75.800 97.000 76.200 ;
        RECT 94.200 75.200 94.500 75.800 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 94.200 74.800 94.600 75.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 89.400 73.200 89.700 73.800 ;
        RECT 89.400 72.800 89.800 73.200 ;
        RECT 91.800 71.800 92.200 72.200 ;
        RECT 91.800 70.200 92.100 71.800 ;
        RECT 91.800 69.800 92.200 70.200 ;
        RECT 88.600 69.100 89.000 69.200 ;
        RECT 89.400 69.100 89.800 69.200 ;
        RECT 80.600 66.800 81.000 67.200 ;
        RECT 78.200 63.800 78.600 64.200 ;
        RECT 78.200 63.200 78.500 63.800 ;
        RECT 78.200 62.800 78.600 63.200 ;
        RECT 81.400 63.100 81.800 68.900 ;
        RECT 83.000 67.800 83.400 68.200 ;
        RECT 83.000 66.200 83.300 67.800 ;
        RECT 83.000 65.800 83.400 66.200 ;
        RECT 86.200 63.100 86.600 68.900 ;
        RECT 88.600 68.800 89.800 69.100 ;
        RECT 91.000 68.100 91.400 68.200 ;
        RECT 91.800 68.100 92.200 68.200 ;
        RECT 91.000 67.800 92.200 68.100 ;
        RECT 89.400 66.800 89.800 67.200 ;
        RECT 89.400 66.200 89.700 66.800 ;
        RECT 93.400 66.200 93.700 74.800 ;
        RECT 95.000 73.800 95.400 74.200 ;
        RECT 95.000 71.200 95.300 73.800 ;
        RECT 95.000 70.800 95.400 71.200 ;
        RECT 96.600 69.200 96.900 75.800 ;
        RECT 101.400 75.200 101.700 93.800 ;
        RECT 103.000 91.200 103.300 105.800 ;
        RECT 103.800 104.200 104.100 106.800 ;
        RECT 103.800 103.800 104.200 104.200 ;
        RECT 103.800 94.800 104.200 95.200 ;
        RECT 103.800 94.200 104.100 94.800 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 105.400 92.100 105.800 97.900 ;
        RECT 106.200 93.800 106.600 94.200 ;
        RECT 106.200 93.200 106.500 93.800 ;
        RECT 106.200 92.800 106.600 93.200 ;
        RECT 107.000 93.100 107.400 95.900 ;
        RECT 108.600 95.200 108.900 120.800 ;
        RECT 109.400 113.800 109.800 114.200 ;
        RECT 109.400 111.200 109.700 113.800 ;
        RECT 110.200 113.200 110.500 123.800 ;
        RECT 114.200 123.200 114.500 125.800 ;
        RECT 115.000 125.100 115.400 125.200 ;
        RECT 115.800 125.100 116.200 125.200 ;
        RECT 115.000 124.800 116.200 125.100 ;
        RECT 118.200 124.800 118.600 125.200 ;
        RECT 119.800 125.100 120.200 125.200 ;
        RECT 120.600 125.100 121.000 125.200 ;
        RECT 119.800 124.800 121.000 125.100 ;
        RECT 118.200 124.200 118.500 124.800 ;
        RECT 118.200 123.800 118.600 124.200 ;
        RECT 119.000 123.800 119.400 124.200 ;
        RECT 119.000 123.200 119.300 123.800 ;
        RECT 114.200 122.800 114.600 123.200 ;
        RECT 119.000 122.800 119.400 123.200 ;
        RECT 112.600 122.100 113.000 122.200 ;
        RECT 113.400 122.100 113.800 122.200 ;
        RECT 112.600 121.800 113.800 122.100 ;
        RECT 111.000 114.800 111.400 115.200 ;
        RECT 110.200 112.800 110.600 113.200 ;
        RECT 109.400 110.800 109.800 111.200 ;
        RECT 111.000 109.200 111.300 114.800 ;
        RECT 112.600 112.100 113.000 117.900 ;
        RECT 115.800 113.100 116.200 115.900 ;
        RECT 116.600 113.800 117.000 114.200 ;
        RECT 115.000 111.800 115.400 112.200 ;
        RECT 111.000 108.800 111.400 109.200 ;
        RECT 111.800 109.100 112.200 109.200 ;
        RECT 112.600 109.100 113.000 109.200 ;
        RECT 111.800 108.800 113.000 109.100 ;
        RECT 110.200 107.800 110.600 108.200 ;
        RECT 110.200 106.200 110.500 107.800 ;
        RECT 115.000 107.100 115.300 111.800 ;
        RECT 115.800 107.800 116.200 108.200 ;
        RECT 115.800 107.200 116.100 107.800 ;
        RECT 115.800 107.100 116.200 107.200 ;
        RECT 115.000 106.800 116.200 107.100 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 110.200 105.800 110.600 106.200 ;
        RECT 111.000 106.100 111.400 106.200 ;
        RECT 111.800 106.100 112.200 106.200 ;
        RECT 111.000 105.800 112.200 106.100 ;
        RECT 109.400 104.200 109.700 105.800 ;
        RECT 109.400 103.800 109.800 104.200 ;
        RECT 108.600 94.800 109.000 95.200 ;
        RECT 110.200 95.100 110.600 95.200 ;
        RECT 111.000 95.100 111.300 105.800 ;
        RECT 115.000 96.800 115.400 97.200 ;
        RECT 110.200 94.800 111.300 95.100 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 103.000 90.800 103.400 91.200 ;
        RECT 104.600 88.100 105.000 88.200 ;
        RECT 105.400 88.100 105.800 88.200 ;
        RECT 102.200 85.100 102.600 87.900 ;
        RECT 104.600 87.800 105.800 88.100 ;
        RECT 103.000 86.800 103.400 87.200 ;
        RECT 103.000 86.200 103.300 86.800 ;
        RECT 103.000 85.800 103.400 86.200 ;
        RECT 103.800 85.800 104.200 86.200 ;
        RECT 106.200 85.800 106.600 86.200 ;
        RECT 100.600 74.800 101.000 75.200 ;
        RECT 101.400 74.800 101.800 75.200 ;
        RECT 100.600 73.200 100.900 74.800 ;
        RECT 103.800 74.200 104.100 85.800 ;
        RECT 106.200 85.200 106.500 85.800 ;
        RECT 106.200 84.800 106.600 85.200 ;
        RECT 108.600 81.200 108.900 94.800 ;
        RECT 113.400 94.200 113.700 94.800 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 115.000 93.200 115.300 96.800 ;
        RECT 115.000 92.800 115.400 93.200 ;
        RECT 115.800 93.100 116.200 95.900 ;
        RECT 115.000 89.800 115.400 90.200 ;
        RECT 109.400 85.100 109.800 87.900 ;
        RECT 110.200 86.800 110.600 87.200 ;
        RECT 108.600 80.800 109.000 81.200 ;
        RECT 110.200 79.200 110.500 86.800 ;
        RECT 111.000 83.100 111.400 88.900 ;
        RECT 112.600 86.800 113.000 87.200 ;
        RECT 112.600 86.200 112.900 86.800 ;
        RECT 112.600 85.800 113.000 86.200 ;
        RECT 110.200 78.800 110.600 79.200 ;
        RECT 108.600 75.800 109.000 76.200 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 106.200 74.800 106.600 75.200 ;
        RECT 101.400 73.800 101.800 74.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 100.600 72.800 101.000 73.200 ;
        RECT 95.000 68.800 95.400 69.200 ;
        RECT 96.600 68.800 97.000 69.200 ;
        RECT 95.000 68.200 95.300 68.800 ;
        RECT 95.000 67.800 95.400 68.200 ;
        RECT 98.200 67.800 98.600 68.200 ;
        RECT 98.200 67.200 98.500 67.800 ;
        RECT 95.000 67.100 95.400 67.200 ;
        RECT 94.200 66.800 95.400 67.100 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 89.400 65.800 89.800 66.200 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 93.400 65.800 93.800 66.200 ;
        RECT 90.200 65.200 90.500 65.800 ;
        RECT 90.200 64.800 90.600 65.200 ;
        RECT 91.800 63.800 92.200 64.200 ;
        RECT 91.800 59.200 92.100 63.800 ;
        RECT 94.200 59.200 94.500 66.800 ;
        RECT 95.000 66.100 95.400 66.200 ;
        RECT 95.800 66.100 96.200 66.200 ;
        RECT 95.000 65.800 96.200 66.100 ;
        RECT 100.600 65.800 101.000 66.200 ;
        RECT 96.600 64.800 97.000 65.200 ;
        RECT 96.600 59.200 96.900 64.800 ;
        RECT 100.600 64.200 100.900 65.800 ;
        RECT 100.600 63.800 101.000 64.200 ;
        RECT 91.800 58.800 92.200 59.200 ;
        RECT 94.200 58.800 94.600 59.200 ;
        RECT 96.600 58.800 97.000 59.200 ;
        RECT 73.400 56.800 73.800 57.200 ;
        RECT 74.200 57.100 74.600 57.200 ;
        RECT 75.000 57.100 75.400 57.200 ;
        RECT 74.200 56.800 75.400 57.100 ;
        RECT 73.400 56.200 73.700 56.800 ;
        RECT 73.400 55.800 73.800 56.200 ;
        RECT 76.600 52.100 77.000 57.900 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 79.800 54.800 81.000 55.100 ;
        RECT 80.600 54.700 81.000 54.800 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 72.600 46.800 73.000 47.200 ;
        RECT 74.200 43.100 74.600 48.900 ;
        RECT 78.200 45.900 78.600 46.300 ;
        RECT 78.200 45.200 78.500 45.900 ;
        RECT 78.200 44.800 78.600 45.200 ;
        RECT 79.000 43.100 79.400 48.900 ;
        RECT 79.800 48.200 80.100 53.800 ;
        RECT 81.400 52.100 81.800 57.900 ;
        RECT 83.800 57.800 84.200 58.200 ;
        RECT 88.600 57.800 89.000 58.200 ;
        RECT 83.000 53.100 83.400 55.900 ;
        RECT 83.800 55.200 84.100 57.800 ;
        RECT 87.000 56.800 87.400 57.200 ;
        RECT 83.800 54.800 84.200 55.200 ;
        RECT 84.600 55.100 85.000 55.200 ;
        RECT 85.400 55.100 85.800 55.200 ;
        RECT 84.600 54.800 85.800 55.100 ;
        RECT 87.000 54.200 87.300 56.800 ;
        RECT 88.600 56.200 88.900 57.800 ;
        RECT 90.200 56.800 90.600 57.200 ;
        RECT 88.600 55.800 89.000 56.200 ;
        RECT 90.200 55.200 90.500 56.800 ;
        RECT 94.200 55.800 94.600 56.200 ;
        RECT 94.200 55.200 94.500 55.800 ;
        RECT 88.600 55.100 89.000 55.200 ;
        RECT 89.400 55.100 89.800 55.200 ;
        RECT 88.600 54.800 89.800 55.100 ;
        RECT 90.200 54.800 90.600 55.200 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 95.000 54.800 95.400 55.200 ;
        RECT 98.200 54.800 98.600 55.200 ;
        RECT 92.600 54.200 92.900 54.800 ;
        RECT 83.800 53.800 84.200 54.200 ;
        RECT 86.200 53.800 86.600 54.200 ;
        RECT 87.000 53.800 87.400 54.200 ;
        RECT 92.600 53.800 93.000 54.200 ;
        RECT 79.800 47.800 80.200 48.200 ;
        RECT 79.800 47.200 80.100 47.800 ;
        RECT 79.800 46.800 80.200 47.200 ;
        RECT 80.600 45.100 81.000 47.900 ;
        RECT 83.800 47.200 84.100 53.800 ;
        RECT 86.200 49.200 86.500 53.800 ;
        RECT 91.000 51.800 91.400 52.200 ;
        RECT 86.200 48.800 86.600 49.200 ;
        RECT 86.200 47.200 86.500 48.800 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 82.200 47.100 82.600 47.200 ;
        RECT 81.400 46.800 82.600 47.100 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 86.200 46.800 86.600 47.200 ;
        RECT 71.800 37.800 72.200 38.200 ;
        RECT 71.800 36.200 72.100 37.800 ;
        RECT 73.400 36.800 73.800 37.200 ;
        RECT 71.800 35.800 72.200 36.200 ;
        RECT 71.800 34.800 72.200 35.200 ;
        RECT 71.800 34.200 72.100 34.800 ;
        RECT 73.400 34.200 73.700 36.800 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 73.400 33.800 73.800 34.200 ;
        RECT 74.200 33.100 74.600 35.900 ;
        RECT 70.200 31.800 70.600 32.200 ;
        RECT 75.800 32.100 76.200 37.900 ;
        RECT 76.600 35.800 77.000 36.200 ;
        RECT 79.800 35.800 80.200 36.200 ;
        RECT 76.600 35.100 76.900 35.800 ;
        RECT 79.800 35.200 80.100 35.800 ;
        RECT 76.600 34.700 77.000 35.100 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 78.200 33.800 78.600 34.200 ;
        RECT 72.600 29.100 73.000 29.200 ;
        RECT 73.400 29.100 73.800 29.200 ;
        RECT 72.600 28.800 73.800 29.100 ;
        RECT 71.800 26.800 72.200 27.200 ;
        RECT 71.800 26.200 72.100 26.800 ;
        RECT 67.800 25.800 68.200 26.200 ;
        RECT 71.800 25.800 72.200 26.200 ;
        RECT 67.800 25.200 68.100 25.800 ;
        RECT 67.800 24.800 68.200 25.200 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 70.200 25.100 70.600 25.200 ;
        RECT 69.400 24.800 70.600 25.100 ;
        RECT 75.000 23.100 75.400 28.900 ;
        RECT 78.200 27.200 78.500 33.800 ;
        RECT 80.600 32.100 81.000 37.900 ;
        RECT 81.400 34.200 81.700 46.800 ;
        RECT 82.200 46.100 82.600 46.200 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 82.200 45.800 83.400 46.100 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 84.600 45.200 84.900 45.800 ;
        RECT 82.200 44.800 82.600 45.200 ;
        RECT 84.600 45.100 85.000 45.200 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 87.000 45.100 87.400 47.900 ;
        RECT 87.800 47.800 88.200 48.200 ;
        RECT 87.800 47.200 88.100 47.800 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 84.600 44.800 85.800 45.100 ;
        RECT 82.200 44.200 82.500 44.800 ;
        RECT 82.200 43.800 82.600 44.200 ;
        RECT 83.800 40.800 84.200 41.200 ;
        RECT 82.200 37.100 82.600 37.200 ;
        RECT 83.000 37.100 83.400 37.200 ;
        RECT 82.200 36.800 83.400 37.100 ;
        RECT 83.800 35.200 84.100 40.800 ;
        RECT 86.200 39.800 86.600 40.200 ;
        RECT 86.200 39.200 86.500 39.800 ;
        RECT 86.200 38.800 86.600 39.200 ;
        RECT 87.000 36.800 87.400 37.200 ;
        RECT 87.000 35.200 87.300 36.800 ;
        RECT 83.800 34.800 84.200 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 83.800 33.800 84.200 34.200 ;
        RECT 83.800 29.200 84.100 33.800 ;
        RECT 79.000 27.800 79.400 28.200 ;
        RECT 78.200 26.800 78.600 27.200 ;
        RECT 79.000 26.300 79.300 27.800 ;
        RECT 79.000 25.900 79.400 26.300 ;
        RECT 79.800 23.100 80.200 28.900 ;
        RECT 83.800 28.800 84.200 29.200 ;
        RECT 81.400 25.100 81.800 27.900 ;
        RECT 83.000 26.800 83.400 27.200 ;
        RECT 83.000 26.200 83.300 26.800 ;
        RECT 83.000 25.800 83.400 26.200 ;
        RECT 67.000 21.800 67.400 22.200 ;
        RECT 67.800 21.800 68.200 22.200 ;
        RECT 75.000 21.800 75.400 22.200 ;
        RECT 63.800 20.800 64.200 21.200 ;
        RECT 67.800 19.200 68.100 21.800 ;
        RECT 75.000 19.200 75.300 21.800 ;
        RECT 83.000 19.200 83.300 25.800 ;
        RECT 84.600 25.200 84.900 34.800 ;
        RECT 86.200 27.800 86.600 28.200 ;
        RECT 87.000 27.800 87.400 28.200 ;
        RECT 86.200 26.200 86.500 27.800 ;
        RECT 87.000 27.200 87.300 27.800 ;
        RECT 87.000 26.800 87.400 27.200 ;
        RECT 85.400 25.800 85.800 26.200 ;
        RECT 86.200 25.800 86.600 26.200 ;
        RECT 84.600 24.800 85.000 25.200 ;
        RECT 67.800 18.800 68.200 19.200 ;
        RECT 75.000 18.800 75.400 19.200 ;
        RECT 80.600 18.800 81.000 19.200 ;
        RECT 83.000 18.800 83.400 19.200 ;
        RECT 63.000 16.800 63.400 17.200 ;
        RECT 61.400 15.800 61.800 16.200 ;
        RECT 62.200 15.800 62.600 16.200 ;
        RECT 61.400 15.200 61.700 15.800 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 58.200 14.100 58.600 14.200 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 58.200 13.800 59.400 14.100 ;
        RECT 60.600 13.800 61.000 14.200 ;
        RECT 61.400 13.800 61.800 14.200 ;
        RECT 61.400 13.200 61.700 13.800 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 50.200 11.800 50.600 12.200 ;
        RECT 55.800 11.800 56.200 12.200 ;
        RECT 50.200 9.200 50.500 11.800 ;
        RECT 55.800 9.200 56.100 11.800 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 55.800 8.800 56.200 9.200 ;
        RECT 29.400 6.800 29.800 7.200 ;
        RECT 31.000 7.100 31.400 7.200 ;
        RECT 31.800 7.100 32.200 7.200 ;
        RECT 31.000 6.800 32.200 7.100 ;
        RECT 34.200 7.100 34.600 7.200 ;
        RECT 35.000 7.100 35.400 7.200 ;
        RECT 34.200 6.800 35.400 7.100 ;
        RECT 38.200 6.800 38.600 7.200 ;
        RECT 40.600 7.100 41.000 7.200 ;
        RECT 41.400 7.100 41.800 7.200 ;
        RECT 40.600 6.800 41.800 7.100 ;
        RECT 48.600 7.100 49.000 7.200 ;
        RECT 49.400 7.100 49.800 7.200 ;
        RECT 48.600 6.800 49.800 7.100 ;
        RECT 55.800 6.800 56.200 7.200 ;
        RECT 55.800 6.200 56.100 6.800 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 32.600 6.100 33.000 6.200 ;
        RECT 33.400 6.100 33.800 6.200 ;
        RECT 32.600 5.800 33.800 6.100 ;
        RECT 35.000 5.800 35.400 6.200 ;
        RECT 55.800 5.800 56.200 6.200 ;
        RECT 31.000 5.200 31.300 5.800 ;
        RECT 35.000 5.200 35.300 5.800 ;
        RECT 31.000 4.800 31.400 5.200 ;
        RECT 35.000 4.800 35.400 5.200 ;
        RECT 62.200 4.200 62.500 15.800 ;
        RECT 63.000 14.200 63.300 16.800 ;
        RECT 63.000 13.800 63.400 14.200 ;
        RECT 63.800 13.100 64.200 15.900 ;
        RECT 64.600 13.800 65.000 14.200 ;
        RECT 64.600 8.200 64.900 13.800 ;
        RECT 65.400 12.100 65.800 17.900 ;
        RECT 66.200 14.700 66.600 15.100 ;
        RECT 66.200 14.200 66.500 14.700 ;
        RECT 66.200 13.800 66.600 14.200 ;
        RECT 70.200 12.100 70.600 17.900 ;
        RECT 72.600 17.100 73.000 17.200 ;
        RECT 73.400 17.100 73.800 17.200 ;
        RECT 72.600 16.800 73.800 17.100 ;
        RECT 74.200 16.800 74.600 17.200 ;
        RECT 73.400 15.800 73.800 16.200 ;
        RECT 73.400 15.200 73.700 15.800 ;
        RECT 74.200 15.200 74.500 16.800 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 74.200 14.800 74.600 15.200 ;
        RECT 76.600 14.800 77.000 15.200 ;
        RECT 65.400 10.800 65.800 11.200 ;
        RECT 64.600 7.800 65.000 8.200 ;
        RECT 64.600 7.200 64.900 7.800 ;
        RECT 64.600 6.800 65.000 7.200 ;
        RECT 65.400 6.200 65.700 10.800 ;
        RECT 76.600 10.200 76.900 14.800 ;
        RECT 78.200 13.100 78.600 15.900 ;
        RECT 79.800 12.100 80.200 17.900 ;
        RECT 80.600 15.100 80.900 18.800 ;
        RECT 83.800 15.800 84.200 16.200 ;
        RECT 83.800 15.200 84.100 15.800 ;
        RECT 80.600 14.700 81.000 15.100 ;
        RECT 83.800 14.800 84.200 15.200 ;
        RECT 84.600 12.100 85.000 17.900 ;
        RECT 85.400 17.200 85.700 25.800 ;
        RECT 86.200 19.100 86.600 19.200 ;
        RECT 87.000 19.100 87.400 19.200 ;
        RECT 86.200 18.800 87.400 19.100 ;
        RECT 87.800 18.100 88.100 46.800 ;
        RECT 88.600 43.100 89.000 48.900 ;
        RECT 90.200 47.800 90.600 48.200 ;
        RECT 90.200 46.200 90.500 47.800 ;
        RECT 90.200 45.800 90.600 46.200 ;
        RECT 91.000 39.200 91.300 51.800 ;
        RECT 92.600 45.800 93.000 46.200 ;
        RECT 92.600 44.200 92.900 45.800 ;
        RECT 92.600 43.800 93.000 44.200 ;
        RECT 92.600 42.800 93.000 43.200 ;
        RECT 93.400 43.100 93.800 48.900 ;
        RECT 95.000 47.200 95.300 54.800 ;
        RECT 98.200 50.200 98.500 54.800 ;
        RECT 99.000 53.100 99.400 55.900 ;
        RECT 100.600 52.100 101.000 57.900 ;
        RECT 101.400 54.200 101.700 73.800 ;
        RECT 104.600 72.200 104.900 74.800 ;
        RECT 106.200 74.200 106.500 74.800 ;
        RECT 106.200 73.800 106.600 74.200 ;
        RECT 108.600 72.200 108.900 75.800 ;
        RECT 110.200 73.800 110.600 74.200 ;
        RECT 110.200 73.200 110.500 73.800 ;
        RECT 110.200 72.800 110.600 73.200 ;
        RECT 111.000 73.100 111.400 75.900 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 111.800 74.200 112.100 74.800 ;
        RECT 111.800 73.800 112.200 74.200 ;
        RECT 102.200 71.800 102.600 72.200 ;
        RECT 104.600 71.800 105.000 72.200 ;
        RECT 108.600 71.800 109.000 72.200 ;
        RECT 112.600 72.100 113.000 77.900 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 113.400 74.800 114.600 75.100 ;
        RECT 113.400 74.700 113.800 74.800 ;
        RECT 102.200 57.200 102.500 71.800 ;
        RECT 103.000 65.800 103.400 66.200 ;
        RECT 103.800 65.800 104.200 66.200 ;
        RECT 103.000 65.200 103.300 65.800 ;
        RECT 103.000 64.800 103.400 65.200 ;
        RECT 103.800 62.200 104.100 65.800 ;
        RECT 103.800 61.800 104.200 62.200 ;
        RECT 103.000 60.800 103.400 61.200 ;
        RECT 102.200 56.800 102.600 57.200 ;
        RECT 102.200 54.800 102.600 55.200 ;
        RECT 102.200 54.200 102.500 54.800 ;
        RECT 101.400 53.800 101.800 54.200 ;
        RECT 102.200 53.800 102.600 54.200 ;
        RECT 98.200 49.800 98.600 50.200 ;
        RECT 99.000 48.800 99.400 49.200 ;
        RECT 99.000 48.200 99.300 48.800 ;
        RECT 99.000 47.800 99.400 48.200 ;
        RECT 95.000 46.800 95.400 47.200 ;
        RECT 99.000 46.800 99.400 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 101.400 47.100 101.800 47.200 ;
        RECT 100.600 46.800 101.800 47.100 ;
        RECT 98.200 45.800 98.600 46.200 ;
        RECT 98.200 45.200 98.500 45.800 ;
        RECT 98.200 44.800 98.600 45.200 ;
        RECT 91.000 38.800 91.400 39.200 ;
        RECT 92.600 35.200 92.900 42.800 ;
        RECT 88.600 34.800 89.000 35.200 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 92.600 34.800 93.000 35.200 ;
        RECT 88.600 34.200 88.900 34.800 ;
        RECT 88.600 33.800 89.000 34.200 ;
        RECT 91.800 31.200 92.100 34.800 ;
        RECT 92.600 33.800 93.000 34.200 ;
        RECT 91.800 30.800 92.200 31.200 ;
        RECT 88.600 27.100 89.000 27.200 ;
        RECT 89.400 27.100 89.800 27.200 ;
        RECT 88.600 26.800 89.800 27.100 ;
        RECT 92.600 26.200 92.900 33.800 ;
        RECT 93.400 33.100 93.800 35.900 ;
        RECT 95.000 32.100 95.400 37.900 ;
        RECT 95.800 35.800 96.200 36.200 ;
        RECT 95.000 30.800 95.400 31.200 ;
        RECT 95.000 29.200 95.300 30.800 ;
        RECT 95.000 28.800 95.400 29.200 ;
        RECT 94.200 27.800 94.600 28.200 ;
        RECT 94.200 26.200 94.500 27.800 ;
        RECT 91.800 25.800 92.200 26.200 ;
        RECT 92.600 25.800 93.000 26.200 ;
        RECT 93.400 25.800 93.800 26.200 ;
        RECT 94.200 25.800 94.600 26.200 ;
        RECT 91.800 25.100 92.100 25.800 ;
        RECT 93.400 25.200 93.700 25.800 ;
        RECT 91.800 24.800 92.900 25.100 ;
        RECT 93.400 24.800 93.800 25.200 ;
        RECT 87.000 17.800 88.100 18.100 ;
        RECT 85.400 16.800 85.800 17.200 ;
        RECT 76.600 9.800 77.000 10.200 ;
        RECT 81.400 9.800 81.800 10.200 ;
        RECT 81.400 9.200 81.700 9.800 ;
        RECT 66.200 8.800 66.600 9.200 ;
        RECT 71.000 8.800 71.400 9.200 ;
        RECT 79.800 9.100 80.200 9.200 ;
        RECT 80.600 9.100 81.000 9.200 ;
        RECT 66.200 6.200 66.500 8.800 ;
        RECT 71.000 8.200 71.300 8.800 ;
        RECT 71.000 7.800 71.400 8.200 ;
        RECT 68.600 7.100 69.000 7.200 ;
        RECT 69.400 7.100 69.800 7.200 ;
        RECT 68.600 6.800 69.800 7.100 ;
        RECT 65.400 5.800 65.800 6.200 ;
        RECT 66.200 5.800 66.600 6.200 ;
        RECT 71.800 5.100 72.200 7.900 ;
        RECT 72.600 7.800 73.000 8.200 ;
        RECT 72.600 7.200 72.900 7.800 ;
        RECT 72.600 6.800 73.000 7.200 ;
        RECT 62.200 3.800 62.600 4.200 ;
        RECT 73.400 3.100 73.800 8.900 ;
        RECT 74.200 6.800 74.600 7.200 ;
        RECT 74.200 6.300 74.500 6.800 ;
        RECT 74.200 5.900 74.600 6.300 ;
        RECT 78.200 3.100 78.600 8.900 ;
        RECT 79.800 8.800 81.000 9.100 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 83.800 3.100 84.200 8.900 ;
        RECT 87.000 7.200 87.300 17.800 ;
        RECT 87.800 16.800 88.200 17.200 ;
        RECT 87.800 13.200 88.100 16.800 ;
        RECT 91.000 16.100 91.400 16.200 ;
        RECT 91.800 16.100 92.200 16.200 ;
        RECT 91.000 15.800 92.200 16.100 ;
        RECT 92.600 15.200 92.900 24.800 ;
        RECT 93.400 17.100 93.800 17.200 ;
        RECT 94.200 17.100 94.600 17.200 ;
        RECT 93.400 16.800 94.600 17.100 ;
        RECT 93.400 15.800 93.800 16.200 ;
        RECT 93.400 15.200 93.700 15.800 ;
        RECT 95.800 15.200 96.100 35.800 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 97.400 34.200 97.700 34.800 ;
        RECT 96.600 33.800 97.000 34.200 ;
        RECT 97.400 33.800 97.800 34.200 ;
        RECT 96.600 19.200 96.900 33.800 ;
        RECT 99.000 29.200 99.300 46.800 ;
        RECT 103.000 46.200 103.300 60.800 ;
        RECT 104.600 58.200 104.900 71.800 ;
        RECT 113.400 69.800 113.800 70.200 ;
        RECT 107.000 68.800 107.400 69.200 ;
        RECT 106.200 66.800 106.600 67.200 ;
        RECT 106.200 66.200 106.500 66.800 ;
        RECT 107.000 66.200 107.300 68.800 ;
        RECT 111.000 66.800 111.400 67.200 ;
        RECT 112.600 66.800 113.000 67.200 ;
        RECT 111.000 66.200 111.300 66.800 ;
        RECT 106.200 65.800 106.600 66.200 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 109.400 66.100 109.800 66.200 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 109.400 65.800 110.600 66.100 ;
        RECT 111.000 65.800 111.400 66.200 ;
        RECT 111.000 64.800 111.400 65.200 ;
        RECT 107.800 63.800 108.200 64.200 ;
        RECT 107.800 59.200 108.100 63.800 ;
        RECT 107.800 58.800 108.200 59.200 ;
        RECT 104.600 57.800 105.000 58.200 ;
        RECT 104.600 53.800 105.000 54.200 ;
        RECT 103.800 52.800 104.200 53.200 ;
        RECT 103.800 50.200 104.100 52.800 ;
        RECT 103.800 49.800 104.200 50.200 ;
        RECT 103.800 49.200 104.100 49.800 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 103.000 45.800 103.400 46.200 ;
        RECT 99.800 32.100 100.200 37.900 ;
        RECT 104.600 36.200 104.900 53.800 ;
        RECT 105.400 52.100 105.800 57.900 ;
        RECT 110.200 55.800 110.600 56.200 ;
        RECT 110.200 55.200 110.500 55.800 ;
        RECT 111.000 55.200 111.300 64.800 ;
        RECT 112.600 64.200 112.900 66.800 ;
        RECT 113.400 66.200 113.700 69.800 ;
        RECT 114.200 66.800 114.600 67.200 ;
        RECT 114.200 66.200 114.500 66.800 ;
        RECT 113.400 65.800 113.800 66.200 ;
        RECT 114.200 65.800 114.600 66.200 ;
        RECT 112.600 63.800 113.000 64.200 ;
        RECT 111.800 61.800 112.200 62.200 ;
        RECT 111.800 56.200 112.100 61.800 ;
        RECT 113.400 56.800 113.800 57.200 ;
        RECT 111.800 55.800 112.200 56.200 ;
        RECT 108.600 55.100 109.000 55.200 ;
        RECT 109.400 55.100 109.800 55.200 ;
        RECT 108.600 54.800 109.800 55.100 ;
        RECT 110.200 54.800 110.600 55.200 ;
        RECT 111.000 54.800 111.400 55.200 ;
        RECT 111.800 55.100 112.200 55.200 ;
        RECT 112.600 55.100 113.000 55.200 ;
        RECT 111.800 54.800 113.000 55.100 ;
        RECT 109.400 50.800 109.800 51.200 ;
        RECT 106.200 43.100 106.600 48.900 ;
        RECT 109.400 46.200 109.700 50.800 ;
        RECT 110.200 46.800 110.600 47.200 ;
        RECT 109.400 45.800 109.800 46.200 ;
        RECT 110.200 44.200 110.500 46.800 ;
        RECT 110.200 43.800 110.600 44.200 ;
        RECT 111.000 43.100 111.400 48.900 ;
        RECT 111.800 45.200 112.100 54.800 ;
        RECT 113.400 54.200 113.700 56.800 ;
        RECT 115.000 55.200 115.300 89.800 ;
        RECT 115.800 83.100 116.200 88.900 ;
        RECT 116.600 75.200 116.900 113.800 ;
        RECT 117.400 112.100 117.800 117.900 ;
        RECT 121.400 115.200 121.700 126.800 ;
        RECT 119.000 115.100 119.400 115.200 ;
        RECT 119.800 115.100 120.200 115.200 ;
        RECT 119.000 114.800 120.200 115.100 ;
        RECT 121.400 114.800 121.800 115.200 ;
        RECT 122.200 112.100 122.600 117.900 ;
        RECT 123.000 116.800 123.400 117.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 117.400 110.800 117.800 111.200 ;
        RECT 117.400 109.200 117.700 110.800 ;
        RECT 117.400 108.800 117.800 109.200 ;
        RECT 123.000 107.200 123.300 116.800 ;
        RECT 124.600 116.200 124.900 116.800 ;
        RECT 124.600 115.800 125.000 116.200 ;
        RECT 125.400 114.200 125.700 130.800 ;
        RECT 127.800 128.200 128.100 131.800 ;
        RECT 127.800 127.800 128.200 128.200 ;
        RECT 127.800 127.200 128.100 127.800 ;
        RECT 127.800 126.800 128.200 127.200 ;
        RECT 128.600 125.200 128.900 133.800 ;
        RECT 129.400 130.800 129.800 131.200 ;
        RECT 129.400 126.200 129.700 130.800 ;
        RECT 130.200 129.200 130.500 154.800 ;
        RECT 131.000 154.200 131.300 154.800 ;
        RECT 131.000 153.800 131.400 154.200 ;
        RECT 131.800 153.800 132.200 154.200 ;
        RECT 131.800 148.200 132.100 153.800 ;
        RECT 132.600 153.100 133.000 155.900 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 133.400 153.200 133.700 153.800 ;
        RECT 133.400 152.800 133.800 153.200 ;
        RECT 134.200 152.100 134.600 157.900 ;
        RECT 135.800 155.800 136.200 156.200 ;
        RECT 135.800 155.200 136.100 155.800 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 136.600 154.800 137.000 155.200 ;
        RECT 136.600 152.200 136.900 154.800 ;
        RECT 136.600 151.800 137.000 152.200 ;
        RECT 136.600 149.200 136.900 151.800 ;
        RECT 138.200 150.200 138.500 165.800 ;
        RECT 141.400 162.200 141.700 166.800 ;
        RECT 142.200 166.200 142.500 176.800 ;
        RECT 148.600 175.800 149.000 176.200 ;
        RECT 148.600 175.200 148.900 175.800 ;
        RECT 147.000 175.100 147.400 175.200 ;
        RECT 147.800 175.100 148.200 175.200 ;
        RECT 147.000 174.800 148.200 175.100 ;
        RECT 148.600 174.800 149.000 175.200 ;
        RECT 149.400 175.100 149.800 175.200 ;
        RECT 150.200 175.100 150.600 175.200 ;
        RECT 149.400 174.800 150.600 175.100 ;
        RECT 152.600 174.800 153.000 175.200 ;
        RECT 144.600 174.100 145.000 174.200 ;
        RECT 145.400 174.100 145.800 174.200 ;
        RECT 144.600 173.800 145.800 174.100 ;
        RECT 146.200 169.800 146.600 170.200 ;
        RECT 143.000 167.800 143.400 168.200 ;
        RECT 143.000 167.200 143.300 167.800 ;
        RECT 143.000 166.800 143.400 167.200 ;
        RECT 144.600 166.800 145.000 167.200 ;
        RECT 142.200 165.800 142.600 166.200 ;
        RECT 143.800 165.800 144.200 166.200 ;
        RECT 143.000 164.800 143.400 165.200 ;
        RECT 141.400 161.800 141.800 162.200 ;
        RECT 139.800 159.800 140.200 160.200 ;
        RECT 139.000 152.100 139.400 157.900 ;
        RECT 138.200 149.800 138.600 150.200 ;
        RECT 139.800 149.200 140.100 159.800 ;
        RECT 143.000 159.200 143.300 164.800 ;
        RECT 143.000 158.800 143.400 159.200 ;
        RECT 141.400 157.100 141.800 157.200 ;
        RECT 142.200 157.100 142.600 157.200 ;
        RECT 141.400 156.800 142.600 157.100 ;
        RECT 142.200 155.800 142.600 156.200 ;
        RECT 142.200 155.200 142.500 155.800 ;
        RECT 142.200 154.800 142.600 155.200 ;
        RECT 143.800 154.200 144.100 165.800 ;
        RECT 144.600 165.200 144.900 166.800 ;
        RECT 146.200 166.200 146.500 169.800 ;
        RECT 146.200 165.800 146.600 166.200 ;
        RECT 144.600 164.800 145.000 165.200 ;
        RECT 144.600 162.800 145.000 163.200 ;
        RECT 144.600 157.200 144.900 162.800 ;
        RECT 147.000 157.200 147.300 174.800 ;
        RECT 148.600 174.200 148.900 174.800 ;
        RECT 152.600 174.200 152.900 174.800 ;
        RECT 148.600 173.800 149.000 174.200 ;
        RECT 150.200 173.800 150.600 174.200 ;
        RECT 152.600 173.800 153.000 174.200 ;
        RECT 150.200 173.200 150.500 173.800 ;
        RECT 147.800 172.800 148.200 173.200 ;
        RECT 150.200 172.800 150.600 173.200 ;
        RECT 151.800 173.100 152.200 173.200 ;
        RECT 152.600 173.100 153.000 173.200 ;
        RECT 156.600 173.100 157.000 175.900 ;
        RECT 151.800 172.800 153.000 173.100 ;
        RECT 147.800 169.200 148.100 172.800 ;
        RECT 158.200 172.100 158.600 177.900 ;
        RECT 160.600 177.200 160.900 193.800 ;
        RECT 161.400 183.100 161.800 188.900 ;
        RECT 162.200 186.200 162.500 206.800 ;
        RECT 163.000 204.800 163.400 205.200 ;
        RECT 163.000 204.200 163.300 204.800 ;
        RECT 164.600 204.200 164.900 206.800 ;
        RECT 163.000 203.800 163.400 204.200 ;
        RECT 164.600 203.800 165.000 204.200 ;
        RECT 163.800 192.100 164.200 197.900 ;
        RECT 164.600 191.200 164.900 203.800 ;
        RECT 167.800 203.100 168.200 208.900 ;
        RECT 171.800 208.200 172.100 213.800 ;
        RECT 175.000 212.100 175.400 217.900 ;
        RECT 177.400 216.800 177.800 217.200 ;
        RECT 175.800 215.800 176.200 216.200 ;
        RECT 175.800 214.200 176.100 215.800 ;
        RECT 175.800 213.800 176.200 214.200 ;
        RECT 176.600 213.100 177.000 215.900 ;
        RECT 177.400 214.200 177.700 216.800 ;
        RECT 177.400 213.800 177.800 214.200 ;
        RECT 178.200 213.200 178.500 225.800 ;
        RECT 179.000 223.800 179.400 224.200 ;
        RECT 181.400 223.800 181.800 224.200 ;
        RECT 179.000 216.200 179.300 223.800 ;
        RECT 179.000 215.800 179.400 216.200 ;
        RECT 181.400 215.200 181.700 223.800 ;
        RECT 182.200 223.200 182.500 225.800 ;
        RECT 183.000 224.800 183.400 225.200 ;
        RECT 184.600 224.800 185.000 225.200 ;
        RECT 183.000 224.200 183.300 224.800 ;
        RECT 183.000 223.800 183.400 224.200 ;
        RECT 182.200 222.800 182.600 223.200 ;
        RECT 183.800 221.800 184.200 222.200 ;
        RECT 183.000 216.100 183.400 216.200 ;
        RECT 183.800 216.100 184.100 221.800 ;
        RECT 184.600 219.200 184.900 224.800 ;
        RECT 187.000 219.200 187.300 233.800 ;
        RECT 187.800 232.100 188.200 237.900 ;
        RECT 188.600 235.800 189.000 236.200 ;
        RECT 188.600 235.100 188.900 235.800 ;
        RECT 188.600 234.700 189.000 235.100 ;
        RECT 192.600 232.100 193.000 237.900 ;
        RECT 194.200 237.100 194.600 237.200 ;
        RECT 195.000 237.100 195.400 237.200 ;
        RECT 194.200 236.800 195.400 237.100 ;
        RECT 195.800 231.800 196.200 232.200 ;
        RECT 198.200 232.100 198.600 237.900 ;
        RECT 199.800 234.800 200.200 235.200 ;
        RECT 187.800 223.100 188.200 228.900 ;
        RECT 191.000 226.800 191.400 227.200 ;
        RECT 190.200 225.800 190.600 226.200 ;
        RECT 190.200 225.200 190.500 225.800 ;
        RECT 190.200 224.800 190.600 225.200 ;
        RECT 184.600 218.800 185.000 219.200 ;
        RECT 187.000 218.800 187.400 219.200 ;
        RECT 183.000 215.800 184.100 216.100 ;
        RECT 187.000 216.200 187.300 218.800 ;
        RECT 187.000 215.800 187.400 216.200 ;
        RECT 179.000 214.800 179.400 215.200 ;
        RECT 181.400 214.800 181.800 215.200 ;
        RECT 183.800 215.100 184.200 215.200 ;
        RECT 184.600 215.100 185.000 215.200 ;
        RECT 183.800 214.800 185.000 215.100 ;
        RECT 179.000 214.200 179.300 214.800 ;
        RECT 179.000 213.800 179.400 214.200 ;
        RECT 182.200 213.800 182.600 214.200 ;
        RECT 185.400 213.800 185.800 214.200 ;
        RECT 182.200 213.200 182.500 213.800 ;
        RECT 178.200 212.800 178.600 213.200 ;
        RECT 182.200 212.800 182.600 213.200 ;
        RECT 171.800 207.800 172.200 208.200 ;
        RECT 171.000 206.800 171.400 207.200 ;
        RECT 171.000 206.200 171.300 206.800 ;
        RECT 169.400 205.800 169.800 206.200 ;
        RECT 171.000 205.800 171.400 206.200 ;
        RECT 167.000 195.800 167.400 196.200 ;
        RECT 167.000 195.200 167.300 195.800 ;
        RECT 167.000 194.800 167.400 195.200 ;
        RECT 168.600 192.100 169.000 197.900 ;
        RECT 169.400 194.200 169.700 205.800 ;
        RECT 172.600 203.100 173.000 208.900 ;
        RECT 174.200 205.100 174.600 207.900 ;
        RECT 177.400 203.100 177.800 208.900 ;
        RECT 179.000 206.100 179.400 206.200 ;
        RECT 178.200 205.800 179.400 206.100 ;
        RECT 180.600 205.800 181.000 206.200 ;
        RECT 175.000 202.100 175.400 202.200 ;
        RECT 174.200 201.800 175.400 202.100 ;
        RECT 173.400 197.800 173.800 198.200 ;
        RECT 169.400 193.800 169.800 194.200 ;
        RECT 170.200 193.100 170.600 195.900 ;
        RECT 173.400 195.200 173.700 197.800 ;
        RECT 173.400 194.800 173.800 195.200 ;
        RECT 174.200 193.200 174.500 201.800 ;
        RECT 178.200 199.200 178.500 205.800 ;
        RECT 179.000 200.800 179.400 201.200 ;
        RECT 178.200 198.800 178.600 199.200 ;
        RECT 179.000 195.200 179.300 200.800 ;
        RECT 179.000 194.800 179.400 195.200 ;
        RECT 179.800 194.800 180.200 195.200 ;
        RECT 179.000 193.200 179.300 194.800 ;
        RECT 179.800 194.200 180.100 194.800 ;
        RECT 180.600 194.200 180.900 205.800 ;
        RECT 182.200 203.100 182.600 208.900 ;
        RECT 184.600 208.800 185.000 209.200 ;
        RECT 183.000 207.800 183.400 208.200 ;
        RECT 183.000 207.200 183.300 207.800 ;
        RECT 183.000 206.800 183.400 207.200 ;
        RECT 183.800 205.100 184.200 207.900 ;
        RECT 184.600 206.200 184.900 208.800 ;
        RECT 184.600 205.800 185.000 206.200 ;
        RECT 184.600 203.800 185.000 204.200 ;
        RECT 184.600 199.200 184.900 203.800 ;
        RECT 185.400 201.200 185.700 213.800 ;
        RECT 187.000 203.100 187.400 208.900 ;
        RECT 191.000 208.200 191.300 226.800 ;
        RECT 192.600 223.100 193.000 228.900 ;
        RECT 195.800 228.200 196.100 231.800 ;
        RECT 196.600 229.800 197.000 230.200 ;
        RECT 196.600 228.200 196.900 229.800 ;
        RECT 199.800 229.200 200.100 234.800 ;
        RECT 203.000 232.100 203.400 237.900 ;
        RECT 203.800 234.800 204.200 235.200 ;
        RECT 203.800 234.200 204.100 234.800 ;
        RECT 203.800 233.800 204.200 234.200 ;
        RECT 198.200 229.100 198.600 229.200 ;
        RECT 199.000 229.100 199.400 229.200 ;
        RECT 198.200 228.800 199.400 229.100 ;
        RECT 199.800 228.800 200.200 229.200 ;
        RECT 200.600 229.100 201.000 229.200 ;
        RECT 201.400 229.100 201.800 229.200 ;
        RECT 200.600 228.800 201.800 229.100 ;
        RECT 195.000 228.100 195.400 228.200 ;
        RECT 195.800 228.100 196.200 228.200 ;
        RECT 193.400 226.800 193.800 227.200 ;
        RECT 193.400 226.200 193.700 226.800 ;
        RECT 193.400 225.800 193.800 226.200 ;
        RECT 194.200 225.100 194.600 227.900 ;
        RECT 195.000 227.800 196.200 228.100 ;
        RECT 196.600 227.800 197.000 228.200 ;
        RECT 199.000 227.800 199.400 228.200 ;
        RECT 196.600 226.200 196.900 227.800 ;
        RECT 199.000 227.200 199.300 227.800 ;
        RECT 199.000 226.800 199.400 227.200 ;
        RECT 196.600 225.800 197.000 226.200 ;
        RECT 199.800 225.800 200.200 226.200 ;
        RECT 199.800 222.200 200.100 225.800 ;
        RECT 203.000 223.100 203.400 228.900 ;
        RECT 203.800 227.200 204.100 233.800 ;
        RECT 204.600 233.100 205.000 235.900 ;
        RECT 224.600 235.800 225.000 236.200 ;
        RECT 206.200 235.100 206.600 235.200 ;
        RECT 207.000 235.100 207.400 235.200 ;
        RECT 206.200 234.800 207.400 235.100 ;
        RECT 221.400 234.800 221.800 235.200 ;
        RECT 222.200 234.800 222.600 235.200 ;
        RECT 221.400 234.200 221.700 234.800 ;
        RECT 222.200 234.200 222.500 234.800 ;
        RECT 224.600 234.200 224.900 235.800 ;
        RECT 213.400 233.800 213.800 234.200 ;
        RECT 214.200 233.800 214.600 234.200 ;
        RECT 220.600 233.800 221.000 234.200 ;
        RECT 221.400 233.800 221.800 234.200 ;
        RECT 222.200 233.800 222.600 234.200 ;
        RECT 224.600 233.800 225.000 234.200 ;
        RECT 226.200 233.800 226.600 234.200 ;
        RECT 227.000 233.800 227.400 234.200 ;
        RECT 213.400 233.200 213.700 233.800 ;
        RECT 213.400 232.800 213.800 233.200 ;
        RECT 204.600 228.800 205.000 229.200 ;
        RECT 203.800 226.800 204.200 227.200 ;
        RECT 195.000 221.800 195.400 222.200 ;
        RECT 199.800 221.800 200.200 222.200 ;
        RECT 192.600 217.800 193.000 218.200 ;
        RECT 192.600 214.200 192.900 217.800 ;
        RECT 194.200 214.800 194.600 215.200 ;
        RECT 192.600 213.800 193.000 214.200 ;
        RECT 193.400 213.800 193.800 214.200 ;
        RECT 193.400 213.200 193.700 213.800 ;
        RECT 193.400 212.800 193.800 213.200 ;
        RECT 194.200 212.200 194.500 214.800 ;
        RECT 194.200 211.800 194.600 212.200 ;
        RECT 191.000 207.800 191.400 208.200 ;
        RECT 190.200 205.800 190.600 206.200 ;
        RECT 190.200 204.200 190.500 205.800 ;
        RECT 190.200 203.800 190.600 204.200 ;
        RECT 191.800 203.100 192.200 208.900 ;
        RECT 193.400 205.100 193.800 207.900 ;
        RECT 194.200 206.800 194.600 207.200 ;
        RECT 194.200 202.200 194.500 206.800 ;
        RECT 195.000 206.200 195.300 221.800 ;
        RECT 198.200 216.800 198.600 217.200 ;
        RECT 196.600 215.800 197.000 216.200 ;
        RECT 195.800 214.800 196.200 215.200 ;
        RECT 195.800 214.200 196.100 214.800 ;
        RECT 195.800 213.800 196.200 214.200 ;
        RECT 196.600 212.200 196.900 215.800 ;
        RECT 198.200 214.200 198.500 216.800 ;
        RECT 198.200 213.800 198.600 214.200 ;
        RECT 196.600 211.800 197.000 212.200 ;
        RECT 199.000 211.800 199.400 212.200 ;
        RECT 201.400 212.100 201.800 217.900 ;
        RECT 203.000 214.800 203.400 215.200 ;
        RECT 199.000 211.200 199.300 211.800 ;
        RECT 197.400 210.800 197.800 211.200 ;
        RECT 199.000 210.800 199.400 211.200 ;
        RECT 196.600 209.800 197.000 210.200 ;
        RECT 196.600 209.200 196.900 209.800 ;
        RECT 196.600 208.800 197.000 209.200 ;
        RECT 195.000 205.800 195.400 206.200 ;
        RECT 194.200 201.800 194.600 202.200 ;
        RECT 185.400 200.800 185.800 201.200 ;
        RECT 188.600 200.800 189.000 201.200 ;
        RECT 184.600 198.800 185.000 199.200 ;
        RECT 187.000 198.800 187.400 199.200 ;
        RECT 182.200 195.800 182.600 196.200 ;
        RECT 182.200 195.200 182.500 195.800 ;
        RECT 187.000 195.200 187.300 198.800 ;
        RECT 182.200 194.800 182.600 195.200 ;
        RECT 183.800 195.100 184.200 195.200 ;
        RECT 184.600 195.100 185.000 195.200 ;
        RECT 183.800 194.800 185.000 195.100 ;
        RECT 186.200 194.800 186.600 195.200 ;
        RECT 187.000 194.800 187.400 195.200 ;
        RECT 179.800 193.800 180.200 194.200 ;
        RECT 180.600 193.800 181.000 194.200 ;
        RECT 171.800 192.800 172.200 193.200 ;
        RECT 174.200 192.800 174.600 193.200 ;
        RECT 179.000 192.800 179.400 193.200 ;
        RECT 171.800 192.200 172.100 192.800 ;
        RECT 169.400 191.800 169.800 192.200 ;
        RECT 171.800 191.800 172.200 192.200 ;
        RECT 164.600 190.800 165.000 191.200 ;
        RECT 163.800 188.800 164.200 189.200 ;
        RECT 163.800 188.200 164.100 188.800 ;
        RECT 163.800 187.800 164.200 188.200 ;
        RECT 164.600 188.100 165.000 188.200 ;
        RECT 165.400 188.100 165.800 188.200 ;
        RECT 164.600 187.800 165.800 188.100 ;
        RECT 165.400 187.100 165.800 187.200 ;
        RECT 166.200 187.100 166.600 187.200 ;
        RECT 165.400 186.800 166.600 187.100 ;
        RECT 169.400 186.200 169.700 191.800 ;
        RECT 171.000 187.800 171.400 188.200 ;
        RECT 171.000 186.200 171.300 187.800 ;
        RECT 174.200 186.200 174.500 192.800 ;
        RECT 175.000 188.800 175.400 189.200 ;
        RECT 175.000 186.200 175.300 188.800 ;
        RECT 179.000 187.800 179.400 188.200 ;
        RECT 179.000 186.200 179.300 187.800 ;
        RECT 162.200 185.800 162.600 186.200 ;
        RECT 169.400 185.800 169.800 186.200 ;
        RECT 170.200 185.800 170.600 186.200 ;
        RECT 171.000 185.800 171.400 186.200 ;
        RECT 174.200 185.800 174.600 186.200 ;
        RECT 175.000 185.800 175.400 186.200 ;
        RECT 175.800 185.800 176.200 186.200 ;
        RECT 176.600 185.800 177.000 186.200 ;
        RECT 179.000 185.800 179.400 186.200 ;
        RECT 179.800 185.800 180.200 186.200 ;
        RECT 180.600 186.100 180.900 193.800 ;
        RECT 181.400 186.100 181.800 186.200 ;
        RECT 180.600 185.800 181.800 186.100 ;
        RECT 183.800 185.800 184.200 186.200 ;
        RECT 162.200 183.800 162.600 184.200 ;
        RECT 162.200 179.200 162.500 183.800 ;
        RECT 165.400 180.800 165.800 181.200 ;
        RECT 165.400 179.200 165.700 180.800 ;
        RECT 162.200 178.800 162.600 179.200 ;
        RECT 165.400 178.800 165.800 179.200 ;
        RECT 160.600 176.800 161.000 177.200 ;
        RECT 159.800 175.100 160.200 175.200 ;
        RECT 160.600 175.100 161.000 175.200 ;
        RECT 159.800 174.800 161.000 175.100 ;
        RECT 159.000 172.800 159.400 173.200 ;
        RECT 159.000 172.200 159.300 172.800 ;
        RECT 159.000 171.800 159.400 172.200 ;
        RECT 163.000 172.100 163.400 177.900 ;
        RECT 169.400 177.200 169.700 185.800 ;
        RECT 164.600 176.800 165.000 177.200 ;
        RECT 169.400 176.800 169.800 177.200 ;
        RECT 158.200 169.800 158.600 170.200 ;
        RECT 147.800 168.800 148.200 169.200 ;
        RECT 152.600 168.800 153.000 169.200 ;
        RECT 149.400 167.800 149.800 168.200 ;
        RECT 149.400 167.200 149.700 167.800 ;
        RECT 152.600 167.200 152.900 168.800 ;
        RECT 149.400 166.800 149.800 167.200 ;
        RECT 150.200 166.800 150.600 167.200 ;
        RECT 152.600 166.800 153.000 167.200 ;
        RECT 150.200 166.200 150.500 166.800 ;
        RECT 158.200 166.200 158.500 169.800 ;
        RECT 147.800 166.100 148.200 166.200 ;
        RECT 148.600 166.100 149.000 166.200 ;
        RECT 147.800 165.800 149.000 166.100 ;
        RECT 150.200 165.800 150.600 166.200 ;
        RECT 151.800 165.800 152.200 166.200 ;
        RECT 153.400 165.800 153.800 166.200 ;
        RECT 154.200 165.800 154.600 166.200 ;
        RECT 155.800 166.100 156.200 166.200 ;
        RECT 156.600 166.100 157.000 166.200 ;
        RECT 155.800 165.800 157.000 166.100 ;
        RECT 158.200 165.800 158.600 166.200 ;
        RECT 147.800 164.800 148.200 165.200 ;
        RECT 147.800 164.200 148.100 164.800 ;
        RECT 147.800 163.800 148.200 164.200 ;
        RECT 151.800 162.200 152.100 165.800 ;
        RECT 152.600 164.800 153.000 165.200 ;
        RECT 151.800 161.800 152.200 162.200 ;
        RECT 144.600 156.800 145.000 157.200 ;
        RECT 147.000 156.800 147.400 157.200 ;
        RECT 148.600 156.800 149.000 157.200 ;
        RECT 144.600 154.200 144.900 156.800 ;
        RECT 145.400 155.800 145.800 156.200 ;
        RECT 146.200 156.100 146.600 156.200 ;
        RECT 147.000 156.100 147.400 156.200 ;
        RECT 146.200 155.800 147.400 156.100 ;
        RECT 145.400 155.100 145.700 155.800 ;
        RECT 145.400 154.800 146.500 155.100 ;
        RECT 146.200 154.200 146.500 154.800 ;
        RECT 143.800 153.800 144.200 154.200 ;
        RECT 144.600 153.800 145.000 154.200 ;
        RECT 146.200 153.800 146.600 154.200 ;
        RECT 148.600 154.100 148.900 156.800 ;
        RECT 149.400 155.800 149.800 156.200 ;
        RECT 150.200 155.800 150.600 156.200 ;
        RECT 149.400 155.200 149.700 155.800 ;
        RECT 150.200 155.200 150.500 155.800 ;
        RECT 149.400 154.800 149.800 155.200 ;
        RECT 150.200 154.800 150.600 155.200 ;
        RECT 151.800 154.200 152.100 161.800 ;
        RECT 149.400 154.100 149.800 154.200 ;
        RECT 148.600 153.800 149.800 154.100 ;
        RECT 151.800 153.800 152.200 154.200 ;
        RECT 143.800 153.200 144.100 153.800 ;
        RECT 143.800 152.800 144.200 153.200 ;
        RECT 141.400 151.800 141.800 152.200 ;
        RECT 133.400 148.800 133.800 149.200 ;
        RECT 136.600 148.800 137.000 149.200 ;
        RECT 139.800 148.800 140.200 149.200 ;
        RECT 131.000 145.100 131.400 147.900 ;
        RECT 131.800 147.800 132.200 148.200 ;
        RECT 133.400 147.200 133.700 148.800 ;
        RECT 131.800 147.100 132.200 147.200 ;
        RECT 132.600 147.100 133.000 147.200 ;
        RECT 131.800 146.800 133.000 147.100 ;
        RECT 133.400 146.800 133.800 147.200 ;
        RECT 134.200 147.100 134.600 147.200 ;
        RECT 135.000 147.100 135.400 147.200 ;
        RECT 134.200 146.800 135.400 147.100 ;
        RECT 140.600 146.800 141.000 147.200 ;
        RECT 135.000 146.100 135.400 146.200 ;
        RECT 135.800 146.100 136.200 146.200 ;
        RECT 135.000 145.800 136.200 146.100 ;
        RECT 137.400 145.800 137.800 146.200 ;
        RECT 138.200 145.800 138.600 146.200 ;
        RECT 135.000 145.200 135.300 145.800 ;
        RECT 131.800 144.800 132.200 145.200 ;
        RECT 135.000 144.800 135.400 145.200 ;
        RECT 131.800 144.100 132.100 144.800 ;
        RECT 131.000 143.800 132.100 144.100 ;
        RECT 131.000 129.200 131.300 143.800 ;
        RECT 134.200 141.800 134.600 142.200 ;
        RECT 131.800 139.800 132.200 140.200 ;
        RECT 131.800 139.200 132.100 139.800 ;
        RECT 134.200 139.200 134.500 141.800 ;
        RECT 135.800 140.800 136.200 141.200 ;
        RECT 131.800 138.800 132.200 139.200 ;
        RECT 134.200 138.800 134.600 139.200 ;
        RECT 135.800 135.200 136.100 140.800 ;
        RECT 137.400 139.200 137.700 145.800 ;
        RECT 138.200 141.200 138.500 145.800 ;
        RECT 139.000 143.800 139.400 144.200 ;
        RECT 138.200 140.800 138.600 141.200 ;
        RECT 139.000 139.200 139.300 143.800 ;
        RECT 139.800 141.800 140.200 142.200 ;
        RECT 137.400 138.800 137.800 139.200 ;
        RECT 139.000 138.800 139.400 139.200 ;
        RECT 139.800 138.200 140.100 141.800 ;
        RECT 139.800 137.800 140.200 138.200 ;
        RECT 140.600 137.200 140.900 146.800 ;
        RECT 141.400 139.200 141.700 151.800 ;
        RECT 143.800 150.800 144.200 151.200 ;
        RECT 149.400 150.800 149.800 151.200 ;
        RECT 142.200 146.100 142.600 146.200 ;
        RECT 143.000 146.100 143.400 146.200 ;
        RECT 142.200 145.800 143.400 146.100 ;
        RECT 143.000 145.200 143.300 145.800 ;
        RECT 143.000 144.800 143.400 145.200 ;
        RECT 142.200 144.100 142.600 144.200 ;
        RECT 143.000 144.100 143.400 144.200 ;
        RECT 142.200 143.800 143.400 144.100 ;
        RECT 143.000 142.800 143.400 143.200 ;
        RECT 143.000 142.200 143.300 142.800 ;
        RECT 143.000 141.800 143.400 142.200 ;
        RECT 143.800 139.200 144.100 150.800 ;
        RECT 146.200 147.800 146.600 148.200 ;
        RECT 147.800 147.800 148.200 148.200 ;
        RECT 145.400 146.800 145.800 147.200 ;
        RECT 145.400 146.200 145.700 146.800 ;
        RECT 144.600 145.800 145.000 146.200 ;
        RECT 145.400 145.800 145.800 146.200 ;
        RECT 144.600 145.200 144.900 145.800 ;
        RECT 144.600 144.800 145.000 145.200 ;
        RECT 141.400 138.800 141.800 139.200 ;
        RECT 143.800 138.800 144.200 139.200 ;
        RECT 140.600 136.800 141.000 137.200 ;
        RECT 138.200 135.800 138.600 136.200 ;
        RECT 135.800 134.800 136.200 135.200 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 138.200 134.200 138.500 135.800 ;
        RECT 140.600 134.200 140.900 136.800 ;
        RECT 143.000 135.800 143.400 136.200 ;
        RECT 135.800 134.100 136.200 134.200 ;
        RECT 136.600 134.100 137.000 134.200 ;
        RECT 135.800 133.800 137.000 134.100 ;
        RECT 138.200 133.800 138.600 134.200 ;
        RECT 139.800 133.800 140.200 134.200 ;
        RECT 140.600 133.800 141.000 134.200 ;
        RECT 139.800 133.200 140.100 133.800 ;
        RECT 143.000 133.200 143.300 135.800 ;
        RECT 144.600 135.200 144.900 144.800 ;
        RECT 145.400 141.800 145.800 142.200 ;
        RECT 145.400 140.200 145.700 141.800 ;
        RECT 145.400 139.800 145.800 140.200 ;
        RECT 146.200 139.200 146.500 147.800 ;
        RECT 147.800 145.200 148.100 147.800 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 148.600 145.200 148.900 145.800 ;
        RECT 149.400 145.200 149.700 150.800 ;
        RECT 151.000 145.800 151.400 146.200 ;
        RECT 147.000 145.100 147.400 145.200 ;
        RECT 147.800 145.100 148.200 145.200 ;
        RECT 147.000 144.800 148.200 145.100 ;
        RECT 148.600 144.800 149.000 145.200 ;
        RECT 149.400 144.800 149.800 145.200 ;
        RECT 148.600 141.800 149.000 142.200 ;
        RECT 146.200 138.800 146.600 139.200 ;
        RECT 147.800 138.800 148.200 139.200 ;
        RECT 145.400 136.800 145.800 137.200 ;
        RECT 144.600 134.800 145.000 135.200 ;
        RECT 145.400 134.200 145.700 136.800 ;
        RECT 147.000 135.800 147.400 136.200 ;
        RECT 147.000 135.200 147.300 135.800 ;
        RECT 147.800 135.200 148.100 138.800 ;
        RECT 148.600 136.200 148.900 141.800 ;
        RECT 149.400 141.200 149.700 144.800 ;
        RECT 151.000 144.200 151.300 145.800 ;
        RECT 151.000 143.800 151.400 144.200 ;
        RECT 149.400 140.800 149.800 141.200 ;
        RECT 150.200 138.800 150.600 139.200 ;
        RECT 148.600 135.800 149.000 136.200 ;
        RECT 150.200 135.200 150.500 138.800 ;
        RECT 151.000 137.200 151.300 143.800 ;
        RECT 151.800 142.200 152.100 153.800 ;
        RECT 152.600 149.200 152.900 164.800 ;
        RECT 153.400 163.200 153.700 165.800 ;
        RECT 154.200 165.200 154.500 165.800 ;
        RECT 154.200 164.800 154.600 165.200 ;
        RECT 153.400 162.800 153.800 163.200 ;
        RECT 154.200 158.100 154.600 158.200 ;
        RECT 155.000 158.100 155.400 158.200 ;
        RECT 154.200 157.800 155.400 158.100 ;
        RECT 156.600 152.100 157.000 157.900 ;
        RECT 157.400 156.800 157.800 157.200 ;
        RECT 153.400 150.800 153.800 151.200 ;
        RECT 152.600 148.800 153.000 149.200 ;
        RECT 151.800 141.800 152.200 142.200 ;
        RECT 152.600 141.800 153.000 142.200 ;
        RECT 151.000 136.800 151.400 137.200 ;
        RECT 147.000 134.800 147.400 135.200 ;
        RECT 147.800 134.800 148.200 135.200 ;
        RECT 150.200 134.800 150.600 135.200 ;
        RECT 152.600 134.200 152.900 141.800 ;
        RECT 153.400 139.200 153.700 150.800 ;
        RECT 157.400 149.200 157.700 156.800 ;
        RECT 158.200 151.200 158.500 165.800 ;
        RECT 159.000 159.200 159.300 171.800 ;
        RECT 160.600 169.100 161.000 169.200 ;
        RECT 161.400 169.100 161.800 169.200 ;
        RECT 160.600 168.800 161.800 169.100 ;
        RECT 164.600 166.200 164.900 176.800 ;
        RECT 167.800 174.800 168.200 175.200 ;
        RECT 167.800 174.200 168.100 174.800 ;
        RECT 167.800 173.800 168.200 174.200 ;
        RECT 168.600 166.800 169.000 167.200 ;
        RECT 168.600 166.200 168.900 166.800 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 162.200 165.800 162.600 166.200 ;
        RECT 163.000 165.800 163.400 166.200 ;
        RECT 163.800 165.800 164.200 166.200 ;
        RECT 164.600 165.800 165.000 166.200 ;
        RECT 167.800 165.800 168.200 166.200 ;
        RECT 168.600 165.800 169.000 166.200 ;
        RECT 169.400 165.800 169.800 166.200 ;
        RECT 159.800 165.200 160.100 165.800 ;
        RECT 159.800 164.800 160.200 165.200 ;
        RECT 162.200 163.200 162.500 165.800 ;
        RECT 162.200 162.800 162.600 163.200 ;
        RECT 163.000 160.200 163.300 165.800 ;
        RECT 163.800 165.200 164.100 165.800 ;
        RECT 163.800 164.800 164.200 165.200 ;
        RECT 165.400 163.100 165.800 163.200 ;
        RECT 166.200 163.100 166.600 163.200 ;
        RECT 165.400 162.800 166.600 163.100 ;
        RECT 163.000 159.800 163.400 160.200 ;
        RECT 159.000 158.800 159.400 159.200 ;
        RECT 159.800 155.000 160.200 155.100 ;
        RECT 160.600 155.000 161.000 155.100 ;
        RECT 159.800 154.700 161.000 155.000 ;
        RECT 159.800 151.800 160.200 152.200 ;
        RECT 161.400 152.100 161.800 157.900 ;
        RECT 165.400 157.800 165.800 158.200 ;
        RECT 163.800 156.100 164.200 156.200 ;
        RECT 164.600 156.100 165.000 156.200 ;
        RECT 162.200 153.800 162.600 154.200 ;
        RECT 158.200 150.800 158.600 151.200 ;
        RECT 159.800 149.200 160.100 151.800 ;
        RECT 157.400 148.800 157.800 149.200 ;
        RECT 159.800 148.800 160.200 149.200 ;
        RECT 162.200 148.200 162.500 153.800 ;
        RECT 163.000 153.100 163.400 155.900 ;
        RECT 163.800 155.800 165.000 156.100 ;
        RECT 165.400 154.200 165.700 157.800 ;
        RECT 166.200 155.100 166.600 155.200 ;
        RECT 167.000 155.100 167.400 155.200 ;
        RECT 166.200 154.800 167.400 155.100 ;
        RECT 165.400 153.800 165.800 154.200 ;
        RECT 167.000 153.800 167.400 154.200 ;
        RECT 164.600 152.800 165.000 153.200 ;
        RECT 164.600 149.200 164.900 152.800 ;
        RECT 164.600 148.800 165.000 149.200 ;
        RECT 154.200 147.800 154.600 148.200 ;
        RECT 162.200 147.800 162.600 148.200 ;
        RECT 154.200 147.200 154.500 147.800 ;
        RECT 167.000 147.200 167.300 153.800 ;
        RECT 167.800 149.200 168.100 165.800 ;
        RECT 169.400 165.200 169.700 165.800 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 169.400 160.800 169.800 161.200 ;
        RECT 168.600 155.800 169.000 156.200 ;
        RECT 168.600 155.200 168.900 155.800 ;
        RECT 168.600 154.800 169.000 155.200 ;
        RECT 169.400 154.200 169.700 160.800 ;
        RECT 169.400 153.800 169.800 154.200 ;
        RECT 170.200 154.100 170.500 185.800 ;
        RECT 171.800 182.800 172.200 183.200 ;
        RECT 171.000 176.800 171.400 177.200 ;
        RECT 171.000 175.200 171.300 176.800 ;
        RECT 171.800 175.200 172.100 182.800 ;
        RECT 175.800 182.200 176.100 185.800 ;
        RECT 173.400 181.800 173.800 182.200 ;
        RECT 175.800 181.800 176.200 182.200 ;
        RECT 171.000 174.800 171.400 175.200 ;
        RECT 171.800 174.800 172.200 175.200 ;
        RECT 171.000 173.800 171.400 174.200 ;
        RECT 171.000 169.200 171.300 173.800 ;
        RECT 171.800 169.200 172.100 174.800 ;
        RECT 172.600 173.100 173.000 175.900 ;
        RECT 171.000 168.800 171.400 169.200 ;
        RECT 171.800 168.800 172.200 169.200 ;
        RECT 171.800 165.800 172.200 166.200 ;
        RECT 172.600 166.100 173.000 166.200 ;
        RECT 173.400 166.100 173.700 181.800 ;
        RECT 176.600 181.200 176.900 185.800 ;
        RECT 178.200 181.800 178.600 182.200 ;
        RECT 176.600 180.800 177.000 181.200 ;
        RECT 174.200 172.100 174.600 177.900 ;
        RECT 175.800 174.800 176.200 175.200 ;
        RECT 175.800 174.200 176.100 174.800 ;
        RECT 175.800 173.800 176.200 174.200 ;
        RECT 175.000 172.800 175.400 173.200 ;
        RECT 177.400 172.800 177.800 173.200 ;
        RECT 175.000 172.200 175.300 172.800 ;
        RECT 175.000 171.800 175.400 172.200 ;
        RECT 175.000 168.800 175.400 169.200 ;
        RECT 175.000 166.200 175.300 168.800 ;
        RECT 177.400 166.200 177.700 172.800 ;
        RECT 178.200 169.200 178.500 181.800 ;
        RECT 179.000 172.100 179.400 177.900 ;
        RECT 179.800 170.200 180.100 185.800 ;
        RECT 182.200 181.800 182.600 182.200 ;
        RECT 181.400 180.800 181.800 181.200 ;
        RECT 181.400 179.200 181.700 180.800 ;
        RECT 181.400 178.800 181.800 179.200 ;
        RECT 182.200 173.200 182.500 181.800 ;
        RECT 183.800 176.200 184.100 185.800 ;
        RECT 184.600 180.200 184.900 194.800 ;
        RECT 185.400 193.800 185.800 194.200 ;
        RECT 185.400 190.200 185.700 193.800 ;
        RECT 185.400 189.800 185.800 190.200 ;
        RECT 185.400 186.800 185.800 187.200 ;
        RECT 185.400 186.200 185.700 186.800 ;
        RECT 185.400 185.800 185.800 186.200 ;
        RECT 184.600 179.800 185.000 180.200 ;
        RECT 185.400 178.800 185.800 179.200 ;
        RECT 183.800 175.800 184.200 176.200 ;
        RECT 183.000 174.800 183.400 175.200 ;
        RECT 182.200 172.800 182.600 173.200 ;
        RECT 181.400 171.800 181.800 172.200 ;
        RECT 182.200 171.800 182.600 172.200 ;
        RECT 179.800 169.800 180.200 170.200 ;
        RECT 178.200 168.800 178.600 169.200 ;
        RECT 179.000 169.100 179.400 169.200 ;
        RECT 179.800 169.100 180.200 169.200 ;
        RECT 179.000 168.800 180.200 169.100 ;
        RECT 181.400 168.100 181.700 171.800 ;
        RECT 182.200 171.200 182.500 171.800 ;
        RECT 182.200 170.800 182.600 171.200 ;
        RECT 183.000 169.200 183.300 174.800 ;
        RECT 184.600 172.100 185.000 177.900 ;
        RECT 185.400 175.200 185.700 178.800 ;
        RECT 186.200 176.200 186.500 194.800 ;
        RECT 187.000 189.800 187.400 190.200 ;
        RECT 187.000 189.200 187.300 189.800 ;
        RECT 187.000 188.800 187.400 189.200 ;
        RECT 188.600 186.200 188.900 200.800 ;
        RECT 195.000 199.200 195.300 205.800 ;
        RECT 197.400 205.200 197.700 210.800 ;
        RECT 203.000 209.200 203.300 214.800 ;
        RECT 203.800 214.200 204.100 226.800 ;
        RECT 203.800 213.800 204.200 214.200 ;
        RECT 203.000 208.800 203.400 209.200 ;
        RECT 199.000 207.100 199.400 207.200 ;
        RECT 199.800 207.100 200.200 207.200 ;
        RECT 199.000 206.800 200.200 207.100 ;
        RECT 204.600 206.200 204.900 228.800 ;
        RECT 207.000 227.800 207.400 228.200 ;
        RECT 207.000 226.300 207.300 227.800 ;
        RECT 207.000 225.900 207.400 226.300 ;
        RECT 207.800 223.100 208.200 228.900 ;
        RECT 210.200 228.800 210.600 229.200 ;
        RECT 210.200 228.200 210.500 228.800 ;
        RECT 208.600 226.800 209.000 227.200 ;
        RECT 208.600 226.200 208.900 226.800 ;
        RECT 208.600 225.800 209.000 226.200 ;
        RECT 209.400 225.100 209.800 227.900 ;
        RECT 210.200 227.800 210.600 228.200 ;
        RECT 214.200 227.200 214.500 233.800 ;
        RECT 220.600 233.200 220.900 233.800 ;
        RECT 220.600 232.800 221.000 233.200 ;
        RECT 215.000 228.800 215.400 229.200 ;
        RECT 215.000 228.200 215.300 228.800 ;
        RECT 215.000 227.800 215.400 228.200 ;
        RECT 214.200 227.100 214.600 227.200 ;
        RECT 214.200 226.800 215.300 227.100 ;
        RECT 213.400 226.100 213.800 226.200 ;
        RECT 214.200 226.100 214.600 226.200 ;
        RECT 213.400 225.800 214.600 226.100 ;
        RECT 205.400 212.800 205.800 213.200 ;
        RECT 205.400 208.200 205.700 212.800 ;
        RECT 206.200 212.100 206.600 217.900 ;
        RECT 207.800 213.100 208.200 215.900 ;
        RECT 208.600 213.800 209.000 214.200 ;
        RECT 208.600 212.200 208.900 213.800 ;
        RECT 210.200 213.100 210.600 215.900 ;
        RECT 207.000 211.800 207.400 212.200 ;
        RECT 208.600 211.800 209.000 212.200 ;
        RECT 211.800 212.100 212.200 217.900 ;
        RECT 212.600 215.800 213.000 216.200 ;
        RECT 212.600 215.100 212.900 215.800 ;
        RECT 215.000 215.200 215.300 226.800 ;
        RECT 215.800 226.800 216.200 227.200 ;
        RECT 215.800 226.200 216.100 226.800 ;
        RECT 215.800 225.800 216.200 226.200 ;
        RECT 216.600 225.800 217.000 226.200 ;
        RECT 212.600 214.700 213.000 215.100 ;
        RECT 215.000 214.800 215.400 215.200 ;
        RECT 213.400 211.800 213.800 212.200 ;
        RECT 205.400 207.800 205.800 208.200 ;
        RECT 205.400 206.200 205.700 207.800 ;
        RECT 199.000 205.800 199.400 206.200 ;
        RECT 200.600 205.800 201.000 206.200 ;
        RECT 201.400 206.100 201.800 206.200 ;
        RECT 202.200 206.100 202.600 206.200 ;
        RECT 201.400 205.800 202.600 206.100 ;
        RECT 204.600 205.800 205.000 206.200 ;
        RECT 205.400 205.800 205.800 206.200 ;
        RECT 197.400 204.800 197.800 205.200 ;
        RECT 197.400 200.200 197.700 204.800 ;
        RECT 199.000 203.200 199.300 205.800 ;
        RECT 200.600 205.200 200.900 205.800 ;
        RECT 200.600 204.800 201.000 205.200 ;
        RECT 199.000 202.800 199.400 203.200 ;
        RECT 202.200 201.800 202.600 202.200 ;
        RECT 197.400 199.800 197.800 200.200 ;
        RECT 199.000 199.800 199.400 200.200 ;
        RECT 195.000 198.800 195.400 199.200 ;
        RECT 190.200 194.800 190.600 195.200 ;
        RECT 190.200 194.200 190.500 194.800 ;
        RECT 190.200 193.800 190.600 194.200 ;
        RECT 191.800 192.800 192.200 193.200 ;
        RECT 191.800 186.200 192.100 192.800 ;
        RECT 195.000 192.100 195.400 197.900 ;
        RECT 197.400 195.100 197.800 195.200 ;
        RECT 198.200 195.100 198.600 195.200 ;
        RECT 197.400 194.800 198.600 195.100 ;
        RECT 196.600 192.800 197.000 193.200 ;
        RECT 192.600 189.800 193.000 190.200 ;
        RECT 188.600 185.800 189.000 186.200 ;
        RECT 189.400 185.800 189.800 186.200 ;
        RECT 191.800 185.800 192.200 186.200 ;
        RECT 188.600 185.200 188.900 185.800 ;
        RECT 188.600 184.800 189.000 185.200 ;
        RECT 186.200 175.800 186.600 176.200 ;
        RECT 185.400 174.800 185.800 175.200 ;
        RECT 187.000 175.100 187.400 175.200 ;
        RECT 187.800 175.100 188.200 175.200 ;
        RECT 187.000 174.800 188.200 175.100 ;
        RECT 184.600 170.800 185.000 171.200 ;
        RECT 183.000 168.800 183.400 169.200 ;
        RECT 180.600 167.800 181.700 168.100 ;
        RECT 184.600 168.200 184.900 170.800 ;
        RECT 184.600 167.800 185.000 168.200 ;
        RECT 187.800 167.800 188.200 168.200 ;
        RECT 172.600 165.800 173.700 166.100 ;
        RECT 174.200 165.800 174.600 166.200 ;
        RECT 175.000 165.800 175.400 166.200 ;
        RECT 176.600 165.800 177.000 166.200 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 171.800 165.200 172.100 165.800 ;
        RECT 174.200 165.200 174.500 165.800 ;
        RECT 176.600 165.200 176.900 165.800 ;
        RECT 171.000 164.800 171.400 165.200 ;
        RECT 171.800 164.800 172.200 165.200 ;
        RECT 174.200 164.800 174.600 165.200 ;
        RECT 176.600 164.800 177.000 165.200 ;
        RECT 177.400 164.800 177.800 165.200 ;
        RECT 171.000 159.200 171.300 164.800 ;
        RECT 171.000 158.800 171.400 159.200 ;
        RECT 175.800 159.100 176.200 159.200 ;
        RECT 176.600 159.100 177.000 159.200 ;
        RECT 175.800 158.800 177.000 159.100 ;
        RECT 177.400 157.200 177.700 164.800 ;
        RECT 179.800 159.200 180.100 165.800 ;
        RECT 180.600 165.200 180.900 167.800 ;
        RECT 187.800 167.200 188.100 167.800 ;
        RECT 182.200 167.100 182.600 167.200 ;
        RECT 183.000 167.100 183.400 167.200 ;
        RECT 182.200 166.800 183.400 167.100 ;
        RECT 186.200 166.800 186.600 167.200 ;
        RECT 187.000 166.800 187.400 167.200 ;
        RECT 187.800 166.800 188.200 167.200 ;
        RECT 186.200 166.200 186.500 166.800 ;
        RECT 187.000 166.200 187.300 166.800 ;
        RECT 181.400 165.800 181.800 166.200 ;
        RECT 186.200 165.800 186.600 166.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 180.600 164.800 181.000 165.200 ;
        RECT 181.400 163.200 181.700 165.800 ;
        RECT 181.400 162.800 181.800 163.200 ;
        RECT 181.400 161.200 181.700 162.800 ;
        RECT 181.400 160.800 181.800 161.200 ;
        RECT 182.200 160.800 182.600 161.200 ;
        RECT 179.800 158.800 180.200 159.200 ;
        RECT 179.000 157.800 179.400 158.200 ;
        RECT 177.400 156.800 177.800 157.200 ;
        RECT 172.600 155.800 173.000 156.200 ;
        RECT 171.000 155.100 171.400 155.200 ;
        RECT 171.800 155.100 172.200 155.200 ;
        RECT 171.000 154.800 172.200 155.100 ;
        RECT 172.600 154.200 172.900 155.800 ;
        RECT 179.000 155.200 179.300 157.800 ;
        RECT 182.200 155.200 182.500 160.800 ;
        RECT 175.800 155.100 176.200 155.200 ;
        RECT 176.600 155.100 177.000 155.200 ;
        RECT 175.800 154.800 177.000 155.100 ;
        RECT 179.000 154.800 179.400 155.200 ;
        RECT 181.400 154.800 181.800 155.200 ;
        RECT 182.200 154.800 182.600 155.200 ;
        RECT 170.200 153.800 171.300 154.100 ;
        RECT 172.600 153.800 173.000 154.200 ;
        RECT 174.200 154.100 174.600 154.200 ;
        RECT 175.000 154.100 175.400 154.200 ;
        RECT 174.200 153.800 175.400 154.100 ;
        RECT 169.400 152.800 169.800 153.200 ;
        RECT 170.200 152.800 170.600 153.200 ;
        RECT 169.400 149.200 169.700 152.800 ;
        RECT 170.200 152.200 170.500 152.800 ;
        RECT 170.200 151.800 170.600 152.200 ;
        RECT 167.800 149.100 168.200 149.200 ;
        RECT 168.600 149.100 169.000 149.200 ;
        RECT 167.800 148.800 169.000 149.100 ;
        RECT 169.400 148.800 169.800 149.200 ;
        RECT 154.200 146.800 154.600 147.200 ;
        RECT 158.200 147.100 158.600 147.200 ;
        RECT 159.000 147.100 159.400 147.200 ;
        RECT 158.200 146.800 159.400 147.100 ;
        RECT 160.600 146.800 161.000 147.200 ;
        RECT 161.400 146.800 161.800 147.200 ;
        RECT 167.000 147.100 167.400 147.200 ;
        RECT 167.800 147.100 168.200 147.200 ;
        RECT 167.000 146.800 168.200 147.100 ;
        RECT 158.200 144.800 158.600 145.200 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 159.800 145.100 160.200 145.200 ;
        RECT 159.000 144.800 160.200 145.100 ;
        RECT 154.200 141.800 154.600 142.200 ;
        RECT 155.000 141.800 155.400 142.200 ;
        RECT 153.400 138.800 153.800 139.200 ;
        RECT 154.200 134.200 154.500 141.800 ;
        RECT 155.000 140.200 155.300 141.800 ;
        RECT 155.000 139.800 155.400 140.200 ;
        RECT 155.800 138.800 156.200 139.200 ;
        RECT 155.800 138.200 156.100 138.800 ;
        RECT 155.000 137.800 155.400 138.200 ;
        RECT 155.800 137.800 156.200 138.200 ;
        RECT 155.000 137.100 155.300 137.800 ;
        RECT 155.000 136.800 156.100 137.100 ;
        RECT 155.000 135.800 155.400 136.200 ;
        RECT 155.000 135.200 155.300 135.800 ;
        RECT 155.000 134.800 155.400 135.200 ;
        RECT 144.600 133.800 145.000 134.200 ;
        RECT 145.400 133.800 145.800 134.200 ;
        RECT 147.800 133.800 148.200 134.200 ;
        RECT 149.400 134.100 149.800 134.200 ;
        RECT 150.200 134.100 150.600 134.200 ;
        RECT 149.400 133.800 150.600 134.100 ;
        RECT 152.600 133.800 153.000 134.200 ;
        RECT 154.200 133.800 154.600 134.200 ;
        RECT 139.800 132.800 140.200 133.200 ;
        RECT 143.000 132.800 143.400 133.200 ;
        RECT 134.200 131.800 134.600 132.200 ;
        RECT 139.000 131.800 139.400 132.200 ;
        RECT 142.200 131.800 142.600 132.200 ;
        RECT 143.000 132.100 143.400 132.200 ;
        RECT 143.800 132.100 144.200 132.200 ;
        RECT 143.000 131.800 144.200 132.100 ;
        RECT 130.200 128.800 130.600 129.200 ;
        RECT 131.000 128.800 131.400 129.200 ;
        RECT 130.200 126.800 130.600 127.200 ;
        RECT 129.400 125.800 129.800 126.200 ;
        RECT 129.400 125.200 129.700 125.800 ;
        RECT 127.800 125.100 128.200 125.200 ;
        RECT 128.600 125.100 129.000 125.200 ;
        RECT 127.800 124.800 129.000 125.100 ;
        RECT 129.400 124.800 129.800 125.200 ;
        RECT 130.200 124.200 130.500 126.800 ;
        RECT 131.800 125.100 132.200 127.900 ;
        RECT 132.600 127.800 133.000 128.200 ;
        RECT 132.600 127.200 132.900 127.800 ;
        RECT 132.600 126.800 133.000 127.200 ;
        RECT 130.200 124.100 130.600 124.200 ;
        RECT 131.000 124.100 131.400 124.200 ;
        RECT 130.200 123.800 131.400 124.100 ;
        RECT 133.400 123.100 133.800 128.900 ;
        RECT 131.000 121.800 131.400 122.200 ;
        RECT 126.200 117.800 126.600 118.200 ;
        RECT 126.200 115.200 126.500 117.800 ;
        RECT 127.800 116.100 128.200 116.200 ;
        RECT 127.000 115.800 128.200 116.100 ;
        RECT 129.400 115.800 129.800 116.200 ;
        RECT 126.200 114.800 126.600 115.200 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 124.600 113.800 125.800 114.100 ;
        RECT 124.600 109.200 124.900 113.800 ;
        RECT 124.600 108.800 125.000 109.200 ;
        RECT 123.000 106.800 123.400 107.200 ;
        RECT 124.600 106.200 124.900 108.800 ;
        RECT 126.200 107.100 126.500 114.800 ;
        RECT 127.000 109.200 127.300 115.800 ;
        RECT 129.400 115.200 129.700 115.800 ;
        RECT 127.800 115.100 128.200 115.200 ;
        RECT 128.600 115.100 129.000 115.200 ;
        RECT 127.800 114.800 129.000 115.100 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 127.800 114.100 128.200 114.200 ;
        RECT 128.600 114.100 129.000 114.200 ;
        RECT 127.800 113.800 129.000 114.100 ;
        RECT 128.600 110.800 129.000 111.200 ;
        RECT 127.000 108.800 127.400 109.200 ;
        RECT 128.600 107.200 128.900 110.800 ;
        RECT 126.200 106.800 127.300 107.100 ;
        RECT 124.600 105.800 125.000 106.200 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 126.200 105.200 126.500 105.800 ;
        RECT 127.000 105.200 127.300 106.800 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 126.200 104.800 126.600 105.200 ;
        RECT 127.000 104.800 127.400 105.200 ;
        RECT 117.400 101.800 117.800 102.200 ;
        RECT 125.400 101.800 125.800 102.200 ;
        RECT 117.400 100.200 117.700 101.800 ;
        RECT 124.600 100.800 125.000 101.200 ;
        RECT 117.400 99.800 117.800 100.200 ;
        RECT 117.400 92.100 117.800 97.900 ;
        RECT 118.200 94.700 118.600 95.100 ;
        RECT 118.200 94.200 118.500 94.700 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 119.800 93.800 120.200 94.200 ;
        RECT 119.800 93.200 120.100 93.800 ;
        RECT 119.800 92.800 120.200 93.200 ;
        RECT 119.000 91.800 119.400 92.200 ;
        RECT 119.000 88.200 119.300 91.800 ;
        RECT 119.800 91.200 120.100 92.800 ;
        RECT 122.200 92.100 122.600 97.900 ;
        RECT 124.600 97.200 124.900 100.800 ;
        RECT 123.800 97.100 124.200 97.200 ;
        RECT 124.600 97.100 125.000 97.200 ;
        RECT 123.800 96.800 125.000 97.100 ;
        RECT 125.400 93.200 125.700 101.800 ;
        RECT 126.200 97.200 126.500 104.800 ;
        RECT 127.000 103.800 127.400 104.200 ;
        RECT 126.200 96.800 126.600 97.200 ;
        RECT 127.000 95.200 127.300 103.800 ;
        RECT 127.800 99.800 128.200 100.200 ;
        RECT 127.000 94.800 127.400 95.200 ;
        RECT 125.400 92.800 125.800 93.200 ;
        RECT 119.800 90.800 120.200 91.200 ;
        RECT 119.000 87.800 119.400 88.200 ;
        RECT 119.800 86.200 120.100 90.800 ;
        RECT 123.800 88.800 124.200 89.200 ;
        RECT 120.600 87.100 121.000 87.200 ;
        RECT 121.400 87.100 121.800 87.200 ;
        RECT 120.600 86.800 121.800 87.100 ;
        RECT 123.800 86.200 124.100 88.800 ;
        RECT 124.600 86.800 125.000 87.200 ;
        RECT 124.600 86.200 124.900 86.800 ;
        RECT 119.800 85.800 120.200 86.200 ;
        RECT 121.400 85.800 121.800 86.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 124.600 85.800 125.000 86.200 ;
        RECT 121.400 79.200 121.700 85.800 ;
        RECT 125.400 85.100 125.800 87.900 ;
        RECT 127.000 83.100 127.400 88.900 ;
        RECT 127.800 88.200 128.100 99.800 ;
        RECT 128.600 98.200 128.900 106.800 ;
        RECT 129.400 105.800 129.800 106.200 ;
        RECT 130.200 105.800 130.600 106.200 ;
        RECT 129.400 99.200 129.700 105.800 ;
        RECT 130.200 101.200 130.500 105.800 ;
        RECT 131.000 101.200 131.300 121.800 ;
        RECT 133.400 118.800 133.800 119.200 ;
        RECT 131.800 116.100 132.200 116.200 ;
        RECT 132.600 116.100 133.000 116.200 ;
        RECT 131.800 115.800 133.000 116.100 ;
        RECT 131.800 115.200 132.100 115.800 ;
        RECT 131.800 114.800 132.200 115.200 ;
        RECT 132.600 114.800 133.000 115.200 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 132.600 114.100 132.900 114.800 ;
        RECT 131.800 113.800 132.900 114.100 ;
        RECT 133.400 114.200 133.700 118.800 ;
        RECT 134.200 117.100 134.500 131.800 ;
        RECT 135.000 126.100 135.400 126.200 ;
        RECT 135.800 126.100 136.200 126.200 ;
        RECT 135.000 125.800 136.200 126.100 ;
        RECT 138.200 123.100 138.600 128.900 ;
        RECT 136.600 118.800 137.000 119.200 ;
        RECT 135.000 117.100 135.400 117.200 ;
        RECT 134.200 116.800 135.400 117.100 ;
        RECT 133.400 113.800 133.800 114.200 ;
        RECT 134.200 113.100 134.600 115.900 ;
        RECT 135.800 112.100 136.200 117.900 ;
        RECT 136.600 117.200 136.900 118.800 ;
        RECT 136.600 116.800 137.000 117.200 ;
        RECT 137.400 115.100 137.800 115.200 ;
        RECT 136.600 114.800 137.800 115.100 ;
        RECT 136.600 114.700 137.000 114.800 ;
        RECT 138.200 113.800 138.600 114.200 ;
        RECT 138.200 110.200 138.500 113.800 ;
        RECT 138.200 109.800 138.600 110.200 ;
        RECT 132.600 106.800 133.000 107.200 ;
        RECT 134.200 106.800 134.600 107.200 ;
        RECT 138.200 106.800 138.600 107.200 ;
        RECT 132.600 106.200 132.900 106.800 ;
        RECT 134.200 106.200 134.500 106.800 ;
        RECT 138.200 106.200 138.500 106.800 ;
        RECT 131.800 105.800 132.200 106.200 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 135.000 105.800 135.400 106.200 ;
        RECT 137.400 105.800 137.800 106.200 ;
        RECT 138.200 105.800 138.600 106.200 ;
        RECT 131.800 105.200 132.100 105.800 ;
        RECT 135.000 105.200 135.300 105.800 ;
        RECT 131.800 104.800 132.200 105.200 ;
        RECT 135.000 104.800 135.400 105.200 ;
        RECT 137.400 104.200 137.700 105.800 ;
        RECT 131.800 103.800 132.200 104.200 ;
        RECT 137.400 103.800 137.800 104.200 ;
        RECT 130.200 100.800 130.600 101.200 ;
        RECT 131.000 100.800 131.400 101.200 ;
        RECT 129.400 98.800 129.800 99.200 ;
        RECT 128.600 97.800 129.000 98.200 ;
        RECT 128.600 95.800 129.000 96.200 ;
        RECT 128.600 95.200 128.900 95.800 ;
        RECT 128.600 94.800 129.000 95.200 ;
        RECT 129.400 94.800 129.800 95.200 ;
        RECT 130.200 94.800 130.600 95.200 ;
        RECT 127.800 87.800 128.200 88.200 ;
        RECT 128.600 86.800 129.000 87.200 ;
        RECT 128.600 86.200 128.900 86.800 ;
        RECT 128.600 85.800 129.000 86.200 ;
        RECT 129.400 85.200 129.700 94.800 ;
        RECT 130.200 92.200 130.500 94.800 ;
        RECT 130.200 91.800 130.600 92.200 ;
        RECT 129.400 84.800 129.800 85.200 ;
        RECT 127.000 79.800 127.400 80.200 ;
        RECT 121.400 78.800 121.800 79.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 117.400 72.100 117.800 77.900 ;
        RECT 127.000 75.200 127.300 79.800 ;
        RECT 127.800 77.100 128.200 77.200 ;
        RECT 128.600 77.100 129.000 77.200 ;
        RECT 127.800 76.800 129.000 77.100 ;
        RECT 129.400 75.800 129.800 76.200 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 127.000 73.800 127.400 74.200 ;
        RECT 119.000 72.800 119.400 73.200 ;
        RECT 119.000 72.100 119.300 72.800 ;
        RECT 119.800 72.100 120.200 72.200 ;
        RECT 119.000 71.800 120.200 72.100 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 117.400 66.200 117.700 66.800 ;
        RECT 119.000 66.200 119.300 71.800 ;
        RECT 124.600 69.200 124.900 73.800 ;
        RECT 127.000 73.200 127.300 73.800 ;
        RECT 127.000 72.800 127.400 73.200 ;
        RECT 129.400 72.100 129.700 75.800 ;
        RECT 130.200 73.100 130.600 75.900 ;
        RECT 129.400 71.800 130.500 72.100 ;
        RECT 130.200 69.200 130.500 71.800 ;
        RECT 124.600 68.800 125.000 69.200 ;
        RECT 129.400 68.800 129.800 69.200 ;
        RECT 130.200 68.800 130.600 69.200 ;
        RECT 128.600 67.800 129.000 68.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 122.200 67.100 122.600 67.200 ;
        RECT 121.400 66.800 122.600 67.100 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 125.400 67.100 125.800 67.200 ;
        RECT 126.200 67.100 126.600 67.200 ;
        RECT 125.400 66.800 126.600 67.100 ;
        RECT 127.000 67.100 127.400 67.200 ;
        RECT 127.800 67.100 128.200 67.200 ;
        RECT 127.000 66.800 128.200 67.100 ;
        RECT 116.600 66.100 117.000 66.200 ;
        RECT 115.800 65.800 117.000 66.100 ;
        RECT 117.400 65.800 117.800 66.200 ;
        RECT 118.200 65.800 118.600 66.200 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 121.400 65.800 121.800 66.200 ;
        RECT 115.000 54.800 115.400 55.200 ;
        RECT 115.000 54.200 115.300 54.800 ;
        RECT 113.400 53.800 113.800 54.200 ;
        RECT 115.000 53.800 115.400 54.200 ;
        RECT 112.600 53.100 113.000 53.200 ;
        RECT 113.400 53.100 113.800 53.200 ;
        RECT 112.600 52.800 113.800 53.100 ;
        RECT 111.800 44.800 112.200 45.200 ;
        RECT 112.600 45.100 113.000 47.900 ;
        RECT 113.400 45.100 113.800 47.900 ;
        RECT 114.200 46.800 114.600 47.200 ;
        RECT 111.800 43.800 112.200 44.200 ;
        RECT 111.800 39.200 112.100 43.800 ;
        RECT 111.800 38.800 112.200 39.200 ;
        RECT 110.200 36.800 110.600 37.200 ;
        RECT 104.600 35.800 105.000 36.200 ;
        RECT 110.200 35.200 110.500 36.800 ;
        RECT 101.400 34.800 101.800 35.200 ;
        RECT 109.400 34.800 109.800 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 97.400 28.800 97.800 29.200 ;
        RECT 99.000 28.800 99.400 29.200 ;
        RECT 96.600 18.800 97.000 19.200 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 93.400 14.800 93.800 15.200 ;
        RECT 95.800 14.800 96.200 15.200 ;
        RECT 87.800 12.800 88.200 13.200 ;
        RECT 91.000 9.800 91.400 10.200 ;
        RECT 87.000 6.800 87.400 7.200 ;
        RECT 87.800 6.800 88.200 7.200 ;
        RECT 87.800 6.300 88.100 6.800 ;
        RECT 87.800 5.900 88.200 6.300 ;
        RECT 88.600 3.100 89.000 8.900 ;
        RECT 90.200 5.100 90.600 7.900 ;
        RECT 91.000 7.200 91.300 9.800 ;
        RECT 92.600 9.200 92.900 14.800 ;
        RECT 93.400 11.200 93.700 14.800 ;
        RECT 96.600 12.100 97.000 17.900 ;
        RECT 97.400 15.200 97.700 28.800 ;
        RECT 101.400 27.200 101.700 34.800 ;
        RECT 103.000 33.800 103.400 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 104.600 33.800 105.800 34.100 ;
        RECT 103.000 33.200 103.300 33.800 ;
        RECT 103.000 32.800 103.400 33.200 ;
        RECT 107.800 28.800 108.200 29.200 ;
        RECT 107.800 27.200 108.100 28.800 ;
        RECT 101.400 26.800 101.800 27.200 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 107.800 26.800 108.200 27.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 100.600 25.800 101.000 26.200 ;
        RECT 97.400 14.800 97.800 15.200 ;
        RECT 97.400 12.200 97.700 14.800 ;
        RECT 98.200 12.200 98.500 25.800 ;
        RECT 100.600 18.200 100.900 25.800 ;
        RECT 101.400 20.200 101.700 26.800 ;
        RECT 104.600 26.200 104.900 26.800 ;
        RECT 102.200 25.800 102.600 26.200 ;
        RECT 104.600 25.800 105.000 26.200 ;
        RECT 102.200 25.200 102.500 25.800 ;
        RECT 102.200 24.800 102.600 25.200 ;
        RECT 103.800 25.100 104.200 25.200 ;
        RECT 104.600 25.100 105.000 25.200 ;
        RECT 103.800 24.800 105.000 25.100 ;
        RECT 101.400 19.800 101.800 20.200 ;
        RECT 100.600 17.800 101.000 18.200 ;
        RECT 100.600 17.200 100.900 17.800 ;
        RECT 100.600 16.800 101.000 17.200 ;
        RECT 99.000 15.100 99.400 15.200 ;
        RECT 99.800 15.100 100.200 15.200 ;
        RECT 99.000 14.800 100.200 15.100 ;
        RECT 97.400 11.800 97.800 12.200 ;
        RECT 98.200 11.800 98.600 12.200 ;
        RECT 101.400 12.100 101.800 17.900 ;
        RECT 93.400 10.800 93.800 11.200 ;
        RECT 92.600 8.800 93.000 9.200 ;
        RECT 95.800 8.800 96.200 9.200 ;
        RECT 95.800 7.200 96.100 8.800 ;
        RECT 91.000 6.800 91.400 7.200 ;
        RECT 92.600 7.100 93.000 7.200 ;
        RECT 93.400 7.100 93.800 7.200 ;
        RECT 92.600 6.800 93.800 7.100 ;
        RECT 95.800 6.800 96.200 7.200 ;
        RECT 92.600 5.800 93.000 6.200 ;
        RECT 94.200 6.100 94.600 6.200 ;
        RECT 95.000 6.100 95.400 6.200 ;
        RECT 94.200 5.800 95.400 6.100 ;
        RECT 92.600 5.200 92.900 5.800 ;
        RECT 92.600 4.800 93.000 5.200 ;
        RECT 96.600 5.100 97.000 7.900 ;
        RECT 97.400 7.800 97.800 8.200 ;
        RECT 97.400 7.200 97.700 7.800 ;
        RECT 97.400 6.800 97.800 7.200 ;
        RECT 98.200 3.100 98.600 8.900 ;
        RECT 101.400 6.800 101.800 7.200 ;
        RECT 101.400 6.200 101.700 6.800 ;
        RECT 102.200 6.200 102.500 24.800 ;
        RECT 109.400 24.200 109.700 34.800 ;
        RECT 114.200 29.200 114.500 46.800 ;
        RECT 115.000 43.100 115.400 48.900 ;
        RECT 115.800 40.200 116.100 65.800 ;
        RECT 118.200 65.200 118.500 65.800 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 121.400 64.200 121.700 65.800 ;
        RECT 121.400 63.800 121.800 64.200 ;
        RECT 123.000 63.200 123.300 66.800 ;
        RECT 128.600 66.200 128.900 67.800 ;
        RECT 129.400 67.200 129.700 68.800 ;
        RECT 129.400 66.800 129.800 67.200 ;
        RECT 125.400 66.100 125.800 66.200 ;
        RECT 126.200 66.100 126.600 66.200 ;
        RECT 125.400 65.800 126.600 66.100 ;
        RECT 128.600 65.800 129.000 66.200 ;
        RECT 129.400 66.100 129.800 66.200 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 129.400 65.800 130.600 66.100 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 124.600 64.200 124.900 64.800 ;
        RECT 124.600 63.800 125.000 64.200 ;
        RECT 126.200 63.800 126.600 64.200 ;
        RECT 126.200 63.200 126.500 63.800 ;
        RECT 123.000 62.800 123.400 63.200 ;
        RECT 126.200 62.800 126.600 63.200 ;
        RECT 131.000 61.200 131.300 100.800 ;
        RECT 131.800 99.200 132.100 103.800 ;
        RECT 131.800 98.800 132.200 99.200 ;
        RECT 132.600 97.800 133.000 98.200 ;
        RECT 137.400 97.800 137.800 98.200 ;
        RECT 132.600 95.200 132.900 97.800 ;
        RECT 134.200 96.800 134.600 97.200 ;
        RECT 134.200 95.200 134.500 96.800 ;
        RECT 137.400 95.200 137.700 97.800 ;
        RECT 139.000 96.200 139.300 131.800 ;
        RECT 140.600 129.100 141.000 129.200 ;
        RECT 141.400 129.100 141.800 129.200 ;
        RECT 140.600 128.800 141.800 129.100 ;
        RECT 142.200 128.200 142.500 131.800 ;
        RECT 144.600 131.200 144.900 133.800 ;
        RECT 147.800 133.200 148.100 133.800 ;
        RECT 147.800 132.800 148.200 133.200 ;
        RECT 149.400 133.100 149.800 133.200 ;
        RECT 150.200 133.100 150.600 133.200 ;
        RECT 149.400 132.800 150.600 133.100 ;
        RECT 151.800 132.800 152.200 133.200 ;
        RECT 144.600 130.800 145.000 131.200 ;
        RECT 146.200 128.800 146.600 129.200 ;
        RECT 147.800 128.800 148.200 129.200 ;
        RECT 142.200 127.800 142.600 128.200 ;
        RECT 144.600 127.800 145.000 128.200 ;
        RECT 145.400 127.800 145.800 128.200 ;
        RECT 141.400 126.800 141.800 127.200 ;
        RECT 139.800 112.800 140.200 113.200 ;
        RECT 139.800 109.200 140.100 112.800 ;
        RECT 140.600 112.100 141.000 117.900 ;
        RECT 141.400 114.200 141.700 126.800 ;
        RECT 142.200 126.200 142.500 127.800 ;
        RECT 142.200 125.800 142.600 126.200 ;
        RECT 143.000 126.100 143.400 126.200 ;
        RECT 143.800 126.100 144.200 126.200 ;
        RECT 143.000 125.800 144.200 126.100 ;
        RECT 144.600 125.200 144.900 127.800 ;
        RECT 144.600 124.800 145.000 125.200 ;
        RECT 143.000 117.100 143.400 117.200 ;
        RECT 143.800 117.100 144.200 117.200 ;
        RECT 143.000 116.800 144.200 117.100 ;
        RECT 144.600 114.200 144.900 124.800 ;
        RECT 145.400 115.200 145.700 127.800 ;
        RECT 146.200 127.200 146.500 128.800 ;
        RECT 146.200 126.800 146.600 127.200 ;
        RECT 147.800 126.200 148.100 128.800 ;
        RECT 151.800 127.200 152.100 132.800 ;
        RECT 154.200 128.200 154.500 133.800 ;
        RECT 155.000 131.800 155.400 132.200 ;
        RECT 155.000 129.200 155.300 131.800 ;
        RECT 155.000 128.800 155.400 129.200 ;
        RECT 154.200 127.800 154.600 128.200 ;
        RECT 150.200 126.800 150.600 127.200 ;
        RECT 151.800 126.800 152.200 127.200 ;
        RECT 150.200 126.200 150.500 126.800 ;
        RECT 155.800 126.200 156.100 136.800 ;
        RECT 158.200 136.200 158.500 144.800 ;
        RECT 159.800 142.800 160.200 143.200 ;
        RECT 159.800 139.200 160.100 142.800 ;
        RECT 159.800 138.800 160.200 139.200 ;
        RECT 158.200 135.800 158.600 136.200 ;
        RECT 156.600 133.800 157.000 134.200 ;
        RECT 156.600 133.200 156.900 133.800 ;
        RECT 156.600 132.800 157.000 133.200 ;
        RECT 157.400 129.800 157.800 130.200 ;
        RECT 157.400 127.200 157.700 129.800 ;
        RECT 158.200 129.200 158.500 135.800 ;
        RECT 160.600 135.200 160.900 146.800 ;
        RECT 161.400 146.200 161.700 146.800 ;
        RECT 161.400 145.800 161.800 146.200 ;
        RECT 163.000 145.800 163.400 146.200 ;
        RECT 163.000 145.200 163.300 145.800 ;
        RECT 163.000 144.800 163.400 145.200 ;
        RECT 161.400 143.800 161.800 144.200 ;
        RECT 162.200 143.800 162.600 144.200 ;
        RECT 161.400 142.200 161.700 143.800 ;
        RECT 162.200 143.200 162.500 143.800 ;
        RECT 162.200 142.800 162.600 143.200 ;
        RECT 170.200 143.100 170.600 148.900 ;
        RECT 171.000 143.200 171.300 153.800 ;
        RECT 175.000 153.200 175.300 153.800 ;
        RECT 173.400 153.100 173.800 153.200 ;
        RECT 174.200 153.100 174.600 153.200 ;
        RECT 173.400 152.800 174.600 153.100 ;
        RECT 175.000 152.800 175.400 153.200 ;
        RECT 173.400 151.800 173.800 152.200 ;
        RECT 173.400 146.200 173.700 151.800 ;
        RECT 181.400 150.200 181.700 154.800 ;
        RECT 181.400 149.800 181.800 150.200 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 173.400 145.800 173.800 146.200 ;
        RECT 172.600 143.800 173.000 144.200 ;
        RECT 171.000 142.800 171.400 143.200 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 166.200 141.800 166.600 142.200 ;
        RECT 165.400 138.800 165.800 139.200 ;
        RECT 163.800 136.100 164.200 136.200 ;
        RECT 164.600 136.100 165.000 136.200 ;
        RECT 163.800 135.800 165.000 136.100 ;
        RECT 160.600 134.800 161.000 135.200 ;
        RECT 163.800 134.800 164.200 135.200 ;
        RECT 160.600 133.800 161.000 134.200 ;
        RECT 160.600 133.200 160.900 133.800 ;
        RECT 160.600 132.800 161.000 133.200 ;
        RECT 161.400 133.100 161.800 133.200 ;
        RECT 162.200 133.100 162.600 133.200 ;
        RECT 161.400 132.800 162.600 133.100 ;
        RECT 159.800 131.800 160.200 132.200 ;
        RECT 159.000 130.800 159.400 131.200 ;
        RECT 159.000 129.200 159.300 130.800 ;
        RECT 158.200 128.800 158.600 129.200 ;
        RECT 159.000 128.800 159.400 129.200 ;
        RECT 157.400 127.100 157.800 127.200 ;
        RECT 158.200 127.100 158.600 127.200 ;
        RECT 157.400 126.800 158.600 127.100 ;
        RECT 146.200 126.100 146.600 126.200 ;
        RECT 147.000 126.100 147.400 126.200 ;
        RECT 146.200 125.800 147.400 126.100 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 152.600 125.800 153.000 126.200 ;
        RECT 155.000 125.800 155.400 126.200 ;
        RECT 155.800 125.800 156.200 126.200 ;
        RECT 158.200 125.800 158.600 126.200 ;
        RECT 147.000 122.800 147.400 123.200 ;
        RECT 147.000 116.200 147.300 122.800 ;
        RECT 149.400 121.800 149.800 122.200 ;
        RECT 147.800 119.100 148.200 119.200 ;
        RECT 148.600 119.100 149.000 119.200 ;
        RECT 147.800 118.800 149.000 119.100 ;
        RECT 149.400 118.200 149.700 121.800 ;
        RECT 152.600 119.200 152.900 125.800 ;
        RECT 153.400 125.100 153.800 125.200 ;
        RECT 154.200 125.100 154.600 125.200 ;
        RECT 153.400 124.800 154.600 125.100 ;
        RECT 152.600 118.800 153.000 119.200 ;
        RECT 149.400 117.800 149.800 118.200 ;
        RECT 154.200 117.800 154.600 118.200 ;
        RECT 151.800 116.800 152.200 117.200 ;
        RECT 147.000 115.800 147.400 116.200 ;
        RECT 151.800 115.200 152.100 116.800 ;
        RECT 145.400 114.800 145.800 115.200 ;
        RECT 148.600 115.100 149.000 115.200 ;
        RECT 149.400 115.100 149.800 115.200 ;
        RECT 148.600 114.800 149.800 115.100 ;
        RECT 150.200 115.100 150.600 115.200 ;
        RECT 151.000 115.100 151.400 115.200 ;
        RECT 150.200 114.800 151.400 115.100 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 141.400 113.800 141.800 114.200 ;
        RECT 143.800 113.800 144.200 114.200 ;
        RECT 144.600 113.800 145.000 114.200 ;
        RECT 139.800 108.800 140.200 109.200 ;
        RECT 141.400 98.200 141.700 113.800 ;
        RECT 143.800 113.200 144.100 113.800 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 143.800 111.800 144.200 112.200 ;
        RECT 144.600 111.800 145.000 112.200 ;
        RECT 143.800 109.200 144.100 111.800 ;
        RECT 143.800 108.800 144.200 109.200 ;
        RECT 144.600 107.200 144.900 111.800 ;
        RECT 143.000 106.800 143.400 107.200 ;
        RECT 144.600 106.800 145.000 107.200 ;
        RECT 143.000 105.200 143.300 106.800 ;
        RECT 144.600 106.100 145.000 106.200 ;
        RECT 145.400 106.100 145.700 114.800 ;
        RECT 146.200 113.100 146.600 113.200 ;
        RECT 147.000 113.100 147.400 113.200 ;
        RECT 146.200 112.800 147.400 113.100 ;
        RECT 150.200 112.800 150.600 113.200 ;
        RECT 147.000 107.200 147.300 112.800 ;
        RECT 150.200 112.200 150.500 112.800 ;
        RECT 150.200 111.800 150.600 112.200 ;
        RECT 150.200 108.200 150.500 111.800 ;
        RECT 148.600 107.800 149.000 108.200 ;
        RECT 150.200 107.800 150.600 108.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 148.600 106.200 148.900 107.800 ;
        RECT 144.600 105.800 146.500 106.100 ;
        RECT 148.600 105.800 149.000 106.200 ;
        RECT 150.200 105.800 150.600 106.200 ;
        RECT 143.000 104.800 143.400 105.200 ;
        RECT 144.600 105.100 145.000 105.200 ;
        RECT 145.400 105.100 145.800 105.200 ;
        RECT 144.600 104.800 145.800 105.100 ;
        RECT 145.400 102.800 145.800 103.200 ;
        RECT 145.400 100.200 145.700 102.800 ;
        RECT 145.400 99.800 145.800 100.200 ;
        RECT 141.400 97.800 141.800 98.200 ;
        RECT 139.000 95.800 139.400 96.200 ;
        RECT 132.600 94.800 133.000 95.200 ;
        RECT 134.200 94.800 134.600 95.200 ;
        RECT 137.400 94.800 137.800 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 139.800 95.100 140.200 95.200 ;
        RECT 139.000 94.800 140.200 95.100 ;
        RECT 138.200 93.800 138.600 94.200 ;
        RECT 139.800 93.800 140.200 94.200 ;
        RECT 138.200 93.200 138.500 93.800 ;
        RECT 139.800 93.200 140.100 93.800 ;
        RECT 138.200 92.800 138.600 93.200 ;
        RECT 139.800 92.800 140.200 93.200 ;
        RECT 140.600 93.100 141.000 95.900 ;
        RECT 141.400 95.800 141.800 96.200 ;
        RECT 135.800 91.800 136.200 92.200 ;
        RECT 135.800 89.200 136.100 91.800 ;
        RECT 138.200 90.200 138.500 92.800 ;
        RECT 138.200 89.800 138.600 90.200 ;
        RECT 131.800 83.100 132.200 88.900 ;
        RECT 135.800 88.800 136.200 89.200 ;
        RECT 135.000 87.800 135.400 88.200 ;
        RECT 135.000 87.200 135.300 87.800 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 135.800 86.200 136.100 88.800 ;
        RECT 136.600 87.100 137.000 87.200 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 136.600 86.800 137.800 87.100 ;
        RECT 141.400 86.200 141.700 95.800 ;
        RECT 142.200 92.100 142.600 97.900 ;
        RECT 143.800 95.100 144.200 95.200 ;
        RECT 143.000 94.800 144.200 95.100 ;
        RECT 143.000 94.700 143.400 94.800 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 143.000 91.200 143.300 92.800 ;
        RECT 143.000 90.800 143.400 91.200 ;
        RECT 144.600 87.800 145.000 88.200 ;
        RECT 144.600 86.200 144.900 87.800 ;
        RECT 145.400 86.200 145.700 99.800 ;
        RECT 146.200 88.200 146.500 105.800 ;
        RECT 148.600 102.100 149.000 102.200 ;
        RECT 149.400 102.100 149.800 102.200 ;
        RECT 148.600 101.800 149.800 102.100 ;
        RECT 147.000 92.100 147.400 97.900 ;
        RECT 150.200 97.200 150.500 105.800 ;
        RECT 151.000 100.200 151.300 114.800 ;
        RECT 152.600 110.800 153.000 111.200 ;
        RECT 152.600 109.200 152.900 110.800 ;
        RECT 152.600 108.800 153.000 109.200 ;
        RECT 154.200 106.200 154.500 117.800 ;
        RECT 154.200 105.800 154.600 106.200 ;
        RECT 154.200 100.800 154.600 101.200 ;
        RECT 151.000 99.800 151.400 100.200 ;
        RECT 149.400 96.800 149.800 97.200 ;
        RECT 150.200 96.800 150.600 97.200 ;
        RECT 151.000 96.800 151.400 97.200 ;
        RECT 149.400 95.100 149.700 96.800 ;
        RECT 151.000 96.200 151.300 96.800 ;
        RECT 154.200 96.200 154.500 100.800 ;
        RECT 155.000 99.200 155.300 125.800 ;
        RECT 155.800 116.800 156.200 117.200 ;
        RECT 155.800 114.200 156.100 116.800 ;
        RECT 156.600 116.100 157.000 116.200 ;
        RECT 157.400 116.100 157.800 116.200 ;
        RECT 156.600 115.800 157.800 116.100 ;
        RECT 155.800 113.800 156.200 114.200 ;
        RECT 155.800 105.800 156.200 106.200 ;
        RECT 157.400 105.800 157.800 106.200 ;
        RECT 155.800 105.200 156.100 105.800 ;
        RECT 155.800 104.800 156.200 105.200 ;
        RECT 157.400 102.200 157.700 105.800 ;
        RECT 157.400 101.800 157.800 102.200 ;
        RECT 155.000 98.800 155.400 99.200 ;
        RECT 151.000 95.800 151.400 96.200 ;
        RECT 154.200 95.800 154.600 96.200 ;
        RECT 158.200 95.200 158.500 125.800 ;
        RECT 159.800 124.200 160.100 131.800 ;
        RECT 160.600 131.200 160.900 132.800 ;
        RECT 160.600 130.800 161.000 131.200 ;
        RECT 162.200 129.100 162.600 129.200 ;
        RECT 163.000 129.100 163.400 129.200 ;
        RECT 162.200 128.800 163.400 129.100 ;
        RECT 163.800 126.200 164.100 134.800 ;
        RECT 165.400 134.200 165.700 138.800 ;
        RECT 166.200 135.200 166.500 141.800 ;
        RECT 168.600 140.800 169.000 141.200 ;
        RECT 168.600 139.200 168.900 140.800 ;
        RECT 167.800 138.800 168.200 139.200 ;
        RECT 168.600 138.800 169.000 139.200 ;
        RECT 167.800 135.200 168.100 138.800 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 167.800 134.800 168.200 135.200 ;
        RECT 166.200 134.200 166.500 134.800 ;
        RECT 165.400 133.800 165.800 134.200 ;
        RECT 166.200 133.800 166.600 134.200 ;
        RECT 164.600 132.800 165.000 133.200 ;
        RECT 166.200 133.100 166.600 133.200 ;
        RECT 167.000 133.100 167.400 133.200 ;
        RECT 166.200 132.800 167.400 133.100 ;
        RECT 164.600 130.200 164.900 132.800 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 171.000 132.100 171.400 137.900 ;
        RECT 171.800 133.800 172.200 134.200 ;
        RECT 167.000 131.200 167.300 131.800 ;
        RECT 167.000 130.800 167.400 131.200 ;
        RECT 164.600 129.800 165.000 130.200 ;
        RECT 171.800 129.200 172.100 133.800 ;
        RECT 165.400 128.800 165.800 129.200 ;
        RECT 170.200 128.800 170.600 129.200 ;
        RECT 171.800 128.800 172.200 129.200 ;
        RECT 165.400 128.200 165.700 128.800 ;
        RECT 165.400 127.800 165.800 128.200 ;
        RECT 169.400 127.800 169.800 128.200 ;
        RECT 164.600 126.800 165.000 127.200 ;
        RECT 165.400 126.800 165.800 127.200 ;
        RECT 167.000 127.100 167.400 127.200 ;
        RECT 166.200 126.800 167.400 127.100 ;
        RECT 164.600 126.200 164.900 126.800 ;
        RECT 165.400 126.200 165.700 126.800 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 164.600 125.800 165.000 126.200 ;
        RECT 165.400 125.800 165.800 126.200 ;
        RECT 159.800 123.800 160.200 124.200 ;
        RECT 160.600 122.800 161.000 123.200 ;
        RECT 160.600 122.200 160.900 122.800 ;
        RECT 160.600 121.800 161.000 122.200 ;
        RECT 162.200 117.100 162.600 117.200 ;
        RECT 163.000 117.100 163.400 117.200 ;
        RECT 162.200 116.800 163.400 117.100 ;
        RECT 161.400 115.800 161.800 116.200 ;
        RECT 161.400 115.200 161.700 115.800 ;
        RECT 161.400 114.800 161.800 115.200 ;
        RECT 159.800 114.100 160.200 114.200 ;
        RECT 160.600 114.100 161.000 114.200 ;
        RECT 159.800 113.800 161.000 114.100 ;
        RECT 162.200 113.800 162.600 114.200 ;
        RECT 162.200 111.200 162.500 113.800 ;
        RECT 162.200 110.800 162.600 111.200 ;
        RECT 160.600 107.100 161.000 107.200 ;
        RECT 161.400 107.100 161.800 107.200 ;
        RECT 160.600 106.800 161.800 107.100 ;
        RECT 159.000 105.800 159.400 106.200 ;
        RECT 159.800 106.100 160.200 106.200 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 159.800 105.800 161.000 106.100 ;
        RECT 159.000 104.200 159.300 105.800 ;
        RECT 159.000 103.800 159.400 104.200 ;
        RECT 159.800 96.100 160.200 96.200 ;
        RECT 160.600 96.100 161.000 96.200 ;
        RECT 159.800 95.800 161.000 96.100 ;
        RECT 150.200 95.100 150.600 95.200 ;
        RECT 149.400 94.800 150.600 95.100 ;
        RECT 151.800 94.800 152.200 95.200 ;
        RECT 152.600 94.800 153.000 95.200 ;
        RECT 155.800 95.100 156.200 95.200 ;
        RECT 156.600 95.100 157.000 95.200 ;
        RECT 155.800 94.800 157.000 95.100 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 158.200 94.800 158.600 95.200 ;
        RECT 150.200 93.200 150.500 94.800 ;
        RECT 151.000 93.800 151.400 94.200 ;
        RECT 148.600 92.800 149.000 93.200 ;
        RECT 150.200 92.800 150.600 93.200 ;
        RECT 147.800 91.800 148.200 92.200 ;
        RECT 146.200 87.800 146.600 88.200 ;
        RECT 146.200 86.800 146.600 87.200 ;
        RECT 147.000 86.800 147.400 87.200 ;
        RECT 135.800 85.800 136.200 86.200 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 139.000 86.100 139.400 86.200 ;
        RECT 139.800 86.100 140.200 86.200 ;
        RECT 139.000 85.800 140.200 86.100 ;
        RECT 141.400 85.800 141.800 86.200 ;
        RECT 142.200 85.800 142.600 86.200 ;
        RECT 143.800 85.800 144.200 86.200 ;
        RECT 144.600 85.800 145.000 86.200 ;
        RECT 145.400 85.800 145.800 86.200 ;
        RECT 131.800 72.100 132.200 77.900 ;
        RECT 133.400 75.100 133.800 75.200 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 133.400 74.800 134.600 75.100 ;
        RECT 132.600 73.100 133.000 73.200 ;
        RECT 133.400 73.100 133.800 73.200 ;
        RECT 132.600 72.800 133.800 73.100 ;
        RECT 136.600 72.100 137.000 77.900 ;
        RECT 131.800 68.800 132.200 69.200 ;
        RECT 131.800 67.200 132.100 68.800 ;
        RECT 131.800 66.800 132.200 67.200 ;
        RECT 136.600 66.800 137.000 67.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 136.600 66.200 136.900 66.800 ;
        RECT 137.400 66.200 137.700 66.800 ;
        RECT 138.200 66.200 138.500 85.800 ;
        RECT 139.000 83.800 139.400 84.200 ;
        RECT 139.000 79.200 139.300 83.800 ;
        RECT 141.400 82.200 141.700 85.800 ;
        RECT 142.200 84.200 142.500 85.800 ;
        RECT 142.200 83.800 142.600 84.200 ;
        RECT 141.400 81.800 141.800 82.200 ;
        RECT 143.000 81.800 143.400 82.200 ;
        RECT 141.400 81.200 141.700 81.800 ;
        RECT 141.400 80.800 141.800 81.200 ;
        RECT 139.000 78.800 139.400 79.200 ;
        RECT 139.000 75.800 139.400 76.200 ;
        RECT 141.400 75.800 141.800 76.200 ;
        RECT 142.200 75.800 142.600 76.200 ;
        RECT 139.000 67.200 139.300 75.800 ;
        RECT 141.400 75.200 141.700 75.800 ;
        RECT 142.200 75.200 142.500 75.800 ;
        RECT 143.000 75.200 143.300 81.800 ;
        RECT 139.800 74.800 140.200 75.200 ;
        RECT 141.400 74.800 141.800 75.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 139.800 69.200 140.100 74.800 ;
        RECT 142.200 72.800 142.600 73.200 ;
        RECT 140.600 71.800 141.000 72.200 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 140.600 68.200 140.900 71.800 ;
        RECT 142.200 70.200 142.500 72.800 ;
        RECT 142.200 69.800 142.600 70.200 ;
        RECT 142.200 69.200 142.500 69.800 ;
        RECT 142.200 68.800 142.600 69.200 ;
        RECT 140.600 67.800 141.000 68.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 133.400 66.100 133.800 66.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 133.400 65.800 134.600 66.100 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 138.200 65.800 138.600 66.200 ;
        RECT 131.000 60.800 131.400 61.200 ;
        RECT 136.600 60.800 137.000 61.200 ;
        RECT 136.600 59.200 136.900 60.800 ;
        RECT 139.000 60.200 139.300 66.800 ;
        RECT 141.400 64.800 141.800 65.200 ;
        RECT 139.000 59.800 139.400 60.200 ;
        RECT 141.400 59.200 141.700 64.800 ;
        RECT 136.600 58.800 137.000 59.200 ;
        RECT 141.400 58.800 141.800 59.200 ;
        RECT 143.000 58.800 143.400 59.200 ;
        RECT 127.800 58.100 128.200 58.200 ;
        RECT 128.600 58.100 129.000 58.200 ;
        RECT 117.400 54.800 117.800 55.200 ;
        RECT 118.200 54.800 118.600 55.200 ;
        RECT 117.400 54.200 117.700 54.800 ;
        RECT 117.400 53.800 117.800 54.200 ;
        RECT 116.600 51.800 117.000 52.200 ;
        RECT 116.600 51.200 116.900 51.800 ;
        RECT 116.600 50.800 117.000 51.200 ;
        RECT 117.400 46.800 117.800 47.200 ;
        RECT 117.400 46.200 117.700 46.800 ;
        RECT 117.400 45.800 117.800 46.200 ;
        RECT 115.800 39.800 116.200 40.200 ;
        RECT 118.200 37.200 118.500 54.800 ;
        RECT 119.000 53.100 119.400 55.900 ;
        RECT 119.800 53.800 120.200 54.200 ;
        RECT 119.800 52.100 120.100 53.800 ;
        RECT 120.600 52.100 121.000 57.900 ;
        RECT 123.000 55.100 123.400 55.200 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 123.000 54.800 124.200 55.100 ;
        RECT 125.400 52.100 125.800 57.900 ;
        RECT 127.800 57.800 129.000 58.100 ;
        RECT 139.800 57.800 140.200 58.200 ;
        RECT 130.200 56.800 130.600 57.200 ;
        RECT 134.200 56.800 134.600 57.200 ;
        RECT 139.000 56.800 139.400 57.200 ;
        RECT 130.200 56.200 130.500 56.800 ;
        RECT 130.200 55.800 130.600 56.200 ;
        RECT 132.600 55.800 133.000 56.200 ;
        RECT 132.600 55.200 132.900 55.800 ;
        RECT 131.000 55.100 131.400 55.200 ;
        RECT 131.800 55.100 132.200 55.200 ;
        RECT 131.000 54.800 132.200 55.100 ;
        RECT 132.600 54.800 133.000 55.200 ;
        RECT 133.400 53.800 133.800 54.200 ;
        RECT 119.000 51.800 120.100 52.100 ;
        RECT 119.000 39.200 119.300 51.800 ;
        RECT 120.600 50.800 121.000 51.200 ;
        RECT 119.800 43.100 120.200 48.900 ;
        RECT 119.000 38.800 119.400 39.200 ;
        RECT 119.000 38.200 119.300 38.800 ;
        RECT 119.000 37.800 119.400 38.200 ;
        RECT 118.200 36.800 118.600 37.200 ;
        RECT 117.400 35.800 117.800 36.200 ;
        RECT 117.400 34.200 117.700 35.800 ;
        RECT 117.400 33.800 117.800 34.200 ;
        RECT 120.600 29.200 120.900 50.800 ;
        RECT 125.400 49.800 125.800 50.200 ;
        RECT 125.400 47.200 125.700 49.800 ;
        RECT 128.600 47.800 129.000 48.200 ;
        RECT 128.600 47.200 128.900 47.800 ;
        RECT 123.000 46.800 123.400 47.200 ;
        RECT 125.400 46.800 125.800 47.200 ;
        RECT 126.200 46.800 126.600 47.200 ;
        RECT 128.600 46.800 129.000 47.200 ;
        RECT 123.000 46.200 123.300 46.800 ;
        RECT 123.000 45.800 123.400 46.200 ;
        RECT 124.600 45.800 125.000 46.200 ;
        RECT 123.000 45.100 123.400 45.200 ;
        RECT 123.800 45.100 124.200 45.200 ;
        RECT 123.000 44.800 124.200 45.100 ;
        RECT 124.600 44.200 124.900 45.800 ;
        RECT 126.200 45.200 126.500 46.800 ;
        RECT 127.800 46.100 128.200 46.200 ;
        RECT 128.600 46.100 129.000 46.200 ;
        RECT 127.800 45.800 129.000 46.100 ;
        RECT 126.200 44.800 126.600 45.200 ;
        RECT 127.800 44.800 128.200 45.200 ;
        RECT 129.400 45.100 129.800 47.900 ;
        RECT 124.600 43.800 125.000 44.200 ;
        RECT 126.200 43.800 126.600 44.200 ;
        RECT 126.200 42.200 126.500 43.800 ;
        RECT 122.200 42.100 122.600 42.200 ;
        RECT 123.000 42.100 123.400 42.200 ;
        RECT 122.200 41.800 123.400 42.100 ;
        RECT 126.200 41.800 126.600 42.200 ;
        RECT 123.000 38.800 123.400 39.200 ;
        RECT 104.600 23.800 105.000 24.200 ;
        RECT 109.400 23.800 109.800 24.200 ;
        RECT 104.600 19.200 104.900 23.800 ;
        RECT 111.000 23.100 111.400 28.900 ;
        RECT 114.200 28.800 114.600 29.200 ;
        RECT 113.400 26.100 113.800 26.200 ;
        RECT 114.200 26.100 114.600 26.200 ;
        RECT 113.400 25.800 114.600 26.100 ;
        RECT 115.800 23.100 116.200 28.900 ;
        RECT 120.600 28.800 121.000 29.200 ;
        RECT 116.600 27.800 117.000 28.200 ;
        RECT 116.600 27.200 116.900 27.800 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 116.600 25.800 117.000 26.200 ;
        RECT 108.600 21.800 109.000 22.200 ;
        RECT 108.600 21.200 108.900 21.800 ;
        RECT 106.200 20.800 106.600 21.200 ;
        RECT 108.600 20.800 109.000 21.200 ;
        RECT 106.200 19.200 106.500 20.800 ;
        RECT 108.600 19.800 109.000 20.200 ;
        RECT 114.200 19.800 114.600 20.200 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 106.200 18.800 106.600 19.200 ;
        RECT 103.000 13.100 103.400 15.900 ;
        RECT 106.200 15.200 106.500 18.800 ;
        RECT 108.600 15.200 108.900 19.800 ;
        RECT 106.200 14.800 106.600 15.200 ;
        RECT 108.600 14.800 109.000 15.200 ;
        RECT 111.000 14.800 111.400 15.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 113.400 14.800 113.800 15.200 ;
        RECT 111.000 14.200 111.300 14.800 ;
        RECT 111.800 14.200 112.100 14.800 ;
        RECT 108.600 14.100 109.000 14.200 ;
        RECT 109.400 14.100 109.800 14.200 ;
        RECT 108.600 13.800 109.800 14.100 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 111.800 13.800 112.200 14.200 ;
        RECT 113.400 13.200 113.700 14.800 ;
        RECT 113.400 12.800 113.800 13.200 ;
        RECT 113.400 12.200 113.700 12.800 ;
        RECT 104.600 11.800 105.000 12.200 ;
        RECT 107.800 11.800 108.200 12.200 ;
        RECT 113.400 11.800 113.800 12.200 ;
        RECT 104.600 9.200 104.900 11.800 ;
        RECT 101.400 5.800 101.800 6.200 ;
        RECT 102.200 5.800 102.600 6.200 ;
        RECT 103.000 3.100 103.400 8.900 ;
        RECT 104.600 8.800 105.000 9.200 ;
        RECT 104.600 6.200 104.900 8.800 ;
        RECT 107.800 8.200 108.100 11.800 ;
        RECT 107.800 7.800 108.200 8.200 ;
        RECT 114.200 7.200 114.500 19.800 ;
        RECT 116.600 19.200 116.900 25.800 ;
        RECT 117.400 25.100 117.800 27.900 ;
        RECT 118.200 26.800 118.600 27.200 ;
        RECT 118.200 26.200 118.500 26.800 ;
        RECT 123.000 26.200 123.300 38.800 ;
        RECT 126.200 35.200 126.500 41.800 ;
        RECT 127.800 39.200 128.100 44.800 ;
        RECT 131.000 43.100 131.400 48.900 ;
        RECT 131.800 48.800 132.200 49.200 ;
        RECT 131.800 48.200 132.100 48.800 ;
        RECT 131.800 47.800 132.200 48.200 ;
        RECT 132.600 45.800 133.000 46.200 ;
        RECT 131.800 43.800 132.200 44.200 ;
        RECT 131.800 39.200 132.100 43.800 ;
        RECT 132.600 43.200 132.900 45.800 ;
        RECT 133.400 44.200 133.700 53.800 ;
        RECT 133.400 43.800 133.800 44.200 ;
        RECT 132.600 42.800 133.000 43.200 ;
        RECT 127.800 38.800 128.200 39.200 ;
        RECT 131.800 38.800 132.200 39.200 ;
        RECT 134.200 36.100 134.500 56.800 ;
        RECT 138.200 55.800 138.600 56.200 ;
        RECT 138.200 55.200 138.500 55.800 ;
        RECT 139.000 55.200 139.300 56.800 ;
        RECT 139.800 55.200 140.100 57.800 ;
        RECT 143.000 55.200 143.300 58.800 ;
        RECT 143.800 57.200 144.100 85.800 ;
        RECT 144.600 83.800 145.000 84.200 ;
        RECT 144.600 79.200 144.900 83.800 ;
        RECT 144.600 78.800 145.000 79.200 ;
        RECT 146.200 78.200 146.500 86.800 ;
        RECT 147.000 86.200 147.300 86.800 ;
        RECT 147.000 85.800 147.400 86.200 ;
        RECT 147.800 79.200 148.100 91.800 ;
        RECT 148.600 89.200 148.900 92.800 ;
        RECT 151.000 89.200 151.300 93.800 ;
        RECT 151.800 93.200 152.100 94.800 ;
        RECT 152.600 94.200 152.900 94.800 ;
        RECT 155.800 94.200 156.100 94.800 ;
        RECT 157.400 94.200 157.700 94.800 ;
        RECT 152.600 93.800 153.000 94.200 ;
        RECT 155.800 93.800 156.200 94.200 ;
        RECT 157.400 93.800 157.800 94.200 ;
        RECT 151.800 92.800 152.200 93.200 ;
        RECT 148.600 88.800 149.000 89.200 ;
        RECT 151.000 88.800 151.400 89.200 ;
        RECT 149.400 87.800 149.800 88.200 ;
        RECT 149.400 87.200 149.700 87.800 ;
        RECT 149.400 86.800 149.800 87.200 ;
        RECT 150.200 81.800 150.600 82.200 ;
        RECT 147.800 78.800 148.200 79.200 ;
        RECT 146.200 77.800 146.600 78.200 ;
        RECT 145.400 74.800 145.800 75.200 ;
        RECT 145.400 59.200 145.700 74.800 ;
        RECT 147.000 73.100 147.400 75.900 ;
        RECT 147.800 74.200 148.100 78.800 ;
        RECT 150.200 78.200 150.500 81.800 ;
        RECT 147.800 73.800 148.200 74.200 ;
        RECT 148.600 72.100 149.000 77.900 ;
        RECT 150.200 77.800 150.600 78.200 ;
        RECT 151.800 75.200 152.100 92.800 ;
        RECT 159.800 90.200 160.100 95.800 ;
        RECT 161.400 93.100 161.800 95.900 ;
        RECT 162.200 94.200 162.500 110.800 ;
        RECT 164.600 108.200 164.900 125.800 ;
        RECT 165.400 112.100 165.800 117.900 ;
        RECT 166.200 109.200 166.500 126.800 ;
        RECT 167.000 126.100 167.400 126.200 ;
        RECT 167.800 126.100 168.200 126.200 ;
        RECT 167.000 125.800 168.200 126.100 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 168.600 125.200 168.900 125.800 ;
        RECT 168.600 124.800 169.000 125.200 ;
        RECT 167.800 114.800 168.200 115.200 ;
        RECT 167.800 114.200 168.100 114.800 ;
        RECT 167.800 113.800 168.200 114.200 ;
        RECT 169.400 111.100 169.700 127.800 ;
        RECT 170.200 125.200 170.500 128.800 ;
        RECT 171.000 127.800 171.400 128.200 ;
        RECT 171.000 127.200 171.300 127.800 ;
        RECT 171.000 126.800 171.400 127.200 ;
        RECT 170.200 125.100 170.600 125.200 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 170.200 124.800 171.400 125.100 ;
        RECT 171.000 122.800 171.400 123.200 ;
        RECT 170.200 112.100 170.600 117.900 ;
        RECT 171.000 114.200 171.300 122.800 ;
        RECT 171.000 113.800 171.400 114.200 ;
        RECT 171.800 113.100 172.200 115.900 ;
        RECT 169.400 110.800 170.500 111.100 ;
        RECT 166.200 108.800 166.600 109.200 ;
        RECT 163.000 107.800 163.400 108.200 ;
        RECT 164.600 107.800 165.000 108.200 ;
        RECT 167.800 107.800 168.200 108.200 ;
        RECT 163.000 107.200 163.300 107.800 ;
        RECT 167.800 107.200 168.100 107.800 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 164.600 106.800 165.000 107.200 ;
        RECT 167.800 106.800 168.200 107.200 ;
        RECT 169.400 106.800 169.800 107.200 ;
        RECT 163.800 106.200 164.100 106.800 ;
        RECT 164.600 106.200 164.900 106.800 ;
        RECT 163.000 105.800 163.400 106.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 164.600 105.800 165.000 106.200 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 167.000 106.100 167.400 106.200 ;
        RECT 166.200 105.800 167.400 106.100 ;
        RECT 168.600 105.800 169.000 106.200 ;
        RECT 163.000 105.200 163.300 105.800 ;
        RECT 168.600 105.200 168.900 105.800 ;
        RECT 169.400 105.200 169.700 106.800 ;
        RECT 170.200 106.200 170.500 110.800 ;
        RECT 170.200 105.800 170.600 106.200 ;
        RECT 163.000 104.800 163.400 105.200 ;
        RECT 166.200 105.100 166.600 105.200 ;
        RECT 167.000 105.100 167.400 105.200 ;
        RECT 166.200 104.800 167.400 105.100 ;
        RECT 168.600 104.800 169.000 105.200 ;
        RECT 169.400 104.800 169.800 105.200 ;
        RECT 170.200 101.200 170.500 105.800 ;
        RECT 171.000 104.100 171.400 104.200 ;
        RECT 171.800 104.100 172.200 104.200 ;
        RECT 171.000 103.800 172.200 104.100 ;
        RECT 170.200 100.800 170.600 101.200 ;
        RECT 162.200 93.800 162.600 94.200 ;
        RECT 160.600 91.800 161.000 92.200 ;
        RECT 163.000 92.100 163.400 97.900 ;
        RECT 164.600 95.100 165.000 95.200 ;
        RECT 165.400 95.100 165.800 95.200 ;
        RECT 164.600 94.800 165.800 95.100 ;
        RECT 164.600 93.800 165.000 94.200 ;
        RECT 163.800 92.800 164.200 93.200 ;
        RECT 163.800 92.200 164.100 92.800 ;
        RECT 163.800 91.800 164.200 92.200 ;
        RECT 159.800 89.800 160.200 90.200 ;
        RECT 153.400 83.100 153.800 88.900 ;
        RECT 157.400 86.800 157.800 87.200 ;
        RECT 157.400 86.300 157.700 86.800 ;
        RECT 154.200 85.800 154.600 86.200 ;
        RECT 157.400 85.900 157.800 86.300 ;
        RECT 151.000 74.800 151.400 75.200 ;
        RECT 151.800 74.800 152.200 75.200 ;
        RECT 151.000 69.200 151.300 74.800 ;
        RECT 153.400 72.100 153.800 77.900 ;
        RECT 151.000 68.800 151.400 69.200 ;
        RECT 151.000 67.800 151.400 68.200 ;
        RECT 148.600 66.800 149.000 67.200 ;
        RECT 149.400 66.800 149.800 67.200 ;
        RECT 148.600 66.200 148.900 66.800 ;
        RECT 149.400 66.200 149.700 66.800 ;
        RECT 146.200 65.800 146.600 66.200 ;
        RECT 148.600 65.800 149.000 66.200 ;
        RECT 149.400 65.800 149.800 66.200 ;
        RECT 145.400 58.800 145.800 59.200 ;
        RECT 143.800 56.800 144.200 57.200 ;
        RECT 135.000 54.800 135.400 55.200 ;
        RECT 137.400 54.800 137.800 55.200 ;
        RECT 138.200 54.800 138.600 55.200 ;
        RECT 139.000 54.800 139.400 55.200 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 142.200 54.800 142.600 55.200 ;
        RECT 143.000 54.800 143.400 55.200 ;
        RECT 144.600 54.800 145.000 55.200 ;
        RECT 135.000 45.200 135.300 54.800 ;
        RECT 135.000 44.800 135.400 45.200 ;
        RECT 135.800 43.100 136.200 48.900 ;
        RECT 137.400 42.200 137.700 54.800 ;
        RECT 142.200 53.200 142.500 54.800 ;
        RECT 142.200 52.800 142.600 53.200 ;
        RECT 144.600 51.200 144.900 54.800 ;
        RECT 143.000 50.800 143.400 51.200 ;
        RECT 144.600 50.800 145.000 51.200 ;
        RECT 139.800 48.800 140.200 49.200 ;
        RECT 139.000 47.800 139.400 48.200 ;
        RECT 139.000 47.200 139.300 47.800 ;
        RECT 139.000 46.800 139.400 47.200 ;
        RECT 139.800 46.200 140.100 48.800 ;
        RECT 139.800 45.800 140.200 46.200 ;
        RECT 143.000 45.200 143.300 50.800 ;
        RECT 146.200 49.200 146.500 65.800 ;
        RECT 151.000 65.200 151.300 67.800 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 151.800 66.200 152.100 66.800 ;
        RECT 151.800 65.800 152.200 66.200 ;
        RECT 152.600 65.800 153.000 66.200 ;
        RECT 152.600 65.200 152.900 65.800 ;
        RECT 151.000 64.800 151.400 65.200 ;
        RECT 152.600 64.800 153.000 65.200 ;
        RECT 147.000 54.800 147.400 55.200 ;
        RECT 147.000 52.200 147.300 54.800 ;
        RECT 148.600 53.100 149.000 55.900 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 147.000 51.800 147.400 52.200 ;
        RECT 146.200 48.800 146.600 49.200 ;
        RECT 143.800 47.100 144.200 47.200 ;
        RECT 144.600 47.100 145.000 47.200 ;
        RECT 143.800 46.800 145.000 47.100 ;
        RECT 143.800 45.800 144.200 46.200 ;
        RECT 143.800 45.200 144.100 45.800 ;
        RECT 138.200 44.800 138.600 45.200 ;
        RECT 142.200 45.100 142.600 45.200 ;
        RECT 143.000 45.100 143.400 45.200 ;
        RECT 142.200 44.800 143.400 45.100 ;
        RECT 143.800 44.800 144.200 45.200 ;
        RECT 138.200 44.200 138.500 44.800 ;
        RECT 138.200 43.800 138.600 44.200 ;
        RECT 143.000 43.800 143.400 44.200 ;
        RECT 143.000 43.200 143.300 43.800 ;
        RECT 139.800 42.800 140.200 43.200 ;
        RECT 143.000 42.800 143.400 43.200 ;
        RECT 139.800 42.200 140.100 42.800 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 137.400 41.800 137.800 42.200 ;
        RECT 139.800 41.800 140.200 42.200 ;
        RECT 135.800 39.200 136.100 41.800 ;
        RECT 135.800 38.800 136.200 39.200 ;
        RECT 133.400 35.800 134.500 36.100 ;
        RECT 133.400 35.200 133.700 35.800 ;
        RECT 143.000 35.200 143.300 42.800 ;
        RECT 143.800 38.200 144.100 44.800 ;
        RECT 144.600 40.200 144.900 46.800 ;
        RECT 146.200 46.200 146.500 48.800 ;
        RECT 145.400 45.800 145.800 46.200 ;
        RECT 146.200 45.800 146.600 46.200 ;
        RECT 145.400 42.200 145.700 45.800 ;
        RECT 145.400 41.800 145.800 42.200 ;
        RECT 147.000 41.800 147.400 42.200 ;
        RECT 144.600 39.800 145.000 40.200 ;
        RECT 145.400 39.200 145.700 41.800 ;
        RECT 145.400 38.800 145.800 39.200 ;
        RECT 143.800 37.800 144.200 38.200 ;
        RECT 125.400 34.800 125.800 35.200 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 133.400 35.100 133.800 35.200 ;
        RECT 132.600 34.800 133.800 35.100 ;
        RECT 134.200 34.800 134.600 35.200 ;
        RECT 138.200 34.800 138.600 35.200 ;
        RECT 139.800 35.100 140.200 35.200 ;
        RECT 140.600 35.100 141.000 35.200 ;
        RECT 139.800 34.800 141.000 35.100 ;
        RECT 142.200 34.800 142.600 35.200 ;
        RECT 143.000 34.800 143.400 35.200 ;
        RECT 123.800 34.100 124.200 34.200 ;
        RECT 124.600 34.100 125.000 34.200 ;
        RECT 123.800 33.800 125.000 34.100 ;
        RECT 118.200 25.800 118.600 26.200 ;
        RECT 119.000 25.800 119.400 26.200 ;
        RECT 121.400 25.800 121.800 26.200 ;
        RECT 123.000 25.800 123.400 26.200 ;
        RECT 123.800 25.800 124.200 26.200 ;
        RECT 119.000 25.200 119.300 25.800 ;
        RECT 119.000 24.800 119.400 25.200 ;
        RECT 119.800 20.800 120.200 21.200 ;
        RECT 116.600 18.800 117.000 19.200 ;
        RECT 118.200 17.800 118.600 18.200 ;
        RECT 118.200 15.200 118.500 17.800 ;
        RECT 119.800 15.200 120.100 20.800 ;
        RECT 121.400 19.200 121.700 25.800 ;
        RECT 123.800 24.200 124.100 25.800 ;
        RECT 123.800 23.800 124.200 24.200 ;
        RECT 121.400 18.800 121.800 19.200 ;
        RECT 125.400 16.200 125.700 34.800 ;
        RECT 128.600 28.200 128.900 34.800 ;
        RECT 130.200 31.200 130.500 34.800 ;
        RECT 130.200 30.800 130.600 31.200 ;
        RECT 128.600 27.800 129.000 28.200 ;
        RECT 127.000 26.800 127.400 27.200 ;
        RECT 127.000 26.200 127.300 26.800 ;
        RECT 127.000 25.800 127.400 26.200 ;
        RECT 130.200 19.200 130.500 30.800 ;
        RECT 131.800 23.100 132.200 28.900 ;
        RECT 130.200 18.800 130.600 19.200 ;
        RECT 132.600 18.200 132.900 34.800 ;
        RECT 133.400 33.800 133.800 34.200 ;
        RECT 123.000 15.800 123.400 16.200 ;
        RECT 125.400 15.800 125.800 16.200 ;
        RECT 123.000 15.200 123.300 15.800 ;
        RECT 117.400 14.800 117.800 15.200 ;
        RECT 118.200 14.800 118.600 15.200 ;
        RECT 119.800 14.800 120.200 15.200 ;
        RECT 122.200 14.800 122.600 15.200 ;
        RECT 123.000 14.800 123.400 15.200 ;
        RECT 117.400 9.200 117.700 14.800 ;
        RECT 122.200 10.200 122.500 14.800 ;
        RECT 123.000 12.100 123.400 12.200 ;
        RECT 123.800 12.100 124.200 12.200 ;
        RECT 126.200 12.100 126.600 17.900 ;
        RECT 128.600 15.100 129.000 15.200 ;
        RECT 129.400 15.100 129.800 15.200 ;
        RECT 128.600 14.800 129.800 15.100 ;
        RECT 131.000 12.100 131.400 17.900 ;
        RECT 132.600 17.800 133.000 18.200 ;
        RECT 131.800 13.800 132.200 14.200 ;
        RECT 123.000 11.800 124.200 12.100 ;
        RECT 122.200 9.800 122.600 10.200 ;
        RECT 129.400 9.800 129.800 10.200 ;
        RECT 117.400 8.800 117.800 9.200 ;
        RECT 119.800 8.800 120.200 9.200 ;
        RECT 119.800 8.200 120.100 8.800 ;
        RECT 119.800 7.800 120.200 8.200 ;
        RECT 109.400 7.100 109.800 7.200 ;
        RECT 110.200 7.100 110.600 7.200 ;
        RECT 109.400 6.800 110.600 7.100 ;
        RECT 113.400 6.800 113.800 7.200 ;
        RECT 114.200 6.800 114.600 7.200 ;
        RECT 117.400 6.800 117.800 7.200 ;
        RECT 113.400 6.200 113.700 6.800 ;
        RECT 117.400 6.200 117.700 6.800 ;
        RECT 104.600 5.800 105.000 6.200 ;
        RECT 111.800 6.100 112.200 6.200 ;
        RECT 112.600 6.100 113.000 6.200 ;
        RECT 111.800 5.800 113.000 6.100 ;
        RECT 113.400 5.800 113.800 6.200 ;
        RECT 115.000 5.800 115.400 6.200 ;
        RECT 117.400 5.800 117.800 6.200 ;
        RECT 115.000 4.200 115.300 5.800 ;
        RECT 117.400 4.800 117.800 5.200 ;
        RECT 117.400 4.200 117.700 4.800 ;
        RECT 115.000 3.800 115.400 4.200 ;
        RECT 117.400 3.800 117.800 4.200 ;
        RECT 122.200 3.100 122.600 8.900 ;
        RECT 124.600 6.100 125.000 6.200 ;
        RECT 125.400 6.100 125.800 6.200 ;
        RECT 124.600 5.800 125.800 6.100 ;
        RECT 127.000 3.100 127.400 8.900 ;
        RECT 127.800 7.800 128.200 8.200 ;
        RECT 127.800 7.200 128.100 7.800 ;
        RECT 127.800 6.800 128.200 7.200 ;
        RECT 128.600 5.100 129.000 7.900 ;
        RECT 129.400 7.200 129.700 9.800 ;
        RECT 131.800 8.200 132.100 13.800 ;
        RECT 132.600 13.100 133.000 15.900 ;
        RECT 133.400 14.200 133.700 33.800 ;
        RECT 134.200 33.200 134.500 34.800 ;
        RECT 138.200 33.200 138.500 34.800 ;
        RECT 142.200 34.200 142.500 34.800 ;
        RECT 142.200 33.800 142.600 34.200 ;
        RECT 134.200 32.800 134.600 33.200 ;
        RECT 138.200 32.800 138.600 33.200 ;
        RECT 143.800 33.100 144.200 35.900 ;
        RECT 144.600 34.800 145.000 35.200 ;
        RECT 144.600 34.200 144.900 34.800 ;
        RECT 144.600 33.800 145.000 34.200 ;
        RECT 138.200 29.100 138.500 32.800 ;
        RECT 141.400 31.800 141.800 32.200 ;
        RECT 145.400 32.100 145.800 37.900 ;
        RECT 147.000 35.200 147.300 41.800 ;
        RECT 149.400 35.200 149.700 53.800 ;
        RECT 150.200 52.100 150.600 57.900 ;
        RECT 151.800 55.100 152.200 55.200 ;
        RECT 152.600 55.100 153.000 55.200 ;
        RECT 151.800 54.800 153.000 55.100 ;
        RECT 151.800 52.800 152.200 53.200 ;
        RECT 151.000 51.800 151.400 52.200 ;
        RECT 151.000 48.200 151.300 51.800 ;
        RECT 151.800 49.200 152.100 52.800 ;
        RECT 151.800 48.800 152.200 49.200 ;
        RECT 151.000 47.800 151.400 48.200 ;
        RECT 151.000 39.200 151.300 47.800 ;
        RECT 151.800 47.200 152.100 48.800 ;
        RECT 151.800 46.800 152.200 47.200 ;
        RECT 153.400 45.800 153.800 46.200 ;
        RECT 153.400 45.200 153.700 45.800 ;
        RECT 153.400 44.800 153.800 45.200 ;
        RECT 153.400 39.800 153.800 40.200 ;
        RECT 151.000 38.800 151.400 39.200 ;
        RECT 151.800 39.100 152.200 39.200 ;
        RECT 152.600 39.100 153.000 39.200 ;
        RECT 151.800 38.800 153.000 39.100 ;
        RECT 147.000 34.800 147.400 35.200 ;
        RECT 149.400 34.800 149.800 35.200 ;
        RECT 150.200 32.100 150.600 37.900 ;
        RECT 153.400 33.200 153.700 39.800 ;
        RECT 154.200 39.200 154.500 85.800 ;
        RECT 158.200 83.100 158.600 88.900 ;
        RECT 159.000 88.800 159.400 89.200 ;
        RECT 159.000 87.200 159.300 88.800 ;
        RECT 159.000 86.800 159.400 87.200 ;
        RECT 159.800 85.100 160.200 87.900 ;
        RECT 160.600 85.200 160.900 91.800 ;
        RECT 163.800 89.800 164.200 90.200 ;
        RECT 161.400 87.800 161.800 88.200 ;
        RECT 161.400 87.200 161.700 87.800 ;
        RECT 161.400 86.800 161.800 87.200 ;
        RECT 163.800 86.200 164.100 89.800 ;
        RECT 164.600 87.200 164.900 93.800 ;
        RECT 167.800 92.100 168.200 97.900 ;
        RECT 172.600 96.200 172.900 143.800 ;
        RECT 173.400 136.800 173.800 137.200 ;
        RECT 173.400 126.200 173.700 136.800 ;
        RECT 174.200 134.200 174.500 146.800 ;
        RECT 175.000 143.100 175.400 148.900 ;
        RECT 176.600 145.100 177.000 147.900 ;
        RECT 177.400 145.800 177.800 146.200 ;
        RECT 178.200 146.100 178.600 146.200 ;
        RECT 179.000 146.100 179.400 146.200 ;
        RECT 178.200 145.800 179.400 146.100 ;
        RECT 177.400 143.200 177.700 145.800 ;
        RECT 182.200 145.200 182.500 154.800 ;
        RECT 183.000 153.100 183.400 155.900 ;
        RECT 184.600 152.100 185.000 157.900 ;
        RECT 186.200 157.200 186.500 165.800 ;
        RECT 188.600 160.200 188.900 184.800 ;
        RECT 189.400 181.200 189.700 185.800 ;
        RECT 189.400 180.800 189.800 181.200 ;
        RECT 189.400 172.100 189.800 177.900 ;
        RECT 190.200 174.800 190.600 175.200 ;
        RECT 190.200 174.200 190.500 174.800 ;
        RECT 190.200 173.800 190.600 174.200 ;
        RECT 191.000 173.100 191.400 175.900 ;
        RECT 191.800 175.800 192.200 176.200 ;
        RECT 191.800 175.200 192.100 175.800 ;
        RECT 192.600 175.200 192.900 189.800 ;
        RECT 196.600 186.200 196.900 192.800 ;
        RECT 199.000 186.200 199.300 199.800 ;
        RECT 199.800 192.100 200.200 197.900 ;
        RECT 200.600 194.800 201.000 195.200 ;
        RECT 200.600 194.200 200.900 194.800 ;
        RECT 200.600 193.800 201.000 194.200 ;
        RECT 201.400 193.100 201.800 195.900 ;
        RECT 202.200 193.200 202.500 201.800 ;
        RECT 202.200 192.800 202.600 193.200 ;
        RECT 201.400 191.800 201.800 192.200 ;
        RECT 202.200 192.100 202.600 192.200 ;
        RECT 203.000 192.100 203.400 192.200 ;
        RECT 204.600 192.100 205.000 197.900 ;
        RECT 207.000 195.200 207.300 211.800 ;
        RECT 211.000 209.800 211.400 210.200 ;
        RECT 211.000 209.200 211.300 209.800 ;
        RECT 211.000 208.800 211.400 209.200 ;
        RECT 213.400 208.200 213.700 211.800 ;
        RECT 211.800 207.800 212.200 208.200 ;
        RECT 213.400 207.800 213.800 208.200 ;
        RECT 211.800 206.200 212.100 207.800 ;
        RECT 211.800 205.800 212.200 206.200 ;
        RECT 212.600 205.800 213.000 206.200 ;
        RECT 210.200 198.800 210.600 199.200 ;
        RECT 208.600 195.800 209.000 196.200 ;
        RECT 207.000 194.800 207.400 195.200 ;
        RECT 208.600 195.100 208.900 195.800 ;
        RECT 207.000 194.200 207.300 194.800 ;
        RECT 208.600 194.700 209.000 195.100 ;
        RECT 207.000 193.800 207.400 194.200 ;
        RECT 209.400 192.100 209.800 197.900 ;
        RECT 202.200 191.800 203.400 192.100 ;
        RECT 200.600 187.800 201.000 188.200 ;
        RECT 200.600 187.200 200.900 187.800 ;
        RECT 200.600 186.800 201.000 187.200 ;
        RECT 201.400 186.200 201.700 191.800 ;
        RECT 206.200 187.800 206.600 188.200 ;
        RECT 203.800 186.800 204.200 187.200 ;
        RECT 203.800 186.200 204.100 186.800 ;
        RECT 206.200 186.200 206.500 187.800 ;
        RECT 210.200 186.200 210.500 198.800 ;
        RECT 211.800 197.200 212.100 205.800 ;
        RECT 212.600 205.200 212.900 205.800 ;
        RECT 212.600 204.800 213.000 205.200 ;
        RECT 211.800 196.800 212.200 197.200 ;
        RECT 211.000 193.100 211.400 195.900 ;
        RECT 211.800 193.800 212.200 194.200 ;
        RECT 211.800 192.200 212.100 193.800 ;
        RECT 211.800 191.800 212.200 192.200 ;
        RECT 213.400 188.100 213.700 207.800 ;
        RECT 215.800 206.200 216.100 225.800 ;
        RECT 216.600 222.200 216.900 225.800 ;
        RECT 217.400 225.100 217.800 227.900 ;
        RECT 219.000 223.100 219.400 228.900 ;
        RECT 220.600 227.200 220.900 232.800 ;
        RECT 223.800 231.800 224.200 232.200 ;
        RECT 223.800 230.200 224.100 231.800 ;
        RECT 221.400 229.800 221.800 230.200 ;
        RECT 223.800 229.800 224.200 230.200 ;
        RECT 220.600 226.800 221.000 227.200 ;
        RECT 216.600 221.800 217.000 222.200 ;
        RECT 220.600 218.200 220.900 226.800 ;
        RECT 221.400 226.200 221.700 229.800 ;
        RECT 226.200 229.200 226.500 233.800 ;
        RECT 227.000 233.200 227.300 233.800 ;
        RECT 227.000 232.800 227.400 233.200 ;
        RECT 234.200 233.100 234.600 235.900 ;
        RECT 235.800 232.100 236.200 237.900 ;
        RECT 238.200 234.800 238.600 235.200 ;
        RECT 237.400 233.800 237.800 234.200 ;
        RECT 221.400 225.800 221.800 226.200 ;
        RECT 223.800 223.100 224.200 228.900 ;
        RECT 226.200 228.800 226.600 229.200 ;
        RECT 231.800 227.800 232.200 228.200 ;
        RECT 231.800 226.200 232.100 227.800 ;
        RECT 234.200 226.800 234.600 227.200 ;
        RECT 235.800 227.100 236.200 227.200 ;
        RECT 236.600 227.100 237.000 227.200 ;
        RECT 235.800 226.800 237.000 227.100 ;
        RECT 234.200 226.200 234.500 226.800 ;
        RECT 231.800 225.800 232.200 226.200 ;
        RECT 234.200 225.800 234.600 226.200 ;
        RECT 235.000 225.800 235.400 226.200 ;
        RECT 236.600 225.800 237.000 226.200 ;
        RECT 235.000 225.200 235.300 225.800 ;
        RECT 236.600 225.200 236.900 225.800 ;
        RECT 235.000 224.800 235.400 225.200 ;
        RECT 236.600 224.800 237.000 225.200 ;
        RECT 223.800 221.800 224.200 222.200 ;
        RECT 226.200 221.800 226.600 222.200 ;
        RECT 227.800 221.800 228.200 222.200 ;
        RECT 232.600 221.800 233.000 222.200 ;
        RECT 223.800 219.200 224.100 221.800 ;
        RECT 223.800 218.800 224.200 219.200 ;
        RECT 225.400 218.800 225.800 219.200 ;
        RECT 216.600 212.100 217.000 217.900 ;
        RECT 220.600 217.800 221.000 218.200 ;
        RECT 218.200 217.100 218.600 217.200 ;
        RECT 219.000 217.100 219.400 217.200 ;
        RECT 218.200 216.800 219.400 217.100 ;
        RECT 225.400 215.200 225.700 218.800 ;
        RECT 226.200 217.200 226.500 221.800 ;
        RECT 227.800 219.200 228.100 221.800 ;
        RECT 227.800 218.800 228.200 219.200 ;
        RECT 226.200 216.800 226.600 217.200 ;
        RECT 217.400 214.800 217.800 215.200 ;
        RECT 219.800 214.800 220.200 215.200 ;
        RECT 225.400 214.800 225.800 215.200 ;
        RECT 217.400 211.100 217.700 214.800 ;
        RECT 219.800 214.200 220.100 214.800 ;
        RECT 219.800 213.800 220.200 214.200 ;
        RECT 222.200 213.800 222.600 214.200 ;
        RECT 221.400 211.800 221.800 212.200 ;
        RECT 216.600 210.800 217.700 211.100 ;
        RECT 219.800 210.800 220.200 211.200 ;
        RECT 216.600 209.200 216.900 210.800 ;
        RECT 216.600 208.800 217.000 209.200 ;
        RECT 217.400 206.800 217.800 207.200 ;
        RECT 218.200 206.800 218.600 207.200 ;
        RECT 217.400 206.200 217.700 206.800 ;
        RECT 218.200 206.200 218.500 206.800 ;
        RECT 219.800 206.200 220.100 210.800 ;
        RECT 221.400 208.200 221.700 211.800 ;
        RECT 221.400 207.800 221.800 208.200 ;
        RECT 221.400 206.200 221.700 207.800 ;
        RECT 214.200 206.100 214.600 206.200 ;
        RECT 215.000 206.100 215.400 206.200 ;
        RECT 214.200 205.800 215.400 206.100 ;
        RECT 215.800 205.800 216.200 206.200 ;
        RECT 217.400 205.800 217.800 206.200 ;
        RECT 218.200 205.800 218.600 206.200 ;
        RECT 219.000 205.800 219.400 206.200 ;
        RECT 219.800 205.800 220.200 206.200 ;
        RECT 221.400 205.800 221.800 206.200 ;
        RECT 219.000 201.200 219.300 205.800 ;
        RECT 220.600 201.800 221.000 202.200 ;
        RECT 219.000 200.800 219.400 201.200 ;
        RECT 218.200 196.800 218.600 197.200 ;
        RECT 214.200 196.100 214.600 196.200 ;
        RECT 215.000 196.100 215.400 196.200 ;
        RECT 214.200 195.800 215.400 196.100 ;
        RECT 217.400 195.800 217.800 196.200 ;
        RECT 217.400 195.200 217.700 195.800 ;
        RECT 215.000 194.800 215.400 195.200 ;
        RECT 217.400 194.800 217.800 195.200 ;
        RECT 215.000 194.200 215.300 194.800 ;
        RECT 218.200 194.200 218.500 196.800 ;
        RECT 219.000 194.800 219.400 195.200 ;
        RECT 219.800 195.100 220.200 195.200 ;
        RECT 220.600 195.100 220.900 201.800 ;
        RECT 219.800 194.800 220.900 195.100 ;
        RECT 222.200 195.200 222.500 213.800 ;
        RECT 223.000 207.100 223.400 207.200 ;
        RECT 223.800 207.100 224.200 207.200 ;
        RECT 223.000 206.800 224.200 207.100 ;
        RECT 223.000 206.100 223.400 206.200 ;
        RECT 223.800 206.100 224.200 206.200 ;
        RECT 223.000 205.800 224.200 206.100 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 224.600 203.200 224.900 205.800 ;
        RECT 224.600 202.800 225.000 203.200 ;
        RECT 225.400 198.200 225.700 214.800 ;
        RECT 226.200 212.100 226.600 212.200 ;
        RECT 227.000 212.100 227.400 212.200 ;
        RECT 228.600 212.100 229.000 217.900 ;
        RECT 231.000 215.100 231.400 215.200 ;
        RECT 231.800 215.100 232.200 215.200 ;
        RECT 231.000 214.800 232.200 215.100 ;
        RECT 232.600 214.200 232.900 221.800 ;
        RECT 232.600 213.800 233.000 214.200 ;
        RECT 233.400 212.100 233.800 217.900 ;
        RECT 234.200 214.800 234.600 215.200 ;
        RECT 234.200 214.200 234.500 214.800 ;
        RECT 234.200 213.800 234.600 214.200 ;
        RECT 235.000 213.100 235.400 215.900 ;
        RECT 235.800 212.800 236.200 213.200 ;
        RECT 235.800 212.200 236.100 212.800 ;
        RECT 226.200 211.800 227.400 212.100 ;
        RECT 235.800 211.800 236.200 212.200 ;
        RECT 236.600 211.100 236.900 224.800 ;
        RECT 237.400 217.200 237.700 233.800 ;
        RECT 238.200 229.200 238.500 234.800 ;
        RECT 240.600 232.100 241.000 237.900 ;
        RECT 241.400 236.800 241.800 237.200 ;
        RECT 243.000 237.100 243.400 237.200 ;
        RECT 243.800 237.100 244.200 237.200 ;
        RECT 243.000 236.800 244.200 237.100 ;
        RECT 238.200 228.800 238.600 229.200 ;
        RECT 240.600 227.800 241.000 228.200 ;
        RECT 240.600 227.200 240.900 227.800 ;
        RECT 241.400 227.200 241.700 236.800 ;
        RECT 243.800 234.800 244.200 235.200 ;
        RECT 243.000 231.800 243.400 232.200 ;
        RECT 243.000 228.200 243.300 231.800 ;
        RECT 243.800 229.200 244.100 234.800 ;
        RECT 246.200 232.100 246.600 237.900 ;
        RECT 247.800 235.100 248.200 235.200 ;
        RECT 248.600 235.100 249.000 235.200 ;
        RECT 247.800 234.800 249.000 235.100 ;
        RECT 250.200 232.800 250.600 233.200 ;
        RECT 243.800 228.800 244.200 229.200 ;
        RECT 243.000 227.800 243.400 228.200 ;
        RECT 249.400 227.800 249.800 228.200 ;
        RECT 240.600 226.800 241.000 227.200 ;
        RECT 241.400 226.800 241.800 227.200 ;
        RECT 246.200 226.800 246.600 227.200 ;
        RECT 241.400 226.200 241.700 226.800 ;
        RECT 241.400 225.800 241.800 226.200 ;
        RECT 245.400 225.800 245.800 226.200 ;
        RECT 245.400 225.200 245.700 225.800 ;
        RECT 238.200 225.100 238.600 225.200 ;
        RECT 239.000 225.100 239.400 225.200 ;
        RECT 238.200 224.800 239.400 225.100 ;
        RECT 243.000 225.100 243.400 225.200 ;
        RECT 243.800 225.100 244.200 225.200 ;
        RECT 243.000 224.800 244.200 225.100 ;
        RECT 245.400 224.800 245.800 225.200 ;
        RECT 237.400 216.800 237.800 217.200 ;
        RECT 238.200 212.100 238.600 217.900 ;
        RECT 241.400 214.800 241.800 215.200 ;
        RECT 239.000 213.800 239.400 214.200 ;
        RECT 239.000 213.200 239.300 213.800 ;
        RECT 239.000 212.800 239.400 213.200 ;
        RECT 241.400 212.200 241.700 214.800 ;
        RECT 241.400 211.800 241.800 212.200 ;
        RECT 243.000 212.100 243.400 217.900 ;
        RECT 243.800 215.800 244.200 216.200 ;
        RECT 243.800 214.200 244.100 215.800 ;
        RECT 243.800 213.800 244.200 214.200 ;
        RECT 244.600 213.100 245.000 215.900 ;
        RECT 245.400 213.100 245.800 215.900 ;
        RECT 235.800 210.800 236.900 211.100 ;
        RECT 228.600 209.800 229.000 210.200 ;
        RECT 226.200 208.800 226.600 209.200 ;
        RECT 226.200 206.200 226.500 208.800 ;
        RECT 228.600 208.200 228.900 209.800 ;
        RECT 229.400 209.100 229.800 209.200 ;
        RECT 230.200 209.100 230.600 209.200 ;
        RECT 229.400 208.800 230.600 209.100 ;
        RECT 228.600 207.800 229.000 208.200 ;
        RECT 228.600 206.200 228.900 207.800 ;
        RECT 229.400 207.100 229.800 207.200 ;
        RECT 230.200 207.100 230.600 207.200 ;
        RECT 229.400 206.800 230.600 207.100 ;
        RECT 226.200 205.800 226.600 206.200 ;
        RECT 227.000 206.100 227.400 206.200 ;
        RECT 227.800 206.100 228.200 206.200 ;
        RECT 227.000 205.800 228.200 206.100 ;
        RECT 228.600 205.800 229.000 206.200 ;
        RECT 226.200 205.200 226.500 205.800 ;
        RECT 226.200 204.800 226.600 205.200 ;
        RECT 232.600 203.100 233.000 208.900 ;
        RECT 234.200 206.100 234.600 206.200 ;
        RECT 235.000 206.100 235.400 206.200 ;
        RECT 234.200 205.800 235.400 206.100 ;
        RECT 227.000 199.800 227.400 200.200 ;
        RECT 230.200 199.800 230.600 200.200 ;
        RECT 223.800 197.800 224.200 198.200 ;
        RECT 225.400 197.800 225.800 198.200 ;
        RECT 223.800 195.200 224.100 197.800 ;
        RECT 224.600 196.800 225.000 197.200 ;
        RECT 222.200 194.800 222.600 195.200 ;
        RECT 223.800 194.800 224.200 195.200 ;
        RECT 219.000 194.200 219.300 194.800 ;
        RECT 215.000 193.800 215.400 194.200 ;
        RECT 218.200 193.800 218.600 194.200 ;
        RECT 219.000 193.800 219.400 194.200 ;
        RECT 220.600 191.800 221.000 192.200 ;
        RECT 220.600 190.100 220.900 191.800 ;
        RECT 212.600 187.800 213.700 188.100 ;
        RECT 219.800 189.800 220.900 190.100 ;
        RECT 212.600 186.200 212.900 187.800 ;
        RECT 213.400 186.800 213.800 187.200 ;
        RECT 215.000 186.800 215.400 187.200 ;
        RECT 213.400 186.200 213.700 186.800 ;
        RECT 215.000 186.200 215.300 186.800 ;
        RECT 196.600 185.800 197.000 186.200 ;
        RECT 197.400 185.800 197.800 186.200 ;
        RECT 199.000 185.800 199.400 186.200 ;
        RECT 201.400 185.800 201.800 186.200 ;
        RECT 202.200 185.800 202.600 186.200 ;
        RECT 203.000 185.800 203.400 186.200 ;
        RECT 203.800 185.800 204.200 186.200 ;
        RECT 206.200 185.800 206.600 186.200 ;
        RECT 209.400 185.800 209.800 186.200 ;
        RECT 210.200 185.800 210.600 186.200 ;
        RECT 212.600 185.800 213.000 186.200 ;
        RECT 213.400 185.800 213.800 186.200 ;
        RECT 214.200 185.800 214.600 186.200 ;
        RECT 215.000 185.800 215.400 186.200 ;
        RECT 217.400 186.100 217.800 186.200 ;
        RECT 218.200 186.100 218.600 186.200 ;
        RECT 217.400 185.800 218.600 186.100 ;
        RECT 195.800 181.800 196.200 182.200 ;
        RECT 195.800 181.200 196.100 181.800 ;
        RECT 195.800 180.800 196.200 181.200 ;
        RECT 197.400 179.200 197.700 185.800 ;
        RECT 197.400 178.800 197.800 179.200 ;
        RECT 194.200 176.800 194.600 177.200 ;
        RECT 195.000 176.800 195.400 177.200 ;
        RECT 194.200 176.200 194.500 176.800 ;
        RECT 194.200 175.800 194.600 176.200 ;
        RECT 195.000 175.200 195.300 176.800 ;
        RECT 191.800 174.800 192.200 175.200 ;
        RECT 192.600 174.800 193.000 175.200 ;
        RECT 195.000 174.800 195.400 175.200 ;
        RECT 192.600 170.100 192.900 174.800 ;
        RECT 196.600 173.100 197.000 175.900 ;
        RECT 197.400 174.800 197.800 175.200 ;
        RECT 197.400 174.200 197.700 174.800 ;
        RECT 197.400 173.800 197.800 174.200 ;
        RECT 198.200 172.100 198.600 177.900 ;
        RECT 199.000 175.800 199.400 176.200 ;
        RECT 199.000 175.100 199.300 175.800 ;
        RECT 199.000 174.700 199.400 175.100 ;
        RECT 199.000 172.800 199.400 173.200 ;
        RECT 192.600 169.800 193.700 170.100 ;
        RECT 189.400 168.800 189.800 169.200 ;
        RECT 192.600 168.800 193.000 169.200 ;
        RECT 189.400 167.200 189.700 168.800 ;
        RECT 192.600 167.200 192.900 168.800 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 192.600 166.800 193.000 167.200 ;
        RECT 189.400 166.100 189.800 166.200 ;
        RECT 190.200 166.100 190.600 166.200 ;
        RECT 189.400 165.800 190.600 166.100 ;
        RECT 189.400 165.100 189.800 165.200 ;
        RECT 191.000 165.100 191.400 165.200 ;
        RECT 189.400 164.800 191.400 165.100 ;
        RECT 193.400 163.200 193.700 169.800 ;
        RECT 199.000 169.200 199.300 172.800 ;
        RECT 202.200 171.200 202.500 185.800 ;
        RECT 203.000 185.200 203.300 185.800 ;
        RECT 203.000 184.800 203.400 185.200 ;
        RECT 209.400 182.200 209.700 185.800 ;
        RECT 205.400 181.800 205.800 182.200 ;
        RECT 209.400 181.800 209.800 182.200 ;
        RECT 205.400 178.200 205.700 181.800 ;
        RECT 213.400 180.800 213.800 181.200 ;
        RECT 203.000 172.100 203.400 177.900 ;
        RECT 205.400 177.800 205.800 178.200 ;
        RECT 211.000 177.800 211.400 178.200 ;
        RECT 206.200 177.100 206.600 177.200 ;
        RECT 207.000 177.100 207.400 177.200 ;
        RECT 206.200 176.800 207.400 177.100 ;
        RECT 207.000 175.800 207.400 176.200 ;
        RECT 209.400 175.800 209.800 176.200 ;
        RECT 207.000 173.200 207.300 175.800 ;
        RECT 209.400 173.200 209.700 175.800 ;
        RECT 211.000 175.200 211.300 177.800 ;
        RECT 211.000 174.800 211.400 175.200 ;
        RECT 211.000 173.800 211.400 174.200 ;
        RECT 211.800 174.100 212.200 174.200 ;
        RECT 212.600 174.100 213.000 174.200 ;
        RECT 211.800 173.800 213.000 174.100 ;
        RECT 213.400 174.100 213.700 180.800 ;
        RECT 214.200 179.200 214.500 185.800 ;
        RECT 219.000 185.100 219.400 187.900 ;
        RECT 216.600 181.800 217.000 182.200 ;
        RECT 214.200 178.800 214.600 179.200 ;
        RECT 214.200 175.100 214.600 175.200 ;
        RECT 215.000 175.100 215.400 175.200 ;
        RECT 214.200 174.800 215.400 175.100 ;
        RECT 216.600 174.200 216.900 181.800 ;
        RECT 219.000 178.800 219.400 179.200 ;
        RECT 214.200 174.100 214.600 174.200 ;
        RECT 213.400 173.800 214.600 174.100 ;
        RECT 216.600 173.800 217.000 174.200 ;
        RECT 218.200 173.800 218.600 174.200 ;
        RECT 211.000 173.200 211.300 173.800 ;
        RECT 218.200 173.200 218.500 173.800 ;
        RECT 207.000 172.800 207.400 173.200 ;
        RECT 209.400 172.800 209.800 173.200 ;
        RECT 211.000 172.800 211.400 173.200 ;
        RECT 213.400 173.100 213.800 173.200 ;
        RECT 214.200 173.100 214.600 173.200 ;
        RECT 213.400 172.800 214.600 173.100 ;
        RECT 218.200 172.800 218.600 173.200 ;
        RECT 207.000 172.200 207.300 172.800 ;
        RECT 205.400 172.100 205.800 172.200 ;
        RECT 206.200 172.100 206.600 172.200 ;
        RECT 205.400 171.800 206.600 172.100 ;
        RECT 207.000 171.800 207.400 172.200 ;
        RECT 210.200 171.800 210.600 172.200 ;
        RECT 216.600 171.800 217.000 172.200 ;
        RECT 202.200 170.800 202.600 171.200 ;
        RECT 195.800 169.100 196.200 169.200 ;
        RECT 196.600 169.100 197.000 169.200 ;
        RECT 195.800 168.800 197.000 169.100 ;
        RECT 199.000 168.800 199.400 169.200 ;
        RECT 205.400 168.800 205.800 169.200 ;
        RECT 205.400 168.200 205.700 168.800 ;
        RECT 196.600 167.800 197.000 168.200 ;
        RECT 205.400 167.800 205.800 168.200 ;
        RECT 196.600 167.200 196.900 167.800 ;
        RECT 196.600 166.800 197.000 167.200 ;
        RECT 199.000 166.800 199.400 167.200 ;
        RECT 199.800 166.800 200.200 167.200 ;
        RECT 203.000 167.100 203.400 167.200 ;
        RECT 203.800 167.100 204.200 167.200 ;
        RECT 203.000 166.800 204.200 167.100 ;
        RECT 194.200 165.800 194.600 166.200 ;
        RECT 195.000 166.100 195.400 166.200 ;
        RECT 195.800 166.100 196.200 166.200 ;
        RECT 195.000 165.800 196.200 166.100 ;
        RECT 194.200 165.200 194.500 165.800 ;
        RECT 194.200 164.800 194.600 165.200 ;
        RECT 195.000 165.100 195.400 165.200 ;
        RECT 195.800 165.100 196.200 165.200 ;
        RECT 195.000 164.800 196.200 165.100 ;
        RECT 196.600 163.200 196.900 166.800 ;
        RECT 193.400 162.800 193.800 163.200 ;
        RECT 196.600 162.800 197.000 163.200 ;
        RECT 188.600 159.800 189.000 160.200 ;
        RECT 191.800 159.100 192.200 159.200 ;
        RECT 192.600 159.100 193.000 159.200 ;
        RECT 191.800 158.800 193.000 159.100 ;
        RECT 193.400 158.200 193.700 162.800 ;
        RECT 199.000 162.200 199.300 166.800 ;
        RECT 199.800 166.200 200.100 166.800 ;
        RECT 199.800 165.800 200.200 166.200 ;
        RECT 200.600 165.800 201.000 166.200 ;
        RECT 201.400 166.100 201.800 166.200 ;
        RECT 202.200 166.100 202.600 166.200 ;
        RECT 201.400 165.800 202.600 166.100 ;
        RECT 199.800 164.200 200.100 165.800 ;
        RECT 200.600 165.200 200.900 165.800 ;
        RECT 200.600 164.800 201.000 165.200 ;
        RECT 199.800 163.800 200.200 164.200 ;
        RECT 207.800 163.100 208.200 168.900 ;
        RECT 210.200 167.200 210.500 171.800 ;
        RECT 216.600 170.200 216.900 171.800 ;
        RECT 216.600 169.800 217.000 170.200 ;
        RECT 210.200 166.800 210.600 167.200 ;
        RECT 211.800 166.800 212.200 167.200 ;
        RECT 211.800 166.300 212.100 166.800 ;
        RECT 211.800 165.900 212.200 166.300 ;
        RECT 211.000 163.800 211.400 164.200 ;
        RECT 211.800 163.800 212.200 164.200 ;
        RECT 199.000 161.800 199.400 162.200 ;
        RECT 202.200 161.800 202.600 162.200 ;
        RECT 205.400 161.800 205.800 162.200 ;
        RECT 201.400 158.800 201.800 159.200 ;
        RECT 186.200 156.800 186.600 157.200 ;
        RECT 186.200 155.100 186.600 155.200 ;
        RECT 187.000 155.100 187.400 155.200 ;
        RECT 186.200 154.800 187.400 155.100 ;
        RECT 187.000 153.800 187.400 154.200 ;
        RECT 187.000 152.200 187.300 153.800 ;
        RECT 187.000 151.800 187.400 152.200 ;
        RECT 189.400 152.100 189.800 157.900 ;
        RECT 193.400 157.800 193.800 158.200 ;
        RECT 195.800 157.800 196.200 158.200 ;
        RECT 193.400 155.200 193.700 157.800 ;
        RECT 195.000 156.800 195.400 157.200 ;
        RECT 195.000 156.200 195.300 156.800 ;
        RECT 195.000 155.800 195.400 156.200 ;
        RECT 193.400 154.800 193.800 155.200 ;
        RECT 194.200 155.100 194.600 155.200 ;
        RECT 195.000 155.100 195.400 155.200 ;
        RECT 194.200 154.800 195.400 155.100 ;
        RECT 195.800 154.200 196.100 157.800 ;
        RECT 201.400 157.200 201.700 158.800 ;
        RECT 202.200 158.200 202.500 161.800 ;
        RECT 202.200 157.800 202.600 158.200 ;
        RECT 201.400 156.800 201.800 157.200 ;
        RECT 205.400 156.200 205.700 161.800 ;
        RECT 200.600 155.800 201.000 156.200 ;
        RECT 201.400 155.800 201.800 156.200 ;
        RECT 205.400 155.800 205.800 156.200 ;
        RECT 207.800 155.800 208.200 156.200 ;
        RECT 200.600 155.200 200.900 155.800 ;
        RECT 201.400 155.200 201.700 155.800 ;
        RECT 207.800 155.200 208.100 155.800 ;
        RECT 211.000 155.200 211.300 163.800 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 200.600 154.800 201.000 155.200 ;
        RECT 201.400 154.800 201.800 155.200 ;
        RECT 203.000 155.100 203.400 155.200 ;
        RECT 202.200 154.800 203.400 155.100 ;
        RECT 204.600 154.800 205.000 155.200 ;
        RECT 206.200 155.100 206.600 155.200 ;
        RECT 207.000 155.100 207.400 155.200 ;
        RECT 206.200 154.800 207.400 155.100 ;
        RECT 207.800 154.800 208.200 155.200 ;
        RECT 208.600 154.800 209.000 155.200 ;
        RECT 211.000 154.800 211.400 155.200 ;
        RECT 192.600 153.800 193.000 154.200 ;
        RECT 195.800 153.800 196.200 154.200 ;
        RECT 191.800 151.800 192.200 152.200 ;
        RECT 187.000 149.800 187.400 150.200 ;
        RECT 187.000 149.200 187.300 149.800 ;
        RECT 183.000 148.800 183.400 149.200 ;
        RECT 187.000 148.800 187.400 149.200 ;
        RECT 183.000 148.200 183.300 148.800 ;
        RECT 183.000 147.800 183.400 148.200 ;
        RECT 182.200 144.800 182.600 145.200 ;
        RECT 177.400 142.800 177.800 143.200 ;
        RECT 175.000 141.800 175.400 142.200 ;
        RECT 179.000 142.100 179.400 142.200 ;
        RECT 179.800 142.100 180.200 142.200 ;
        RECT 179.000 141.800 180.200 142.100 ;
        RECT 175.000 135.100 175.300 141.800 ;
        RECT 183.000 141.200 183.300 147.800 ;
        RECT 185.400 146.800 185.800 147.200 ;
        RECT 185.400 146.200 185.700 146.800 ;
        RECT 183.800 145.800 184.200 146.200 ;
        RECT 185.400 145.800 185.800 146.200 ;
        RECT 183.000 140.800 183.400 141.200 ;
        RECT 179.000 139.800 179.400 140.200 ;
        RECT 175.000 134.700 175.400 135.100 ;
        RECT 174.200 133.800 174.600 134.200 ;
        RECT 175.800 132.100 176.200 137.900 ;
        RECT 176.600 133.800 177.000 134.200 ;
        RECT 175.800 130.800 176.200 131.200 ;
        RECT 175.800 129.200 176.100 130.800 ;
        RECT 175.800 128.800 176.200 129.200 ;
        RECT 173.400 125.800 173.800 126.200 ;
        RECT 176.600 124.200 176.900 133.800 ;
        RECT 177.400 133.100 177.800 135.900 ;
        RECT 178.200 135.800 178.600 136.200 ;
        RECT 178.200 135.200 178.500 135.800 ;
        RECT 179.000 135.200 179.300 139.800 ;
        RECT 182.200 137.800 182.600 138.200 ;
        RECT 178.200 134.800 178.600 135.200 ;
        RECT 179.000 134.800 179.400 135.200 ;
        RECT 180.600 131.800 181.000 132.200 ;
        RECT 181.400 131.800 181.800 132.200 ;
        RECT 180.600 131.200 180.900 131.800 ;
        RECT 180.600 130.800 181.000 131.200 ;
        RECT 180.600 127.800 181.000 128.200 ;
        RECT 180.600 127.200 180.900 127.800 ;
        RECT 180.600 126.800 181.000 127.200 ;
        RECT 178.200 125.800 178.600 126.200 ;
        RECT 179.000 125.800 179.400 126.200 ;
        RECT 180.600 125.800 181.000 126.200 ;
        RECT 178.200 125.200 178.500 125.800 ;
        RECT 178.200 124.800 178.600 125.200 ;
        RECT 179.000 125.100 179.300 125.800 ;
        RECT 180.600 125.100 180.900 125.800 ;
        RECT 179.000 124.800 180.900 125.100 ;
        RECT 176.600 123.800 177.000 124.200 ;
        RECT 175.800 121.800 176.200 122.200 ;
        RECT 173.400 111.800 173.800 112.200 ;
        RECT 173.400 110.100 173.700 111.800 ;
        RECT 174.200 110.100 174.600 110.200 ;
        RECT 173.400 109.800 174.600 110.100 ;
        RECT 173.400 103.100 173.800 108.900 ;
        RECT 175.800 97.200 176.100 121.800 ;
        RECT 179.000 113.800 179.400 114.200 ;
        RECT 177.400 108.800 177.800 109.200 ;
        RECT 177.400 106.300 177.700 108.800 ;
        RECT 177.400 105.900 177.800 106.300 ;
        RECT 178.200 103.100 178.600 108.900 ;
        RECT 179.000 108.200 179.300 113.800 ;
        RECT 179.000 107.800 179.400 108.200 ;
        RECT 179.000 107.200 179.300 107.800 ;
        RECT 179.000 106.800 179.400 107.200 ;
        RECT 179.800 105.100 180.200 107.900 ;
        RECT 180.600 106.800 181.000 107.200 ;
        RECT 180.600 104.200 180.900 106.800 ;
        RECT 181.400 105.100 181.700 131.800 ;
        RECT 182.200 129.200 182.500 137.800 ;
        RECT 183.800 137.200 184.100 145.800 ;
        RECT 189.400 143.100 189.800 148.900 ;
        RECT 191.800 148.200 192.100 151.800 ;
        RECT 192.600 151.200 192.900 153.800 ;
        RECT 192.600 150.800 193.000 151.200 ;
        RECT 192.600 148.200 192.900 150.800 ;
        RECT 191.800 147.800 192.200 148.200 ;
        RECT 192.600 147.800 193.000 148.200 ;
        RECT 191.800 147.200 192.100 147.800 ;
        RECT 191.800 146.800 192.200 147.200 ;
        RECT 183.800 136.800 184.200 137.200 ;
        RECT 183.800 135.800 184.200 136.200 ;
        RECT 183.800 133.200 184.100 135.800 ;
        RECT 183.800 132.800 184.200 133.200 ;
        RECT 184.600 133.100 185.000 135.900 ;
        RECT 186.200 132.100 186.600 137.900 ;
        RECT 187.000 134.700 187.400 135.100 ;
        RECT 190.200 134.800 190.600 135.200 ;
        RECT 187.000 131.200 187.300 134.700 ;
        RECT 190.200 131.200 190.500 134.800 ;
        RECT 191.000 132.100 191.400 137.900 ;
        RECT 187.000 130.800 187.400 131.200 ;
        RECT 190.200 130.800 190.600 131.200 ;
        RECT 191.800 131.100 192.100 146.800 ;
        RECT 192.600 146.200 193.000 146.300 ;
        RECT 193.400 146.200 193.800 146.300 ;
        RECT 192.600 145.900 193.800 146.200 ;
        RECT 193.400 144.800 193.800 145.200 ;
        RECT 193.400 137.200 193.700 144.800 ;
        RECT 194.200 143.100 194.600 148.900 ;
        RECT 195.800 145.100 196.200 147.900 ;
        RECT 196.600 144.200 196.900 154.800 ;
        RECT 199.000 153.800 199.400 154.200 ;
        RECT 198.200 151.800 198.600 152.200 ;
        RECT 198.200 146.200 198.500 151.800 ;
        RECT 199.000 150.200 199.300 153.800 ;
        RECT 201.400 152.800 201.800 153.200 ;
        RECT 199.000 149.800 199.400 150.200 ;
        RECT 201.400 147.200 201.700 152.800 ;
        RECT 199.800 146.800 200.200 147.200 ;
        RECT 201.400 146.800 201.800 147.200 ;
        RECT 199.800 146.200 200.100 146.800 ;
        RECT 202.200 146.200 202.500 154.800 ;
        RECT 203.800 153.800 204.200 154.200 ;
        RECT 203.800 153.200 204.100 153.800 ;
        RECT 203.800 152.800 204.200 153.200 ;
        RECT 204.600 149.200 204.900 154.800 ;
        RECT 208.600 153.200 208.900 154.800 ;
        RECT 211.800 154.200 212.100 163.800 ;
        RECT 212.600 163.100 213.000 168.900 ;
        RECT 213.400 168.800 213.800 169.200 ;
        RECT 213.400 167.200 213.700 168.800 ;
        RECT 213.400 166.800 213.800 167.200 ;
        RECT 214.200 165.100 214.600 167.900 ;
        RECT 215.000 167.800 215.400 168.200 ;
        RECT 215.000 167.200 215.300 167.800 ;
        RECT 215.000 166.800 215.400 167.200 ;
        RECT 216.600 166.800 217.000 167.200 ;
        RECT 216.600 166.200 216.900 166.800 ;
        RECT 216.600 165.800 217.000 166.200 ;
        RECT 213.400 162.800 213.800 163.200 ;
        RECT 213.400 154.200 213.700 162.800 ;
        RECT 215.000 156.800 215.400 157.200 ;
        RECT 215.000 155.200 215.300 156.800 ;
        RECT 215.800 155.800 216.200 156.200 ;
        RECT 215.800 155.200 216.100 155.800 ;
        RECT 219.000 155.200 219.300 178.800 ;
        RECT 219.800 175.200 220.100 189.800 ;
        RECT 220.600 183.100 221.000 188.900 ;
        RECT 222.200 186.800 222.600 187.200 ;
        RECT 221.400 185.800 221.800 186.200 ;
        RECT 221.400 179.200 221.700 185.800 ;
        RECT 221.400 178.800 221.800 179.200 ;
        RECT 220.600 175.800 221.000 176.200 ;
        RECT 220.600 175.200 220.900 175.800 ;
        RECT 219.800 174.800 220.200 175.200 ;
        RECT 220.600 174.800 221.000 175.200 ;
        RECT 219.800 171.800 220.200 172.200 ;
        RECT 219.800 166.200 220.100 171.800 ;
        RECT 222.200 169.200 222.500 186.800 ;
        RECT 224.600 186.200 224.900 196.800 ;
        RECT 227.000 195.200 227.300 199.800 ;
        RECT 230.200 196.200 230.500 199.800 ;
        RECT 231.800 196.800 232.200 197.200 ;
        RECT 230.200 195.800 230.600 196.200 ;
        RECT 227.000 194.800 227.400 195.200 ;
        RECT 230.200 194.800 230.600 195.200 ;
        RECT 230.200 194.200 230.500 194.800 ;
        RECT 231.800 194.200 232.100 196.800 ;
        RECT 227.000 193.800 227.400 194.200 ;
        RECT 230.200 193.800 230.600 194.200 ;
        RECT 231.800 193.800 232.200 194.200 ;
        RECT 225.400 191.800 225.800 192.200 ;
        RECT 225.400 191.200 225.700 191.800 ;
        RECT 225.400 190.800 225.800 191.200 ;
        RECT 223.800 185.800 224.200 186.200 ;
        RECT 224.600 185.800 225.000 186.200 ;
        RECT 223.800 177.200 224.100 185.800 ;
        RECT 225.400 183.100 225.800 188.900 ;
        RECT 223.800 176.800 224.200 177.200 ;
        RECT 223.000 174.800 223.400 175.200 ;
        RECT 223.800 174.800 224.200 175.200 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 225.400 175.100 225.800 175.200 ;
        RECT 226.200 175.100 226.600 175.200 ;
        RECT 225.400 174.800 226.600 175.100 ;
        RECT 223.000 174.200 223.300 174.800 ;
        RECT 223.000 173.800 223.400 174.200 ;
        RECT 222.200 168.800 222.600 169.200 ;
        RECT 220.600 166.800 221.000 167.200 ;
        RECT 220.600 166.200 220.900 166.800 ;
        RECT 219.800 165.800 220.200 166.200 ;
        RECT 220.600 165.800 221.000 166.200 ;
        RECT 222.200 165.800 222.600 166.200 ;
        RECT 214.200 154.800 214.600 155.200 ;
        RECT 215.000 154.800 215.400 155.200 ;
        RECT 215.800 154.800 216.200 155.200 ;
        RECT 219.000 154.800 219.400 155.200 ;
        RECT 211.800 153.800 212.200 154.200 ;
        RECT 213.400 153.800 213.800 154.200 ;
        RECT 214.200 153.200 214.500 154.800 ;
        RECT 219.800 154.100 220.100 165.800 ;
        RECT 222.200 162.200 222.500 165.800 ;
        RECT 223.000 164.800 223.400 165.200 ;
        RECT 223.800 165.100 224.100 174.800 ;
        RECT 224.600 174.200 224.900 174.800 ;
        RECT 224.600 173.800 225.000 174.200 ;
        RECT 227.000 172.200 227.300 193.800 ;
        RECT 231.800 187.200 232.100 193.800 ;
        RECT 235.000 192.100 235.400 197.900 ;
        RECT 232.600 189.800 233.000 190.200 ;
        RECT 229.400 186.800 229.800 187.200 ;
        RECT 231.800 186.800 232.200 187.200 ;
        RECT 229.400 186.200 229.700 186.800 ;
        RECT 229.400 185.800 229.800 186.200 ;
        RECT 231.800 186.100 232.200 186.200 ;
        RECT 232.600 186.100 232.900 189.800 ;
        RECT 233.400 187.800 233.800 188.200 ;
        RECT 233.400 187.200 233.700 187.800 ;
        RECT 233.400 186.800 233.800 187.200 ;
        RECT 231.800 185.800 232.900 186.100 ;
        RECT 233.400 185.800 233.800 186.200 ;
        RECT 234.200 185.800 234.600 186.200 ;
        RECT 233.400 185.200 233.700 185.800 ;
        RECT 233.400 184.800 233.800 185.200 ;
        RECT 228.600 183.800 229.000 184.200 ;
        RECT 227.800 181.800 228.200 182.200 ;
        RECT 227.800 175.200 228.100 181.800 ;
        RECT 227.800 174.800 228.200 175.200 ;
        RECT 226.200 171.800 226.600 172.200 ;
        RECT 227.000 171.800 227.400 172.200 ;
        RECT 224.600 166.800 225.000 167.200 ;
        RECT 224.600 166.200 224.900 166.800 ;
        RECT 224.600 165.800 225.000 166.200 ;
        RECT 225.400 165.800 225.800 166.200 ;
        RECT 223.800 164.800 224.900 165.100 ;
        RECT 223.000 164.200 223.300 164.800 ;
        RECT 223.000 163.800 223.400 164.200 ;
        RECT 221.400 161.800 221.800 162.200 ;
        RECT 222.200 161.800 222.600 162.200 ;
        RECT 221.400 159.200 221.700 161.800 ;
        RECT 221.400 158.800 221.800 159.200 ;
        RECT 220.600 156.800 221.000 157.200 ;
        RECT 220.600 155.200 220.900 156.800 ;
        RECT 223.800 155.800 224.200 156.200 ;
        RECT 223.800 155.200 224.100 155.800 ;
        RECT 224.600 155.200 224.900 164.800 ;
        RECT 225.400 156.200 225.700 165.800 ;
        RECT 226.200 163.200 226.500 171.800 ;
        RECT 227.000 165.800 227.400 166.200 ;
        RECT 227.000 163.200 227.300 165.800 ;
        RECT 226.200 162.800 226.600 163.200 ;
        RECT 227.000 162.800 227.400 163.200 ;
        RECT 226.200 161.800 226.600 162.200 ;
        RECT 227.800 161.800 228.200 162.200 ;
        RECT 226.200 159.200 226.500 161.800 ;
        RECT 226.200 158.800 226.600 159.200 ;
        RECT 227.800 157.200 228.100 161.800 ;
        RECT 227.800 156.800 228.200 157.200 ;
        RECT 225.400 155.800 225.800 156.200 ;
        RECT 220.600 154.800 221.000 155.200 ;
        RECT 223.000 154.800 223.400 155.200 ;
        RECT 223.800 154.800 224.200 155.200 ;
        RECT 224.600 154.800 225.000 155.200 ;
        RECT 225.400 154.800 225.800 155.200 ;
        RECT 227.800 154.800 228.200 155.200 ;
        RECT 219.800 153.800 220.900 154.100 ;
        RECT 208.600 152.800 209.000 153.200 ;
        RECT 214.200 152.800 214.600 153.200 ;
        RECT 216.600 153.100 217.000 153.200 ;
        RECT 217.400 153.100 217.800 153.200 ;
        RECT 216.600 152.800 217.800 153.100 ;
        RECT 212.600 151.800 213.000 152.200 ;
        RECT 204.600 148.800 205.000 149.200 ;
        RECT 207.000 147.800 207.400 148.200 ;
        RECT 207.000 147.200 207.300 147.800 ;
        RECT 203.800 146.800 204.200 147.200 ;
        RECT 204.600 147.100 205.000 147.200 ;
        RECT 205.400 147.100 205.800 147.200 ;
        RECT 204.600 146.800 205.800 147.100 ;
        RECT 207.000 146.800 207.400 147.200 ;
        RECT 203.800 146.200 204.100 146.800 ;
        RECT 197.400 145.800 197.800 146.200 ;
        RECT 198.200 145.800 198.600 146.200 ;
        RECT 199.800 145.800 200.200 146.200 ;
        RECT 200.600 145.800 201.000 146.200 ;
        RECT 202.200 145.800 202.600 146.200 ;
        RECT 203.000 145.800 203.400 146.200 ;
        RECT 203.800 145.800 204.200 146.200 ;
        RECT 204.600 145.800 205.000 146.200 ;
        RECT 206.200 145.800 206.600 146.200 ;
        RECT 210.200 145.800 210.600 146.200 ;
        RECT 197.400 145.200 197.700 145.800 ;
        RECT 200.600 145.200 200.900 145.800 ;
        RECT 197.400 144.800 197.800 145.200 ;
        RECT 200.600 144.800 201.000 145.200 ;
        RECT 196.600 143.800 197.000 144.200 ;
        RECT 198.200 141.800 198.600 142.200 ;
        RECT 198.200 141.200 198.500 141.800 ;
        RECT 196.600 140.800 197.000 141.200 ;
        RECT 198.200 140.800 198.600 141.200 ;
        RECT 195.000 139.800 195.400 140.200 ;
        RECT 195.000 139.200 195.300 139.800 ;
        RECT 195.000 138.800 195.400 139.200 ;
        RECT 193.400 136.800 193.800 137.200 ;
        RECT 193.400 136.200 193.700 136.800 ;
        RECT 193.400 135.800 193.800 136.200 ;
        RECT 194.200 135.800 194.600 136.200 ;
        RECT 194.200 134.200 194.500 135.800 ;
        RECT 196.600 135.200 196.900 140.800 ;
        RECT 199.800 135.800 200.200 136.200 ;
        RECT 199.800 135.200 200.100 135.800 ;
        RECT 202.200 135.200 202.500 145.800 ;
        RECT 203.000 145.200 203.300 145.800 ;
        RECT 203.800 145.200 204.100 145.800 ;
        RECT 204.600 145.200 204.900 145.800 ;
        RECT 203.000 144.800 203.400 145.200 ;
        RECT 203.800 144.800 204.200 145.200 ;
        RECT 204.600 144.800 205.000 145.200 ;
        RECT 206.200 142.200 206.500 145.800 ;
        RECT 209.400 144.800 209.800 145.200 ;
        RECT 209.400 144.200 209.700 144.800 ;
        RECT 209.400 143.800 209.800 144.200 ;
        RECT 206.200 141.800 206.600 142.200 ;
        RECT 206.200 141.200 206.500 141.800 ;
        RECT 206.200 140.800 206.600 141.200 ;
        RECT 207.000 139.100 207.400 139.200 ;
        RECT 207.800 139.100 208.200 139.200 ;
        RECT 207.000 138.800 208.200 139.100 ;
        RECT 210.200 137.200 210.500 145.800 ;
        RECT 211.800 143.100 212.200 148.900 ;
        RECT 211.800 140.800 212.200 141.200 ;
        RECT 211.000 139.800 211.400 140.200 ;
        RECT 211.000 137.200 211.300 139.800 ;
        RECT 211.800 139.200 212.100 140.800 ;
        RECT 211.800 138.800 212.200 139.200 ;
        RECT 210.200 136.800 210.600 137.200 ;
        RECT 211.000 136.800 211.400 137.200 ;
        RECT 206.200 136.100 206.600 136.200 ;
        RECT 207.000 136.100 207.400 136.200 ;
        RECT 206.200 135.800 207.400 136.100 ;
        RECT 210.200 135.200 210.500 136.800 ;
        RECT 212.600 136.200 212.900 151.800 ;
        RECT 220.600 149.200 220.900 153.800 ;
        RECT 215.000 146.800 215.400 147.200 ;
        RECT 215.000 146.200 215.300 146.800 ;
        RECT 215.000 145.800 215.400 146.200 ;
        RECT 216.600 143.100 217.000 148.900 ;
        RECT 220.600 148.800 221.000 149.200 ;
        RECT 217.400 147.800 217.800 148.200 ;
        RECT 217.400 147.200 217.700 147.800 ;
        RECT 217.400 146.800 217.800 147.200 ;
        RECT 218.200 145.100 218.600 147.900 ;
        RECT 223.000 147.200 223.300 154.800 ;
        RECT 224.600 152.200 224.900 154.800 ;
        RECT 224.600 151.800 225.000 152.200 ;
        RECT 225.400 151.200 225.700 154.800 ;
        RECT 226.200 151.800 226.600 152.200 ;
        RECT 223.800 150.800 224.200 151.200 ;
        RECT 225.400 150.800 225.800 151.200 ;
        RECT 223.000 146.800 223.400 147.200 ;
        RECT 219.000 145.800 219.400 146.200 ;
        RECT 223.000 145.800 223.400 146.200 ;
        RECT 219.000 145.200 219.300 145.800 ;
        RECT 219.000 144.800 219.400 145.200 ;
        RECT 219.000 141.200 219.300 144.800 ;
        RECT 219.000 140.800 219.400 141.200 ;
        RECT 212.600 135.800 213.000 136.200 ;
        RECT 215.800 136.100 216.200 136.200 ;
        RECT 215.800 135.800 216.900 136.100 ;
        RECT 216.600 135.200 216.900 135.800 ;
        RECT 217.400 135.800 217.800 136.200 ;
        RECT 220.600 135.800 221.000 136.200 ;
        RECT 217.400 135.200 217.700 135.800 ;
        RECT 220.600 135.200 220.900 135.800 ;
        RECT 196.600 134.800 197.000 135.200 ;
        RECT 199.000 134.800 199.400 135.200 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 200.600 135.100 201.000 135.200 ;
        RECT 201.400 135.100 201.800 135.200 ;
        RECT 200.600 134.800 201.800 135.100 ;
        RECT 202.200 134.800 202.600 135.200 ;
        RECT 204.600 135.100 205.000 135.200 ;
        RECT 205.400 135.100 205.800 135.200 ;
        RECT 204.600 134.800 205.800 135.100 ;
        RECT 210.200 134.800 210.600 135.200 ;
        RECT 212.600 134.800 213.000 135.200 ;
        RECT 214.200 134.800 214.600 135.200 ;
        RECT 216.600 134.800 217.000 135.200 ;
        RECT 217.400 134.800 217.800 135.200 ;
        RECT 219.800 134.800 220.200 135.200 ;
        RECT 220.600 134.800 221.000 135.200 ;
        RECT 194.200 133.800 194.600 134.200 ;
        RECT 194.200 133.200 194.500 133.800 ;
        RECT 194.200 132.800 194.600 133.200 ;
        RECT 197.400 133.100 197.800 133.200 ;
        RECT 198.200 133.100 198.600 133.200 ;
        RECT 197.400 132.800 198.600 133.100 ;
        RECT 191.000 130.800 192.100 131.100 ;
        RECT 182.200 128.800 182.600 129.200 ;
        RECT 182.200 128.200 182.500 128.800 ;
        RECT 182.200 127.800 182.600 128.200 ;
        RECT 183.800 126.800 184.200 127.200 ;
        RECT 184.600 126.800 185.000 127.200 ;
        RECT 183.800 126.200 184.100 126.800 ;
        RECT 183.800 125.800 184.200 126.200 ;
        RECT 184.600 125.200 184.900 126.800 ;
        RECT 184.600 124.800 185.000 125.200 ;
        RECT 185.400 125.100 185.800 127.900 ;
        RECT 185.400 123.800 185.800 124.200 ;
        RECT 185.400 122.200 185.700 123.800 ;
        RECT 187.000 123.100 187.400 128.900 ;
        RECT 191.000 127.200 191.300 130.800 ;
        RECT 191.000 126.800 191.400 127.200 ;
        RECT 187.800 125.900 188.200 126.300 ;
        RECT 191.000 126.200 191.300 126.800 ;
        RECT 182.200 121.800 182.600 122.200 ;
        RECT 185.400 121.800 185.800 122.200 ;
        RECT 182.200 121.200 182.500 121.800 ;
        RECT 182.200 120.800 182.600 121.200 ;
        RECT 185.400 119.200 185.700 121.800 ;
        RECT 187.800 121.200 188.100 125.900 ;
        RECT 191.000 125.800 191.400 126.200 ;
        RECT 191.800 123.100 192.200 128.900 ;
        RECT 194.200 128.800 194.600 129.200 ;
        RECT 194.200 128.200 194.500 128.800 ;
        RECT 194.200 127.800 194.600 128.200 ;
        RECT 195.000 126.100 195.400 126.200 ;
        RECT 195.800 126.100 196.200 126.200 ;
        RECT 195.000 125.800 196.200 126.100 ;
        RECT 199.000 124.200 199.300 134.800 ;
        RECT 212.600 134.200 212.900 134.800 ;
        RECT 214.200 134.200 214.500 134.800 ;
        RECT 219.800 134.200 220.100 134.800 ;
        RECT 201.400 133.800 201.800 134.200 ;
        RECT 202.200 134.100 202.600 134.200 ;
        RECT 203.000 134.100 203.400 134.200 ;
        RECT 202.200 133.800 203.400 134.100 ;
        RECT 204.600 133.800 205.000 134.200 ;
        RECT 207.800 134.100 208.200 134.200 ;
        RECT 208.600 134.100 209.000 134.200 ;
        RECT 207.800 133.800 209.000 134.100 ;
        RECT 212.600 133.800 213.000 134.200 ;
        RECT 214.200 133.800 214.600 134.200 ;
        RECT 219.800 133.800 220.200 134.200 ;
        RECT 201.400 133.200 201.700 133.800 ;
        RECT 204.600 133.200 204.900 133.800 ;
        RECT 223.000 133.200 223.300 145.800 ;
        RECT 223.800 139.200 224.100 150.800 ;
        RECT 225.400 146.800 225.800 147.200 ;
        RECT 225.400 146.200 225.700 146.800 ;
        RECT 226.200 146.200 226.500 151.800 ;
        RECT 227.000 150.800 227.400 151.200 ;
        RECT 227.000 147.200 227.300 150.800 ;
        RECT 227.800 150.200 228.100 154.800 ;
        RECT 227.800 149.800 228.200 150.200 ;
        RECT 227.000 146.800 227.400 147.200 ;
        RECT 225.400 145.800 225.800 146.200 ;
        RECT 226.200 145.800 226.600 146.200 ;
        RECT 226.200 143.200 226.500 145.800 ;
        RECT 228.600 145.200 228.900 183.800 ;
        RECT 230.200 181.800 230.600 182.200 ;
        RECT 230.200 179.200 230.500 181.800 ;
        RECT 234.200 181.200 234.500 185.800 ;
        RECT 234.200 180.800 234.600 181.200 ;
        RECT 230.200 178.800 230.600 179.200 ;
        RECT 229.400 177.800 229.800 178.200 ;
        RECT 229.400 166.200 229.700 177.800 ;
        RECT 233.400 176.800 233.800 177.200 ;
        RECT 231.000 176.100 231.400 176.200 ;
        RECT 231.800 176.100 232.200 176.200 ;
        RECT 232.600 176.100 233.000 176.200 ;
        RECT 231.000 175.800 233.000 176.100 ;
        RECT 233.400 175.200 233.700 176.800 ;
        RECT 235.800 176.200 236.100 210.800 ;
        RECT 246.200 210.200 246.500 226.800 ;
        RECT 247.800 221.800 248.200 222.200 ;
        RECT 247.000 212.100 247.400 217.900 ;
        RECT 247.800 216.200 248.100 221.800 ;
        RECT 247.800 215.800 248.200 216.200 ;
        RECT 247.800 214.700 248.200 215.100 ;
        RECT 240.600 209.800 241.000 210.200 ;
        RECT 246.200 210.100 246.600 210.200 ;
        RECT 246.200 209.800 247.300 210.100 ;
        RECT 237.400 203.100 237.800 208.900 ;
        RECT 238.200 207.800 238.600 208.200 ;
        RECT 238.200 207.200 238.500 207.800 ;
        RECT 238.200 206.800 238.600 207.200 ;
        RECT 239.000 205.100 239.400 207.900 ;
        RECT 240.600 206.200 240.900 209.800 ;
        RECT 243.800 206.800 244.200 207.200 ;
        RECT 243.800 206.200 244.100 206.800 ;
        RECT 239.800 205.800 240.200 206.200 ;
        RECT 240.600 205.800 241.000 206.200 ;
        RECT 243.800 205.800 244.200 206.200 ;
        RECT 239.800 205.200 240.100 205.800 ;
        RECT 239.800 204.800 240.200 205.200 ;
        RECT 246.200 201.800 246.600 202.200 ;
        RECT 246.200 199.200 246.500 201.800 ;
        RECT 246.200 198.800 246.600 199.200 ;
        RECT 237.400 195.100 237.800 195.200 ;
        RECT 238.200 195.100 238.600 195.200 ;
        RECT 237.400 194.800 238.600 195.100 ;
        RECT 239.800 192.100 240.200 197.900 ;
        RECT 240.600 193.800 241.000 194.200 ;
        RECT 240.600 192.200 240.900 193.800 ;
        RECT 241.400 193.100 241.800 195.900 ;
        RECT 242.200 194.800 242.600 195.200 ;
        RECT 243.000 194.800 243.400 195.200 ;
        RECT 245.400 195.100 245.800 195.200 ;
        RECT 246.200 195.100 246.600 195.200 ;
        RECT 245.400 194.800 246.600 195.100 ;
        RECT 240.600 191.800 241.000 192.200 ;
        RECT 242.200 192.100 242.500 194.800 ;
        RECT 243.000 194.200 243.300 194.800 ;
        RECT 247.000 194.200 247.300 209.800 ;
        RECT 247.800 199.200 248.100 214.700 ;
        RECT 248.600 203.100 249.000 208.900 ;
        RECT 247.800 198.800 248.200 199.200 ;
        RECT 249.400 196.200 249.700 227.800 ;
        RECT 250.200 197.200 250.500 232.800 ;
        RECT 251.000 232.100 251.400 237.900 ;
        RECT 251.800 233.800 252.200 234.200 ;
        RECT 251.800 233.200 252.100 233.800 ;
        RECT 251.800 232.800 252.200 233.200 ;
        RECT 252.600 233.100 253.000 235.900 ;
        RECT 253.400 235.800 253.800 236.200 ;
        RECT 253.400 234.200 253.700 235.800 ;
        RECT 253.400 233.800 253.800 234.200 ;
        RECT 255.000 233.800 255.400 234.200 ;
        RECT 253.400 231.800 253.800 232.200 ;
        RECT 253.400 228.200 253.700 231.800 ;
        RECT 253.400 227.800 253.800 228.200 ;
        RECT 253.400 227.100 253.800 227.200 ;
        RECT 254.200 227.100 254.600 227.200 ;
        RECT 253.400 226.800 254.600 227.100 ;
        RECT 253.400 225.100 253.800 225.200 ;
        RECT 254.200 225.100 254.600 225.200 ;
        RECT 253.400 224.800 254.600 225.100 ;
        RECT 255.000 223.100 255.300 233.800 ;
        RECT 262.200 232.800 262.600 233.200 ;
        RECT 261.400 231.800 261.800 232.200 ;
        RECT 261.400 227.200 261.700 231.800 ;
        RECT 262.200 229.200 262.500 232.800 ;
        RECT 262.200 228.800 262.600 229.200 ;
        RECT 254.200 222.800 255.300 223.100 ;
        RECT 255.800 226.800 256.200 227.200 ;
        RECT 256.600 226.800 257.000 227.200 ;
        RECT 261.400 226.800 261.800 227.200 ;
        RECT 254.200 219.200 254.500 222.800 ;
        RECT 255.800 222.200 256.100 226.800 ;
        RECT 255.000 221.800 255.400 222.200 ;
        RECT 255.800 221.800 256.200 222.200 ;
        RECT 254.200 218.800 254.600 219.200 ;
        RECT 251.800 212.100 252.200 217.900 ;
        RECT 255.000 217.200 255.300 221.800 ;
        RECT 256.600 221.100 256.900 226.800 ;
        RECT 255.800 220.800 256.900 221.100 ;
        RECT 255.000 216.800 255.400 217.200 ;
        RECT 252.600 212.800 253.000 213.200 ;
        RECT 255.000 213.100 255.400 215.900 ;
        RECT 252.600 211.200 252.900 212.800 ;
        RECT 252.600 210.800 253.000 211.200 ;
        RECT 251.000 206.100 251.400 206.200 ;
        RECT 251.800 206.100 252.200 206.200 ;
        RECT 251.000 205.800 252.200 206.100 ;
        RECT 253.400 203.100 253.800 208.900 ;
        RECT 254.200 206.800 254.600 207.200 ;
        RECT 254.200 202.100 254.500 206.800 ;
        RECT 255.000 205.100 255.400 207.900 ;
        RECT 255.800 207.200 256.100 220.800 ;
        RECT 256.600 212.100 257.000 217.900 ;
        RECT 258.200 215.100 258.600 215.200 ;
        RECT 259.000 215.100 259.400 215.200 ;
        RECT 258.200 214.800 259.400 215.100 ;
        RECT 259.000 213.800 259.400 214.200 ;
        RECT 259.000 211.200 259.300 213.800 ;
        RECT 261.400 212.100 261.800 217.900 ;
        RECT 262.200 214.800 262.600 215.200 ;
        RECT 259.000 210.800 259.400 211.200 ;
        RECT 261.400 210.800 261.800 211.200 ;
        RECT 261.400 209.200 261.700 210.800 ;
        RECT 261.400 208.800 261.800 209.200 ;
        RECT 255.800 206.800 256.200 207.200 ;
        RECT 253.400 201.800 254.500 202.100 ;
        RECT 253.400 197.200 253.700 201.800 ;
        RECT 262.200 199.200 262.500 214.800 ;
        RECT 263.800 211.800 264.200 212.200 ;
        RECT 262.200 198.800 262.600 199.200 ;
        RECT 250.200 196.800 250.600 197.200 ;
        RECT 253.400 196.800 253.800 197.200 ;
        RECT 247.800 195.800 248.200 196.200 ;
        RECT 249.400 195.800 249.800 196.200 ;
        RECT 247.800 195.200 248.100 195.800 ;
        RECT 247.800 194.800 248.200 195.200 ;
        RECT 249.400 195.100 249.800 195.200 ;
        RECT 250.200 195.100 250.600 195.200 ;
        RECT 249.400 194.800 250.600 195.100 ;
        RECT 243.000 193.800 243.400 194.200 ;
        RECT 245.400 194.100 245.800 194.200 ;
        RECT 246.200 194.100 246.600 194.200 ;
        RECT 245.400 193.800 246.600 194.100 ;
        RECT 247.000 193.800 247.400 194.200 ;
        RECT 241.400 191.800 242.500 192.100 ;
        RECT 243.000 192.800 243.400 193.200 ;
        RECT 251.000 192.800 251.400 193.200 ;
        RECT 236.600 186.800 237.000 187.200 ;
        RECT 238.200 186.800 238.600 187.200 ;
        RECT 236.600 186.200 236.900 186.800 ;
        RECT 238.200 186.200 238.500 186.800 ;
        RECT 236.600 185.800 237.000 186.200 ;
        RECT 237.400 185.800 237.800 186.200 ;
        RECT 238.200 185.800 238.600 186.200 ;
        RECT 239.800 185.800 240.200 186.200 ;
        RECT 237.400 185.200 237.700 185.800 ;
        RECT 239.800 185.200 240.100 185.800 ;
        RECT 237.400 184.800 237.800 185.200 ;
        RECT 239.800 184.800 240.200 185.200 ;
        RECT 241.400 183.200 241.700 191.800 ;
        RECT 243.000 191.200 243.300 192.800 ;
        RECT 243.000 190.800 243.400 191.200 ;
        RECT 243.000 187.200 243.300 190.800 ;
        RECT 251.000 190.200 251.300 192.800 ;
        RECT 253.400 191.800 253.800 192.200 ;
        RECT 254.200 192.100 254.600 197.900 ;
        RECT 257.400 194.800 257.800 195.200 ;
        RECT 257.400 194.200 257.700 194.800 ;
        RECT 257.400 193.800 257.800 194.200 ;
        RECT 259.000 192.100 259.400 197.900 ;
        RECT 259.800 193.800 260.200 194.200 ;
        RECT 251.000 189.800 251.400 190.200 ;
        RECT 243.800 188.800 244.200 189.200 ;
        RECT 243.800 187.200 244.100 188.800 ;
        RECT 243.000 186.800 243.400 187.200 ;
        RECT 243.800 186.800 244.200 187.200 ;
        RECT 243.000 186.100 243.400 186.200 ;
        RECT 243.800 186.100 244.200 186.200 ;
        RECT 243.000 185.800 244.200 186.100 ;
        RECT 242.200 185.100 242.600 185.200 ;
        RECT 243.000 185.100 243.400 185.200 ;
        RECT 242.200 184.800 243.400 185.100 ;
        RECT 241.400 182.800 241.800 183.200 ;
        RECT 246.200 183.100 246.600 188.900 ;
        RECT 249.400 185.800 249.800 186.200 ;
        RECT 249.400 185.200 249.700 185.800 ;
        RECT 249.400 184.800 249.800 185.200 ;
        RECT 251.000 183.100 251.400 188.900 ;
        RECT 251.800 187.800 252.200 188.200 ;
        RECT 251.800 187.200 252.100 187.800 ;
        RECT 251.800 186.800 252.200 187.200 ;
        RECT 252.600 185.100 253.000 187.900 ;
        RECT 253.400 187.200 253.700 191.800 ;
        RECT 259.800 187.200 260.100 193.800 ;
        RECT 260.600 193.100 261.000 195.900 ;
        RECT 262.200 194.800 262.600 195.200 ;
        RECT 261.400 193.800 261.800 194.200 ;
        RECT 261.400 193.200 261.700 193.800 ;
        RECT 261.400 192.800 261.800 193.200 ;
        RECT 261.400 191.800 261.800 192.200 ;
        RECT 261.400 189.200 261.700 191.800 ;
        RECT 261.400 188.800 261.800 189.200 ;
        RECT 253.400 186.800 253.800 187.200 ;
        RECT 259.800 186.800 260.200 187.200 ;
        RECT 253.400 184.100 253.700 186.800 ;
        RECT 252.600 183.800 253.700 184.100 ;
        RECT 260.600 184.800 261.000 185.200 ;
        RECT 260.600 184.200 260.900 184.800 ;
        RECT 262.200 184.200 262.500 194.800 ;
        RECT 263.800 187.200 264.100 211.800 ;
        RECT 264.600 195.800 265.000 196.200 ;
        RECT 264.600 192.200 264.900 195.800 ;
        RECT 264.600 191.800 265.000 192.200 ;
        RECT 263.800 186.800 264.200 187.200 ;
        RECT 260.600 183.800 261.000 184.200 ;
        RECT 262.200 183.800 262.600 184.200 ;
        RECT 237.400 180.800 237.800 181.200 ;
        RECT 237.400 177.200 237.700 180.800 ;
        RECT 249.400 179.800 249.800 180.200 ;
        RECT 237.400 176.800 237.800 177.200 ;
        RECT 235.800 175.800 236.200 176.200 ;
        RECT 230.200 175.100 230.600 175.200 ;
        RECT 231.000 175.100 231.400 175.200 ;
        RECT 230.200 174.800 231.400 175.100 ;
        RECT 233.400 174.800 233.800 175.200 ;
        RECT 234.200 174.800 234.600 175.200 ;
        RECT 231.000 174.100 231.400 174.200 ;
        RECT 231.800 174.100 232.200 174.200 ;
        RECT 231.000 173.800 232.200 174.100 ;
        RECT 234.200 172.200 234.500 174.800 ;
        RECT 235.000 173.800 235.400 174.200 ;
        RECT 235.000 173.200 235.300 173.800 ;
        RECT 235.800 173.200 236.100 175.800 ;
        RECT 236.600 174.800 237.000 175.200 ;
        RECT 235.000 172.800 235.400 173.200 ;
        RECT 235.800 172.800 236.200 173.200 ;
        RECT 234.200 171.800 234.600 172.200 ;
        RECT 235.800 171.800 236.200 172.200 ;
        RECT 234.200 169.800 234.600 170.200 ;
        RECT 231.000 168.800 231.400 169.200 ;
        RECT 231.000 166.200 231.300 168.800 ;
        RECT 231.800 166.800 232.200 167.200 ;
        RECT 231.800 166.200 232.100 166.800 ;
        RECT 234.200 166.200 234.500 169.800 ;
        RECT 229.400 165.800 229.800 166.200 ;
        RECT 230.200 165.800 230.600 166.200 ;
        RECT 231.000 165.800 231.400 166.200 ;
        RECT 231.800 165.800 232.200 166.200 ;
        RECT 234.200 165.800 234.600 166.200 ;
        RECT 235.000 165.800 235.400 166.200 ;
        RECT 229.400 163.800 229.800 164.200 ;
        RECT 229.400 153.200 229.700 163.800 ;
        RECT 230.200 160.200 230.500 165.800 ;
        RECT 235.000 165.200 235.300 165.800 ;
        RECT 235.800 165.200 236.100 171.800 ;
        RECT 236.600 167.200 236.900 174.800 ;
        RECT 237.400 174.200 237.700 176.800 ;
        RECT 237.400 173.800 237.800 174.200 ;
        RECT 237.400 171.800 237.800 172.200 ;
        RECT 240.600 172.100 241.000 177.900 ;
        RECT 243.000 175.100 243.400 175.200 ;
        RECT 243.800 175.100 244.200 175.200 ;
        RECT 243.000 174.800 244.200 175.100 ;
        RECT 243.800 173.800 244.200 174.200 ;
        RECT 236.600 166.800 237.000 167.200 ;
        RECT 237.400 166.200 237.700 171.800 ;
        RECT 243.800 171.200 244.100 173.800 ;
        RECT 244.600 172.800 245.000 173.200 ;
        RECT 244.600 172.200 244.900 172.800 ;
        RECT 244.600 171.800 245.000 172.200 ;
        RECT 245.400 172.100 245.800 177.900 ;
        RECT 246.200 175.800 246.600 176.200 ;
        RECT 243.800 170.800 244.200 171.200 ;
        RECT 244.600 170.800 245.000 171.200 ;
        RECT 240.600 168.800 241.000 169.200 ;
        RECT 240.600 168.200 240.900 168.800 ;
        RECT 238.200 167.800 238.600 168.200 ;
        RECT 240.600 167.800 241.000 168.200 ;
        RECT 238.200 167.200 238.500 167.800 ;
        RECT 238.200 166.800 238.600 167.200 ;
        RECT 239.000 166.800 239.400 167.200 ;
        RECT 242.200 167.100 242.600 167.200 ;
        RECT 243.000 167.100 243.400 167.200 ;
        RECT 242.200 166.800 243.400 167.100 ;
        RECT 239.000 166.200 239.300 166.800 ;
        RECT 243.800 166.200 244.100 170.800 ;
        RECT 244.600 170.200 244.900 170.800 ;
        RECT 244.600 169.800 245.000 170.200 ;
        RECT 244.600 167.200 244.900 169.800 ;
        RECT 246.200 169.200 246.500 175.800 ;
        RECT 247.000 173.100 247.400 175.900 ;
        RECT 247.800 175.800 248.200 176.200 ;
        RECT 248.600 175.800 249.000 176.200 ;
        RECT 247.800 175.200 248.100 175.800 ;
        RECT 248.600 175.200 248.900 175.800 ;
        RECT 249.400 175.200 249.700 179.800 ;
        RECT 247.800 174.800 248.200 175.200 ;
        RECT 248.600 174.800 249.000 175.200 ;
        RECT 249.400 174.800 249.800 175.200 ;
        RECT 249.400 174.100 249.800 174.200 ;
        RECT 250.200 174.100 250.600 174.200 ;
        RECT 249.400 173.800 250.600 174.100 ;
        RECT 251.000 171.800 251.400 172.200 ;
        RECT 251.000 171.200 251.300 171.800 ;
        RECT 251.000 170.800 251.400 171.200 ;
        RECT 246.200 168.800 246.600 169.200 ;
        RECT 247.000 168.800 247.400 169.200 ;
        RECT 247.000 168.200 247.300 168.800 ;
        RECT 247.000 167.800 247.400 168.200 ;
        RECT 244.600 166.800 245.000 167.200 ;
        RECT 237.400 165.800 237.800 166.200 ;
        RECT 239.000 166.100 239.400 166.200 ;
        RECT 238.200 165.800 239.400 166.100 ;
        RECT 242.200 166.100 242.600 166.200 ;
        RECT 243.000 166.100 243.400 166.200 ;
        RECT 242.200 165.800 243.400 166.100 ;
        RECT 243.800 165.800 244.200 166.200 ;
        RECT 235.000 164.800 235.400 165.200 ;
        RECT 235.800 164.800 236.200 165.200 ;
        RECT 230.200 159.800 230.600 160.200 ;
        RECT 231.000 157.800 231.400 158.200 ;
        RECT 230.200 155.800 230.600 156.200 ;
        RECT 230.200 155.200 230.500 155.800 ;
        RECT 230.200 154.800 230.600 155.200 ;
        RECT 231.000 154.200 231.300 157.800 ;
        RECT 231.800 154.800 232.200 155.200 ;
        RECT 231.800 154.200 232.100 154.800 ;
        RECT 231.000 153.800 231.400 154.200 ;
        RECT 231.800 153.800 232.200 154.200 ;
        RECT 229.400 152.800 229.800 153.200 ;
        RECT 232.600 153.100 233.000 155.900 ;
        RECT 233.400 153.800 233.800 154.200 ;
        RECT 228.600 144.800 229.000 145.200 ;
        RECT 228.600 144.200 228.900 144.800 ;
        RECT 228.600 143.800 229.000 144.200 ;
        RECT 226.200 142.800 226.600 143.200 ;
        RECT 223.800 138.800 224.200 139.200 ;
        RECT 229.400 138.200 229.700 152.800 ;
        RECT 233.400 148.200 233.700 153.800 ;
        RECT 234.200 152.100 234.600 157.900 ;
        RECT 235.000 155.800 235.400 156.200 ;
        RECT 235.000 155.100 235.300 155.800 ;
        RECT 235.000 154.700 235.400 155.100 ;
        RECT 235.800 150.800 236.200 151.200 ;
        RECT 231.000 147.100 231.400 147.200 ;
        RECT 231.800 147.100 232.200 147.200 ;
        RECT 231.000 146.800 232.200 147.100 ;
        RECT 230.200 145.800 230.600 146.200 ;
        RECT 231.000 145.800 231.400 146.200 ;
        RECT 201.400 132.800 201.800 133.200 ;
        RECT 202.200 133.100 202.600 133.200 ;
        RECT 203.000 133.100 203.400 133.200 ;
        RECT 202.200 132.800 203.400 133.100 ;
        RECT 204.600 132.800 205.000 133.200 ;
        RECT 218.200 133.100 218.600 133.200 ;
        RECT 219.000 133.100 219.400 133.200 ;
        RECT 218.200 132.800 219.400 133.100 ;
        RECT 221.400 133.100 221.800 133.200 ;
        RECT 222.200 133.100 222.600 133.200 ;
        RECT 221.400 132.800 222.600 133.100 ;
        RECT 223.000 132.800 223.400 133.200 ;
        RECT 205.400 131.800 205.800 132.200 ;
        RECT 211.800 131.800 212.200 132.200 ;
        RECT 219.000 131.800 219.400 132.200 ;
        RECT 199.800 130.800 200.200 131.200 ;
        RECT 203.000 130.800 203.400 131.200 ;
        RECT 199.800 127.200 200.100 130.800 ;
        RECT 202.200 127.800 202.600 128.200 ;
        RECT 199.800 126.800 200.200 127.200 ;
        RECT 200.600 127.100 201.000 127.200 ;
        RECT 201.400 127.100 201.800 127.200 ;
        RECT 200.600 126.800 201.800 127.100 ;
        RECT 199.000 123.800 199.400 124.200 ;
        RECT 187.800 120.800 188.200 121.200 ;
        RECT 199.000 120.800 199.400 121.200 ;
        RECT 199.000 119.200 199.300 120.800 ;
        RECT 185.400 118.800 185.800 119.200 ;
        RECT 199.000 118.800 199.400 119.200 ;
        RECT 187.000 113.800 187.400 114.200 ;
        RECT 187.000 112.200 187.300 113.800 ;
        RECT 187.800 112.800 188.200 113.200 ;
        RECT 187.800 112.200 188.100 112.800 ;
        RECT 187.000 111.800 187.400 112.200 ;
        RECT 187.800 111.800 188.200 112.200 ;
        RECT 188.600 111.800 189.000 112.200 ;
        RECT 191.000 112.100 191.400 117.900 ;
        RECT 191.800 115.800 192.200 116.200 ;
        RECT 191.800 115.200 192.100 115.800 ;
        RECT 191.800 114.800 192.200 115.200 ;
        RECT 195.000 114.700 195.400 115.100 ;
        RECT 195.000 113.200 195.300 114.700 ;
        RECT 195.000 112.800 195.400 113.200 ;
        RECT 195.800 112.100 196.200 117.900 ;
        RECT 197.400 113.100 197.800 115.900 ;
        RECT 199.000 111.800 199.400 112.200 ;
        RECT 183.000 108.800 183.400 109.200 ;
        RECT 183.000 108.200 183.300 108.800 ;
        RECT 187.000 108.200 187.300 111.800 ;
        RECT 188.600 108.200 188.900 111.800 ;
        RECT 199.000 111.200 199.300 111.800 ;
        RECT 199.000 110.800 199.400 111.200 ;
        RECT 183.000 107.800 183.400 108.200 ;
        RECT 187.000 107.800 187.400 108.200 ;
        RECT 188.600 107.800 189.000 108.200 ;
        RECT 187.000 106.800 187.400 107.200 ;
        RECT 188.600 106.800 189.000 107.200 ;
        RECT 182.200 105.800 182.600 106.200 ;
        RECT 183.800 106.100 184.200 106.200 ;
        RECT 184.600 106.100 185.000 106.200 ;
        RECT 183.800 105.800 185.000 106.100 ;
        RECT 186.200 105.800 186.600 106.200 ;
        RECT 182.200 105.200 182.500 105.800 ;
        RECT 182.200 105.100 182.600 105.200 ;
        RECT 181.400 104.800 182.600 105.100 ;
        RECT 183.000 104.800 183.400 105.200 ;
        RECT 180.600 103.800 181.000 104.200 ;
        RECT 178.200 101.800 178.600 102.200 ;
        RECT 178.200 99.200 178.500 101.800 ;
        RECT 178.200 98.800 178.600 99.200 ;
        RECT 180.600 98.100 180.900 103.800 ;
        RECT 183.000 99.200 183.300 104.800 ;
        RECT 183.000 98.800 183.400 99.200 ;
        RECT 179.800 97.800 180.900 98.100 ;
        RECT 175.800 96.800 176.200 97.200 ;
        RECT 172.600 95.800 173.000 96.200 ;
        RECT 175.000 95.800 175.400 96.200 ;
        RECT 175.000 95.200 175.300 95.800 ;
        RECT 179.800 95.200 180.100 97.800 ;
        RECT 180.600 95.800 181.000 96.200 ;
        RECT 180.600 95.200 180.900 95.800 ;
        RECT 172.600 94.800 173.000 95.200 ;
        RECT 175.000 95.100 175.400 95.200 ;
        RECT 175.000 94.800 176.100 95.100 ;
        RECT 172.600 94.200 172.900 94.800 ;
        RECT 172.600 93.800 173.000 94.200 ;
        RECT 168.600 92.800 169.000 93.200 ;
        RECT 167.800 90.800 168.200 91.200 ;
        RECT 167.800 89.200 168.100 90.800 ;
        RECT 167.800 88.800 168.200 89.200 ;
        RECT 164.600 86.800 165.000 87.200 ;
        RECT 168.600 86.200 168.900 92.800 ;
        RECT 169.400 86.800 169.800 87.200 ;
        RECT 169.400 86.200 169.700 86.800 ;
        RECT 163.800 85.800 164.200 86.200 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 168.600 85.800 169.000 86.200 ;
        RECT 169.400 85.800 169.800 86.200 ;
        RECT 160.600 84.800 161.000 85.200 ;
        RECT 159.000 82.800 159.400 83.200 ;
        RECT 159.000 79.200 159.300 82.800 ;
        RECT 163.000 80.800 163.400 81.200 ;
        RECT 163.000 79.200 163.300 80.800 ;
        RECT 163.800 79.200 164.100 85.800 ;
        RECT 159.000 78.800 159.400 79.200 ;
        RECT 163.000 78.800 163.400 79.200 ;
        RECT 163.800 78.800 164.200 79.200 ;
        RECT 159.800 77.800 160.200 78.200 ;
        RECT 159.800 76.200 160.100 77.800 ;
        RECT 163.000 76.800 163.400 77.200 ;
        RECT 163.800 76.800 164.200 77.200 ;
        RECT 158.200 75.800 158.600 76.200 ;
        RECT 159.800 75.800 160.200 76.200 ;
        RECT 158.200 74.200 158.500 75.800 ;
        RECT 159.800 74.200 160.100 75.800 ;
        RECT 158.200 73.800 158.600 74.200 ;
        RECT 159.800 73.800 160.200 74.200 ;
        RECT 161.400 74.000 161.800 74.400 ;
        RECT 161.400 72.200 161.700 74.000 ;
        RECT 155.800 71.800 156.200 72.200 ;
        RECT 161.400 71.800 161.800 72.200 ;
        RECT 155.800 69.200 156.100 71.800 ;
        RECT 159.800 70.800 160.200 71.200 ;
        RECT 155.800 68.800 156.200 69.200 ;
        RECT 157.400 68.100 157.800 68.200 ;
        RECT 158.200 68.100 158.600 68.200 ;
        RECT 157.400 67.800 158.600 68.100 ;
        RECT 159.800 66.200 160.100 70.800 ;
        RECT 160.600 68.800 161.000 69.200 ;
        RECT 160.600 67.200 160.900 68.800 ;
        RECT 162.200 67.800 162.600 68.200 ;
        RECT 162.200 67.200 162.500 67.800 ;
        RECT 163.000 67.200 163.300 76.800 ;
        RECT 163.800 76.200 164.100 76.800 ;
        RECT 163.800 75.800 164.200 76.200 ;
        RECT 163.800 73.800 164.200 74.200 ;
        RECT 160.600 66.800 161.000 67.200 ;
        RECT 161.400 66.800 161.800 67.200 ;
        RECT 162.200 66.800 162.600 67.200 ;
        RECT 163.000 66.800 163.400 67.200 ;
        RECT 155.000 65.800 155.400 66.200 ;
        RECT 155.800 65.800 156.200 66.200 ;
        RECT 158.200 65.800 158.600 66.200 ;
        RECT 159.800 65.800 160.200 66.200 ;
        RECT 155.000 63.200 155.300 65.800 ;
        RECT 155.800 64.200 156.100 65.800 ;
        RECT 158.200 65.200 158.500 65.800 ;
        RECT 158.200 64.800 158.600 65.200 ;
        RECT 155.800 63.800 156.200 64.200 ;
        RECT 155.000 62.800 155.400 63.200 ;
        RECT 158.200 60.200 158.500 64.800 ;
        RECT 161.400 62.200 161.700 66.800 ;
        RECT 163.800 66.200 164.100 73.800 ;
        RECT 164.600 69.200 164.900 85.800 ;
        RECT 170.200 85.100 170.600 87.900 ;
        RECT 171.800 83.100 172.200 88.900 ;
        RECT 173.400 88.800 173.800 89.200 ;
        RECT 173.400 87.200 173.700 88.800 ;
        RECT 173.400 86.800 173.800 87.200 ;
        RECT 175.000 86.800 175.400 87.200 ;
        RECT 175.000 86.200 175.300 86.800 ;
        RECT 175.000 85.800 175.400 86.200 ;
        RECT 165.400 81.800 165.800 82.200 ;
        RECT 165.400 79.200 165.700 81.800 ;
        RECT 171.000 79.800 171.400 80.200 ;
        RECT 165.400 78.800 165.800 79.200 ;
        RECT 165.400 75.800 165.800 76.200 ;
        RECT 170.200 75.800 170.600 76.200 ;
        RECT 165.400 75.200 165.700 75.800 ;
        RECT 170.200 75.200 170.500 75.800 ;
        RECT 171.000 75.200 171.300 79.800 ;
        RECT 171.800 77.800 172.200 78.200 ;
        RECT 171.800 75.200 172.100 77.800 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 167.000 74.800 167.400 75.200 ;
        RECT 170.200 74.800 170.600 75.200 ;
        RECT 171.000 74.800 171.400 75.200 ;
        RECT 171.800 74.800 172.200 75.200 ;
        RECT 172.600 74.800 173.000 75.200 ;
        RECT 166.200 74.100 166.600 74.200 ;
        RECT 165.400 73.800 166.600 74.100 ;
        RECT 165.400 69.200 165.700 73.800 ;
        RECT 167.000 73.200 167.300 74.800 ;
        RECT 167.800 74.100 168.200 74.200 ;
        RECT 168.600 74.100 169.000 74.200 ;
        RECT 167.800 73.800 169.000 74.100 ;
        RECT 167.000 72.800 167.400 73.200 ;
        RECT 172.600 69.200 172.900 74.800 ;
        RECT 173.400 71.800 173.800 72.200 ;
        RECT 173.400 71.200 173.700 71.800 ;
        RECT 173.400 70.800 173.800 71.200 ;
        RECT 174.200 69.800 174.600 70.200 ;
        RECT 164.600 68.800 165.000 69.200 ;
        RECT 165.400 68.800 165.800 69.200 ;
        RECT 166.200 68.800 166.600 69.200 ;
        RECT 168.600 69.100 169.000 69.200 ;
        RECT 169.400 69.100 169.800 69.200 ;
        RECT 168.600 68.800 169.800 69.100 ;
        RECT 171.000 69.100 171.400 69.200 ;
        RECT 171.800 69.100 172.200 69.200 ;
        RECT 171.000 68.800 172.200 69.100 ;
        RECT 172.600 68.800 173.000 69.200 ;
        RECT 164.600 67.800 165.000 68.200 ;
        RECT 164.600 67.200 164.900 67.800 ;
        RECT 164.600 66.800 165.000 67.200 ;
        RECT 163.800 65.800 164.200 66.200 ;
        RECT 166.200 65.200 166.500 68.800 ;
        RECT 167.800 67.800 168.200 68.200 ;
        RECT 167.800 67.200 168.100 67.800 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 170.200 66.800 170.600 67.200 ;
        RECT 169.400 66.200 169.700 66.800 ;
        RECT 170.200 66.200 170.500 66.800 ;
        RECT 167.000 66.100 167.400 66.200 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 167.000 65.800 168.200 66.100 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 166.200 64.800 166.600 65.200 ;
        RECT 167.000 63.800 167.400 64.200 ;
        RECT 161.400 61.800 161.800 62.200 ;
        RECT 159.000 60.800 159.400 61.200 ;
        RECT 158.200 59.800 158.600 60.200 ;
        RECT 159.000 59.200 159.300 60.800 ;
        RECT 167.000 59.200 167.300 63.800 ;
        RECT 171.800 62.800 172.200 63.200 ;
        RECT 173.400 63.100 173.800 68.900 ;
        RECT 174.200 66.200 174.500 69.800 ;
        RECT 174.200 65.800 174.600 66.200 ;
        RECT 171.800 59.200 172.100 62.800 ;
        RECT 159.000 58.800 159.400 59.200 ;
        RECT 167.000 58.800 167.400 59.200 ;
        RECT 171.800 58.800 172.200 59.200 ;
        RECT 175.800 58.200 176.100 94.800 ;
        RECT 176.600 94.800 177.000 95.200 ;
        RECT 177.400 94.800 177.800 95.200 ;
        RECT 179.800 94.800 180.200 95.200 ;
        RECT 180.600 94.800 181.000 95.200 ;
        RECT 182.200 94.800 182.600 95.200 ;
        RECT 176.600 94.200 176.900 94.800 ;
        RECT 176.600 93.800 177.000 94.200 ;
        RECT 176.600 92.200 176.900 93.800 ;
        RECT 176.600 91.800 177.000 92.200 ;
        RECT 177.400 89.200 177.700 94.800 ;
        RECT 182.200 91.200 182.500 94.800 ;
        RECT 182.200 90.800 182.600 91.200 ;
        RECT 176.600 83.100 177.000 88.900 ;
        RECT 177.400 88.800 177.800 89.200 ;
        RECT 178.200 89.100 178.600 89.200 ;
        RECT 179.000 89.100 179.400 89.200 ;
        RECT 178.200 88.800 179.400 89.100 ;
        RECT 182.200 87.800 182.600 88.200 ;
        RECT 182.200 87.200 182.500 87.800 ;
        RECT 182.200 86.800 182.600 87.200 ;
        RECT 183.000 86.800 183.400 87.200 ;
        RECT 183.000 86.200 183.300 86.800 ;
        RECT 182.200 85.800 182.600 86.200 ;
        RECT 183.000 85.800 183.400 86.200 ;
        RECT 182.200 85.200 182.500 85.800 ;
        RECT 181.400 84.800 181.800 85.200 ;
        RECT 182.200 84.800 182.600 85.200 ;
        RECT 183.000 84.800 183.400 85.200 ;
        RECT 181.400 84.200 181.700 84.800 ;
        RECT 183.000 84.200 183.300 84.800 ;
        RECT 181.400 83.800 181.800 84.200 ;
        RECT 183.000 83.800 183.400 84.200 ;
        RECT 183.800 80.200 184.100 105.800 ;
        RECT 186.200 103.200 186.500 105.800 ;
        RECT 187.000 104.200 187.300 106.800 ;
        RECT 188.600 106.200 188.900 106.800 ;
        RECT 188.600 105.800 189.000 106.200 ;
        RECT 189.400 105.800 189.800 106.200 ;
        RECT 189.400 104.200 189.700 105.800 ;
        RECT 187.000 103.800 187.400 104.200 ;
        RECT 189.400 103.800 189.800 104.200 ;
        RECT 186.200 102.800 186.600 103.200 ;
        RECT 194.200 103.100 194.600 108.900 ;
        RECT 196.600 106.100 197.000 106.200 ;
        RECT 197.400 106.100 197.800 106.200 ;
        RECT 196.600 105.800 197.800 106.100 ;
        RECT 199.000 103.100 199.400 108.900 ;
        RECT 199.800 107.200 200.100 126.800 ;
        RECT 202.200 126.200 202.500 127.800 ;
        RECT 202.200 125.800 202.600 126.200 ;
        RECT 201.400 114.800 201.800 115.200 ;
        RECT 202.200 114.800 202.600 115.200 ;
        RECT 201.400 114.200 201.700 114.800 ;
        RECT 202.200 114.200 202.500 114.800 ;
        RECT 201.400 113.800 201.800 114.200 ;
        RECT 202.200 113.800 202.600 114.200 ;
        RECT 199.800 106.800 200.200 107.200 ;
        RECT 191.800 101.800 192.200 102.200 ;
        RECT 194.200 101.800 194.600 102.200 ;
        RECT 185.400 96.800 185.800 97.200 ;
        RECT 185.400 95.200 185.700 96.800 ;
        RECT 191.800 95.200 192.100 101.800 ;
        RECT 194.200 99.200 194.500 101.800 ;
        RECT 194.200 98.800 194.600 99.200 ;
        RECT 197.400 98.800 197.800 99.200 ;
        RECT 197.400 98.200 197.700 98.800 ;
        RECT 197.400 97.800 197.800 98.200 ;
        RECT 192.600 96.100 193.000 96.200 ;
        RECT 193.400 96.100 193.800 96.200 ;
        RECT 192.600 95.800 193.800 96.100 ;
        RECT 184.600 94.800 185.000 95.200 ;
        RECT 185.400 94.800 185.800 95.200 ;
        RECT 186.200 94.800 186.600 95.200 ;
        RECT 187.000 95.100 187.400 95.200 ;
        RECT 187.800 95.100 188.200 95.200 ;
        RECT 187.000 94.800 188.200 95.100 ;
        RECT 189.400 94.800 189.800 95.200 ;
        RECT 190.200 94.800 190.600 95.200 ;
        RECT 191.000 94.800 191.400 95.200 ;
        RECT 191.800 94.800 192.200 95.200 ;
        RECT 184.600 94.200 184.900 94.800 ;
        RECT 186.200 94.200 186.500 94.800 ;
        RECT 189.400 94.200 189.700 94.800 ;
        RECT 184.600 93.800 185.000 94.200 ;
        RECT 186.200 93.800 186.600 94.200 ;
        RECT 189.400 93.800 189.800 94.200 ;
        RECT 184.600 91.800 185.000 92.200 ;
        RECT 184.600 86.200 184.900 91.800 ;
        RECT 189.400 89.200 189.700 93.800 ;
        RECT 190.200 92.200 190.500 94.800 ;
        RECT 191.000 94.200 191.300 94.800 ;
        RECT 191.000 93.800 191.400 94.200 ;
        RECT 190.200 91.800 190.600 92.200 ;
        RECT 191.800 91.800 192.200 92.200 ;
        RECT 191.800 90.200 192.100 91.800 ;
        RECT 191.800 89.800 192.200 90.200 ;
        RECT 189.400 88.800 189.800 89.200 ;
        RECT 188.600 88.100 189.000 88.200 ;
        RECT 188.600 87.800 189.700 88.100 ;
        RECT 185.400 86.800 185.800 87.200 ;
        RECT 188.600 86.800 189.000 87.200 ;
        RECT 189.400 87.100 189.700 87.800 ;
        RECT 190.200 87.100 190.600 87.200 ;
        RECT 189.400 86.800 190.600 87.100 ;
        RECT 184.600 85.800 185.000 86.200 ;
        RECT 185.400 83.200 185.700 86.800 ;
        RECT 187.000 86.100 187.400 86.200 ;
        RECT 187.800 86.100 188.200 86.200 ;
        RECT 187.000 85.800 188.200 86.100 ;
        RECT 188.600 85.200 188.900 86.800 ;
        RECT 188.600 84.800 189.000 85.200 ;
        RECT 185.400 82.800 185.800 83.200 ;
        RECT 191.800 83.100 192.200 88.900 ;
        RECT 192.600 86.200 192.900 95.800 ;
        RECT 195.800 95.100 196.200 95.200 ;
        RECT 196.600 95.100 197.000 95.200 ;
        RECT 195.800 94.800 197.000 95.100 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 199.000 95.100 199.400 95.200 ;
        RECT 198.200 94.800 199.400 95.100 ;
        RECT 194.200 91.800 194.600 92.200 ;
        RECT 197.400 91.800 197.800 92.200 ;
        RECT 194.200 91.200 194.500 91.800 ;
        RECT 194.200 90.800 194.600 91.200 ;
        RECT 195.800 89.800 196.200 90.200 ;
        RECT 194.200 88.800 194.600 89.200 ;
        RECT 192.600 85.800 193.000 86.200 ;
        RECT 192.600 83.800 193.000 84.200 ;
        RECT 185.400 81.200 185.700 82.800 ;
        RECT 192.600 82.100 192.900 83.800 ;
        RECT 191.800 81.800 192.900 82.100 ;
        RECT 185.400 80.800 185.800 81.200 ;
        RECT 183.800 79.800 184.200 80.200 ;
        RECT 182.200 78.800 182.600 79.200 ;
        RECT 177.400 74.100 177.800 74.200 ;
        RECT 178.200 74.100 178.600 74.200 ;
        RECT 177.400 73.800 178.600 74.100 ;
        RECT 179.000 72.100 179.400 77.900 ;
        RECT 177.400 66.800 177.800 67.200 ;
        RECT 177.400 66.300 177.700 66.800 ;
        RECT 177.400 65.900 177.800 66.300 ;
        RECT 178.200 63.100 178.600 68.900 ;
        RECT 180.600 68.800 181.000 69.200 ;
        RECT 179.800 65.100 180.200 67.900 ;
        RECT 180.600 67.200 180.900 68.800 ;
        RECT 180.600 66.800 181.000 67.200 ;
        RECT 182.200 66.200 182.500 78.800 ;
        RECT 183.000 74.700 183.400 75.100 ;
        RECT 183.000 72.200 183.300 74.700 ;
        RECT 183.000 71.800 183.400 72.200 ;
        RECT 183.800 72.100 184.200 77.900 ;
        RECT 184.600 73.800 185.000 74.200 ;
        RECT 184.600 73.200 184.900 73.800 ;
        RECT 184.600 72.800 185.000 73.200 ;
        RECT 185.400 73.100 185.800 75.900 ;
        RECT 191.800 75.200 192.100 81.800 ;
        RECT 192.600 75.800 193.000 76.200 ;
        RECT 187.000 75.100 187.400 75.200 ;
        RECT 187.800 75.100 188.200 75.200 ;
        RECT 187.000 74.800 188.200 75.100 ;
        RECT 190.200 74.800 190.600 75.200 ;
        RECT 191.000 74.800 191.400 75.200 ;
        RECT 191.800 74.800 192.200 75.200 ;
        RECT 190.200 74.200 190.500 74.800 ;
        RECT 186.200 73.800 186.600 74.200 ;
        RECT 188.600 74.100 189.000 74.200 ;
        RECT 189.400 74.100 189.800 74.200 ;
        RECT 188.600 73.800 189.800 74.100 ;
        RECT 190.200 73.800 190.600 74.200 ;
        RECT 186.200 73.200 186.500 73.800 ;
        RECT 186.200 72.800 186.600 73.200 ;
        RECT 191.000 72.200 191.300 74.800 ;
        RECT 192.600 74.200 192.900 75.800 ;
        RECT 192.600 73.800 193.000 74.200 ;
        RECT 187.000 71.800 187.400 72.200 ;
        RECT 191.000 71.800 191.400 72.200 ;
        RECT 187.000 69.200 187.300 71.800 ;
        RECT 188.600 70.800 189.000 71.200 ;
        RECT 187.000 68.800 187.400 69.200 ;
        RECT 183.000 67.100 183.400 67.200 ;
        RECT 183.800 67.100 184.200 67.200 ;
        RECT 183.000 66.800 184.200 67.100 ;
        RECT 188.600 66.200 188.900 70.800 ;
        RECT 189.400 69.800 189.800 70.200 ;
        RECT 189.400 67.200 189.700 69.800 ;
        RECT 189.400 66.800 189.800 67.200 ;
        RECT 182.200 65.800 182.600 66.200 ;
        RECT 183.800 66.100 184.200 66.200 ;
        RECT 184.600 66.100 185.000 66.200 ;
        RECT 183.800 65.800 185.000 66.100 ;
        RECT 188.600 65.800 189.000 66.200 ;
        RECT 182.200 65.200 182.500 65.800 ;
        RECT 182.200 64.800 182.600 65.200 ;
        RECT 179.800 61.800 180.200 62.200 ;
        RECT 155.000 52.100 155.400 57.900 ;
        RECT 175.800 57.800 176.200 58.200 ;
        RECT 157.400 56.800 157.800 57.200 ;
        RECT 160.600 56.800 161.000 57.200 ;
        RECT 163.000 56.800 163.400 57.200 ;
        RECT 169.400 56.800 169.800 57.200 ;
        RECT 174.200 56.800 174.600 57.200 ;
        RECT 157.400 56.200 157.700 56.800 ;
        RECT 157.400 55.800 157.800 56.200 ;
        RECT 160.600 55.200 160.900 56.800 ;
        RECT 163.000 56.200 163.300 56.800 ;
        RECT 163.000 55.800 163.400 56.200 ;
        RECT 164.600 55.800 165.000 56.200 ;
        RECT 160.600 54.800 161.000 55.200 ;
        RECT 161.400 55.100 161.800 55.200 ;
        RECT 162.200 55.100 162.600 55.200 ;
        RECT 161.400 54.800 162.600 55.100 ;
        RECT 164.600 54.200 164.900 55.800 ;
        RECT 169.400 55.200 169.700 56.800 ;
        RECT 174.200 55.200 174.500 56.800 ;
        RECT 176.600 55.800 177.000 56.200 ;
        RECT 179.000 55.800 179.400 56.200 ;
        RECT 176.600 55.200 176.900 55.800 ;
        RECT 168.600 54.800 169.000 55.200 ;
        RECT 169.400 54.800 169.800 55.200 ;
        RECT 170.200 55.100 170.600 55.200 ;
        RECT 171.000 55.100 171.400 55.200 ;
        RECT 170.200 54.800 171.400 55.100 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 174.200 54.800 174.600 55.200 ;
        RECT 175.000 54.800 175.400 55.200 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 177.400 55.100 177.800 55.200 ;
        RECT 178.200 55.100 178.600 55.200 ;
        RECT 177.400 54.800 178.600 55.100 ;
        RECT 159.800 53.800 160.200 54.200 ;
        RECT 164.600 53.800 165.000 54.200 ;
        RECT 158.200 49.100 158.600 49.200 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 158.200 48.800 159.400 49.100 ;
        RECT 155.000 47.800 155.400 48.200 ;
        RECT 154.200 38.800 154.600 39.200 ;
        RECT 155.000 39.100 155.300 47.800 ;
        RECT 155.800 46.800 156.200 47.200 ;
        RECT 156.600 46.800 157.000 47.200 ;
        RECT 155.800 46.200 156.100 46.800 ;
        RECT 155.800 45.800 156.200 46.200 ;
        RECT 155.800 44.800 156.200 45.200 ;
        RECT 155.800 44.200 156.100 44.800 ;
        RECT 155.800 43.800 156.200 44.200 ;
        RECT 156.600 43.200 156.900 46.800 ;
        RECT 159.800 43.200 160.100 53.800 ;
        RECT 168.600 51.200 168.900 54.800 ;
        RECT 169.400 54.200 169.700 54.800 ;
        RECT 169.400 53.800 169.800 54.200 ;
        RECT 170.200 53.800 170.600 54.200 ;
        RECT 168.600 50.800 169.000 51.200 ;
        RECT 170.200 49.200 170.500 53.800 ;
        RECT 173.400 53.200 173.700 54.800 ;
        RECT 175.000 53.200 175.300 54.800 ;
        RECT 179.000 54.200 179.300 55.800 ;
        RECT 179.800 55.200 180.100 61.800 ;
        RECT 179.800 54.800 180.200 55.200 ;
        RECT 179.800 54.200 180.100 54.800 ;
        RECT 179.000 53.800 179.400 54.200 ;
        RECT 179.800 53.800 180.200 54.200 ;
        RECT 173.400 52.800 173.800 53.200 ;
        RECT 175.000 52.800 175.400 53.200 ;
        RECT 177.400 52.800 177.800 53.200 ;
        RECT 175.000 52.200 175.300 52.800 ;
        RECT 175.000 51.800 175.400 52.200 ;
        RECT 171.000 50.800 171.400 51.200 ;
        RECT 156.600 42.800 157.000 43.200 ;
        RECT 159.800 42.800 160.200 43.200 ;
        RECT 161.400 43.100 161.800 48.900 ;
        RECT 164.600 45.800 165.000 46.200 ;
        RECT 164.600 45.200 164.900 45.800 ;
        RECT 164.600 44.800 165.000 45.200 ;
        RECT 165.400 42.800 165.800 43.200 ;
        RECT 166.200 43.100 166.600 48.900 ;
        RECT 170.200 48.800 170.600 49.200 ;
        RECT 167.000 47.800 167.400 48.200 ;
        RECT 167.000 47.200 167.300 47.800 ;
        RECT 167.000 46.800 167.400 47.200 ;
        RECT 167.800 45.100 168.200 47.900 ;
        RECT 168.600 45.800 169.000 46.200 ;
        RECT 155.800 39.100 156.200 39.200 ;
        RECT 155.000 38.800 156.200 39.100 ;
        RECT 156.600 38.800 157.000 39.200 ;
        RECT 155.800 38.200 156.100 38.800 ;
        RECT 154.200 37.800 154.600 38.200 ;
        RECT 155.800 37.800 156.200 38.200 ;
        RECT 154.200 34.200 154.500 37.800 ;
        RECT 154.200 33.800 154.600 34.200 ;
        RECT 153.400 32.800 153.800 33.200 ;
        RECT 141.400 30.200 141.700 31.800 ;
        RECT 141.400 29.800 141.800 30.200 ;
        RECT 144.600 29.800 145.000 30.200 ;
        RECT 139.000 29.100 139.400 29.200 ;
        RECT 134.200 26.100 134.600 26.200 ;
        RECT 135.000 26.100 135.400 26.200 ;
        RECT 134.200 25.800 135.400 26.100 ;
        RECT 136.600 23.100 137.000 28.900 ;
        RECT 138.200 28.800 139.400 29.100 ;
        RECT 137.400 26.800 137.800 27.200 ;
        RECT 137.400 26.200 137.700 26.800 ;
        RECT 137.400 25.800 137.800 26.200 ;
        RECT 138.200 25.100 138.600 27.900 ;
        RECT 139.000 23.800 139.400 24.200 ;
        RECT 140.600 23.800 141.000 24.200 ;
        RECT 139.000 19.200 139.300 23.800 ;
        RECT 139.000 18.800 139.400 19.200 ;
        RECT 140.600 15.200 140.900 23.800 ;
        RECT 141.400 23.100 141.800 28.900 ;
        RECT 142.200 26.800 142.600 27.200 ;
        RECT 142.200 26.200 142.500 26.800 ;
        RECT 144.600 26.200 144.900 29.800 ;
        RECT 142.200 25.800 142.600 26.200 ;
        RECT 144.600 25.800 145.000 26.200 ;
        RECT 146.200 23.100 146.600 28.900 ;
        RECT 155.000 28.800 155.400 29.200 ;
        RECT 147.800 25.100 148.200 27.900 ;
        RECT 155.000 27.200 155.300 28.800 ;
        RECT 156.600 28.200 156.900 38.800 ;
        RECT 158.200 33.100 158.600 35.900 ;
        RECT 159.000 33.800 159.400 34.200 ;
        RECT 159.000 32.200 159.300 33.800 ;
        RECT 159.000 31.800 159.400 32.200 ;
        RECT 159.800 32.100 160.200 37.900 ;
        RECT 161.400 34.800 161.800 35.200 ;
        RECT 161.400 33.200 161.700 34.800 ;
        RECT 161.400 32.800 161.800 33.200 ;
        RECT 164.600 32.100 165.000 37.900 ;
        RECT 148.600 26.800 149.000 27.200 ;
        RECT 149.400 26.800 149.800 27.200 ;
        RECT 151.000 26.800 151.400 27.200 ;
        RECT 155.000 26.800 155.400 27.200 ;
        RECT 134.200 14.800 134.600 15.200 ;
        RECT 140.600 14.800 141.000 15.200 ;
        RECT 133.400 13.800 133.800 14.200 ;
        RECT 131.800 7.800 132.200 8.200 ;
        RECT 134.200 7.200 134.500 14.800 ;
        RECT 140.600 14.200 140.900 14.800 ;
        RECT 140.600 13.800 141.000 14.200 ;
        RECT 144.600 13.800 145.000 14.200 ;
        RECT 135.000 9.800 135.400 10.200 ;
        RECT 135.000 9.200 135.300 9.800 ;
        RECT 135.000 8.800 135.400 9.200 ;
        RECT 129.400 6.800 129.800 7.200 ;
        RECT 134.200 6.800 134.600 7.200 ;
        RECT 131.000 5.800 131.400 6.200 ;
        RECT 132.600 5.800 133.000 6.200 ;
        RECT 133.400 6.100 133.800 6.200 ;
        RECT 134.200 6.100 134.600 6.200 ;
        RECT 133.400 5.800 134.600 6.100 ;
        RECT 131.000 5.200 131.300 5.800 ;
        RECT 132.600 5.200 132.900 5.800 ;
        RECT 130.200 5.100 130.600 5.200 ;
        RECT 131.000 5.100 131.400 5.200 ;
        RECT 130.200 4.800 131.400 5.100 ;
        RECT 132.600 4.800 133.000 5.200 ;
        RECT 137.400 3.100 137.800 8.900 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 139.000 5.200 139.300 5.800 ;
        RECT 139.000 4.800 139.400 5.200 ;
        RECT 142.200 3.100 142.600 8.900 ;
        RECT 143.000 7.800 143.400 8.200 ;
        RECT 143.000 7.200 143.300 7.800 ;
        RECT 143.000 6.800 143.400 7.200 ;
        RECT 143.800 5.100 144.200 7.900 ;
        RECT 144.600 7.200 144.900 13.800 ;
        RECT 147.800 13.100 148.200 15.900 ;
        RECT 148.600 15.200 148.900 26.800 ;
        RECT 149.400 26.200 149.700 26.800 ;
        RECT 149.400 25.800 149.800 26.200 ;
        RECT 151.000 25.200 151.300 26.800 ;
        RECT 151.800 25.800 152.200 26.200 ;
        RECT 151.800 25.200 152.100 25.800 ;
        RECT 151.000 24.800 151.400 25.200 ;
        RECT 151.800 24.800 152.200 25.200 ;
        RECT 155.800 25.100 156.200 27.900 ;
        RECT 156.600 27.800 157.000 28.200 ;
        RECT 156.600 27.200 156.900 27.800 ;
        RECT 156.600 26.800 157.000 27.200 ;
        RECT 157.400 23.100 157.800 28.900 ;
        RECT 158.200 25.900 158.600 26.300 ;
        RECT 158.200 25.200 158.500 25.900 ;
        RECT 158.200 24.800 158.600 25.200 ;
        RECT 159.000 24.200 159.300 31.800 ;
        RECT 163.800 29.100 164.200 29.200 ;
        RECT 164.600 29.100 165.000 29.200 ;
        RECT 159.000 23.800 159.400 24.200 ;
        RECT 162.200 23.100 162.600 28.900 ;
        RECT 163.800 28.800 165.000 29.100 ;
        RECT 165.400 27.200 165.700 42.800 ;
        RECT 167.000 39.100 167.400 39.200 ;
        RECT 167.800 39.100 168.200 39.200 ;
        RECT 167.000 38.800 168.200 39.100 ;
        RECT 168.600 38.200 168.900 45.800 ;
        RECT 170.200 39.800 170.600 40.200 ;
        RECT 170.200 39.200 170.500 39.800 ;
        RECT 170.200 38.800 170.600 39.200 ;
        RECT 168.600 37.800 169.000 38.200 ;
        RECT 170.200 37.800 170.600 38.200 ;
        RECT 167.000 35.100 167.400 35.200 ;
        RECT 167.800 35.100 168.200 35.200 ;
        RECT 167.000 34.800 168.200 35.100 ;
        RECT 168.600 34.800 169.000 35.200 ;
        RECT 168.600 34.100 168.900 34.800 ;
        RECT 167.800 33.800 168.900 34.100 ;
        RECT 165.400 26.800 165.800 27.200 ;
        RECT 165.400 26.100 165.800 26.200 ;
        RECT 166.200 26.100 166.600 26.200 ;
        RECT 165.400 25.800 166.600 26.100 ;
        RECT 166.200 24.800 166.600 25.200 ;
        RECT 166.200 24.200 166.500 24.800 ;
        RECT 166.200 23.800 166.600 24.200 ;
        RECT 165.400 19.800 165.800 20.200 ;
        RECT 148.600 14.800 149.000 15.200 ;
        RECT 148.600 13.800 149.000 14.200 ;
        RECT 148.600 13.200 148.900 13.800 ;
        RECT 148.600 12.800 149.000 13.200 ;
        RECT 149.400 12.100 149.800 17.900 ;
        RECT 151.000 14.800 151.400 15.200 ;
        RECT 152.600 14.800 153.000 15.200 ;
        RECT 151.000 13.200 151.300 14.800 ;
        RECT 151.000 12.800 151.400 13.200 ;
        RECT 152.600 9.200 152.900 14.800 ;
        RECT 154.200 12.100 154.600 17.900 ;
        RECT 159.000 17.800 159.400 18.200 ;
        RECT 159.000 15.200 159.300 17.800 ;
        RECT 165.400 16.200 165.700 19.800 ;
        RECT 167.800 19.200 168.100 33.800 ;
        RECT 170.200 31.200 170.500 37.800 ;
        RECT 170.200 30.800 170.600 31.200 ;
        RECT 168.600 25.800 169.000 26.200 ;
        RECT 168.600 25.200 168.900 25.800 ;
        RECT 168.600 24.800 169.000 25.200 ;
        RECT 167.800 18.800 168.200 19.200 ;
        RECT 170.200 19.100 170.500 30.800 ;
        RECT 171.000 29.200 171.300 50.800 ;
        RECT 177.400 49.200 177.700 52.800 ;
        RECT 179.800 52.100 180.200 52.200 ;
        RECT 180.600 52.100 181.000 52.200 ;
        RECT 179.800 51.800 181.000 52.100 ;
        RECT 177.400 48.800 177.800 49.200 ;
        RECT 171.800 46.800 172.200 47.200 ;
        RECT 174.200 47.100 174.600 47.200 ;
        RECT 175.000 47.100 175.400 47.200 ;
        RECT 174.200 46.800 175.400 47.100 ;
        RECT 171.800 43.200 172.100 46.800 ;
        RECT 172.600 45.800 173.000 46.200 ;
        RECT 176.600 45.800 177.000 46.200 ;
        RECT 172.600 45.200 172.900 45.800 ;
        RECT 172.600 44.800 173.000 45.200 ;
        RECT 175.000 45.100 175.400 45.200 ;
        RECT 175.800 45.100 176.200 45.200 ;
        RECT 175.000 44.800 176.200 45.100 ;
        RECT 171.800 42.800 172.200 43.200 ;
        RECT 172.600 38.800 173.000 39.200 ;
        RECT 171.800 34.800 172.200 35.200 ;
        RECT 171.000 28.800 171.400 29.200 ;
        RECT 171.800 22.200 172.100 34.800 ;
        RECT 172.600 33.200 172.900 38.800 ;
        RECT 176.600 36.200 176.900 45.800 ;
        RECT 179.800 43.100 180.200 48.900 ;
        RECT 182.200 45.200 182.500 64.800 ;
        RECT 191.000 63.200 191.300 71.800 ;
        RECT 191.000 62.800 191.400 63.200 ;
        RECT 190.200 58.800 190.600 59.200 ;
        RECT 183.000 52.100 183.400 57.900 ;
        RECT 184.600 55.100 185.000 55.200 ;
        RECT 185.400 55.100 185.800 55.200 ;
        RECT 184.600 54.800 185.800 55.100 ;
        RECT 185.400 53.800 185.800 54.200 ;
        RECT 183.000 46.800 183.400 47.200 ;
        RECT 183.000 46.200 183.300 46.800 ;
        RECT 183.000 45.800 183.400 46.200 ;
        RECT 182.200 44.800 182.600 45.200 ;
        RECT 184.600 43.100 185.000 48.900 ;
        RECT 185.400 48.200 185.700 53.800 ;
        RECT 187.800 52.100 188.200 57.900 ;
        RECT 189.400 53.100 189.800 55.900 ;
        RECT 190.200 55.200 190.500 58.800 ;
        RECT 190.200 54.800 190.600 55.200 ;
        RECT 191.000 54.800 191.400 55.200 ;
        RECT 185.400 47.800 185.800 48.200 ;
        RECT 185.400 47.200 185.700 47.800 ;
        RECT 185.400 46.800 185.800 47.200 ;
        RECT 185.400 44.800 185.800 45.200 ;
        RECT 186.200 45.100 186.600 47.900 ;
        RECT 187.000 45.100 187.400 47.900 ;
        RECT 187.800 46.800 188.200 47.200 ;
        RECT 187.800 45.200 188.100 46.800 ;
        RECT 187.800 44.800 188.200 45.200 ;
        RECT 174.200 35.800 174.600 36.200 ;
        RECT 176.600 35.800 177.000 36.200 ;
        RECT 174.200 35.200 174.500 35.800 ;
        RECT 174.200 34.800 174.600 35.200 ;
        RECT 176.600 34.200 176.900 35.800 ;
        RECT 177.400 34.800 177.800 35.200 ;
        RECT 177.400 34.200 177.700 34.800 ;
        RECT 175.800 33.800 176.200 34.200 ;
        RECT 176.600 33.800 177.000 34.200 ;
        RECT 177.400 33.800 177.800 34.200 ;
        RECT 175.800 33.200 176.100 33.800 ;
        RECT 172.600 32.800 173.000 33.200 ;
        RECT 175.800 32.800 176.200 33.200 ;
        RECT 178.200 33.100 178.600 35.900 ;
        RECT 179.000 33.800 179.400 34.200 ;
        RECT 179.000 32.200 179.300 33.800 ;
        RECT 179.000 31.800 179.400 32.200 ;
        RECT 179.800 32.100 180.200 37.900 ;
        RECT 183.800 35.800 184.200 36.200 ;
        RECT 181.400 35.100 181.800 35.200 ;
        RECT 182.200 35.100 182.600 35.200 ;
        RECT 181.400 34.800 182.600 35.100 ;
        RECT 181.400 29.100 181.800 29.200 ;
        RECT 182.200 29.100 182.600 29.200 ;
        RECT 173.400 23.100 173.800 28.900 ;
        RECT 175.800 25.800 176.200 26.200 ;
        RECT 175.800 24.200 176.100 25.800 ;
        RECT 175.800 23.800 176.200 24.200 ;
        RECT 175.000 22.800 175.400 23.200 ;
        RECT 178.200 23.100 178.600 28.900 ;
        RECT 181.400 28.800 182.600 29.100 ;
        RECT 179.000 26.800 179.400 27.200 ;
        RECT 171.800 21.800 172.200 22.200 ;
        RECT 171.000 19.100 171.400 19.200 ;
        RECT 170.200 18.800 171.400 19.100 ;
        RECT 175.000 16.200 175.300 22.800 ;
        RECT 165.400 15.800 165.800 16.200 ;
        RECT 175.000 15.800 175.400 16.200 ;
        RECT 176.600 16.100 177.000 16.200 ;
        RECT 177.400 16.100 177.800 16.200 ;
        RECT 176.600 15.800 177.800 16.100 ;
        RECT 165.400 15.200 165.700 15.800 ;
        RECT 175.000 15.200 175.300 15.800 ;
        RECT 159.000 14.800 159.400 15.200 ;
        RECT 159.800 15.100 160.200 15.200 ;
        RECT 160.600 15.100 161.000 15.200 ;
        RECT 159.800 14.800 161.000 15.100 ;
        RECT 165.400 14.800 165.800 15.200 ;
        RECT 166.200 14.800 166.600 15.200 ;
        RECT 168.600 14.800 169.000 15.200 ;
        RECT 171.000 14.800 171.400 15.200 ;
        RECT 174.200 14.800 174.600 15.200 ;
        RECT 175.000 14.800 175.400 15.200 ;
        RECT 166.200 14.200 166.500 14.800 ;
        RECT 156.600 13.800 157.000 14.200 ;
        RECT 164.600 13.800 165.000 14.200 ;
        RECT 166.200 13.800 166.600 14.200 ;
        RECT 156.600 12.200 156.900 13.800 ;
        RECT 164.600 13.200 164.900 13.800 ;
        RECT 160.600 13.100 161.000 13.200 ;
        RECT 161.400 13.100 161.800 13.200 ;
        RECT 160.600 12.800 161.800 13.100 ;
        RECT 164.600 12.800 165.000 13.200 ;
        RECT 156.600 11.800 157.000 12.200 ;
        RECT 168.600 9.200 168.900 14.800 ;
        RECT 152.600 8.800 153.000 9.200 ;
        RECT 165.400 9.100 165.800 9.200 ;
        RECT 166.200 9.100 166.600 9.200 ;
        RECT 151.000 7.800 151.400 8.200 ;
        RECT 151.000 7.200 151.300 7.800 ;
        RECT 144.600 6.800 145.000 7.200 ;
        RECT 151.000 6.800 151.400 7.200 ;
        RECT 154.200 6.100 154.600 6.200 ;
        RECT 155.000 6.100 155.400 6.200 ;
        RECT 154.200 5.800 155.400 6.100 ;
        RECT 156.600 5.100 157.000 7.900 ;
        RECT 157.400 7.800 157.800 8.200 ;
        RECT 157.400 7.200 157.700 7.800 ;
        RECT 157.400 6.800 157.800 7.200 ;
        RECT 158.200 3.100 158.600 8.900 ;
        RECT 161.400 7.800 161.800 8.200 ;
        RECT 161.400 6.200 161.700 7.800 ;
        RECT 161.400 5.800 161.800 6.200 ;
        RECT 163.000 3.100 163.400 8.900 ;
        RECT 165.400 8.800 166.600 9.100 ;
        RECT 168.600 8.800 169.000 9.200 ;
        RECT 171.000 8.200 171.300 14.800 ;
        RECT 174.200 14.200 174.500 14.800 ;
        RECT 174.200 13.800 174.600 14.200 ;
        RECT 176.600 14.100 177.000 14.200 ;
        RECT 177.400 14.100 177.800 14.200 ;
        RECT 176.600 13.800 177.800 14.100 ;
        RECT 175.000 9.100 175.400 9.200 ;
        RECT 175.800 9.100 176.200 9.200 ;
        RECT 175.000 8.800 176.200 9.100 ;
        RECT 179.000 8.200 179.300 26.800 ;
        RECT 179.800 25.100 180.200 27.900 ;
        RECT 183.800 26.200 184.100 35.800 ;
        RECT 184.600 32.100 185.000 37.900 ;
        RECT 185.400 37.200 185.700 44.800 ;
        RECT 188.600 43.100 189.000 48.900 ;
        RECT 191.000 37.200 191.300 54.800 ;
        RECT 194.200 54.200 194.500 88.800 ;
        RECT 195.000 86.800 195.400 87.200 ;
        RECT 195.000 86.200 195.300 86.800 ;
        RECT 195.000 85.800 195.400 86.200 ;
        RECT 195.000 78.800 195.400 79.200 ;
        RECT 195.000 75.200 195.300 78.800 ;
        RECT 195.800 78.200 196.100 89.800 ;
        RECT 197.400 89.200 197.700 91.800 ;
        RECT 196.600 83.100 197.000 88.900 ;
        RECT 197.400 88.800 197.800 89.200 ;
        RECT 199.000 88.800 199.400 89.200 ;
        RECT 197.400 86.800 197.800 87.200 ;
        RECT 197.400 86.200 197.700 86.800 ;
        RECT 197.400 85.800 197.800 86.200 ;
        RECT 198.200 85.100 198.600 87.900 ;
        RECT 199.000 87.200 199.300 88.800 ;
        RECT 199.000 86.800 199.400 87.200 ;
        RECT 199.800 87.100 200.100 106.800 ;
        RECT 200.600 105.100 201.000 107.900 ;
        RECT 201.400 106.200 201.700 113.800 ;
        RECT 203.000 109.200 203.300 130.800 ;
        RECT 204.600 127.100 205.000 127.200 ;
        RECT 205.400 127.100 205.700 131.800 ;
        RECT 204.600 126.800 205.700 127.100 ;
        RECT 209.400 128.800 209.800 129.200 ;
        RECT 209.400 126.200 209.700 128.800 ;
        RECT 211.800 126.200 212.100 131.800 ;
        RECT 215.000 127.800 215.400 128.200 ;
        RECT 213.400 126.800 213.800 127.200 ;
        RECT 213.400 126.200 213.700 126.800 ;
        RECT 204.600 126.100 205.000 126.200 ;
        RECT 205.400 126.100 205.800 126.200 ;
        RECT 204.600 125.800 205.800 126.100 ;
        RECT 209.400 125.800 209.800 126.200 ;
        RECT 210.200 126.100 210.600 126.200 ;
        RECT 211.000 126.100 211.400 126.200 ;
        RECT 210.200 125.800 211.400 126.100 ;
        RECT 211.800 125.800 212.200 126.200 ;
        RECT 213.400 125.800 213.800 126.200 ;
        RECT 206.200 125.100 206.600 125.200 ;
        RECT 207.000 125.100 207.400 125.200 ;
        RECT 206.200 124.800 207.400 125.100 ;
        RECT 206.200 123.800 206.600 124.200 ;
        RECT 205.400 121.800 205.800 122.200 ;
        RECT 205.400 117.200 205.700 121.800 ;
        RECT 206.200 119.200 206.500 123.800 ;
        RECT 209.400 120.200 209.700 125.800 ;
        RECT 209.400 119.800 209.800 120.200 ;
        RECT 211.800 119.800 212.200 120.200 ;
        RECT 211.800 119.200 212.100 119.800 ;
        RECT 215.000 119.200 215.300 127.800 ;
        RECT 215.800 125.100 216.200 127.900 ;
        RECT 217.400 123.100 217.800 128.900 ;
        RECT 219.000 126.200 219.300 131.800 ;
        RECT 223.000 129.200 223.300 132.800 ;
        RECT 226.200 132.100 226.600 137.900 ;
        RECT 229.400 137.800 229.800 138.200 ;
        RECT 230.200 135.100 230.500 145.800 ;
        RECT 231.000 144.200 231.300 145.800 ;
        RECT 232.600 145.100 233.000 147.900 ;
        RECT 233.400 147.800 233.800 148.200 ;
        RECT 233.400 147.200 233.700 147.800 ;
        RECT 233.400 146.800 233.800 147.200 ;
        RECT 231.000 143.800 231.400 144.200 ;
        RECT 230.200 134.700 230.600 135.100 ;
        RECT 227.000 133.800 227.400 134.200 ;
        RECT 227.000 129.200 227.300 133.800 ;
        RECT 231.000 132.100 231.400 137.900 ;
        RECT 231.800 134.800 232.200 135.200 ;
        RECT 231.800 134.200 232.100 134.800 ;
        RECT 231.800 133.800 232.200 134.200 ;
        RECT 232.600 133.100 233.000 135.900 ;
        RECT 233.400 135.200 233.700 146.800 ;
        RECT 234.200 143.100 234.600 148.900 ;
        RECT 235.800 146.200 236.100 150.800 ;
        RECT 235.800 145.800 236.200 146.200 ;
        RECT 233.400 134.800 233.800 135.200 ;
        RECT 233.400 134.200 233.700 134.800 ;
        RECT 233.400 133.800 233.800 134.200 ;
        RECT 219.000 125.800 219.400 126.200 ;
        RECT 221.400 125.800 221.800 126.200 ;
        RECT 218.200 124.800 218.600 125.200 ;
        RECT 206.200 118.800 206.600 119.200 ;
        RECT 211.800 118.800 212.200 119.200 ;
        RECT 215.000 118.800 215.400 119.200 ;
        RECT 208.600 117.800 209.000 118.200 ;
        RECT 205.400 116.800 205.800 117.200 ;
        RECT 207.800 115.800 208.200 116.200 ;
        RECT 207.800 115.200 208.100 115.800 ;
        RECT 208.600 115.200 208.900 117.800 ;
        RECT 215.000 116.200 215.300 118.800 ;
        RECT 212.600 115.800 213.000 116.200 ;
        RECT 215.000 115.800 215.400 116.200 ;
        RECT 203.800 114.800 204.200 115.200 ;
        RECT 205.400 114.800 205.800 115.200 ;
        RECT 207.800 114.800 208.200 115.200 ;
        RECT 208.600 114.800 209.000 115.200 ;
        RECT 211.000 114.800 211.400 115.200 ;
        RECT 203.800 114.200 204.100 114.800 ;
        RECT 205.400 114.200 205.700 114.800 ;
        RECT 203.800 113.800 204.200 114.200 ;
        RECT 205.400 113.800 205.800 114.200 ;
        RECT 210.200 113.800 210.600 114.200 ;
        RECT 210.200 112.200 210.500 113.800 ;
        RECT 210.200 111.800 210.600 112.200 ;
        RECT 205.400 110.800 205.800 111.200 ;
        RECT 205.400 109.200 205.700 110.800 ;
        RECT 203.000 108.800 203.400 109.200 ;
        RECT 205.400 108.800 205.800 109.200 ;
        RECT 210.200 108.200 210.500 111.800 ;
        RECT 204.600 107.800 205.000 108.200 ;
        RECT 206.200 108.100 206.600 108.200 ;
        RECT 207.000 108.100 207.400 108.200 ;
        RECT 206.200 107.800 207.400 108.100 ;
        RECT 210.200 107.800 210.600 108.200 ;
        RECT 204.600 107.200 204.900 107.800 ;
        RECT 204.600 106.800 205.000 107.200 ;
        RECT 201.400 105.800 201.800 106.200 ;
        RECT 206.200 105.800 206.600 106.200 ;
        RECT 208.600 106.100 209.000 106.200 ;
        RECT 209.400 106.100 209.800 106.200 ;
        RECT 208.600 105.800 209.800 106.100 ;
        RECT 201.400 98.200 201.700 105.800 ;
        RECT 206.200 105.200 206.500 105.800 ;
        RECT 206.200 104.800 206.600 105.200 ;
        RECT 207.000 102.800 207.400 103.200 ;
        RECT 203.000 101.800 203.400 102.200 ;
        RECT 201.400 97.800 201.800 98.200 ;
        RECT 201.400 95.200 201.700 97.800 ;
        RECT 201.400 95.100 201.800 95.200 ;
        RECT 202.200 95.100 202.600 95.200 ;
        RECT 201.400 94.800 202.600 95.100 ;
        RECT 200.600 92.800 201.000 93.200 ;
        RECT 200.600 92.200 200.900 92.800 ;
        RECT 200.600 91.800 201.000 92.200 ;
        RECT 200.600 87.100 201.000 87.200 ;
        RECT 199.800 86.800 201.000 87.100 ;
        RECT 199.000 86.200 199.300 86.800 ;
        RECT 199.000 85.800 199.400 86.200 ;
        RECT 198.200 81.800 198.600 82.200 ;
        RECT 198.200 79.200 198.500 81.800 ;
        RECT 200.600 79.200 200.900 86.800 ;
        RECT 198.200 78.800 198.600 79.200 ;
        RECT 200.600 78.800 201.000 79.200 ;
        RECT 195.800 77.800 196.200 78.200 ;
        RECT 195.800 75.200 196.100 77.800 ;
        RECT 196.600 76.800 197.000 77.200 ;
        RECT 196.600 76.200 196.900 76.800 ;
        RECT 196.600 75.800 197.000 76.200 ;
        RECT 195.000 74.800 195.400 75.200 ;
        RECT 195.800 74.800 196.200 75.200 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 198.200 75.100 198.600 75.200 ;
        RECT 197.400 74.800 198.600 75.100 ;
        RECT 198.200 74.100 198.600 74.200 ;
        RECT 199.000 74.100 199.400 74.200 ;
        RECT 198.200 73.800 199.400 74.100 ;
        RECT 199.800 73.800 200.200 74.200 ;
        RECT 200.600 73.800 201.000 74.200 ;
        RECT 199.800 73.200 200.100 73.800 ;
        RECT 199.800 72.800 200.200 73.200 ;
        RECT 197.400 69.800 197.800 70.200 ;
        RECT 197.400 68.200 197.700 69.800 ;
        RECT 200.600 69.200 200.900 73.800 ;
        RECT 203.000 69.200 203.300 101.800 ;
        RECT 204.600 91.800 205.000 92.200 ;
        RECT 204.600 90.200 204.900 91.800 ;
        RECT 204.600 89.800 205.000 90.200 ;
        RECT 207.000 89.200 207.300 102.800 ;
        RECT 211.000 102.200 211.300 114.800 ;
        RECT 212.600 110.200 212.900 115.800 ;
        RECT 218.200 115.200 218.500 124.800 ;
        RECT 221.400 123.200 221.700 125.800 ;
        RECT 221.400 122.800 221.800 123.200 ;
        RECT 222.200 123.100 222.600 128.900 ;
        RECT 223.000 128.800 223.400 129.200 ;
        RECT 223.800 129.100 224.200 129.200 ;
        RECT 224.600 129.100 225.000 129.200 ;
        RECT 223.800 128.800 225.000 129.100 ;
        RECT 226.200 128.800 226.600 129.200 ;
        RECT 227.000 128.800 227.400 129.200 ;
        RECT 226.200 126.200 226.500 128.800 ;
        RECT 230.200 127.800 230.600 128.200 ;
        RECT 232.600 127.800 233.000 128.200 ;
        RECT 230.200 127.200 230.500 127.800 ;
        RECT 230.200 126.800 230.600 127.200 ;
        RECT 225.400 125.800 225.800 126.200 ;
        RECT 226.200 125.800 226.600 126.200 ;
        RECT 228.600 125.800 229.000 126.200 ;
        RECT 229.400 125.800 229.800 126.200 ;
        RECT 225.400 121.200 225.700 125.800 ;
        RECT 225.400 120.800 225.800 121.200 ;
        RECT 214.200 115.100 214.600 115.200 ;
        RECT 215.000 115.100 215.400 115.200 ;
        RECT 214.200 114.800 215.400 115.100 ;
        RECT 217.400 114.800 217.800 115.200 ;
        RECT 218.200 114.800 218.600 115.200 ;
        RECT 217.400 114.200 217.700 114.800 ;
        RECT 218.200 114.200 218.500 114.800 ;
        RECT 213.400 113.800 213.800 114.200 ;
        RECT 217.400 113.800 217.800 114.200 ;
        RECT 218.200 113.800 218.600 114.200 ;
        RECT 213.400 113.200 213.700 113.800 ;
        RECT 213.400 112.800 213.800 113.200 ;
        RECT 219.000 113.100 219.400 115.900 ;
        RECT 212.600 109.800 213.000 110.200 ;
        RECT 213.400 109.200 213.700 112.800 ;
        RECT 216.600 111.800 217.000 112.200 ;
        RECT 220.600 112.100 221.000 117.900 ;
        RECT 222.200 115.100 222.600 115.200 ;
        RECT 223.000 115.100 223.400 115.200 ;
        RECT 222.200 114.800 223.400 115.100 ;
        RECT 221.400 112.800 221.800 113.200 ;
        RECT 213.400 108.800 213.800 109.200 ;
        RECT 212.600 106.800 213.000 107.200 ;
        RECT 212.600 106.200 212.900 106.800 ;
        RECT 212.600 105.800 213.000 106.200 ;
        RECT 212.600 104.200 212.900 105.800 ;
        RECT 212.600 103.800 213.000 104.200 ;
        RECT 215.800 103.100 216.200 108.900 ;
        RECT 216.600 106.100 216.900 111.800 ;
        RECT 218.200 107.100 218.600 107.200 ;
        RECT 219.000 107.100 219.400 107.200 ;
        RECT 218.200 106.800 219.400 107.100 ;
        RECT 217.400 106.100 217.800 106.200 ;
        RECT 216.600 105.800 217.800 106.100 ;
        RECT 220.600 103.100 221.000 108.900 ;
        RECT 221.400 107.200 221.700 112.800 ;
        RECT 225.400 112.100 225.800 117.900 ;
        RECT 228.600 117.200 228.900 125.800 ;
        RECT 228.600 116.800 229.000 117.200 ;
        RECT 228.600 114.200 228.900 116.800 ;
        RECT 228.600 113.800 229.000 114.200 ;
        RECT 223.000 108.800 223.400 109.200 ;
        RECT 223.000 108.200 223.300 108.800 ;
        RECT 221.400 106.800 221.800 107.200 ;
        RECT 222.200 105.100 222.600 107.900 ;
        RECT 223.000 107.800 223.400 108.200 ;
        RECT 225.400 108.100 225.800 108.200 ;
        RECT 226.200 108.100 226.600 108.200 ;
        RECT 225.400 107.800 226.600 108.100 ;
        RECT 227.800 107.800 228.200 108.200 ;
        RECT 227.800 107.200 228.100 107.800 ;
        RECT 227.800 106.800 228.200 107.200 ;
        RECT 223.000 105.800 223.400 106.200 ;
        RECT 226.200 106.100 226.600 106.200 ;
        RECT 227.000 106.100 227.400 106.200 ;
        RECT 226.200 105.800 227.400 106.100 ;
        RECT 223.000 105.200 223.300 105.800 ;
        RECT 223.000 104.800 223.400 105.200 ;
        RECT 225.400 105.100 225.800 105.200 ;
        RECT 226.200 105.100 226.600 105.200 ;
        RECT 225.400 104.800 226.600 105.100 ;
        RECT 207.800 102.100 208.200 102.200 ;
        RECT 208.600 102.100 209.000 102.200 ;
        RECT 207.800 101.800 209.000 102.100 ;
        RECT 211.000 101.800 211.400 102.200 ;
        RECT 211.800 101.800 212.200 102.200 ;
        RECT 213.400 101.800 213.800 102.200 ;
        RECT 211.800 101.200 212.100 101.800 ;
        RECT 211.800 100.800 212.200 101.200 ;
        RECT 207.800 92.100 208.200 92.200 ;
        RECT 208.600 92.100 209.000 92.200 ;
        RECT 210.200 92.100 210.600 97.900 ;
        RECT 207.800 91.800 209.000 92.100 ;
        RECT 211.800 91.800 212.200 92.200 ;
        RECT 207.000 88.800 207.400 89.200 ;
        RECT 204.600 87.100 205.000 87.200 ;
        RECT 205.400 87.100 205.800 87.200 ;
        RECT 204.600 86.800 205.800 87.100 ;
        RECT 206.200 86.800 206.600 87.200 ;
        RECT 206.200 86.200 206.500 86.800 ;
        RECT 205.400 85.800 205.800 86.200 ;
        RECT 206.200 85.800 206.600 86.200 ;
        RECT 200.600 68.800 201.000 69.200 ;
        RECT 203.000 68.800 203.400 69.200 ;
        RECT 205.400 68.200 205.700 85.800 ;
        RECT 211.800 85.200 212.100 91.800 ;
        RECT 212.600 86.800 213.000 87.200 ;
        RECT 211.800 84.800 212.200 85.200 ;
        RECT 211.800 84.200 212.100 84.800 ;
        RECT 211.800 83.800 212.200 84.200 ;
        RECT 210.200 77.800 210.600 78.200 ;
        RECT 210.200 77.200 210.500 77.800 ;
        RECT 210.200 76.800 210.600 77.200 ;
        RECT 207.800 76.100 208.200 76.200 ;
        RECT 208.600 76.100 209.000 76.200 ;
        RECT 207.800 75.800 209.000 76.100 ;
        RECT 209.400 75.100 209.800 75.200 ;
        RECT 210.200 75.100 210.600 75.200 ;
        RECT 209.400 74.800 210.600 75.100 ;
        RECT 211.000 73.800 211.400 74.200 ;
        RECT 211.000 73.200 211.300 73.800 ;
        RECT 211.000 72.800 211.400 73.200 ;
        RECT 211.800 73.100 212.200 75.900 ;
        RECT 212.600 74.200 212.900 86.800 ;
        RECT 213.400 86.200 213.700 101.800 ;
        RECT 227.800 101.200 228.100 106.800 ;
        RECT 229.400 105.200 229.700 125.800 ;
        RECT 231.800 121.800 232.200 122.200 ;
        RECT 231.800 119.200 232.100 121.800 ;
        RECT 231.800 118.800 232.200 119.200 ;
        RECT 232.600 116.200 232.900 127.800 ;
        RECT 233.400 123.800 233.800 124.200 ;
        RECT 230.200 116.100 230.600 116.200 ;
        RECT 231.000 116.100 231.400 116.200 ;
        RECT 230.200 115.800 231.400 116.100 ;
        RECT 232.600 115.800 233.000 116.200 ;
        RECT 232.600 115.200 232.900 115.800 ;
        RECT 230.200 114.800 230.600 115.200 ;
        RECT 232.600 114.800 233.000 115.200 ;
        RECT 230.200 114.200 230.500 114.800 ;
        RECT 233.400 114.200 233.700 123.800 ;
        RECT 234.200 123.100 234.600 128.900 ;
        RECT 237.400 128.200 237.700 165.800 ;
        RECT 238.200 153.200 238.500 165.800 ;
        RECT 243.000 164.800 243.400 165.200 ;
        RECT 245.400 165.100 245.800 165.200 ;
        RECT 246.200 165.100 246.600 165.200 ;
        RECT 245.400 164.800 246.600 165.100 ;
        RECT 241.400 161.800 241.800 162.200 ;
        RECT 239.800 160.800 240.200 161.200 ;
        RECT 238.200 152.800 238.600 153.200 ;
        RECT 239.000 152.100 239.400 157.900 ;
        RECT 239.000 143.100 239.400 148.900 ;
        RECT 239.800 134.200 240.100 160.800 ;
        RECT 241.400 159.200 241.700 161.800 ;
        RECT 241.400 158.800 241.800 159.200 ;
        RECT 242.200 154.800 242.600 155.200 ;
        RECT 242.200 154.200 242.500 154.800 ;
        RECT 242.200 153.800 242.600 154.200 ;
        RECT 242.200 152.800 242.600 153.200 ;
        RECT 241.400 149.800 241.800 150.200 ;
        RECT 241.400 149.200 241.700 149.800 ;
        RECT 241.400 148.800 241.800 149.200 ;
        RECT 242.200 147.200 242.500 152.800 ;
        RECT 241.400 147.100 241.800 147.200 ;
        RECT 242.200 147.100 242.600 147.200 ;
        RECT 241.400 146.800 242.600 147.100 ;
        RECT 243.000 146.200 243.300 164.800 ;
        RECT 249.400 163.100 249.800 168.900 ;
        RECT 252.600 167.200 252.900 183.800 ;
        RECT 259.000 181.800 259.400 182.200 ;
        RECT 253.400 172.100 253.800 177.900 ;
        RECT 255.800 175.100 256.200 175.200 ;
        RECT 256.600 175.100 257.000 175.200 ;
        RECT 255.800 174.800 257.000 175.100 ;
        RECT 258.200 172.100 258.600 177.900 ;
        RECT 259.000 174.200 259.300 181.800 ;
        RECT 263.800 178.200 264.100 186.800 ;
        RECT 263.800 177.800 264.200 178.200 ;
        RECT 259.000 173.800 259.400 174.200 ;
        RECT 259.800 173.100 260.200 175.900 ;
        RECT 260.600 175.800 261.000 176.200 ;
        RECT 252.600 166.800 253.000 167.200 ;
        RECT 251.000 165.800 251.400 166.200 ;
        RECT 251.800 166.100 252.200 166.200 ;
        RECT 252.600 166.100 253.000 166.200 ;
        RECT 251.800 165.800 253.000 166.100 ;
        RECT 250.200 162.800 250.600 163.200 ;
        RECT 250.200 157.200 250.500 162.800 ;
        RECT 251.000 161.200 251.300 165.800 ;
        RECT 254.200 163.100 254.600 168.900 ;
        RECT 259.000 168.800 259.400 169.200 ;
        RECT 255.800 165.100 256.200 167.900 ;
        RECT 256.600 167.800 257.000 168.200 ;
        RECT 256.600 164.200 256.900 167.800 ;
        RECT 257.400 167.100 257.800 167.200 ;
        RECT 258.200 167.100 258.600 167.200 ;
        RECT 257.400 166.800 258.600 167.100 ;
        RECT 259.000 166.200 259.300 168.800 ;
        RECT 259.000 165.800 259.400 166.200 ;
        RECT 259.800 166.100 260.200 166.200 ;
        RECT 260.600 166.100 260.900 175.800 ;
        RECT 261.400 171.800 261.800 172.200 ;
        RECT 261.400 169.200 261.700 171.800 ;
        RECT 261.400 168.800 261.800 169.200 ;
        RECT 259.800 165.800 260.900 166.100 ;
        RECT 256.600 163.800 257.000 164.200 ;
        RECT 256.600 161.800 257.000 162.200 ;
        RECT 251.000 160.800 251.400 161.200 ;
        RECT 250.200 156.800 250.600 157.200 ;
        RECT 255.000 157.100 255.400 157.200 ;
        RECT 255.800 157.100 256.200 157.200 ;
        RECT 255.000 156.800 256.200 157.100 ;
        RECT 246.200 155.800 246.600 156.200 ;
        RECT 246.200 155.200 246.500 155.800 ;
        RECT 246.200 154.800 246.600 155.200 ;
        RECT 248.600 155.100 249.000 155.200 ;
        RECT 249.400 155.100 249.800 155.200 ;
        RECT 248.600 154.800 249.800 155.100 ;
        RECT 250.200 154.200 250.500 156.800 ;
        RECT 251.800 155.800 252.200 156.200 ;
        RECT 251.800 155.200 252.100 155.800 ;
        RECT 251.800 154.800 252.200 155.200 ;
        RECT 254.200 155.100 254.600 155.200 ;
        RECT 255.000 155.100 255.400 155.200 ;
        RECT 254.200 154.800 255.400 155.100 ;
        RECT 244.600 153.800 245.000 154.200 ;
        RECT 248.600 154.100 249.000 154.200 ;
        RECT 249.400 154.100 249.800 154.200 ;
        RECT 248.600 153.800 249.800 154.100 ;
        RECT 250.200 153.800 250.600 154.200 ;
        RECT 252.600 154.100 253.000 154.200 ;
        RECT 253.400 154.100 253.800 154.200 ;
        RECT 252.600 153.800 253.800 154.100 ;
        RECT 255.000 153.800 255.400 154.200 ;
        RECT 244.600 149.200 244.900 153.800 ;
        RECT 255.000 153.200 255.300 153.800 ;
        RECT 255.000 152.800 255.400 153.200 ;
        RECT 247.000 151.800 247.400 152.200 ;
        RECT 247.000 151.200 247.300 151.800 ;
        RECT 247.000 150.800 247.400 151.200 ;
        RECT 244.600 148.800 245.000 149.200 ;
        RECT 247.000 148.800 247.400 149.200 ;
        RECT 249.400 149.100 249.800 149.200 ;
        RECT 250.200 149.100 250.600 149.200 ;
        RECT 249.400 148.800 250.600 149.100 ;
        RECT 247.000 147.200 247.300 148.800 ;
        RECT 244.600 147.100 245.000 147.200 ;
        RECT 245.400 147.100 245.800 147.200 ;
        RECT 244.600 146.800 245.800 147.100 ;
        RECT 247.000 146.800 247.400 147.200 ;
        RECT 247.000 146.200 247.300 146.800 ;
        RECT 243.000 145.800 243.400 146.200 ;
        RECT 247.000 145.800 247.400 146.200 ;
        RECT 243.000 145.200 243.300 145.800 ;
        RECT 243.000 144.800 243.400 145.200 ;
        RECT 244.600 145.100 245.000 145.200 ;
        RECT 245.400 145.100 245.800 145.200 ;
        RECT 244.600 144.800 245.800 145.100 ;
        RECT 249.400 143.800 249.800 144.200 ;
        RECT 251.800 143.800 252.200 144.200 ;
        RECT 242.200 141.800 242.600 142.200 ;
        RECT 248.600 141.800 249.000 142.200 ;
        RECT 241.400 136.800 241.800 137.200 ;
        RECT 241.400 134.200 241.700 136.800 ;
        RECT 242.200 135.200 242.500 141.800 ;
        RECT 243.000 135.800 243.400 136.200 ;
        RECT 242.200 134.800 242.600 135.200 ;
        RECT 239.800 133.800 240.200 134.200 ;
        RECT 241.400 133.800 241.800 134.200 ;
        RECT 242.200 133.800 242.600 134.200 ;
        RECT 237.400 127.800 237.800 128.200 ;
        RECT 235.000 125.800 235.400 126.200 ;
        RECT 236.600 126.100 237.000 126.200 ;
        RECT 237.400 126.100 237.800 126.200 ;
        RECT 236.600 125.800 237.800 126.100 ;
        RECT 235.000 122.200 235.300 125.800 ;
        RECT 237.400 124.800 237.800 125.200 ;
        RECT 235.000 121.800 235.400 122.200 ;
        RECT 237.400 115.200 237.700 124.800 ;
        RECT 239.000 123.100 239.400 128.900 ;
        RECT 239.800 128.200 240.100 133.800 ;
        RECT 242.200 129.200 242.500 133.800 ;
        RECT 243.000 133.200 243.300 135.800 ;
        RECT 243.000 132.800 243.400 133.200 ;
        RECT 243.800 131.800 244.200 132.200 ;
        RECT 246.200 132.100 246.600 137.900 ;
        RECT 242.200 128.800 242.600 129.200 ;
        RECT 239.800 127.800 240.200 128.200 ;
        RECT 240.600 125.100 241.000 127.900 ;
        RECT 243.800 126.200 244.100 131.800 ;
        RECT 244.600 126.800 245.000 127.200 ;
        RECT 247.800 126.800 248.200 127.200 ;
        RECT 243.800 125.800 244.200 126.200 ;
        RECT 243.800 125.200 244.100 125.800 ;
        RECT 243.800 124.800 244.200 125.200 ;
        RECT 244.600 124.200 244.900 126.800 ;
        RECT 247.800 126.200 248.100 126.800 ;
        RECT 245.400 125.800 245.800 126.200 ;
        RECT 247.800 125.800 248.200 126.200 ;
        RECT 245.400 125.200 245.700 125.800 ;
        RECT 245.400 124.800 245.800 125.200 ;
        RECT 247.000 125.100 247.400 125.200 ;
        RECT 247.800 125.100 248.200 125.200 ;
        RECT 247.000 124.800 248.200 125.100 ;
        RECT 244.600 123.800 245.000 124.200 ;
        RECT 247.000 122.800 247.400 123.200 ;
        RECT 238.200 121.800 238.600 122.200 ;
        RECT 242.200 121.800 242.600 122.200 ;
        RECT 237.400 114.800 237.800 115.200 ;
        RECT 230.200 113.800 230.600 114.200 ;
        RECT 232.600 114.100 233.000 114.200 ;
        RECT 233.400 114.100 233.800 114.200 ;
        RECT 232.600 113.800 233.800 114.100 ;
        RECT 235.000 113.800 235.400 114.200 ;
        RECT 235.800 113.800 236.200 114.200 ;
        RECT 236.600 113.800 237.000 114.200 ;
        RECT 235.000 112.200 235.300 113.800 ;
        RECT 235.800 113.200 236.100 113.800 ;
        RECT 236.600 113.200 236.900 113.800 ;
        RECT 235.800 112.800 236.200 113.200 ;
        RECT 236.600 112.800 237.000 113.200 ;
        RECT 235.000 111.800 235.400 112.200 ;
        RECT 231.000 110.800 231.400 111.200 ;
        RECT 231.000 109.200 231.300 110.800 ;
        RECT 231.000 108.800 231.400 109.200 ;
        RECT 232.600 108.800 233.000 109.200 ;
        RECT 232.600 108.200 232.900 108.800 ;
        RECT 230.200 107.800 230.600 108.200 ;
        RECT 232.600 107.800 233.000 108.200 ;
        RECT 230.200 107.200 230.500 107.800 ;
        RECT 230.200 106.800 230.600 107.200 ;
        RECT 230.200 106.200 230.500 106.800 ;
        RECT 230.200 105.800 230.600 106.200 ;
        RECT 229.400 105.100 229.800 105.200 ;
        RECT 230.200 105.100 230.600 105.200 ;
        RECT 229.400 104.800 230.600 105.100 ;
        RECT 231.800 104.800 232.200 105.200 ;
        RECT 228.600 104.100 229.000 104.200 ;
        RECT 229.400 104.100 229.800 104.200 ;
        RECT 228.600 103.800 229.800 104.100 ;
        RECT 230.200 102.800 230.600 103.200 ;
        RECT 227.800 100.800 228.200 101.200 ;
        RECT 230.200 99.200 230.500 102.800 ;
        RECT 231.000 101.800 231.400 102.200 ;
        RECT 230.200 98.800 230.600 99.200 ;
        RECT 214.200 94.700 214.600 95.100 ;
        RECT 214.200 89.100 214.500 94.700 ;
        RECT 215.000 92.100 215.400 97.900 ;
        RECT 219.000 97.100 219.400 97.200 ;
        RECT 219.800 97.100 220.200 97.200 ;
        RECT 219.000 96.800 220.200 97.100 ;
        RECT 215.800 93.800 216.200 94.200 ;
        RECT 215.800 91.200 216.100 93.800 ;
        RECT 216.600 93.100 217.000 95.900 ;
        RECT 219.800 93.100 220.200 95.900 ;
        RECT 220.600 92.800 221.000 93.200 ;
        RECT 218.200 91.800 218.600 92.200 ;
        RECT 215.800 90.800 216.200 91.200 ;
        RECT 215.000 89.100 215.400 89.200 ;
        RECT 214.200 88.800 215.400 89.100 ;
        RECT 214.200 87.800 214.600 88.200 ;
        RECT 214.200 87.200 214.500 87.800 ;
        RECT 214.200 86.800 214.600 87.200 ;
        RECT 217.400 86.800 217.800 87.200 ;
        RECT 213.400 85.800 213.800 86.200 ;
        RECT 215.800 86.100 216.200 86.200 ;
        RECT 216.600 86.100 217.000 86.200 ;
        RECT 215.800 85.800 217.000 86.100 ;
        RECT 215.000 84.800 215.400 85.200 ;
        RECT 215.000 84.200 215.300 84.800 ;
        RECT 213.400 83.800 213.800 84.200 ;
        RECT 215.000 83.800 215.400 84.200 ;
        RECT 213.400 83.200 213.700 83.800 ;
        RECT 213.400 82.800 213.800 83.200 ;
        RECT 217.400 81.200 217.700 86.800 ;
        RECT 218.200 86.200 218.500 91.800 ;
        RECT 219.800 89.800 220.200 90.200 ;
        RECT 219.800 89.200 220.100 89.800 ;
        RECT 219.800 88.800 220.200 89.200 ;
        RECT 220.600 88.200 220.900 92.800 ;
        RECT 221.400 92.100 221.800 97.900 ;
        RECT 223.000 94.800 223.400 95.200 ;
        RECT 222.200 92.800 222.600 93.200 ;
        RECT 220.600 87.800 221.000 88.200 ;
        RECT 219.000 86.800 219.400 87.200 ;
        RECT 219.000 86.200 219.300 86.800 ;
        RECT 218.200 85.800 218.600 86.200 ;
        RECT 219.000 85.800 219.400 86.200 ;
        RECT 221.400 85.100 221.800 85.200 ;
        RECT 220.600 84.800 221.800 85.100 ;
        RECT 217.400 80.800 217.800 81.200 ;
        RECT 220.600 79.200 220.900 84.800 ;
        RECT 222.200 82.200 222.500 92.800 ;
        RECT 223.000 90.200 223.300 94.800 ;
        RECT 226.200 92.100 226.600 97.900 ;
        RECT 227.000 97.800 227.400 98.200 ;
        RECT 227.000 95.200 227.300 97.800 ;
        RECT 227.800 97.100 228.200 97.200 ;
        RECT 228.600 97.100 229.000 97.200 ;
        RECT 227.800 96.800 229.000 97.100 ;
        RECT 231.000 95.200 231.300 101.800 ;
        RECT 231.800 100.200 232.100 104.800 ;
        RECT 235.000 103.100 235.400 108.900 ;
        RECT 237.400 102.200 237.700 114.800 ;
        RECT 238.200 107.200 238.500 121.800 ;
        RECT 239.000 118.800 239.400 119.200 ;
        RECT 239.000 118.200 239.300 118.800 ;
        RECT 242.200 118.200 242.500 121.800 ;
        RECT 243.000 120.800 243.400 121.200 ;
        RECT 239.000 117.800 239.400 118.200 ;
        RECT 242.200 117.800 242.600 118.200 ;
        RECT 243.000 115.200 243.300 120.800 ;
        RECT 246.200 119.800 246.600 120.200 ;
        RECT 246.200 119.200 246.500 119.800 ;
        RECT 246.200 118.800 246.600 119.200 ;
        RECT 243.800 116.800 244.200 117.200 ;
        RECT 245.400 116.800 245.800 117.200 ;
        RECT 243.000 114.800 243.400 115.200 ;
        RECT 243.800 114.200 244.100 116.800 ;
        RECT 245.400 116.200 245.700 116.800 ;
        RECT 245.400 115.800 245.800 116.200 ;
        RECT 243.800 113.800 244.200 114.200 ;
        RECT 241.400 113.100 241.800 113.200 ;
        RECT 242.200 113.100 242.600 113.200 ;
        RECT 241.400 112.800 242.600 113.100 ;
        RECT 245.400 112.800 245.800 113.200 ;
        RECT 245.400 112.200 245.700 112.800 ;
        RECT 245.400 111.800 245.800 112.200 ;
        RECT 238.200 106.800 238.600 107.200 ;
        RECT 238.200 106.200 238.600 106.300 ;
        RECT 239.000 106.200 239.400 106.300 ;
        RECT 238.200 105.900 239.400 106.200 ;
        RECT 239.800 103.100 240.200 108.900 ;
        RECT 241.400 105.100 241.800 107.900 ;
        RECT 244.600 107.800 245.000 108.200 ;
        RECT 243.000 106.800 243.400 107.200 ;
        RECT 243.000 105.200 243.300 106.800 ;
        RECT 244.600 106.200 244.900 107.800 ;
        RECT 243.800 105.800 244.200 106.200 ;
        RECT 244.600 105.800 245.000 106.200 ;
        RECT 243.800 105.200 244.100 105.800 ;
        RECT 243.000 104.800 243.400 105.200 ;
        RECT 243.800 104.800 244.200 105.200 ;
        RECT 237.400 101.800 237.800 102.200 ;
        RECT 239.800 100.800 240.200 101.200 ;
        RECT 231.800 99.800 232.200 100.200 ;
        RECT 238.200 99.800 238.600 100.200 ;
        RECT 237.400 95.800 237.800 96.200 ;
        RECT 227.000 94.800 227.400 95.200 ;
        RECT 231.000 95.100 231.400 95.200 ;
        RECT 231.800 95.100 232.200 95.200 ;
        RECT 231.000 94.800 232.200 95.100 ;
        RECT 223.000 89.800 223.400 90.200 ;
        RECT 223.800 87.800 224.200 88.200 ;
        RECT 223.800 87.200 224.100 87.800 ;
        RECT 223.800 86.800 224.200 87.200 ;
        RECT 227.000 86.200 227.300 94.800 ;
        RECT 234.200 93.800 234.600 94.200 ;
        RECT 232.600 93.100 233.000 93.200 ;
        RECT 233.400 93.100 233.800 93.200 ;
        RECT 232.600 92.800 233.800 93.100 ;
        RECT 234.200 92.200 234.500 93.800 ;
        RECT 233.400 91.800 233.800 92.200 ;
        RECT 234.200 91.800 234.600 92.200 ;
        RECT 231.800 88.800 232.200 89.200 ;
        RECT 227.800 87.800 228.200 88.200 ;
        RECT 227.800 87.200 228.100 87.800 ;
        RECT 227.800 86.800 228.200 87.200 ;
        RECT 223.000 85.800 223.400 86.200 ;
        RECT 227.000 85.800 227.400 86.200 ;
        RECT 228.600 85.800 229.000 86.200 ;
        RECT 229.400 85.800 229.800 86.200 ;
        RECT 223.000 85.200 223.300 85.800 ;
        RECT 228.600 85.200 228.900 85.800 ;
        RECT 223.000 84.800 223.400 85.200 ;
        RECT 228.600 84.800 229.000 85.200 ;
        RECT 222.200 81.800 222.600 82.200 ;
        RECT 223.000 81.800 223.400 82.200 ;
        RECT 225.400 81.800 225.800 82.200 ;
        RECT 220.600 78.800 221.000 79.200 ;
        RECT 212.600 73.800 213.000 74.200 ;
        RECT 212.600 72.800 213.000 73.200 ;
        RECT 207.000 69.800 207.400 70.200 ;
        RECT 197.400 67.800 197.800 68.200 ;
        RECT 203.800 68.100 204.200 68.200 ;
        RECT 203.000 67.800 204.200 68.100 ;
        RECT 205.400 67.800 205.800 68.200 ;
        RECT 197.400 67.200 197.700 67.800 ;
        RECT 203.000 67.200 203.300 67.800 ;
        RECT 205.400 67.200 205.700 67.800 ;
        RECT 207.000 67.200 207.300 69.800 ;
        RECT 212.600 69.200 212.900 72.800 ;
        RECT 213.400 72.100 213.800 77.900 ;
        RECT 215.800 75.100 216.200 75.200 ;
        RECT 216.600 75.100 217.000 75.200 ;
        RECT 215.800 74.800 217.000 75.100 ;
        RECT 218.200 72.100 218.600 77.900 ;
        RECT 223.000 76.200 223.300 81.800 ;
        RECT 225.400 81.200 225.700 81.800 ;
        RECT 223.800 80.800 224.200 81.200 ;
        RECT 225.400 80.800 225.800 81.200 ;
        RECT 221.400 76.100 221.800 76.200 ;
        RECT 222.200 76.100 222.600 76.200 ;
        RECT 221.400 75.800 222.600 76.100 ;
        RECT 223.000 75.800 223.400 76.200 ;
        RECT 223.800 75.200 224.100 80.800 ;
        RECT 226.200 79.800 226.600 80.200 ;
        RECT 224.600 77.800 225.000 78.200 ;
        RECT 220.600 75.100 221.000 75.200 ;
        RECT 221.400 75.100 221.800 75.200 ;
        RECT 220.600 74.800 221.800 75.100 ;
        RECT 223.000 74.800 223.400 75.200 ;
        RECT 223.800 74.800 224.200 75.200 ;
        RECT 223.000 72.200 223.300 74.800 ;
        RECT 223.800 74.200 224.100 74.800 ;
        RECT 224.600 74.200 224.900 77.800 ;
        RECT 226.200 76.200 226.500 79.800 ;
        RECT 227.000 76.800 227.400 77.200 ;
        RECT 226.200 75.800 226.600 76.200 ;
        RECT 227.000 75.200 227.300 76.800 ;
        RECT 229.400 76.200 229.700 85.800 ;
        RECT 230.200 84.800 230.600 85.200 ;
        RECT 231.000 85.100 231.400 87.900 ;
        RECT 231.800 87.200 232.100 88.800 ;
        RECT 231.800 86.800 232.200 87.200 ;
        RECT 230.200 83.200 230.500 84.800 ;
        RECT 230.200 82.800 230.600 83.200 ;
        RECT 232.600 83.100 233.000 88.900 ;
        RECT 233.400 86.300 233.700 91.800 ;
        RECT 237.400 90.200 237.700 95.800 ;
        RECT 238.200 95.200 238.500 99.800 ;
        RECT 239.800 99.200 240.100 100.800 ;
        RECT 239.800 98.800 240.200 99.200 ;
        RECT 238.200 95.100 238.600 95.200 ;
        RECT 239.000 95.100 239.400 95.200 ;
        RECT 238.200 94.800 239.400 95.100 ;
        RECT 242.200 92.100 242.600 97.900 ;
        RECT 243.000 94.800 243.400 95.200 ;
        RECT 241.400 90.800 241.800 91.200 ;
        RECT 237.400 89.800 237.800 90.200 ;
        RECT 239.800 89.800 240.200 90.200 ;
        RECT 239.800 89.200 240.100 89.800 ;
        RECT 241.400 89.200 241.700 90.800 ;
        RECT 233.400 85.900 233.800 86.300 ;
        RECT 234.200 82.800 234.600 83.200 ;
        RECT 237.400 83.100 237.800 88.900 ;
        RECT 239.800 88.800 240.200 89.200 ;
        RECT 241.400 88.800 241.800 89.200 ;
        RECT 241.400 84.800 241.800 85.200 ;
        RECT 238.200 83.800 238.600 84.200 ;
        RECT 231.000 81.800 231.400 82.200 ;
        RECT 230.200 76.800 230.600 77.200 ;
        RECT 230.200 76.200 230.500 76.800 ;
        RECT 229.400 75.800 229.800 76.200 ;
        RECT 230.200 75.800 230.600 76.200 ;
        RECT 226.200 74.800 226.600 75.200 ;
        RECT 227.000 74.800 227.400 75.200 ;
        RECT 227.800 74.800 228.200 75.200 ;
        RECT 226.200 74.200 226.500 74.800 ;
        RECT 223.800 73.800 224.200 74.200 ;
        RECT 224.600 73.800 225.000 74.200 ;
        RECT 226.200 73.800 226.600 74.200 ;
        RECT 220.600 71.800 221.000 72.200 ;
        RECT 223.000 71.800 223.400 72.200 ;
        RECT 212.600 68.800 213.000 69.200 ;
        RECT 219.800 68.800 220.200 69.200 ;
        RECT 215.800 68.100 216.200 68.200 ;
        RECT 210.200 67.800 212.900 68.100 ;
        RECT 197.400 66.800 197.800 67.200 ;
        RECT 199.800 66.800 200.200 67.200 ;
        RECT 200.600 67.100 201.000 67.200 ;
        RECT 200.600 66.800 201.700 67.100 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 203.800 66.800 204.200 67.200 ;
        RECT 205.400 66.800 205.800 67.200 ;
        RECT 207.000 66.800 207.400 67.200 ;
        RECT 210.200 67.100 210.500 67.800 ;
        RECT 212.600 67.200 212.900 67.800 ;
        RECT 215.000 67.800 216.200 68.100 ;
        RECT 217.400 67.800 217.800 68.200 ;
        RECT 215.000 67.200 215.300 67.800 ;
        RECT 217.400 67.200 217.700 67.800 ;
        RECT 207.800 66.800 210.500 67.100 ;
        RECT 211.000 66.800 211.400 67.200 ;
        RECT 211.800 66.800 212.200 67.200 ;
        RECT 212.600 66.800 213.000 67.200 ;
        RECT 215.000 66.800 215.400 67.200 ;
        RECT 215.800 66.800 216.200 67.200 ;
        RECT 217.400 66.800 217.800 67.200 ;
        RECT 199.800 66.200 200.100 66.800 ;
        RECT 195.800 66.100 196.200 66.200 ;
        RECT 196.600 66.100 197.000 66.200 ;
        RECT 195.800 65.800 197.000 66.100 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 199.000 65.100 199.400 65.200 ;
        RECT 200.600 65.100 201.000 65.200 ;
        RECT 199.000 64.800 201.000 65.100 ;
        RECT 195.000 61.800 195.400 62.200 ;
        RECT 194.200 53.800 194.600 54.200 ;
        RECT 191.800 51.800 192.200 52.200 ;
        RECT 191.800 46.200 192.100 51.800 ;
        RECT 191.800 45.800 192.200 46.200 ;
        RECT 193.400 43.100 193.800 48.900 ;
        RECT 185.400 36.800 185.800 37.200 ;
        RECT 191.000 36.800 191.400 37.200 ;
        RECT 184.600 30.800 185.000 31.200 ;
        RECT 184.600 29.200 184.900 30.800 ;
        RECT 184.600 28.800 185.000 29.200 ;
        RECT 184.600 26.200 184.900 28.800 ;
        RECT 183.000 25.800 183.400 26.200 ;
        RECT 183.800 25.800 184.200 26.200 ;
        RECT 184.600 25.800 185.000 26.200 ;
        RECT 183.000 22.200 183.300 25.800 ;
        RECT 181.400 21.800 181.800 22.200 ;
        RECT 183.000 21.800 183.400 22.200 ;
        RECT 181.400 19.200 181.700 21.800 ;
        RECT 181.400 18.800 181.800 19.200 ;
        RECT 183.000 17.200 183.300 21.800 ;
        RECT 183.000 16.800 183.400 17.200 ;
        RECT 183.800 15.800 184.200 16.200 ;
        RECT 183.800 15.200 184.100 15.800 ;
        RECT 183.000 14.800 183.400 15.200 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 179.800 13.800 180.200 14.200 ;
        RECT 179.800 12.200 180.100 13.800 ;
        RECT 179.800 11.800 180.200 12.200 ;
        RECT 183.000 9.200 183.300 14.800 ;
        RECT 184.600 13.100 185.000 15.900 ;
        RECT 185.400 14.200 185.700 36.800 ;
        RECT 187.800 35.800 188.200 36.200 ;
        RECT 187.800 35.200 188.100 35.800 ;
        RECT 187.800 34.800 188.200 35.200 ;
        RECT 188.600 34.800 189.000 35.200 ;
        RECT 189.400 34.800 189.800 35.200 ;
        RECT 188.600 34.200 188.900 34.800 ;
        RECT 188.600 33.800 189.000 34.200 ;
        RECT 187.000 32.800 187.400 33.200 ;
        RECT 187.000 32.200 187.300 32.800 ;
        RECT 187.000 31.800 187.400 32.200 ;
        RECT 186.200 21.800 186.600 22.200 ;
        RECT 186.200 19.200 186.500 21.800 ;
        RECT 186.200 18.800 186.600 19.200 ;
        RECT 185.400 13.800 185.800 14.200 ;
        RECT 186.200 12.100 186.600 17.900 ;
        RECT 187.000 15.800 187.400 16.200 ;
        RECT 187.000 15.100 187.300 15.800 ;
        RECT 188.600 15.200 188.900 33.800 ;
        RECT 189.400 28.200 189.700 34.800 ;
        RECT 190.200 33.800 190.600 34.200 ;
        RECT 190.200 33.200 190.500 33.800 ;
        RECT 190.200 32.800 190.600 33.200 ;
        RECT 191.000 31.200 191.300 36.800 ;
        RECT 194.200 35.200 194.500 53.800 ;
        RECT 195.000 53.200 195.300 61.800 ;
        RECT 196.600 60.800 197.000 61.200 ;
        RECT 196.600 55.200 196.900 60.800 ;
        RECT 201.400 57.200 201.700 66.800 ;
        RECT 202.200 66.100 202.600 66.200 ;
        RECT 203.000 66.100 203.400 66.200 ;
        RECT 202.200 65.800 203.400 66.100 ;
        RECT 203.800 59.200 204.100 66.800 ;
        RECT 207.800 66.200 208.100 66.800 ;
        RECT 207.800 65.800 208.200 66.200 ;
        RECT 208.600 65.800 209.000 66.200 ;
        RECT 208.600 65.200 208.900 65.800 ;
        RECT 208.600 64.800 209.000 65.200 ;
        RECT 211.000 65.100 211.300 66.800 ;
        RECT 211.800 66.200 212.100 66.800 ;
        RECT 211.800 65.800 212.200 66.200 ;
        RECT 214.200 66.100 214.600 66.200 ;
        RECT 215.000 66.100 215.400 66.200 ;
        RECT 214.200 65.800 215.400 66.100 ;
        RECT 211.000 64.800 212.100 65.100 ;
        RECT 211.000 63.800 211.400 64.200 ;
        RECT 211.000 63.200 211.300 63.800 ;
        RECT 211.800 63.200 212.100 64.800 ;
        RECT 212.600 64.800 213.000 65.200 ;
        RECT 212.600 64.200 212.900 64.800 ;
        RECT 212.600 63.800 213.000 64.200 ;
        RECT 205.400 62.800 205.800 63.200 ;
        RECT 211.000 62.800 211.400 63.200 ;
        RECT 211.800 62.800 212.200 63.200 ;
        RECT 203.800 58.800 204.200 59.200 ;
        RECT 199.000 56.800 199.400 57.200 ;
        RECT 201.400 56.800 201.800 57.200 ;
        RECT 199.000 56.200 199.300 56.800 ;
        RECT 199.000 55.800 199.400 56.200 ;
        RECT 202.200 55.800 202.600 56.200 ;
        RECT 202.200 55.200 202.500 55.800 ;
        RECT 196.600 54.800 197.000 55.200 ;
        RECT 197.400 54.800 197.800 55.200 ;
        RECT 199.800 54.800 200.200 55.200 ;
        RECT 200.600 55.100 201.000 55.200 ;
        RECT 201.400 55.100 201.800 55.200 ;
        RECT 200.600 54.800 201.800 55.100 ;
        RECT 202.200 54.800 202.600 55.200 ;
        RECT 204.600 54.800 205.000 55.200 ;
        RECT 195.000 52.800 195.400 53.200 ;
        RECT 195.800 52.800 196.200 53.200 ;
        RECT 195.800 52.200 196.100 52.800 ;
        RECT 197.400 52.200 197.700 54.800 ;
        RECT 199.800 52.200 200.100 54.800 ;
        RECT 195.800 51.800 196.200 52.200 ;
        RECT 197.400 51.800 197.800 52.200 ;
        RECT 199.800 51.800 200.200 52.200 ;
        RECT 195.800 49.200 196.100 51.800 ;
        RECT 195.800 48.800 196.200 49.200 ;
        RECT 196.600 45.100 197.000 47.900 ;
        RECT 196.600 43.800 197.000 44.200 ;
        RECT 196.600 39.200 196.900 43.800 ;
        RECT 198.200 43.100 198.600 48.900 ;
        RECT 199.800 47.800 200.200 48.200 ;
        RECT 199.000 46.800 199.400 47.200 ;
        RECT 199.000 42.100 199.300 46.800 ;
        RECT 199.800 46.200 200.100 47.800 ;
        RECT 201.400 47.200 201.700 54.800 ;
        RECT 202.200 51.800 202.600 52.200 ;
        RECT 202.200 48.200 202.500 51.800 ;
        RECT 202.200 47.800 202.600 48.200 ;
        RECT 201.400 46.800 201.800 47.200 ;
        RECT 199.800 45.800 200.200 46.200 ;
        RECT 198.200 41.800 199.300 42.100 ;
        RECT 201.400 44.800 201.800 45.200 ;
        RECT 196.600 38.800 197.000 39.200 ;
        RECT 194.200 34.800 194.600 35.200 ;
        RECT 195.000 34.800 195.400 35.200 ;
        RECT 196.600 35.100 197.000 35.200 ;
        RECT 197.400 35.100 197.800 35.200 ;
        RECT 196.600 34.800 197.800 35.100 ;
        RECT 195.000 34.200 195.300 34.800 ;
        RECT 193.400 33.800 193.800 34.200 ;
        RECT 195.000 33.800 195.400 34.200 ;
        RECT 193.400 33.200 193.700 33.800 ;
        RECT 193.400 32.800 193.800 33.200 ;
        RECT 191.000 30.800 191.400 31.200 ;
        RECT 195.000 29.200 195.300 33.800 ;
        RECT 190.200 29.100 190.600 29.200 ;
        RECT 191.000 29.100 191.400 29.200 ;
        RECT 190.200 28.800 191.400 29.100 ;
        RECT 189.400 27.800 189.800 28.200 ;
        RECT 187.000 14.700 187.400 15.100 ;
        RECT 188.600 14.800 189.000 15.200 ;
        RECT 189.400 9.200 189.700 27.800 ;
        RECT 192.600 23.100 193.000 28.900 ;
        RECT 195.000 28.800 195.400 29.200 ;
        RECT 195.800 28.800 196.200 29.200 ;
        RECT 195.800 26.200 196.100 28.800 ;
        RECT 196.600 26.800 197.000 27.200 ;
        RECT 195.800 25.800 196.200 26.200 ;
        RECT 196.600 24.200 196.900 26.800 ;
        RECT 196.600 23.800 197.000 24.200 ;
        RECT 197.400 23.100 197.800 28.900 ;
        RECT 198.200 19.200 198.500 41.800 ;
        RECT 201.400 39.200 201.700 44.800 ;
        RECT 203.000 43.100 203.400 48.900 ;
        RECT 204.600 44.200 204.900 54.800 ;
        RECT 205.400 54.200 205.700 62.800 ;
        RECT 206.200 57.800 206.600 58.200 ;
        RECT 206.200 55.200 206.500 57.800 ;
        RECT 208.600 56.100 209.000 56.200 ;
        RECT 209.400 56.100 209.800 56.200 ;
        RECT 208.600 55.800 209.800 56.100 ;
        RECT 206.200 54.800 206.600 55.200 ;
        RECT 209.400 55.100 209.800 55.200 ;
        RECT 210.200 55.100 210.600 55.200 ;
        RECT 209.400 54.800 210.600 55.100 ;
        RECT 205.400 53.800 205.800 54.200 ;
        RECT 206.200 49.200 206.500 54.800 ;
        RECT 211.000 53.100 211.400 55.900 ;
        RECT 211.800 53.800 212.200 54.200 ;
        RECT 211.800 53.200 212.100 53.800 ;
        RECT 211.800 52.800 212.200 53.200 ;
        RECT 212.600 52.100 213.000 57.900 ;
        RECT 213.400 55.000 213.800 55.100 ;
        RECT 214.200 55.000 214.600 55.100 ;
        RECT 213.400 54.700 214.600 55.000 ;
        RECT 215.800 49.200 216.100 66.800 ;
        RECT 219.000 65.800 219.400 66.200 ;
        RECT 219.000 65.200 219.300 65.800 ;
        RECT 219.000 64.800 219.400 65.200 ;
        RECT 217.400 52.100 217.800 57.900 ;
        RECT 218.200 55.800 218.600 56.200 ;
        RECT 218.200 49.200 218.500 55.800 ;
        RECT 219.800 53.100 220.100 68.800 ;
        RECT 220.600 55.200 220.900 71.800 ;
        RECT 223.800 70.800 224.200 71.200 ;
        RECT 223.800 66.200 224.100 70.800 ;
        RECT 227.800 69.200 228.100 74.800 ;
        RECT 229.400 71.800 229.800 72.200 ;
        RECT 229.400 71.200 229.700 71.800 ;
        RECT 229.400 70.800 229.800 71.200 ;
        RECT 227.800 68.800 228.200 69.200 ;
        RECT 224.600 67.800 225.000 68.200 ;
        RECT 225.400 67.800 225.800 68.200 ;
        RECT 224.600 66.200 224.900 67.800 ;
        RECT 225.400 67.200 225.700 67.800 ;
        RECT 225.400 66.800 225.800 67.200 ;
        RECT 222.200 65.800 222.600 66.200 ;
        RECT 223.800 65.800 224.200 66.200 ;
        RECT 224.600 65.800 225.000 66.200 ;
        RECT 227.800 65.800 228.200 66.200 ;
        RECT 222.200 59.200 222.500 65.800 ;
        RECT 227.000 62.800 227.400 63.200 ;
        RECT 227.000 59.200 227.300 62.800 ;
        RECT 222.200 58.800 222.600 59.200 ;
        RECT 225.400 58.800 225.800 59.200 ;
        RECT 227.000 58.800 227.400 59.200 ;
        RECT 225.400 55.200 225.700 58.800 ;
        RECT 227.000 56.800 227.400 57.200 ;
        RECT 220.600 54.800 221.000 55.200 ;
        RECT 223.000 54.800 223.400 55.200 ;
        RECT 223.800 54.800 224.200 55.200 ;
        RECT 224.600 54.800 225.000 55.200 ;
        RECT 225.400 54.800 225.800 55.200 ;
        RECT 226.200 54.800 226.600 55.200 ;
        RECT 219.800 52.800 220.900 53.100 ;
        RECT 219.800 51.800 220.200 52.200 ;
        RECT 206.200 48.800 206.600 49.200 ;
        RECT 215.800 48.800 216.200 49.200 ;
        RECT 217.400 48.800 217.800 49.200 ;
        RECT 218.200 48.800 218.600 49.200 ;
        RECT 211.000 48.100 211.400 48.200 ;
        RECT 211.800 48.100 212.200 48.200 ;
        RECT 211.000 47.800 212.200 48.100 ;
        RECT 211.800 46.800 212.200 47.200 ;
        RECT 213.400 46.800 213.800 47.200 ;
        RECT 211.800 46.200 212.100 46.800 ;
        RECT 213.400 46.200 213.700 46.800 ;
        RECT 217.400 46.200 217.700 48.800 ;
        RECT 219.800 47.200 220.100 51.800 ;
        RECT 219.800 46.800 220.200 47.200 ;
        RECT 220.600 46.200 220.900 52.800 ;
        RECT 223.000 49.200 223.300 54.800 ;
        RECT 223.800 49.200 224.100 54.800 ;
        RECT 224.600 54.200 224.900 54.800 ;
        RECT 224.600 53.800 225.000 54.200 ;
        RECT 223.000 48.800 223.400 49.200 ;
        RECT 223.800 48.800 224.200 49.200 ;
        RECT 225.400 46.200 225.700 54.800 ;
        RECT 226.200 54.200 226.500 54.800 ;
        RECT 226.200 53.800 226.600 54.200 ;
        RECT 227.000 49.200 227.300 56.800 ;
        RECT 227.000 48.800 227.400 49.200 ;
        RECT 207.000 46.100 207.400 46.200 ;
        RECT 207.800 46.100 208.200 46.200 ;
        RECT 207.000 45.800 208.200 46.100 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 212.600 45.800 213.000 46.200 ;
        RECT 213.400 45.800 213.800 46.200 ;
        RECT 214.200 45.800 214.600 46.200 ;
        RECT 216.600 45.800 217.000 46.200 ;
        RECT 217.400 45.800 217.800 46.200 ;
        RECT 220.600 45.800 221.000 46.200 ;
        RECT 221.400 45.800 221.800 46.200 ;
        RECT 223.800 45.800 224.200 46.200 ;
        RECT 225.400 45.800 225.800 46.200 ;
        RECT 226.200 45.800 226.600 46.200 ;
        RECT 204.600 43.800 205.000 44.200 ;
        RECT 204.600 41.800 205.000 42.200 ;
        RECT 203.800 40.800 204.200 41.200 ;
        RECT 201.400 38.800 201.800 39.200 ;
        RECT 203.000 35.800 203.400 36.200 ;
        RECT 203.000 35.200 203.300 35.800 ;
        RECT 203.800 35.200 204.100 40.800 ;
        RECT 204.600 36.200 204.900 41.800 ;
        RECT 212.600 41.200 212.900 45.800 ;
        RECT 214.200 45.100 214.500 45.800 ;
        RECT 213.400 44.800 214.500 45.100 ;
        RECT 216.600 45.200 216.900 45.800 ;
        RECT 216.600 44.800 217.000 45.200 ;
        RECT 212.600 40.800 213.000 41.200 ;
        RECT 213.400 39.200 213.700 44.800 ;
        RECT 217.400 40.200 217.700 45.800 ;
        RECT 221.400 45.200 221.700 45.800 ;
        RECT 221.400 44.800 221.800 45.200 ;
        RECT 218.200 43.800 218.600 44.200 ;
        RECT 217.400 39.800 217.800 40.200 ;
        RECT 218.200 39.200 218.500 43.800 ;
        RECT 211.800 38.800 212.200 39.200 ;
        RECT 213.400 38.800 213.800 39.200 ;
        RECT 218.200 38.800 218.600 39.200 ;
        RECT 204.600 35.800 205.000 36.200 ;
        RECT 207.000 35.800 207.400 36.200 ;
        RECT 199.000 34.800 199.400 35.200 ;
        RECT 202.200 34.800 202.600 35.200 ;
        RECT 203.000 34.800 203.400 35.200 ;
        RECT 203.800 34.800 204.200 35.200 ;
        RECT 199.000 33.200 199.300 34.800 ;
        RECT 202.200 33.200 202.500 34.800 ;
        RECT 199.000 32.800 199.400 33.200 ;
        RECT 202.200 32.800 202.600 33.200 ;
        RECT 203.800 31.200 204.100 34.800 ;
        RECT 204.600 34.200 204.900 35.800 ;
        RECT 207.000 35.200 207.300 35.800 ;
        RECT 211.800 35.200 212.100 38.800 ;
        RECT 215.000 37.800 215.400 38.200 ;
        RECT 215.000 35.200 215.300 37.800 ;
        RECT 219.800 35.800 220.200 36.200 ;
        RECT 219.800 35.200 220.100 35.800 ;
        RECT 207.000 34.800 207.400 35.200 ;
        RECT 211.800 34.800 212.200 35.200 ;
        RECT 214.200 34.800 214.600 35.200 ;
        RECT 215.000 34.800 215.400 35.200 ;
        RECT 215.800 34.800 216.200 35.200 ;
        RECT 219.000 34.800 219.400 35.200 ;
        RECT 219.800 34.800 220.200 35.200 ;
        RECT 220.600 34.800 221.000 35.200 ;
        RECT 207.000 34.200 207.300 34.800 ;
        RECT 204.600 33.800 205.000 34.200 ;
        RECT 207.000 33.800 207.400 34.200 ;
        RECT 207.000 32.800 207.400 33.200 ;
        RECT 209.400 33.100 209.800 33.200 ;
        RECT 210.200 33.100 210.600 33.200 ;
        RECT 209.400 32.800 210.600 33.100 ;
        RECT 205.400 31.800 205.800 32.200 ;
        RECT 201.400 30.800 201.800 31.200 ;
        RECT 203.800 30.800 204.200 31.200 ;
        RECT 199.000 25.100 199.400 27.900 ;
        RECT 199.800 27.100 200.200 27.200 ;
        RECT 200.600 27.100 201.000 27.200 ;
        RECT 199.800 26.800 201.000 27.100 ;
        RECT 195.800 18.800 196.200 19.200 ;
        RECT 198.200 18.800 198.600 19.200 ;
        RECT 191.000 12.100 191.400 17.900 ;
        RECT 194.200 14.800 194.600 15.200 ;
        RECT 194.200 13.200 194.500 14.800 ;
        RECT 194.200 12.800 194.600 13.200 ;
        RECT 192.600 12.100 193.000 12.200 ;
        RECT 193.400 12.100 193.800 12.200 ;
        RECT 192.600 11.800 193.800 12.100 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 168.600 7.800 169.000 8.200 ;
        RECT 171.000 7.800 171.400 8.200 ;
        RECT 177.400 7.800 177.800 8.200 ;
        RECT 179.000 7.800 179.400 8.200 ;
        RECT 168.600 7.200 168.900 7.800 ;
        RECT 168.600 6.800 169.000 7.200 ;
        RECT 171.000 6.200 171.300 7.800 ;
        RECT 171.800 6.800 172.200 7.200 ;
        RECT 171.800 6.200 172.100 6.800 ;
        RECT 177.400 6.200 177.700 7.800 ;
        RECT 180.600 6.800 181.000 7.200 ;
        RECT 180.600 6.200 180.900 6.800 ;
        RECT 171.000 5.800 171.400 6.200 ;
        RECT 171.800 5.800 172.200 6.200 ;
        RECT 172.600 6.100 173.000 6.200 ;
        RECT 173.400 6.100 173.800 6.200 ;
        RECT 172.600 5.800 173.800 6.100 ;
        RECT 175.800 6.100 176.200 6.200 ;
        RECT 176.600 6.100 177.000 6.200 ;
        RECT 175.800 5.800 177.000 6.100 ;
        RECT 177.400 5.800 177.800 6.200 ;
        RECT 180.600 5.800 181.000 6.200 ;
        RECT 185.400 3.100 185.800 8.900 ;
        RECT 189.400 8.800 189.800 9.200 ;
        RECT 187.800 6.100 188.200 6.200 ;
        RECT 188.600 6.100 189.000 6.200 ;
        RECT 187.800 5.800 189.000 6.100 ;
        RECT 190.200 3.100 190.600 8.900 ;
        RECT 191.000 7.800 191.400 8.200 ;
        RECT 191.000 7.200 191.300 7.800 ;
        RECT 191.000 6.800 191.400 7.200 ;
        RECT 191.800 5.100 192.200 7.900 ;
        RECT 192.600 5.100 193.000 7.900 ;
        RECT 194.200 3.100 194.600 8.900 ;
        RECT 195.800 6.200 196.100 18.800 ;
        RECT 196.600 14.800 197.000 15.200 ;
        RECT 196.600 14.200 196.900 14.800 ;
        RECT 199.800 14.200 200.100 26.800 ;
        RECT 200.600 26.100 201.000 26.200 ;
        RECT 201.400 26.100 201.700 30.800 ;
        RECT 205.400 29.200 205.700 31.800 ;
        RECT 202.200 29.100 202.600 29.200 ;
        RECT 203.000 29.100 203.400 29.200 ;
        RECT 202.200 28.800 203.400 29.100 ;
        RECT 205.400 28.800 205.800 29.200 ;
        RECT 205.400 27.800 205.800 28.200 ;
        RECT 205.400 27.200 205.700 27.800 ;
        RECT 200.600 25.800 201.700 26.100 ;
        RECT 203.000 26.800 203.400 27.200 ;
        RECT 205.400 26.800 205.800 27.200 ;
        RECT 203.000 25.200 203.300 26.800 ;
        RECT 203.800 26.100 204.200 26.200 ;
        RECT 204.600 26.100 205.000 26.200 ;
        RECT 203.800 25.800 205.000 26.100 ;
        RECT 203.000 24.800 203.400 25.200 ;
        RECT 204.600 15.200 204.900 25.800 ;
        RECT 204.600 14.800 205.000 15.200 ;
        RECT 196.600 13.800 197.000 14.200 ;
        RECT 199.800 13.800 200.200 14.200 ;
        RECT 203.800 13.800 204.200 14.200 ;
        RECT 204.600 14.100 205.000 14.200 ;
        RECT 205.400 14.100 205.700 26.800 ;
        RECT 207.000 17.200 207.300 32.800 ;
        RECT 214.200 32.200 214.500 34.800 ;
        RECT 215.800 33.200 216.100 34.800 ;
        RECT 219.000 33.200 219.300 34.800 ;
        RECT 215.800 33.100 216.200 33.200 ;
        RECT 215.800 32.800 216.900 33.100 ;
        RECT 219.000 32.800 219.400 33.200 ;
        RECT 214.200 31.800 214.600 32.200 ;
        RECT 216.600 29.200 216.900 32.800 ;
        RECT 219.000 29.800 219.400 30.200 ;
        RECT 219.000 29.200 219.300 29.800 ;
        RECT 220.600 29.200 220.900 34.800 ;
        RECT 221.400 34.100 221.800 34.200 ;
        RECT 222.200 34.100 222.600 34.200 ;
        RECT 221.400 33.800 222.600 34.100 ;
        RECT 223.800 33.200 224.100 45.800 ;
        RECT 226.200 44.200 226.500 45.800 ;
        RECT 226.200 43.800 226.600 44.200 ;
        RECT 225.400 41.800 225.800 42.200 ;
        RECT 225.400 35.200 225.700 41.800 ;
        RECT 227.800 39.200 228.100 65.800 ;
        RECT 228.600 65.100 229.000 67.900 ;
        RECT 229.400 66.800 229.800 67.200 ;
        RECT 229.400 55.200 229.700 66.800 ;
        RECT 230.200 63.100 230.600 68.900 ;
        RECT 231.000 68.200 231.300 81.800 ;
        RECT 232.600 78.100 233.000 78.200 ;
        RECT 233.400 78.100 233.800 78.200 ;
        RECT 232.600 77.800 233.800 78.100 ;
        RECT 231.800 77.100 232.200 77.200 ;
        RECT 232.600 77.100 233.000 77.200 ;
        RECT 231.800 76.800 233.000 77.100 ;
        RECT 231.800 75.800 232.200 76.200 ;
        RECT 231.800 75.200 232.100 75.800 ;
        RECT 231.800 74.800 232.200 75.200 ;
        RECT 232.600 74.800 233.000 75.200 ;
        RECT 232.600 74.200 232.900 74.800 ;
        RECT 232.600 73.800 233.000 74.200 ;
        RECT 231.800 70.800 232.200 71.200 ;
        RECT 231.000 67.800 231.400 68.200 ;
        RECT 231.800 66.200 232.100 70.800 ;
        RECT 231.800 65.800 232.200 66.200 ;
        RECT 232.600 62.200 232.900 73.800 ;
        RECT 234.200 68.200 234.500 82.800 ;
        RECT 238.200 79.200 238.500 83.800 ;
        RECT 238.200 78.800 238.600 79.200 ;
        RECT 235.800 72.100 236.200 77.900 ;
        RECT 238.200 76.800 238.600 77.200 ;
        RECT 238.200 75.200 238.500 76.800 ;
        RECT 238.200 74.800 238.600 75.200 ;
        RECT 240.600 72.100 241.000 77.900 ;
        RECT 241.400 74.200 241.700 84.800 ;
        RECT 243.000 80.200 243.300 94.800 ;
        RECT 245.400 93.200 245.700 111.800 ;
        RECT 247.000 109.200 247.300 122.800 ;
        RECT 248.600 121.200 248.900 141.800 ;
        RECT 249.400 127.200 249.700 143.800 ;
        RECT 250.200 134.700 250.600 135.100 ;
        RECT 250.200 134.200 250.500 134.700 ;
        RECT 250.200 133.800 250.600 134.200 ;
        RECT 251.000 132.100 251.400 137.900 ;
        RECT 251.800 134.200 252.100 143.800 ;
        RECT 252.600 143.100 253.000 148.900 ;
        RECT 255.800 146.800 256.200 147.200 ;
        RECT 255.800 146.200 256.100 146.800 ;
        RECT 255.800 145.800 256.200 146.200 ;
        RECT 254.200 138.800 254.600 139.200 ;
        RECT 251.800 133.800 252.200 134.200 ;
        RECT 252.600 133.100 253.000 135.900 ;
        RECT 254.200 134.200 254.500 138.800 ;
        RECT 256.600 137.200 256.900 161.800 ;
        RECT 258.200 152.100 258.600 157.900 ;
        RECT 259.000 155.800 259.400 156.200 ;
        RECT 259.000 155.200 259.300 155.800 ;
        RECT 259.000 154.800 259.400 155.200 ;
        RECT 259.800 154.800 260.200 155.200 ;
        RECT 259.000 149.100 259.300 154.800 ;
        RECT 259.800 154.200 260.100 154.800 ;
        RECT 259.800 153.800 260.200 154.200 ;
        RECT 257.400 143.100 257.800 148.900 ;
        RECT 258.200 148.800 259.300 149.100 ;
        RECT 258.200 147.200 258.500 148.800 ;
        RECT 258.200 146.800 258.600 147.200 ;
        RECT 259.000 145.100 259.400 147.900 ;
        RECT 260.600 143.200 260.900 165.800 ;
        RECT 262.200 165.800 262.600 166.200 ;
        RECT 262.200 162.200 262.500 165.800 ;
        RECT 262.200 161.800 262.600 162.200 ;
        RECT 263.000 152.100 263.400 157.900 ;
        RECT 264.600 153.100 265.000 155.900 ;
        RECT 260.600 142.800 261.000 143.200 ;
        RECT 260.600 141.800 261.000 142.200 ;
        RECT 260.600 141.200 260.900 141.800 ;
        RECT 260.600 140.800 261.000 141.200 ;
        RECT 256.600 136.800 257.000 137.200 ;
        RECT 257.400 135.800 257.800 136.200 ;
        RECT 257.400 135.200 257.700 135.800 ;
        RECT 255.000 134.800 255.400 135.200 ;
        RECT 257.400 134.800 257.800 135.200 ;
        RECT 261.400 134.800 261.800 135.200 ;
        RECT 255.000 134.200 255.300 134.800 ;
        RECT 254.200 133.800 254.600 134.200 ;
        RECT 255.000 133.800 255.400 134.200 ;
        RECT 255.800 133.800 256.200 134.200 ;
        RECT 259.000 134.100 259.400 134.200 ;
        RECT 259.800 134.100 260.200 134.200 ;
        RECT 259.000 133.800 260.200 134.100 ;
        RECT 255.800 133.200 256.100 133.800 ;
        RECT 255.800 132.800 256.200 133.200 ;
        RECT 261.400 130.100 261.700 134.800 ;
        RECT 260.600 129.800 261.700 130.100 ;
        RECT 250.200 128.800 250.600 129.200 ;
        RECT 250.200 128.200 250.500 128.800 ;
        RECT 250.200 127.800 250.600 128.200 ;
        RECT 249.400 126.800 249.800 127.200 ;
        RECT 248.600 120.800 249.000 121.200 ;
        RECT 249.400 119.200 249.700 126.800 ;
        RECT 252.600 123.100 253.000 128.900 ;
        RECT 254.200 125.800 254.600 126.200 ;
        RECT 255.000 126.100 255.400 126.200 ;
        RECT 255.800 126.100 256.200 126.200 ;
        RECT 255.000 125.800 256.200 126.100 ;
        RECT 249.400 118.800 249.800 119.200 ;
        RECT 248.600 112.100 249.000 117.900 ;
        RECT 251.800 115.800 252.200 116.200 ;
        RECT 251.800 115.200 252.100 115.800 ;
        RECT 251.800 114.800 252.200 115.200 ;
        RECT 253.400 112.100 253.800 117.900 ;
        RECT 254.200 114.200 254.500 125.800 ;
        RECT 257.400 123.100 257.800 128.900 ;
        RECT 259.000 125.100 259.400 127.900 ;
        RECT 259.800 126.800 260.200 127.200 ;
        RECT 259.800 126.200 260.100 126.800 ;
        RECT 259.800 125.800 260.200 126.200 ;
        RECT 256.600 116.800 257.000 117.200 ;
        RECT 254.200 113.800 254.600 114.200 ;
        RECT 254.200 113.200 254.500 113.800 ;
        RECT 254.200 112.800 254.600 113.200 ;
        RECT 255.000 113.100 255.400 115.900 ;
        RECT 255.800 113.100 256.200 115.900 ;
        RECT 256.600 114.200 256.900 116.800 ;
        RECT 256.600 113.800 257.000 114.200 ;
        RECT 257.400 112.100 257.800 117.900 ;
        RECT 258.200 115.000 258.600 115.100 ;
        RECT 259.000 115.000 259.400 115.100 ;
        RECT 258.200 114.700 259.400 115.000 ;
        RECT 246.200 109.100 246.600 109.200 ;
        RECT 247.000 109.100 247.400 109.200 ;
        RECT 246.200 108.800 247.400 109.100 ;
        RECT 253.400 108.800 253.800 109.200 ;
        RECT 251.000 107.100 251.400 107.200 ;
        RECT 251.800 107.100 252.200 107.200 ;
        RECT 251.000 106.800 252.200 107.100 ;
        RECT 252.600 105.100 253.000 107.900 ;
        RECT 253.400 107.200 253.700 108.800 ;
        RECT 253.400 106.800 253.800 107.200 ;
        RECT 254.200 103.100 254.600 108.900 ;
        RECT 255.800 105.800 256.200 106.200 ;
        RECT 246.200 94.700 246.600 95.100 ;
        RECT 246.200 93.200 246.500 94.700 ;
        RECT 245.400 92.800 245.800 93.200 ;
        RECT 246.200 92.800 246.600 93.200 ;
        RECT 247.000 92.100 247.400 97.900 ;
        RECT 255.000 96.800 255.400 97.200 ;
        RECT 250.200 96.100 250.600 96.200 ;
        RECT 251.000 96.100 251.400 96.200 ;
        RECT 248.600 93.100 249.000 95.900 ;
        RECT 250.200 95.800 251.400 96.100 ;
        RECT 249.400 93.800 249.800 94.200 ;
        RECT 247.000 86.800 247.400 87.200 ;
        RECT 247.000 85.200 247.300 86.800 ;
        RECT 247.000 84.800 247.400 85.200 ;
        RECT 243.000 79.800 243.400 80.200 ;
        RECT 241.400 73.800 241.800 74.200 ;
        RECT 242.200 73.100 242.600 75.900 ;
        RECT 243.000 75.100 243.400 75.200 ;
        RECT 243.800 75.100 244.200 75.200 ;
        RECT 243.000 74.800 244.200 75.100 ;
        RECT 245.400 74.800 245.800 75.200 ;
        RECT 243.000 69.200 243.300 74.800 ;
        RECT 245.400 74.200 245.700 74.800 ;
        RECT 243.800 73.800 244.200 74.200 ;
        RECT 245.400 73.800 245.800 74.200 ;
        RECT 243.800 73.200 244.100 73.800 ;
        RECT 243.800 72.800 244.200 73.200 ;
        RECT 245.400 73.100 245.800 73.200 ;
        RECT 246.200 73.100 246.600 73.200 ;
        RECT 245.400 72.800 246.600 73.100 ;
        RECT 246.200 72.100 246.600 72.200 ;
        RECT 247.000 72.100 247.400 72.200 ;
        RECT 248.600 72.100 249.000 77.900 ;
        RECT 249.400 76.200 249.700 93.800 ;
        RECT 250.200 76.200 250.500 95.800 ;
        RECT 255.000 95.200 255.300 96.800 ;
        RECT 251.000 94.800 251.400 95.200 ;
        RECT 255.000 94.800 255.400 95.200 ;
        RECT 251.000 94.200 251.300 94.800 ;
        RECT 251.000 93.800 251.400 94.200 ;
        RECT 253.400 92.800 253.800 93.200 ;
        RECT 254.200 93.100 254.600 93.200 ;
        RECT 255.000 93.100 255.400 93.200 ;
        RECT 254.200 92.800 255.400 93.100 ;
        RECT 253.400 92.200 253.700 92.800 ;
        RECT 251.000 91.800 251.400 92.200 ;
        RECT 253.400 91.800 253.800 92.200 ;
        RECT 249.400 75.800 249.800 76.200 ;
        RECT 250.200 75.800 250.600 76.200 ;
        RECT 249.400 75.100 249.800 75.200 ;
        RECT 250.200 75.100 250.600 75.200 ;
        RECT 249.400 74.800 250.600 75.100 ;
        RECT 246.200 71.800 247.400 72.100 ;
        RECT 249.400 71.800 249.800 72.200 ;
        RECT 234.200 67.800 234.600 68.200 ;
        RECT 233.400 65.800 233.800 66.200 ;
        RECT 232.600 61.800 233.000 62.200 ;
        RECT 230.200 55.800 230.600 56.200 ;
        RECT 228.600 54.800 229.000 55.200 ;
        RECT 229.400 54.800 229.800 55.200 ;
        RECT 228.600 54.200 228.900 54.800 ;
        RECT 228.600 53.800 229.000 54.200 ;
        RECT 230.200 47.200 230.500 55.800 ;
        RECT 231.000 54.800 231.400 55.200 ;
        RECT 231.000 52.200 231.300 54.800 ;
        RECT 231.800 53.800 232.200 54.200 ;
        RECT 231.800 53.200 232.100 53.800 ;
        RECT 233.400 53.200 233.700 65.800 ;
        RECT 235.000 63.100 235.400 68.900 ;
        RECT 243.000 68.800 243.400 69.200 ;
        RECT 238.200 67.800 238.600 68.200 ;
        RECT 244.600 68.100 245.000 68.200 ;
        RECT 245.400 68.100 245.800 68.200 ;
        RECT 244.600 67.800 245.800 68.100 ;
        RECT 238.200 67.200 238.500 67.800 ;
        RECT 238.200 66.800 238.600 67.200 ;
        RECT 247.800 66.800 248.200 67.200 ;
        RECT 248.600 66.800 249.000 67.200 ;
        RECT 247.800 66.200 248.100 66.800 ;
        RECT 248.600 66.200 248.900 66.800 ;
        RECT 241.400 65.800 241.800 66.200 ;
        RECT 242.200 65.800 242.600 66.200 ;
        RECT 243.000 65.800 243.400 66.200 ;
        RECT 243.800 65.800 244.200 66.200 ;
        RECT 246.200 65.800 246.600 66.200 ;
        RECT 247.800 65.800 248.200 66.200 ;
        RECT 248.600 65.800 249.000 66.200 ;
        RECT 235.800 59.800 236.200 60.200 ;
        RECT 234.200 55.800 234.600 56.200 ;
        RECT 234.200 54.200 234.500 55.800 ;
        RECT 235.800 55.200 236.100 59.800 ;
        RECT 236.600 55.800 237.000 56.200 ;
        RECT 237.400 55.800 237.800 56.200 ;
        RECT 236.600 55.200 236.900 55.800 ;
        RECT 235.000 54.800 235.400 55.200 ;
        RECT 235.800 54.800 236.200 55.200 ;
        RECT 236.600 54.800 237.000 55.200 ;
        RECT 234.200 53.800 234.600 54.200 ;
        RECT 231.800 52.800 232.200 53.200 ;
        RECT 233.400 52.800 233.800 53.200 ;
        RECT 235.000 52.200 235.300 54.800 ;
        RECT 231.000 51.800 231.400 52.200 ;
        RECT 235.000 51.800 235.400 52.200 ;
        RECT 235.800 52.100 236.100 54.800 ;
        RECT 235.800 51.800 236.900 52.100 ;
        RECT 235.000 51.100 235.300 51.800 ;
        RECT 235.000 50.800 236.100 51.100 ;
        RECT 235.000 48.800 235.400 49.200 ;
        RECT 235.000 47.200 235.300 48.800 ;
        RECT 235.800 47.200 236.100 50.800 ;
        RECT 230.200 46.800 230.600 47.200 ;
        RECT 231.000 46.800 231.400 47.200 ;
        RECT 232.600 47.100 233.000 47.200 ;
        RECT 233.400 47.100 233.800 47.200 ;
        RECT 232.600 46.800 233.800 47.100 ;
        RECT 235.000 46.800 235.400 47.200 ;
        RECT 235.800 46.800 236.200 47.200 ;
        RECT 231.000 46.200 231.300 46.800 ;
        RECT 228.600 45.800 229.000 46.200 ;
        RECT 231.000 45.800 231.400 46.200 ;
        RECT 233.400 45.800 233.800 46.200 ;
        RECT 228.600 43.200 228.900 45.800 ;
        RECT 233.400 45.200 233.700 45.800 ;
        RECT 233.400 44.800 233.800 45.200 ;
        RECT 236.600 45.100 236.900 51.800 ;
        RECT 237.400 49.200 237.700 55.800 ;
        RECT 238.200 53.100 238.600 55.900 ;
        RECT 239.000 53.800 239.400 54.200 ;
        RECT 239.000 53.200 239.300 53.800 ;
        RECT 239.000 52.800 239.400 53.200 ;
        RECT 239.800 52.100 240.200 57.900 ;
        RECT 240.600 55.800 241.000 56.200 ;
        RECT 240.600 55.100 240.900 55.800 ;
        RECT 240.600 54.700 241.000 55.100 ;
        RECT 241.400 51.200 241.700 65.800 ;
        RECT 242.200 65.200 242.500 65.800 ;
        RECT 242.200 64.800 242.600 65.200 ;
        RECT 242.200 57.200 242.500 64.800 ;
        RECT 243.000 59.200 243.300 65.800 ;
        RECT 243.800 65.200 244.100 65.800 ;
        RECT 243.800 64.800 244.200 65.200 ;
        RECT 246.200 63.200 246.500 65.800 ;
        RECT 246.200 62.800 246.600 63.200 ;
        RECT 249.400 62.200 249.700 71.800 ;
        RECT 251.000 68.200 251.300 91.800 ;
        RECT 251.800 90.800 252.200 91.200 ;
        RECT 251.000 67.800 251.400 68.200 ;
        RECT 250.200 65.800 250.600 66.200 ;
        RECT 251.000 65.800 251.400 66.200 ;
        RECT 250.200 65.200 250.500 65.800 ;
        RECT 250.200 64.800 250.600 65.200 ;
        RECT 251.000 62.200 251.300 65.800 ;
        RECT 249.400 61.800 249.800 62.200 ;
        RECT 251.000 61.800 251.400 62.200 ;
        RECT 243.000 58.800 243.400 59.200 ;
        RECT 242.200 56.800 242.600 57.200 ;
        RECT 244.600 52.100 245.000 57.900 ;
        RECT 247.800 55.100 248.200 55.200 ;
        RECT 248.600 55.100 249.000 55.200 ;
        RECT 247.800 54.800 249.000 55.100 ;
        RECT 247.800 53.800 248.200 54.200 ;
        RECT 248.600 53.800 249.000 54.200 ;
        RECT 246.200 52.100 246.600 52.200 ;
        RECT 247.000 52.100 247.400 52.200 ;
        RECT 246.200 51.800 247.400 52.100 ;
        RECT 241.400 50.800 241.800 51.200 ;
        RECT 247.800 49.200 248.100 53.800 ;
        RECT 248.600 49.200 248.900 53.800 ;
        RECT 237.400 48.800 237.800 49.200 ;
        RECT 238.200 48.800 238.600 49.200 ;
        RECT 238.200 48.200 238.500 48.800 ;
        RECT 238.200 47.800 238.600 48.200 ;
        RECT 237.400 45.100 237.800 45.200 ;
        RECT 236.600 44.800 237.800 45.100 ;
        RECT 230.200 43.800 230.600 44.200 ;
        RECT 228.600 42.800 229.000 43.200 ;
        RECT 227.800 38.800 228.200 39.200 ;
        RECT 226.200 35.800 226.600 36.200 ;
        RECT 226.200 35.200 226.500 35.800 ;
        RECT 225.400 34.800 225.800 35.200 ;
        RECT 226.200 34.800 226.600 35.200 ;
        RECT 227.000 34.800 227.400 35.200 ;
        RECT 225.400 34.200 225.700 34.800 ;
        RECT 225.400 33.800 225.800 34.200 ;
        RECT 223.800 32.800 224.200 33.200 ;
        RECT 222.200 31.800 222.600 32.200 ;
        RECT 222.200 30.200 222.500 31.800 ;
        RECT 222.200 29.800 222.600 30.200 ;
        RECT 223.800 29.200 224.100 32.800 ;
        RECT 226.200 29.800 226.600 30.200 ;
        RECT 207.800 25.100 208.200 27.900 ;
        RECT 209.400 23.100 209.800 28.900 ;
        RECT 210.200 28.800 210.600 29.200 ;
        RECT 210.200 26.300 210.500 28.800 ;
        RECT 213.400 27.800 213.800 28.200 ;
        RECT 210.200 25.900 210.600 26.300 ;
        RECT 213.400 26.200 213.700 27.800 ;
        RECT 213.400 25.800 213.800 26.200 ;
        RECT 214.200 23.100 214.600 28.900 ;
        RECT 216.600 28.800 217.000 29.200 ;
        RECT 219.000 28.800 219.400 29.200 ;
        RECT 220.600 28.800 221.000 29.200 ;
        RECT 222.200 29.100 222.600 29.200 ;
        RECT 223.000 29.100 223.400 29.200 ;
        RECT 222.200 28.800 223.400 29.100 ;
        RECT 223.800 28.800 224.200 29.200 ;
        RECT 218.200 26.800 218.600 27.200 ;
        RECT 218.200 26.200 218.500 26.800 ;
        RECT 216.600 26.100 217.000 26.200 ;
        RECT 217.400 26.100 217.800 26.200 ;
        RECT 216.600 25.800 217.800 26.100 ;
        RECT 218.200 25.800 218.600 26.200 ;
        RECT 220.600 25.800 221.000 26.200 ;
        RECT 207.000 17.100 207.400 17.200 ;
        RECT 208.600 17.100 209.000 17.200 ;
        RECT 207.000 16.800 209.000 17.100 ;
        RECT 211.800 17.100 212.200 17.200 ;
        RECT 212.600 17.100 213.000 17.200 ;
        RECT 211.800 16.800 213.000 17.100 ;
        RECT 211.000 16.100 211.400 16.200 ;
        RECT 211.800 16.100 212.200 16.200 ;
        RECT 211.000 15.800 212.200 16.100 ;
        RECT 210.200 15.100 210.600 15.200 ;
        RECT 211.000 15.100 211.400 15.200 ;
        RECT 210.200 14.800 211.400 15.100 ;
        RECT 213.400 14.800 213.800 15.200 ;
        RECT 204.600 13.800 205.700 14.100 ;
        RECT 211.000 14.100 211.400 14.200 ;
        RECT 211.800 14.100 212.200 14.200 ;
        RECT 211.000 13.800 212.200 14.100 ;
        RECT 203.800 13.100 204.100 13.800 ;
        RECT 203.800 12.800 204.900 13.100 ;
        RECT 198.200 11.800 198.600 12.200 ;
        RECT 198.200 7.200 198.500 11.800 ;
        RECT 204.600 9.200 204.900 12.800 ;
        RECT 206.200 11.800 206.600 12.200 ;
        RECT 200.600 9.100 201.000 9.200 ;
        RECT 201.400 9.100 201.800 9.200 ;
        RECT 198.200 6.800 198.600 7.200 ;
        RECT 195.800 5.800 196.200 6.200 ;
        RECT 199.000 3.100 199.400 8.900 ;
        RECT 200.600 8.800 201.800 9.100 ;
        RECT 202.200 5.100 202.600 7.900 ;
        RECT 203.800 3.100 204.200 8.900 ;
        RECT 204.600 8.800 205.000 9.200 ;
        RECT 206.200 7.200 206.500 11.800 ;
        RECT 206.200 6.800 206.600 7.200 ;
        RECT 205.400 6.100 205.800 6.200 ;
        RECT 206.200 6.100 206.600 6.200 ;
        RECT 205.400 5.800 206.600 6.100 ;
        RECT 208.600 3.100 209.000 8.900 ;
        RECT 211.000 8.800 211.400 9.200 ;
        RECT 211.000 8.200 211.300 8.800 ;
        RECT 211.000 7.800 211.400 8.200 ;
        RECT 213.400 7.200 213.700 14.800 ;
        RECT 215.000 12.100 215.400 17.900 ;
        RECT 218.200 15.800 218.600 16.200 ;
        RECT 218.200 15.200 218.500 15.800 ;
        RECT 218.200 14.800 218.600 15.200 ;
        RECT 219.000 12.800 219.400 13.200 ;
        RECT 219.000 12.200 219.300 12.800 ;
        RECT 219.000 11.800 219.400 12.200 ;
        RECT 219.800 12.100 220.200 17.900 ;
        RECT 218.200 7.800 218.600 8.200 ;
        RECT 218.200 7.200 218.500 7.800 ;
        RECT 219.000 7.200 219.300 11.800 ;
        RECT 220.600 10.200 220.900 25.800 ;
        RECT 224.600 23.100 225.000 28.900 ;
        RECT 226.200 26.200 226.500 29.800 ;
        RECT 227.000 29.200 227.300 34.800 ;
        RECT 227.000 28.800 227.400 29.200 ;
        RECT 226.200 25.800 226.600 26.200 ;
        RECT 229.400 23.100 229.800 28.900 ;
        RECT 230.200 27.200 230.500 43.800 ;
        RECT 240.600 43.100 241.000 48.900 ;
        RECT 244.600 47.800 245.000 48.200 ;
        RECT 243.800 46.800 244.200 47.200 ;
        RECT 243.800 46.200 244.100 46.800 ;
        RECT 241.400 45.800 241.800 46.200 ;
        RECT 243.800 45.800 244.200 46.200 ;
        RECT 241.400 44.200 241.700 45.800 ;
        RECT 241.400 43.800 241.800 44.200 ;
        RECT 232.600 36.800 233.000 37.200 ;
        RECT 235.000 37.100 235.400 37.200 ;
        RECT 235.800 37.100 236.200 37.200 ;
        RECT 235.000 36.800 236.200 37.100 ;
        RECT 236.600 36.800 237.000 37.200 ;
        RECT 232.600 36.200 232.900 36.800 ;
        RECT 232.600 35.800 233.000 36.200 ;
        RECT 235.000 35.800 235.400 36.200 ;
        RECT 235.000 35.200 235.300 35.800 ;
        RECT 236.600 35.200 236.900 36.800 ;
        RECT 231.000 34.800 231.400 35.200 ;
        RECT 235.000 34.800 235.400 35.200 ;
        RECT 236.600 34.800 237.000 35.200 ;
        RECT 231.000 34.200 231.300 34.800 ;
        RECT 231.000 33.800 231.400 34.200 ;
        RECT 235.800 33.800 236.200 34.200 ;
        RECT 232.600 31.800 233.000 32.200 ;
        RECT 232.600 28.200 232.900 31.800 ;
        RECT 235.800 31.200 236.100 33.800 ;
        RECT 239.000 32.100 239.400 37.900 ;
        RECT 241.400 36.800 241.800 37.200 ;
        RECT 241.400 35.200 241.700 36.800 ;
        RECT 241.400 34.800 241.800 35.200 ;
        RECT 239.800 33.800 240.200 34.200 ;
        RECT 235.800 30.800 236.200 31.200 ;
        RECT 233.400 29.100 233.800 29.200 ;
        RECT 234.200 29.100 234.600 29.200 ;
        RECT 233.400 28.800 234.600 29.100 ;
        RECT 230.200 26.800 230.600 27.200 ;
        RECT 222.200 21.800 222.600 22.200 ;
        RECT 221.400 13.100 221.800 15.900 ;
        RECT 222.200 15.200 222.500 21.800 ;
        RECT 227.800 20.800 228.200 21.200 ;
        RECT 227.000 16.800 227.400 17.200 ;
        RECT 227.000 16.200 227.300 16.800 ;
        RECT 227.000 15.800 227.400 16.200 ;
        RECT 222.200 14.800 222.600 15.200 ;
        RECT 224.600 14.800 225.000 15.200 ;
        RECT 224.600 14.200 224.900 14.800 ;
        RECT 224.600 13.800 225.000 14.200 ;
        RECT 225.400 13.800 225.800 14.200 ;
        RECT 225.400 10.200 225.700 13.800 ;
        RECT 226.200 11.800 226.600 12.200 ;
        RECT 220.600 9.800 221.000 10.200 ;
        RECT 225.400 9.800 225.800 10.200 ;
        RECT 225.400 8.800 225.800 9.200 ;
        RECT 225.400 7.200 225.700 8.800 ;
        RECT 213.400 6.800 213.800 7.200 ;
        RECT 215.000 6.800 215.400 7.200 ;
        RECT 218.200 6.800 218.600 7.200 ;
        RECT 219.000 6.800 219.400 7.200 ;
        RECT 225.400 6.800 225.800 7.200 ;
        RECT 215.000 6.200 215.300 6.800 ;
        RECT 214.200 5.800 214.600 6.200 ;
        RECT 215.000 5.800 215.400 6.200 ;
        RECT 214.200 5.200 214.500 5.800 ;
        RECT 226.200 5.200 226.500 11.800 ;
        RECT 227.000 8.100 227.300 15.800 ;
        RECT 227.800 15.200 228.100 20.800 ;
        RECT 228.600 15.800 229.000 16.200 ;
        RECT 228.600 15.200 228.900 15.800 ;
        RECT 227.800 14.800 228.200 15.200 ;
        RECT 228.600 14.800 229.000 15.200 ;
        RECT 227.000 7.800 228.100 8.100 ;
        RECT 227.000 6.800 227.400 7.200 ;
        RECT 227.000 6.200 227.300 6.800 ;
        RECT 227.800 6.200 228.100 7.800 ;
        RECT 228.600 7.200 228.900 14.800 ;
        RECT 230.200 10.200 230.500 26.800 ;
        RECT 231.000 25.100 231.400 27.900 ;
        RECT 232.600 27.800 233.000 28.200 ;
        RECT 231.800 21.800 232.200 22.200 ;
        RECT 231.800 15.200 232.100 21.800 ;
        RECT 232.600 19.200 232.900 27.800 ;
        RECT 235.800 23.100 236.200 28.900 ;
        RECT 239.800 28.200 240.100 33.800 ;
        RECT 243.800 32.100 244.200 37.900 ;
        RECT 244.600 34.200 244.900 47.800 ;
        RECT 245.400 43.100 245.800 48.900 ;
        RECT 246.200 48.800 246.600 49.200 ;
        RECT 247.800 48.800 248.200 49.200 ;
        RECT 248.600 48.800 249.000 49.200 ;
        RECT 244.600 33.800 245.000 34.200 ;
        RECT 245.400 33.100 245.800 35.900 ;
        RECT 246.200 34.200 246.500 48.800 ;
        RECT 249.400 48.200 249.700 61.800 ;
        RECT 251.000 55.800 251.400 56.200 ;
        RECT 251.000 55.200 251.300 55.800 ;
        RECT 251.000 54.800 251.400 55.200 ;
        RECT 250.200 51.800 250.600 52.200 ;
        RECT 250.200 49.100 250.500 51.800 ;
        RECT 251.800 50.100 252.100 90.800 ;
        RECT 255.800 89.200 256.100 105.800 ;
        RECT 259.000 103.100 259.400 108.900 ;
        RECT 260.600 107.200 260.900 129.800 ;
        RECT 262.200 129.100 262.600 129.200 ;
        RECT 263.000 129.100 263.400 129.200 ;
        RECT 262.200 128.800 263.400 129.100 ;
        RECT 263.800 119.100 264.200 119.200 ;
        RECT 264.600 119.100 265.000 119.200 ;
        RECT 263.800 118.800 265.000 119.100 ;
        RECT 262.200 112.100 262.600 117.900 ;
        RECT 263.800 113.800 264.200 114.200 ;
        RECT 260.600 106.800 261.000 107.200 ;
        RECT 262.200 106.800 262.600 107.200 ;
        RECT 262.200 106.200 262.500 106.800 ;
        RECT 262.200 105.800 262.600 106.200 ;
        RECT 261.400 101.800 261.800 102.200 ;
        RECT 261.400 97.200 261.700 101.800 ;
        RECT 261.400 96.800 261.800 97.200 ;
        RECT 262.200 94.800 262.600 95.200 ;
        RECT 258.200 93.100 258.600 93.200 ;
        RECT 259.000 93.100 259.400 93.200 ;
        RECT 258.200 92.800 259.400 93.100 ;
        RECT 260.600 91.800 261.000 92.200 ;
        RECT 255.800 88.800 256.200 89.200 ;
        RECT 255.000 88.100 255.400 88.200 ;
        RECT 255.800 88.100 256.200 88.200 ;
        RECT 255.000 87.800 256.200 88.100 ;
        RECT 255.800 87.100 256.200 87.200 ;
        RECT 256.600 87.100 257.000 87.200 ;
        RECT 255.800 86.800 257.000 87.100 ;
        RECT 257.400 86.800 257.800 87.200 ;
        RECT 258.200 86.800 258.600 87.200 ;
        RECT 257.400 86.200 257.700 86.800 ;
        RECT 257.400 85.800 257.800 86.200 ;
        RECT 258.200 85.200 258.500 86.800 ;
        RECT 260.600 86.200 260.900 91.800 ;
        RECT 262.200 90.200 262.500 94.800 ;
        RECT 262.200 89.800 262.600 90.200 ;
        RECT 263.800 89.200 264.100 113.800 ;
        RECT 263.800 88.800 264.200 89.200 ;
        RECT 260.600 85.800 261.000 86.200 ;
        RECT 253.400 84.800 253.800 85.200 ;
        RECT 258.200 84.800 258.600 85.200 ;
        RECT 253.400 82.200 253.700 84.800 ;
        RECT 253.400 82.100 253.800 82.200 ;
        RECT 252.600 81.800 253.800 82.100 ;
        RECT 263.800 81.800 264.200 82.200 ;
        RECT 252.600 74.200 252.900 81.800 ;
        RECT 252.600 73.800 253.000 74.200 ;
        RECT 253.400 72.100 253.800 77.900 ;
        RECT 254.200 75.800 254.600 76.200 ;
        RECT 252.600 67.800 253.000 68.200 ;
        RECT 252.600 65.200 252.900 67.800 ;
        RECT 254.200 66.200 254.500 75.800 ;
        RECT 255.000 73.100 255.400 75.900 ;
        RECT 255.800 72.100 256.200 72.200 ;
        RECT 256.600 72.100 257.000 72.200 ;
        RECT 255.800 71.800 257.000 72.100 ;
        RECT 257.400 71.800 257.800 72.200 ;
        RECT 258.200 72.100 258.600 77.900 ;
        RECT 261.400 74.800 261.800 75.200 ;
        RECT 255.000 68.800 255.400 69.200 ;
        RECT 255.800 68.800 256.200 69.200 ;
        RECT 255.000 67.200 255.300 68.800 ;
        RECT 255.800 67.200 256.100 68.800 ;
        RECT 255.000 66.800 255.400 67.200 ;
        RECT 255.800 66.800 256.200 67.200 ;
        RECT 254.200 65.800 254.600 66.200 ;
        RECT 252.600 64.800 253.000 65.200 ;
        RECT 254.200 64.800 254.600 65.200 ;
        RECT 254.200 64.200 254.500 64.800 ;
        RECT 254.200 63.800 254.600 64.200 ;
        RECT 255.000 58.200 255.300 66.800 ;
        RECT 255.800 62.800 256.200 63.200 ;
        RECT 255.800 59.200 256.100 62.800 ;
        RECT 255.800 58.800 256.200 59.200 ;
        RECT 255.000 57.800 255.400 58.200 ;
        RECT 253.400 56.800 253.800 57.200 ;
        RECT 253.400 55.200 253.700 56.800 ;
        RECT 257.400 55.200 257.700 71.800 ;
        RECT 258.200 63.100 258.600 68.900 ;
        RECT 260.600 65.800 261.000 66.200 ;
        RECT 260.600 65.200 260.900 65.800 ;
        RECT 260.600 64.800 261.000 65.200 ;
        RECT 261.400 59.200 261.700 74.800 ;
        RECT 263.000 72.100 263.400 77.900 ;
        RECT 263.800 74.200 264.100 81.800 ;
        RECT 263.800 73.800 264.200 74.200 ;
        RECT 262.200 66.800 262.600 67.200 ;
        RECT 261.400 58.800 261.800 59.200 ;
        RECT 260.600 57.800 261.000 58.200 ;
        RECT 258.200 57.100 258.600 57.200 ;
        RECT 259.000 57.100 259.400 57.200 ;
        RECT 258.200 56.800 259.400 57.100 ;
        RECT 259.000 56.100 259.400 56.200 ;
        RECT 259.800 56.100 260.200 56.200 ;
        RECT 259.000 55.800 260.200 56.100 ;
        RECT 253.400 54.800 253.800 55.200 ;
        RECT 254.200 55.100 254.600 55.200 ;
        RECT 255.000 55.100 255.400 55.200 ;
        RECT 254.200 54.800 255.400 55.100 ;
        RECT 256.600 54.800 257.000 55.200 ;
        RECT 257.400 54.800 257.800 55.200 ;
        RECT 256.600 54.200 256.900 54.800 ;
        RECT 257.400 54.200 257.700 54.800 ;
        RECT 260.600 54.200 260.900 57.800 ;
        RECT 252.600 53.800 253.000 54.200 ;
        RECT 256.600 53.800 257.000 54.200 ;
        RECT 257.400 53.800 257.800 54.200 ;
        RECT 259.800 53.800 260.200 54.200 ;
        RECT 260.600 54.100 261.000 54.200 ;
        RECT 260.600 53.800 261.700 54.100 ;
        RECT 252.600 51.200 252.900 53.800 ;
        RECT 252.600 50.800 253.000 51.200 ;
        RECT 259.000 50.800 259.400 51.200 ;
        RECT 251.800 49.800 252.900 50.100 ;
        RECT 250.200 48.800 251.300 49.100 ;
        RECT 247.000 45.100 247.400 47.900 ;
        RECT 249.400 47.800 249.800 48.200 ;
        RECT 247.800 45.800 248.200 46.200 ;
        RECT 247.800 42.200 248.100 45.800 ;
        RECT 250.200 45.100 250.600 47.900 ;
        RECT 251.000 46.200 251.300 48.800 ;
        RECT 251.000 45.800 251.400 46.200 ;
        RECT 250.200 42.800 250.600 43.200 ;
        RECT 251.800 43.100 252.200 48.900 ;
        RECT 252.600 48.200 252.900 49.800 ;
        RECT 259.000 49.200 259.300 50.800 ;
        RECT 252.600 47.800 253.000 48.200 ;
        RECT 252.600 46.800 253.000 47.200 ;
        RECT 252.600 46.300 252.900 46.800 ;
        RECT 252.600 45.900 253.000 46.300 ;
        RECT 253.400 45.800 253.800 46.200 ;
        RECT 247.800 41.800 248.200 42.200 ;
        RECT 247.000 39.800 247.400 40.200 ;
        RECT 249.400 39.800 249.800 40.200 ;
        RECT 247.000 35.200 247.300 39.800 ;
        RECT 249.400 36.200 249.700 39.800 ;
        RECT 249.400 35.800 249.800 36.200 ;
        RECT 247.000 34.800 247.400 35.200 ;
        RECT 249.400 34.800 249.800 35.200 ;
        RECT 249.400 34.200 249.700 34.800 ;
        RECT 246.200 33.800 246.600 34.200 ;
        RECT 249.400 33.800 249.800 34.200 ;
        RECT 246.200 31.200 246.500 33.800 ;
        RECT 246.200 30.800 246.600 31.200 ;
        RECT 247.800 30.800 248.200 31.200 ;
        RECT 239.800 27.800 240.200 28.200 ;
        RECT 238.200 27.100 238.600 27.200 ;
        RECT 239.000 27.100 239.400 27.200 ;
        RECT 238.200 26.800 239.400 27.100 ;
        RECT 239.800 26.800 240.200 27.200 ;
        RECT 232.600 18.800 233.000 19.200 ;
        RECT 231.000 14.800 231.400 15.200 ;
        RECT 231.800 14.800 232.200 15.200 ;
        RECT 231.000 14.200 231.300 14.800 ;
        RECT 231.000 13.800 231.400 14.200 ;
        RECT 235.000 12.100 235.400 17.900 ;
        RECT 237.400 15.100 237.800 15.200 ;
        RECT 238.200 15.100 238.600 15.200 ;
        RECT 237.400 14.800 238.600 15.100 ;
        RECT 239.000 14.200 239.300 26.800 ;
        RECT 239.800 26.300 240.100 26.800 ;
        RECT 239.800 25.900 240.200 26.300 ;
        RECT 240.600 23.100 241.000 28.900 ;
        RECT 243.000 28.800 243.400 29.200 ;
        RECT 242.200 25.100 242.600 27.900 ;
        RECT 243.000 27.200 243.300 28.800 ;
        RECT 247.800 27.200 248.100 30.800 ;
        RECT 248.600 29.800 249.000 30.200 ;
        RECT 243.000 26.800 243.400 27.200 ;
        RECT 244.600 26.800 245.000 27.200 ;
        RECT 247.800 26.800 248.200 27.200 ;
        RECT 244.600 26.200 244.900 26.800 ;
        RECT 244.600 25.800 245.000 26.200 ;
        RECT 247.000 25.800 247.400 26.200 ;
        RECT 247.000 25.200 247.300 25.800 ;
        RECT 243.800 25.100 244.200 25.200 ;
        RECT 244.600 25.100 245.000 25.200 ;
        RECT 243.800 24.800 245.000 25.100 ;
        RECT 247.000 24.800 247.400 25.200 ;
        RECT 239.000 13.800 239.400 14.200 ;
        RECT 239.800 12.100 240.200 17.900 ;
        RECT 241.400 13.100 241.800 15.900 ;
        RECT 247.800 14.200 248.100 26.800 ;
        RECT 248.600 26.200 248.900 29.800 ;
        RECT 250.200 29.200 250.500 42.800 ;
        RECT 251.000 36.800 251.400 37.200 ;
        RECT 251.000 34.200 251.300 36.800 ;
        RECT 251.000 33.800 251.400 34.200 ;
        RECT 250.200 28.800 250.600 29.200 ;
        RECT 251.000 26.200 251.300 33.800 ;
        RECT 253.400 29.200 253.700 45.800 ;
        RECT 256.600 43.100 257.000 48.900 ;
        RECT 259.000 48.800 259.400 49.200 ;
        RECT 259.800 47.200 260.100 53.800 ;
        RECT 261.400 47.200 261.700 53.800 ;
        RECT 259.800 46.800 260.200 47.200 ;
        RECT 261.400 46.800 261.800 47.200 ;
        RECT 259.800 46.200 260.100 46.800 ;
        RECT 259.800 45.800 260.200 46.200 ;
        RECT 260.600 45.100 261.000 45.200 ;
        RECT 261.400 45.100 261.800 45.200 ;
        RECT 260.600 44.800 261.800 45.100 ;
        RECT 259.800 44.100 260.200 44.200 ;
        RECT 260.600 44.100 261.000 44.200 ;
        RECT 259.800 43.800 261.000 44.100 ;
        RECT 254.200 32.100 254.600 37.900 ;
        RECT 256.600 35.100 257.000 35.200 ;
        RECT 257.400 35.100 257.800 35.200 ;
        RECT 256.600 34.800 257.800 35.100 ;
        RECT 256.600 33.800 257.000 34.200 ;
        RECT 253.400 28.800 253.800 29.200 ;
        RECT 253.400 27.800 253.800 28.200 ;
        RECT 248.600 25.800 249.000 26.200 ;
        RECT 249.400 26.100 249.800 26.200 ;
        RECT 250.200 26.100 250.600 26.200 ;
        RECT 249.400 25.800 250.600 26.100 ;
        RECT 251.000 25.800 251.400 26.200 ;
        RECT 252.600 25.800 253.000 26.200 ;
        RECT 250.200 17.800 250.600 18.200 ;
        RECT 250.200 15.200 250.500 17.800 ;
        RECT 251.800 16.800 252.200 17.200 ;
        RECT 251.800 16.200 252.100 16.800 ;
        RECT 251.800 15.800 252.200 16.200 ;
        RECT 250.200 14.800 250.600 15.200 ;
        RECT 251.000 15.100 251.400 15.200 ;
        RECT 251.800 15.100 252.200 15.200 ;
        RECT 251.000 14.800 252.200 15.100 ;
        RECT 242.200 13.800 242.600 14.200 ;
        RECT 247.800 13.800 248.200 14.200 ;
        RECT 248.600 14.100 249.000 14.200 ;
        RECT 249.400 14.100 249.800 14.200 ;
        RECT 248.600 13.800 249.800 14.100 ;
        RECT 229.400 9.800 229.800 10.200 ;
        RECT 230.200 9.800 230.600 10.200 ;
        RECT 237.400 9.800 237.800 10.200 ;
        RECT 229.400 9.200 229.700 9.800 ;
        RECT 229.400 8.800 229.800 9.200 ;
        RECT 228.600 6.800 229.000 7.200 ;
        RECT 227.000 5.800 227.400 6.200 ;
        RECT 227.800 5.800 228.200 6.200 ;
        RECT 214.200 4.800 214.600 5.200 ;
        RECT 216.600 5.100 217.000 5.200 ;
        RECT 217.400 5.100 217.800 5.200 ;
        RECT 216.600 4.800 217.800 5.100 ;
        RECT 226.200 4.800 226.600 5.200 ;
        RECT 231.800 3.100 232.200 8.900 ;
        RECT 234.200 6.100 234.600 6.200 ;
        RECT 235.000 6.100 235.400 6.200 ;
        RECT 234.200 5.800 235.400 6.100 ;
        RECT 236.600 3.100 237.000 8.900 ;
        RECT 237.400 7.200 237.700 9.800 ;
        RECT 242.200 9.200 242.500 13.800 ;
        RECT 247.800 11.800 248.200 12.200 ;
        RECT 247.800 10.200 248.100 11.800 ;
        RECT 247.800 9.800 248.200 10.200 ;
        RECT 242.200 8.800 242.600 9.200 ;
        RECT 243.800 9.100 244.200 9.200 ;
        RECT 244.600 9.100 245.000 9.200 ;
        RECT 243.800 8.800 245.000 9.100 ;
        RECT 246.200 8.800 246.600 9.200 ;
        RECT 237.400 6.800 237.800 7.200 ;
        RECT 238.200 5.100 238.600 7.900 ;
        RECT 246.200 7.200 246.500 8.800 ;
        RECT 246.200 6.800 246.600 7.200 ;
        RECT 250.200 5.200 250.500 14.800 ;
        RECT 252.600 14.200 252.900 25.800 ;
        RECT 253.400 19.200 253.700 27.800 ;
        RECT 255.800 23.100 256.200 28.900 ;
        RECT 256.600 24.200 256.900 33.800 ;
        RECT 259.000 32.100 259.400 37.900 ;
        RECT 259.800 34.800 260.200 35.200 ;
        RECT 259.800 26.300 260.100 34.800 ;
        RECT 260.600 33.100 261.000 35.900 ;
        RECT 261.400 35.200 261.700 44.800 ;
        RECT 261.400 34.800 261.800 35.200 ;
        RECT 261.400 33.800 261.800 34.200 ;
        RECT 261.400 31.200 261.700 33.800 ;
        RECT 261.400 30.800 261.800 31.200 ;
        RECT 262.200 29.100 262.500 66.800 ;
        RECT 263.000 63.100 263.400 68.900 ;
        RECT 263.800 67.200 264.100 73.800 ;
        RECT 264.600 73.100 265.000 75.900 ;
        RECT 263.800 66.800 264.200 67.200 ;
        RECT 264.600 65.100 265.000 67.900 ;
        RECT 263.000 56.800 263.400 57.200 ;
        RECT 263.000 56.200 263.300 56.800 ;
        RECT 263.000 55.800 263.400 56.200 ;
        RECT 264.600 44.800 265.000 45.200 ;
        RECT 264.600 44.200 264.900 44.800 ;
        RECT 264.600 43.800 265.000 44.200 ;
        RECT 263.000 41.800 263.400 42.200 ;
        RECT 263.000 35.200 263.300 41.800 ;
        RECT 263.800 35.800 264.200 36.200 ;
        RECT 263.000 34.800 263.400 35.200 ;
        RECT 259.800 25.900 260.200 26.300 ;
        RECT 256.600 23.800 257.000 24.200 ;
        RECT 255.000 19.800 255.400 20.200 ;
        RECT 255.000 19.200 255.300 19.800 ;
        RECT 253.400 18.800 253.800 19.200 ;
        RECT 255.000 18.800 255.400 19.200 ;
        RECT 254.200 17.800 254.600 18.200 ;
        RECT 254.200 16.200 254.500 17.800 ;
        RECT 256.600 17.200 256.900 23.800 ;
        RECT 260.600 23.100 261.000 28.900 ;
        RECT 261.400 28.800 262.500 29.100 ;
        RECT 263.000 33.800 263.400 34.200 ;
        RECT 261.400 27.200 261.700 28.800 ;
        RECT 261.400 26.800 261.800 27.200 ;
        RECT 262.200 25.100 262.600 27.900 ;
        RECT 256.600 16.800 257.000 17.200 ;
        RECT 254.200 15.800 254.600 16.200 ;
        RECT 252.600 13.800 253.000 14.200 ;
        RECT 252.600 9.100 252.900 13.800 ;
        RECT 257.400 12.100 257.800 17.900 ;
        RECT 259.800 15.100 260.200 15.200 ;
        RECT 260.600 15.100 261.000 15.200 ;
        RECT 259.800 14.800 261.000 15.100 ;
        RECT 261.400 12.800 261.800 13.200 ;
        RECT 253.400 9.100 253.800 9.200 ;
        RECT 252.600 8.800 253.800 9.100 ;
        RECT 251.800 6.100 252.200 6.200 ;
        RECT 252.600 6.100 253.000 6.200 ;
        RECT 251.800 5.800 253.000 6.100 ;
        RECT 250.200 4.800 250.600 5.200 ;
        RECT 255.800 3.100 256.200 8.900 ;
        RECT 256.600 6.800 257.000 7.200 ;
        RECT 259.800 6.800 260.200 7.200 ;
        RECT 256.600 6.200 256.900 6.800 ;
        RECT 259.800 6.300 260.100 6.800 ;
        RECT 256.600 5.800 257.000 6.200 ;
        RECT 259.800 5.900 260.200 6.300 ;
        RECT 260.600 3.100 261.000 8.900 ;
        RECT 261.400 7.200 261.700 12.800 ;
        RECT 262.200 12.100 262.600 17.900 ;
        RECT 261.400 6.800 261.800 7.200 ;
        RECT 262.200 5.100 262.600 7.900 ;
        RECT 263.000 6.200 263.300 33.800 ;
        RECT 263.800 28.200 264.100 35.800 ;
        RECT 263.800 27.800 264.200 28.200 ;
        RECT 263.800 13.100 264.200 15.900 ;
        RECT 263.000 5.800 263.400 6.200 ;
      LAYER via2 ;
        RECT 28.600 236.800 29.000 237.200 ;
        RECT 1.400 211.800 1.800 212.200 ;
        RECT 5.400 205.800 5.800 206.200 ;
        RECT 10.200 208.800 10.600 209.200 ;
        RECT 17.400 223.800 17.800 224.200 ;
        RECT 15.000 213.800 15.400 214.200 ;
        RECT 14.200 206.800 14.600 207.200 ;
        RECT 11.800 205.800 12.200 206.200 ;
        RECT 11.800 194.800 12.200 195.200 ;
        RECT 13.400 189.800 13.800 190.200 ;
        RECT 1.400 171.800 1.800 172.200 ;
        RECT 34.200 225.800 34.600 226.200 ;
        RECT 35.000 223.800 35.400 224.200 ;
        RECT 12.600 166.800 13.000 167.200 ;
        RECT 12.600 155.800 13.000 156.200 ;
        RECT 10.200 148.800 10.600 149.200 ;
        RECT 15.000 165.800 15.400 166.200 ;
        RECT 62.200 234.800 62.600 235.200 ;
        RECT 41.400 208.800 41.800 209.200 ;
        RECT 26.200 188.800 26.600 189.200 ;
        RECT 28.600 187.800 29.000 188.200 ;
        RECT 27.000 184.800 27.400 185.200 ;
        RECT 25.400 168.800 25.800 169.200 ;
        RECT 14.200 146.800 14.600 147.200 ;
        RECT 4.600 134.800 5.000 135.200 ;
        RECT 19.000 146.800 19.400 147.200 ;
        RECT 49.400 205.800 49.800 206.200 ;
        RECT 49.400 193.800 49.800 194.200 ;
        RECT 53.400 191.800 53.800 192.200 ;
        RECT 28.600 174.800 29.000 175.200 ;
        RECT 65.400 233.800 65.800 234.200 ;
        RECT 81.400 234.800 81.800 235.200 ;
        RECT 63.800 228.800 64.200 229.200 ;
        RECT 66.200 226.800 66.600 227.200 ;
        RECT 64.600 194.800 65.000 195.200 ;
        RECT 59.800 185.800 60.200 186.200 ;
        RECT 63.800 185.800 64.200 186.200 ;
        RECT 44.600 174.800 45.000 175.200 ;
        RECT 48.600 174.800 49.000 175.200 ;
        RECT 40.600 173.800 41.000 174.200 ;
        RECT 29.400 151.800 29.800 152.200 ;
        RECT 34.200 164.800 34.600 165.200 ;
        RECT 52.600 166.800 53.000 167.200 ;
        RECT 51.800 165.800 52.200 166.200 ;
        RECT 41.400 154.800 41.800 155.200 ;
        RECT 51.800 153.800 52.200 154.200 ;
        RECT 25.400 134.800 25.800 135.200 ;
        RECT 11.800 125.800 12.200 126.200 ;
        RECT 17.400 128.800 17.800 129.200 ;
        RECT 2.200 102.800 2.600 103.200 ;
        RECT 19.800 124.800 20.200 125.200 ;
        RECT 39.000 145.800 39.400 146.200 ;
        RECT 31.000 133.800 31.400 134.200 ;
        RECT 19.000 116.800 19.400 117.200 ;
        RECT 32.600 125.800 33.000 126.200 ;
        RECT 21.400 115.800 21.800 116.200 ;
        RECT 24.600 114.800 25.000 115.200 ;
        RECT 29.400 113.800 29.800 114.200 ;
        RECT 8.600 105.800 9.000 106.200 ;
        RECT 14.200 108.800 14.600 109.200 ;
        RECT 16.600 105.800 17.000 106.200 ;
        RECT 4.600 85.800 5.000 86.200 ;
        RECT 4.600 74.800 5.000 75.200 ;
        RECT 4.600 45.800 5.000 46.200 ;
        RECT 10.200 96.800 10.600 97.200 ;
        RECT 15.800 93.800 16.200 94.200 ;
        RECT 17.400 88.800 17.800 89.200 ;
        RECT 16.600 85.800 17.000 86.200 ;
        RECT 27.000 86.800 27.400 87.200 ;
        RECT 39.800 125.800 40.200 126.200 ;
        RECT 53.400 145.800 53.800 146.200 ;
        RECT 12.600 75.800 13.000 76.200 ;
        RECT 25.400 71.800 25.800 72.200 ;
        RECT 26.200 66.800 26.600 67.200 ;
        RECT 23.800 54.800 24.200 55.200 ;
        RECT 17.400 48.800 17.800 49.200 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 1.400 18.800 1.800 19.200 ;
        RECT 11.000 15.800 11.400 16.200 ;
        RECT 29.400 51.800 29.800 52.200 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 39.800 85.800 40.200 86.200 ;
        RECT 39.000 83.800 39.400 84.200 ;
        RECT 66.200 174.800 66.600 175.200 ;
        RECT 68.600 175.800 69.000 176.200 ;
        RECT 67.000 173.800 67.400 174.200 ;
        RECT 90.200 226.800 90.600 227.200 ;
        RECT 85.400 205.800 85.800 206.200 ;
        RECT 98.200 234.800 98.600 235.200 ;
        RECT 103.800 235.800 104.200 236.200 ;
        RECT 103.000 231.800 103.400 232.200 ;
        RECT 100.600 213.800 101.000 214.200 ;
        RECT 105.400 211.800 105.800 212.200 ;
        RECT 82.200 194.800 82.600 195.200 ;
        RECT 82.200 174.800 82.600 175.200 ;
        RECT 83.800 171.800 84.200 172.200 ;
        RECT 68.600 165.800 69.000 166.200 ;
        RECT 67.000 164.800 67.400 165.200 ;
        RECT 75.000 156.800 75.400 157.200 ;
        RECT 111.800 225.800 112.200 226.200 ;
        RECT 119.800 221.800 120.200 222.200 ;
        RECT 132.600 234.800 133.000 235.200 ;
        RECT 147.000 235.800 147.400 236.200 ;
        RECT 107.000 188.800 107.400 189.200 ;
        RECT 94.200 165.800 94.600 166.200 ;
        RECT 96.600 165.800 97.000 166.200 ;
        RECT 63.000 145.800 63.400 146.200 ;
        RECT 66.200 133.800 66.600 134.200 ;
        RECT 63.000 127.800 63.400 128.200 ;
        RECT 107.000 175.800 107.400 176.200 ;
        RECT 109.400 175.800 109.800 176.200 ;
        RECT 111.800 174.800 112.200 175.200 ;
        RECT 101.400 154.800 101.800 155.200 ;
        RECT 92.600 145.800 93.000 146.200 ;
        RECT 98.200 145.800 98.600 146.200 ;
        RECT 100.600 145.800 101.000 146.200 ;
        RECT 99.800 143.800 100.200 144.200 ;
        RECT 91.000 138.800 91.400 139.200 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 33.400 62.800 33.800 63.200 ;
        RECT 65.400 114.800 65.800 115.200 ;
        RECT 72.600 127.800 73.000 128.200 ;
        RECT 82.200 134.800 82.600 135.200 ;
        RECT 103.800 143.800 104.200 144.200 ;
        RECT 133.400 225.800 133.800 226.200 ;
        RECT 153.400 225.800 153.800 226.200 ;
        RECT 133.400 211.800 133.800 212.200 ;
        RECT 150.200 211.800 150.600 212.200 ;
        RECT 118.200 186.800 118.600 187.200 ;
        RECT 131.800 195.800 132.200 196.200 ;
        RECT 118.200 184.800 118.600 185.200 ;
        RECT 114.200 175.800 114.600 176.200 ;
        RECT 118.200 174.800 118.600 175.200 ;
        RECT 132.600 185.800 133.000 186.200 ;
        RECT 141.400 208.800 141.800 209.200 ;
        RECT 175.800 236.800 176.200 237.200 ;
        RECT 185.400 235.800 185.800 236.200 ;
        RECT 175.800 225.800 176.200 226.200 ;
        RECT 168.600 216.800 169.000 217.200 ;
        RECT 163.800 206.800 164.200 207.200 ;
        RECT 155.800 194.800 156.200 195.200 ;
        RECT 111.000 154.800 111.400 155.200 ;
        RECT 131.000 173.800 131.400 174.200 ;
        RECT 147.800 185.800 148.200 186.200 ;
        RECT 139.800 165.800 140.200 166.200 ;
        RECT 113.400 151.800 113.800 152.200 ;
        RECT 113.400 145.800 113.800 146.200 ;
        RECT 126.200 157.800 126.600 158.200 ;
        RECT 127.800 156.800 128.200 157.200 ;
        RECT 115.000 134.800 115.400 135.200 ;
        RECT 115.800 133.800 116.200 134.200 ;
        RECT 73.400 113.800 73.800 114.200 ;
        RECT 71.000 105.800 71.400 106.200 ;
        RECT 64.600 95.800 65.000 96.200 ;
        RECT 33.400 48.800 33.800 49.200 ;
        RECT 32.600 45.800 33.000 46.200 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 34.200 34.800 34.600 35.200 ;
        RECT 17.400 15.800 17.800 16.200 ;
        RECT 8.600 6.800 9.000 7.200 ;
        RECT 20.600 8.800 21.000 9.200 ;
        RECT 59.000 71.800 59.400 72.200 ;
        RECT 103.800 128.800 104.200 129.200 ;
        RECT 105.400 124.800 105.800 125.200 ;
        RECT 109.400 124.800 109.800 125.200 ;
        RECT 124.600 135.800 125.000 136.200 ;
        RECT 123.000 134.800 123.400 135.200 ;
        RECT 117.400 126.800 117.800 127.200 ;
        RECT 118.200 125.800 118.600 126.200 ;
        RECT 82.200 93.800 82.600 94.200 ;
        RECT 76.600 85.800 77.000 86.200 ;
        RECT 71.000 72.800 71.400 73.200 ;
        RECT 59.000 68.800 59.400 69.200 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 62.200 52.800 62.600 53.200 ;
        RECT 63.000 48.800 63.400 49.200 ;
        RECT 63.800 35.800 64.200 36.200 ;
        RECT 61.400 34.800 61.800 35.200 ;
        RECT 61.400 26.800 61.800 27.200 ;
        RECT 37.400 11.800 37.800 12.200 ;
        RECT 52.600 17.800 53.000 18.200 ;
        RECT 66.200 26.800 66.600 27.200 ;
        RECT 69.400 33.800 69.800 34.200 ;
        RECT 92.600 84.800 93.000 85.200 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 95.800 75.800 96.200 76.200 ;
        RECT 89.400 68.800 89.800 69.200 ;
        RECT 91.800 67.800 92.200 68.200 ;
        RECT 115.800 124.800 116.200 125.200 ;
        RECT 120.600 124.800 121.000 125.200 ;
        RECT 113.400 121.800 113.800 122.200 ;
        RECT 115.800 106.800 116.200 107.200 ;
        RECT 111.800 105.800 112.200 106.200 ;
        RECT 105.400 87.800 105.800 88.200 ;
        RECT 75.000 56.800 75.400 57.200 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 73.400 28.800 73.800 29.200 ;
        RECT 83.000 45.800 83.400 46.200 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 59.000 13.800 59.400 14.200 ;
        RECT 31.800 6.800 32.200 7.200 ;
        RECT 35.000 6.800 35.400 7.200 ;
        RECT 49.400 6.800 49.800 7.200 ;
        RECT 73.400 16.800 73.800 17.200 ;
        RECT 114.200 74.800 114.600 75.200 ;
        RECT 89.400 26.800 89.800 27.200 ;
        RECT 91.800 15.800 92.200 16.200 ;
        RECT 112.600 54.800 113.000 55.200 ;
        RECT 119.800 114.800 120.200 115.200 ;
        RECT 150.200 174.800 150.600 175.200 ;
        RECT 145.400 173.800 145.800 174.200 ;
        RECT 142.200 156.800 142.600 157.200 ;
        RECT 152.600 172.800 153.000 173.200 ;
        RECT 199.000 228.800 199.400 229.200 ;
        RECT 201.400 228.800 201.800 229.200 ;
        RECT 195.800 227.800 196.200 228.200 ;
        RECT 207.000 234.800 207.400 235.200 ;
        RECT 165.400 187.800 165.800 188.200 ;
        RECT 160.600 174.800 161.000 175.200 ;
        RECT 156.600 165.800 157.000 166.200 ;
        RECT 147.000 155.800 147.400 156.200 ;
        RECT 132.600 146.800 133.000 147.200 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 155.000 157.800 155.400 158.200 ;
        RECT 161.400 168.800 161.800 169.200 ;
        RECT 166.200 162.800 166.600 163.200 ;
        RECT 164.600 155.800 165.000 156.200 ;
        RECT 167.000 154.800 167.400 155.200 ;
        RECT 179.800 168.800 180.200 169.200 ;
        RECT 214.200 225.800 214.600 226.200 ;
        RECT 202.200 205.800 202.600 206.200 ;
        RECT 176.600 158.800 177.000 159.200 ;
        RECT 183.000 166.800 183.400 167.200 ;
        RECT 176.600 154.800 177.000 155.200 ;
        RECT 168.600 148.800 169.000 149.200 ;
        RECT 159.000 146.800 159.400 147.200 ;
        RECT 167.800 146.800 168.200 147.200 ;
        RECT 131.000 123.800 131.400 124.200 ;
        RECT 125.400 113.800 125.800 114.200 ;
        RECT 121.400 86.800 121.800 87.200 ;
        RECT 132.600 115.800 133.000 116.200 ;
        RECT 135.800 125.800 136.200 126.200 ;
        RECT 135.000 116.800 135.400 117.200 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 93.400 6.800 93.800 7.200 ;
        RECT 126.200 65.800 126.600 66.200 ;
        RECT 130.200 65.800 130.600 66.200 ;
        RECT 141.400 128.800 141.800 129.200 ;
        RECT 143.800 125.800 144.200 126.200 ;
        RECT 143.800 116.800 144.200 117.200 ;
        RECT 164.600 135.800 165.000 136.200 ;
        RECT 162.200 132.800 162.600 133.200 ;
        RECT 154.200 124.800 154.600 125.200 ;
        RECT 149.400 114.800 149.800 115.200 ;
        RECT 147.000 112.800 147.400 113.200 ;
        RECT 137.400 86.800 137.800 87.200 ;
        RECT 143.800 94.800 144.200 95.200 ;
        RECT 149.400 101.800 149.800 102.200 ;
        RECT 163.000 128.800 163.400 129.200 ;
        RECT 167.000 132.800 167.400 133.200 ;
        RECT 150.200 94.800 150.600 95.200 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 134.200 74.800 134.600 75.200 ;
        RECT 133.400 72.800 133.800 73.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 128.600 57.800 129.000 58.200 ;
        RECT 123.800 44.800 124.200 45.200 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 123.000 41.800 123.400 42.200 ;
        RECT 167.800 125.800 168.200 126.200 ;
        RECT 171.000 124.800 171.400 125.200 ;
        RECT 167.000 104.800 167.400 105.200 ;
        RECT 171.800 103.800 172.200 104.200 ;
        RECT 165.400 94.800 165.800 95.200 ;
        RECT 143.000 44.800 143.400 45.200 ;
        RECT 140.600 34.800 141.000 35.200 ;
        RECT 152.600 54.800 153.000 55.200 ;
        RECT 179.000 145.800 179.400 146.200 ;
        RECT 203.000 191.800 203.400 192.200 ;
        RECT 236.600 226.800 237.000 227.200 ;
        RECT 223.800 205.800 224.200 206.200 ;
        RECT 227.000 211.800 227.400 212.200 ;
        RECT 243.800 224.800 244.200 225.200 ;
        RECT 230.200 206.800 230.600 207.200 ;
        RECT 218.200 185.800 218.600 186.200 ;
        RECT 214.200 172.800 214.600 173.200 ;
        RECT 206.200 171.800 206.600 172.200 ;
        RECT 196.600 168.800 197.000 169.200 ;
        RECT 203.800 166.800 204.200 167.200 ;
        RECT 192.600 158.800 193.000 159.200 ;
        RECT 187.000 154.800 187.400 155.200 ;
        RECT 203.000 154.800 203.400 155.200 ;
        RECT 207.000 154.800 207.400 155.200 ;
        RECT 174.200 109.800 174.600 110.200 ;
        RECT 226.200 174.800 226.600 175.200 ;
        RECT 217.400 152.800 217.800 153.200 ;
        RECT 207.800 138.800 208.200 139.200 ;
        RECT 207.000 135.800 207.400 136.200 ;
        RECT 201.400 134.800 201.800 135.200 ;
        RECT 205.400 134.800 205.800 135.200 ;
        RECT 195.800 125.800 196.200 126.200 ;
        RECT 208.600 133.800 209.000 134.200 ;
        RECT 231.800 175.800 232.200 176.200 ;
        RECT 246.200 194.800 246.600 195.200 ;
        RECT 254.200 226.800 254.600 227.200 ;
        RECT 259.000 214.800 259.400 215.200 ;
        RECT 250.200 194.800 250.600 195.200 ;
        RECT 243.800 185.800 244.200 186.200 ;
        RECT 243.000 184.800 243.400 185.200 ;
        RECT 243.000 165.800 243.400 166.200 ;
        RECT 203.000 132.800 203.400 133.200 ;
        RECT 219.000 132.800 219.400 133.200 ;
        RECT 222.200 132.800 222.600 133.200 ;
        RECT 158.200 67.800 158.600 68.200 ;
        RECT 168.600 73.800 169.000 74.200 ;
        RECT 169.400 68.800 169.800 69.200 ;
        RECT 171.800 68.800 172.200 69.200 ;
        RECT 167.800 65.800 168.200 66.200 ;
        RECT 193.400 95.800 193.800 96.200 ;
        RECT 187.800 94.800 188.200 95.200 ;
        RECT 190.200 86.800 190.600 87.200 ;
        RECT 187.800 85.800 188.200 86.200 ;
        RECT 196.600 94.800 197.000 95.200 ;
        RECT 183.800 66.800 184.200 67.200 ;
        RECT 162.200 54.800 162.600 55.200 ;
        RECT 171.000 54.800 171.400 55.200 ;
        RECT 134.200 5.800 134.600 6.200 ;
        RECT 167.800 38.800 168.200 39.200 ;
        RECT 175.800 44.800 176.200 45.200 ;
        RECT 182.200 34.800 182.600 35.200 ;
        RECT 182.200 28.800 182.600 29.200 ;
        RECT 160.600 14.800 161.000 15.200 ;
        RECT 161.400 12.800 161.800 13.200 ;
        RECT 155.000 5.800 155.400 6.200 ;
        RECT 166.200 8.800 166.600 9.200 ;
        RECT 175.800 8.800 176.200 9.200 ;
        RECT 211.000 125.800 211.400 126.200 ;
        RECT 209.400 105.800 209.800 106.200 ;
        RECT 200.600 86.800 201.000 87.200 ;
        RECT 223.000 114.800 223.400 115.200 ;
        RECT 219.000 106.800 219.400 107.200 ;
        RECT 226.200 107.800 226.600 108.200 ;
        RECT 208.600 91.800 209.000 92.200 ;
        RECT 231.000 115.800 231.400 116.200 ;
        RECT 249.400 154.800 249.800 155.200 ;
        RECT 255.000 154.800 255.400 155.200 ;
        RECT 230.200 104.800 230.600 105.200 ;
        RECT 229.400 103.800 229.800 104.200 ;
        RECT 219.800 96.800 220.200 97.200 ;
        RECT 233.400 92.800 233.800 93.200 ;
        RECT 216.600 74.800 217.000 75.200 ;
        RECT 222.200 75.800 222.600 76.200 ;
        RECT 239.000 94.800 239.400 95.200 ;
        RECT 191.000 28.800 191.400 29.200 ;
        RECT 209.400 55.800 209.800 56.200 ;
        RECT 210.200 54.800 210.600 55.200 ;
        RECT 214.200 54.700 214.600 55.100 ;
        RECT 211.800 47.800 212.200 48.200 ;
        RECT 210.200 32.800 210.600 33.200 ;
        RECT 200.600 26.800 201.000 27.200 ;
        RECT 173.400 5.800 173.800 6.200 ;
        RECT 203.000 28.800 203.400 29.200 ;
        RECT 222.200 33.800 222.600 34.200 ;
        RECT 232.600 76.800 233.000 77.200 ;
        RECT 259.800 133.800 260.200 134.200 ;
        RECT 259.000 114.700 259.400 115.100 ;
        RECT 247.000 108.800 247.400 109.200 ;
        RECT 243.800 74.800 244.200 75.200 ;
        RECT 246.200 72.800 246.600 73.200 ;
        RECT 247.000 71.800 247.400 72.200 ;
        RECT 255.000 92.800 255.400 93.200 ;
        RECT 245.400 67.800 245.800 68.200 ;
        RECT 237.400 44.800 237.800 45.200 ;
        RECT 223.000 28.800 223.400 29.200 ;
        RECT 208.600 16.800 209.000 17.200 ;
        RECT 211.800 15.800 212.200 16.200 ;
        RECT 206.200 5.800 206.600 6.200 ;
        RECT 235.800 36.800 236.200 37.200 ;
        RECT 234.200 28.800 234.600 29.200 ;
        RECT 255.800 87.800 256.200 88.200 ;
        RECT 256.600 71.800 257.000 72.200 ;
        RECT 259.000 56.800 259.400 57.200 ;
        RECT 255.000 54.800 255.400 55.200 ;
        RECT 239.000 26.800 239.400 27.200 ;
        RECT 260.600 43.800 261.000 44.200 ;
        RECT 250.200 25.800 250.600 26.200 ;
        RECT 217.400 4.800 217.800 5.200 ;
      LAYER metal3 ;
        RECT 21.400 237.100 21.800 237.200 ;
        RECT 28.600 237.100 29.000 237.200 ;
        RECT 29.400 237.100 29.800 237.200 ;
        RECT 36.600 237.100 37.000 237.200 ;
        RECT 53.400 237.100 53.800 237.200 ;
        RECT 21.400 236.800 53.800 237.100 ;
        RECT 118.200 237.100 118.600 237.200 ;
        RECT 124.600 237.100 125.000 237.200 ;
        RECT 118.200 236.800 125.000 237.100 ;
        RECT 126.200 237.100 126.600 237.200 ;
        RECT 160.600 237.100 161.000 237.200 ;
        RECT 126.200 236.800 161.000 237.100 ;
        RECT 162.200 237.100 162.600 237.200 ;
        RECT 175.800 237.100 176.200 237.200 ;
        RECT 176.600 237.100 177.000 237.200 ;
        RECT 162.200 236.800 177.000 237.100 ;
        RECT 180.600 237.100 181.000 237.200 ;
        RECT 194.200 237.100 194.600 237.200 ;
        RECT 180.600 236.800 194.600 237.100 ;
        RECT 241.400 237.100 241.800 237.200 ;
        RECT 243.000 237.100 243.400 237.200 ;
        RECT 241.400 236.800 243.400 237.100 ;
        RECT 32.600 236.100 33.000 236.200 ;
        RECT 92.600 236.100 93.000 236.200 ;
        RECT 32.600 235.800 93.000 236.100 ;
        RECT 103.800 236.100 104.200 236.200 ;
        RECT 108.600 236.100 109.000 236.200 ;
        RECT 103.800 235.800 109.000 236.100 ;
        RECT 114.200 236.100 114.600 236.200 ;
        RECT 139.000 236.100 139.400 236.200 ;
        RECT 142.200 236.100 142.600 236.200 ;
        RECT 114.200 235.800 142.600 236.100 ;
        RECT 147.000 236.100 147.400 236.200 ;
        RECT 153.400 236.100 153.800 236.200 ;
        RECT 147.000 235.800 153.800 236.100 ;
        RECT 163.800 236.100 164.200 236.200 ;
        RECT 168.600 236.100 169.000 236.200 ;
        RECT 185.400 236.100 185.800 236.200 ;
        RECT 188.600 236.100 189.000 236.200 ;
        RECT 163.800 235.800 169.000 236.100 ;
        RECT 184.600 235.800 189.000 236.100 ;
        RECT 35.800 234.800 36.200 235.200 ;
        RECT 44.600 234.800 45.000 235.200 ;
        RECT 62.200 235.100 62.600 235.200 ;
        RECT 65.400 235.100 65.800 235.200 ;
        RECT 62.200 234.800 65.800 235.100 ;
        RECT 81.400 235.100 81.800 235.200 ;
        RECT 88.600 235.100 89.000 235.200 ;
        RECT 81.400 234.800 89.000 235.100 ;
        RECT 98.200 235.100 98.600 235.200 ;
        RECT 102.200 235.100 102.600 235.200 ;
        RECT 98.200 234.800 102.600 235.100 ;
        RECT 107.800 235.100 108.200 235.200 ;
        RECT 123.800 235.100 124.200 235.200 ;
        RECT 126.200 235.100 126.600 235.200 ;
        RECT 107.800 234.800 126.600 235.100 ;
        RECT 132.600 235.100 133.000 235.200 ;
        RECT 139.800 235.100 140.200 235.200 ;
        RECT 132.600 234.800 140.200 235.100 ;
        RECT 142.200 235.100 142.600 235.200 ;
        RECT 182.200 235.100 182.600 235.200 ;
        RECT 183.800 235.100 184.200 235.200 ;
        RECT 142.200 234.800 184.200 235.100 ;
        RECT 203.800 235.100 204.200 235.200 ;
        RECT 207.000 235.100 207.400 235.200 ;
        RECT 203.800 234.800 207.400 235.100 ;
        RECT 221.400 234.800 221.800 235.200 ;
        RECT 243.800 235.100 244.200 235.200 ;
        RECT 247.800 235.100 248.200 235.200 ;
        RECT 243.800 234.800 248.200 235.100 ;
        RECT 23.800 234.100 24.200 234.200 ;
        RECT 35.800 234.100 36.100 234.800 ;
        RECT 44.600 234.100 44.900 234.800 ;
        RECT 23.800 233.800 44.900 234.100 ;
        RECT 65.400 234.100 65.800 234.200 ;
        RECT 71.000 234.100 71.400 234.200 ;
        RECT 65.400 233.800 71.400 234.100 ;
        RECT 111.000 234.100 111.400 234.200 ;
        RECT 114.200 234.100 114.600 234.200 ;
        RECT 111.000 233.800 114.600 234.100 ;
        RECT 115.800 234.100 116.200 234.200 ;
        RECT 160.600 234.100 161.000 234.200 ;
        RECT 164.600 234.100 165.000 234.200 ;
        RECT 115.800 233.800 129.700 234.100 ;
        RECT 160.600 233.800 165.000 234.100 ;
        RECT 175.800 234.100 176.200 234.200 ;
        RECT 182.200 234.100 182.600 234.200 ;
        RECT 175.800 233.800 182.600 234.100 ;
        RECT 185.400 234.100 185.800 234.200 ;
        RECT 221.400 234.100 221.700 234.800 ;
        RECT 185.400 233.800 221.700 234.100 ;
        RECT 222.200 234.100 222.600 234.200 ;
        RECT 223.000 234.100 223.400 234.200 ;
        RECT 224.600 234.100 225.000 234.200 ;
        RECT 253.400 234.100 253.800 234.200 ;
        RECT 222.200 233.800 253.800 234.100 ;
        RECT 129.400 233.200 129.700 233.800 ;
        RECT 68.600 233.100 69.000 233.200 ;
        RECT 79.800 233.100 80.200 233.200 ;
        RECT 60.600 232.800 80.200 233.100 ;
        RECT 100.600 233.100 101.000 233.200 ;
        RECT 111.800 233.100 112.200 233.200 ;
        RECT 100.600 232.800 112.200 233.100 ;
        RECT 129.400 232.800 129.800 233.200 ;
        RECT 136.600 233.100 137.000 233.200 ;
        RECT 146.200 233.100 146.600 233.200 ;
        RECT 149.400 233.100 149.800 233.200 ;
        RECT 136.600 232.800 149.800 233.100 ;
        RECT 165.400 233.100 165.800 233.200 ;
        RECT 185.400 233.100 185.800 233.200 ;
        RECT 165.400 232.800 185.800 233.100 ;
        RECT 213.400 233.100 213.800 233.200 ;
        RECT 220.600 233.100 221.000 233.200 ;
        RECT 227.000 233.100 227.400 233.200 ;
        RECT 213.400 232.800 227.400 233.100 ;
        RECT 251.800 233.100 252.200 233.200 ;
        RECT 262.200 233.100 262.600 233.200 ;
        RECT 251.800 232.800 262.600 233.100 ;
        RECT 60.600 232.200 60.900 232.800 ;
        RECT 0.600 232.100 1.000 232.200 ;
        RECT 5.400 232.100 5.800 232.200 ;
        RECT 0.600 231.800 5.800 232.100 ;
        RECT 60.600 231.800 61.000 232.200 ;
        RECT 67.000 232.100 67.400 232.200 ;
        RECT 72.600 232.100 73.000 232.200 ;
        RECT 75.800 232.100 76.200 232.200 ;
        RECT 67.000 231.800 76.200 232.100 ;
        RECT 103.000 232.100 103.400 232.200 ;
        RECT 108.600 232.100 109.000 232.200 ;
        RECT 103.000 231.800 109.000 232.100 ;
        RECT 120.600 232.100 121.000 232.200 ;
        RECT 123.000 232.100 123.400 232.200 ;
        RECT 143.000 232.100 143.400 232.200 ;
        RECT 120.600 231.800 143.400 232.100 ;
        RECT 83.000 231.100 83.400 231.200 ;
        RECT 95.000 231.100 95.400 231.200 ;
        RECT 83.000 230.800 95.400 231.100 ;
        RECT 122.200 231.100 122.600 231.200 ;
        RECT 127.800 231.100 128.200 231.200 ;
        RECT 122.200 230.800 128.200 231.100 ;
        RECT 49.400 230.100 49.800 230.200 ;
        RECT 75.000 230.100 75.400 230.200 ;
        RECT 49.400 229.800 75.400 230.100 ;
        RECT 87.000 230.100 87.400 230.200 ;
        RECT 94.200 230.100 94.600 230.200 ;
        RECT 87.000 229.800 94.600 230.100 ;
        RECT 107.800 230.100 108.200 230.200 ;
        RECT 110.200 230.100 110.600 230.200 ;
        RECT 116.600 230.100 117.000 230.200 ;
        RECT 107.800 229.800 117.000 230.100 ;
        RECT 129.400 230.100 129.800 230.200 ;
        RECT 144.600 230.100 145.000 230.200 ;
        RECT 148.600 230.100 149.000 230.200 ;
        RECT 174.200 230.100 174.600 230.200 ;
        RECT 176.600 230.100 177.000 230.200 ;
        RECT 196.600 230.100 197.000 230.200 ;
        RECT 129.400 229.800 197.000 230.100 ;
        RECT 221.400 230.100 221.800 230.200 ;
        RECT 223.800 230.100 224.200 230.200 ;
        RECT 221.400 229.800 224.200 230.100 ;
        RECT 6.200 229.100 6.600 229.200 ;
        RECT 15.800 229.100 16.200 229.200 ;
        RECT 25.400 229.100 25.800 229.200 ;
        RECT 6.200 228.800 25.800 229.100 ;
        RECT 63.800 229.100 64.200 229.200 ;
        RECT 68.600 229.100 69.000 229.200 ;
        RECT 63.800 228.800 69.000 229.100 ;
        RECT 88.600 229.100 89.000 229.200 ;
        RECT 102.200 229.100 102.600 229.200 ;
        RECT 107.800 229.100 108.100 229.800 ;
        RECT 88.600 228.800 108.100 229.100 ;
        RECT 109.400 229.100 109.800 229.200 ;
        RECT 122.200 229.100 122.600 229.200 ;
        RECT 109.400 228.800 122.600 229.100 ;
        RECT 135.800 229.100 136.200 229.200 ;
        RECT 141.400 229.100 141.800 229.200 ;
        RECT 135.800 228.800 141.800 229.100 ;
        RECT 148.600 229.100 149.000 229.200 ;
        RECT 152.600 229.100 153.000 229.200 ;
        RECT 148.600 228.800 153.000 229.100 ;
        RECT 155.000 229.100 155.400 229.200 ;
        RECT 177.400 229.100 177.800 229.200 ;
        RECT 155.000 228.800 177.800 229.100 ;
        RECT 199.000 229.100 199.400 229.200 ;
        RECT 199.800 229.100 200.200 229.200 ;
        RECT 199.000 228.800 200.200 229.100 ;
        RECT 201.400 229.100 201.800 229.200 ;
        RECT 204.600 229.100 205.000 229.200 ;
        RECT 210.200 229.100 210.600 229.200 ;
        RECT 201.400 228.800 210.600 229.100 ;
        RECT 215.000 228.800 215.400 229.200 ;
        RECT 19.000 227.800 19.400 228.200 ;
        RECT 42.200 228.100 42.600 228.200 ;
        RECT 59.800 228.100 60.200 228.200 ;
        RECT 42.200 227.800 60.200 228.100 ;
        RECT 75.000 228.100 75.400 228.200 ;
        RECT 166.200 228.100 166.600 228.200 ;
        RECT 75.000 227.800 166.600 228.100 ;
        RECT 179.000 228.100 179.400 228.200 ;
        RECT 195.800 228.100 196.200 228.200 ;
        RECT 179.000 227.800 196.200 228.100 ;
        RECT 196.600 228.100 197.000 228.200 ;
        RECT 199.000 228.100 199.400 228.200 ;
        RECT 196.600 227.800 199.400 228.100 ;
        RECT 207.000 228.100 207.400 228.200 ;
        RECT 215.000 228.100 215.300 228.800 ;
        RECT 207.000 227.800 215.300 228.100 ;
        RECT 231.800 228.100 232.200 228.200 ;
        RECT 240.600 228.100 241.000 228.200 ;
        RECT 243.000 228.100 243.400 228.200 ;
        RECT 231.800 227.800 243.400 228.100 ;
        RECT 249.400 228.100 249.800 228.200 ;
        RECT 253.400 228.100 253.800 228.200 ;
        RECT 249.400 227.800 253.800 228.100 ;
        RECT 12.600 227.100 13.000 227.200 ;
        RECT 19.000 227.100 19.300 227.800 ;
        RECT 7.000 226.800 8.900 227.100 ;
        RECT 12.600 226.800 19.300 227.100 ;
        RECT 31.800 227.100 32.200 227.200 ;
        RECT 38.200 227.100 38.600 227.200 ;
        RECT 39.800 227.100 40.200 227.200 ;
        RECT 31.800 226.800 40.200 227.100 ;
        RECT 42.200 227.100 42.600 227.200 ;
        RECT 47.800 227.100 48.200 227.200 ;
        RECT 52.600 227.100 53.000 227.200 ;
        RECT 42.200 226.800 53.000 227.100 ;
        RECT 57.400 227.100 57.800 227.200 ;
        RECT 66.200 227.100 66.600 227.200 ;
        RECT 57.400 226.800 66.600 227.100 ;
        RECT 80.600 227.100 81.000 227.200 ;
        RECT 86.200 227.100 86.600 227.200 ;
        RECT 80.600 226.800 86.600 227.100 ;
        RECT 90.200 227.100 90.600 227.200 ;
        RECT 110.200 227.100 110.600 227.200 ;
        RECT 115.800 227.100 116.200 227.200 ;
        RECT 90.200 226.800 116.200 227.100 ;
        RECT 125.400 226.800 125.800 227.200 ;
        RECT 130.200 227.100 130.600 227.200 ;
        RECT 138.200 227.100 138.600 227.200 ;
        RECT 130.200 226.800 138.600 227.100 ;
        RECT 141.400 226.800 141.800 227.200 ;
        RECT 159.000 227.100 159.400 227.200 ;
        RECT 163.000 227.100 163.400 227.200 ;
        RECT 172.600 227.100 173.000 227.200 ;
        RECT 159.000 226.800 173.000 227.100 ;
        RECT 173.400 227.100 173.800 227.200 ;
        RECT 177.400 227.100 177.800 227.200 ;
        RECT 173.400 226.800 177.800 227.100 ;
        RECT 181.400 227.100 181.800 227.200 ;
        RECT 184.600 227.100 185.000 227.200 ;
        RECT 203.800 227.100 204.200 227.200 ;
        RECT 214.200 227.100 214.600 227.200 ;
        RECT 181.400 226.800 185.000 227.100 ;
        RECT 193.400 226.800 204.200 227.100 ;
        RECT 208.600 226.800 214.600 227.100 ;
        RECT 234.200 226.800 234.600 227.200 ;
        RECT 236.600 227.100 237.000 227.200 ;
        RECT 246.200 227.100 246.600 227.200 ;
        RECT 236.600 226.800 246.600 227.100 ;
        RECT 254.200 227.100 254.600 227.200 ;
        RECT 256.600 227.100 257.000 227.200 ;
        RECT 261.400 227.100 261.800 227.200 ;
        RECT 254.200 226.800 261.800 227.100 ;
        RECT 7.000 226.200 7.300 226.800 ;
        RECT 8.600 226.200 8.900 226.800 ;
        RECT 125.400 226.200 125.700 226.800 ;
        RECT 141.400 226.200 141.700 226.800 ;
        RECT 193.400 226.200 193.700 226.800 ;
        RECT 208.600 226.200 208.900 226.800 ;
        RECT 7.000 225.800 7.400 226.200 ;
        RECT 8.600 225.800 9.000 226.200 ;
        RECT 18.200 226.100 18.600 226.200 ;
        RECT 20.600 226.100 21.000 226.200 ;
        RECT 18.200 225.800 21.000 226.100 ;
        RECT 31.800 226.100 32.200 226.200 ;
        RECT 32.600 226.100 33.000 226.200 ;
        RECT 31.800 225.800 33.000 226.100 ;
        RECT 34.200 226.100 34.600 226.200 ;
        RECT 43.000 226.100 43.400 226.200 ;
        RECT 34.200 225.800 43.400 226.100 ;
        RECT 45.400 226.100 45.800 226.200 ;
        RECT 50.200 226.100 50.600 226.200 ;
        RECT 45.400 225.800 50.600 226.100 ;
        RECT 51.800 226.100 52.200 226.200 ;
        RECT 84.600 226.100 85.000 226.200 ;
        RECT 87.800 226.100 88.200 226.200 ;
        RECT 51.800 225.800 88.200 226.100 ;
        RECT 107.000 226.100 107.400 226.200 ;
        RECT 111.800 226.100 112.200 226.200 ;
        RECT 107.000 225.800 112.200 226.100 ;
        RECT 125.400 225.800 125.800 226.200 ;
        RECT 131.000 226.100 131.400 226.200 ;
        RECT 131.800 226.100 132.200 226.200 ;
        RECT 131.000 225.800 132.200 226.100 ;
        RECT 133.400 226.100 133.800 226.200 ;
        RECT 135.800 226.100 136.200 226.200 ;
        RECT 133.400 225.800 136.200 226.100 ;
        RECT 138.200 226.100 138.600 226.200 ;
        RECT 139.800 226.100 140.200 226.200 ;
        RECT 138.200 225.800 140.200 226.100 ;
        RECT 141.400 225.800 141.800 226.200 ;
        RECT 142.200 226.100 142.600 226.200 ;
        RECT 147.000 226.100 147.400 226.200 ;
        RECT 142.200 225.800 147.400 226.100 ;
        RECT 153.400 226.100 153.800 226.200 ;
        RECT 155.800 226.100 156.200 226.200 ;
        RECT 153.400 225.800 156.200 226.100 ;
        RECT 168.600 226.100 169.000 226.200 ;
        RECT 175.800 226.100 176.200 226.200 ;
        RECT 168.600 225.800 176.200 226.100 ;
        RECT 178.200 226.100 178.600 226.200 ;
        RECT 185.400 226.100 185.800 226.200 ;
        RECT 178.200 225.800 185.800 226.100 ;
        RECT 193.400 225.800 193.800 226.200 ;
        RECT 208.600 225.800 209.000 226.200 ;
        RECT 214.200 226.100 214.600 226.200 ;
        RECT 215.800 226.100 216.200 226.200 ;
        RECT 214.200 225.800 216.200 226.100 ;
        RECT 234.200 226.100 234.500 226.800 ;
        RECT 241.400 226.100 241.800 226.200 ;
        RECT 247.000 226.100 247.400 226.200 ;
        RECT 234.200 225.800 241.800 226.100 ;
        RECT 245.400 225.800 247.400 226.100 ;
        RECT 245.400 225.200 245.700 225.800 ;
        RECT 15.000 225.100 15.400 225.200 ;
        RECT 17.400 225.100 17.800 225.200 ;
        RECT 21.400 225.100 21.800 225.200 ;
        RECT 33.400 225.100 33.800 225.200 ;
        RECT 15.000 224.800 33.800 225.100 ;
        RECT 64.600 225.100 65.000 225.200 ;
        RECT 67.000 225.100 67.400 225.200 ;
        RECT 64.600 224.800 67.400 225.100 ;
        RECT 73.400 225.100 73.800 225.200 ;
        RECT 107.800 225.100 108.200 225.200 ;
        RECT 117.400 225.100 117.800 225.200 ;
        RECT 73.400 224.800 89.700 225.100 ;
        RECT 107.800 224.800 117.800 225.100 ;
        RECT 126.200 225.100 126.600 225.200 ;
        RECT 135.000 225.100 135.400 225.200 ;
        RECT 151.800 225.100 152.200 225.200 ;
        RECT 126.200 224.800 152.200 225.100 ;
        RECT 184.600 225.100 185.000 225.200 ;
        RECT 190.200 225.100 190.600 225.200 ;
        RECT 184.600 224.800 190.600 225.100 ;
        RECT 234.200 225.100 234.600 225.200 ;
        RECT 235.000 225.100 235.400 225.200 ;
        RECT 234.200 224.800 235.400 225.100 ;
        RECT 236.600 225.100 237.000 225.200 ;
        RECT 238.200 225.100 238.600 225.200 ;
        RECT 236.600 224.800 238.600 225.100 ;
        RECT 243.800 225.100 244.200 225.200 ;
        RECT 245.400 225.100 245.800 225.200 ;
        RECT 243.800 224.800 245.800 225.100 ;
        RECT 246.200 225.100 246.600 225.200 ;
        RECT 253.400 225.100 253.800 225.200 ;
        RECT 246.200 224.800 253.800 225.100 ;
        RECT 17.400 224.100 17.800 224.200 ;
        RECT 22.200 224.100 22.600 224.200 ;
        RECT 17.400 223.800 22.600 224.100 ;
        RECT 26.200 224.100 26.600 224.200 ;
        RECT 35.000 224.100 35.400 224.200 ;
        RECT 26.200 223.800 35.400 224.100 ;
        RECT 62.200 224.100 62.600 224.200 ;
        RECT 63.800 224.100 64.200 224.200 ;
        RECT 88.600 224.100 89.000 224.200 ;
        RECT 62.200 223.800 89.000 224.100 ;
        RECT 89.400 224.100 89.700 224.800 ;
        RECT 127.000 224.100 127.400 224.200 ;
        RECT 89.400 223.800 127.400 224.100 ;
        RECT 135.800 224.100 136.200 224.200 ;
        RECT 138.200 224.100 138.600 224.200 ;
        RECT 179.000 224.100 179.400 224.200 ;
        RECT 181.400 224.100 181.800 224.200 ;
        RECT 183.000 224.100 183.400 224.200 ;
        RECT 135.800 223.800 183.400 224.100 ;
        RECT 59.800 223.100 60.200 223.200 ;
        RECT 97.400 223.100 97.800 223.200 ;
        RECT 59.800 222.800 97.800 223.100 ;
        RECT 140.600 223.100 141.000 223.200 ;
        RECT 143.000 223.100 143.400 223.200 ;
        RECT 140.600 222.800 143.400 223.100 ;
        RECT 182.200 223.100 182.600 223.200 ;
        RECT 237.400 223.100 237.800 223.200 ;
        RECT 182.200 222.800 237.800 223.100 ;
        RECT 51.800 222.100 52.200 222.200 ;
        RECT 73.400 222.100 73.800 222.200 ;
        RECT 83.800 222.100 84.200 222.200 ;
        RECT 51.800 221.800 84.200 222.100 ;
        RECT 119.800 222.100 120.200 222.200 ;
        RECT 121.400 222.100 121.800 222.200 ;
        RECT 138.200 222.100 138.600 222.200 ;
        RECT 119.800 221.800 138.600 222.100 ;
        RECT 195.000 222.100 195.400 222.200 ;
        RECT 199.800 222.100 200.200 222.200 ;
        RECT 211.800 222.100 212.200 222.200 ;
        RECT 216.600 222.100 217.000 222.200 ;
        RECT 223.800 222.100 224.200 222.200 ;
        RECT 195.000 221.800 224.200 222.100 ;
        RECT 255.000 222.100 255.400 222.200 ;
        RECT 255.800 222.100 256.200 222.200 ;
        RECT 255.000 221.800 256.200 222.100 ;
        RECT 74.200 221.100 74.600 221.200 ;
        RECT 107.800 221.100 108.200 221.200 ;
        RECT 74.200 220.800 108.200 221.100 ;
        RECT 111.000 221.100 111.400 221.200 ;
        RECT 123.800 221.100 124.200 221.200 ;
        RECT 111.000 220.800 124.200 221.100 ;
        RECT 127.000 221.100 127.400 221.200 ;
        RECT 127.800 221.100 128.200 221.200 ;
        RECT 127.000 220.800 128.200 221.100 ;
        RECT 111.800 220.100 112.200 220.200 ;
        RECT 153.400 220.100 153.800 220.200 ;
        RECT 111.800 219.800 153.800 220.100 ;
        RECT 30.200 219.100 30.600 219.200 ;
        RECT 81.400 219.100 81.800 219.200 ;
        RECT 30.200 218.800 81.800 219.100 ;
        RECT 108.600 219.100 109.000 219.200 ;
        RECT 115.000 219.100 115.400 219.200 ;
        RECT 108.600 218.800 115.400 219.100 ;
        RECT 225.400 219.100 225.800 219.200 ;
        RECT 227.800 219.100 228.200 219.200 ;
        RECT 225.400 218.800 228.200 219.100 ;
        RECT 45.400 218.100 45.800 218.200 ;
        RECT 126.200 218.100 126.600 218.200 ;
        RECT 45.400 217.800 126.600 218.100 ;
        RECT 192.600 218.100 193.000 218.200 ;
        RECT 220.600 218.100 221.000 218.200 ;
        RECT 192.600 217.800 221.000 218.100 ;
        RECT 26.200 217.100 26.600 217.200 ;
        RECT 74.200 217.100 74.600 217.200 ;
        RECT 26.200 216.800 74.600 217.100 ;
        RECT 79.800 217.100 80.200 217.200 ;
        RECT 83.800 217.100 84.200 217.200 ;
        RECT 79.800 216.800 84.200 217.100 ;
        RECT 112.600 217.100 113.000 217.200 ;
        RECT 120.600 217.100 121.000 217.200 ;
        RECT 112.600 216.800 121.000 217.100 ;
        RECT 161.400 217.100 161.800 217.200 ;
        RECT 168.600 217.100 169.000 217.200 ;
        RECT 177.400 217.100 177.800 217.200 ;
        RECT 161.400 216.800 177.800 217.100 ;
        RECT 179.000 217.100 179.400 217.200 ;
        RECT 198.200 217.100 198.600 217.200 ;
        RECT 218.200 217.100 218.600 217.200 ;
        RECT 179.000 216.800 218.600 217.100 ;
        RECT 226.200 216.800 226.600 217.200 ;
        RECT 252.600 217.100 253.000 217.200 ;
        RECT 255.000 217.100 255.400 217.200 ;
        RECT 252.600 216.800 255.400 217.100 ;
        RECT 226.200 216.200 226.500 216.800 ;
        RECT 7.000 215.800 7.400 216.200 ;
        RECT 31.800 216.100 32.200 216.200 ;
        RECT 37.400 216.100 37.800 216.200 ;
        RECT 31.800 215.800 37.800 216.100 ;
        RECT 43.000 216.100 43.400 216.200 ;
        RECT 45.400 216.100 45.800 216.200 ;
        RECT 43.000 215.800 45.800 216.100 ;
        RECT 66.200 216.100 66.600 216.200 ;
        RECT 67.000 216.100 67.400 216.200 ;
        RECT 67.800 216.100 68.200 216.200 ;
        RECT 66.200 215.800 68.200 216.100 ;
        RECT 77.400 216.100 77.800 216.200 ;
        RECT 95.000 216.100 95.400 216.200 ;
        RECT 107.800 216.100 108.200 216.200 ;
        RECT 77.400 215.800 108.200 216.100 ;
        RECT 114.200 216.100 114.600 216.200 ;
        RECT 115.000 216.100 115.400 216.200 ;
        RECT 114.200 215.800 115.400 216.100 ;
        RECT 152.600 215.800 153.000 216.200 ;
        RECT 174.200 215.800 174.600 216.200 ;
        RECT 175.800 216.100 176.200 216.200 ;
        RECT 187.000 216.100 187.400 216.200 ;
        RECT 175.800 215.800 187.400 216.100 ;
        RECT 212.600 215.800 213.000 216.200 ;
        RECT 226.200 215.800 226.600 216.200 ;
        RECT 243.800 216.100 244.200 216.200 ;
        RECT 247.800 216.100 248.200 216.200 ;
        RECT 243.800 215.800 248.200 216.100 ;
        RECT 7.000 215.100 7.300 215.800 ;
        RECT 12.600 215.100 13.000 215.200 ;
        RECT 7.000 214.800 13.000 215.100 ;
        RECT 36.600 215.100 37.000 215.200 ;
        RECT 39.000 215.100 39.400 215.200 ;
        RECT 36.600 214.800 39.400 215.100 ;
        RECT 41.400 215.100 41.800 215.200 ;
        RECT 61.400 215.100 61.800 215.200 ;
        RECT 63.800 215.100 64.200 215.200 ;
        RECT 41.400 214.800 44.900 215.100 ;
        RECT 61.400 214.800 64.200 215.100 ;
        RECT 68.600 215.100 69.000 215.200 ;
        RECT 75.800 215.100 76.200 215.200 ;
        RECT 68.600 214.800 76.200 215.100 ;
        RECT 79.000 215.100 79.400 215.200 ;
        RECT 116.600 215.100 117.000 215.200 ;
        RECT 119.800 215.100 120.200 215.200 ;
        RECT 79.000 214.800 120.200 215.100 ;
        RECT 129.400 215.100 129.800 215.200 ;
        RECT 131.000 215.100 131.400 215.200 ;
        RECT 129.400 214.800 131.400 215.100 ;
        RECT 135.000 214.800 135.400 215.200 ;
        RECT 148.600 215.100 149.000 215.200 ;
        RECT 152.600 215.100 152.900 215.800 ;
        RECT 159.800 215.100 160.200 215.200 ;
        RECT 148.600 214.800 160.200 215.100 ;
        RECT 174.200 215.100 174.500 215.800 ;
        RECT 179.000 215.100 179.400 215.200 ;
        RECT 174.200 214.800 179.400 215.100 ;
        RECT 181.400 215.100 181.800 215.200 ;
        RECT 183.800 215.100 184.200 215.200 ;
        RECT 181.400 214.800 184.200 215.100 ;
        RECT 195.800 215.100 196.200 215.200 ;
        RECT 212.600 215.100 212.900 215.800 ;
        RECT 195.800 214.800 212.900 215.100 ;
        RECT 217.400 215.100 217.800 215.200 ;
        RECT 231.000 215.100 231.400 215.200 ;
        RECT 217.400 214.800 231.400 215.100 ;
        RECT 234.200 214.800 234.600 215.200 ;
        RECT 259.000 215.100 259.400 215.200 ;
        RECT 262.200 215.100 262.600 215.200 ;
        RECT 259.000 214.800 262.600 215.100 ;
        RECT 44.600 214.200 44.900 214.800 ;
        RECT 63.800 214.200 64.100 214.800 ;
        RECT 135.000 214.200 135.300 214.800 ;
        RECT 11.800 214.100 12.200 214.200 ;
        RECT 15.000 214.100 15.400 214.200 ;
        RECT 19.000 214.100 19.400 214.200 ;
        RECT 11.800 213.800 19.400 214.100 ;
        RECT 44.600 214.100 45.000 214.200 ;
        RECT 51.000 214.100 51.400 214.200 ;
        RECT 44.600 213.800 51.400 214.100 ;
        RECT 53.400 214.100 53.800 214.200 ;
        RECT 61.400 214.100 61.800 214.200 ;
        RECT 53.400 213.800 61.800 214.100 ;
        RECT 63.800 213.800 64.200 214.200 ;
        RECT 93.400 214.100 93.800 214.200 ;
        RECT 100.600 214.100 101.000 214.200 ;
        RECT 93.400 213.800 101.000 214.100 ;
        RECT 111.000 214.100 111.400 214.200 ;
        RECT 117.400 214.100 117.800 214.200 ;
        RECT 111.000 213.800 117.800 214.100 ;
        RECT 135.000 213.800 135.400 214.200 ;
        RECT 182.200 213.800 182.600 214.200 ;
        RECT 185.400 214.100 185.800 214.200 ;
        RECT 199.800 214.100 200.200 214.200 ;
        RECT 219.800 214.100 220.200 214.200 ;
        RECT 185.400 213.800 193.700 214.100 ;
        RECT 199.800 213.800 220.200 214.100 ;
        RECT 222.200 214.100 222.600 214.200 ;
        RECT 232.600 214.100 233.000 214.200 ;
        RECT 222.200 213.800 233.000 214.100 ;
        RECT 234.200 214.100 234.500 214.800 ;
        RECT 239.000 214.100 239.400 214.200 ;
        RECT 234.200 213.800 239.400 214.100 ;
        RECT 182.200 213.200 182.500 213.800 ;
        RECT 193.400 213.200 193.700 213.800 ;
        RECT 0.600 213.100 1.000 213.200 ;
        RECT 6.200 213.100 6.600 213.200 ;
        RECT 0.600 212.800 6.600 213.100 ;
        RECT 25.400 213.100 25.800 213.200 ;
        RECT 35.000 213.100 35.400 213.200 ;
        RECT 25.400 212.800 35.400 213.100 ;
        RECT 37.400 213.100 37.800 213.200 ;
        RECT 49.400 213.100 49.800 213.200 ;
        RECT 37.400 212.800 49.800 213.100 ;
        RECT 51.000 213.100 51.400 213.200 ;
        RECT 64.600 213.100 65.000 213.200 ;
        RECT 51.000 212.800 65.000 213.100 ;
        RECT 111.000 213.100 111.400 213.200 ;
        RECT 114.200 213.100 114.600 213.200 ;
        RECT 121.400 213.100 121.800 213.200 ;
        RECT 111.000 212.800 121.800 213.100 ;
        RECT 129.400 213.100 129.800 213.200 ;
        RECT 130.200 213.100 130.600 213.200 ;
        RECT 142.200 213.100 142.600 213.200 ;
        RECT 129.400 212.800 142.600 213.100 ;
        RECT 178.200 213.100 178.600 213.200 ;
        RECT 182.200 213.100 182.600 213.200 ;
        RECT 178.200 212.800 182.600 213.100 ;
        RECT 193.400 212.800 193.800 213.200 ;
        RECT 205.400 213.100 205.800 213.200 ;
        RECT 235.800 213.100 236.200 213.200 ;
        RECT 205.400 212.800 236.200 213.100 ;
        RECT 1.400 212.100 1.800 212.200 ;
        RECT 10.200 212.100 10.600 212.200 ;
        RECT 30.200 212.100 30.600 212.200 ;
        RECT 1.400 211.800 30.600 212.100 ;
        RECT 31.000 212.100 31.400 212.200 ;
        RECT 38.200 212.100 38.600 212.200 ;
        RECT 79.800 212.100 80.200 212.200 ;
        RECT 31.000 211.800 80.200 212.100 ;
        RECT 105.400 212.100 105.800 212.200 ;
        RECT 107.800 212.100 108.200 212.200 ;
        RECT 115.800 212.100 116.200 212.200 ;
        RECT 105.400 211.800 116.200 212.100 ;
        RECT 118.200 212.100 118.600 212.200 ;
        RECT 133.400 212.100 133.800 212.200 ;
        RECT 118.200 211.800 133.800 212.100 ;
        RECT 150.200 212.100 150.600 212.200 ;
        RECT 151.000 212.100 151.400 212.200 ;
        RECT 150.200 211.800 151.400 212.100 ;
        RECT 170.200 212.100 170.600 212.200 ;
        RECT 194.200 212.100 194.600 212.200 ;
        RECT 196.600 212.100 197.000 212.200 ;
        RECT 206.200 212.100 206.600 212.200 ;
        RECT 170.200 211.800 206.600 212.100 ;
        RECT 207.000 212.100 207.400 212.200 ;
        RECT 208.600 212.100 209.000 212.200 ;
        RECT 207.000 211.800 209.000 212.100 ;
        RECT 213.400 212.100 213.800 212.200 ;
        RECT 227.000 212.100 227.400 212.200 ;
        RECT 213.400 211.800 227.400 212.100 ;
        RECT 227.800 212.100 228.200 212.200 ;
        RECT 241.400 212.100 241.800 212.200 ;
        RECT 227.800 211.800 241.800 212.100 ;
        RECT 20.600 211.100 21.000 211.200 ;
        RECT 51.800 211.100 52.200 211.200 ;
        RECT 20.600 210.800 52.200 211.100 ;
        RECT 78.200 211.100 78.600 211.200 ;
        RECT 86.200 211.100 86.600 211.200 ;
        RECT 78.200 210.800 86.600 211.100 ;
        RECT 114.200 211.100 114.600 211.200 ;
        RECT 127.000 211.100 127.400 211.200 ;
        RECT 114.200 210.800 127.400 211.100 ;
        RECT 197.400 211.100 197.800 211.200 ;
        RECT 199.000 211.100 199.400 211.200 ;
        RECT 197.400 210.800 199.400 211.100 ;
        RECT 219.800 211.100 220.200 211.200 ;
        RECT 252.600 211.100 253.000 211.200 ;
        RECT 219.800 210.800 253.000 211.100 ;
        RECT 259.000 211.100 259.400 211.200 ;
        RECT 261.400 211.100 261.800 211.200 ;
        RECT 259.000 210.800 261.800 211.100 ;
        RECT 35.800 210.100 36.200 210.200 ;
        RECT 40.600 210.100 41.000 210.200 ;
        RECT 35.800 209.800 41.000 210.100 ;
        RECT 55.800 210.100 56.200 210.200 ;
        RECT 58.200 210.100 58.600 210.200 ;
        RECT 55.800 209.800 58.600 210.100 ;
        RECT 75.000 210.100 75.400 210.200 ;
        RECT 80.600 210.100 81.000 210.200 ;
        RECT 75.000 209.800 81.000 210.100 ;
        RECT 99.800 210.100 100.200 210.200 ;
        RECT 101.400 210.100 101.800 210.200 ;
        RECT 122.200 210.100 122.600 210.200 ;
        RECT 99.800 209.800 101.800 210.100 ;
        RECT 107.800 209.800 122.600 210.100 ;
        RECT 196.600 209.800 197.000 210.200 ;
        RECT 211.000 210.100 211.400 210.200 ;
        RECT 227.800 210.100 228.200 210.200 ;
        RECT 211.000 209.800 228.200 210.100 ;
        RECT 228.600 210.100 229.000 210.200 ;
        RECT 240.600 210.100 241.000 210.200 ;
        RECT 246.200 210.100 246.600 210.200 ;
        RECT 228.600 209.800 246.600 210.100 ;
        RECT 10.200 209.100 10.600 209.200 ;
        RECT 15.000 209.100 15.400 209.200 ;
        RECT 30.200 209.100 30.600 209.200 ;
        RECT 10.200 208.800 30.600 209.100 ;
        RECT 41.400 209.100 41.800 209.200 ;
        RECT 45.400 209.100 45.800 209.200 ;
        RECT 47.000 209.100 47.400 209.200 ;
        RECT 41.400 208.800 47.400 209.100 ;
        RECT 103.800 209.100 104.200 209.200 ;
        RECT 107.800 209.100 108.100 209.800 ;
        RECT 103.800 208.800 108.100 209.100 ;
        RECT 119.000 208.800 119.400 209.200 ;
        RECT 141.400 209.100 141.800 209.200 ;
        RECT 196.600 209.100 196.900 209.800 ;
        RECT 203.000 209.100 203.400 209.200 ;
        RECT 141.400 208.800 146.500 209.100 ;
        RECT 196.600 208.800 203.400 209.100 ;
        RECT 211.800 208.800 212.200 209.200 ;
        RECT 226.200 209.100 226.600 209.200 ;
        RECT 229.400 209.100 229.800 209.200 ;
        RECT 226.200 208.800 229.800 209.100 ;
        RECT 13.400 208.100 13.800 208.200 ;
        RECT 17.400 208.100 17.800 208.200 ;
        RECT 13.400 207.800 17.800 208.100 ;
        RECT 19.000 208.100 19.400 208.200 ;
        RECT 35.000 208.100 35.400 208.200 ;
        RECT 42.200 208.100 42.600 208.200 ;
        RECT 63.800 208.100 64.200 208.200 ;
        RECT 71.000 208.100 71.400 208.200 ;
        RECT 19.000 207.800 34.500 208.100 ;
        RECT 35.000 207.800 43.300 208.100 ;
        RECT 63.800 207.800 71.400 208.100 ;
        RECT 73.400 208.100 73.800 208.200 ;
        RECT 75.000 208.100 75.400 208.200 ;
        RECT 73.400 207.800 75.400 208.100 ;
        RECT 98.200 208.100 98.600 208.200 ;
        RECT 101.400 208.100 101.800 208.200 ;
        RECT 98.200 207.800 101.800 208.100 ;
        RECT 102.200 208.100 102.600 208.200 ;
        RECT 116.600 208.100 117.000 208.200 ;
        RECT 102.200 207.800 117.000 208.100 ;
        RECT 119.000 208.100 119.300 208.800 ;
        RECT 146.200 208.200 146.500 208.800 ;
        RECT 211.800 208.200 212.100 208.800 ;
        RECT 127.800 208.100 128.200 208.200 ;
        RECT 119.000 207.800 128.200 208.100 ;
        RECT 136.600 208.100 137.000 208.200 ;
        RECT 141.400 208.100 141.800 208.200 ;
        RECT 136.600 207.800 141.800 208.100 ;
        RECT 146.200 208.100 146.600 208.200 ;
        RECT 147.800 208.100 148.200 208.200 ;
        RECT 146.200 207.800 148.200 208.100 ;
        RECT 154.200 208.100 154.600 208.200 ;
        RECT 158.200 208.100 158.600 208.200 ;
        RECT 183.000 208.100 183.400 208.200 ;
        RECT 191.000 208.100 191.400 208.200 ;
        RECT 154.200 207.800 182.500 208.100 ;
        RECT 183.000 207.800 191.400 208.100 ;
        RECT 211.800 207.800 212.200 208.200 ;
        RECT 221.400 208.100 221.800 208.200 ;
        RECT 228.600 208.100 229.000 208.200 ;
        RECT 221.400 207.800 229.000 208.100 ;
        RECT 238.200 207.800 238.600 208.200 ;
        RECT 10.200 207.100 10.600 207.200 ;
        RECT 14.200 207.100 14.600 207.200 ;
        RECT 10.200 206.800 14.600 207.100 ;
        RECT 34.200 207.100 34.500 207.800 ;
        RECT 76.600 207.100 77.000 207.200 ;
        RECT 78.200 207.100 78.600 207.200 ;
        RECT 34.200 206.800 78.600 207.100 ;
        RECT 79.800 207.100 80.200 207.200 ;
        RECT 107.000 207.100 107.400 207.200 ;
        RECT 162.200 207.100 162.600 207.200 ;
        RECT 163.800 207.100 164.200 207.200 ;
        RECT 171.000 207.100 171.400 207.200 ;
        RECT 79.800 206.800 162.600 207.100 ;
        RECT 163.000 206.800 171.400 207.100 ;
        RECT 182.200 207.100 182.500 207.800 ;
        RECT 199.000 207.100 199.400 207.200 ;
        RECT 223.000 207.100 223.400 207.200 ;
        RECT 227.800 207.100 228.200 207.200 ;
        RECT 182.200 206.800 228.200 207.100 ;
        RECT 229.400 207.100 229.800 207.200 ;
        RECT 230.200 207.100 230.600 207.200 ;
        RECT 229.400 206.800 230.600 207.100 ;
        RECT 238.200 207.100 238.500 207.800 ;
        RECT 255.800 207.100 256.200 207.200 ;
        RECT 238.200 206.800 256.200 207.100 ;
        RECT 5.400 206.100 5.800 206.200 ;
        RECT 11.800 206.100 12.200 206.200 ;
        RECT 5.400 205.800 12.200 206.100 ;
        RECT 16.600 206.100 17.000 206.200 ;
        RECT 27.000 206.100 27.400 206.200 ;
        RECT 16.600 205.800 27.400 206.100 ;
        RECT 31.800 206.100 32.200 206.200 ;
        RECT 40.600 206.100 41.000 206.200 ;
        RECT 43.800 206.100 44.200 206.200 ;
        RECT 31.800 205.800 44.200 206.100 ;
        RECT 45.400 206.100 45.800 206.200 ;
        RECT 49.400 206.100 49.800 206.200 ;
        RECT 45.400 205.800 49.800 206.100 ;
        RECT 56.600 206.100 57.000 206.200 ;
        RECT 65.400 206.100 65.800 206.200 ;
        RECT 56.600 205.800 65.800 206.100 ;
        RECT 67.800 206.100 68.200 206.200 ;
        RECT 78.200 206.100 78.600 206.200 ;
        RECT 79.000 206.100 79.400 206.200 ;
        RECT 67.800 205.800 79.400 206.100 ;
        RECT 85.400 206.100 85.800 206.200 ;
        RECT 90.200 206.100 90.600 206.200 ;
        RECT 85.400 205.800 90.600 206.100 ;
        RECT 92.600 206.100 93.000 206.200 ;
        RECT 112.600 206.100 113.000 206.200 ;
        RECT 92.600 205.800 113.000 206.100 ;
        RECT 116.600 205.800 117.000 206.200 ;
        RECT 117.400 206.100 117.800 206.200 ;
        RECT 146.200 206.100 146.600 206.200 ;
        RECT 180.600 206.100 181.000 206.200 ;
        RECT 184.600 206.100 185.000 206.200 ;
        RECT 117.400 205.800 164.100 206.100 ;
        RECT 180.600 205.800 185.000 206.100 ;
        RECT 200.600 205.800 201.000 206.200 ;
        RECT 202.200 206.100 202.600 206.200 ;
        RECT 205.400 206.100 205.800 206.200 ;
        RECT 202.200 205.800 205.800 206.100 ;
        RECT 211.800 206.100 212.200 206.200 ;
        RECT 214.200 206.100 214.600 206.200 ;
        RECT 215.800 206.100 216.200 206.200 ;
        RECT 217.400 206.100 217.800 206.200 ;
        RECT 211.800 205.800 217.800 206.100 ;
        RECT 218.200 206.100 218.600 206.200 ;
        RECT 221.400 206.100 221.800 206.200 ;
        RECT 218.200 205.800 221.800 206.100 ;
        RECT 223.800 206.100 224.200 206.200 ;
        RECT 226.200 206.100 226.600 206.200 ;
        RECT 223.800 205.800 226.600 206.100 ;
        RECT 227.000 206.100 227.400 206.200 ;
        RECT 234.200 206.100 234.600 206.200 ;
        RECT 227.000 205.800 234.600 206.100 ;
        RECT 243.800 206.100 244.200 206.200 ;
        RECT 251.000 206.100 251.400 206.200 ;
        RECT 243.800 205.800 251.400 206.100 ;
        RECT 116.600 205.200 116.900 205.800 ;
        RECT 8.600 205.100 9.000 205.200 ;
        RECT 32.600 205.100 33.000 205.200 ;
        RECT 8.600 204.800 33.000 205.100 ;
        RECT 33.400 205.100 33.800 205.200 ;
        RECT 47.800 205.100 48.200 205.200 ;
        RECT 93.400 205.100 93.800 205.200 ;
        RECT 33.400 204.800 93.800 205.100 ;
        RECT 116.600 205.100 117.000 205.200 ;
        RECT 119.000 205.100 119.400 205.200 ;
        RECT 116.600 204.800 119.400 205.100 ;
        RECT 142.200 205.100 142.600 205.200 ;
        RECT 144.600 205.100 145.000 205.200 ;
        RECT 160.600 205.100 161.000 205.200 ;
        RECT 163.000 205.100 163.400 205.200 ;
        RECT 142.200 204.800 145.000 205.100 ;
        RECT 153.400 204.800 155.300 205.100 ;
        RECT 160.600 204.800 163.400 205.100 ;
        RECT 163.800 205.100 164.100 205.800 ;
        RECT 200.600 205.200 200.900 205.800 ;
        RECT 200.600 205.100 201.000 205.200 ;
        RECT 163.800 204.800 201.000 205.100 ;
        RECT 210.200 205.100 210.600 205.200 ;
        RECT 212.600 205.100 213.000 205.200 ;
        RECT 239.800 205.100 240.200 205.200 ;
        RECT 210.200 204.800 240.200 205.100 ;
        RECT 144.600 204.200 144.900 204.800 ;
        RECT 153.400 204.200 153.700 204.800 ;
        RECT 155.000 204.200 155.300 204.800 ;
        RECT 163.000 204.200 163.300 204.800 ;
        RECT 13.400 204.100 13.800 204.200 ;
        RECT 39.000 204.100 39.400 204.200 ;
        RECT 13.400 203.800 39.400 204.100 ;
        RECT 86.200 204.100 86.600 204.200 ;
        RECT 90.200 204.100 90.600 204.200 ;
        RECT 86.200 203.800 90.600 204.100 ;
        RECT 135.000 204.100 135.400 204.200 ;
        RECT 135.000 203.800 142.500 204.100 ;
        RECT 144.600 203.800 145.000 204.200 ;
        RECT 153.400 203.800 153.800 204.200 ;
        RECT 155.000 203.800 155.400 204.200 ;
        RECT 163.000 203.800 163.400 204.200 ;
        RECT 184.600 204.100 185.000 204.200 ;
        RECT 190.200 204.100 190.600 204.200 ;
        RECT 184.600 203.800 190.600 204.100 ;
        RECT 142.200 203.200 142.500 203.800 ;
        RECT 17.400 203.100 17.800 203.200 ;
        RECT 21.400 203.100 21.800 203.200 ;
        RECT 69.400 203.100 69.800 203.200 ;
        RECT 111.800 203.100 112.200 203.200 ;
        RECT 17.400 202.800 112.200 203.100 ;
        RECT 142.200 202.800 142.600 203.200 ;
        RECT 154.200 203.100 154.600 203.200 ;
        RECT 199.000 203.100 199.400 203.200 ;
        RECT 224.600 203.100 225.000 203.200 ;
        RECT 231.000 203.100 231.400 203.200 ;
        RECT 154.200 202.800 231.400 203.100 ;
        RECT 154.200 202.200 154.500 202.800 ;
        RECT 31.000 202.100 31.400 202.200 ;
        RECT 52.600 202.100 53.000 202.200 ;
        RECT 31.000 201.800 53.000 202.100 ;
        RECT 90.200 202.100 90.600 202.200 ;
        RECT 104.600 202.100 105.000 202.200 ;
        RECT 131.800 202.100 132.200 202.200 ;
        RECT 142.200 202.100 142.600 202.200 ;
        RECT 90.200 201.800 142.600 202.100 ;
        RECT 154.200 201.800 154.600 202.200 ;
        RECT 157.400 202.100 157.800 202.200 ;
        RECT 194.200 202.100 194.600 202.200 ;
        RECT 229.400 202.100 229.800 202.200 ;
        RECT 157.400 201.800 229.800 202.100 ;
        RECT 87.000 201.100 87.400 201.200 ;
        RECT 89.400 201.100 89.800 201.200 ;
        RECT 87.000 200.800 89.800 201.100 ;
        RECT 179.000 201.100 179.400 201.200 ;
        RECT 185.400 201.100 185.800 201.200 ;
        RECT 179.000 200.800 185.800 201.100 ;
        RECT 188.600 201.100 189.000 201.200 ;
        RECT 219.000 201.100 219.400 201.200 ;
        RECT 188.600 200.800 219.400 201.100 ;
        RECT 67.000 200.100 67.400 200.200 ;
        RECT 99.800 200.100 100.200 200.200 ;
        RECT 67.000 199.800 100.200 200.100 ;
        RECT 197.400 200.100 197.800 200.200 ;
        RECT 199.000 200.100 199.400 200.200 ;
        RECT 197.400 199.800 199.400 200.100 ;
        RECT 206.200 200.100 206.600 200.200 ;
        RECT 227.000 200.100 227.400 200.200 ;
        RECT 230.200 200.100 230.600 200.200 ;
        RECT 206.200 199.800 230.600 200.100 ;
        RECT 43.800 199.100 44.200 199.200 ;
        RECT 87.800 199.100 88.200 199.200 ;
        RECT 43.800 198.800 88.200 199.100 ;
        RECT 88.600 199.100 89.000 199.200 ;
        RECT 95.000 199.100 95.400 199.200 ;
        RECT 88.600 198.800 95.400 199.100 ;
        RECT 187.000 199.100 187.400 199.200 ;
        RECT 195.000 199.100 195.400 199.200 ;
        RECT 187.000 198.800 195.400 199.100 ;
        RECT 210.200 199.100 210.600 199.200 ;
        RECT 246.200 199.100 246.600 199.200 ;
        RECT 210.200 198.800 246.600 199.100 ;
        RECT 32.600 198.100 33.000 198.200 ;
        RECT 49.400 198.100 49.800 198.200 ;
        RECT 32.600 197.800 49.800 198.100 ;
        RECT 65.400 198.100 65.800 198.200 ;
        RECT 70.200 198.100 70.600 198.200 ;
        RECT 65.400 197.800 70.600 198.100 ;
        RECT 71.800 198.100 72.200 198.200 ;
        RECT 95.000 198.100 95.400 198.200 ;
        RECT 71.800 197.800 95.400 198.100 ;
        RECT 107.800 198.100 108.200 198.200 ;
        RECT 173.400 198.100 173.800 198.200 ;
        RECT 223.800 198.100 224.200 198.200 ;
        RECT 225.400 198.100 225.800 198.200 ;
        RECT 107.800 197.800 225.800 198.100 ;
        RECT 27.000 196.800 27.400 197.200 ;
        RECT 39.000 197.100 39.400 197.200 ;
        RECT 69.400 197.100 69.800 197.200 ;
        RECT 39.000 196.800 69.800 197.100 ;
        RECT 83.800 197.100 84.200 197.200 ;
        RECT 108.600 197.100 109.000 197.200 ;
        RECT 83.800 196.800 109.000 197.100 ;
        RECT 128.600 197.100 129.000 197.200 ;
        RECT 140.600 197.100 141.000 197.200 ;
        RECT 145.400 197.100 145.800 197.200 ;
        RECT 128.600 196.800 145.800 197.100 ;
        RECT 211.800 197.100 212.200 197.200 ;
        RECT 218.200 197.100 218.600 197.200 ;
        RECT 211.800 196.800 218.600 197.100 ;
        RECT 224.600 197.100 225.000 197.200 ;
        RECT 250.200 197.100 250.600 197.200 ;
        RECT 255.800 197.100 256.200 197.200 ;
        RECT 224.600 196.800 256.200 197.100 ;
        RECT 19.000 196.100 19.400 196.200 ;
        RECT 26.200 196.100 26.600 196.200 ;
        RECT 19.000 195.800 26.600 196.100 ;
        RECT 27.000 196.100 27.300 196.800 ;
        RECT 34.200 196.100 34.600 196.200 ;
        RECT 27.000 195.800 34.600 196.100 ;
        RECT 57.400 195.800 57.800 196.200 ;
        RECT 68.600 195.800 69.000 196.200 ;
        RECT 84.600 196.100 85.000 196.200 ;
        RECT 85.400 196.100 85.800 196.200 ;
        RECT 91.800 196.100 92.200 196.200 ;
        RECT 84.600 195.800 92.200 196.100 ;
        RECT 93.400 196.100 93.800 196.200 ;
        RECT 112.600 196.100 113.000 196.200 ;
        RECT 93.400 195.800 113.000 196.100 ;
        RECT 115.000 196.100 115.400 196.200 ;
        RECT 121.400 196.100 121.800 196.200 ;
        RECT 131.800 196.100 132.200 196.200 ;
        RECT 135.000 196.100 135.400 196.200 ;
        RECT 115.000 195.800 121.800 196.100 ;
        RECT 131.000 195.800 135.400 196.100 ;
        RECT 158.200 196.100 158.600 196.200 ;
        RECT 167.000 196.100 167.400 196.200 ;
        RECT 158.200 195.800 167.400 196.100 ;
        RECT 208.600 195.800 209.000 196.200 ;
        RECT 213.400 196.100 213.800 196.200 ;
        RECT 214.200 196.100 214.600 196.200 ;
        RECT 217.400 196.100 217.800 196.200 ;
        RECT 222.200 196.100 222.600 196.200 ;
        RECT 247.800 196.100 248.200 196.200 ;
        RECT 213.400 195.800 248.200 196.100 ;
        RECT 8.600 194.800 9.000 195.200 ;
        RECT 11.800 195.100 12.200 195.200 ;
        RECT 19.800 195.100 20.200 195.200 ;
        RECT 11.800 194.800 20.200 195.100 ;
        RECT 27.800 194.800 28.200 195.200 ;
        RECT 36.600 195.100 37.000 195.200 ;
        RECT 52.600 195.100 53.000 195.200 ;
        RECT 36.600 194.800 53.000 195.100 ;
        RECT 57.400 195.100 57.700 195.800 ;
        RECT 64.600 195.100 65.000 195.200 ;
        RECT 57.400 194.800 65.000 195.100 ;
        RECT 68.600 195.100 68.900 195.800 ;
        RECT 75.800 195.100 76.200 195.200 ;
        RECT 68.600 194.800 76.200 195.100 ;
        RECT 82.200 195.100 82.600 195.200 ;
        RECT 88.600 195.100 89.000 195.200 ;
        RECT 82.200 194.800 89.000 195.100 ;
        RECT 91.800 195.100 92.200 195.200 ;
        RECT 99.000 195.100 99.400 195.200 ;
        RECT 91.800 194.800 99.400 195.100 ;
        RECT 100.600 194.800 101.000 195.200 ;
        RECT 119.800 195.100 120.200 195.200 ;
        RECT 122.200 195.100 122.600 195.200 ;
        RECT 119.800 194.800 122.600 195.100 ;
        RECT 127.000 195.100 127.400 195.200 ;
        RECT 131.000 195.100 131.400 195.200 ;
        RECT 127.000 194.800 131.400 195.100 ;
        RECT 131.800 194.800 132.200 195.200 ;
        RECT 155.000 195.100 155.400 195.200 ;
        RECT 155.800 195.100 156.200 195.200 ;
        RECT 159.000 195.100 159.400 195.200 ;
        RECT 182.200 195.100 182.600 195.200 ;
        RECT 183.800 195.100 184.200 195.200 ;
        RECT 155.000 194.800 184.200 195.100 ;
        RECT 190.200 195.100 190.600 195.200 ;
        RECT 197.400 195.100 197.800 195.200 ;
        RECT 190.200 194.800 197.800 195.100 ;
        RECT 200.600 195.100 201.000 195.200 ;
        RECT 207.000 195.100 207.400 195.200 ;
        RECT 200.600 194.800 207.400 195.100 ;
        RECT 208.600 195.100 208.900 195.800 ;
        RECT 215.000 195.100 215.400 195.200 ;
        RECT 208.600 194.800 215.400 195.100 ;
        RECT 230.200 195.100 230.600 195.200 ;
        RECT 237.400 195.100 237.800 195.200 ;
        RECT 230.200 194.800 237.800 195.100 ;
        RECT 246.200 195.100 246.600 195.200 ;
        RECT 250.200 195.100 250.600 195.200 ;
        RECT 246.200 194.800 250.600 195.100 ;
        RECT 0.600 194.100 1.000 194.200 ;
        RECT 6.200 194.100 6.600 194.200 ;
        RECT 8.600 194.100 8.900 194.800 ;
        RECT 0.600 193.800 8.900 194.100 ;
        RECT 20.600 194.100 21.000 194.200 ;
        RECT 27.800 194.100 28.100 194.800 ;
        RECT 20.600 193.800 28.100 194.100 ;
        RECT 41.400 194.100 41.800 194.200 ;
        RECT 49.400 194.100 49.800 194.200 ;
        RECT 41.400 193.800 49.800 194.100 ;
        RECT 51.000 194.100 51.400 194.200 ;
        RECT 62.200 194.100 62.600 194.200 ;
        RECT 51.000 193.800 62.600 194.100 ;
        RECT 70.200 194.100 70.600 194.200 ;
        RECT 88.600 194.100 89.000 194.200 ;
        RECT 70.200 193.800 89.000 194.100 ;
        RECT 100.600 194.100 100.900 194.800 ;
        RECT 131.000 194.200 131.300 194.800 ;
        RECT 130.200 194.100 130.600 194.200 ;
        RECT 100.600 193.800 130.600 194.100 ;
        RECT 131.000 193.800 131.400 194.200 ;
        RECT 131.800 194.100 132.100 194.800 ;
        RECT 136.600 194.100 137.000 194.200 ;
        RECT 153.400 194.100 153.800 194.200 ;
        RECT 159.800 194.100 160.200 194.200 ;
        RECT 131.800 193.800 160.200 194.100 ;
        RECT 166.200 194.100 166.600 194.200 ;
        RECT 179.800 194.100 180.200 194.200 ;
        RECT 166.200 193.800 180.200 194.100 ;
        RECT 203.800 194.100 204.200 194.200 ;
        RECT 215.800 194.100 216.200 194.200 ;
        RECT 219.000 194.100 219.400 194.200 ;
        RECT 203.800 193.800 219.400 194.100 ;
        RECT 227.000 194.100 227.400 194.200 ;
        RECT 243.000 194.100 243.400 194.200 ;
        RECT 227.000 193.800 243.400 194.100 ;
        RECT 245.400 194.100 245.800 194.200 ;
        RECT 257.400 194.100 257.800 194.200 ;
        RECT 245.400 193.800 257.800 194.100 ;
        RECT 19.000 193.100 19.400 193.200 ;
        RECT 21.400 193.100 21.800 193.200 ;
        RECT 19.000 192.800 21.800 193.100 ;
        RECT 23.000 193.100 23.400 193.200 ;
        RECT 28.600 193.100 29.000 193.200 ;
        RECT 23.000 192.800 29.000 193.100 ;
        RECT 43.800 193.100 44.200 193.200 ;
        RECT 63.000 193.100 63.400 193.200 ;
        RECT 67.000 193.100 67.400 193.200 ;
        RECT 43.800 192.800 67.400 193.100 ;
        RECT 79.800 193.100 80.200 193.200 ;
        RECT 80.600 193.100 81.000 193.200 ;
        RECT 79.800 192.800 81.000 193.100 ;
        RECT 130.200 193.100 130.600 193.200 ;
        RECT 132.600 193.100 133.000 193.200 ;
        RECT 155.800 193.100 156.200 193.200 ;
        RECT 130.200 192.800 156.200 193.100 ;
        RECT 171.800 193.100 172.200 193.200 ;
        RECT 179.000 193.100 179.400 193.200 ;
        RECT 171.800 192.800 179.400 193.100 ;
        RECT 196.600 193.100 197.000 193.200 ;
        RECT 202.200 193.100 202.600 193.200 ;
        RECT 196.600 192.800 202.600 193.100 ;
        RECT 243.000 193.100 243.400 193.200 ;
        RECT 261.400 193.100 261.800 193.200 ;
        RECT 243.000 192.800 261.800 193.100 ;
        RECT 19.000 192.100 19.400 192.200 ;
        RECT 23.000 192.100 23.300 192.800 ;
        RECT 19.000 191.800 23.300 192.100 ;
        RECT 24.600 192.100 25.000 192.200 ;
        RECT 27.000 192.100 27.400 192.200 ;
        RECT 34.200 192.100 34.600 192.200 ;
        RECT 24.600 191.800 34.600 192.100 ;
        RECT 53.400 192.100 53.800 192.200 ;
        RECT 65.400 192.100 65.800 192.200 ;
        RECT 53.400 191.800 65.800 192.100 ;
        RECT 66.200 192.100 66.600 192.200 ;
        RECT 87.800 192.100 88.200 192.200 ;
        RECT 66.200 191.800 88.200 192.100 ;
        RECT 103.000 192.100 103.400 192.200 ;
        RECT 107.800 192.100 108.200 192.200 ;
        RECT 118.200 192.100 118.600 192.200 ;
        RECT 103.000 191.800 118.600 192.100 ;
        RECT 169.400 192.100 169.800 192.200 ;
        RECT 171.800 192.100 172.100 192.800 ;
        RECT 169.400 191.800 172.100 192.100 ;
        RECT 201.400 192.100 201.800 192.200 ;
        RECT 203.000 192.100 203.400 192.200 ;
        RECT 211.800 192.100 212.200 192.200 ;
        RECT 201.400 191.800 212.200 192.100 ;
        RECT 240.600 192.100 241.000 192.200 ;
        RECT 253.400 192.100 253.800 192.200 ;
        RECT 240.600 191.800 253.800 192.100 ;
        RECT 261.400 192.100 261.800 192.200 ;
        RECT 264.600 192.100 265.000 192.200 ;
        RECT 261.400 191.800 265.000 192.100 ;
        RECT 6.200 191.100 6.600 191.200 ;
        RECT 39.000 191.100 39.400 191.200 ;
        RECT 6.200 190.800 39.400 191.100 ;
        RECT 53.400 191.100 53.800 191.200 ;
        RECT 65.400 191.100 65.800 191.200 ;
        RECT 71.000 191.100 71.400 191.200 ;
        RECT 53.400 190.800 71.400 191.100 ;
        RECT 83.000 191.100 83.400 191.200 ;
        RECT 84.600 191.100 85.000 191.200 ;
        RECT 83.000 190.800 85.000 191.100 ;
        RECT 159.000 191.100 159.400 191.200 ;
        RECT 164.600 191.100 165.000 191.200 ;
        RECT 159.000 190.800 165.000 191.100 ;
        RECT 225.400 191.100 225.800 191.200 ;
        RECT 238.200 191.100 238.600 191.200 ;
        RECT 243.000 191.100 243.400 191.200 ;
        RECT 225.400 190.800 243.400 191.100 ;
        RECT 13.400 190.100 13.800 190.200 ;
        RECT 22.200 190.100 22.600 190.200 ;
        RECT 27.000 190.100 27.400 190.200 ;
        RECT 36.600 190.100 37.000 190.200 ;
        RECT 42.200 190.100 42.600 190.200 ;
        RECT 104.600 190.100 105.000 190.200 ;
        RECT 13.400 189.800 105.000 190.100 ;
        RECT 126.200 190.100 126.600 190.200 ;
        RECT 167.000 190.100 167.400 190.200 ;
        RECT 126.200 189.800 167.400 190.100 ;
        RECT 185.400 190.100 185.800 190.200 ;
        RECT 187.000 190.100 187.400 190.200 ;
        RECT 192.600 190.100 193.000 190.200 ;
        RECT 185.400 189.800 193.000 190.100 ;
        RECT 232.600 190.100 233.000 190.200 ;
        RECT 251.000 190.100 251.400 190.200 ;
        RECT 232.600 189.800 251.400 190.100 ;
        RECT 26.200 189.100 26.600 189.200 ;
        RECT 31.800 189.100 32.200 189.200 ;
        RECT 43.000 189.100 43.400 189.200 ;
        RECT 26.200 188.800 43.400 189.100 ;
        RECT 59.000 189.100 59.400 189.200 ;
        RECT 61.400 189.100 61.800 189.200 ;
        RECT 59.000 188.800 61.800 189.100 ;
        RECT 73.400 189.100 73.800 189.200 ;
        RECT 82.200 189.100 82.600 189.200 ;
        RECT 84.600 189.100 85.000 189.200 ;
        RECT 73.400 188.800 85.000 189.100 ;
        RECT 100.600 189.100 101.000 189.200 ;
        RECT 107.000 189.100 107.400 189.200 ;
        RECT 115.800 189.100 116.200 189.200 ;
        RECT 100.600 188.800 116.200 189.100 ;
        RECT 131.000 189.100 131.400 189.200 ;
        RECT 146.200 189.100 146.600 189.200 ;
        RECT 131.000 188.800 146.600 189.100 ;
        RECT 173.400 189.100 173.800 189.200 ;
        RECT 175.000 189.100 175.400 189.200 ;
        RECT 234.200 189.100 234.600 189.200 ;
        RECT 173.400 188.800 234.600 189.100 ;
        RECT 19.800 188.100 20.200 188.200 ;
        RECT 28.600 188.100 29.000 188.200 ;
        RECT 19.800 187.800 29.000 188.100 ;
        RECT 67.000 188.100 67.400 188.200 ;
        RECT 69.400 188.100 69.800 188.200 ;
        RECT 67.000 187.800 69.800 188.100 ;
        RECT 93.400 188.100 93.800 188.200 ;
        RECT 110.200 188.100 110.600 188.200 ;
        RECT 120.600 188.100 121.000 188.200 ;
        RECT 93.400 187.800 121.000 188.100 ;
        RECT 130.200 188.100 130.600 188.200 ;
        RECT 131.000 188.100 131.300 188.800 ;
        RECT 130.200 187.800 131.300 188.100 ;
        RECT 137.400 188.100 137.800 188.200 ;
        RECT 143.000 188.100 143.400 188.200 ;
        RECT 137.400 187.800 143.400 188.100 ;
        RECT 163.800 188.100 164.200 188.200 ;
        RECT 165.400 188.100 165.800 188.200 ;
        RECT 171.000 188.100 171.400 188.200 ;
        RECT 163.800 187.800 171.400 188.100 ;
        RECT 179.000 188.100 179.400 188.200 ;
        RECT 179.800 188.100 180.200 188.200 ;
        RECT 179.000 187.800 180.200 188.100 ;
        RECT 206.200 188.100 206.600 188.200 ;
        RECT 233.400 188.100 233.800 188.200 ;
        RECT 206.200 187.800 233.800 188.100 ;
        RECT 251.800 187.800 252.200 188.200 ;
        RECT 14.200 187.100 14.600 187.200 ;
        RECT 38.200 187.100 38.600 187.200 ;
        RECT 14.200 186.800 38.600 187.100 ;
        RECT 40.600 187.100 41.000 187.200 ;
        RECT 43.800 187.100 44.200 187.200 ;
        RECT 40.600 186.800 44.200 187.100 ;
        RECT 50.200 186.800 50.600 187.200 ;
        RECT 55.800 186.800 56.200 187.200 ;
        RECT 60.600 187.100 61.000 187.200 ;
        RECT 60.600 186.800 84.100 187.100 ;
        RECT 10.200 186.100 10.600 186.200 ;
        RECT 11.800 186.100 12.200 186.200 ;
        RECT 23.000 186.100 23.400 186.200 ;
        RECT 10.200 185.800 12.200 186.100 ;
        RECT 15.800 185.800 23.400 186.100 ;
        RECT 29.400 186.100 29.800 186.200 ;
        RECT 35.000 186.100 35.400 186.200 ;
        RECT 35.800 186.100 36.200 186.200 ;
        RECT 29.400 185.800 33.700 186.100 ;
        RECT 35.000 185.800 36.200 186.100 ;
        RECT 41.400 186.100 41.800 186.200 ;
        RECT 47.000 186.100 47.400 186.200 ;
        RECT 50.200 186.100 50.500 186.800 ;
        RECT 41.400 185.800 42.500 186.100 ;
        RECT 47.000 185.800 50.500 186.100 ;
        RECT 55.800 186.100 56.100 186.800 ;
        RECT 56.600 186.100 57.000 186.200 ;
        RECT 55.800 185.800 57.000 186.100 ;
        RECT 59.800 186.100 60.200 186.200 ;
        RECT 63.800 186.100 64.200 186.200 ;
        RECT 59.800 185.800 64.200 186.100 ;
        RECT 68.600 186.100 69.000 186.200 ;
        RECT 70.200 186.100 70.600 186.200 ;
        RECT 68.600 185.800 70.600 186.100 ;
        RECT 71.800 186.100 72.200 186.200 ;
        RECT 83.800 186.100 84.100 186.800 ;
        RECT 98.200 186.800 98.600 187.200 ;
        RECT 112.600 187.100 113.000 187.200 ;
        RECT 118.200 187.100 118.600 187.200 ;
        RECT 112.600 186.800 118.600 187.100 ;
        RECT 120.600 187.100 120.900 187.800 ;
        RECT 123.000 187.100 123.400 187.200 ;
        RECT 120.600 186.800 123.400 187.100 ;
        RECT 139.800 186.800 140.200 187.200 ;
        RECT 159.800 187.100 160.200 187.200 ;
        RECT 165.400 187.100 165.800 187.200 ;
        RECT 159.800 186.800 165.800 187.100 ;
        RECT 167.000 187.100 167.400 187.200 ;
        RECT 185.400 187.100 185.800 187.200 ;
        RECT 199.800 187.100 200.200 187.200 ;
        RECT 167.000 186.800 200.200 187.100 ;
        RECT 200.600 187.100 201.000 187.200 ;
        RECT 203.800 187.100 204.200 187.200 ;
        RECT 200.600 186.800 204.200 187.100 ;
        RECT 215.000 186.800 215.400 187.200 ;
        RECT 229.400 187.100 229.800 187.200 ;
        RECT 231.800 187.100 232.200 187.200 ;
        RECT 229.400 186.800 232.200 187.100 ;
        RECT 236.600 187.100 237.000 187.200 ;
        RECT 238.200 187.100 238.600 187.200 ;
        RECT 243.800 187.100 244.200 187.200 ;
        RECT 236.600 186.800 244.200 187.100 ;
        RECT 251.800 187.100 252.100 187.800 ;
        RECT 259.800 187.100 260.200 187.200 ;
        RECT 251.800 186.800 260.200 187.100 ;
        RECT 91.000 186.100 91.400 186.200 ;
        RECT 71.800 185.800 76.900 186.100 ;
        RECT 15.800 185.200 16.100 185.800 ;
        RECT 33.400 185.200 33.700 185.800 ;
        RECT 42.200 185.200 42.500 185.800 ;
        RECT 68.600 185.200 68.900 185.800 ;
        RECT 76.600 185.200 76.900 185.800 ;
        RECT 83.800 185.800 91.400 186.100 ;
        RECT 93.400 186.100 93.800 186.200 ;
        RECT 98.200 186.100 98.500 186.800 ;
        RECT 102.200 186.100 102.600 186.200 ;
        RECT 93.400 185.800 94.500 186.100 ;
        RECT 98.200 185.800 102.600 186.100 ;
        RECT 114.200 186.100 114.600 186.200 ;
        RECT 121.400 186.100 121.800 186.200 ;
        RECT 126.200 186.100 126.600 186.200 ;
        RECT 114.200 185.800 126.600 186.100 ;
        RECT 132.600 186.100 133.000 186.200 ;
        RECT 139.800 186.100 140.100 186.800 ;
        RECT 132.600 185.800 140.100 186.100 ;
        RECT 147.800 186.100 148.200 186.200 ;
        RECT 151.800 186.100 152.200 186.200 ;
        RECT 147.800 185.800 152.200 186.100 ;
        RECT 162.200 186.100 162.600 186.200 ;
        RECT 202.200 186.100 202.600 186.200 ;
        RECT 162.200 185.800 202.600 186.100 ;
        RECT 213.400 186.100 213.800 186.200 ;
        RECT 215.000 186.100 215.300 186.800 ;
        RECT 213.400 185.800 215.300 186.100 ;
        RECT 218.200 186.100 218.600 186.200 ;
        RECT 221.400 186.100 221.800 186.200 ;
        RECT 234.200 186.100 234.600 186.200 ;
        RECT 218.200 185.800 221.800 186.100 ;
        RECT 233.400 185.800 234.600 186.100 ;
        RECT 237.400 185.800 237.800 186.200 ;
        RECT 239.800 186.100 240.200 186.200 ;
        RECT 243.800 186.100 244.200 186.200 ;
        RECT 247.000 186.100 247.400 186.200 ;
        RECT 239.800 185.800 247.400 186.100 ;
        RECT 83.800 185.200 84.100 185.800 ;
        RECT 94.200 185.200 94.500 185.800 ;
        RECT 233.400 185.200 233.700 185.800 ;
        RECT 237.400 185.200 237.700 185.800 ;
        RECT 3.800 185.100 4.200 185.200 ;
        RECT 11.800 185.100 12.200 185.200 ;
        RECT 3.800 184.800 12.200 185.100 ;
        RECT 15.800 184.800 16.200 185.200 ;
        RECT 27.000 185.100 27.400 185.200 ;
        RECT 32.600 185.100 33.000 185.200 ;
        RECT 27.000 184.800 33.000 185.100 ;
        RECT 33.400 184.800 33.800 185.200 ;
        RECT 42.200 184.800 42.600 185.200 ;
        RECT 55.000 185.100 55.400 185.200 ;
        RECT 56.600 185.100 57.000 185.200 ;
        RECT 55.000 184.800 57.000 185.100 ;
        RECT 64.600 185.100 65.000 185.200 ;
        RECT 66.200 185.100 66.600 185.200 ;
        RECT 64.600 184.800 66.600 185.100 ;
        RECT 68.600 184.800 69.000 185.200 ;
        RECT 76.600 184.800 77.000 185.200 ;
        RECT 83.800 184.800 84.200 185.200 ;
        RECT 94.200 184.800 94.600 185.200 ;
        RECT 114.200 185.100 114.600 185.200 ;
        RECT 118.200 185.100 118.600 185.200 ;
        RECT 119.800 185.100 120.200 185.200 ;
        RECT 114.200 184.800 120.200 185.100 ;
        RECT 122.200 185.100 122.600 185.200 ;
        RECT 139.800 185.100 140.200 185.200 ;
        RECT 122.200 184.800 140.200 185.100 ;
        RECT 142.200 185.100 142.600 185.200 ;
        RECT 188.600 185.100 189.000 185.200 ;
        RECT 142.200 184.800 189.000 185.100 ;
        RECT 198.200 185.100 198.600 185.200 ;
        RECT 203.000 185.100 203.400 185.200 ;
        RECT 203.800 185.100 204.200 185.200 ;
        RECT 198.200 184.800 204.200 185.100 ;
        RECT 233.400 184.800 233.800 185.200 ;
        RECT 237.400 184.800 237.800 185.200 ;
        RECT 243.000 185.100 243.400 185.200 ;
        RECT 249.400 185.100 249.800 185.200 ;
        RECT 242.200 184.800 249.800 185.100 ;
        RECT 36.600 184.100 37.000 184.200 ;
        RECT 41.400 184.100 41.800 184.200 ;
        RECT 42.200 184.100 42.600 184.200 ;
        RECT 36.600 183.800 42.600 184.100 ;
        RECT 48.600 184.100 49.000 184.200 ;
        RECT 51.800 184.100 52.200 184.200 ;
        RECT 61.400 184.100 61.800 184.200 ;
        RECT 48.600 183.800 61.800 184.100 ;
        RECT 93.400 184.100 93.800 184.200 ;
        RECT 109.400 184.100 109.800 184.200 ;
        RECT 93.400 183.800 109.800 184.100 ;
        RECT 228.600 184.100 229.000 184.200 ;
        RECT 260.600 184.100 261.000 184.200 ;
        RECT 262.200 184.100 262.600 184.200 ;
        RECT 228.600 183.800 262.600 184.100 ;
        RECT 67.800 183.100 68.200 183.200 ;
        RECT 97.400 183.100 97.800 183.200 ;
        RECT 67.800 182.800 97.800 183.100 ;
        RECT 139.000 183.100 139.400 183.200 ;
        RECT 141.400 183.100 141.800 183.200 ;
        RECT 139.000 182.800 141.800 183.100 ;
        RECT 151.000 183.100 151.400 183.200 ;
        RECT 151.800 183.100 152.200 183.200 ;
        RECT 151.000 182.800 152.200 183.100 ;
        RECT 171.800 183.100 172.200 183.200 ;
        RECT 241.400 183.100 241.800 183.200 ;
        RECT 171.800 182.800 241.800 183.100 ;
        RECT 141.400 182.200 141.700 182.800 ;
        RECT 49.400 182.100 49.800 182.200 ;
        RECT 79.000 182.100 79.400 182.200 ;
        RECT 49.400 181.800 79.400 182.100 ;
        RECT 141.400 181.800 141.800 182.200 ;
        RECT 142.200 182.100 142.600 182.200 ;
        RECT 175.800 182.100 176.200 182.200 ;
        RECT 209.400 182.100 209.800 182.200 ;
        RECT 235.000 182.100 235.400 182.200 ;
        RECT 142.200 181.800 235.400 182.100 ;
        RECT 71.800 181.100 72.200 181.200 ;
        RECT 104.600 181.100 105.000 181.200 ;
        RECT 142.200 181.100 142.600 181.200 ;
        RECT 71.800 180.800 142.600 181.100 ;
        RECT 165.400 181.100 165.800 181.200 ;
        RECT 176.600 181.100 177.000 181.200 ;
        RECT 165.400 180.800 177.000 181.100 ;
        RECT 181.400 181.100 181.800 181.200 ;
        RECT 189.400 181.100 189.800 181.200 ;
        RECT 181.400 180.800 189.800 181.100 ;
        RECT 195.800 181.100 196.200 181.200 ;
        RECT 213.400 181.100 213.800 181.200 ;
        RECT 195.800 180.800 213.800 181.100 ;
        RECT 234.200 181.100 234.600 181.200 ;
        RECT 237.400 181.100 237.800 181.200 ;
        RECT 234.200 180.800 237.800 181.100 ;
        RECT 85.400 180.100 85.800 180.200 ;
        RECT 88.600 180.100 89.000 180.200 ;
        RECT 90.200 180.100 90.600 180.200 ;
        RECT 85.400 179.800 90.600 180.100 ;
        RECT 184.600 180.100 185.000 180.200 ;
        RECT 246.200 180.100 246.600 180.200 ;
        RECT 249.400 180.100 249.800 180.200 ;
        RECT 184.600 179.800 249.800 180.100 ;
        RECT 56.600 179.100 57.000 179.200 ;
        RECT 99.000 179.100 99.400 179.200 ;
        RECT 56.600 178.800 99.400 179.100 ;
        RECT 162.200 179.100 162.600 179.200 ;
        RECT 185.400 179.100 185.800 179.200 ;
        RECT 162.200 178.800 185.800 179.100 ;
        RECT 197.400 179.100 197.800 179.200 ;
        RECT 214.200 179.100 214.600 179.200 ;
        RECT 197.400 178.800 214.600 179.100 ;
        RECT 219.000 179.100 219.400 179.200 ;
        RECT 230.200 179.100 230.600 179.200 ;
        RECT 219.000 178.800 230.600 179.100 ;
        RECT 197.400 178.200 197.700 178.800 ;
        RECT 21.400 178.100 21.800 178.200 ;
        RECT 25.400 178.100 25.800 178.200 ;
        RECT 21.400 177.800 25.800 178.100 ;
        RECT 31.000 178.100 31.400 178.200 ;
        RECT 43.000 178.100 43.400 178.200 ;
        RECT 31.000 177.800 43.400 178.100 ;
        RECT 58.200 178.100 58.600 178.200 ;
        RECT 95.800 178.100 96.200 178.200 ;
        RECT 58.200 177.800 96.200 178.100 ;
        RECT 127.000 178.100 127.400 178.200 ;
        RECT 133.400 178.100 133.800 178.200 ;
        RECT 134.200 178.100 134.600 178.200 ;
        RECT 127.000 177.800 134.600 178.100 ;
        RECT 197.400 177.800 197.800 178.200 ;
        RECT 205.400 178.100 205.800 178.200 ;
        RECT 211.000 178.100 211.400 178.200 ;
        RECT 205.400 177.800 211.400 178.100 ;
        RECT 229.400 178.100 229.800 178.200 ;
        RECT 263.800 178.100 264.200 178.200 ;
        RECT 229.400 177.800 264.200 178.100 ;
        RECT 14.200 177.100 14.600 177.200 ;
        RECT 17.400 177.100 17.800 177.200 ;
        RECT 14.200 176.800 17.800 177.100 ;
        RECT 26.200 176.800 26.600 177.200 ;
        RECT 29.400 177.100 29.800 177.200 ;
        RECT 31.000 177.100 31.400 177.200 ;
        RECT 29.400 176.800 31.400 177.100 ;
        RECT 39.000 177.100 39.400 177.200 ;
        RECT 55.800 177.100 56.200 177.200 ;
        RECT 39.000 176.800 56.200 177.100 ;
        RECT 67.000 177.100 67.400 177.200 ;
        RECT 71.000 177.100 71.400 177.200 ;
        RECT 67.000 176.800 71.400 177.100 ;
        RECT 97.400 177.100 97.800 177.200 ;
        RECT 105.400 177.100 105.800 177.200 ;
        RECT 97.400 176.800 105.800 177.100 ;
        RECT 115.000 176.800 115.400 177.200 ;
        RECT 142.200 177.100 142.600 177.200 ;
        RECT 148.600 177.100 149.000 177.200 ;
        RECT 142.200 176.800 149.000 177.100 ;
        RECT 160.600 177.100 161.000 177.200 ;
        RECT 164.600 177.100 165.000 177.200 ;
        RECT 160.600 176.800 165.000 177.100 ;
        RECT 169.400 177.100 169.800 177.200 ;
        RECT 171.000 177.100 171.400 177.200 ;
        RECT 169.400 176.800 171.400 177.100 ;
        RECT 194.200 176.800 194.600 177.200 ;
        RECT 195.000 177.100 195.400 177.200 ;
        RECT 206.200 177.100 206.600 177.200 ;
        RECT 195.000 176.800 206.600 177.100 ;
        RECT 223.800 177.100 224.200 177.200 ;
        RECT 233.400 177.100 233.800 177.200 ;
        RECT 223.800 176.800 233.800 177.100 ;
        RECT 26.200 176.100 26.500 176.800 ;
        RECT 30.200 176.100 30.600 176.200 ;
        RECT 26.200 175.800 30.600 176.100 ;
        RECT 33.400 176.100 33.800 176.200 ;
        RECT 38.200 176.100 38.600 176.200 ;
        RECT 68.600 176.100 69.000 176.200 ;
        RECT 70.200 176.100 70.600 176.200 ;
        RECT 71.000 176.100 71.400 176.200 ;
        RECT 33.400 175.800 71.400 176.100 ;
        RECT 99.800 176.100 100.200 176.200 ;
        RECT 101.400 176.100 101.800 176.200 ;
        RECT 99.800 175.800 101.800 176.100 ;
        RECT 107.000 176.100 107.400 176.200 ;
        RECT 109.400 176.100 109.800 176.200 ;
        RECT 107.000 175.800 109.800 176.100 ;
        RECT 114.200 176.100 114.600 176.200 ;
        RECT 115.000 176.100 115.300 176.800 ;
        RECT 114.200 175.800 115.300 176.100 ;
        RECT 148.600 176.100 149.000 176.200 ;
        RECT 178.200 176.100 178.600 176.200 ;
        RECT 186.200 176.100 186.600 176.200 ;
        RECT 191.800 176.100 192.200 176.200 ;
        RECT 148.600 175.800 192.200 176.100 ;
        RECT 194.200 176.100 194.500 176.800 ;
        RECT 199.000 176.100 199.400 176.200 ;
        RECT 194.200 175.800 199.400 176.100 ;
        RECT 207.000 176.100 207.400 176.200 ;
        RECT 220.600 176.100 221.000 176.200 ;
        RECT 207.000 175.800 221.000 176.100 ;
        RECT 226.200 175.800 226.600 176.200 ;
        RECT 231.800 176.100 232.200 176.200 ;
        RECT 231.000 175.800 232.200 176.100 ;
        RECT 246.200 176.100 246.600 176.200 ;
        RECT 246.200 175.800 248.100 176.100 ;
        RECT 226.200 175.200 226.500 175.800 ;
        RECT 247.800 175.200 248.100 175.800 ;
        RECT 248.600 175.800 249.000 176.200 ;
        RECT 8.600 174.800 9.000 175.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 31.800 175.100 32.200 175.200 ;
        RECT 28.600 174.800 32.200 175.100 ;
        RECT 39.000 175.100 39.400 175.200 ;
        RECT 44.600 175.100 45.000 175.200 ;
        RECT 45.400 175.100 45.800 175.200 ;
        RECT 39.000 174.800 45.800 175.100 ;
        RECT 47.000 174.800 47.400 175.200 ;
        RECT 48.600 175.100 49.000 175.200 ;
        RECT 51.800 175.100 52.200 175.200 ;
        RECT 48.600 174.800 52.200 175.100 ;
        RECT 52.600 175.100 53.000 175.200 ;
        RECT 56.600 175.100 57.000 175.200 ;
        RECT 52.600 174.800 57.000 175.100 ;
        RECT 66.200 175.100 66.600 175.200 ;
        RECT 75.000 175.100 75.400 175.200 ;
        RECT 66.200 174.800 75.400 175.100 ;
        RECT 79.800 174.800 80.200 175.200 ;
        RECT 81.400 175.100 81.800 175.200 ;
        RECT 82.200 175.100 82.600 175.200 ;
        RECT 81.400 174.800 82.600 175.100 ;
        RECT 83.800 175.100 84.200 175.200 ;
        RECT 84.600 175.100 85.000 175.200 ;
        RECT 83.800 174.800 85.000 175.100 ;
        RECT 97.400 175.100 97.800 175.200 ;
        RECT 110.200 175.100 110.600 175.200 ;
        RECT 97.400 174.800 110.600 175.100 ;
        RECT 111.000 175.100 111.400 175.200 ;
        RECT 111.800 175.100 112.200 175.200 ;
        RECT 111.000 174.800 112.200 175.100 ;
        RECT 118.200 175.100 118.600 175.200 ;
        RECT 119.000 175.100 119.400 175.200 ;
        RECT 118.200 174.800 119.400 175.100 ;
        RECT 123.000 175.100 123.400 175.200 ;
        RECT 131.800 175.100 132.200 175.200 ;
        RECT 138.200 175.100 138.600 175.200 ;
        RECT 147.000 175.100 147.400 175.200 ;
        RECT 123.000 174.800 147.400 175.100 ;
        RECT 150.200 175.100 150.600 175.200 ;
        RECT 152.600 175.100 153.000 175.200 ;
        RECT 150.200 174.800 153.000 175.100 ;
        RECT 160.600 175.100 161.000 175.200 ;
        RECT 167.800 175.100 168.200 175.200 ;
        RECT 160.600 174.800 168.200 175.100 ;
        RECT 183.000 175.100 183.400 175.200 ;
        RECT 187.000 175.100 187.400 175.200 ;
        RECT 183.000 174.800 187.400 175.100 ;
        RECT 190.200 174.800 190.600 175.200 ;
        RECT 197.400 174.800 197.800 175.200 ;
        RECT 199.800 175.100 200.200 175.200 ;
        RECT 214.200 175.100 214.600 175.200 ;
        RECT 199.800 174.800 214.600 175.100 ;
        RECT 223.000 174.800 223.400 175.200 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 226.200 174.800 226.600 175.200 ;
        RECT 230.200 175.100 230.600 175.200 ;
        RECT 231.000 175.100 231.400 175.200 ;
        RECT 230.200 174.800 231.400 175.100 ;
        RECT 236.600 175.100 237.000 175.200 ;
        RECT 243.000 175.100 243.400 175.200 ;
        RECT 236.600 174.800 243.400 175.100 ;
        RECT 247.800 174.800 248.200 175.200 ;
        RECT 248.600 175.100 248.900 175.800 ;
        RECT 255.800 175.100 256.200 175.200 ;
        RECT 248.600 174.800 256.200 175.100 ;
        RECT 8.600 174.100 8.900 174.800 ;
        RECT 47.000 174.200 47.300 174.800 ;
        RECT 13.400 174.100 13.800 174.200 ;
        RECT 17.400 174.100 17.800 174.200 ;
        RECT 8.600 173.800 17.800 174.100 ;
        RECT 23.800 174.100 24.200 174.200 ;
        RECT 31.000 174.100 31.400 174.200 ;
        RECT 33.400 174.100 33.800 174.200 ;
        RECT 39.000 174.100 39.400 174.200 ;
        RECT 23.800 173.800 39.400 174.100 ;
        RECT 39.800 174.100 40.200 174.200 ;
        RECT 40.600 174.100 41.000 174.200 ;
        RECT 39.800 173.800 41.000 174.100 ;
        RECT 47.000 173.800 47.400 174.200 ;
        RECT 52.600 174.100 53.000 174.200 ;
        RECT 54.200 174.100 54.600 174.200 ;
        RECT 52.600 173.800 54.600 174.100 ;
        RECT 62.200 174.100 62.600 174.200 ;
        RECT 67.000 174.100 67.400 174.200 ;
        RECT 62.200 173.800 67.400 174.100 ;
        RECT 68.600 174.100 69.000 174.200 ;
        RECT 76.600 174.100 77.000 174.200 ;
        RECT 68.600 173.800 77.000 174.100 ;
        RECT 79.800 174.100 80.100 174.800 ;
        RECT 85.400 174.100 85.800 174.200 ;
        RECT 79.800 173.800 85.800 174.100 ;
        RECT 95.000 174.100 95.400 174.200 ;
        RECT 107.800 174.100 108.200 174.200 ;
        RECT 113.400 174.100 113.800 174.200 ;
        RECT 95.000 173.800 113.800 174.100 ;
        RECT 124.600 174.100 125.000 174.200 ;
        RECT 131.000 174.100 131.400 174.200 ;
        RECT 124.600 173.800 131.400 174.100 ;
        RECT 136.600 174.100 137.000 174.200 ;
        RECT 145.400 174.100 145.800 174.200 ;
        RECT 136.600 173.800 145.800 174.100 ;
        RECT 147.800 174.100 148.200 174.200 ;
        RECT 148.600 174.100 149.000 174.200 ;
        RECT 147.800 173.800 149.000 174.100 ;
        RECT 171.000 174.100 171.400 174.200 ;
        RECT 175.800 174.100 176.200 174.200 ;
        RECT 171.000 173.800 176.200 174.100 ;
        RECT 190.200 174.100 190.500 174.800 ;
        RECT 191.800 174.100 192.200 174.200 ;
        RECT 197.400 174.100 197.700 174.800 ;
        RECT 223.000 174.200 223.300 174.800 ;
        RECT 224.600 174.200 224.900 174.800 ;
        RECT 190.200 173.800 197.700 174.100 ;
        RECT 199.000 174.100 199.400 174.200 ;
        RECT 211.800 174.100 212.200 174.200 ;
        RECT 199.000 173.800 218.500 174.100 ;
        RECT 223.000 173.800 223.400 174.200 ;
        RECT 224.600 173.800 225.000 174.200 ;
        RECT 227.800 174.100 228.200 174.200 ;
        RECT 231.000 174.100 231.400 174.200 ;
        RECT 227.800 173.800 231.400 174.100 ;
        RECT 243.800 174.100 244.200 174.200 ;
        RECT 248.600 174.100 249.000 174.200 ;
        RECT 249.400 174.100 249.800 174.200 ;
        RECT 243.800 173.800 249.800 174.100 ;
        RECT 218.200 173.200 218.500 173.800 ;
        RECT 21.400 173.100 21.800 173.200 ;
        RECT 35.800 173.100 36.200 173.200 ;
        RECT 21.400 172.800 36.200 173.100 ;
        RECT 37.400 173.100 37.800 173.200 ;
        RECT 41.400 173.100 41.800 173.200 ;
        RECT 84.600 173.100 85.000 173.200 ;
        RECT 37.400 172.800 85.000 173.100 ;
        RECT 103.000 173.100 103.400 173.200 ;
        RECT 103.800 173.100 104.200 173.200 ;
        RECT 103.000 172.800 104.200 173.100 ;
        RECT 110.200 173.100 110.600 173.200 ;
        RECT 115.800 173.100 116.200 173.200 ;
        RECT 116.600 173.100 117.000 173.200 ;
        RECT 110.200 172.800 117.000 173.100 ;
        RECT 118.200 173.100 118.600 173.200 ;
        RECT 127.800 173.100 128.200 173.200 ;
        RECT 118.200 172.800 128.200 173.100 ;
        RECT 129.400 173.100 129.800 173.200 ;
        RECT 132.600 173.100 133.000 173.200 ;
        RECT 136.600 173.100 137.000 173.200 ;
        RECT 129.400 172.800 137.000 173.100 ;
        RECT 147.800 173.100 148.200 173.200 ;
        RECT 150.200 173.100 150.600 173.200 ;
        RECT 147.800 172.800 150.600 173.100 ;
        RECT 152.600 173.100 153.000 173.200 ;
        RECT 167.800 173.100 168.200 173.200 ;
        RECT 152.600 172.800 168.200 173.100 ;
        RECT 177.400 173.100 177.800 173.200 ;
        RECT 182.200 173.100 182.600 173.200 ;
        RECT 177.400 172.800 182.600 173.100 ;
        RECT 199.000 173.100 199.400 173.200 ;
        RECT 209.400 173.100 209.800 173.200 ;
        RECT 199.000 172.800 209.800 173.100 ;
        RECT 211.000 173.100 211.400 173.200 ;
        RECT 214.200 173.100 214.600 173.200 ;
        RECT 211.000 172.800 214.600 173.100 ;
        RECT 218.200 172.800 218.600 173.200 ;
        RECT 223.800 173.100 224.200 173.200 ;
        RECT 229.400 173.100 229.800 173.200 ;
        RECT 235.000 173.100 235.400 173.200 ;
        RECT 223.800 172.800 235.400 173.100 ;
        RECT 235.800 172.800 236.200 173.200 ;
        RECT 244.600 172.800 245.000 173.200 ;
        RECT 1.400 172.100 1.800 172.200 ;
        RECT 27.800 172.100 28.200 172.200 ;
        RECT 1.400 171.800 28.200 172.100 ;
        RECT 42.200 172.100 42.600 172.200 ;
        RECT 48.600 172.100 49.000 172.200 ;
        RECT 42.200 171.800 49.000 172.100 ;
        RECT 49.400 172.100 49.800 172.200 ;
        RECT 55.000 172.100 55.400 172.200 ;
        RECT 49.400 171.800 55.400 172.100 ;
        RECT 58.200 172.100 58.600 172.200 ;
        RECT 82.200 172.100 82.600 172.200 ;
        RECT 83.800 172.100 84.200 172.200 ;
        RECT 111.800 172.100 112.200 172.200 ;
        RECT 58.200 171.800 82.600 172.100 ;
        RECT 83.000 171.800 112.200 172.100 ;
        RECT 159.000 172.100 159.400 172.200 ;
        RECT 175.000 172.100 175.400 172.200 ;
        RECT 159.000 171.800 175.400 172.100 ;
        RECT 206.200 172.100 206.600 172.200 ;
        RECT 207.000 172.100 207.400 172.200 ;
        RECT 206.200 171.800 207.400 172.100 ;
        RECT 219.800 172.100 220.200 172.200 ;
        RECT 227.000 172.100 227.400 172.200 ;
        RECT 234.200 172.100 234.600 172.200 ;
        RECT 219.800 171.800 234.600 172.100 ;
        RECT 235.800 172.100 236.100 172.800 ;
        RECT 244.600 172.200 244.900 172.800 ;
        RECT 237.400 172.100 237.800 172.200 ;
        RECT 235.800 171.800 237.800 172.100 ;
        RECT 244.600 171.800 245.000 172.200 ;
        RECT 9.400 171.100 9.800 171.200 ;
        RECT 15.800 171.100 16.200 171.200 ;
        RECT 9.400 170.800 16.200 171.100 ;
        RECT 25.400 171.100 25.800 171.200 ;
        RECT 36.600 171.100 37.000 171.200 ;
        RECT 40.600 171.100 41.000 171.200 ;
        RECT 25.400 170.800 41.000 171.100 ;
        RECT 45.400 171.100 45.800 171.200 ;
        RECT 53.400 171.100 53.800 171.200 ;
        RECT 68.600 171.100 69.000 171.200 ;
        RECT 69.400 171.100 69.800 171.200 ;
        RECT 71.000 171.100 71.400 171.200 ;
        RECT 45.400 170.800 71.400 171.100 ;
        RECT 80.600 171.100 81.000 171.200 ;
        RECT 88.600 171.100 89.000 171.200 ;
        RECT 80.600 170.800 89.000 171.100 ;
        RECT 104.600 170.800 105.000 171.200 ;
        RECT 124.600 171.100 125.000 171.200 ;
        RECT 127.000 171.100 127.400 171.200 ;
        RECT 173.400 171.100 173.800 171.200 ;
        RECT 181.400 171.100 181.800 171.200 ;
        RECT 124.600 170.800 181.800 171.100 ;
        RECT 182.200 171.100 182.600 171.200 ;
        RECT 184.600 171.100 185.000 171.200 ;
        RECT 182.200 170.800 185.000 171.100 ;
        RECT 202.200 170.800 202.600 171.200 ;
        RECT 234.200 171.100 234.500 171.800 ;
        RECT 243.800 171.100 244.200 171.200 ;
        RECT 234.200 170.800 244.200 171.100 ;
        RECT 244.600 171.100 245.000 171.200 ;
        RECT 251.000 171.100 251.400 171.200 ;
        RECT 244.600 170.800 251.400 171.100 ;
        RECT 104.600 170.200 104.900 170.800 ;
        RECT 202.200 170.200 202.500 170.800 ;
        RECT 15.000 170.100 15.400 170.200 ;
        RECT 15.800 170.100 16.200 170.200 ;
        RECT 60.600 170.100 61.000 170.200 ;
        RECT 15.000 169.800 61.000 170.100 ;
        RECT 70.200 169.800 70.600 170.200 ;
        RECT 71.000 170.100 71.400 170.200 ;
        RECT 72.600 170.100 73.000 170.200 ;
        RECT 71.000 169.800 73.000 170.100 ;
        RECT 104.600 169.800 105.000 170.200 ;
        RECT 113.400 170.100 113.800 170.200 ;
        RECT 146.200 170.100 146.600 170.200 ;
        RECT 113.400 169.800 146.600 170.100 ;
        RECT 158.200 170.100 158.600 170.200 ;
        RECT 179.800 170.100 180.200 170.200 ;
        RECT 158.200 169.800 180.200 170.100 ;
        RECT 202.200 169.800 202.600 170.200 ;
        RECT 212.600 170.100 213.000 170.200 ;
        RECT 216.600 170.100 217.000 170.200 ;
        RECT 212.600 169.800 217.000 170.100 ;
        RECT 234.200 170.100 234.600 170.200 ;
        RECT 244.600 170.100 245.000 170.200 ;
        RECT 234.200 169.800 245.000 170.100 ;
        RECT 25.400 169.100 25.800 169.200 ;
        RECT 39.000 169.100 39.400 169.200 ;
        RECT 25.400 168.800 39.400 169.100 ;
        RECT 48.600 169.100 49.000 169.200 ;
        RECT 50.200 169.100 50.600 169.200 ;
        RECT 48.600 168.800 50.600 169.100 ;
        RECT 64.600 169.100 65.000 169.200 ;
        RECT 70.200 169.100 70.500 169.800 ;
        RECT 64.600 168.800 70.500 169.100 ;
        RECT 85.400 169.100 85.800 169.200 ;
        RECT 117.400 169.100 117.800 169.200 ;
        RECT 85.400 168.800 117.800 169.100 ;
        RECT 119.800 169.100 120.200 169.200 ;
        RECT 120.600 169.100 121.000 169.200 ;
        RECT 119.800 168.800 121.000 169.100 ;
        RECT 121.400 168.800 121.800 169.200 ;
        RECT 152.600 169.100 153.000 169.200 ;
        RECT 161.400 169.100 161.800 169.200 ;
        RECT 152.600 168.800 161.800 169.100 ;
        RECT 167.000 169.100 167.400 169.200 ;
        RECT 171.800 169.100 172.200 169.200 ;
        RECT 167.000 168.800 172.200 169.100 ;
        RECT 175.000 169.100 175.400 169.200 ;
        RECT 178.200 169.100 178.600 169.200 ;
        RECT 179.800 169.100 180.200 169.200 ;
        RECT 189.400 169.100 189.800 169.200 ;
        RECT 175.000 168.800 178.600 169.100 ;
        RECT 179.000 168.800 189.800 169.100 ;
        RECT 192.600 169.100 193.000 169.200 ;
        RECT 193.400 169.100 193.800 169.200 ;
        RECT 196.600 169.100 197.000 169.200 ;
        RECT 211.000 169.100 211.400 169.200 ;
        RECT 192.600 168.800 193.800 169.100 ;
        RECT 195.800 168.800 211.400 169.100 ;
        RECT 213.400 169.100 213.800 169.200 ;
        RECT 222.200 169.100 222.600 169.200 ;
        RECT 213.400 168.800 222.600 169.100 ;
        RECT 231.000 169.100 231.400 169.200 ;
        RECT 240.600 169.100 241.000 169.200 ;
        RECT 259.000 169.100 259.400 169.200 ;
        RECT 261.400 169.100 261.800 169.200 ;
        RECT 231.000 168.800 247.300 169.100 ;
        RECT 259.000 168.800 261.800 169.100 ;
        RECT 121.400 168.200 121.700 168.800 ;
        RECT 247.000 168.200 247.300 168.800 ;
        RECT 7.800 168.100 8.200 168.200 ;
        RECT 36.600 168.100 37.000 168.200 ;
        RECT 37.400 168.100 37.800 168.200 ;
        RECT 7.800 167.800 34.500 168.100 ;
        RECT 36.600 167.800 37.800 168.100 ;
        RECT 39.000 168.100 39.400 168.200 ;
        RECT 86.200 168.100 86.600 168.200 ;
        RECT 92.600 168.100 93.000 168.200 ;
        RECT 39.000 167.800 85.700 168.100 ;
        RECT 86.200 167.800 93.000 168.100 ;
        RECT 96.600 168.100 97.000 168.200 ;
        RECT 98.200 168.100 98.600 168.200 ;
        RECT 96.600 167.800 98.600 168.100 ;
        RECT 104.600 168.100 105.000 168.200 ;
        RECT 119.000 168.100 119.400 168.200 ;
        RECT 104.600 167.800 119.400 168.100 ;
        RECT 121.400 167.800 121.800 168.200 ;
        RECT 123.000 167.800 123.400 168.200 ;
        RECT 135.800 168.100 136.200 168.200 ;
        RECT 139.800 168.100 140.200 168.200 ;
        RECT 135.800 167.800 140.200 168.100 ;
        RECT 140.600 167.800 141.000 168.200 ;
        RECT 143.000 167.800 143.400 168.200 ;
        RECT 149.400 168.100 149.800 168.200 ;
        RECT 159.800 168.100 160.200 168.200 ;
        RECT 187.800 168.100 188.200 168.200 ;
        RECT 196.600 168.100 197.000 168.200 ;
        RECT 149.400 167.800 197.000 168.100 ;
        RECT 205.400 168.100 205.800 168.200 ;
        RECT 215.000 168.100 215.400 168.200 ;
        RECT 205.400 167.800 215.400 168.100 ;
        RECT 238.200 167.800 238.600 168.200 ;
        RECT 247.000 167.800 247.400 168.200 ;
        RECT 34.200 167.200 34.500 167.800 ;
        RECT 3.800 167.100 4.200 167.200 ;
        RECT 12.600 167.100 13.000 167.200 ;
        RECT 3.800 166.800 13.000 167.100 ;
        RECT 14.200 167.100 14.600 167.200 ;
        RECT 20.600 167.100 21.000 167.200 ;
        RECT 30.200 167.100 30.600 167.200 ;
        RECT 14.200 166.800 30.600 167.100 ;
        RECT 34.200 166.800 34.600 167.200 ;
        RECT 37.400 167.100 37.700 167.800 ;
        RECT 39.000 167.100 39.400 167.200 ;
        RECT 37.400 166.800 39.400 167.100 ;
        RECT 51.800 167.100 52.200 167.200 ;
        RECT 52.600 167.100 53.000 167.200 ;
        RECT 51.800 166.800 53.000 167.100 ;
        RECT 85.400 167.100 85.700 167.800 ;
        RECT 95.800 167.100 96.200 167.200 ;
        RECT 85.400 166.800 96.200 167.100 ;
        RECT 108.600 167.100 109.000 167.200 ;
        RECT 115.800 167.100 116.200 167.200 ;
        RECT 119.800 167.100 120.200 167.200 ;
        RECT 123.000 167.100 123.300 167.800 ;
        RECT 127.000 167.100 127.400 167.200 ;
        RECT 108.600 166.800 116.900 167.100 ;
        RECT 119.800 166.800 127.400 167.100 ;
        RECT 132.600 167.100 133.000 167.200 ;
        RECT 139.000 167.100 139.400 167.200 ;
        RECT 132.600 166.800 139.400 167.100 ;
        RECT 140.600 167.100 140.900 167.800 ;
        RECT 143.000 167.100 143.300 167.800 ;
        RECT 238.200 167.200 238.500 167.800 ;
        RECT 140.600 166.800 143.300 167.100 ;
        RECT 144.600 167.100 145.000 167.200 ;
        RECT 183.000 167.100 183.400 167.200 ;
        RECT 186.200 167.100 186.600 167.200 ;
        RECT 144.600 166.800 150.500 167.100 ;
        RECT 183.000 166.800 186.600 167.100 ;
        RECT 187.000 166.800 187.400 167.200 ;
        RECT 199.800 167.100 200.200 167.200 ;
        RECT 190.200 166.800 200.200 167.100 ;
        RECT 201.400 166.800 201.800 167.200 ;
        RECT 203.800 167.100 204.200 167.200 ;
        RECT 210.200 167.100 210.600 167.200 ;
        RECT 203.800 166.800 210.600 167.100 ;
        RECT 211.800 166.800 212.200 167.200 ;
        RECT 220.600 166.800 221.000 167.200 ;
        RECT 224.600 166.800 225.000 167.200 ;
        RECT 238.200 166.800 238.600 167.200 ;
        RECT 239.000 167.100 239.400 167.200 ;
        RECT 242.200 167.100 242.600 167.200 ;
        RECT 239.000 166.800 242.600 167.100 ;
        RECT 257.400 167.100 257.800 167.200 ;
        RECT 258.200 167.100 258.600 167.200 ;
        RECT 257.400 166.800 258.600 167.100 ;
        RECT 150.200 166.200 150.500 166.800 ;
        RECT 187.000 166.200 187.300 166.800 ;
        RECT 190.200 166.200 190.500 166.800 ;
        RECT 201.400 166.200 201.700 166.800 ;
        RECT 11.800 166.100 12.200 166.200 ;
        RECT 15.000 166.100 15.400 166.200 ;
        RECT 33.400 166.100 33.800 166.200 ;
        RECT 11.800 165.800 33.800 166.100 ;
        RECT 35.000 166.100 35.400 166.200 ;
        RECT 37.400 166.100 37.800 166.200 ;
        RECT 35.000 165.800 37.800 166.100 ;
        RECT 39.800 166.100 40.200 166.200 ;
        RECT 45.400 166.100 45.800 166.200 ;
        RECT 39.800 165.800 45.800 166.100 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 59.000 166.100 59.400 166.200 ;
        RECT 68.600 166.100 69.000 166.200 ;
        RECT 75.000 166.100 75.400 166.200 ;
        RECT 51.800 165.800 59.400 166.100 ;
        RECT 67.800 165.800 75.400 166.100 ;
        RECT 76.600 166.100 77.000 166.200 ;
        RECT 87.000 166.100 87.400 166.200 ;
        RECT 76.600 165.800 87.400 166.100 ;
        RECT 88.600 165.800 89.000 166.200 ;
        RECT 94.200 166.100 94.600 166.200 ;
        RECT 95.000 166.100 95.400 166.200 ;
        RECT 93.400 165.800 95.400 166.100 ;
        RECT 96.600 166.100 97.000 166.200 ;
        RECT 99.800 166.100 100.200 166.200 ;
        RECT 96.600 165.800 100.200 166.100 ;
        RECT 100.600 166.100 101.000 166.200 ;
        RECT 114.200 166.100 114.600 166.200 ;
        RECT 100.600 165.800 114.600 166.100 ;
        RECT 115.000 166.100 115.400 166.200 ;
        RECT 128.600 166.100 129.000 166.200 ;
        RECT 136.600 166.100 137.000 166.200 ;
        RECT 115.000 165.800 125.700 166.100 ;
        RECT 128.600 165.800 137.000 166.100 ;
        RECT 139.800 166.100 140.200 166.200 ;
        RECT 143.800 166.100 144.200 166.200 ;
        RECT 139.800 165.800 144.200 166.100 ;
        RECT 147.000 166.100 147.400 166.200 ;
        RECT 147.800 166.100 148.200 166.200 ;
        RECT 147.000 165.800 148.200 166.100 ;
        RECT 150.200 165.800 150.600 166.200 ;
        RECT 154.200 165.800 154.600 166.200 ;
        RECT 156.600 166.100 157.000 166.200 ;
        RECT 159.000 166.100 159.400 166.200 ;
        RECT 156.600 165.800 159.400 166.100 ;
        RECT 163.800 165.800 164.200 166.200 ;
        RECT 168.600 165.800 169.000 166.200 ;
        RECT 169.400 165.800 169.800 166.200 ;
        RECT 171.800 165.800 172.200 166.200 ;
        RECT 174.200 165.800 174.600 166.200 ;
        RECT 176.600 165.800 177.000 166.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 189.400 166.100 189.800 166.200 ;
        RECT 190.200 166.100 190.600 166.200 ;
        RECT 189.400 165.800 190.600 166.100 ;
        RECT 194.200 165.800 194.600 166.200 ;
        RECT 195.000 166.100 195.400 166.200 ;
        RECT 195.800 166.100 196.200 166.200 ;
        RECT 195.000 165.800 196.200 166.100 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 211.800 166.100 212.100 166.800 ;
        RECT 216.600 166.100 217.000 166.200 ;
        RECT 211.800 165.800 217.000 166.100 ;
        RECT 217.400 166.100 217.800 166.200 ;
        RECT 220.600 166.100 220.900 166.800 ;
        RECT 217.400 165.800 220.900 166.100 ;
        RECT 224.600 166.100 224.900 166.800 ;
        RECT 231.800 166.100 232.200 166.200 ;
        RECT 224.600 165.800 232.200 166.100 ;
        RECT 235.000 165.800 235.400 166.200 ;
        RECT 243.000 166.100 243.400 166.200 ;
        RECT 251.800 166.100 252.200 166.200 ;
        RECT 242.200 165.800 252.200 166.100 ;
        RECT 6.200 165.100 6.600 165.200 ;
        RECT 16.600 165.100 17.000 165.200 ;
        RECT 6.200 164.800 17.000 165.100 ;
        RECT 20.600 165.100 21.000 165.200 ;
        RECT 27.800 165.100 28.200 165.200 ;
        RECT 20.600 164.800 28.200 165.100 ;
        RECT 34.200 165.100 34.600 165.200 ;
        RECT 35.800 165.100 36.200 165.200 ;
        RECT 38.200 165.100 38.600 165.200 ;
        RECT 67.000 165.100 67.400 165.200 ;
        RECT 69.400 165.100 69.800 165.200 ;
        RECT 34.200 164.800 69.800 165.100 ;
        RECT 76.600 165.100 77.000 165.200 ;
        RECT 84.600 165.100 85.000 165.200 ;
        RECT 76.600 164.800 85.000 165.100 ;
        RECT 88.600 165.100 88.900 165.800 ;
        RECT 99.000 165.200 99.300 165.800 ;
        RECT 125.400 165.200 125.700 165.800 ;
        RECT 88.600 164.800 98.500 165.100 ;
        RECT 99.000 164.800 99.400 165.200 ;
        RECT 120.600 165.100 121.000 165.200 ;
        RECT 122.200 165.100 122.600 165.200 ;
        RECT 120.600 164.800 122.600 165.100 ;
        RECT 125.400 164.800 125.800 165.200 ;
        RECT 143.000 165.100 143.400 165.200 ;
        RECT 148.600 165.100 149.000 165.200 ;
        RECT 143.000 164.800 149.000 165.100 ;
        RECT 151.000 165.100 151.400 165.200 ;
        RECT 152.600 165.100 153.000 165.200 ;
        RECT 151.000 164.800 153.000 165.100 ;
        RECT 154.200 165.100 154.500 165.800 ;
        RECT 163.800 165.200 164.100 165.800 ;
        RECT 168.600 165.200 168.900 165.800 ;
        RECT 169.400 165.200 169.700 165.800 ;
        RECT 171.800 165.200 172.100 165.800 ;
        RECT 159.800 165.100 160.200 165.200 ;
        RECT 154.200 164.800 160.200 165.100 ;
        RECT 163.800 164.800 164.200 165.200 ;
        RECT 168.600 164.800 169.000 165.200 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 171.800 164.800 172.200 165.200 ;
        RECT 174.200 165.100 174.500 165.800 ;
        RECT 176.600 165.200 176.900 165.800 ;
        RECT 194.200 165.200 194.500 165.800 ;
        RECT 235.000 165.200 235.300 165.800 ;
        RECT 175.000 165.100 175.400 165.200 ;
        RECT 174.200 164.800 175.400 165.100 ;
        RECT 176.600 164.800 177.000 165.200 ;
        RECT 177.400 165.100 177.800 165.200 ;
        RECT 180.600 165.100 181.000 165.200 ;
        RECT 177.400 164.800 181.000 165.100 ;
        RECT 194.200 164.800 194.600 165.200 ;
        RECT 195.000 165.100 195.400 165.200 ;
        RECT 200.600 165.100 201.000 165.200 ;
        RECT 206.200 165.100 206.600 165.200 ;
        RECT 195.000 164.800 206.600 165.100 ;
        RECT 223.000 164.800 223.400 165.200 ;
        RECT 235.000 164.800 235.400 165.200 ;
        RECT 243.000 165.100 243.400 165.200 ;
        RECT 245.400 165.100 245.800 165.200 ;
        RECT 246.200 165.100 246.600 165.200 ;
        RECT 243.000 164.800 246.600 165.100 ;
        RECT 97.400 163.800 97.800 164.200 ;
        RECT 98.200 164.100 98.500 164.800 ;
        RECT 99.800 164.100 100.200 164.200 ;
        RECT 98.200 163.800 100.200 164.100 ;
        RECT 129.400 164.100 129.800 164.200 ;
        RECT 142.200 164.100 142.600 164.200 ;
        RECT 129.400 163.800 142.600 164.100 ;
        RECT 147.800 164.100 148.200 164.200 ;
        RECT 195.000 164.100 195.300 164.800 ;
        RECT 147.800 163.800 195.300 164.100 ;
        RECT 199.800 164.100 200.200 164.200 ;
        RECT 211.000 164.100 211.400 164.200 ;
        RECT 199.800 163.800 211.400 164.100 ;
        RECT 211.800 164.100 212.200 164.200 ;
        RECT 223.000 164.100 223.300 164.800 ;
        RECT 211.800 163.800 223.300 164.100 ;
        RECT 229.400 164.100 229.800 164.200 ;
        RECT 256.600 164.100 257.000 164.200 ;
        RECT 257.400 164.100 257.800 164.200 ;
        RECT 229.400 163.800 257.800 164.100 ;
        RECT 76.600 163.100 77.000 163.200 ;
        RECT 95.000 163.100 95.400 163.200 ;
        RECT 76.600 162.800 95.400 163.100 ;
        RECT 97.400 163.100 97.700 163.800 ;
        RECT 143.000 163.100 143.400 163.200 ;
        RECT 97.400 162.800 143.400 163.100 ;
        RECT 144.600 163.100 145.000 163.200 ;
        RECT 153.400 163.100 153.800 163.200 ;
        RECT 144.600 162.800 153.800 163.100 ;
        RECT 162.200 163.100 162.600 163.200 ;
        RECT 166.200 163.100 166.600 163.200 ;
        RECT 162.200 162.800 166.600 163.100 ;
        RECT 181.400 163.100 181.800 163.200 ;
        RECT 193.400 163.100 193.800 163.200 ;
        RECT 181.400 162.800 193.800 163.100 ;
        RECT 196.600 163.100 197.000 163.200 ;
        RECT 213.400 163.100 213.800 163.200 ;
        RECT 196.600 162.800 213.800 163.100 ;
        RECT 216.600 163.100 217.000 163.200 ;
        RECT 226.200 163.100 226.600 163.200 ;
        RECT 216.600 162.800 226.600 163.100 ;
        RECT 227.000 163.100 227.400 163.200 ;
        RECT 250.200 163.100 250.600 163.200 ;
        RECT 227.000 162.800 250.600 163.100 ;
        RECT 58.200 162.100 58.600 162.200 ;
        RECT 106.200 162.100 106.600 162.200 ;
        RECT 58.200 161.800 106.600 162.100 ;
        RECT 141.400 162.100 141.800 162.200 ;
        RECT 145.400 162.100 145.800 162.200 ;
        RECT 141.400 161.800 145.800 162.100 ;
        RECT 151.800 162.100 152.200 162.200 ;
        RECT 190.200 162.100 190.600 162.200 ;
        RECT 151.800 161.800 190.600 162.100 ;
        RECT 199.000 162.100 199.400 162.200 ;
        RECT 221.400 162.100 221.800 162.200 ;
        RECT 199.000 161.800 221.800 162.100 ;
        RECT 222.200 162.100 222.600 162.200 ;
        RECT 226.200 162.100 226.600 162.200 ;
        RECT 222.200 161.800 226.600 162.100 ;
        RECT 241.400 162.100 241.800 162.200 ;
        RECT 262.200 162.100 262.600 162.200 ;
        RECT 241.400 161.800 262.600 162.100 ;
        RECT 84.600 161.100 85.000 161.200 ;
        RECT 103.800 161.100 104.200 161.200 ;
        RECT 84.600 160.800 104.200 161.100 ;
        RECT 169.400 161.100 169.800 161.200 ;
        RECT 181.400 161.100 181.800 161.200 ;
        RECT 169.400 160.800 181.800 161.100 ;
        RECT 182.200 161.100 182.600 161.200 ;
        RECT 224.600 161.100 225.000 161.200 ;
        RECT 182.200 160.800 225.000 161.100 ;
        RECT 239.800 161.100 240.200 161.200 ;
        RECT 251.000 161.100 251.400 161.200 ;
        RECT 239.800 160.800 251.400 161.100 ;
        RECT 69.400 160.100 69.800 160.200 ;
        RECT 98.200 160.100 98.600 160.200 ;
        RECT 69.400 159.800 98.600 160.100 ;
        RECT 103.000 160.100 103.400 160.200 ;
        RECT 135.000 160.100 135.400 160.200 ;
        RECT 139.800 160.100 140.200 160.200 ;
        RECT 103.000 159.800 140.200 160.100 ;
        RECT 163.000 160.100 163.400 160.200 ;
        RECT 176.600 160.100 177.000 160.200 ;
        RECT 163.000 159.800 177.000 160.100 ;
        RECT 188.600 160.100 189.000 160.200 ;
        RECT 207.000 160.100 207.400 160.200 ;
        RECT 188.600 159.800 207.400 160.100 ;
        RECT 211.000 160.100 211.400 160.200 ;
        RECT 230.200 160.100 230.600 160.200 ;
        RECT 211.000 159.800 230.600 160.100 ;
        RECT 48.600 159.100 49.000 159.200 ;
        RECT 59.000 159.100 59.400 159.200 ;
        RECT 159.000 159.100 159.400 159.200 ;
        RECT 48.600 158.800 159.400 159.100 ;
        RECT 171.000 159.100 171.400 159.200 ;
        RECT 176.600 159.100 177.000 159.200 ;
        RECT 171.000 158.800 177.000 159.100 ;
        RECT 192.600 159.100 193.000 159.200 ;
        RECT 201.400 159.100 201.800 159.200 ;
        RECT 223.000 159.100 223.400 159.200 ;
        RECT 192.600 158.800 223.400 159.100 ;
        RECT 25.400 158.100 25.800 158.200 ;
        RECT 56.600 158.100 57.000 158.200 ;
        RECT 58.200 158.100 58.600 158.200 ;
        RECT 25.400 157.800 58.600 158.100 ;
        RECT 88.600 158.100 89.000 158.200 ;
        RECT 91.000 158.100 91.400 158.200 ;
        RECT 88.600 157.800 91.400 158.100 ;
        RECT 99.800 158.100 100.200 158.200 ;
        RECT 124.600 158.100 125.000 158.200 ;
        RECT 99.800 157.800 125.000 158.100 ;
        RECT 126.200 158.100 126.600 158.200 ;
        RECT 129.400 158.100 129.800 158.200 ;
        RECT 126.200 157.800 129.800 158.100 ;
        RECT 155.000 158.100 155.400 158.200 ;
        RECT 165.400 158.100 165.800 158.200 ;
        RECT 179.000 158.100 179.400 158.200 ;
        RECT 155.000 157.800 179.400 158.100 ;
        RECT 193.400 158.100 193.800 158.200 ;
        RECT 195.800 158.100 196.200 158.200 ;
        RECT 193.400 157.800 196.200 158.100 ;
        RECT 202.200 158.100 202.600 158.200 ;
        RECT 231.000 158.100 231.400 158.200 ;
        RECT 202.200 157.800 231.400 158.100 ;
        RECT 45.400 156.800 45.800 157.200 ;
        RECT 75.000 157.100 75.400 157.200 ;
        RECT 79.800 157.100 80.200 157.200 ;
        RECT 75.000 156.800 80.200 157.100 ;
        RECT 87.000 157.100 87.400 157.200 ;
        RECT 102.200 157.100 102.600 157.200 ;
        RECT 87.000 156.800 102.600 157.100 ;
        RECT 120.600 157.100 121.000 157.200 ;
        RECT 127.800 157.100 128.200 157.200 ;
        RECT 120.600 156.800 128.200 157.100 ;
        RECT 142.200 157.100 142.600 157.200 ;
        RECT 144.600 157.100 145.000 157.200 ;
        RECT 142.200 156.800 145.000 157.100 ;
        RECT 147.000 157.100 147.400 157.200 ;
        RECT 148.600 157.100 149.000 157.200 ;
        RECT 156.600 157.100 157.000 157.200 ;
        RECT 147.000 156.800 157.000 157.100 ;
        RECT 157.400 157.100 157.800 157.200 ;
        RECT 170.200 157.100 170.600 157.200 ;
        RECT 157.400 156.800 170.600 157.100 ;
        RECT 186.200 157.100 186.600 157.200 ;
        RECT 187.000 157.100 187.400 157.200 ;
        RECT 186.200 156.800 187.400 157.100 ;
        RECT 195.000 156.800 195.400 157.200 ;
        RECT 196.600 157.100 197.000 157.200 ;
        RECT 215.000 157.100 215.400 157.200 ;
        RECT 196.600 156.800 215.400 157.100 ;
        RECT 220.600 157.100 221.000 157.200 ;
        RECT 227.800 157.100 228.200 157.200 ;
        RECT 220.600 156.800 228.200 157.100 ;
        RECT 250.200 157.100 250.600 157.200 ;
        RECT 255.000 157.100 255.400 157.200 ;
        RECT 250.200 156.800 255.400 157.100 ;
        RECT 12.600 156.100 13.000 156.200 ;
        RECT 38.200 156.100 38.600 156.200 ;
        RECT 12.600 155.800 38.600 156.100 ;
        RECT 45.400 156.100 45.700 156.800 ;
        RECT 48.600 156.100 49.000 156.200 ;
        RECT 59.800 156.100 60.200 156.200 ;
        RECT 45.400 155.800 60.200 156.100 ;
        RECT 68.600 156.100 69.000 156.200 ;
        RECT 82.200 156.100 82.600 156.200 ;
        RECT 68.600 155.800 82.600 156.100 ;
        RECT 127.000 156.100 127.400 156.200 ;
        RECT 127.800 156.100 128.200 156.200 ;
        RECT 127.000 155.800 128.200 156.100 ;
        RECT 135.800 156.100 136.200 156.200 ;
        RECT 145.400 156.100 145.800 156.200 ;
        RECT 135.800 155.800 145.800 156.100 ;
        RECT 147.000 156.100 147.400 156.200 ;
        RECT 149.400 156.100 149.800 156.200 ;
        RECT 164.600 156.100 165.000 156.200 ;
        RECT 168.600 156.100 169.000 156.200 ;
        RECT 147.000 155.800 169.000 156.100 ;
        RECT 172.600 156.100 173.000 156.200 ;
        RECT 186.200 156.100 186.500 156.800 ;
        RECT 172.600 155.800 186.500 156.100 ;
        RECT 195.000 156.100 195.300 156.800 ;
        RECT 201.400 156.100 201.800 156.200 ;
        RECT 195.000 155.800 201.800 156.100 ;
        RECT 205.400 156.100 205.800 156.200 ;
        RECT 207.800 156.100 208.200 156.200 ;
        RECT 205.400 155.800 208.200 156.100 ;
        RECT 215.800 155.800 216.200 156.200 ;
        RECT 223.800 156.100 224.200 156.200 ;
        RECT 225.400 156.100 225.800 156.200 ;
        RECT 223.800 155.800 225.800 156.100 ;
        RECT 230.200 156.100 230.600 156.200 ;
        RECT 235.000 156.100 235.400 156.200 ;
        RECT 230.200 155.800 235.400 156.100 ;
        RECT 259.000 155.800 259.400 156.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 20.600 154.800 21.000 155.200 ;
        RECT 41.400 155.100 41.800 155.200 ;
        RECT 43.000 155.100 43.400 155.200 ;
        RECT 43.800 155.100 44.200 155.200 ;
        RECT 49.400 155.100 49.800 155.200 ;
        RECT 41.400 154.800 44.200 155.100 ;
        RECT 47.800 154.800 49.800 155.100 ;
        RECT 53.400 155.100 53.800 155.200 ;
        RECT 64.600 155.100 65.000 155.200 ;
        RECT 75.000 155.100 75.400 155.200 ;
        RECT 53.400 154.800 75.400 155.100 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 81.400 155.100 81.800 155.200 ;
        RECT 83.800 155.100 84.200 155.200 ;
        RECT 85.400 155.100 85.800 155.200 ;
        RECT 81.400 154.800 85.800 155.100 ;
        RECT 89.400 154.800 89.800 155.200 ;
        RECT 99.000 155.100 99.400 155.200 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 103.800 155.100 104.200 155.200 ;
        RECT 99.000 154.800 104.200 155.100 ;
        RECT 106.200 155.100 106.600 155.200 ;
        RECT 111.000 155.100 111.400 155.200 ;
        RECT 130.200 155.100 130.600 155.200 ;
        RECT 135.800 155.100 136.200 155.200 ;
        RECT 106.200 154.800 136.200 155.100 ;
        RECT 136.600 155.100 137.000 155.200 ;
        RECT 142.200 155.100 142.600 155.200 ;
        RECT 150.200 155.100 150.600 155.200 ;
        RECT 167.000 155.100 167.400 155.200 ;
        RECT 136.600 154.800 150.600 155.100 ;
        RECT 159.800 154.800 167.400 155.100 ;
        RECT 170.200 155.100 170.600 155.200 ;
        RECT 171.000 155.100 171.400 155.200 ;
        RECT 170.200 154.800 171.400 155.100 ;
        RECT 175.800 155.100 176.200 155.200 ;
        RECT 176.600 155.100 177.000 155.200 ;
        RECT 175.800 154.800 177.000 155.100 ;
        RECT 187.000 155.100 187.400 155.200 ;
        RECT 194.200 155.100 194.600 155.200 ;
        RECT 187.000 154.800 194.600 155.100 ;
        RECT 196.600 155.100 197.000 155.200 ;
        RECT 200.600 155.100 201.000 155.200 ;
        RECT 196.600 154.800 201.000 155.100 ;
        RECT 203.000 155.100 203.400 155.200 ;
        RECT 203.800 155.100 204.200 155.200 ;
        RECT 207.000 155.100 207.400 155.200 ;
        RECT 215.800 155.100 216.100 155.800 ;
        RECT 223.800 155.100 224.100 155.800 ;
        RECT 259.000 155.200 259.300 155.800 ;
        RECT 242.200 155.100 242.600 155.200 ;
        RECT 203.000 154.800 204.200 155.100 ;
        RECT 206.200 154.800 216.100 155.100 ;
        RECT 216.600 154.800 224.100 155.100 ;
        RECT 231.800 154.800 242.600 155.100 ;
        RECT 246.200 155.100 246.600 155.200 ;
        RECT 249.400 155.100 249.800 155.200 ;
        RECT 251.800 155.100 252.200 155.200 ;
        RECT 254.200 155.100 254.600 155.200 ;
        RECT 255.000 155.100 255.400 155.200 ;
        RECT 246.200 154.800 255.400 155.100 ;
        RECT 259.000 154.800 259.400 155.200 ;
        RECT 19.000 154.100 19.300 154.800 ;
        RECT 20.600 154.100 20.900 154.800 ;
        RECT 47.800 154.200 48.100 154.800 ;
        RECT 79.000 154.200 79.300 154.800 ;
        RECT 89.400 154.200 89.700 154.800 ;
        RECT 159.800 154.700 160.200 154.800 ;
        RECT 19.000 153.800 20.900 154.100 ;
        RECT 31.800 154.100 32.200 154.200 ;
        RECT 47.800 154.100 48.200 154.200 ;
        RECT 31.800 153.800 48.200 154.100 ;
        RECT 51.800 154.100 52.200 154.200 ;
        RECT 58.200 154.100 58.600 154.200 ;
        RECT 51.800 153.800 58.600 154.100 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 79.800 154.100 80.200 154.200 ;
        RECT 86.200 154.100 86.600 154.200 ;
        RECT 79.800 153.800 86.600 154.100 ;
        RECT 89.400 153.800 89.800 154.200 ;
        RECT 93.400 154.100 93.800 154.200 ;
        RECT 106.200 154.100 106.600 154.200 ;
        RECT 93.400 153.800 106.600 154.100 ;
        RECT 109.400 154.100 109.800 154.200 ;
        RECT 110.200 154.100 110.600 154.200 ;
        RECT 114.200 154.100 114.600 154.200 ;
        RECT 109.400 153.800 110.600 154.100 ;
        RECT 112.600 153.800 114.600 154.100 ;
        RECT 115.800 154.100 116.200 154.200 ;
        RECT 120.600 154.100 121.000 154.200 ;
        RECT 129.400 154.100 129.800 154.200 ;
        RECT 115.800 153.800 129.800 154.100 ;
        RECT 131.000 154.100 131.400 154.200 ;
        RECT 142.200 154.100 142.600 154.200 ;
        RECT 167.000 154.100 167.400 154.200 ;
        RECT 131.000 153.800 167.400 154.100 ;
        RECT 170.200 154.100 170.600 154.200 ;
        RECT 174.200 154.100 174.600 154.200 ;
        RECT 170.200 153.800 174.600 154.100 ;
        RECT 176.600 154.100 177.000 154.200 ;
        RECT 216.600 154.100 216.900 154.800 ;
        RECT 176.600 153.800 216.900 154.100 ;
        RECT 231.800 154.200 232.100 154.800 ;
        RECT 231.800 153.800 232.200 154.200 ;
        RECT 247.800 154.100 248.200 154.200 ;
        RECT 248.600 154.100 249.000 154.200 ;
        RECT 247.800 153.800 249.000 154.100 ;
        RECT 252.600 154.100 253.000 154.200 ;
        RECT 259.800 154.100 260.200 154.200 ;
        RECT 252.600 153.800 260.200 154.100 ;
        RECT 23.000 153.100 23.400 153.200 ;
        RECT 80.600 153.100 81.000 153.200 ;
        RECT 91.000 153.100 91.400 153.200 ;
        RECT 23.000 152.800 42.500 153.100 ;
        RECT 80.600 152.800 91.400 153.100 ;
        RECT 104.600 153.100 105.000 153.200 ;
        RECT 112.600 153.100 112.900 153.800 ;
        RECT 104.600 152.800 112.900 153.100 ;
        RECT 113.400 153.100 113.800 153.200 ;
        RECT 122.200 153.100 122.600 153.200 ;
        RECT 133.400 153.100 133.800 153.200 ;
        RECT 113.400 152.800 114.500 153.100 ;
        RECT 122.200 152.800 133.800 153.100 ;
        RECT 141.400 152.800 141.800 153.200 ;
        RECT 143.800 153.100 144.200 153.200 ;
        RECT 164.600 153.100 165.000 153.200 ;
        RECT 173.400 153.100 173.800 153.200 ;
        RECT 143.800 152.800 165.000 153.100 ;
        RECT 170.200 152.800 173.800 153.100 ;
        RECT 175.000 153.100 175.400 153.200 ;
        RECT 201.400 153.100 201.800 153.200 ;
        RECT 203.800 153.100 204.200 153.200 ;
        RECT 175.000 152.800 204.200 153.100 ;
        RECT 207.000 153.100 207.400 153.200 ;
        RECT 208.600 153.100 209.000 153.200 ;
        RECT 207.000 152.800 209.000 153.100 ;
        RECT 214.200 153.100 214.600 153.200 ;
        RECT 217.400 153.100 217.800 153.200 ;
        RECT 214.200 152.800 217.800 153.100 ;
        RECT 219.800 153.100 220.200 153.200 ;
        RECT 238.200 153.100 238.600 153.200 ;
        RECT 219.800 152.800 238.600 153.100 ;
        RECT 242.200 153.100 242.600 153.200 ;
        RECT 255.000 153.100 255.400 153.200 ;
        RECT 242.200 152.800 255.400 153.100 ;
        RECT 42.200 152.200 42.500 152.800 ;
        RECT 29.400 152.100 29.800 152.200 ;
        RECT 39.000 152.100 39.400 152.200 ;
        RECT 29.400 151.800 39.400 152.100 ;
        RECT 42.200 151.800 42.600 152.200 ;
        RECT 59.800 152.100 60.200 152.200 ;
        RECT 69.400 152.100 69.800 152.200 ;
        RECT 90.200 152.100 90.600 152.200 ;
        RECT 59.800 151.800 90.600 152.100 ;
        RECT 91.800 152.100 92.200 152.200 ;
        RECT 113.400 152.100 113.800 152.200 ;
        RECT 91.800 151.800 113.800 152.100 ;
        RECT 114.200 152.100 114.500 152.800 ;
        RECT 141.400 152.200 141.700 152.800 ;
        RECT 170.200 152.200 170.500 152.800 ;
        RECT 136.600 152.100 137.000 152.200 ;
        RECT 114.200 151.800 137.000 152.100 ;
        RECT 141.400 151.800 141.800 152.200 ;
        RECT 143.000 152.100 143.400 152.200 ;
        RECT 159.800 152.100 160.200 152.200 ;
        RECT 167.000 152.100 167.400 152.200 ;
        RECT 143.000 151.800 167.400 152.100 ;
        RECT 170.200 151.800 170.600 152.200 ;
        RECT 187.000 152.100 187.400 152.200 ;
        RECT 191.800 152.100 192.200 152.200 ;
        RECT 187.000 151.800 192.200 152.100 ;
        RECT 224.600 152.100 225.000 152.200 ;
        RECT 226.200 152.100 226.600 152.200 ;
        RECT 224.600 151.800 226.600 152.100 ;
        RECT 45.400 151.100 45.800 151.200 ;
        RECT 66.200 151.100 66.600 151.200 ;
        RECT 45.400 150.800 66.600 151.100 ;
        RECT 84.600 151.100 85.000 151.200 ;
        RECT 96.600 151.100 97.000 151.200 ;
        RECT 84.600 150.800 97.000 151.100 ;
        RECT 111.000 151.100 111.400 151.200 ;
        RECT 121.400 151.100 121.800 151.200 ;
        RECT 111.000 150.800 121.800 151.100 ;
        RECT 126.200 151.100 126.600 151.200 ;
        RECT 131.800 151.100 132.200 151.200 ;
        RECT 126.200 150.800 132.200 151.100 ;
        RECT 143.800 151.100 144.200 151.200 ;
        RECT 144.600 151.100 145.000 151.200 ;
        RECT 143.800 150.800 145.000 151.100 ;
        RECT 145.400 151.100 145.800 151.200 ;
        RECT 149.400 151.100 149.800 151.200 ;
        RECT 145.400 150.800 149.800 151.100 ;
        RECT 153.400 151.100 153.800 151.200 ;
        RECT 155.000 151.100 155.400 151.200 ;
        RECT 153.400 150.800 155.400 151.100 ;
        RECT 158.200 151.100 158.600 151.200 ;
        RECT 162.200 151.100 162.600 151.200 ;
        RECT 158.200 150.800 162.600 151.100 ;
        RECT 168.600 151.100 169.000 151.200 ;
        RECT 192.600 151.100 193.000 151.200 ;
        RECT 168.600 150.800 193.000 151.100 ;
        RECT 223.800 151.100 224.200 151.200 ;
        RECT 225.400 151.100 225.800 151.200 ;
        RECT 227.000 151.100 227.400 151.200 ;
        RECT 223.800 150.800 227.400 151.100 ;
        RECT 235.800 151.100 236.200 151.200 ;
        RECT 247.000 151.100 247.400 151.200 ;
        RECT 235.800 150.800 247.400 151.100 ;
        RECT 10.200 150.100 10.600 150.200 ;
        RECT 15.800 150.100 16.200 150.200 ;
        RECT 10.200 149.800 16.200 150.100 ;
        RECT 39.000 150.100 39.400 150.200 ;
        RECT 74.200 150.100 74.600 150.200 ;
        RECT 39.000 149.800 74.600 150.100 ;
        RECT 75.800 150.100 76.200 150.200 ;
        RECT 78.200 150.100 78.600 150.200 ;
        RECT 85.400 150.100 85.800 150.200 ;
        RECT 75.800 149.800 85.800 150.100 ;
        RECT 88.600 150.100 89.000 150.200 ;
        RECT 91.800 150.100 92.200 150.200 ;
        RECT 88.600 149.800 92.200 150.100 ;
        RECT 114.200 150.100 114.600 150.200 ;
        RECT 122.200 150.100 122.600 150.200 ;
        RECT 114.200 149.800 122.600 150.100 ;
        RECT 138.200 150.100 138.600 150.200 ;
        RECT 167.000 150.100 167.400 150.200 ;
        RECT 138.200 149.800 167.400 150.100 ;
        RECT 181.400 150.100 181.800 150.200 ;
        RECT 187.000 150.100 187.400 150.200 ;
        RECT 199.000 150.100 199.400 150.200 ;
        RECT 181.400 149.800 199.400 150.100 ;
        RECT 227.800 150.100 228.200 150.200 ;
        RECT 241.400 150.100 241.800 150.200 ;
        RECT 227.800 149.800 241.800 150.100 ;
        RECT 10.200 149.100 10.600 149.200 ;
        RECT 18.200 149.100 18.600 149.200 ;
        RECT 10.200 148.800 18.600 149.100 ;
        RECT 39.000 149.100 39.400 149.200 ;
        RECT 67.000 149.100 67.400 149.200 ;
        RECT 39.000 148.800 67.400 149.100 ;
        RECT 84.600 149.100 85.000 149.200 ;
        RECT 110.200 149.100 110.600 149.200 ;
        RECT 84.600 148.800 110.600 149.100 ;
        RECT 112.600 149.100 113.000 149.200 ;
        RECT 133.400 149.100 133.800 149.200 ;
        RECT 160.600 149.100 161.000 149.200 ;
        RECT 112.600 148.800 161.000 149.100 ;
        RECT 168.600 149.100 169.000 149.200 ;
        RECT 169.400 149.100 169.800 149.200 ;
        RECT 168.600 148.800 169.800 149.100 ;
        RECT 183.000 149.100 183.400 149.200 ;
        RECT 204.600 149.100 205.000 149.200 ;
        RECT 183.000 148.800 205.000 149.100 ;
        RECT 241.400 149.100 241.700 149.800 ;
        RECT 244.600 149.100 245.000 149.200 ;
        RECT 241.400 148.800 245.000 149.100 ;
        RECT 247.000 149.100 247.400 149.200 ;
        RECT 249.400 149.100 249.800 149.200 ;
        RECT 247.000 148.800 249.800 149.100 ;
        RECT 3.800 148.100 4.200 148.200 ;
        RECT 13.400 148.100 13.800 148.200 ;
        RECT 23.800 148.100 24.200 148.200 ;
        RECT 3.800 147.800 10.500 148.100 ;
        RECT 13.400 147.800 24.200 148.100 ;
        RECT 51.800 148.100 52.200 148.200 ;
        RECT 99.800 148.100 100.200 148.200 ;
        RECT 51.800 147.800 100.200 148.100 ;
        RECT 103.800 148.100 104.200 148.200 ;
        RECT 111.800 148.100 112.200 148.200 ;
        RECT 103.800 147.800 112.200 148.100 ;
        RECT 115.000 148.100 115.400 148.200 ;
        RECT 118.200 148.100 118.600 148.200 ;
        RECT 115.000 147.800 118.600 148.100 ;
        RECT 126.200 148.100 126.600 148.200 ;
        RECT 127.000 148.100 127.400 148.200 ;
        RECT 126.200 147.800 127.400 148.100 ;
        RECT 128.600 148.100 129.000 148.200 ;
        RECT 131.800 148.100 132.200 148.200 ;
        RECT 146.200 148.100 146.600 148.200 ;
        RECT 147.000 148.100 147.400 148.200 ;
        RECT 128.600 147.800 147.400 148.100 ;
        RECT 147.800 148.100 148.200 148.200 ;
        RECT 154.200 148.100 154.600 148.200 ;
        RECT 147.800 147.800 154.600 148.100 ;
        RECT 162.200 148.100 162.600 148.200 ;
        RECT 191.800 148.100 192.200 148.200 ;
        RECT 162.200 147.800 192.200 148.100 ;
        RECT 192.600 148.100 193.000 148.200 ;
        RECT 207.000 148.100 207.400 148.200 ;
        RECT 192.600 147.800 207.400 148.100 ;
        RECT 217.400 148.100 217.800 148.200 ;
        RECT 233.400 148.100 233.800 148.200 ;
        RECT 217.400 147.800 233.800 148.100 ;
        RECT 10.200 147.200 10.500 147.800 ;
        RECT 10.200 146.800 10.600 147.200 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 15.000 147.100 15.400 147.200 ;
        RECT 19.000 147.100 19.400 147.200 ;
        RECT 19.800 147.100 20.200 147.200 ;
        RECT 14.200 146.800 15.400 147.100 ;
        RECT 18.200 146.800 20.200 147.100 ;
        RECT 23.800 147.100 24.200 147.200 ;
        RECT 41.400 147.100 41.800 147.200 ;
        RECT 47.000 147.100 47.400 147.200 ;
        RECT 58.200 147.100 58.600 147.200 ;
        RECT 65.400 147.100 65.800 147.200 ;
        RECT 71.800 147.100 72.200 147.200 ;
        RECT 23.800 146.800 47.400 147.100 ;
        RECT 48.600 146.800 50.500 147.100 ;
        RECT 58.200 146.800 72.200 147.100 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 80.600 147.100 81.000 147.200 ;
        RECT 79.800 146.800 81.000 147.100 ;
        RECT 82.200 146.800 82.600 147.200 ;
        RECT 96.600 147.100 97.000 147.200 ;
        RECT 109.400 147.100 109.800 147.200 ;
        RECT 96.600 146.800 109.800 147.100 ;
        RECT 132.600 147.100 133.000 147.200 ;
        RECT 134.200 147.100 134.600 147.200 ;
        RECT 132.600 146.800 134.600 147.100 ;
        RECT 140.600 147.100 141.000 147.200 ;
        RECT 145.400 147.100 145.800 147.200 ;
        RECT 159.000 147.100 159.400 147.200 ;
        RECT 160.600 147.100 161.000 147.200 ;
        RECT 161.400 147.100 161.800 147.200 ;
        RECT 140.600 146.800 161.800 147.100 ;
        RECT 167.800 147.100 168.200 147.200 ;
        RECT 175.000 147.100 175.400 147.200 ;
        RECT 167.800 146.800 175.400 147.100 ;
        RECT 199.800 147.100 200.200 147.200 ;
        RECT 203.800 147.100 204.200 147.200 ;
        RECT 199.800 146.800 204.200 147.100 ;
        RECT 204.600 147.100 205.000 147.200 ;
        RECT 215.000 147.100 215.400 147.200 ;
        RECT 204.600 146.800 215.400 147.100 ;
        RECT 225.400 146.800 225.800 147.200 ;
        RECT 231.000 147.100 231.400 147.200 ;
        RECT 231.800 147.100 232.200 147.200 ;
        RECT 231.000 146.800 232.200 147.100 ;
        RECT 238.200 147.100 238.600 147.200 ;
        RECT 241.400 147.100 241.800 147.200 ;
        RECT 238.200 146.800 241.800 147.100 ;
        RECT 244.600 147.100 245.000 147.200 ;
        RECT 255.800 147.100 256.200 147.200 ;
        RECT 244.600 146.800 256.200 147.100 ;
        RECT 48.600 146.200 48.900 146.800 ;
        RECT 50.200 146.200 50.500 146.800 ;
        RECT 13.400 146.100 13.800 146.200 ;
        RECT 16.600 146.100 17.000 146.200 ;
        RECT 13.400 145.800 17.000 146.100 ;
        RECT 18.200 146.100 18.600 146.200 ;
        RECT 19.000 146.100 19.400 146.200 ;
        RECT 18.200 145.800 19.400 146.100 ;
        RECT 36.600 146.100 37.000 146.200 ;
        RECT 39.000 146.100 39.400 146.200 ;
        RECT 36.600 145.800 39.400 146.100 ;
        RECT 48.600 145.800 49.000 146.200 ;
        RECT 50.200 145.800 50.600 146.200 ;
        RECT 53.400 146.100 53.800 146.200 ;
        RECT 63.000 146.100 63.400 146.200 ;
        RECT 71.800 146.100 72.200 146.200 ;
        RECT 75.000 146.100 75.400 146.200 ;
        RECT 53.400 145.800 63.400 146.100 ;
        RECT 71.000 145.800 75.400 146.100 ;
        RECT 82.200 146.100 82.500 146.800 ;
        RECT 87.000 146.100 87.400 146.200 ;
        RECT 82.200 145.800 87.400 146.100 ;
        RECT 92.600 146.100 93.000 146.200 ;
        RECT 93.400 146.100 93.800 146.200 ;
        RECT 92.600 145.800 93.800 146.100 ;
        RECT 97.400 146.100 97.800 146.200 ;
        RECT 98.200 146.100 98.600 146.200 ;
        RECT 97.400 145.800 98.600 146.100 ;
        RECT 100.600 146.100 101.000 146.200 ;
        RECT 101.400 146.100 101.800 146.200 ;
        RECT 100.600 145.800 101.800 146.100 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 113.400 146.100 113.800 146.200 ;
        RECT 112.600 145.800 113.800 146.100 ;
        RECT 119.000 146.100 119.400 146.200 ;
        RECT 126.200 146.100 126.600 146.200 ;
        RECT 119.000 145.800 126.600 146.100 ;
        RECT 135.800 146.100 136.200 146.200 ;
        RECT 142.200 146.100 142.600 146.200 ;
        RECT 135.800 145.800 142.600 146.100 ;
        RECT 144.600 146.100 145.000 146.200 ;
        RECT 163.000 146.100 163.400 146.200 ;
        RECT 144.600 145.800 163.400 146.100 ;
        RECT 179.000 146.100 179.400 146.200 ;
        RECT 182.200 146.100 182.600 146.200 ;
        RECT 185.400 146.100 185.800 146.200 ;
        RECT 179.000 145.800 185.800 146.100 ;
        RECT 192.600 146.100 193.000 146.300 ;
        RECT 198.200 146.100 198.600 146.200 ;
        RECT 192.600 145.800 198.600 146.100 ;
        RECT 200.600 145.800 201.000 146.200 ;
        RECT 204.600 146.100 205.000 146.200 ;
        RECT 203.000 145.800 205.000 146.100 ;
        RECT 210.200 146.100 210.600 146.200 ;
        RECT 225.400 146.100 225.700 146.800 ;
        RECT 247.000 146.100 247.400 146.200 ;
        RECT 210.200 145.800 219.300 146.100 ;
        RECT 225.400 145.800 247.400 146.100 ;
        RECT 71.000 145.200 71.300 145.800 ;
        RECT 148.600 145.200 148.900 145.800 ;
        RECT 200.600 145.200 200.900 145.800 ;
        RECT 203.000 145.200 203.300 145.800 ;
        RECT 219.000 145.200 219.300 145.800 ;
        RECT 3.800 145.100 4.200 145.200 ;
        RECT 35.000 145.100 35.400 145.200 ;
        RECT 40.600 145.100 41.000 145.200 ;
        RECT 3.800 144.800 14.500 145.100 ;
        RECT 35.000 144.800 41.000 145.100 ;
        RECT 61.400 145.100 61.800 145.200 ;
        RECT 63.800 145.100 64.200 145.200 ;
        RECT 61.400 144.800 64.200 145.100 ;
        RECT 66.200 145.100 66.600 145.200 ;
        RECT 70.200 145.100 70.600 145.200 ;
        RECT 66.200 144.800 70.600 145.100 ;
        RECT 71.000 144.800 71.400 145.200 ;
        RECT 75.000 145.100 75.400 145.200 ;
        RECT 100.600 145.100 101.000 145.200 ;
        RECT 75.000 144.800 101.000 145.100 ;
        RECT 102.200 145.100 102.600 145.200 ;
        RECT 107.000 145.100 107.400 145.200 ;
        RECT 135.000 145.100 135.400 145.200 ;
        RECT 102.200 144.800 135.400 145.100 ;
        RECT 143.000 145.100 143.400 145.200 ;
        RECT 147.000 145.100 147.400 145.200 ;
        RECT 143.000 144.800 147.400 145.100 ;
        RECT 148.600 144.800 149.000 145.200 ;
        RECT 158.200 145.100 158.600 145.200 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 158.200 144.800 159.400 145.100 ;
        RECT 160.600 145.100 161.000 145.200 ;
        RECT 182.200 145.100 182.600 145.200 ;
        RECT 187.800 145.100 188.200 145.200 ;
        RECT 160.600 144.800 188.200 145.100 ;
        RECT 193.400 145.100 193.800 145.200 ;
        RECT 197.400 145.100 197.800 145.200 ;
        RECT 193.400 144.800 197.800 145.100 ;
        RECT 200.600 144.800 201.000 145.200 ;
        RECT 203.000 144.800 203.400 145.200 ;
        RECT 203.800 145.100 204.200 145.200 ;
        RECT 209.400 145.100 209.800 145.200 ;
        RECT 203.800 144.800 209.800 145.100 ;
        RECT 219.000 144.800 219.400 145.200 ;
        RECT 243.000 145.100 243.400 145.200 ;
        RECT 244.600 145.100 245.000 145.200 ;
        RECT 248.600 145.100 249.000 145.200 ;
        RECT 243.000 144.800 249.000 145.100 ;
        RECT 14.200 144.200 14.500 144.800 ;
        RECT 14.200 143.800 14.600 144.200 ;
        RECT 16.600 144.100 17.000 144.200 ;
        RECT 61.400 144.100 61.700 144.800 ;
        RECT 16.600 143.800 61.700 144.100 ;
        RECT 81.400 144.100 81.800 144.200 ;
        RECT 99.800 144.100 100.200 144.200 ;
        RECT 103.800 144.100 104.200 144.200 ;
        RECT 107.800 144.100 108.200 144.200 ;
        RECT 81.400 143.800 108.200 144.100 ;
        RECT 120.600 144.100 121.000 144.200 ;
        RECT 121.400 144.100 121.800 144.200 ;
        RECT 120.600 143.800 121.800 144.100 ;
        RECT 122.200 144.100 122.600 144.200 ;
        RECT 139.000 144.100 139.400 144.200 ;
        RECT 122.200 143.800 139.400 144.100 ;
        RECT 142.200 144.100 142.600 144.200 ;
        RECT 143.000 144.100 143.400 144.200 ;
        RECT 142.200 143.800 143.400 144.100 ;
        RECT 146.200 144.100 146.600 144.200 ;
        RECT 151.000 144.100 151.400 144.200 ;
        RECT 146.200 143.800 151.400 144.100 ;
        RECT 162.200 144.100 162.600 144.200 ;
        RECT 163.000 144.100 163.400 144.200 ;
        RECT 172.600 144.100 173.000 144.200 ;
        RECT 196.600 144.100 197.000 144.200 ;
        RECT 228.600 144.100 229.000 144.200 ;
        RECT 231.000 144.100 231.400 144.200 ;
        RECT 162.200 143.800 231.400 144.100 ;
        RECT 37.400 143.100 37.800 143.200 ;
        RECT 52.600 143.100 53.000 143.200 ;
        RECT 60.600 143.100 61.000 143.200 ;
        RECT 37.400 142.800 61.000 143.100 ;
        RECT 71.000 143.100 71.400 143.200 ;
        RECT 102.200 143.100 102.600 143.200 ;
        RECT 71.000 142.800 102.600 143.100 ;
        RECT 120.600 143.100 121.000 143.200 ;
        RECT 143.000 143.100 143.400 143.200 ;
        RECT 120.600 142.800 143.400 143.100 ;
        RECT 159.800 143.100 160.200 143.200 ;
        RECT 171.000 143.100 171.400 143.200 ;
        RECT 177.400 143.100 177.800 143.200 ;
        RECT 159.800 142.800 177.800 143.100 ;
        RECT 203.000 143.100 203.400 143.200 ;
        RECT 226.200 143.100 226.600 143.200 ;
        RECT 203.000 142.800 226.600 143.100 ;
        RECT 260.600 143.100 261.000 143.200 ;
        RECT 263.000 143.100 263.400 143.200 ;
        RECT 260.600 142.800 263.400 143.100 ;
        RECT 16.600 142.100 17.000 142.200 ;
        RECT 27.000 142.100 27.400 142.200 ;
        RECT 31.000 142.100 31.400 142.200 ;
        RECT 72.600 142.100 73.000 142.200 ;
        RECT 16.600 141.800 73.000 142.100 ;
        RECT 83.800 142.100 84.200 142.200 ;
        RECT 84.600 142.100 85.000 142.200 ;
        RECT 83.800 141.800 85.000 142.100 ;
        RECT 99.800 142.100 100.200 142.200 ;
        RECT 134.200 142.100 134.600 142.200 ;
        RECT 140.600 142.100 141.000 142.200 ;
        RECT 99.800 141.800 141.000 142.100 ;
        RECT 143.000 142.100 143.300 142.800 ;
        RECT 148.600 142.100 149.000 142.200 ;
        RECT 143.000 141.800 149.000 142.100 ;
        RECT 151.800 142.100 152.200 142.200 ;
        RECT 154.200 142.100 154.600 142.200 ;
        RECT 161.400 142.100 161.800 142.200 ;
        RECT 151.800 141.800 161.800 142.100 ;
        RECT 175.000 142.100 175.400 142.200 ;
        RECT 179.000 142.100 179.400 142.200 ;
        RECT 175.000 141.800 179.400 142.100 ;
        RECT 180.600 142.100 181.000 142.200 ;
        RECT 206.200 142.100 206.600 142.200 ;
        RECT 180.600 141.800 206.600 142.100 ;
        RECT 207.800 142.100 208.200 142.200 ;
        RECT 242.200 142.100 242.600 142.200 ;
        RECT 207.800 141.800 242.600 142.100 ;
        RECT 9.400 141.100 9.800 141.200 ;
        RECT 22.200 141.100 22.600 141.200 ;
        RECT 9.400 140.800 22.600 141.100 ;
        RECT 102.200 141.100 102.600 141.200 ;
        RECT 118.200 141.100 118.600 141.200 ;
        RECT 135.800 141.100 136.200 141.200 ;
        RECT 138.200 141.100 138.600 141.200 ;
        RECT 146.200 141.100 146.600 141.200 ;
        RECT 102.200 140.800 146.600 141.100 ;
        RECT 149.400 141.100 149.800 141.200 ;
        RECT 155.000 141.100 155.400 141.200 ;
        RECT 149.400 140.800 155.400 141.100 ;
        RECT 168.600 141.100 169.000 141.200 ;
        RECT 183.000 141.100 183.400 141.200 ;
        RECT 168.600 140.800 183.400 141.100 ;
        RECT 196.600 141.100 197.000 141.200 ;
        RECT 198.200 141.100 198.600 141.200 ;
        RECT 196.600 140.800 198.600 141.100 ;
        RECT 206.200 141.100 206.600 141.200 ;
        RECT 211.800 141.100 212.200 141.200 ;
        RECT 206.200 140.800 212.200 141.100 ;
        RECT 219.000 141.100 219.400 141.200 ;
        RECT 260.600 141.100 261.000 141.200 ;
        RECT 219.000 140.800 261.000 141.100 ;
        RECT 87.800 140.100 88.200 140.200 ;
        RECT 107.000 140.100 107.400 140.200 ;
        RECT 87.800 139.800 107.400 140.100 ;
        RECT 131.800 140.100 132.200 140.200 ;
        RECT 132.600 140.100 133.000 140.200 ;
        RECT 131.800 139.800 133.000 140.100 ;
        RECT 139.800 140.100 140.200 140.200 ;
        RECT 145.400 140.100 145.800 140.200 ;
        RECT 139.800 139.800 145.800 140.100 ;
        RECT 146.200 140.100 146.600 140.200 ;
        RECT 155.000 140.100 155.400 140.200 ;
        RECT 146.200 139.800 155.400 140.100 ;
        RECT 179.000 140.100 179.400 140.200 ;
        RECT 180.600 140.100 181.000 140.200 ;
        RECT 179.000 139.800 181.000 140.100 ;
        RECT 182.200 140.100 182.600 140.200 ;
        RECT 195.000 140.100 195.400 140.200 ;
        RECT 211.000 140.100 211.400 140.200 ;
        RECT 182.200 139.800 211.400 140.100 ;
        RECT 88.600 139.100 89.000 139.200 ;
        RECT 91.000 139.100 91.400 139.200 ;
        RECT 88.600 138.800 91.400 139.100 ;
        RECT 103.800 138.800 104.200 139.200 ;
        RECT 137.400 139.100 137.800 139.200 ;
        RECT 147.800 139.100 148.200 139.200 ;
        RECT 150.200 139.100 150.600 139.200 ;
        RECT 158.200 139.100 158.600 139.200 ;
        RECT 137.400 138.800 150.600 139.100 ;
        RECT 155.800 138.800 158.600 139.100 ;
        RECT 165.400 139.100 165.800 139.200 ;
        RECT 167.800 139.100 168.200 139.200 ;
        RECT 207.800 139.100 208.200 139.200 ;
        RECT 254.200 139.100 254.600 139.200 ;
        RECT 165.400 138.800 254.600 139.100 ;
        RECT 19.800 138.100 20.200 138.200 ;
        RECT 33.400 138.100 33.800 138.200 ;
        RECT 19.800 137.800 33.800 138.100 ;
        RECT 72.600 138.100 73.000 138.200 ;
        RECT 103.800 138.100 104.100 138.800 ;
        RECT 155.800 138.200 156.100 138.800 ;
        RECT 72.600 137.800 104.100 138.100 ;
        RECT 137.400 138.100 137.800 138.200 ;
        RECT 139.800 138.100 140.200 138.200 ;
        RECT 155.000 138.100 155.400 138.200 ;
        RECT 137.400 137.800 155.400 138.100 ;
        RECT 155.800 137.800 156.200 138.200 ;
        RECT 179.000 137.800 179.400 138.200 ;
        RECT 182.200 138.100 182.600 138.200 ;
        RECT 229.400 138.100 229.800 138.200 ;
        RECT 182.200 137.800 229.800 138.100 ;
        RECT 27.800 137.100 28.200 137.200 ;
        RECT 28.600 137.100 29.000 137.200 ;
        RECT 27.800 136.800 29.000 137.100 ;
        RECT 29.400 137.100 29.800 137.200 ;
        RECT 33.400 137.100 33.800 137.200 ;
        RECT 29.400 136.800 33.800 137.100 ;
        RECT 56.600 136.800 57.000 137.200 ;
        RECT 60.600 137.100 61.000 137.200 ;
        RECT 86.200 137.100 86.600 137.200 ;
        RECT 90.200 137.100 90.600 137.200 ;
        RECT 60.600 136.800 90.600 137.100 ;
        RECT 99.800 136.800 100.200 137.200 ;
        RECT 104.600 137.100 105.000 137.200 ;
        RECT 105.400 137.100 105.800 137.200 ;
        RECT 104.600 136.800 105.800 137.100 ;
        RECT 119.800 137.100 120.200 137.200 ;
        RECT 140.600 137.100 141.000 137.200 ;
        RECT 145.400 137.100 145.800 137.200 ;
        RECT 119.800 136.800 145.800 137.100 ;
        RECT 151.000 137.100 151.400 137.200 ;
        RECT 173.400 137.100 173.800 137.200 ;
        RECT 151.000 136.800 173.800 137.100 ;
        RECT 178.200 136.800 178.600 137.200 ;
        RECT 179.000 137.100 179.300 137.800 ;
        RECT 183.800 137.100 184.200 137.200 ;
        RECT 210.200 137.100 210.600 137.200 ;
        RECT 179.000 136.800 210.600 137.100 ;
        RECT 211.000 137.100 211.400 137.200 ;
        RECT 241.400 137.100 241.800 137.200 ;
        RECT 211.000 136.800 241.800 137.100 ;
        RECT 256.600 137.100 257.000 137.200 ;
        RECT 258.200 137.100 258.600 137.200 ;
        RECT 256.600 136.800 258.600 137.100 ;
        RECT 11.800 136.100 12.200 136.200 ;
        RECT 14.200 136.100 14.600 136.200 ;
        RECT 43.000 136.100 43.400 136.200 ;
        RECT 11.800 135.800 43.400 136.100 ;
        RECT 47.800 136.100 48.200 136.200 ;
        RECT 56.600 136.100 56.900 136.800 ;
        RECT 47.800 135.800 56.900 136.100 ;
        RECT 85.400 136.100 85.800 136.200 ;
        RECT 86.200 136.100 86.600 136.200 ;
        RECT 85.400 135.800 86.600 136.100 ;
        RECT 88.600 136.100 89.000 136.200 ;
        RECT 99.800 136.100 100.100 136.800 ;
        RECT 178.200 136.200 178.500 136.800 ;
        RECT 88.600 135.800 100.100 136.100 ;
        RECT 100.600 136.100 101.000 136.200 ;
        RECT 107.000 136.100 107.400 136.200 ;
        RECT 107.800 136.100 108.200 136.200 ;
        RECT 110.200 136.100 110.600 136.200 ;
        RECT 100.600 135.800 110.600 136.100 ;
        RECT 121.400 136.100 121.800 136.200 ;
        RECT 124.600 136.100 125.000 136.200 ;
        RECT 131.000 136.100 131.400 136.200 ;
        RECT 148.600 136.100 149.000 136.200 ;
        RECT 152.600 136.100 153.000 136.200 ;
        RECT 121.400 135.800 153.000 136.100 ;
        RECT 164.600 136.100 165.000 136.200 ;
        RECT 168.600 136.100 169.000 136.200 ;
        RECT 164.600 135.800 169.000 136.100 ;
        RECT 178.200 136.100 178.600 136.200 ;
        RECT 180.600 136.100 181.000 136.200 ;
        RECT 178.200 135.800 181.000 136.100 ;
        RECT 183.800 136.100 184.200 136.200 ;
        RECT 193.400 136.100 193.800 136.200 ;
        RECT 183.800 135.800 193.800 136.100 ;
        RECT 194.200 136.100 194.600 136.200 ;
        RECT 197.400 136.100 197.800 136.200 ;
        RECT 199.800 136.100 200.200 136.200 ;
        RECT 194.200 135.800 200.200 136.100 ;
        RECT 207.000 136.100 207.400 136.200 ;
        RECT 212.600 136.100 213.000 136.200 ;
        RECT 207.000 135.800 213.000 136.100 ;
        RECT 215.800 136.100 216.200 136.200 ;
        RECT 216.600 136.100 217.000 136.200 ;
        RECT 215.800 135.800 217.000 136.100 ;
        RECT 217.400 135.800 217.800 136.200 ;
        RECT 220.600 136.100 221.000 136.200 ;
        RECT 238.200 136.100 238.600 136.200 ;
        RECT 220.600 135.800 238.600 136.100 ;
        RECT 243.000 136.100 243.400 136.200 ;
        RECT 243.000 135.800 257.700 136.100 ;
        RECT 4.600 135.100 5.000 135.200 ;
        RECT 12.600 135.100 13.000 135.200 ;
        RECT 4.600 134.800 13.000 135.100 ;
        RECT 21.400 135.100 21.800 135.200 ;
        RECT 23.000 135.100 23.400 135.200 ;
        RECT 21.400 134.800 23.400 135.100 ;
        RECT 25.400 135.100 25.800 135.200 ;
        RECT 56.600 135.100 57.000 135.200 ;
        RECT 63.000 135.100 63.400 135.200 ;
        RECT 72.600 135.100 73.000 135.200 ;
        RECT 25.400 134.800 73.000 135.100 ;
        RECT 82.200 135.100 82.600 135.200 ;
        RECT 86.200 135.100 86.600 135.200 ;
        RECT 82.200 134.800 86.600 135.100 ;
        RECT 100.600 135.100 101.000 135.200 ;
        RECT 101.400 135.100 101.800 135.200 ;
        RECT 100.600 134.800 101.800 135.100 ;
        RECT 102.200 135.100 102.600 135.200 ;
        RECT 106.200 135.100 106.600 135.200 ;
        RECT 108.600 135.100 109.000 135.200 ;
        RECT 102.200 134.800 109.000 135.100 ;
        RECT 109.400 135.100 109.800 135.200 ;
        RECT 111.800 135.100 112.200 135.200 ;
        RECT 109.400 134.800 112.200 135.100 ;
        RECT 115.000 135.100 115.400 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 115.000 134.800 123.400 135.100 ;
        RECT 125.400 135.100 125.800 135.200 ;
        RECT 132.600 135.100 133.000 135.200 ;
        RECT 125.400 134.800 133.000 135.100 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 144.600 135.100 145.000 135.200 ;
        RECT 147.000 135.100 147.400 135.200 ;
        RECT 155.000 135.100 155.400 135.200 ;
        RECT 163.800 135.100 164.200 135.200 ;
        RECT 136.600 134.800 164.200 135.100 ;
        RECT 166.200 135.100 166.600 135.200 ;
        RECT 199.800 135.100 200.200 135.200 ;
        RECT 201.400 135.100 201.800 135.200 ;
        RECT 166.200 134.800 201.800 135.100 ;
        RECT 202.200 135.100 202.600 135.200 ;
        RECT 203.800 135.100 204.200 135.200 ;
        RECT 202.200 134.800 204.200 135.100 ;
        RECT 205.400 135.100 205.800 135.200 ;
        RECT 212.600 135.100 213.000 135.200 ;
        RECT 205.400 134.800 213.000 135.100 ;
        RECT 215.800 135.100 216.200 135.200 ;
        RECT 217.400 135.100 217.700 135.800 ;
        RECT 257.400 135.200 257.700 135.800 ;
        RECT 215.800 134.800 217.700 135.100 ;
        RECT 219.000 135.100 219.400 135.200 ;
        RECT 219.800 135.100 220.200 135.200 ;
        RECT 219.000 134.800 220.200 135.100 ;
        RECT 231.800 134.800 232.200 135.200 ;
        RECT 250.200 134.800 255.300 135.100 ;
        RECT 257.400 134.800 257.800 135.200 ;
        RECT 30.200 134.100 30.600 134.200 ;
        RECT 31.000 134.100 31.400 134.200 ;
        RECT 30.200 133.800 31.400 134.100 ;
        RECT 31.800 134.100 32.200 134.200 ;
        RECT 38.200 134.100 38.600 134.200 ;
        RECT 53.400 134.100 53.800 134.200 ;
        RECT 55.000 134.100 55.400 134.200 ;
        RECT 31.800 133.800 55.400 134.100 ;
        RECT 66.200 134.100 66.600 134.200 ;
        RECT 115.800 134.100 116.200 134.200 ;
        RECT 121.400 134.100 121.800 134.200 ;
        RECT 128.600 134.100 129.000 134.200 ;
        RECT 135.800 134.100 136.200 134.200 ;
        RECT 66.200 133.800 126.500 134.100 ;
        RECT 128.600 133.800 136.200 134.100 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 139.000 134.100 139.400 134.200 ;
        RECT 143.800 134.100 144.200 134.200 ;
        RECT 138.200 133.800 139.400 134.100 ;
        RECT 139.800 133.800 144.200 134.100 ;
        RECT 145.400 134.100 145.800 134.200 ;
        RECT 149.400 134.100 149.800 134.200 ;
        RECT 145.400 133.800 149.800 134.100 ;
        RECT 152.600 134.100 153.000 134.200 ;
        RECT 165.400 134.100 165.800 134.200 ;
        RECT 166.200 134.100 166.600 134.200 ;
        RECT 152.600 133.800 164.900 134.100 ;
        RECT 165.400 133.800 166.600 134.100 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 171.800 134.100 172.200 134.200 ;
        RECT 199.800 134.100 200.200 134.200 ;
        RECT 202.200 134.100 202.600 134.200 ;
        RECT 167.000 133.800 183.300 134.100 ;
        RECT 199.800 133.800 202.600 134.100 ;
        RECT 208.600 134.100 209.000 134.200 ;
        RECT 211.000 134.100 211.400 134.200 ;
        RECT 208.600 133.800 211.400 134.100 ;
        RECT 214.200 134.100 214.600 134.200 ;
        RECT 227.000 134.100 227.400 134.200 ;
        RECT 214.200 133.800 227.400 134.100 ;
        RECT 231.800 134.100 232.100 134.800 ;
        RECT 250.200 134.200 250.500 134.800 ;
        RECT 255.000 134.200 255.300 134.800 ;
        RECT 233.400 134.100 233.800 134.200 ;
        RECT 231.800 133.800 233.800 134.100 ;
        RECT 234.200 134.100 234.600 134.200 ;
        RECT 242.200 134.100 242.600 134.200 ;
        RECT 234.200 133.800 242.600 134.100 ;
        RECT 250.200 133.800 250.600 134.200 ;
        RECT 255.000 133.800 255.400 134.200 ;
        RECT 255.800 134.100 256.200 134.200 ;
        RECT 259.800 134.100 260.200 134.200 ;
        RECT 255.800 133.800 260.200 134.100 ;
        RECT 126.200 133.200 126.500 133.800 ;
        RECT 139.800 133.200 140.100 133.800 ;
        RECT 164.600 133.200 164.900 133.800 ;
        RECT 22.200 133.100 22.600 133.200 ;
        RECT 28.600 133.100 29.000 133.200 ;
        RECT 22.200 132.800 29.000 133.100 ;
        RECT 30.200 133.100 30.600 133.200 ;
        RECT 40.600 133.100 41.000 133.200 ;
        RECT 30.200 132.800 41.000 133.100 ;
        RECT 59.000 133.100 59.400 133.200 ;
        RECT 71.800 133.100 72.200 133.200 ;
        RECT 78.200 133.100 78.600 133.200 ;
        RECT 59.000 132.800 78.600 133.100 ;
        RECT 103.000 133.100 103.400 133.200 ;
        RECT 103.800 133.100 104.200 133.200 ;
        RECT 103.000 132.800 104.200 133.100 ;
        RECT 107.000 133.100 107.400 133.200 ;
        RECT 107.800 133.100 108.200 133.200 ;
        RECT 107.000 132.800 108.200 133.100 ;
        RECT 109.400 133.100 109.800 133.200 ;
        RECT 115.800 133.100 116.200 133.200 ;
        RECT 116.600 133.100 117.000 133.200 ;
        RECT 109.400 132.800 117.000 133.100 ;
        RECT 119.800 133.100 120.200 133.200 ;
        RECT 125.400 133.100 125.800 133.200 ;
        RECT 119.800 132.800 125.800 133.100 ;
        RECT 126.200 132.800 126.600 133.200 ;
        RECT 139.800 132.800 140.200 133.200 ;
        RECT 143.000 133.100 143.400 133.200 ;
        RECT 147.800 133.100 148.200 133.200 ;
        RECT 143.000 132.800 148.200 133.100 ;
        RECT 149.400 133.100 149.800 133.200 ;
        RECT 154.200 133.100 154.600 133.200 ;
        RECT 149.400 132.800 154.600 133.100 ;
        RECT 156.600 133.100 157.000 133.200 ;
        RECT 160.600 133.100 161.000 133.200 ;
        RECT 156.600 132.800 161.000 133.100 ;
        RECT 161.400 133.100 161.800 133.200 ;
        RECT 162.200 133.100 162.600 133.200 ;
        RECT 163.800 133.100 164.200 133.200 ;
        RECT 161.400 132.800 164.200 133.100 ;
        RECT 164.600 133.100 165.000 133.200 ;
        RECT 167.000 133.100 167.400 133.200 ;
        RECT 164.600 132.800 167.400 133.100 ;
        RECT 183.000 133.100 183.300 133.800 ;
        RECT 194.200 133.100 194.600 133.200 ;
        RECT 183.000 132.800 194.600 133.100 ;
        RECT 197.400 133.100 197.800 133.200 ;
        RECT 201.400 133.100 201.800 133.200 ;
        RECT 203.000 133.100 203.400 133.200 ;
        RECT 204.600 133.100 205.000 133.200 ;
        RECT 197.400 132.800 201.800 133.100 ;
        RECT 202.200 132.800 205.000 133.100 ;
        RECT 219.000 133.100 219.400 133.200 ;
        RECT 222.200 133.100 222.600 133.200 ;
        RECT 219.000 132.800 222.600 133.100 ;
        RECT 30.200 132.100 30.600 132.200 ;
        RECT 45.400 132.100 45.800 132.200 ;
        RECT 30.200 131.800 45.800 132.100 ;
        RECT 98.200 132.100 98.600 132.200 ;
        RECT 127.800 132.100 128.200 132.200 ;
        RECT 98.200 131.800 128.200 132.100 ;
        RECT 143.000 132.100 143.400 132.200 ;
        RECT 181.400 132.100 181.800 132.200 ;
        RECT 143.000 131.800 181.800 132.100 ;
        RECT 31.800 131.100 32.200 131.200 ;
        RECT 32.600 131.100 33.000 131.200 ;
        RECT 31.800 130.800 33.000 131.100 ;
        RECT 41.400 131.100 41.800 131.200 ;
        RECT 98.200 131.100 98.600 131.200 ;
        RECT 41.400 130.800 98.600 131.100 ;
        RECT 107.800 131.100 108.200 131.200 ;
        RECT 110.200 131.100 110.600 131.200 ;
        RECT 107.800 130.800 110.600 131.100 ;
        RECT 120.600 131.100 121.000 131.200 ;
        RECT 125.400 131.100 125.800 131.200 ;
        RECT 120.600 130.800 125.800 131.100 ;
        RECT 129.400 131.100 129.800 131.200 ;
        RECT 144.600 131.100 145.000 131.200 ;
        RECT 159.000 131.100 159.400 131.200 ;
        RECT 129.400 130.800 159.400 131.100 ;
        RECT 160.600 131.100 161.000 131.200 ;
        RECT 167.000 131.100 167.400 131.200 ;
        RECT 160.600 130.800 167.400 131.100 ;
        RECT 175.800 131.100 176.200 131.200 ;
        RECT 176.600 131.100 177.000 131.200 ;
        RECT 175.800 130.800 177.000 131.100 ;
        RECT 180.600 131.100 181.000 131.200 ;
        RECT 187.000 131.100 187.400 131.200 ;
        RECT 180.600 130.800 187.400 131.100 ;
        RECT 190.200 131.100 190.600 131.200 ;
        RECT 199.800 131.100 200.200 131.200 ;
        RECT 190.200 130.800 200.200 131.100 ;
        RECT 203.000 131.100 203.400 131.200 ;
        RECT 207.000 131.100 207.400 131.200 ;
        RECT 203.000 130.800 207.400 131.100 ;
        RECT 21.400 130.100 21.800 130.200 ;
        RECT 38.200 130.100 38.600 130.200 ;
        RECT 21.400 129.800 38.600 130.100 ;
        RECT 42.200 130.100 42.600 130.200 ;
        RECT 44.600 130.100 45.000 130.200 ;
        RECT 70.200 130.100 70.600 130.200 ;
        RECT 42.200 129.800 70.600 130.100 ;
        RECT 72.600 130.100 73.000 130.200 ;
        RECT 90.200 130.100 90.600 130.200 ;
        RECT 72.600 129.800 90.600 130.100 ;
        RECT 103.000 130.100 103.400 130.200 ;
        RECT 103.800 130.100 104.200 130.200 ;
        RECT 103.000 129.800 104.200 130.100 ;
        RECT 109.400 130.100 109.800 130.200 ;
        RECT 119.800 130.100 120.200 130.200 ;
        RECT 109.400 129.800 120.200 130.100 ;
        RECT 157.400 130.100 157.800 130.200 ;
        RECT 164.600 130.100 165.000 130.200 ;
        RECT 157.400 129.800 165.000 130.100 ;
        RECT 17.400 129.100 17.800 129.200 ;
        RECT 19.000 129.100 19.400 129.200 ;
        RECT 16.600 128.800 19.400 129.100 ;
        RECT 24.600 129.100 25.000 129.200 ;
        RECT 29.400 129.100 29.800 129.200 ;
        RECT 24.600 128.800 29.800 129.100 ;
        RECT 30.200 128.800 30.600 129.200 ;
        RECT 31.000 129.100 31.400 129.200 ;
        RECT 47.000 129.100 47.400 129.200 ;
        RECT 55.800 129.100 56.200 129.200 ;
        RECT 67.000 129.100 67.400 129.200 ;
        RECT 31.000 128.800 67.400 129.100 ;
        RECT 68.600 129.100 69.000 129.200 ;
        RECT 71.800 129.100 72.200 129.200 ;
        RECT 101.400 129.100 101.800 129.200 ;
        RECT 102.200 129.100 102.600 129.200 ;
        RECT 103.800 129.100 104.200 129.200 ;
        RECT 131.000 129.100 131.400 129.200 ;
        RECT 68.600 128.800 102.600 129.100 ;
        RECT 103.000 128.800 131.400 129.100 ;
        RECT 141.400 129.100 141.800 129.200 ;
        RECT 146.200 129.100 146.600 129.200 ;
        RECT 147.800 129.100 148.200 129.200 ;
        RECT 155.000 129.100 155.400 129.200 ;
        RECT 141.400 128.800 148.200 129.100 ;
        RECT 153.400 128.800 155.400 129.100 ;
        RECT 158.200 129.100 158.600 129.200 ;
        RECT 163.000 129.100 163.400 129.200 ;
        RECT 158.200 128.800 163.400 129.100 ;
        RECT 165.400 129.100 165.800 129.200 ;
        RECT 170.200 129.100 170.600 129.200 ;
        RECT 165.400 128.800 170.600 129.100 ;
        RECT 171.800 129.100 172.200 129.200 ;
        RECT 182.200 129.100 182.600 129.200 ;
        RECT 171.800 128.800 182.600 129.100 ;
        RECT 209.400 129.100 209.800 129.200 ;
        RECT 210.200 129.100 210.600 129.200 ;
        RECT 209.400 128.800 210.600 129.100 ;
        RECT 223.000 129.100 223.400 129.200 ;
        RECT 223.800 129.100 224.200 129.200 ;
        RECT 223.000 128.800 224.200 129.100 ;
        RECT 226.200 129.100 226.600 129.200 ;
        RECT 257.400 129.100 257.800 129.200 ;
        RECT 262.200 129.100 262.600 129.200 ;
        RECT 226.200 128.800 250.500 129.100 ;
        RECT 257.400 128.800 262.600 129.100 ;
        RECT 30.200 128.200 30.500 128.800 ;
        RECT 15.000 128.100 15.400 128.200 ;
        RECT 17.400 128.100 17.800 128.200 ;
        RECT 22.200 128.100 22.600 128.200 ;
        RECT 26.200 128.100 26.600 128.200 ;
        RECT 15.000 127.800 26.600 128.100 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 36.600 128.100 37.000 128.200 ;
        RECT 42.200 128.100 42.600 128.200 ;
        RECT 36.600 127.800 42.600 128.100 ;
        RECT 44.600 128.100 45.000 128.200 ;
        RECT 45.400 128.100 45.800 128.200 ;
        RECT 44.600 127.800 45.800 128.100 ;
        RECT 55.000 128.100 55.400 128.200 ;
        RECT 63.000 128.100 63.400 128.200 ;
        RECT 55.000 127.800 63.400 128.100 ;
        RECT 67.000 127.800 67.400 128.200 ;
        RECT 71.800 128.100 72.200 128.200 ;
        RECT 72.600 128.100 73.000 128.200 ;
        RECT 71.800 127.800 73.000 128.100 ;
        RECT 78.200 128.100 78.600 128.200 ;
        RECT 80.600 128.100 81.000 128.200 ;
        RECT 82.200 128.100 82.600 128.200 ;
        RECT 78.200 127.800 82.600 128.100 ;
        RECT 84.600 128.100 85.000 128.200 ;
        RECT 86.200 128.100 86.600 128.200 ;
        RECT 87.800 128.100 88.200 128.200 ;
        RECT 84.600 127.800 88.200 128.100 ;
        RECT 92.600 128.100 93.000 128.200 ;
        RECT 115.000 128.100 115.400 128.200 ;
        RECT 92.600 127.800 115.400 128.100 ;
        RECT 127.800 128.100 128.200 128.200 ;
        RECT 132.600 128.100 133.000 128.200 ;
        RECT 127.800 127.800 133.000 128.100 ;
        RECT 142.200 128.100 142.600 128.200 ;
        RECT 144.600 128.100 145.000 128.200 ;
        RECT 142.200 127.800 145.000 128.100 ;
        RECT 145.400 128.100 145.800 128.200 ;
        RECT 153.400 128.100 153.700 128.800 ;
        RECT 250.200 128.200 250.500 128.800 ;
        RECT 145.400 127.800 153.700 128.100 ;
        RECT 154.200 128.100 154.600 128.200 ;
        RECT 169.400 128.100 169.800 128.200 ;
        RECT 154.200 127.800 169.800 128.100 ;
        RECT 171.000 128.100 171.400 128.200 ;
        RECT 180.600 128.100 181.000 128.200 ;
        RECT 194.200 128.100 194.600 128.200 ;
        RECT 202.200 128.100 202.600 128.200 ;
        RECT 171.000 127.800 181.000 128.100 ;
        RECT 190.200 127.800 202.600 128.100 ;
        RECT 230.200 127.800 230.600 128.200 ;
        RECT 232.600 128.100 233.000 128.200 ;
        RECT 237.400 128.100 237.800 128.200 ;
        RECT 232.600 127.800 237.800 128.100 ;
        RECT 239.800 127.800 240.200 128.200 ;
        RECT 250.200 127.800 250.600 128.200 ;
        RECT 18.200 127.100 18.600 127.200 ;
        RECT 23.000 127.100 23.400 127.200 ;
        RECT 18.200 126.800 23.400 127.100 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 38.200 127.100 38.600 127.200 ;
        RECT 39.000 127.100 39.400 127.200 ;
        RECT 40.600 127.100 41.000 127.200 ;
        RECT 38.200 126.800 41.000 127.100 ;
        RECT 42.200 127.100 42.600 127.200 ;
        RECT 50.200 127.100 50.600 127.200 ;
        RECT 42.200 126.800 50.600 127.100 ;
        RECT 54.200 127.100 54.600 127.200 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 54.200 126.800 65.800 127.100 ;
        RECT 67.000 127.100 67.300 127.800 ;
        RECT 86.200 127.100 86.600 127.200 ;
        RECT 88.600 127.100 89.000 127.200 ;
        RECT 67.000 126.800 85.700 127.100 ;
        RECT 86.200 126.800 89.000 127.100 ;
        RECT 103.800 127.100 104.200 127.200 ;
        RECT 104.600 127.100 105.000 127.200 ;
        RECT 103.800 126.800 105.000 127.100 ;
        RECT 111.000 127.100 111.400 127.200 ;
        RECT 111.800 127.100 112.200 127.200 ;
        RECT 111.000 126.800 112.200 127.100 ;
        RECT 117.400 127.100 117.800 127.200 ;
        RECT 130.200 127.100 130.600 127.200 ;
        RECT 117.400 126.800 130.600 127.100 ;
        RECT 132.600 127.100 133.000 127.200 ;
        RECT 150.200 127.100 150.600 127.200 ;
        RECT 132.600 126.800 150.600 127.100 ;
        RECT 151.800 127.100 152.200 127.200 ;
        RECT 157.400 127.100 157.800 127.200 ;
        RECT 151.800 126.800 157.800 127.100 ;
        RECT 159.800 127.100 160.200 127.200 ;
        RECT 164.600 127.100 165.000 127.200 ;
        RECT 159.800 126.800 165.000 127.100 ;
        RECT 165.400 126.800 165.800 127.200 ;
        RECT 183.800 126.800 184.200 127.200 ;
        RECT 184.600 127.100 185.000 127.200 ;
        RECT 190.200 127.100 190.500 127.800 ;
        RECT 230.200 127.200 230.500 127.800 ;
        RECT 239.800 127.200 240.100 127.800 ;
        RECT 184.600 126.800 190.500 127.100 ;
        RECT 191.000 126.800 191.400 127.200 ;
        RECT 199.800 127.100 200.200 127.200 ;
        RECT 200.600 127.100 201.000 127.200 ;
        RECT 199.800 126.800 201.000 127.100 ;
        RECT 230.200 126.800 230.600 127.200 ;
        RECT 239.800 126.800 240.200 127.200 ;
        RECT 249.400 127.100 249.800 127.200 ;
        RECT 259.800 127.100 260.200 127.200 ;
        RECT 249.400 126.800 260.200 127.100 ;
        RECT 11.800 126.100 12.200 126.200 ;
        RECT 19.000 126.100 19.400 126.200 ;
        RECT 11.800 125.800 19.400 126.100 ;
        RECT 27.000 126.100 27.300 126.800 ;
        RECT 85.400 126.200 85.700 126.800 ;
        RECT 31.000 126.100 31.400 126.200 ;
        RECT 27.000 125.800 31.400 126.100 ;
        RECT 32.600 126.100 33.000 126.200 ;
        RECT 39.800 126.100 40.200 126.200 ;
        RECT 32.600 125.800 40.200 126.100 ;
        RECT 43.800 126.100 44.200 126.200 ;
        RECT 67.800 126.100 68.200 126.200 ;
        RECT 43.800 125.800 68.200 126.100 ;
        RECT 78.200 126.100 78.600 126.200 ;
        RECT 79.000 126.100 79.400 126.200 ;
        RECT 84.600 126.100 85.000 126.200 ;
        RECT 78.200 125.800 85.000 126.100 ;
        RECT 85.400 125.800 85.800 126.200 ;
        RECT 87.000 126.100 87.400 126.200 ;
        RECT 89.400 126.100 89.800 126.200 ;
        RECT 87.000 125.800 89.800 126.100 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 117.400 126.100 117.800 126.200 ;
        RECT 118.200 126.100 118.600 126.200 ;
        RECT 117.400 125.800 118.600 126.100 ;
        RECT 119.800 126.100 120.200 126.200 ;
        RECT 135.800 126.100 136.200 126.200 ;
        RECT 143.800 126.100 144.200 126.200 ;
        RECT 119.800 125.800 129.700 126.100 ;
        RECT 135.800 125.800 144.200 126.100 ;
        RECT 146.200 126.100 146.600 126.200 ;
        RECT 147.800 126.100 148.200 126.200 ;
        RECT 158.200 126.100 158.600 126.200 ;
        RECT 146.200 125.800 158.600 126.100 ;
        RECT 163.800 126.100 164.200 126.200 ;
        RECT 165.400 126.100 165.700 126.800 ;
        RECT 163.800 125.800 165.700 126.100 ;
        RECT 167.800 126.100 168.200 126.200 ;
        RECT 171.800 126.100 172.200 126.200 ;
        RECT 167.800 125.800 172.200 126.100 ;
        RECT 178.200 125.800 178.600 126.200 ;
        RECT 180.600 126.100 181.000 126.200 ;
        RECT 183.800 126.100 184.100 126.800 ;
        RECT 180.600 125.800 184.100 126.100 ;
        RECT 191.000 126.100 191.300 126.800 ;
        RECT 195.800 126.100 196.200 126.200 ;
        RECT 191.000 125.800 196.200 126.100 ;
        RECT 204.600 126.100 205.000 126.200 ;
        RECT 205.400 126.100 205.800 126.200 ;
        RECT 204.600 125.800 205.800 126.100 ;
        RECT 206.200 125.800 206.600 126.200 ;
        RECT 211.000 126.100 211.400 126.200 ;
        RECT 211.800 126.100 212.200 126.200 ;
        RECT 211.000 125.800 212.200 126.100 ;
        RECT 213.400 126.100 213.800 126.200 ;
        RECT 236.600 126.100 237.000 126.200 ;
        RECT 213.400 125.800 237.000 126.100 ;
        RECT 247.800 126.100 248.200 126.200 ;
        RECT 255.000 126.100 255.400 126.200 ;
        RECT 247.800 125.800 255.400 126.100 ;
        RECT 87.000 125.200 87.300 125.800 ;
        RECT 19.800 125.100 20.200 125.200 ;
        RECT 21.400 125.100 21.800 125.200 ;
        RECT 19.800 124.800 21.800 125.100 ;
        RECT 32.600 125.100 33.000 125.200 ;
        RECT 47.800 125.100 48.200 125.200 ;
        RECT 52.600 125.100 53.000 125.200 ;
        RECT 32.600 124.800 48.200 125.100 ;
        RECT 48.600 124.800 53.000 125.100 ;
        RECT 53.400 125.100 53.800 125.200 ;
        RECT 59.800 125.100 60.200 125.200 ;
        RECT 61.400 125.100 61.800 125.200 ;
        RECT 53.400 124.800 61.800 125.100 ;
        RECT 65.400 125.100 65.800 125.200 ;
        RECT 66.200 125.100 66.600 125.200 ;
        RECT 65.400 124.800 66.600 125.100 ;
        RECT 74.200 125.100 74.600 125.200 ;
        RECT 86.200 125.100 86.600 125.200 ;
        RECT 74.200 124.800 86.600 125.100 ;
        RECT 87.000 124.800 87.400 125.200 ;
        RECT 105.400 125.100 105.800 125.200 ;
        RECT 107.800 125.100 108.200 125.200 ;
        RECT 105.400 124.800 108.200 125.100 ;
        RECT 108.600 125.100 109.000 125.200 ;
        RECT 109.400 125.100 109.800 125.200 ;
        RECT 108.600 124.800 109.800 125.100 ;
        RECT 113.400 125.100 113.700 125.800 ;
        RECT 129.400 125.200 129.700 125.800 ;
        RECT 115.800 125.100 116.200 125.200 ;
        RECT 113.400 124.800 116.200 125.100 ;
        RECT 118.200 124.800 118.600 125.200 ;
        RECT 119.800 125.100 120.200 125.200 ;
        RECT 120.600 125.100 121.000 125.200 ;
        RECT 127.800 125.100 128.200 125.200 ;
        RECT 119.800 124.800 128.200 125.100 ;
        RECT 129.400 124.800 129.800 125.200 ;
        RECT 144.600 125.100 145.000 125.200 ;
        RECT 154.200 125.100 154.600 125.200 ;
        RECT 144.600 124.800 154.600 125.100 ;
        RECT 167.800 125.100 168.200 125.200 ;
        RECT 168.600 125.100 169.000 125.200 ;
        RECT 167.800 124.800 169.000 125.100 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 178.200 125.100 178.500 125.800 ;
        RECT 206.200 125.200 206.500 125.800 ;
        RECT 196.600 125.100 197.000 125.200 ;
        RECT 206.200 125.100 206.600 125.200 ;
        RECT 171.000 124.800 206.600 125.100 ;
        RECT 211.800 125.100 212.100 125.800 ;
        RECT 218.200 125.100 218.600 125.200 ;
        RECT 211.800 124.800 218.600 125.100 ;
        RECT 237.400 125.100 237.800 125.200 ;
        RECT 243.800 125.100 244.200 125.200 ;
        RECT 237.400 124.800 244.200 125.100 ;
        RECT 245.400 125.100 245.800 125.200 ;
        RECT 247.000 125.100 247.400 125.200 ;
        RECT 245.400 124.800 247.400 125.100 ;
        RECT 48.600 124.200 48.900 124.800 ;
        RECT 47.800 124.100 48.200 124.200 ;
        RECT 45.400 123.800 48.200 124.100 ;
        RECT 48.600 123.800 49.000 124.200 ;
        RECT 64.600 124.100 65.000 124.200 ;
        RECT 67.000 124.100 67.400 124.200 ;
        RECT 79.800 124.100 80.200 124.200 ;
        RECT 83.800 124.100 84.200 124.200 ;
        RECT 116.600 124.100 117.000 124.200 ;
        RECT 118.200 124.100 118.500 124.800 ;
        RECT 247.000 124.200 247.300 124.800 ;
        RECT 64.600 123.800 118.500 124.100 ;
        RECT 131.000 124.100 131.400 124.200 ;
        RECT 143.000 124.100 143.400 124.200 ;
        RECT 131.000 123.800 143.400 124.100 ;
        RECT 144.600 124.100 145.000 124.200 ;
        RECT 159.800 124.100 160.200 124.200 ;
        RECT 144.600 123.800 160.200 124.100 ;
        RECT 176.600 124.100 177.000 124.200 ;
        RECT 185.400 124.100 185.800 124.200 ;
        RECT 176.600 123.800 185.800 124.100 ;
        RECT 199.000 124.100 199.400 124.200 ;
        RECT 206.200 124.100 206.600 124.200 ;
        RECT 199.000 123.800 206.600 124.100 ;
        RECT 231.800 124.100 232.200 124.200 ;
        RECT 233.400 124.100 233.800 124.200 ;
        RECT 244.600 124.100 245.000 124.200 ;
        RECT 231.800 123.800 245.000 124.100 ;
        RECT 247.000 123.800 247.400 124.200 ;
        RECT 45.400 123.200 45.700 123.800 ;
        RECT 45.400 122.800 45.800 123.200 ;
        RECT 46.200 123.100 46.600 123.200 ;
        RECT 58.200 123.100 58.600 123.200 ;
        RECT 64.600 123.100 65.000 123.200 ;
        RECT 73.400 123.100 73.800 123.200 ;
        RECT 109.400 123.100 109.800 123.200 ;
        RECT 46.200 122.800 109.800 123.100 ;
        RECT 110.200 123.100 110.600 123.200 ;
        RECT 114.200 123.100 114.600 123.200 ;
        RECT 119.000 123.100 119.400 123.200 ;
        RECT 125.400 123.100 125.800 123.200 ;
        RECT 147.000 123.100 147.400 123.200 ;
        RECT 110.200 122.800 147.400 123.100 ;
        RECT 160.600 123.100 161.000 123.200 ;
        RECT 166.200 123.100 166.600 123.200 ;
        RECT 160.600 122.800 166.600 123.100 ;
        RECT 171.000 123.100 171.400 123.200 ;
        RECT 221.400 123.100 221.800 123.200 ;
        RECT 244.600 123.100 245.000 123.200 ;
        RECT 247.000 123.100 247.400 123.200 ;
        RECT 171.000 122.800 247.400 123.100 ;
        RECT 47.000 122.100 47.400 122.200 ;
        RECT 65.400 122.100 65.800 122.200 ;
        RECT 47.000 121.800 65.800 122.100 ;
        RECT 72.600 122.100 73.000 122.200 ;
        RECT 79.000 122.100 79.400 122.200 ;
        RECT 84.600 122.100 85.000 122.200 ;
        RECT 89.400 122.100 89.800 122.200 ;
        RECT 113.400 122.100 113.800 122.200 ;
        RECT 135.000 122.100 135.400 122.200 ;
        RECT 160.600 122.100 160.900 122.800 ;
        RECT 72.600 121.800 80.100 122.100 ;
        RECT 84.600 121.800 89.800 122.100 ;
        RECT 112.600 121.800 135.400 122.100 ;
        RECT 135.800 121.800 160.900 122.100 ;
        RECT 185.400 122.100 185.800 122.200 ;
        RECT 235.000 122.100 235.400 122.200 ;
        RECT 238.200 122.100 238.600 122.200 ;
        RECT 185.400 121.800 238.600 122.100 ;
        RECT 79.800 121.100 80.200 121.200 ;
        RECT 88.600 121.100 89.000 121.200 ;
        RECT 79.800 120.800 89.000 121.100 ;
        RECT 89.400 121.100 89.800 121.200 ;
        RECT 91.800 121.100 92.200 121.200 ;
        RECT 89.400 120.800 92.200 121.100 ;
        RECT 92.600 121.100 93.000 121.200 ;
        RECT 108.600 121.100 109.000 121.200 ;
        RECT 135.800 121.100 136.100 121.800 ;
        RECT 92.600 120.800 136.100 121.100 ;
        RECT 182.200 121.100 182.600 121.200 ;
        RECT 187.800 121.100 188.200 121.200 ;
        RECT 182.200 120.800 188.200 121.100 ;
        RECT 199.000 121.100 199.400 121.200 ;
        RECT 202.200 121.100 202.600 121.200 ;
        RECT 225.400 121.100 225.800 121.200 ;
        RECT 199.000 120.800 225.800 121.100 ;
        RECT 243.000 121.100 243.400 121.200 ;
        RECT 248.600 121.100 249.000 121.200 ;
        RECT 243.000 120.800 249.000 121.100 ;
        RECT 85.400 120.100 85.800 120.200 ;
        RECT 97.400 120.100 97.800 120.200 ;
        RECT 85.400 119.800 97.800 120.100 ;
        RECT 193.400 120.100 193.800 120.200 ;
        RECT 209.400 120.100 209.800 120.200 ;
        RECT 193.400 119.800 209.800 120.100 ;
        RECT 211.800 120.100 212.200 120.200 ;
        RECT 231.000 120.100 231.400 120.200 ;
        RECT 211.800 119.800 231.400 120.100 ;
        RECT 246.200 119.800 246.600 120.200 ;
        RECT 47.000 118.800 47.400 119.200 ;
        RECT 133.400 119.100 133.800 119.200 ;
        RECT 136.600 119.100 137.000 119.200 ;
        RECT 133.400 118.800 137.000 119.100 ;
        RECT 143.000 119.100 143.400 119.200 ;
        RECT 147.800 119.100 148.200 119.200 ;
        RECT 143.000 118.800 148.200 119.100 ;
        RECT 215.000 119.100 215.400 119.200 ;
        RECT 231.800 119.100 232.200 119.200 ;
        RECT 215.000 118.800 232.200 119.100 ;
        RECT 239.000 118.800 239.400 119.200 ;
        RECT 246.200 119.100 246.500 119.800 ;
        RECT 249.400 119.100 249.800 119.200 ;
        RECT 246.200 118.800 249.800 119.100 ;
        RECT 263.000 119.100 263.400 119.200 ;
        RECT 263.800 119.100 264.200 119.200 ;
        RECT 263.000 118.800 264.200 119.100 ;
        RECT 47.000 118.200 47.300 118.800 ;
        RECT 35.800 117.800 36.200 118.200 ;
        RECT 47.000 117.800 47.400 118.200 ;
        RECT 50.200 118.100 50.600 118.200 ;
        RECT 51.800 118.100 52.200 118.200 ;
        RECT 50.200 117.800 52.200 118.100 ;
        RECT 59.000 118.100 59.400 118.200 ;
        RECT 63.800 118.100 64.200 118.200 ;
        RECT 59.000 117.800 64.200 118.100 ;
        RECT 84.600 118.100 85.000 118.200 ;
        RECT 126.200 118.100 126.600 118.200 ;
        RECT 146.200 118.100 146.600 118.200 ;
        RECT 84.600 117.800 146.600 118.100 ;
        RECT 149.400 118.100 149.800 118.200 ;
        RECT 154.200 118.100 154.600 118.200 ;
        RECT 149.400 117.800 154.600 118.100 ;
        RECT 208.600 118.100 209.000 118.200 ;
        RECT 237.400 118.100 237.800 118.200 ;
        RECT 239.000 118.100 239.300 118.800 ;
        RECT 208.600 117.800 239.300 118.100 ;
        RECT 242.200 118.100 242.600 118.200 ;
        RECT 247.800 118.100 248.200 118.200 ;
        RECT 242.200 117.800 248.200 118.100 ;
        RECT 35.800 117.200 36.100 117.800 ;
        RECT 11.800 117.100 12.200 117.200 ;
        RECT 19.000 117.100 19.400 117.200 ;
        RECT 11.800 116.800 19.400 117.100 ;
        RECT 35.800 116.800 36.200 117.200 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 86.200 117.100 86.600 117.200 ;
        RECT 43.000 116.800 86.600 117.100 ;
        RECT 87.800 116.800 88.200 117.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 134.200 117.100 134.600 117.200 ;
        RECT 135.000 117.100 135.400 117.200 ;
        RECT 134.200 116.800 135.400 117.100 ;
        RECT 136.600 117.100 137.000 117.200 ;
        RECT 143.800 117.100 144.200 117.200 ;
        RECT 151.800 117.100 152.200 117.200 ;
        RECT 136.600 116.800 152.200 117.100 ;
        RECT 155.800 117.100 156.200 117.200 ;
        RECT 162.200 117.100 162.600 117.200 ;
        RECT 155.800 116.800 162.600 117.100 ;
        RECT 191.800 116.800 192.200 117.200 ;
        RECT 205.400 117.100 205.800 117.200 ;
        RECT 243.800 117.100 244.200 117.200 ;
        RECT 205.400 116.800 244.200 117.100 ;
        RECT 245.400 116.800 245.800 117.200 ;
        RECT 255.800 117.100 256.200 117.200 ;
        RECT 256.600 117.100 257.000 117.200 ;
        RECT 255.800 116.800 257.000 117.100 ;
        RECT 87.800 116.200 88.100 116.800 ;
        RECT 124.600 116.200 124.900 116.800 ;
        RECT 191.800 116.200 192.100 116.800 ;
        RECT 18.200 116.100 18.600 116.200 ;
        RECT 21.400 116.100 21.800 116.200 ;
        RECT 46.200 116.100 46.600 116.200 ;
        RECT 18.200 115.800 46.600 116.100 ;
        RECT 47.000 116.100 47.400 116.200 ;
        RECT 63.800 116.100 64.200 116.200 ;
        RECT 70.200 116.100 70.600 116.200 ;
        RECT 74.200 116.100 74.600 116.200 ;
        RECT 47.000 115.800 74.600 116.100 ;
        RECT 85.400 116.100 85.800 116.200 ;
        RECT 87.800 116.100 88.200 116.200 ;
        RECT 85.400 115.800 88.200 116.100 ;
        RECT 90.200 116.100 90.600 116.200 ;
        RECT 103.000 116.100 103.400 116.200 ;
        RECT 90.200 115.800 103.400 116.100 ;
        RECT 124.600 115.800 125.000 116.200 ;
        RECT 129.400 115.800 129.800 116.200 ;
        RECT 132.600 116.100 133.000 116.200 ;
        RECT 139.800 116.100 140.200 116.200 ;
        RECT 132.600 115.800 140.200 116.100 ;
        RECT 148.600 116.100 149.000 116.200 ;
        RECT 156.600 116.100 157.000 116.200 ;
        RECT 159.000 116.100 159.400 116.200 ;
        RECT 161.400 116.100 161.800 116.200 ;
        RECT 148.600 115.800 161.800 116.100 ;
        RECT 191.800 115.800 192.200 116.200 ;
        RECT 207.800 116.100 208.200 116.200 ;
        RECT 215.000 116.100 215.400 116.200 ;
        RECT 207.800 115.800 215.400 116.100 ;
        RECT 227.000 116.100 227.400 116.200 ;
        RECT 231.000 116.100 231.400 116.200 ;
        RECT 232.600 116.100 233.000 116.200 ;
        RECT 227.000 115.800 233.000 116.100 ;
        RECT 245.400 116.100 245.700 116.800 ;
        RECT 251.800 116.100 252.200 116.200 ;
        RECT 245.400 115.800 252.200 116.100 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 22.200 115.100 22.600 115.200 ;
        RECT 24.600 115.100 25.000 115.200 ;
        RECT 16.600 114.800 25.000 115.100 ;
        RECT 34.200 115.100 34.600 115.200 ;
        RECT 40.600 115.100 41.000 115.200 ;
        RECT 47.800 115.100 48.200 115.200 ;
        RECT 34.200 114.800 37.700 115.100 ;
        RECT 40.600 114.800 48.200 115.100 ;
        RECT 53.400 115.100 53.800 115.200 ;
        RECT 55.000 115.100 55.400 115.200 ;
        RECT 65.400 115.100 65.800 115.200 ;
        RECT 74.200 115.100 74.600 115.200 ;
        RECT 77.400 115.100 77.800 115.200 ;
        RECT 53.400 114.800 55.400 115.100 ;
        RECT 64.600 114.800 71.300 115.100 ;
        RECT 74.200 114.800 77.800 115.100 ;
        RECT 88.600 115.100 89.000 115.200 ;
        RECT 92.600 115.100 93.000 115.200 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 88.600 114.800 93.000 115.100 ;
        RECT 101.400 114.800 105.000 115.100 ;
        RECT 119.800 115.100 120.200 115.200 ;
        RECT 127.800 115.100 128.200 115.200 ;
        RECT 119.800 114.800 128.200 115.100 ;
        RECT 129.400 115.100 129.700 115.800 ;
        RECT 130.200 115.100 130.600 115.200 ;
        RECT 131.800 115.100 132.200 115.200 ;
        RECT 129.400 114.800 132.200 115.100 ;
        RECT 132.600 115.100 133.000 115.200 ;
        RECT 137.400 115.100 137.800 115.200 ;
        RECT 132.600 114.800 137.800 115.100 ;
        RECT 148.600 115.100 149.000 115.200 ;
        RECT 149.400 115.100 149.800 115.200 ;
        RECT 148.600 114.800 149.800 115.100 ;
        RECT 150.200 115.100 150.600 115.200 ;
        RECT 202.200 115.100 202.600 115.200 ;
        RECT 203.000 115.100 203.400 115.200 ;
        RECT 150.200 114.800 203.400 115.100 ;
        RECT 211.800 115.100 212.200 115.200 ;
        RECT 214.200 115.100 214.600 115.200 ;
        RECT 217.400 115.100 217.800 115.200 ;
        RECT 211.800 114.800 217.800 115.100 ;
        RECT 223.000 115.100 223.400 115.200 ;
        RECT 230.200 115.100 230.600 115.200 ;
        RECT 223.000 114.800 230.600 115.100 ;
        RECT 258.200 115.100 258.600 115.200 ;
        RECT 258.200 114.800 259.400 115.100 ;
        RECT 37.400 114.200 37.700 114.800 ;
        RECT 71.000 114.200 71.300 114.800 ;
        RECT 101.400 114.200 101.700 114.800 ;
        RECT 259.000 114.700 259.400 114.800 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 27.800 114.100 28.200 114.200 ;
        RECT 17.400 113.800 28.200 114.100 ;
        RECT 29.400 114.100 29.800 114.200 ;
        RECT 33.400 114.100 33.800 114.200 ;
        RECT 29.400 113.800 33.800 114.100 ;
        RECT 37.400 114.100 37.800 114.200 ;
        RECT 39.000 114.100 39.400 114.200 ;
        RECT 37.400 113.800 39.400 114.100 ;
        RECT 51.000 114.100 51.400 114.200 ;
        RECT 68.600 114.100 69.000 114.200 ;
        RECT 69.400 114.100 69.800 114.200 ;
        RECT 51.000 113.800 60.900 114.100 ;
        RECT 68.600 113.800 69.800 114.100 ;
        RECT 71.000 113.800 71.400 114.200 ;
        RECT 73.400 114.100 73.800 114.200 ;
        RECT 75.800 114.100 76.200 114.200 ;
        RECT 73.400 113.800 76.200 114.100 ;
        RECT 82.200 114.100 82.600 114.200 ;
        RECT 91.000 114.100 91.400 114.200 ;
        RECT 82.200 113.800 91.400 114.100 ;
        RECT 101.400 113.800 101.800 114.200 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 127.800 114.100 128.200 114.200 ;
        RECT 141.400 114.100 141.800 114.200 ;
        RECT 125.400 113.800 141.800 114.100 ;
        RECT 143.800 113.800 144.200 114.200 ;
        RECT 144.600 114.100 145.000 114.200 ;
        RECT 147.000 114.100 147.400 114.200 ;
        RECT 144.600 113.800 147.400 114.100 ;
        RECT 159.800 114.100 160.200 114.200 ;
        RECT 167.800 114.100 168.200 114.200 ;
        RECT 159.800 113.800 168.200 114.100 ;
        RECT 201.400 114.100 201.800 114.200 ;
        RECT 203.800 114.100 204.200 114.200 ;
        RECT 201.400 113.800 204.200 114.100 ;
        RECT 205.400 114.100 205.800 114.200 ;
        RECT 213.400 114.100 213.800 114.200 ;
        RECT 205.400 113.800 213.800 114.100 ;
        RECT 218.200 114.100 218.600 114.200 ;
        RECT 232.600 114.100 233.000 114.200 ;
        RECT 218.200 113.800 233.000 114.100 ;
        RECT 235.800 113.800 236.200 114.200 ;
        RECT 236.600 113.800 237.000 114.200 ;
        RECT 263.800 114.100 264.200 114.200 ;
        RECT 254.200 113.800 264.200 114.100 ;
        RECT 60.600 113.200 60.900 113.800 ;
        RECT 143.800 113.200 144.100 113.800 ;
        RECT 18.200 113.100 18.600 113.200 ;
        RECT 19.800 113.100 20.200 113.200 ;
        RECT 18.200 112.800 20.200 113.100 ;
        RECT 23.000 112.800 23.400 113.200 ;
        RECT 27.000 113.100 27.400 113.200 ;
        RECT 28.600 113.100 29.000 113.200 ;
        RECT 30.200 113.100 30.600 113.200 ;
        RECT 27.000 112.800 30.600 113.100 ;
        RECT 31.800 113.100 32.200 113.200 ;
        RECT 36.600 113.100 37.000 113.200 ;
        RECT 31.800 112.800 37.000 113.100 ;
        RECT 60.600 112.800 61.000 113.200 ;
        RECT 68.600 113.100 69.000 113.200 ;
        RECT 72.600 113.100 73.000 113.200 ;
        RECT 68.600 112.800 73.000 113.100 ;
        RECT 75.000 113.100 75.400 113.200 ;
        RECT 79.000 113.100 79.400 113.200 ;
        RECT 91.000 113.100 91.400 113.200 ;
        RECT 75.000 112.800 91.400 113.100 ;
        RECT 110.200 113.100 110.600 113.200 ;
        RECT 139.800 113.100 140.200 113.200 ;
        RECT 110.200 112.800 140.200 113.100 ;
        RECT 142.200 113.100 142.600 113.200 ;
        RECT 143.800 113.100 144.200 113.200 ;
        RECT 142.200 112.800 144.200 113.100 ;
        RECT 147.000 113.100 147.400 113.200 ;
        RECT 187.800 113.100 188.200 113.200 ;
        RECT 147.000 112.800 188.200 113.100 ;
        RECT 195.000 113.100 195.400 113.200 ;
        RECT 235.800 113.100 236.100 113.800 ;
        RECT 195.000 112.800 236.100 113.100 ;
        RECT 236.600 113.100 236.900 113.800 ;
        RECT 254.200 113.200 254.500 113.800 ;
        RECT 241.400 113.100 241.800 113.200 ;
        RECT 236.600 112.800 241.800 113.100 ;
        RECT 254.200 112.800 254.600 113.200 ;
        RECT 23.000 112.200 23.300 112.800 ;
        RECT 23.000 111.800 23.400 112.200 ;
        RECT 24.600 112.100 25.000 112.200 ;
        RECT 39.800 112.100 40.200 112.200 ;
        RECT 43.000 112.100 43.400 112.200 ;
        RECT 91.800 112.100 92.200 112.200 ;
        RECT 24.600 111.800 29.700 112.100 ;
        RECT 39.800 111.800 92.200 112.100 ;
        RECT 92.600 112.100 93.000 112.200 ;
        RECT 143.800 112.100 144.200 112.200 ;
        RECT 92.600 111.800 144.200 112.100 ;
        RECT 150.200 112.100 150.600 112.200 ;
        RECT 187.000 112.100 187.400 112.200 ;
        RECT 150.200 111.800 187.400 112.100 ;
        RECT 187.800 112.100 188.100 112.800 ;
        RECT 210.200 112.100 210.600 112.200 ;
        RECT 235.000 112.100 235.400 112.200 ;
        RECT 187.800 111.800 235.400 112.100 ;
        RECT 245.400 112.100 245.800 112.200 ;
        RECT 257.400 112.100 257.800 112.200 ;
        RECT 245.400 111.800 257.800 112.100 ;
        RECT 29.400 111.200 29.700 111.800 ;
        RECT 29.400 110.800 29.800 111.200 ;
        RECT 33.400 111.100 33.800 111.200 ;
        RECT 42.200 111.100 42.600 111.200 ;
        RECT 51.800 111.100 52.200 111.200 ;
        RECT 53.400 111.100 53.800 111.200 ;
        RECT 33.400 110.800 53.800 111.100 ;
        RECT 54.200 111.100 54.600 111.200 ;
        RECT 62.200 111.100 62.600 111.200 ;
        RECT 54.200 110.800 62.600 111.100 ;
        RECT 67.800 111.100 68.200 111.200 ;
        RECT 78.200 111.100 78.600 111.200 ;
        RECT 67.800 110.800 78.600 111.100 ;
        RECT 83.000 111.100 83.400 111.200 ;
        RECT 84.600 111.100 85.000 111.200 ;
        RECT 99.000 111.100 99.400 111.200 ;
        RECT 83.000 110.800 99.400 111.100 ;
        RECT 109.400 111.100 109.800 111.200 ;
        RECT 117.400 111.100 117.800 111.200 ;
        RECT 109.400 110.800 117.800 111.100 ;
        RECT 124.600 111.100 125.000 111.200 ;
        RECT 128.600 111.100 129.000 111.200 ;
        RECT 124.600 110.800 129.000 111.100 ;
        RECT 152.600 111.100 153.000 111.200 ;
        RECT 162.200 111.100 162.600 111.200 ;
        RECT 152.600 110.800 162.600 111.100 ;
        RECT 172.600 111.100 173.000 111.200 ;
        RECT 199.000 111.100 199.400 111.200 ;
        RECT 172.600 110.800 199.400 111.100 ;
        RECT 203.800 111.100 204.200 111.200 ;
        RECT 205.400 111.100 205.800 111.200 ;
        RECT 203.800 110.800 205.800 111.100 ;
        RECT 210.200 111.100 210.600 111.200 ;
        RECT 231.000 111.100 231.400 111.200 ;
        RECT 210.200 110.800 231.400 111.100 ;
        RECT 45.400 109.800 45.800 110.200 ;
        RECT 53.400 110.100 53.800 110.200 ;
        RECT 57.400 110.100 57.800 110.200 ;
        RECT 92.600 110.100 93.000 110.200 ;
        RECT 53.400 109.800 93.000 110.100 ;
        RECT 138.200 110.100 138.600 110.200 ;
        RECT 173.400 110.100 173.800 110.200 ;
        RECT 174.200 110.100 174.600 110.200 ;
        RECT 138.200 109.800 174.600 110.100 ;
        RECT 212.600 109.800 213.000 110.200 ;
        RECT 14.200 109.100 14.600 109.200 ;
        RECT 19.000 109.100 19.400 109.200 ;
        RECT 30.200 109.100 30.600 109.200 ;
        RECT 14.200 108.800 30.600 109.100 ;
        RECT 34.200 109.100 34.600 109.200 ;
        RECT 45.400 109.100 45.700 109.800 ;
        RECT 212.600 109.200 212.900 109.800 ;
        RECT 34.200 108.800 45.700 109.100 ;
        RECT 63.800 109.100 64.200 109.200 ;
        RECT 67.800 109.100 68.200 109.200 ;
        RECT 63.800 108.800 68.200 109.100 ;
        RECT 95.000 109.100 95.400 109.200 ;
        RECT 106.200 109.100 106.600 109.200 ;
        RECT 95.000 108.800 106.600 109.100 ;
        RECT 111.000 109.100 111.400 109.200 ;
        RECT 111.800 109.100 112.200 109.200 ;
        RECT 111.000 108.800 112.200 109.100 ;
        RECT 177.400 109.100 177.800 109.200 ;
        RECT 177.400 108.800 183.300 109.100 ;
        RECT 212.600 108.800 213.000 109.200 ;
        RECT 232.600 108.800 233.000 109.200 ;
        RECT 247.000 109.100 247.400 109.200 ;
        RECT 253.400 109.100 253.800 109.200 ;
        RECT 246.200 108.800 253.800 109.100 ;
        RECT 183.000 108.200 183.300 108.800 ;
        RECT 15.000 108.100 15.400 108.200 ;
        RECT 17.400 108.100 17.800 108.200 ;
        RECT 25.400 108.100 25.800 108.200 ;
        RECT 103.800 108.100 104.200 108.200 ;
        RECT 15.000 107.800 104.200 108.100 ;
        RECT 110.200 108.100 110.600 108.200 ;
        RECT 113.400 108.100 113.800 108.200 ;
        RECT 144.600 108.100 145.000 108.200 ;
        RECT 110.200 107.800 145.000 108.100 ;
        RECT 148.600 108.100 149.000 108.200 ;
        RECT 160.600 108.100 161.000 108.200 ;
        RECT 148.600 107.800 161.000 108.100 ;
        RECT 163.000 107.800 163.400 108.200 ;
        RECT 164.600 108.100 165.000 108.200 ;
        RECT 167.800 108.100 168.200 108.200 ;
        RECT 164.600 107.800 168.200 108.100 ;
        RECT 179.000 107.800 179.400 108.200 ;
        RECT 183.000 107.800 183.400 108.200 ;
        RECT 187.000 108.100 187.400 108.200 ;
        RECT 188.600 108.100 189.000 108.200 ;
        RECT 204.600 108.100 205.000 108.200 ;
        RECT 206.200 108.100 206.600 108.200 ;
        RECT 187.000 107.800 206.600 108.100 ;
        RECT 209.400 108.100 209.800 108.200 ;
        RECT 223.000 108.100 223.400 108.200 ;
        RECT 209.400 107.800 223.400 108.100 ;
        RECT 226.200 108.100 226.600 108.200 ;
        RECT 227.800 108.100 228.200 108.200 ;
        RECT 226.200 107.800 228.200 108.100 ;
        RECT 230.200 108.100 230.600 108.200 ;
        RECT 232.600 108.100 232.900 108.800 ;
        RECT 230.200 107.800 232.900 108.100 ;
        RECT 163.000 107.200 163.300 107.800 ;
        RECT 3.000 107.100 3.400 107.200 ;
        RECT 41.400 107.100 41.800 107.200 ;
        RECT 3.000 106.800 20.900 107.100 ;
        RECT 20.600 106.200 20.900 106.800 ;
        RECT 33.400 106.800 41.800 107.100 ;
        RECT 71.800 107.100 72.200 107.200 ;
        RECT 77.400 107.100 77.800 107.200 ;
        RECT 71.800 106.800 77.800 107.100 ;
        RECT 83.800 107.100 84.200 107.200 ;
        RECT 89.400 107.100 89.800 107.200 ;
        RECT 83.800 106.800 89.800 107.100 ;
        RECT 115.800 107.100 116.200 107.200 ;
        RECT 132.600 107.100 133.000 107.200 ;
        RECT 115.800 106.800 133.000 107.100 ;
        RECT 134.200 106.800 134.600 107.200 ;
        RECT 136.600 107.100 137.000 107.200 ;
        RECT 141.400 107.100 141.800 107.200 ;
        RECT 144.600 107.100 145.000 107.200 ;
        RECT 136.600 106.800 145.000 107.100 ;
        RECT 155.000 107.100 155.400 107.200 ;
        RECT 160.600 107.100 161.000 107.200 ;
        RECT 155.000 106.800 161.000 107.100 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 163.800 107.100 164.200 107.200 ;
        RECT 165.400 107.100 165.800 107.200 ;
        RECT 163.800 106.800 165.800 107.100 ;
        RECT 179.000 107.100 179.300 107.800 ;
        RECT 199.800 107.100 200.200 107.200 ;
        RECT 219.000 107.100 219.400 107.200 ;
        RECT 239.800 107.100 240.200 107.200 ;
        RECT 251.000 107.100 251.400 107.200 ;
        RECT 179.000 106.800 251.400 107.100 ;
        RECT 33.400 106.200 33.700 106.800 ;
        RECT 8.600 106.100 9.000 106.200 ;
        RECT 16.600 106.100 17.000 106.200 ;
        RECT 8.600 105.800 17.000 106.100 ;
        RECT 20.600 105.800 21.000 106.200 ;
        RECT 33.400 105.800 33.800 106.200 ;
        RECT 37.400 105.800 37.800 106.200 ;
        RECT 67.000 106.100 67.400 106.200 ;
        RECT 65.400 105.800 67.400 106.100 ;
        RECT 71.000 106.100 71.400 106.200 ;
        RECT 72.600 106.100 73.000 106.200 ;
        RECT 85.400 106.100 85.800 106.200 ;
        RECT 71.000 105.800 85.800 106.100 ;
        RECT 87.000 106.100 87.400 106.200 ;
        RECT 88.600 106.100 89.000 106.200 ;
        RECT 87.000 105.800 89.000 106.100 ;
        RECT 89.400 106.100 89.700 106.800 ;
        RECT 134.200 106.200 134.500 106.800 ;
        RECT 99.800 106.100 100.200 106.200 ;
        RECT 89.400 105.800 100.200 106.100 ;
        RECT 111.800 106.100 112.200 106.200 ;
        RECT 124.600 106.100 125.000 106.200 ;
        RECT 111.800 105.800 125.000 106.100 ;
        RECT 131.800 105.800 132.200 106.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 138.200 106.100 138.600 106.200 ;
        RECT 153.400 106.100 153.800 106.200 ;
        RECT 159.800 106.100 160.200 106.200 ;
        RECT 138.200 105.800 153.800 106.100 ;
        RECT 155.800 105.800 160.200 106.100 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 164.600 106.100 165.000 106.200 ;
        RECT 163.000 105.800 165.000 106.100 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 167.000 106.100 167.400 106.200 ;
        RECT 166.200 105.800 167.400 106.100 ;
        RECT 182.200 106.100 182.600 106.200 ;
        RECT 183.800 106.100 184.200 106.200 ;
        RECT 182.200 105.800 184.200 106.100 ;
        RECT 188.600 106.100 189.000 106.200 ;
        RECT 196.600 106.100 197.000 106.200 ;
        RECT 188.600 105.800 197.000 106.100 ;
        RECT 209.400 106.100 209.800 106.200 ;
        RECT 212.600 106.100 213.000 106.200 ;
        RECT 209.400 105.800 213.000 106.100 ;
        RECT 223.000 106.100 223.400 106.200 ;
        RECT 226.200 106.100 226.600 106.200 ;
        RECT 230.200 106.100 230.600 106.200 ;
        RECT 223.000 105.800 230.600 106.100 ;
        RECT 238.200 106.100 238.600 106.300 ;
        RECT 244.600 106.100 245.000 106.200 ;
        RECT 262.200 106.100 262.600 106.200 ;
        RECT 238.200 105.800 244.100 106.100 ;
        RECT 244.600 105.800 262.600 106.100 ;
        RECT 37.400 105.100 37.700 105.800 ;
        RECT 65.400 105.200 65.700 105.800 ;
        RECT 51.000 105.100 51.400 105.200 ;
        RECT 37.400 104.800 51.400 105.100 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 74.200 105.100 74.600 105.200 ;
        RECT 83.800 105.100 84.200 105.200 ;
        RECT 74.200 104.800 84.200 105.100 ;
        RECT 86.200 105.100 86.600 105.200 ;
        RECT 88.600 105.100 89.000 105.200 ;
        RECT 86.200 104.800 89.000 105.100 ;
        RECT 89.400 105.100 89.800 105.200 ;
        RECT 93.400 105.100 93.800 105.200 ;
        RECT 89.400 104.800 93.800 105.100 ;
        RECT 102.200 105.100 102.600 105.200 ;
        RECT 126.200 105.100 126.600 105.200 ;
        RECT 102.200 104.800 126.600 105.100 ;
        RECT 131.800 105.100 132.100 105.800 ;
        RECT 155.800 105.200 156.100 105.800 ;
        RECT 243.800 105.200 244.100 105.800 ;
        RECT 135.000 105.100 135.400 105.200 ;
        RECT 131.800 104.800 135.400 105.100 ;
        RECT 143.000 105.100 143.400 105.200 ;
        RECT 144.600 105.100 145.000 105.200 ;
        RECT 143.000 104.800 145.000 105.100 ;
        RECT 155.800 104.800 156.200 105.200 ;
        RECT 167.000 105.100 167.400 105.200 ;
        RECT 168.600 105.100 169.000 105.200 ;
        RECT 167.000 104.800 169.000 105.100 ;
        RECT 169.400 105.100 169.800 105.200 ;
        RECT 183.000 105.100 183.400 105.200 ;
        RECT 169.400 104.800 183.400 105.100 ;
        RECT 206.200 105.100 206.600 105.200 ;
        RECT 212.600 105.100 213.000 105.200 ;
        RECT 225.400 105.100 225.800 105.200 ;
        RECT 206.200 104.800 225.800 105.100 ;
        RECT 230.200 105.100 230.600 105.200 ;
        RECT 243.000 105.100 243.400 105.200 ;
        RECT 230.200 104.800 243.400 105.100 ;
        RECT 243.800 104.800 244.200 105.200 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 43.000 104.100 43.400 104.200 ;
        RECT 41.400 103.800 43.400 104.100 ;
        RECT 59.000 104.100 59.400 104.200 ;
        RECT 102.200 104.100 102.500 104.800 ;
        RECT 59.000 103.800 102.500 104.100 ;
        RECT 103.800 104.100 104.200 104.200 ;
        RECT 109.400 104.100 109.800 104.200 ;
        RECT 127.000 104.100 127.400 104.200 ;
        RECT 103.800 103.800 127.400 104.100 ;
        RECT 131.800 104.100 132.200 104.200 ;
        RECT 137.400 104.100 137.800 104.200 ;
        RECT 131.800 103.800 137.800 104.100 ;
        RECT 159.000 104.100 159.400 104.200 ;
        RECT 164.600 104.100 165.000 104.200 ;
        RECT 159.000 103.800 165.000 104.100 ;
        RECT 171.800 104.100 172.200 104.200 ;
        RECT 180.600 104.100 181.000 104.200 ;
        RECT 171.800 103.800 181.000 104.100 ;
        RECT 182.200 104.100 182.600 104.200 ;
        RECT 187.000 104.100 187.400 104.200 ;
        RECT 189.400 104.100 189.800 104.200 ;
        RECT 182.200 103.800 189.800 104.100 ;
        RECT 212.600 104.100 213.000 104.200 ;
        RECT 229.400 104.100 229.800 104.200 ;
        RECT 212.600 103.800 229.800 104.100 ;
        RECT 2.200 103.100 2.600 103.200 ;
        RECT 59.000 103.100 59.300 103.800 ;
        RECT 2.200 102.800 59.300 103.100 ;
        RECT 91.000 103.100 91.400 103.200 ;
        RECT 94.200 103.100 94.600 103.200 ;
        RECT 145.400 103.100 145.800 103.200 ;
        RECT 91.000 102.800 145.800 103.100 ;
        RECT 184.600 103.100 185.000 103.200 ;
        RECT 186.200 103.100 186.600 103.200 ;
        RECT 184.600 102.800 186.600 103.100 ;
        RECT 199.800 103.100 200.200 103.200 ;
        RECT 207.000 103.100 207.400 103.200 ;
        RECT 199.800 102.800 207.400 103.100 ;
        RECT 211.000 103.100 211.400 103.200 ;
        RECT 230.200 103.100 230.600 103.200 ;
        RECT 211.000 102.800 230.600 103.100 ;
        RECT 75.800 102.100 76.200 102.200 ;
        RECT 92.600 102.100 93.000 102.200 ;
        RECT 75.800 101.800 93.000 102.100 ;
        RECT 103.800 102.100 104.200 102.200 ;
        RECT 125.400 102.100 125.800 102.200 ;
        RECT 149.400 102.100 149.800 102.200 ;
        RECT 103.800 101.800 149.800 102.100 ;
        RECT 157.400 102.100 157.800 102.200 ;
        RECT 178.200 102.100 178.600 102.200 ;
        RECT 157.400 101.800 178.600 102.100 ;
        RECT 194.200 102.100 194.600 102.200 ;
        RECT 200.600 102.100 201.000 102.200 ;
        RECT 194.200 101.800 201.000 102.100 ;
        RECT 206.200 102.100 206.600 102.200 ;
        RECT 207.800 102.100 208.200 102.200 ;
        RECT 206.200 101.800 208.200 102.100 ;
        RECT 211.000 102.100 211.400 102.200 ;
        RECT 213.400 102.100 213.800 102.200 ;
        RECT 211.000 101.800 213.800 102.100 ;
        RECT 231.000 102.100 231.400 102.200 ;
        RECT 237.400 102.100 237.800 102.200 ;
        RECT 231.000 101.800 237.800 102.100 ;
        RECT 124.600 101.100 125.000 101.200 ;
        RECT 130.200 101.100 130.600 101.200 ;
        RECT 124.600 100.800 130.600 101.100 ;
        RECT 131.000 101.100 131.400 101.200 ;
        RECT 154.200 101.100 154.600 101.200 ;
        RECT 131.000 100.800 154.600 101.100 ;
        RECT 170.200 101.100 170.600 101.200 ;
        RECT 199.800 101.100 200.200 101.200 ;
        RECT 211.800 101.100 212.200 101.200 ;
        RECT 170.200 100.800 212.200 101.100 ;
        RECT 227.800 101.100 228.200 101.200 ;
        RECT 239.800 101.100 240.200 101.200 ;
        RECT 227.800 100.800 240.200 101.100 ;
        RECT 11.800 100.100 12.200 100.200 ;
        RECT 14.200 100.100 14.600 100.200 ;
        RECT 47.000 100.100 47.400 100.200 ;
        RECT 11.800 99.800 47.400 100.100 ;
        RECT 79.800 100.100 80.200 100.200 ;
        RECT 80.600 100.100 81.000 100.200 ;
        RECT 79.800 99.800 81.000 100.100 ;
        RECT 99.000 100.100 99.400 100.200 ;
        RECT 117.400 100.100 117.800 100.200 ;
        RECT 127.800 100.100 128.200 100.200 ;
        RECT 99.000 99.800 128.200 100.100 ;
        RECT 145.400 100.100 145.800 100.200 ;
        RECT 151.000 100.100 151.400 100.200 ;
        RECT 145.400 99.800 151.400 100.100 ;
        RECT 231.800 100.100 232.200 100.200 ;
        RECT 238.200 100.100 238.600 100.200 ;
        RECT 231.800 99.800 238.600 100.100 ;
        RECT 19.000 99.100 19.400 99.200 ;
        RECT 29.400 99.100 29.800 99.200 ;
        RECT 41.400 99.100 41.800 99.200 ;
        RECT 56.600 99.100 57.000 99.200 ;
        RECT 67.800 99.100 68.200 99.200 ;
        RECT 87.000 99.100 87.400 99.200 ;
        RECT 129.400 99.100 129.800 99.200 ;
        RECT 161.400 99.100 161.800 99.200 ;
        RECT 19.000 98.800 197.700 99.100 ;
        RECT 197.400 98.200 197.700 98.800 ;
        RECT 34.200 98.100 34.600 98.200 ;
        RECT 36.600 98.100 37.000 98.200 ;
        RECT 58.200 98.100 58.600 98.200 ;
        RECT 71.000 98.100 71.400 98.200 ;
        RECT 34.200 97.800 71.400 98.100 ;
        RECT 90.200 98.100 90.600 98.200 ;
        RECT 95.000 98.100 95.400 98.200 ;
        RECT 90.200 97.800 95.400 98.100 ;
        RECT 128.600 98.100 129.000 98.200 ;
        RECT 132.600 98.100 133.000 98.200 ;
        RECT 128.600 97.800 133.000 98.100 ;
        RECT 137.400 98.100 137.800 98.200 ;
        RECT 141.400 98.100 141.800 98.200 ;
        RECT 137.400 97.800 141.800 98.100 ;
        RECT 197.400 97.800 197.800 98.200 ;
        RECT 201.400 98.100 201.800 98.200 ;
        RECT 227.000 98.100 227.400 98.200 ;
        RECT 201.400 97.800 227.400 98.100 ;
        RECT 10.200 97.100 10.600 97.200 ;
        RECT 16.600 97.100 17.000 97.200 ;
        RECT 10.200 96.800 17.000 97.100 ;
        RECT 70.200 97.100 70.600 97.200 ;
        RECT 82.200 97.100 82.600 97.200 ;
        RECT 70.200 96.800 82.600 97.100 ;
        RECT 115.000 97.100 115.400 97.200 ;
        RECT 123.800 97.100 124.200 97.200 ;
        RECT 115.000 96.800 124.200 97.100 ;
        RECT 126.200 97.100 126.600 97.200 ;
        RECT 134.200 97.100 134.600 97.200 ;
        RECT 150.200 97.100 150.600 97.200 ;
        RECT 126.200 96.800 150.600 97.100 ;
        RECT 151.000 96.800 151.400 97.200 ;
        RECT 175.800 97.100 176.200 97.200 ;
        RECT 185.400 97.100 185.800 97.200 ;
        RECT 195.800 97.100 196.200 97.200 ;
        RECT 219.800 97.100 220.200 97.200 ;
        RECT 227.800 97.100 228.200 97.200 ;
        RECT 255.000 97.100 255.400 97.200 ;
        RECT 175.800 96.800 196.200 97.100 ;
        RECT 219.000 96.800 255.400 97.100 ;
        RECT 15.800 95.800 16.200 96.200 ;
        RECT 26.200 96.100 26.600 96.200 ;
        RECT 35.000 96.100 35.400 96.200 ;
        RECT 26.200 95.800 35.400 96.100 ;
        RECT 40.600 96.100 41.000 96.200 ;
        RECT 42.200 96.100 42.600 96.200 ;
        RECT 40.600 95.800 42.600 96.100 ;
        RECT 46.200 96.100 46.600 96.200 ;
        RECT 47.800 96.100 48.200 96.200 ;
        RECT 64.600 96.100 65.000 96.200 ;
        RECT 71.000 96.100 71.400 96.200 ;
        RECT 46.200 95.800 48.200 96.100 ;
        RECT 63.800 95.800 71.400 96.100 ;
        RECT 91.800 95.800 92.200 96.200 ;
        RECT 128.600 95.800 129.000 96.200 ;
        RECT 139.000 96.100 139.400 96.200 ;
        RECT 141.400 96.100 141.800 96.200 ;
        RECT 139.000 95.800 141.800 96.100 ;
        RECT 142.200 96.100 142.600 96.200 ;
        RECT 151.000 96.100 151.300 96.800 ;
        RECT 142.200 95.800 151.300 96.100 ;
        RECT 154.200 96.100 154.600 96.200 ;
        RECT 159.800 96.100 160.200 96.200 ;
        RECT 154.200 95.800 160.200 96.100 ;
        RECT 172.600 96.100 173.000 96.200 ;
        RECT 175.000 96.100 175.400 96.200 ;
        RECT 172.600 95.800 175.400 96.100 ;
        RECT 180.600 95.800 181.000 96.200 ;
        RECT 193.400 96.100 193.800 96.200 ;
        RECT 248.600 96.100 249.000 96.200 ;
        RECT 250.200 96.100 250.600 96.200 ;
        RECT 193.400 95.800 250.600 96.100 ;
        RECT 15.800 95.200 16.100 95.800 ;
        RECT 91.800 95.200 92.100 95.800 ;
        RECT 128.600 95.200 128.900 95.800 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 15.800 95.100 16.200 95.200 ;
        RECT 6.200 94.800 16.200 95.100 ;
        RECT 22.200 95.100 22.600 95.200 ;
        RECT 27.800 95.100 28.200 95.200 ;
        RECT 32.600 95.100 33.000 95.200 ;
        RECT 70.200 95.100 70.600 95.200 ;
        RECT 22.200 94.800 70.600 95.100 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 95.800 95.100 96.200 95.200 ;
        RECT 113.400 95.100 113.800 95.200 ;
        RECT 128.600 95.100 129.000 95.200 ;
        RECT 131.000 95.100 131.400 95.200 ;
        RECT 95.800 94.800 104.100 95.100 ;
        RECT 113.400 94.800 118.500 95.100 ;
        RECT 128.600 94.800 131.400 95.100 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 143.800 95.100 144.200 95.200 ;
        RECT 139.000 94.800 144.200 95.100 ;
        RECT 150.200 95.100 150.600 95.200 ;
        RECT 152.600 95.100 153.000 95.200 ;
        RECT 150.200 94.800 153.000 95.100 ;
        RECT 156.600 95.100 157.000 95.200 ;
        RECT 157.400 95.100 157.800 95.200 ;
        RECT 156.600 94.800 157.800 95.100 ;
        RECT 165.400 95.100 165.800 95.200 ;
        RECT 172.600 95.100 173.000 95.200 ;
        RECT 165.400 94.800 173.000 95.100 ;
        RECT 176.600 94.800 177.000 95.200 ;
        RECT 180.600 95.100 180.900 95.800 ;
        RECT 181.400 95.100 181.800 95.200 ;
        RECT 186.200 95.100 186.600 95.200 ;
        RECT 180.600 94.800 181.800 95.100 ;
        RECT 184.600 94.800 186.600 95.100 ;
        RECT 187.800 95.100 188.200 95.200 ;
        RECT 191.800 95.100 192.200 95.200 ;
        RECT 187.800 94.800 192.200 95.100 ;
        RECT 196.600 95.100 197.000 95.200 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 201.400 95.100 201.800 95.200 ;
        RECT 227.000 95.100 227.400 95.200 ;
        RECT 231.000 95.100 231.400 95.200 ;
        RECT 196.600 94.800 202.500 95.100 ;
        RECT 227.000 94.800 231.400 95.100 ;
        RECT 239.000 95.100 239.400 95.200 ;
        RECT 251.000 95.100 251.400 95.200 ;
        RECT 239.000 94.800 251.400 95.100 ;
        RECT 5.400 94.100 5.800 94.200 ;
        RECT 11.800 94.100 12.200 94.200 ;
        RECT 5.400 93.800 12.200 94.100 ;
        RECT 15.800 94.100 16.200 94.200 ;
        RECT 28.600 94.100 29.000 94.200 ;
        RECT 39.000 94.100 39.400 94.200 ;
        RECT 15.800 93.800 39.400 94.100 ;
        RECT 47.800 94.100 48.200 94.200 ;
        RECT 58.200 94.100 58.600 94.200 ;
        RECT 47.800 93.800 58.600 94.100 ;
        RECT 70.200 94.100 70.600 94.200 ;
        RECT 71.000 94.100 71.400 94.200 ;
        RECT 70.200 93.800 71.400 94.100 ;
        RECT 73.400 94.100 73.700 94.800 ;
        RECT 75.000 94.100 75.300 94.800 ;
        RECT 103.800 94.200 104.100 94.800 ;
        RECT 118.200 94.200 118.500 94.800 ;
        RECT 73.400 93.800 75.300 94.100 ;
        RECT 82.200 94.100 82.600 94.200 ;
        RECT 90.200 94.100 90.600 94.200 ;
        RECT 82.200 93.800 90.600 94.100 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 139.800 94.100 140.200 94.200 ;
        RECT 142.200 94.100 142.600 94.200 ;
        RECT 139.800 93.800 142.600 94.100 ;
        RECT 151.000 94.100 151.400 94.200 ;
        RECT 155.800 94.100 156.200 94.200 ;
        RECT 151.000 93.800 156.200 94.100 ;
        RECT 162.200 94.100 162.600 94.200 ;
        RECT 164.600 94.100 165.000 94.200 ;
        RECT 176.600 94.100 176.900 94.800 ;
        RECT 162.200 93.800 176.900 94.100 ;
        RECT 184.600 94.200 184.900 94.800 ;
        RECT 184.600 93.800 185.000 94.200 ;
        RECT 189.400 94.100 189.800 94.200 ;
        RECT 191.000 94.100 191.400 94.200 ;
        RECT 189.400 93.800 191.400 94.100 ;
        RECT 23.800 93.100 24.200 93.200 ;
        RECT 24.600 93.100 25.000 93.200 ;
        RECT 23.800 92.800 25.000 93.100 ;
        RECT 39.000 93.100 39.400 93.200 ;
        RECT 59.000 93.100 59.400 93.200 ;
        RECT 63.800 93.100 64.200 93.200 ;
        RECT 39.000 92.800 64.200 93.100 ;
        RECT 64.600 93.100 65.000 93.200 ;
        RECT 75.000 93.100 75.400 93.200 ;
        RECT 64.600 92.800 75.400 93.100 ;
        RECT 87.800 93.100 88.200 93.200 ;
        RECT 97.400 93.100 97.800 93.200 ;
        RECT 87.800 92.800 97.800 93.100 ;
        RECT 106.200 93.100 106.600 93.200 ;
        RECT 119.800 93.100 120.200 93.200 ;
        RECT 106.200 92.800 120.200 93.100 ;
        RECT 138.200 93.100 138.600 93.200 ;
        RECT 148.600 93.100 149.000 93.200 ;
        RECT 151.800 93.100 152.200 93.200 ;
        RECT 138.200 92.800 152.200 93.100 ;
        RECT 200.600 92.800 201.000 93.200 ;
        RECT 220.600 93.100 221.000 93.200 ;
        RECT 233.400 93.100 233.800 93.200 ;
        RECT 245.400 93.100 245.800 93.200 ;
        RECT 220.600 92.800 245.800 93.100 ;
        RECT 246.200 93.100 246.600 93.200 ;
        RECT 255.000 93.100 255.400 93.200 ;
        RECT 258.200 93.100 258.600 93.200 ;
        RECT 246.200 92.800 253.700 93.100 ;
        RECT 255.000 92.800 258.600 93.100 ;
        RECT 10.200 92.100 10.600 92.200 ;
        RECT 43.800 92.100 44.200 92.200 ;
        RECT 10.200 91.800 44.200 92.100 ;
        RECT 78.200 92.100 78.600 92.200 ;
        RECT 89.400 92.100 89.800 92.200 ;
        RECT 103.800 92.100 104.200 92.200 ;
        RECT 78.200 91.800 104.200 92.100 ;
        RECT 119.000 92.100 119.400 92.200 ;
        RECT 130.200 92.100 130.600 92.200 ;
        RECT 119.000 91.800 130.600 92.100 ;
        RECT 147.800 92.100 148.200 92.200 ;
        RECT 163.800 92.100 164.200 92.200 ;
        RECT 147.800 91.800 164.200 92.100 ;
        RECT 176.600 92.100 177.000 92.200 ;
        RECT 184.600 92.100 185.000 92.200 ;
        RECT 176.600 91.800 185.000 92.100 ;
        RECT 187.000 92.100 187.400 92.200 ;
        RECT 187.800 92.100 188.200 92.200 ;
        RECT 190.200 92.100 190.600 92.200 ;
        RECT 200.600 92.100 200.900 92.800 ;
        RECT 253.400 92.200 253.700 92.800 ;
        RECT 187.000 91.800 200.900 92.100 ;
        RECT 208.600 92.100 209.000 92.200 ;
        RECT 211.800 92.100 212.200 92.200 ;
        RECT 208.600 91.800 212.200 92.100 ;
        RECT 221.400 92.100 221.800 92.200 ;
        RECT 234.200 92.100 234.600 92.200 ;
        RECT 221.400 91.800 234.600 92.100 ;
        RECT 253.400 91.800 253.800 92.200 ;
        RECT 41.400 91.100 41.800 91.200 ;
        RECT 45.400 91.100 45.800 91.200 ;
        RECT 64.600 91.100 65.000 91.200 ;
        RECT 41.400 90.800 65.000 91.100 ;
        RECT 75.000 91.100 75.400 91.200 ;
        RECT 92.600 91.100 93.000 91.200 ;
        RECT 98.200 91.100 98.600 91.200 ;
        RECT 103.000 91.100 103.400 91.200 ;
        RECT 75.000 90.800 103.400 91.100 ;
        RECT 119.800 91.100 120.200 91.200 ;
        RECT 143.000 91.100 143.400 91.200 ;
        RECT 119.800 90.800 143.400 91.100 ;
        RECT 167.800 91.100 168.200 91.200 ;
        RECT 182.200 91.100 182.600 91.200 ;
        RECT 167.800 90.800 182.600 91.100 ;
        RECT 183.800 91.100 184.200 91.200 ;
        RECT 194.200 91.100 194.600 91.200 ;
        RECT 183.800 90.800 194.600 91.100 ;
        RECT 215.800 91.100 216.200 91.200 ;
        RECT 241.400 91.100 241.800 91.200 ;
        RECT 251.800 91.100 252.200 91.200 ;
        RECT 215.800 90.800 252.200 91.100 ;
        RECT 59.800 90.100 60.200 90.200 ;
        RECT 62.200 90.100 62.600 90.200 ;
        RECT 59.800 89.800 62.600 90.100 ;
        RECT 79.000 90.100 79.400 90.200 ;
        RECT 83.800 90.100 84.200 90.200 ;
        RECT 79.000 89.800 84.200 90.100 ;
        RECT 115.000 90.100 115.400 90.200 ;
        RECT 121.400 90.100 121.800 90.200 ;
        RECT 138.200 90.100 138.600 90.200 ;
        RECT 115.000 89.800 138.600 90.100 ;
        RECT 159.800 90.100 160.200 90.200 ;
        RECT 163.800 90.100 164.200 90.200 ;
        RECT 159.800 89.800 164.200 90.100 ;
        RECT 188.600 90.100 189.000 90.200 ;
        RECT 191.800 90.100 192.200 90.200 ;
        RECT 188.600 89.800 192.200 90.100 ;
        RECT 195.800 90.100 196.200 90.200 ;
        RECT 204.600 90.100 205.000 90.200 ;
        RECT 195.800 89.800 205.000 90.100 ;
        RECT 219.800 90.100 220.200 90.200 ;
        RECT 223.000 90.100 223.400 90.200 ;
        RECT 219.800 89.800 223.400 90.100 ;
        RECT 237.400 90.100 237.800 90.200 ;
        RECT 239.800 90.100 240.200 90.200 ;
        RECT 262.200 90.100 262.600 90.200 ;
        RECT 237.400 89.800 262.600 90.100 ;
        RECT 17.400 89.100 17.800 89.200 ;
        RECT 19.800 89.100 20.200 89.200 ;
        RECT 17.400 88.800 20.200 89.100 ;
        RECT 48.600 89.100 49.000 89.200 ;
        RECT 76.600 89.100 77.000 89.200 ;
        RECT 48.600 88.800 77.000 89.100 ;
        RECT 80.600 88.800 81.000 89.200 ;
        RECT 83.000 89.100 83.400 89.200 ;
        RECT 91.800 89.100 92.200 89.200 ;
        RECT 92.600 89.100 93.000 89.200 ;
        RECT 83.000 88.800 93.000 89.100 ;
        RECT 123.800 89.100 124.200 89.200 ;
        RECT 135.800 89.100 136.200 89.200 ;
        RECT 123.800 88.800 136.200 89.100 ;
        RECT 159.000 89.100 159.400 89.200 ;
        RECT 173.400 89.100 173.800 89.200 ;
        RECT 174.200 89.100 174.600 89.200 ;
        RECT 159.000 88.800 174.600 89.100 ;
        RECT 177.400 89.100 177.800 89.200 ;
        RECT 178.200 89.100 178.600 89.200 ;
        RECT 177.400 88.800 178.600 89.100 ;
        RECT 194.200 89.100 194.600 89.200 ;
        RECT 197.400 89.100 197.800 89.200 ;
        RECT 194.200 88.800 197.800 89.100 ;
        RECT 199.000 89.100 199.400 89.200 ;
        RECT 231.800 89.100 232.200 89.200 ;
        RECT 199.000 88.800 232.200 89.100 ;
        RECT 80.600 88.200 80.900 88.800 ;
        RECT 52.600 88.100 53.000 88.200 ;
        RECT 60.600 88.100 61.000 88.200 ;
        RECT 71.800 88.100 72.200 88.200 ;
        RECT 52.600 87.800 72.200 88.100 ;
        RECT 80.600 87.800 81.000 88.200 ;
        RECT 99.800 88.100 100.200 88.200 ;
        RECT 105.400 88.100 105.800 88.200 ;
        RECT 99.800 87.800 105.800 88.100 ;
        RECT 135.000 88.100 135.400 88.200 ;
        RECT 144.600 88.100 145.000 88.200 ;
        RECT 135.000 87.800 145.000 88.100 ;
        RECT 146.200 88.100 146.600 88.200 ;
        RECT 149.400 88.100 149.800 88.200 ;
        RECT 182.200 88.100 182.600 88.200 ;
        RECT 214.200 88.100 214.600 88.200 ;
        RECT 223.800 88.100 224.200 88.200 ;
        RECT 227.800 88.100 228.200 88.200 ;
        RECT 146.200 87.800 228.200 88.100 ;
        RECT 255.800 88.100 256.200 88.200 ;
        RECT 257.400 88.100 257.800 88.200 ;
        RECT 255.800 87.800 257.800 88.100 ;
        RECT 22.200 87.100 22.600 87.200 ;
        RECT 27.000 87.100 27.400 87.200 ;
        RECT 22.200 86.800 27.400 87.100 ;
        RECT 45.400 86.800 45.800 87.200 ;
        RECT 55.000 86.800 55.400 87.200 ;
        RECT 65.400 87.100 65.800 87.200 ;
        RECT 75.000 87.100 75.400 87.200 ;
        RECT 83.800 87.100 84.200 87.200 ;
        RECT 65.400 86.800 84.200 87.100 ;
        RECT 103.000 86.800 103.400 87.200 ;
        RECT 112.600 87.100 113.000 87.200 ;
        RECT 121.400 87.100 121.800 87.200 ;
        RECT 112.600 86.800 121.800 87.100 ;
        RECT 124.600 86.800 125.000 87.200 ;
        RECT 128.600 87.100 129.000 87.200 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 128.600 86.800 137.800 87.100 ;
        RECT 140.600 87.100 141.000 87.200 ;
        RECT 147.000 87.100 147.400 87.200 ;
        RECT 147.800 87.100 148.200 87.200 ;
        RECT 140.600 86.800 148.200 87.100 ;
        RECT 157.400 87.100 157.800 87.200 ;
        RECT 161.400 87.100 161.800 87.200 ;
        RECT 157.400 86.800 161.800 87.100 ;
        RECT 169.400 86.800 169.800 87.200 ;
        RECT 175.000 87.100 175.400 87.200 ;
        RECT 188.600 87.100 189.000 87.200 ;
        RECT 189.400 87.100 189.800 87.200 ;
        RECT 175.000 86.800 183.300 87.100 ;
        RECT 188.600 86.800 189.800 87.100 ;
        RECT 190.200 87.100 190.600 87.200 ;
        RECT 195.000 87.100 195.400 87.200 ;
        RECT 200.600 87.100 201.000 87.200 ;
        RECT 204.600 87.100 205.000 87.200 ;
        RECT 212.600 87.100 213.000 87.200 ;
        RECT 190.200 86.800 195.400 87.100 ;
        RECT 197.400 86.800 199.300 87.100 ;
        RECT 200.600 86.800 213.000 87.100 ;
        RECT 219.000 86.800 219.400 87.200 ;
        RECT 223.000 87.100 223.400 87.200 ;
        RECT 255.800 87.100 256.200 87.200 ;
        RECT 223.000 86.800 256.200 87.100 ;
        RECT 257.400 86.800 257.800 87.200 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 4.600 85.800 12.200 86.100 ;
        RECT 16.600 86.100 17.000 86.200 ;
        RECT 17.400 86.100 17.800 86.200 ;
        RECT 16.600 85.800 17.800 86.100 ;
        RECT 26.200 85.800 26.600 86.200 ;
        RECT 34.200 86.100 34.600 86.200 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 34.200 85.800 40.200 86.100 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 45.400 86.100 45.700 86.800 ;
        RECT 51.800 86.100 52.200 86.200 ;
        RECT 45.400 85.800 52.200 86.100 ;
        RECT 55.000 86.100 55.300 86.800 ;
        RECT 103.000 86.200 103.300 86.800 ;
        RECT 57.400 86.100 57.800 86.200 ;
        RECT 65.400 86.100 65.800 86.200 ;
        RECT 72.600 86.100 73.000 86.200 ;
        RECT 55.000 85.800 65.800 86.100 ;
        RECT 67.000 85.800 73.000 86.100 ;
        RECT 75.800 86.100 76.200 86.200 ;
        RECT 76.600 86.100 77.000 86.200 ;
        RECT 75.800 85.800 77.000 86.100 ;
        RECT 103.000 85.800 103.400 86.200 ;
        RECT 119.800 86.100 120.200 86.200 ;
        RECT 121.400 86.100 121.800 86.200 ;
        RECT 119.800 85.800 121.800 86.100 ;
        RECT 123.800 86.100 124.200 86.200 ;
        RECT 124.600 86.100 124.900 86.800 ;
        RECT 123.800 85.800 124.900 86.100 ;
        RECT 135.800 86.100 136.200 86.200 ;
        RECT 138.200 86.100 138.600 86.200 ;
        RECT 139.000 86.100 139.400 86.200 ;
        RECT 135.800 85.800 139.400 86.100 ;
        RECT 143.800 86.100 144.200 86.200 ;
        RECT 169.400 86.100 169.700 86.800 ;
        RECT 183.000 86.200 183.300 86.800 ;
        RECT 197.400 86.200 197.700 86.800 ;
        RECT 199.000 86.200 199.300 86.800 ;
        RECT 219.000 86.200 219.300 86.800 ;
        RECT 172.600 86.100 173.000 86.200 ;
        RECT 143.800 85.800 173.000 86.100 ;
        RECT 183.000 85.800 183.400 86.200 ;
        RECT 187.800 86.100 188.200 86.200 ;
        RECT 192.600 86.100 193.000 86.200 ;
        RECT 187.800 85.800 193.000 86.100 ;
        RECT 197.400 85.800 197.800 86.200 ;
        RECT 199.000 85.800 199.400 86.200 ;
        RECT 206.200 86.100 206.600 86.200 ;
        RECT 213.400 86.100 213.800 86.200 ;
        RECT 206.200 85.800 213.800 86.100 ;
        RECT 215.800 86.100 216.200 86.200 ;
        RECT 216.600 86.100 217.000 86.200 ;
        RECT 215.800 85.800 217.000 86.100 ;
        RECT 219.000 85.800 219.400 86.200 ;
        RECT 257.400 86.100 257.700 86.800 ;
        RECT 260.600 86.100 261.000 86.200 ;
        RECT 257.400 85.800 261.000 86.100 ;
        RECT 21.400 85.100 21.800 85.200 ;
        RECT 26.200 85.100 26.500 85.800 ;
        RECT 21.400 84.800 26.500 85.100 ;
        RECT 43.800 85.100 44.100 85.800 ;
        RECT 67.000 85.200 67.300 85.800 ;
        RECT 47.800 85.100 48.200 85.200 ;
        RECT 43.800 84.800 48.200 85.100 ;
        RECT 67.000 84.800 67.400 85.200 ;
        RECT 70.200 85.100 70.600 85.200 ;
        RECT 74.200 85.100 74.600 85.200 ;
        RECT 70.200 84.800 74.600 85.100 ;
        RECT 92.600 85.100 93.000 85.200 ;
        RECT 106.200 85.100 106.600 85.200 ;
        RECT 92.600 84.800 106.600 85.100 ;
        RECT 111.800 85.100 112.200 85.200 ;
        RECT 129.400 85.100 129.800 85.200 ;
        RECT 160.600 85.100 161.000 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 111.800 84.800 162.600 85.100 ;
        RECT 181.400 84.800 181.800 85.200 ;
        RECT 182.200 85.100 182.600 85.200 ;
        RECT 206.200 85.100 206.500 85.800 ;
        RECT 182.200 84.800 206.500 85.100 ;
        RECT 213.400 85.100 213.700 85.800 ;
        RECT 223.000 85.100 223.400 85.200 ;
        RECT 228.600 85.100 229.000 85.200 ;
        RECT 213.400 84.800 229.000 85.100 ;
        RECT 241.400 85.100 241.800 85.200 ;
        RECT 247.000 85.100 247.400 85.200 ;
        RECT 253.400 85.100 253.800 85.200 ;
        RECT 258.200 85.100 258.600 85.200 ;
        RECT 241.400 84.800 258.600 85.100 ;
        RECT 25.400 83.800 25.800 84.200 ;
        RECT 39.000 84.100 39.400 84.200 ;
        RECT 42.200 84.100 42.600 84.200 ;
        RECT 39.000 83.800 42.600 84.100 ;
        RECT 88.600 84.100 89.000 84.200 ;
        RECT 91.800 84.100 92.200 84.200 ;
        RECT 88.600 83.800 92.200 84.100 ;
        RECT 139.000 84.100 139.400 84.200 ;
        RECT 142.200 84.100 142.600 84.200 ;
        RECT 139.000 83.800 142.600 84.100 ;
        RECT 144.600 84.100 145.000 84.200 ;
        RECT 163.000 84.100 163.400 84.200 ;
        RECT 144.600 83.800 163.400 84.100 ;
        RECT 181.400 84.100 181.700 84.800 ;
        RECT 183.000 84.100 183.400 84.200 ;
        RECT 181.400 83.800 183.400 84.100 ;
        RECT 192.600 84.100 193.000 84.200 ;
        RECT 211.800 84.100 212.200 84.200 ;
        RECT 215.000 84.100 215.400 84.200 ;
        RECT 192.600 83.800 212.200 84.100 ;
        RECT 213.400 83.800 215.400 84.100 ;
        RECT 25.400 83.200 25.700 83.800 ;
        RECT 213.400 83.200 213.700 83.800 ;
        RECT 25.400 82.800 25.800 83.200 ;
        RECT 76.600 83.100 77.000 83.200 ;
        RECT 79.000 83.100 79.400 83.200 ;
        RECT 76.600 82.800 79.400 83.100 ;
        RECT 159.000 83.100 159.400 83.200 ;
        RECT 185.400 83.100 185.800 83.200 ;
        RECT 159.000 82.800 185.800 83.100 ;
        RECT 213.400 82.800 213.800 83.200 ;
        RECT 230.200 83.100 230.600 83.200 ;
        RECT 234.200 83.100 234.600 83.200 ;
        RECT 230.200 82.800 234.600 83.100 ;
        RECT 141.400 82.100 141.800 82.200 ;
        RECT 163.800 82.100 164.200 82.200 ;
        RECT 141.400 81.800 164.200 82.100 ;
        RECT 165.400 82.100 165.800 82.200 ;
        RECT 197.400 82.100 197.800 82.200 ;
        RECT 165.400 81.800 197.800 82.100 ;
        RECT 198.200 82.100 198.600 82.200 ;
        RECT 221.400 82.100 221.800 82.200 ;
        RECT 198.200 81.800 221.800 82.100 ;
        RECT 222.200 82.100 222.600 82.200 ;
        RECT 231.000 82.100 231.400 82.200 ;
        RECT 222.200 81.800 231.400 82.100 ;
        RECT 24.600 81.100 25.000 81.200 ;
        RECT 25.400 81.100 25.800 81.200 ;
        RECT 24.600 80.800 25.800 81.100 ;
        RECT 90.200 81.100 90.600 81.200 ;
        RECT 108.600 81.100 109.000 81.200 ;
        RECT 90.200 80.800 109.000 81.100 ;
        RECT 110.200 81.100 110.600 81.200 ;
        RECT 141.400 81.100 141.800 81.200 ;
        RECT 110.200 80.800 141.800 81.100 ;
        RECT 163.000 81.100 163.400 81.200 ;
        RECT 182.200 81.100 182.600 81.200 ;
        RECT 163.000 80.800 182.600 81.100 ;
        RECT 185.400 81.100 185.800 81.200 ;
        RECT 217.400 81.100 217.800 81.200 ;
        RECT 223.800 81.100 224.200 81.200 ;
        RECT 185.400 80.800 224.200 81.100 ;
        RECT 225.400 81.100 225.800 81.200 ;
        RECT 231.800 81.100 232.200 81.200 ;
        RECT 235.000 81.100 235.400 81.200 ;
        RECT 225.400 80.800 235.400 81.100 ;
        RECT 57.400 80.100 57.800 80.200 ;
        RECT 63.800 80.100 64.200 80.200 ;
        RECT 57.400 79.800 64.200 80.100 ;
        RECT 76.600 80.100 77.000 80.200 ;
        RECT 127.000 80.100 127.400 80.200 ;
        RECT 76.600 79.800 127.400 80.100 ;
        RECT 164.600 80.100 165.000 80.200 ;
        RECT 171.000 80.100 171.400 80.200 ;
        RECT 164.600 79.800 171.400 80.100 ;
        RECT 183.800 80.100 184.200 80.200 ;
        RECT 226.200 80.100 226.600 80.200 ;
        RECT 183.800 79.800 226.600 80.100 ;
        RECT 242.200 80.100 242.600 80.200 ;
        RECT 243.000 80.100 243.400 80.200 ;
        RECT 242.200 79.800 243.400 80.100 ;
        RECT 23.800 79.100 24.200 79.200 ;
        RECT 110.200 79.100 110.600 79.200 ;
        RECT 132.600 79.100 133.000 79.200 ;
        RECT 147.800 79.100 148.200 79.200 ;
        RECT 23.800 78.800 148.200 79.100 ;
        RECT 163.800 79.100 164.200 79.200 ;
        RECT 182.200 79.100 182.600 79.200 ;
        RECT 163.800 78.800 182.600 79.100 ;
        RECT 195.000 79.100 195.400 79.200 ;
        RECT 195.000 78.800 224.900 79.100 ;
        RECT 224.600 78.200 224.900 78.800 ;
        RECT 238.200 78.800 238.600 79.200 ;
        RECT 238.200 78.200 238.500 78.800 ;
        RECT 63.800 78.100 64.200 78.200 ;
        RECT 80.600 78.100 81.000 78.200 ;
        RECT 63.800 77.800 81.000 78.100 ;
        RECT 94.200 78.100 94.600 78.200 ;
        RECT 146.200 78.100 146.600 78.200 ;
        RECT 150.200 78.100 150.600 78.200 ;
        RECT 159.800 78.100 160.200 78.200 ;
        RECT 94.200 77.800 160.200 78.100 ;
        RECT 160.600 78.100 161.000 78.200 ;
        RECT 171.800 78.100 172.200 78.200 ;
        RECT 195.800 78.100 196.200 78.200 ;
        RECT 207.000 78.100 207.400 78.200 ;
        RECT 223.000 78.100 223.400 78.200 ;
        RECT 160.600 77.800 207.400 78.100 ;
        RECT 210.200 77.800 223.400 78.100 ;
        RECT 224.600 78.100 225.000 78.200 ;
        RECT 232.600 78.100 233.000 78.200 ;
        RECT 224.600 77.800 233.000 78.100 ;
        RECT 238.200 77.800 238.600 78.200 ;
        RECT 210.200 77.200 210.500 77.800 ;
        RECT 27.800 77.100 28.200 77.200 ;
        RECT 40.600 77.100 41.000 77.200 ;
        RECT 47.000 77.100 47.400 77.200 ;
        RECT 27.800 76.800 47.400 77.100 ;
        RECT 59.800 77.100 60.200 77.200 ;
        RECT 69.400 77.100 69.800 77.200 ;
        RECT 71.800 77.100 72.200 77.200 ;
        RECT 59.800 76.800 72.200 77.100 ;
        RECT 93.400 77.100 93.800 77.200 ;
        RECT 125.400 77.100 125.800 77.200 ;
        RECT 93.400 76.800 125.800 77.100 ;
        RECT 128.600 77.100 129.000 77.200 ;
        RECT 156.600 77.100 157.000 77.200 ;
        RECT 163.000 77.100 163.400 77.200 ;
        RECT 128.600 76.800 157.000 77.100 ;
        RECT 158.200 76.800 163.400 77.100 ;
        RECT 163.800 77.100 164.200 77.200 ;
        RECT 196.600 77.100 197.000 77.200 ;
        RECT 163.800 76.800 197.000 77.100 ;
        RECT 210.200 76.800 210.600 77.200 ;
        RECT 227.000 77.100 227.400 77.200 ;
        RECT 230.200 77.100 230.600 77.200 ;
        RECT 232.600 77.100 233.000 77.200 ;
        RECT 238.200 77.100 238.600 77.200 ;
        RECT 227.000 76.800 230.600 77.100 ;
        RECT 231.800 76.800 238.600 77.100 ;
        RECT 158.200 76.200 158.500 76.800 ;
        RECT 196.600 76.200 196.900 76.800 ;
        RECT 12.600 76.100 13.000 76.200 ;
        RECT 14.200 76.100 14.600 76.200 ;
        RECT 18.200 76.100 18.600 76.200 ;
        RECT 12.600 75.800 18.600 76.100 ;
        RECT 31.800 76.100 32.200 76.200 ;
        RECT 40.600 76.100 41.000 76.200 ;
        RECT 73.400 76.100 73.800 76.200 ;
        RECT 89.400 76.100 89.800 76.200 ;
        RECT 31.800 75.800 89.800 76.100 ;
        RECT 91.800 76.100 92.200 76.200 ;
        RECT 94.200 76.100 94.600 76.200 ;
        RECT 91.800 75.800 94.600 76.100 ;
        RECT 95.800 76.100 96.200 76.200 ;
        RECT 127.800 76.100 128.200 76.200 ;
        RECT 95.800 75.800 128.200 76.100 ;
        RECT 139.000 76.100 139.400 76.200 ;
        RECT 141.400 76.100 141.800 76.200 ;
        RECT 139.000 75.800 141.800 76.100 ;
        RECT 142.200 75.800 142.600 76.200 ;
        RECT 155.000 76.100 155.400 76.200 ;
        RECT 158.200 76.100 158.600 76.200 ;
        RECT 155.000 75.800 158.600 76.100 ;
        RECT 163.000 76.100 163.400 76.200 ;
        RECT 165.400 76.100 165.800 76.200 ;
        RECT 163.000 75.800 165.800 76.100 ;
        RECT 170.200 76.100 170.600 76.200 ;
        RECT 192.600 76.100 193.000 76.200 ;
        RECT 170.200 75.800 193.000 76.100 ;
        RECT 196.600 76.100 197.000 76.200 ;
        RECT 207.800 76.100 208.200 76.200 ;
        RECT 196.600 75.800 208.200 76.100 ;
        RECT 222.200 76.100 222.600 76.200 ;
        RECT 223.000 76.100 223.400 76.200 ;
        RECT 222.200 75.800 223.400 76.100 ;
        RECT 226.200 76.100 226.600 76.200 ;
        RECT 231.000 76.100 231.400 76.200 ;
        RECT 231.800 76.100 232.200 76.200 ;
        RECT 226.200 75.800 232.200 76.100 ;
        RECT 248.600 76.100 249.000 76.200 ;
        RECT 249.400 76.100 249.800 76.200 ;
        RECT 248.600 75.800 249.800 76.100 ;
        RECT 250.200 76.100 250.600 76.200 ;
        RECT 254.200 76.100 254.600 76.200 ;
        RECT 250.200 75.800 254.600 76.100 ;
        RECT 141.400 75.200 141.700 75.800 ;
        RECT 142.200 75.200 142.500 75.800 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 11.800 75.100 12.200 75.200 ;
        RECT 4.600 74.800 12.200 75.100 ;
        RECT 12.600 75.100 13.000 75.200 ;
        RECT 25.400 75.100 25.800 75.200 ;
        RECT 29.400 75.100 29.800 75.200 ;
        RECT 12.600 74.800 29.800 75.100 ;
        RECT 44.600 75.100 45.000 75.200 ;
        RECT 51.800 75.100 52.200 75.200 ;
        RECT 44.600 74.800 52.200 75.100 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 77.400 75.100 77.800 75.200 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 77.400 74.800 85.000 75.100 ;
        RECT 87.800 75.100 88.200 75.200 ;
        RECT 101.400 75.100 101.800 75.200 ;
        RECT 87.800 74.800 101.800 75.100 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 107.000 75.100 107.400 75.200 ;
        RECT 106.200 74.800 107.400 75.100 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 112.600 74.800 114.600 75.100 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 139.800 75.100 140.200 75.200 ;
        RECT 134.200 74.800 140.200 75.100 ;
        RECT 141.400 74.800 141.800 75.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 151.800 75.100 152.200 75.200 ;
        RECT 176.600 75.100 177.000 75.200 ;
        RECT 187.000 75.100 187.400 75.200 ;
        RECT 190.200 75.100 190.600 75.200 ;
        RECT 151.800 74.800 190.600 75.100 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 198.200 75.100 198.600 75.200 ;
        RECT 197.400 74.800 198.600 75.100 ;
        RECT 209.400 75.100 209.800 75.200 ;
        RECT 210.200 75.100 210.600 75.200 ;
        RECT 209.400 74.800 210.600 75.100 ;
        RECT 216.600 75.100 217.000 75.200 ;
        RECT 220.600 75.100 221.000 75.200 ;
        RECT 216.600 74.800 221.000 75.100 ;
        RECT 223.800 75.100 224.200 75.200 ;
        RECT 226.200 75.100 226.600 75.200 ;
        RECT 223.800 74.800 226.600 75.100 ;
        RECT 232.600 75.100 233.000 75.200 ;
        RECT 243.800 75.100 244.200 75.200 ;
        RECT 232.600 74.800 244.200 75.100 ;
        RECT 245.400 75.100 245.800 75.200 ;
        RECT 249.400 75.100 249.800 75.200 ;
        RECT 245.400 74.800 249.800 75.100 ;
        RECT 10.200 74.100 10.600 74.200 ;
        RECT 39.000 74.100 39.400 74.200 ;
        RECT 10.200 73.800 39.400 74.100 ;
        RECT 66.200 74.100 66.500 74.800 ;
        RECT 81.400 74.100 81.800 74.200 ;
        RECT 101.400 74.100 101.800 74.200 ;
        RECT 111.800 74.100 112.100 74.800 ;
        RECT 66.200 73.800 112.100 74.100 ;
        RECT 112.600 74.200 112.900 74.800 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 124.600 74.100 125.000 74.200 ;
        RECT 163.000 74.100 163.400 74.200 ;
        RECT 124.600 73.800 163.400 74.100 ;
        RECT 163.800 74.100 164.200 74.200 ;
        RECT 168.600 74.100 169.000 74.200 ;
        RECT 163.800 73.800 169.000 74.100 ;
        RECT 177.400 74.100 177.800 74.200 ;
        RECT 186.200 74.100 186.600 74.200 ;
        RECT 177.400 73.800 186.600 74.100 ;
        RECT 188.600 74.100 189.000 74.200 ;
        RECT 189.400 74.100 189.800 74.200 ;
        RECT 188.600 73.800 189.800 74.100 ;
        RECT 198.200 74.100 198.600 74.200 ;
        RECT 200.600 74.100 201.000 74.200 ;
        RECT 198.200 73.800 201.000 74.100 ;
        RECT 19.000 73.100 19.400 73.200 ;
        RECT 63.800 73.100 64.200 73.200 ;
        RECT 71.000 73.100 71.400 73.200 ;
        RECT 19.000 72.800 28.900 73.100 ;
        RECT 63.800 72.800 71.400 73.100 ;
        RECT 76.600 73.100 77.000 73.200 ;
        RECT 88.600 73.100 89.000 73.200 ;
        RECT 89.400 73.100 89.800 73.200 ;
        RECT 76.600 72.800 89.800 73.100 ;
        RECT 100.600 73.100 101.000 73.200 ;
        RECT 109.400 73.100 109.800 73.200 ;
        RECT 100.600 72.800 109.800 73.100 ;
        RECT 110.200 73.100 110.600 73.200 ;
        RECT 119.000 73.100 119.400 73.200 ;
        RECT 110.200 72.800 119.400 73.100 ;
        RECT 127.000 73.100 127.400 73.200 ;
        RECT 133.400 73.100 133.800 73.200 ;
        RECT 142.200 73.100 142.600 73.200 ;
        RECT 127.000 72.800 142.600 73.100 ;
        RECT 166.200 73.100 166.600 73.200 ;
        RECT 167.000 73.100 167.400 73.200 ;
        RECT 166.200 72.800 167.400 73.100 ;
        RECT 183.000 72.800 183.400 73.200 ;
        RECT 184.600 73.100 185.000 73.200 ;
        RECT 199.800 73.100 200.200 73.200 ;
        RECT 184.600 72.800 200.200 73.100 ;
        RECT 211.000 73.100 211.400 73.200 ;
        RECT 212.600 73.100 213.000 73.200 ;
        RECT 211.000 72.800 213.000 73.100 ;
        RECT 243.800 72.800 244.200 73.200 ;
        RECT 245.400 73.100 245.800 73.200 ;
        RECT 246.200 73.100 246.600 73.200 ;
        RECT 245.400 72.800 246.600 73.100 ;
        RECT 28.600 72.200 28.900 72.800 ;
        RECT 183.000 72.200 183.300 72.800 ;
        RECT 243.800 72.200 244.100 72.800 ;
        RECT 25.400 72.100 25.800 72.200 ;
        RECT 27.000 72.100 27.400 72.200 ;
        RECT 25.400 71.800 27.400 72.100 ;
        RECT 28.600 71.800 29.000 72.200 ;
        RECT 47.000 72.100 47.400 72.200 ;
        RECT 56.600 72.100 57.000 72.200 ;
        RECT 47.000 71.800 57.000 72.100 ;
        RECT 59.000 72.100 59.400 72.200 ;
        RECT 64.600 72.100 65.000 72.200 ;
        RECT 67.800 72.100 68.200 72.200 ;
        RECT 59.000 71.800 68.200 72.100 ;
        RECT 104.600 72.100 105.000 72.200 ;
        RECT 108.600 72.100 109.000 72.200 ;
        RECT 130.200 72.100 130.600 72.200 ;
        RECT 104.600 71.800 130.600 72.100 ;
        RECT 161.400 72.100 161.800 72.200 ;
        RECT 170.200 72.100 170.600 72.200 ;
        RECT 161.400 71.800 170.600 72.100 ;
        RECT 183.000 71.800 183.400 72.200 ;
        RECT 187.000 72.100 187.400 72.200 ;
        RECT 191.000 72.100 191.400 72.200 ;
        RECT 223.000 72.100 223.400 72.200 ;
        RECT 229.400 72.100 229.800 72.200 ;
        RECT 187.000 71.800 229.800 72.100 ;
        RECT 243.800 71.800 244.200 72.200 ;
        RECT 247.000 72.100 247.400 72.200 ;
        RECT 249.400 72.100 249.800 72.200 ;
        RECT 247.000 71.800 249.800 72.100 ;
        RECT 256.600 72.100 257.000 72.200 ;
        RECT 257.400 72.100 257.800 72.200 ;
        RECT 256.600 71.800 257.800 72.100 ;
        RECT 18.200 71.100 18.600 71.200 ;
        RECT 33.400 71.100 33.800 71.200 ;
        RECT 18.200 70.800 33.800 71.100 ;
        RECT 34.200 71.100 34.600 71.200 ;
        RECT 70.200 71.100 70.600 71.200 ;
        RECT 95.000 71.100 95.400 71.200 ;
        RECT 34.200 70.800 70.600 71.100 ;
        RECT 91.000 70.800 95.400 71.100 ;
        RECT 159.800 71.100 160.200 71.200 ;
        RECT 165.400 71.100 165.800 71.200 ;
        RECT 159.800 70.800 165.800 71.100 ;
        RECT 166.200 71.100 166.600 71.200 ;
        RECT 173.400 71.100 173.800 71.200 ;
        RECT 166.200 70.800 173.800 71.100 ;
        RECT 179.800 71.100 180.200 71.200 ;
        RECT 188.600 71.100 189.000 71.200 ;
        RECT 179.800 70.800 189.000 71.100 ;
        RECT 215.800 71.100 216.200 71.200 ;
        RECT 223.800 71.100 224.200 71.200 ;
        RECT 215.800 70.800 224.200 71.100 ;
        RECT 229.400 71.100 229.800 71.200 ;
        RECT 231.800 71.100 232.200 71.200 ;
        RECT 229.400 70.800 232.200 71.100 ;
        RECT 27.000 70.100 27.400 70.200 ;
        RECT 44.600 70.100 45.000 70.200 ;
        RECT 27.000 69.800 45.000 70.100 ;
        RECT 53.400 70.100 53.800 70.200 ;
        RECT 91.000 70.100 91.300 70.800 ;
        RECT 53.400 69.800 91.300 70.100 ;
        RECT 91.800 70.100 92.200 70.200 ;
        RECT 95.000 70.100 95.400 70.200 ;
        RECT 91.800 69.800 95.400 70.100 ;
        RECT 108.600 70.100 109.000 70.200 ;
        RECT 113.400 70.100 113.800 70.200 ;
        RECT 134.200 70.100 134.600 70.200 ;
        RECT 108.600 69.800 134.600 70.100 ;
        RECT 142.200 70.100 142.600 70.200 ;
        RECT 174.200 70.100 174.600 70.200 ;
        RECT 189.400 70.100 189.800 70.200 ;
        RECT 142.200 69.800 189.800 70.100 ;
        RECT 197.400 70.100 197.800 70.200 ;
        RECT 206.200 70.100 206.600 70.200 ;
        RECT 207.000 70.100 207.400 70.200 ;
        RECT 197.400 69.800 207.400 70.100 ;
        RECT 19.800 69.100 20.200 69.200 ;
        RECT 25.400 69.100 25.800 69.200 ;
        RECT 19.800 68.800 25.800 69.100 ;
        RECT 29.400 69.100 29.800 69.200 ;
        RECT 47.000 69.100 47.400 69.200 ;
        RECT 29.400 68.800 47.400 69.100 ;
        RECT 54.200 69.100 54.600 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 54.200 68.800 59.400 69.100 ;
        RECT 89.400 69.100 89.800 69.200 ;
        RECT 95.000 69.100 95.400 69.200 ;
        RECT 107.000 69.100 107.400 69.200 ;
        RECT 89.400 68.800 107.400 69.100 ;
        RECT 127.800 69.100 128.200 69.200 ;
        RECT 129.400 69.100 129.800 69.200 ;
        RECT 127.800 68.800 129.800 69.100 ;
        RECT 131.800 69.100 132.200 69.200 ;
        RECT 140.600 69.100 141.000 69.200 ;
        RECT 131.800 68.800 141.000 69.100 ;
        RECT 155.800 69.100 156.200 69.200 ;
        RECT 160.600 69.100 161.000 69.200 ;
        RECT 164.600 69.100 165.000 69.200 ;
        RECT 155.800 68.800 165.000 69.100 ;
        RECT 166.200 69.100 166.600 69.200 ;
        RECT 169.400 69.100 169.800 69.200 ;
        RECT 166.200 68.800 169.800 69.100 ;
        RECT 171.800 69.100 172.200 69.200 ;
        RECT 172.600 69.100 173.000 69.200 ;
        RECT 180.600 69.100 181.000 69.200 ;
        RECT 171.800 68.800 181.000 69.100 ;
        RECT 203.000 69.100 203.400 69.200 ;
        RECT 219.800 69.100 220.200 69.200 ;
        RECT 203.000 68.800 220.200 69.100 ;
        RECT 227.800 69.100 228.200 69.200 ;
        RECT 242.200 69.100 242.600 69.200 ;
        RECT 227.800 68.800 242.600 69.100 ;
        RECT 243.000 69.100 243.400 69.200 ;
        RECT 255.000 69.100 255.400 69.200 ;
        RECT 243.000 68.800 255.400 69.100 ;
        RECT 23.800 68.100 24.200 68.200 ;
        RECT 29.400 68.100 29.800 68.200 ;
        RECT 23.800 67.800 29.800 68.100 ;
        RECT 35.800 68.100 36.200 68.200 ;
        RECT 37.400 68.100 37.800 68.200 ;
        RECT 35.800 67.800 37.800 68.100 ;
        RECT 39.800 68.100 40.200 68.200 ;
        RECT 40.600 68.100 41.000 68.200 ;
        RECT 39.800 67.800 41.000 68.100 ;
        RECT 51.800 68.100 52.200 68.200 ;
        RECT 76.600 68.100 77.000 68.200 ;
        RECT 51.800 67.800 77.000 68.100 ;
        RECT 83.000 68.100 83.400 68.200 ;
        RECT 91.800 68.100 92.200 68.200 ;
        RECT 83.000 67.800 92.200 68.100 ;
        RECT 98.200 68.100 98.600 68.200 ;
        RECT 128.600 68.100 129.000 68.200 ;
        RECT 129.400 68.100 129.800 68.200 ;
        RECT 98.200 67.800 127.300 68.100 ;
        RECT 128.600 67.800 129.800 68.100 ;
        RECT 151.000 68.100 151.400 68.200 ;
        RECT 158.200 68.100 158.600 68.200 ;
        RECT 151.000 67.800 158.600 68.100 ;
        RECT 162.200 67.800 162.600 68.200 ;
        RECT 164.600 67.800 165.000 68.200 ;
        RECT 167.800 68.100 168.200 68.200 ;
        RECT 197.400 68.100 197.800 68.200 ;
        RECT 167.800 67.800 197.800 68.100 ;
        RECT 205.400 68.100 205.800 68.200 ;
        RECT 217.400 68.100 217.800 68.200 ;
        RECT 205.400 67.800 217.800 68.100 ;
        RECT 224.600 68.100 225.000 68.200 ;
        RECT 238.200 68.100 238.600 68.200 ;
        RECT 224.600 67.800 238.600 68.100 ;
        RECT 240.600 68.100 241.000 68.200 ;
        RECT 245.400 68.100 245.800 68.200 ;
        RECT 240.600 67.800 245.800 68.100 ;
        RECT 247.800 67.800 248.200 68.200 ;
        RECT 251.000 68.100 251.400 68.200 ;
        RECT 252.600 68.100 253.000 68.200 ;
        RECT 251.000 67.800 253.000 68.100 ;
        RECT 127.000 67.200 127.300 67.800 ;
        RECT 0.600 67.100 1.000 67.200 ;
        RECT 13.400 67.100 13.800 67.200 ;
        RECT 23.800 67.100 24.200 67.200 ;
        RECT 0.600 66.800 8.100 67.100 ;
        RECT 13.400 66.800 24.200 67.100 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 27.800 67.100 28.200 67.200 ;
        RECT 26.200 66.800 28.200 67.100 ;
        RECT 35.000 66.800 35.400 67.200 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 69.400 67.100 69.800 67.200 ;
        RECT 77.400 67.100 77.800 67.200 ;
        RECT 69.400 66.800 77.800 67.100 ;
        RECT 89.400 66.800 89.800 67.200 ;
        RECT 95.800 67.100 96.200 67.200 ;
        RECT 106.200 67.100 106.600 67.200 ;
        RECT 111.800 67.100 112.200 67.200 ;
        RECT 95.800 66.800 112.200 67.100 ;
        RECT 114.200 66.800 114.600 67.200 ;
        RECT 120.600 67.100 121.000 67.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 120.600 66.800 121.800 67.100 ;
        RECT 122.200 67.100 122.600 67.200 ;
        RECT 125.400 67.100 125.800 67.200 ;
        RECT 122.200 66.800 125.800 67.100 ;
        RECT 127.000 67.100 127.400 67.200 ;
        RECT 131.800 67.100 132.200 67.200 ;
        RECT 127.000 66.800 132.200 67.100 ;
        RECT 133.400 66.800 133.800 67.200 ;
        RECT 136.600 66.800 137.000 67.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 149.400 66.800 149.800 67.200 ;
        RECT 150.200 67.100 150.600 67.200 ;
        RECT 151.800 67.100 152.200 67.200 ;
        RECT 150.200 66.800 152.200 67.100 ;
        RECT 162.200 67.100 162.500 67.800 ;
        RECT 164.600 67.100 164.900 67.800 ;
        RECT 162.200 66.800 164.900 67.100 ;
        RECT 167.800 67.200 168.100 67.800 ;
        RECT 247.800 67.200 248.100 67.800 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 170.200 66.800 170.600 67.200 ;
        RECT 177.400 67.100 177.800 67.200 ;
        RECT 183.800 67.100 184.200 67.200 ;
        RECT 177.400 66.800 184.200 67.100 ;
        RECT 199.800 67.100 200.200 67.200 ;
        RECT 211.800 67.100 212.200 67.200 ;
        RECT 199.800 66.800 212.200 67.100 ;
        RECT 212.600 67.100 213.000 67.200 ;
        RECT 225.400 67.100 225.800 67.200 ;
        RECT 212.600 66.800 225.800 67.100 ;
        RECT 229.400 67.100 229.800 67.200 ;
        RECT 247.800 67.100 248.200 67.200 ;
        RECT 229.400 66.800 248.200 67.100 ;
        RECT 248.600 67.100 249.000 67.200 ;
        RECT 255.800 67.100 256.200 67.200 ;
        RECT 248.600 66.800 256.200 67.100 ;
        RECT 7.800 66.200 8.100 66.800 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 50.200 66.200 50.500 66.800 ;
        RECT 64.600 66.200 64.900 66.800 ;
        RECT 65.400 66.200 65.700 66.800 ;
        RECT 66.200 66.200 66.500 66.800 ;
        RECT 7.800 65.800 8.200 66.200 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 28.600 66.100 29.000 66.200 ;
        RECT 8.600 65.800 29.000 66.100 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 39.000 66.100 39.400 66.200 ;
        RECT 48.600 66.100 49.000 66.200 ;
        RECT 39.000 65.800 49.000 66.100 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 55.800 65.800 57.000 66.100 ;
        RECT 57.400 66.100 57.800 66.200 ;
        RECT 58.200 66.100 58.600 66.200 ;
        RECT 57.400 65.800 58.600 66.100 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 73.400 65.800 74.600 66.100 ;
        RECT 89.400 66.100 89.700 66.800 ;
        RECT 90.200 66.100 90.600 66.200 ;
        RECT 91.800 66.100 92.200 66.200 ;
        RECT 89.400 65.800 92.200 66.100 ;
        RECT 93.400 66.100 93.800 66.200 ;
        RECT 95.000 66.100 95.400 66.200 ;
        RECT 93.400 65.800 95.400 66.100 ;
        RECT 96.600 66.100 97.000 66.200 ;
        RECT 109.400 66.100 109.800 66.200 ;
        RECT 96.600 65.800 109.800 66.100 ;
        RECT 111.000 66.100 111.400 66.200 ;
        RECT 114.200 66.100 114.500 66.800 ;
        RECT 133.400 66.200 133.700 66.800 ;
        RECT 136.600 66.200 136.900 66.800 ;
        RECT 137.400 66.200 137.700 66.800 ;
        RECT 149.400 66.200 149.700 66.800 ;
        RECT 169.400 66.200 169.700 66.800 ;
        RECT 170.200 66.200 170.500 66.800 ;
        RECT 199.800 66.200 200.100 66.800 ;
        RECT 248.600 66.200 248.900 66.800 ;
        RECT 111.000 65.800 114.500 66.100 ;
        RECT 117.400 66.100 117.800 66.200 ;
        RECT 124.600 66.100 125.000 66.200 ;
        RECT 117.400 65.800 125.000 66.100 ;
        RECT 125.400 66.100 125.800 66.200 ;
        RECT 126.200 66.100 126.600 66.200 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 125.400 65.800 130.600 66.100 ;
        RECT 133.400 65.800 133.800 66.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 138.200 66.100 138.600 66.200 ;
        RECT 146.200 66.100 146.600 66.200 ;
        RECT 148.600 66.100 149.000 66.200 ;
        RECT 138.200 65.800 149.000 66.100 ;
        RECT 149.400 66.100 149.800 66.200 ;
        RECT 158.200 66.100 158.600 66.200 ;
        RECT 149.400 65.800 158.600 66.100 ;
        RECT 166.200 66.100 166.600 66.200 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 166.200 65.800 168.200 66.100 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 182.200 66.100 182.600 66.200 ;
        RECT 183.800 66.100 184.200 66.200 ;
        RECT 182.200 65.800 184.200 66.100 ;
        RECT 195.800 66.100 196.200 66.200 ;
        RECT 196.600 66.100 197.000 66.200 ;
        RECT 195.800 65.800 197.000 66.100 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 202.200 66.100 202.600 66.200 ;
        RECT 203.000 66.100 203.400 66.200 ;
        RECT 214.200 66.100 214.600 66.200 ;
        RECT 202.200 65.800 214.600 66.100 ;
        RECT 219.000 65.800 219.400 66.200 ;
        RECT 231.800 66.100 232.200 66.200 ;
        RECT 231.800 65.800 242.500 66.100 ;
        RECT 248.600 65.800 249.000 66.200 ;
        RECT 250.200 65.800 250.600 66.200 ;
        RECT 251.800 66.100 252.200 66.200 ;
        RECT 254.200 66.100 254.600 66.200 ;
        RECT 251.800 65.800 254.600 66.100 ;
        RECT 219.000 65.200 219.300 65.800 ;
        RECT 242.200 65.200 242.500 65.800 ;
        RECT 15.800 65.100 16.200 65.200 ;
        RECT 24.600 65.100 25.000 65.200 ;
        RECT 35.800 65.100 36.200 65.200 ;
        RECT 15.800 64.800 36.200 65.100 ;
        RECT 54.200 65.100 54.600 65.200 ;
        RECT 79.000 65.100 79.400 65.200 ;
        RECT 54.200 64.800 79.400 65.100 ;
        RECT 90.200 65.100 90.600 65.200 ;
        RECT 91.000 65.100 91.400 65.200 ;
        RECT 90.200 64.800 91.400 65.100 ;
        RECT 96.600 65.100 97.000 65.200 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 96.600 64.800 103.400 65.100 ;
        RECT 103.800 65.100 104.200 65.200 ;
        RECT 118.200 65.100 118.600 65.200 ;
        RECT 135.800 65.100 136.200 65.200 ;
        RECT 103.800 64.800 136.200 65.100 ;
        RECT 141.400 65.100 141.800 65.200 ;
        RECT 152.600 65.100 153.000 65.200 ;
        RECT 141.400 64.800 153.000 65.100 ;
        RECT 167.000 64.800 167.400 65.200 ;
        RECT 206.200 65.100 206.600 65.200 ;
        RECT 208.600 65.100 209.000 65.200 ;
        RECT 206.200 64.800 209.000 65.100 ;
        RECT 219.000 64.800 219.400 65.200 ;
        RECT 242.200 64.800 242.600 65.200 ;
        RECT 243.800 65.100 244.200 65.200 ;
        RECT 250.200 65.100 250.500 65.800 ;
        RECT 260.600 65.100 261.000 65.200 ;
        RECT 243.800 64.800 250.500 65.100 ;
        RECT 254.200 64.800 261.000 65.100 ;
        RECT 167.000 64.200 167.300 64.800 ;
        RECT 254.200 64.200 254.500 64.800 ;
        RECT 17.400 64.100 17.800 64.200 ;
        RECT 33.400 64.100 33.800 64.200 ;
        RECT 17.400 63.800 33.800 64.100 ;
        RECT 35.800 64.100 36.200 64.200 ;
        RECT 42.200 64.100 42.600 64.200 ;
        RECT 35.800 63.800 42.600 64.100 ;
        RECT 43.000 64.100 43.400 64.200 ;
        RECT 45.400 64.100 45.800 64.200 ;
        RECT 43.000 63.800 45.800 64.100 ;
        RECT 47.800 64.100 48.200 64.200 ;
        RECT 48.600 64.100 49.000 64.200 ;
        RECT 47.800 63.800 49.000 64.100 ;
        RECT 53.400 64.100 53.800 64.200 ;
        RECT 71.800 64.100 72.200 64.200 ;
        RECT 53.400 63.800 72.200 64.100 ;
        RECT 78.200 63.800 78.600 64.200 ;
        RECT 91.800 64.100 92.200 64.200 ;
        RECT 100.600 64.100 101.000 64.200 ;
        RECT 91.800 63.800 101.000 64.100 ;
        RECT 107.800 64.100 108.200 64.200 ;
        RECT 112.600 64.100 113.000 64.200 ;
        RECT 121.400 64.100 121.800 64.200 ;
        RECT 107.800 63.800 121.800 64.100 ;
        RECT 124.600 64.100 125.000 64.200 ;
        RECT 137.400 64.100 137.800 64.200 ;
        RECT 155.800 64.100 156.200 64.200 ;
        RECT 124.600 63.800 126.500 64.100 ;
        RECT 137.400 63.800 156.200 64.100 ;
        RECT 167.000 63.800 167.400 64.200 ;
        RECT 212.600 64.100 213.000 64.200 ;
        RECT 211.000 63.800 213.000 64.100 ;
        RECT 254.200 63.800 254.600 64.200 ;
        RECT 33.400 63.100 33.800 63.200 ;
        RECT 51.000 63.100 51.400 63.200 ;
        RECT 32.600 62.800 51.400 63.100 ;
        RECT 51.800 63.100 52.200 63.200 ;
        RECT 62.200 63.100 62.600 63.200 ;
        RECT 51.800 62.800 62.600 63.100 ;
        RECT 78.200 63.100 78.500 63.800 ;
        RECT 126.200 63.200 126.500 63.800 ;
        RECT 211.000 63.200 211.300 63.800 ;
        RECT 123.000 63.100 123.400 63.200 ;
        RECT 78.200 62.800 123.400 63.100 ;
        RECT 126.200 62.800 126.600 63.200 ;
        RECT 155.000 63.100 155.400 63.200 ;
        RECT 171.800 63.100 172.200 63.200 ;
        RECT 155.000 62.800 172.200 63.100 ;
        RECT 191.000 63.100 191.400 63.200 ;
        RECT 205.400 63.100 205.800 63.200 ;
        RECT 191.000 62.800 205.800 63.100 ;
        RECT 211.000 62.800 211.400 63.200 ;
        RECT 211.800 63.100 212.200 63.200 ;
        RECT 227.000 63.100 227.400 63.200 ;
        RECT 211.800 62.800 227.400 63.100 ;
        RECT 246.200 63.100 246.600 63.200 ;
        RECT 255.800 63.100 256.200 63.200 ;
        RECT 246.200 62.800 256.200 63.100 ;
        RECT 45.400 62.100 45.800 62.200 ;
        RECT 79.800 62.100 80.200 62.200 ;
        RECT 89.400 62.100 89.800 62.200 ;
        RECT 45.400 61.800 89.800 62.100 ;
        RECT 103.800 62.100 104.200 62.200 ;
        RECT 137.400 62.100 137.800 62.200 ;
        RECT 161.400 62.100 161.800 62.200 ;
        RECT 103.800 61.800 137.800 62.100 ;
        RECT 155.000 61.800 161.800 62.100 ;
        RECT 179.800 62.100 180.200 62.200 ;
        RECT 216.600 62.100 217.000 62.200 ;
        RECT 232.600 62.100 233.000 62.200 ;
        RECT 179.800 61.800 233.000 62.100 ;
        RECT 249.400 62.100 249.800 62.200 ;
        RECT 251.000 62.100 251.400 62.200 ;
        RECT 249.400 61.800 251.400 62.100 ;
        RECT 44.600 61.100 45.000 61.200 ;
        RECT 53.400 61.100 53.800 61.200 ;
        RECT 44.600 60.800 53.800 61.100 ;
        RECT 103.000 61.100 103.400 61.200 ;
        RECT 131.000 61.100 131.400 61.200 ;
        RECT 103.000 60.800 131.400 61.100 ;
        RECT 136.600 61.100 137.000 61.200 ;
        RECT 155.000 61.100 155.300 61.800 ;
        RECT 136.600 60.800 155.300 61.100 ;
        RECT 159.000 61.100 159.400 61.200 ;
        RECT 196.600 61.100 197.000 61.200 ;
        RECT 211.000 61.100 211.400 61.200 ;
        RECT 159.000 60.800 211.400 61.100 ;
        RECT 139.000 60.100 139.400 60.200 ;
        RECT 139.800 60.100 140.200 60.200 ;
        RECT 139.000 59.800 140.200 60.100 ;
        RECT 158.200 60.100 158.600 60.200 ;
        RECT 235.800 60.100 236.200 60.200 ;
        RECT 158.200 59.800 236.200 60.100 ;
        RECT 25.400 59.100 25.800 59.200 ;
        RECT 94.200 59.100 94.600 59.200 ;
        RECT 25.400 58.800 94.600 59.100 ;
        RECT 143.000 59.100 143.400 59.200 ;
        RECT 159.000 59.100 159.400 59.200 ;
        RECT 143.000 58.800 159.400 59.100 ;
        RECT 163.800 59.100 164.200 59.200 ;
        RECT 190.200 59.100 190.600 59.200 ;
        RECT 193.400 59.100 193.800 59.200 ;
        RECT 163.800 58.800 193.800 59.100 ;
        RECT 195.800 59.100 196.200 59.200 ;
        RECT 225.400 59.100 225.800 59.200 ;
        RECT 243.000 59.100 243.400 59.200 ;
        RECT 195.800 58.800 243.400 59.100 ;
        RECT 30.200 58.100 30.600 58.200 ;
        RECT 40.600 58.100 41.000 58.200 ;
        RECT 41.400 58.100 41.800 58.200 ;
        RECT 57.400 58.100 57.800 58.200 ;
        RECT 30.200 57.800 57.800 58.100 ;
        RECT 68.600 58.100 69.000 58.200 ;
        RECT 69.400 58.100 69.800 58.200 ;
        RECT 68.600 57.800 69.800 58.100 ;
        RECT 73.400 57.800 73.800 58.200 ;
        RECT 83.800 58.100 84.200 58.200 ;
        RECT 88.600 58.100 89.000 58.200 ;
        RECT 104.600 58.100 105.000 58.200 ;
        RECT 83.800 57.800 105.000 58.100 ;
        RECT 128.600 58.100 129.000 58.200 ;
        RECT 139.800 58.100 140.200 58.200 ;
        RECT 128.600 57.800 140.200 58.100 ;
        RECT 175.800 58.100 176.200 58.200 ;
        RECT 206.200 58.100 206.600 58.200 ;
        RECT 175.800 57.800 206.600 58.100 ;
        RECT 255.000 58.100 255.400 58.200 ;
        RECT 260.600 58.100 261.000 58.200 ;
        RECT 255.000 57.800 261.000 58.100 ;
        RECT 73.400 57.200 73.700 57.800 ;
        RECT 27.000 57.100 27.400 57.200 ;
        RECT 41.400 57.100 41.800 57.200 ;
        RECT 43.000 57.100 43.400 57.200 ;
        RECT 27.000 56.800 43.400 57.100 ;
        RECT 67.800 56.800 68.200 57.200 ;
        RECT 69.400 57.100 69.800 57.200 ;
        RECT 73.400 57.100 73.800 57.200 ;
        RECT 69.400 56.800 73.800 57.100 ;
        RECT 75.000 57.100 75.400 57.200 ;
        RECT 87.000 57.100 87.400 57.200 ;
        RECT 90.200 57.100 90.600 57.200 ;
        RECT 75.000 56.800 90.600 57.100 ;
        RECT 102.200 57.100 102.600 57.200 ;
        RECT 113.400 57.100 113.800 57.200 ;
        RECT 102.200 56.800 113.800 57.100 ;
        RECT 130.200 56.800 130.600 57.200 ;
        RECT 134.200 57.100 134.600 57.200 ;
        RECT 139.000 57.100 139.400 57.200 ;
        RECT 143.800 57.100 144.200 57.200 ;
        RECT 134.200 56.800 144.200 57.100 ;
        RECT 152.600 57.100 153.000 57.200 ;
        RECT 160.600 57.100 161.000 57.200 ;
        RECT 163.000 57.100 163.400 57.200 ;
        RECT 152.600 56.800 163.400 57.100 ;
        RECT 169.400 57.100 169.800 57.200 ;
        RECT 174.200 57.100 174.600 57.200 ;
        RECT 187.000 57.100 187.400 57.200 ;
        RECT 169.400 56.800 187.400 57.100 ;
        RECT 199.000 56.800 199.400 57.200 ;
        RECT 201.400 57.100 201.800 57.200 ;
        RECT 227.000 57.100 227.400 57.200 ;
        RECT 201.400 56.800 227.400 57.100 ;
        RECT 242.200 57.100 242.600 57.200 ;
        RECT 253.400 57.100 253.800 57.200 ;
        RECT 242.200 56.800 253.800 57.100 ;
        RECT 259.000 57.100 259.400 57.200 ;
        RECT 263.000 57.100 263.400 57.200 ;
        RECT 259.000 56.800 263.400 57.100 ;
        RECT 67.800 56.200 68.100 56.800 ;
        RECT 130.200 56.200 130.500 56.800 ;
        RECT 15.000 55.800 15.400 56.200 ;
        RECT 16.600 56.100 17.000 56.200 ;
        RECT 29.400 56.100 29.800 56.200 ;
        RECT 16.600 55.800 29.800 56.100 ;
        RECT 42.200 55.800 42.600 56.200 ;
        RECT 51.000 56.100 51.400 56.200 ;
        RECT 59.800 56.100 60.200 56.200 ;
        RECT 51.000 55.800 60.200 56.100 ;
        RECT 67.800 55.800 68.200 56.200 ;
        RECT 94.200 56.100 94.600 56.200 ;
        RECT 111.800 56.100 112.200 56.200 ;
        RECT 68.600 55.800 94.600 56.100 ;
        RECT 110.200 55.800 112.200 56.100 ;
        RECT 130.200 56.100 130.600 56.200 ;
        RECT 132.600 56.100 133.000 56.200 ;
        RECT 130.200 55.800 133.000 56.100 ;
        RECT 138.200 55.800 138.600 56.200 ;
        RECT 157.400 56.100 157.800 56.200 ;
        RECT 164.600 56.100 165.000 56.200 ;
        RECT 157.400 55.800 165.000 56.100 ;
        RECT 176.600 56.100 177.000 56.200 ;
        RECT 179.000 56.100 179.400 56.200 ;
        RECT 176.600 55.800 179.400 56.100 ;
        RECT 199.000 56.100 199.300 56.800 ;
        RECT 202.200 56.100 202.600 56.200 ;
        RECT 199.000 55.800 202.600 56.100 ;
        RECT 209.400 56.100 209.800 56.200 ;
        RECT 218.200 56.100 218.600 56.200 ;
        RECT 209.400 55.800 218.600 56.100 ;
        RECT 229.400 56.100 229.800 56.200 ;
        RECT 230.200 56.100 230.600 56.200 ;
        RECT 234.200 56.100 234.600 56.200 ;
        RECT 229.400 55.800 234.600 56.100 ;
        RECT 236.600 56.100 237.000 56.200 ;
        RECT 240.600 56.100 241.000 56.200 ;
        RECT 236.600 55.800 241.000 56.100 ;
        RECT 259.000 56.100 259.400 56.200 ;
        RECT 259.800 56.100 260.200 56.200 ;
        RECT 259.000 55.800 260.200 56.100 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 15.000 55.100 15.300 55.800 ;
        RECT 19.800 55.100 20.200 55.200 ;
        RECT 15.000 54.800 20.200 55.100 ;
        RECT 20.600 54.800 21.000 55.200 ;
        RECT 23.800 55.100 24.200 55.200 ;
        RECT 31.000 55.100 31.400 55.200 ;
        RECT 23.800 54.800 31.400 55.100 ;
        RECT 42.200 55.100 42.500 55.800 ;
        RECT 68.600 55.100 68.900 55.800 ;
        RECT 94.200 55.200 94.500 55.800 ;
        RECT 110.200 55.200 110.500 55.800 ;
        RECT 42.200 54.800 68.900 55.100 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 84.600 55.100 85.000 55.200 ;
        RECT 79.800 54.800 85.000 55.100 ;
        RECT 88.600 55.100 89.000 55.200 ;
        RECT 89.400 55.100 89.800 55.200 ;
        RECT 88.600 54.800 89.800 55.100 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 108.600 55.100 109.000 55.200 ;
        RECT 102.200 54.800 109.000 55.100 ;
        RECT 110.200 54.800 110.600 55.200 ;
        RECT 111.000 55.100 111.400 55.200 ;
        RECT 112.600 55.100 113.000 55.200 ;
        RECT 115.000 55.100 115.400 55.200 ;
        RECT 111.000 54.800 115.400 55.100 ;
        RECT 117.400 54.800 117.800 55.200 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 131.000 55.100 131.400 55.200 ;
        RECT 123.800 54.800 131.400 55.100 ;
        RECT 138.200 55.100 138.500 55.800 ;
        RECT 176.600 55.200 176.900 55.800 ;
        RECT 142.200 55.100 142.600 55.200 ;
        RECT 138.200 54.800 142.600 55.100 ;
        RECT 152.600 55.100 153.000 55.200 ;
        RECT 162.200 55.100 162.600 55.200 ;
        RECT 152.600 54.800 162.600 55.100 ;
        RECT 171.000 55.100 171.400 55.200 ;
        RECT 175.000 55.100 175.400 55.200 ;
        RECT 171.000 54.800 175.400 55.100 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 177.400 55.100 177.800 55.200 ;
        RECT 184.600 55.100 185.000 55.200 ;
        RECT 177.400 54.800 185.000 55.100 ;
        RECT 194.200 55.100 194.600 55.200 ;
        RECT 200.600 55.100 201.000 55.200 ;
        RECT 194.200 54.800 201.000 55.100 ;
        RECT 210.200 55.100 210.600 55.200 ;
        RECT 223.000 55.100 223.400 55.200 ;
        RECT 231.000 55.100 231.400 55.200 ;
        RECT 247.800 55.100 248.200 55.200 ;
        RECT 251.000 55.100 251.400 55.200 ;
        RECT 210.200 54.800 214.600 55.100 ;
        RECT 223.000 54.800 226.500 55.100 ;
        RECT 231.000 54.800 251.400 55.100 ;
        RECT 255.000 55.100 255.400 55.200 ;
        RECT 257.400 55.100 257.800 55.200 ;
        RECT 255.000 54.800 257.800 55.100 ;
        RECT 7.000 54.100 7.300 54.800 ;
        RECT 20.600 54.100 20.900 54.800 ;
        RECT 102.200 54.200 102.500 54.800 ;
        RECT 7.000 53.800 20.900 54.100 ;
        RECT 35.000 54.100 35.400 54.200 ;
        RECT 43.000 54.100 43.400 54.200 ;
        RECT 35.000 53.800 43.400 54.100 ;
        RECT 47.000 54.100 47.400 54.200 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 47.000 53.800 63.400 54.100 ;
        RECT 67.000 54.100 67.400 54.200 ;
        RECT 71.800 54.100 72.200 54.200 ;
        RECT 67.000 53.800 72.200 54.100 ;
        RECT 86.200 54.100 86.600 54.200 ;
        RECT 92.600 54.100 93.000 54.200 ;
        RECT 86.200 53.800 93.000 54.100 ;
        RECT 102.200 53.800 102.600 54.200 ;
        RECT 115.000 54.100 115.400 54.200 ;
        RECT 117.400 54.100 117.700 54.800 ;
        RECT 214.200 54.700 214.600 54.800 ;
        RECT 226.200 54.200 226.500 54.800 ;
        RECT 115.000 53.800 117.700 54.100 ;
        RECT 135.800 54.100 136.200 54.200 ;
        RECT 169.400 54.100 169.800 54.200 ;
        RECT 135.800 53.800 169.800 54.100 ;
        RECT 170.200 54.100 170.600 54.200 ;
        RECT 179.800 54.100 180.200 54.200 ;
        RECT 170.200 53.800 180.200 54.100 ;
        RECT 194.200 54.100 194.600 54.200 ;
        RECT 224.600 54.100 225.000 54.200 ;
        RECT 194.200 53.800 225.000 54.100 ;
        RECT 226.200 53.800 226.600 54.200 ;
        RECT 228.600 54.100 229.000 54.200 ;
        RECT 231.800 54.100 232.200 54.200 ;
        RECT 228.600 53.800 232.200 54.100 ;
        RECT 245.400 54.100 245.800 54.200 ;
        RECT 248.600 54.100 249.000 54.200 ;
        RECT 245.400 53.800 249.000 54.100 ;
        RECT 256.600 54.100 257.000 54.200 ;
        RECT 259.800 54.100 260.200 54.200 ;
        RECT 256.600 53.800 260.200 54.100 ;
        RECT 10.200 53.100 10.600 53.200 ;
        RECT 15.800 53.100 16.200 53.200 ;
        RECT 10.200 52.800 16.200 53.100 ;
        RECT 55.800 53.100 56.200 53.200 ;
        RECT 62.200 53.100 62.600 53.200 ;
        RECT 63.800 53.100 64.200 53.200 ;
        RECT 55.800 52.800 64.200 53.100 ;
        RECT 103.800 53.100 104.200 53.200 ;
        RECT 112.600 53.100 113.000 53.200 ;
        RECT 103.800 52.800 113.000 53.100 ;
        RECT 142.200 53.100 142.600 53.200 ;
        RECT 151.800 53.100 152.200 53.200 ;
        RECT 142.200 52.800 152.200 53.100 ;
        RECT 173.400 53.100 173.800 53.200 ;
        RECT 177.400 53.100 177.800 53.200 ;
        RECT 173.400 52.800 177.800 53.100 ;
        RECT 195.000 53.100 195.400 53.200 ;
        RECT 211.800 53.100 212.200 53.200 ;
        RECT 233.400 53.100 233.800 53.200 ;
        RECT 239.000 53.100 239.400 53.200 ;
        RECT 195.000 52.800 239.400 53.100 ;
        RECT 15.000 52.100 15.400 52.200 ;
        RECT 24.600 52.100 25.000 52.200 ;
        RECT 15.000 51.800 25.000 52.100 ;
        RECT 29.400 52.100 29.800 52.200 ;
        RECT 35.000 52.100 35.400 52.200 ;
        RECT 29.400 51.800 35.400 52.100 ;
        RECT 40.600 52.100 41.000 52.200 ;
        RECT 69.400 52.100 69.800 52.200 ;
        RECT 40.600 51.800 69.800 52.100 ;
        RECT 91.000 52.100 91.400 52.200 ;
        RECT 146.200 52.100 146.600 52.200 ;
        RECT 91.000 51.800 146.600 52.100 ;
        RECT 147.000 52.100 147.400 52.200 ;
        RECT 151.000 52.100 151.400 52.200 ;
        RECT 147.000 51.800 151.400 52.100 ;
        RECT 175.000 52.100 175.400 52.200 ;
        RECT 179.800 52.100 180.200 52.200 ;
        RECT 175.000 51.800 180.200 52.100 ;
        RECT 195.800 52.100 196.200 52.200 ;
        RECT 197.400 52.100 197.800 52.200 ;
        RECT 195.800 51.800 197.800 52.100 ;
        RECT 199.800 52.100 200.200 52.200 ;
        RECT 202.200 52.100 202.600 52.200 ;
        RECT 199.800 51.800 202.600 52.100 ;
        RECT 219.800 52.100 220.200 52.200 ;
        RECT 231.000 52.100 231.400 52.200 ;
        RECT 219.800 51.800 231.400 52.100 ;
        RECT 235.000 52.100 235.400 52.200 ;
        RECT 246.200 52.100 246.600 52.200 ;
        RECT 235.000 51.800 246.600 52.100 ;
        RECT 57.400 51.100 57.800 51.200 ;
        RECT 59.800 51.100 60.200 51.200 ;
        RECT 68.600 51.100 69.000 51.200 ;
        RECT 57.400 50.800 69.000 51.100 ;
        RECT 109.400 51.100 109.800 51.200 ;
        RECT 116.600 51.100 117.000 51.200 ;
        RECT 109.400 50.800 117.000 51.100 ;
        RECT 120.600 51.100 121.000 51.200 ;
        RECT 127.800 51.100 128.200 51.200 ;
        RECT 120.600 50.800 128.200 51.100 ;
        RECT 143.000 51.100 143.400 51.200 ;
        RECT 144.600 51.100 145.000 51.200 ;
        RECT 143.000 50.800 145.000 51.100 ;
        RECT 168.600 51.100 169.000 51.200 ;
        RECT 171.000 51.100 171.400 51.200 ;
        RECT 168.600 50.800 171.400 51.100 ;
        RECT 241.400 51.100 241.800 51.200 ;
        RECT 252.600 51.100 253.000 51.200 ;
        RECT 259.000 51.100 259.400 51.200 ;
        RECT 241.400 50.800 259.400 51.100 ;
        RECT 71.800 49.800 72.200 50.200 ;
        RECT 98.200 50.100 98.600 50.200 ;
        RECT 103.800 50.100 104.200 50.200 ;
        RECT 98.200 49.800 104.200 50.100 ;
        RECT 125.400 50.100 125.800 50.200 ;
        RECT 129.400 50.100 129.800 50.200 ;
        RECT 125.400 49.800 129.800 50.100 ;
        RECT 17.400 49.100 17.800 49.200 ;
        RECT 18.200 49.100 18.600 49.200 ;
        RECT 26.200 49.100 26.600 49.200 ;
        RECT 17.400 48.800 26.600 49.100 ;
        RECT 33.400 49.100 33.800 49.200 ;
        RECT 35.800 49.100 36.200 49.200 ;
        RECT 33.400 48.800 36.200 49.100 ;
        RECT 39.000 48.800 39.400 49.200 ;
        RECT 43.000 49.100 43.400 49.200 ;
        RECT 51.800 49.100 52.200 49.200 ;
        RECT 43.000 48.800 52.200 49.100 ;
        RECT 63.000 49.100 63.400 49.200 ;
        RECT 67.000 49.100 67.400 49.200 ;
        RECT 63.000 48.800 67.400 49.100 ;
        RECT 68.600 49.100 69.000 49.200 ;
        RECT 71.000 49.100 71.400 49.200 ;
        RECT 68.600 48.800 71.400 49.100 ;
        RECT 71.800 49.100 72.100 49.800 ;
        RECT 86.200 49.100 86.600 49.200 ;
        RECT 71.800 48.800 86.600 49.100 ;
        RECT 99.000 48.800 99.400 49.200 ;
        RECT 131.800 49.100 132.200 49.200 ;
        RECT 132.600 49.100 133.000 49.200 ;
        RECT 131.800 48.800 133.000 49.100 ;
        RECT 139.800 49.100 140.200 49.200 ;
        RECT 146.200 49.100 146.600 49.200 ;
        RECT 139.800 48.800 146.600 49.100 ;
        RECT 151.800 49.100 152.200 49.200 ;
        RECT 158.200 49.100 158.600 49.200 ;
        RECT 151.800 48.800 158.600 49.100 ;
        RECT 206.200 49.100 206.600 49.200 ;
        RECT 217.400 49.100 217.800 49.200 ;
        RECT 206.200 48.800 217.800 49.100 ;
        RECT 223.800 49.100 224.200 49.200 ;
        RECT 235.000 49.100 235.400 49.200 ;
        RECT 242.200 49.100 242.600 49.200 ;
        RECT 246.200 49.100 246.600 49.200 ;
        RECT 247.800 49.100 248.200 49.200 ;
        RECT 223.800 48.800 238.500 49.100 ;
        RECT 242.200 48.800 248.200 49.100 ;
        RECT 14.200 48.100 14.600 48.200 ;
        RECT 39.000 48.100 39.300 48.800 ;
        RECT 52.600 48.100 53.000 48.200 ;
        RECT 14.200 47.800 53.000 48.100 ;
        RECT 79.800 48.100 80.200 48.200 ;
        RECT 87.800 48.100 88.200 48.200 ;
        RECT 79.800 47.800 88.200 48.100 ;
        RECT 90.200 48.100 90.600 48.200 ;
        RECT 99.000 48.100 99.300 48.800 ;
        RECT 238.200 48.200 238.500 48.800 ;
        RECT 90.200 47.800 99.300 48.100 ;
        RECT 128.600 47.800 129.000 48.200 ;
        RECT 129.400 48.100 129.800 48.200 ;
        RECT 131.800 48.100 132.200 48.200 ;
        RECT 139.000 48.100 139.400 48.200 ;
        RECT 155.000 48.100 155.400 48.200 ;
        RECT 129.400 47.800 155.400 48.100 ;
        RECT 167.000 48.100 167.400 48.200 ;
        RECT 185.400 48.100 185.800 48.200 ;
        RECT 167.000 47.800 185.800 48.100 ;
        RECT 199.800 48.100 200.200 48.200 ;
        RECT 211.800 48.100 212.200 48.200 ;
        RECT 199.800 47.800 212.200 48.100 ;
        RECT 238.200 47.800 238.600 48.200 ;
        RECT 244.600 48.100 245.000 48.200 ;
        RECT 252.600 48.100 253.000 48.200 ;
        RECT 244.600 47.800 253.000 48.100 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 26.200 47.100 26.600 47.200 ;
        RECT 31.800 47.100 32.200 47.200 ;
        RECT 26.200 46.800 32.200 47.100 ;
        RECT 48.600 47.100 49.000 47.200 ;
        RECT 53.400 47.100 53.800 47.200 ;
        RECT 48.600 46.800 53.800 47.100 ;
        RECT 57.400 46.800 57.800 47.200 ;
        RECT 72.600 47.100 73.000 47.200 ;
        RECT 82.200 47.100 82.600 47.200 ;
        RECT 83.800 47.100 84.200 47.200 ;
        RECT 91.000 47.100 91.400 47.200 ;
        RECT 99.000 47.100 99.400 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 72.600 46.800 101.000 47.100 ;
        RECT 117.400 46.800 117.800 47.200 ;
        RECT 128.600 47.100 128.900 47.800 ;
        RECT 131.000 47.100 131.400 47.200 ;
        RECT 143.800 47.100 144.200 47.200 ;
        RECT 128.600 46.800 144.200 47.100 ;
        RECT 155.800 46.800 156.200 47.200 ;
        RECT 174.200 47.100 174.600 47.200 ;
        RECT 183.000 47.100 183.400 47.200 ;
        RECT 174.200 46.800 183.400 47.100 ;
        RECT 185.400 47.100 185.700 47.800 ;
        RECT 199.000 47.100 199.400 47.200 ;
        RECT 185.400 46.800 199.400 47.100 ;
        RECT 201.400 47.100 201.800 47.200 ;
        RECT 213.400 47.100 213.800 47.200 ;
        RECT 201.400 46.800 213.800 47.100 ;
        RECT 231.000 46.800 231.400 47.200 ;
        RECT 232.600 47.100 233.000 47.200 ;
        RECT 243.800 47.100 244.200 47.200 ;
        RECT 232.600 46.800 244.200 47.100 ;
        RECT 252.600 46.800 253.000 47.200 ;
        RECT 16.600 46.200 16.900 46.800 ;
        RECT 4.600 46.100 5.000 46.200 ;
        RECT 11.800 46.100 12.200 46.200 ;
        RECT 4.600 45.800 12.200 46.100 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 22.200 46.100 22.600 46.300 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 22.200 45.800 28.200 46.100 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 31.800 45.800 33.000 46.100 ;
        RECT 35.800 46.100 36.200 46.200 ;
        RECT 53.400 46.100 53.800 46.200 ;
        RECT 57.400 46.100 57.700 46.800 ;
        RECT 58.200 46.100 58.600 46.200 ;
        RECT 35.800 45.800 58.600 46.100 ;
        RECT 83.000 46.100 83.400 46.200 ;
        RECT 84.600 46.100 85.000 46.200 ;
        RECT 83.000 45.800 85.000 46.100 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 98.200 45.800 103.400 46.100 ;
        RECT 117.400 46.100 117.700 46.800 ;
        RECT 123.000 46.100 123.400 46.200 ;
        RECT 117.400 45.800 123.400 46.100 ;
        RECT 128.600 46.100 129.000 46.200 ;
        RECT 143.800 46.100 144.200 46.200 ;
        RECT 128.600 45.800 144.200 46.100 ;
        RECT 153.400 46.100 153.800 46.200 ;
        RECT 155.800 46.100 156.100 46.800 ;
        RECT 231.000 46.200 231.300 46.800 ;
        RECT 159.000 46.100 159.400 46.200 ;
        RECT 153.400 45.800 159.400 46.100 ;
        RECT 176.600 46.100 177.000 46.200 ;
        RECT 207.000 46.100 207.400 46.200 ;
        RECT 211.800 46.100 212.200 46.200 ;
        RECT 176.600 45.800 212.200 46.100 ;
        RECT 219.800 46.100 220.200 46.200 ;
        RECT 231.000 46.100 231.400 46.200 ;
        RECT 233.400 46.100 233.800 46.200 ;
        RECT 219.800 45.800 221.700 46.100 ;
        RECT 231.000 45.800 233.800 46.100 ;
        RECT 251.000 46.100 251.400 46.200 ;
        RECT 252.600 46.100 252.900 46.800 ;
        RECT 251.000 45.800 252.900 46.100 ;
        RECT 253.400 46.100 253.800 46.200 ;
        RECT 259.800 46.100 260.200 46.200 ;
        RECT 253.400 45.800 260.200 46.100 ;
        RECT 143.800 45.200 144.100 45.800 ;
        RECT 221.400 45.200 221.700 45.800 ;
        RECT 31.000 45.100 31.400 45.200 ;
        RECT 58.200 45.100 58.600 45.200 ;
        RECT 31.000 44.800 58.600 45.100 ;
        RECT 61.400 45.100 61.800 45.200 ;
        RECT 62.200 45.100 62.600 45.200 ;
        RECT 61.400 44.800 62.600 45.100 ;
        RECT 78.200 45.100 78.600 45.200 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 111.800 45.100 112.200 45.200 ;
        RECT 78.200 44.800 82.500 45.100 ;
        RECT 85.400 44.800 112.200 45.100 ;
        RECT 123.800 45.100 124.200 45.200 ;
        RECT 126.200 45.100 126.600 45.200 ;
        RECT 123.800 44.800 126.600 45.100 ;
        RECT 127.800 45.100 128.200 45.200 ;
        RECT 135.000 45.100 135.400 45.200 ;
        RECT 127.800 44.800 135.400 45.100 ;
        RECT 138.200 45.100 138.600 45.200 ;
        RECT 143.000 45.100 143.400 45.200 ;
        RECT 138.200 44.800 143.400 45.100 ;
        RECT 143.800 44.800 144.200 45.200 ;
        RECT 164.600 45.100 165.000 45.200 ;
        RECT 155.800 44.800 165.000 45.100 ;
        RECT 172.600 45.100 173.000 45.200 ;
        RECT 175.800 45.100 176.200 45.200 ;
        RECT 182.200 45.100 182.600 45.200 ;
        RECT 172.600 44.800 182.600 45.100 ;
        RECT 185.400 45.100 185.800 45.200 ;
        RECT 187.800 45.100 188.200 45.200 ;
        RECT 185.400 44.800 188.200 45.100 ;
        RECT 201.400 45.100 201.800 45.200 ;
        RECT 216.600 45.100 217.000 45.200 ;
        RECT 201.400 44.800 217.000 45.100 ;
        RECT 221.400 44.800 221.800 45.200 ;
        RECT 237.400 45.100 237.800 45.200 ;
        RECT 254.200 45.100 254.600 45.200 ;
        RECT 260.600 45.100 261.000 45.200 ;
        RECT 237.400 44.800 261.000 45.100 ;
        RECT 82.200 44.200 82.500 44.800 ;
        RECT 155.800 44.200 156.100 44.800 ;
        RECT 82.200 43.800 82.600 44.200 ;
        RECT 92.600 44.100 93.000 44.200 ;
        RECT 110.200 44.100 110.600 44.200 ;
        RECT 111.800 44.100 112.200 44.200 ;
        RECT 92.600 43.800 112.200 44.100 ;
        RECT 124.600 44.100 125.000 44.200 ;
        RECT 131.800 44.100 132.200 44.200 ;
        RECT 133.400 44.100 133.800 44.200 ;
        RECT 143.000 44.100 143.400 44.200 ;
        RECT 124.600 43.800 143.400 44.100 ;
        RECT 155.800 43.800 156.200 44.200 ;
        RECT 196.600 44.100 197.000 44.200 ;
        RECT 204.600 44.100 205.000 44.200 ;
        RECT 196.600 43.800 205.000 44.100 ;
        RECT 218.200 44.100 218.600 44.200 ;
        RECT 226.200 44.100 226.600 44.200 ;
        RECT 218.200 43.800 226.600 44.100 ;
        RECT 230.200 44.100 230.600 44.200 ;
        RECT 241.400 44.100 241.800 44.200 ;
        RECT 243.000 44.100 243.400 44.200 ;
        RECT 230.200 43.800 243.400 44.100 ;
        RECT 260.600 44.100 261.000 44.200 ;
        RECT 264.600 44.100 265.000 44.200 ;
        RECT 260.600 43.800 265.000 44.100 ;
        RECT 92.600 43.100 93.000 43.200 ;
        RECT 108.600 43.100 109.000 43.200 ;
        RECT 92.600 42.800 109.000 43.100 ;
        RECT 132.600 43.100 133.000 43.200 ;
        RECT 143.000 43.100 143.400 43.200 ;
        RECT 156.600 43.100 157.000 43.200 ;
        RECT 159.800 43.100 160.200 43.200 ;
        RECT 165.400 43.100 165.800 43.200 ;
        RECT 171.800 43.100 172.200 43.200 ;
        RECT 132.600 42.800 140.100 43.100 ;
        RECT 143.000 42.800 172.200 43.100 ;
        RECT 228.600 43.100 229.000 43.200 ;
        RECT 250.200 43.100 250.600 43.200 ;
        RECT 228.600 42.800 250.600 43.100 ;
        RECT 139.800 42.200 140.100 42.800 ;
        RECT 38.200 42.100 38.600 42.200 ;
        RECT 95.800 42.100 96.200 42.200 ;
        RECT 38.200 41.800 96.200 42.100 ;
        RECT 123.000 42.100 123.400 42.200 ;
        RECT 126.200 42.100 126.600 42.200 ;
        RECT 123.000 41.800 126.600 42.100 ;
        RECT 135.800 42.100 136.200 42.200 ;
        RECT 137.400 42.100 137.800 42.200 ;
        RECT 135.800 41.800 137.800 42.100 ;
        RECT 139.800 41.800 140.200 42.200 ;
        RECT 145.400 42.100 145.800 42.200 ;
        RECT 180.600 42.100 181.000 42.200 ;
        RECT 145.400 41.800 181.000 42.100 ;
        RECT 182.200 42.100 182.600 42.200 ;
        RECT 204.600 42.100 205.000 42.200 ;
        RECT 182.200 41.800 205.000 42.100 ;
        RECT 225.400 42.100 225.800 42.200 ;
        RECT 243.800 42.100 244.200 42.200 ;
        RECT 247.800 42.100 248.200 42.200 ;
        RECT 225.400 41.800 248.200 42.100 ;
        RECT 83.800 41.100 84.200 41.200 ;
        RECT 103.800 41.100 104.200 41.200 ;
        RECT 83.800 40.800 104.200 41.100 ;
        RECT 203.800 41.100 204.200 41.200 ;
        RECT 212.600 41.100 213.000 41.200 ;
        RECT 203.800 40.800 213.000 41.100 ;
        RECT 86.200 40.100 86.600 40.200 ;
        RECT 115.800 40.100 116.200 40.200 ;
        RECT 86.200 39.800 116.200 40.100 ;
        RECT 144.600 40.100 145.000 40.200 ;
        RECT 153.400 40.100 153.800 40.200 ;
        RECT 144.600 39.800 153.800 40.100 ;
        RECT 170.200 40.100 170.600 40.200 ;
        RECT 206.200 40.100 206.600 40.200 ;
        RECT 170.200 39.800 206.600 40.100 ;
        RECT 217.400 40.100 217.800 40.200 ;
        RECT 247.000 40.100 247.400 40.200 ;
        RECT 249.400 40.100 249.800 40.200 ;
        RECT 259.800 40.100 260.200 40.200 ;
        RECT 217.400 39.800 260.200 40.100 ;
        RECT 0.600 39.100 1.000 39.200 ;
        RECT 13.400 39.100 13.800 39.200 ;
        RECT 15.000 39.100 15.400 39.200 ;
        RECT 122.200 39.100 122.600 39.200 ;
        RECT 0.600 38.800 15.400 39.100 ;
        RECT 66.200 38.800 122.600 39.100 ;
        RECT 123.000 39.100 123.400 39.200 ;
        RECT 145.400 39.100 145.800 39.200 ;
        RECT 123.000 38.800 145.800 39.100 ;
        RECT 151.000 39.100 151.400 39.200 ;
        RECT 151.800 39.100 152.200 39.200 ;
        RECT 151.000 38.800 152.200 39.100 ;
        RECT 154.200 39.100 154.600 39.200 ;
        RECT 156.600 39.100 157.000 39.200 ;
        RECT 154.200 38.800 157.000 39.100 ;
        RECT 167.800 39.100 168.200 39.200 ;
        RECT 172.600 39.100 173.000 39.200 ;
        RECT 211.800 39.100 212.200 39.200 ;
        RECT 167.800 38.800 212.200 39.100 ;
        RECT 66.200 38.200 66.500 38.800 ;
        RECT 66.200 37.800 66.600 38.200 ;
        RECT 69.400 38.100 69.800 38.200 ;
        RECT 71.800 38.100 72.200 38.200 ;
        RECT 84.600 38.100 85.000 38.200 ;
        RECT 88.600 38.100 89.000 38.200 ;
        RECT 69.400 37.800 89.000 38.100 ;
        RECT 89.400 38.100 89.800 38.200 ;
        RECT 119.000 38.100 119.400 38.200 ;
        RECT 89.400 37.800 119.400 38.100 ;
        RECT 143.800 38.100 144.200 38.200 ;
        RECT 154.200 38.100 154.600 38.200 ;
        RECT 143.800 37.800 154.600 38.100 ;
        RECT 155.800 38.100 156.200 38.200 ;
        RECT 167.800 38.100 168.200 38.200 ;
        RECT 155.800 37.800 168.200 38.100 ;
        RECT 168.600 38.100 169.000 38.200 ;
        RECT 170.200 38.100 170.600 38.200 ;
        RECT 168.600 37.800 170.600 38.100 ;
        RECT 187.000 38.100 187.400 38.200 ;
        RECT 215.000 38.100 215.400 38.200 ;
        RECT 187.000 37.800 215.400 38.100 ;
        RECT 1.400 37.100 1.800 37.200 ;
        RECT 3.800 37.100 4.200 37.200 ;
        RECT 12.600 37.100 13.000 37.200 ;
        RECT 1.400 36.800 13.000 37.100 ;
        RECT 73.400 37.100 73.800 37.200 ;
        RECT 82.200 37.100 82.600 37.200 ;
        RECT 87.000 37.100 87.400 37.200 ;
        RECT 73.400 36.800 87.400 37.100 ;
        RECT 110.200 37.100 110.600 37.200 ;
        RECT 111.000 37.100 111.400 37.200 ;
        RECT 110.200 36.800 111.400 37.100 ;
        RECT 118.200 37.100 118.600 37.200 ;
        RECT 191.000 37.100 191.400 37.200 ;
        RECT 118.200 36.800 191.400 37.100 ;
        RECT 226.200 36.800 226.600 37.200 ;
        RECT 232.600 36.800 233.000 37.200 ;
        RECT 235.800 37.100 236.200 37.200 ;
        RECT 241.400 37.100 241.800 37.200 ;
        RECT 235.000 36.800 241.800 37.100 ;
        RECT 226.200 36.200 226.500 36.800 ;
        RECT 232.600 36.200 232.900 36.800 ;
        RECT 11.800 35.800 12.200 36.200 ;
        RECT 27.800 36.100 28.200 36.200 ;
        RECT 29.400 36.100 29.800 36.200 ;
        RECT 39.000 36.100 39.400 36.200 ;
        RECT 27.800 35.800 39.400 36.100 ;
        RECT 62.200 36.100 62.600 36.200 ;
        RECT 63.800 36.100 64.200 36.200 ;
        RECT 67.000 36.100 67.400 36.200 ;
        RECT 62.200 35.800 67.400 36.100 ;
        RECT 76.600 35.800 77.000 36.200 ;
        RECT 79.800 36.100 80.200 36.200 ;
        RECT 80.600 36.100 81.000 36.200 ;
        RECT 79.800 35.800 81.000 36.100 ;
        RECT 95.800 36.100 96.200 36.200 ;
        RECT 104.600 36.100 105.000 36.200 ;
        RECT 117.400 36.100 117.800 36.200 ;
        RECT 174.200 36.100 174.600 36.200 ;
        RECT 176.600 36.100 177.000 36.200 ;
        RECT 95.800 35.800 117.800 36.100 ;
        RECT 142.200 35.800 177.000 36.100 ;
        RECT 180.600 36.100 181.000 36.200 ;
        RECT 183.800 36.100 184.200 36.200 ;
        RECT 187.800 36.100 188.200 36.200 ;
        RECT 180.600 35.800 188.200 36.100 ;
        RECT 203.000 35.800 203.400 36.200 ;
        RECT 204.600 36.100 205.000 36.200 ;
        RECT 207.000 36.100 207.400 36.200 ;
        RECT 204.600 35.800 207.400 36.100 ;
        RECT 219.800 35.800 220.200 36.200 ;
        RECT 226.200 35.800 226.600 36.200 ;
        RECT 232.600 36.100 233.000 36.200 ;
        RECT 235.000 36.100 235.400 36.200 ;
        RECT 232.600 35.800 235.400 36.100 ;
        RECT 11.800 35.100 12.100 35.800 ;
        RECT 22.200 35.100 22.600 35.200 ;
        RECT 11.800 34.800 22.600 35.100 ;
        RECT 34.200 35.100 34.600 35.200 ;
        RECT 35.800 35.100 36.200 35.200 ;
        RECT 34.200 34.800 36.200 35.100 ;
        RECT 37.400 35.100 37.800 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 37.400 34.800 41.000 35.100 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 61.400 35.100 61.800 35.200 ;
        RECT 60.600 34.800 61.800 35.100 ;
        RECT 63.000 35.100 63.400 35.200 ;
        RECT 63.800 35.100 64.200 35.200 ;
        RECT 63.000 34.800 64.200 35.100 ;
        RECT 71.800 35.100 72.200 35.200 ;
        RECT 76.600 35.100 76.900 35.800 ;
        RECT 71.800 34.800 76.900 35.100 ;
        RECT 79.800 35.100 80.100 35.800 ;
        RECT 142.200 35.200 142.500 35.800 ;
        RECT 89.400 35.100 89.800 35.200 ;
        RECT 79.800 34.800 89.800 35.100 ;
        RECT 101.400 35.100 101.800 35.200 ;
        RECT 102.200 35.100 102.600 35.200 ;
        RECT 101.400 34.800 102.600 35.100 ;
        RECT 106.200 35.100 106.600 35.200 ;
        RECT 125.400 35.100 125.800 35.200 ;
        RECT 106.200 34.800 125.800 35.100 ;
        RECT 139.800 35.100 140.200 35.200 ;
        RECT 140.600 35.100 141.000 35.200 ;
        RECT 142.200 35.100 142.600 35.200 ;
        RECT 139.800 34.800 142.600 35.100 ;
        RECT 144.600 34.800 145.000 35.200 ;
        RECT 166.200 35.100 166.600 35.200 ;
        RECT 167.000 35.100 167.400 35.200 ;
        RECT 166.200 34.800 167.400 35.100 ;
        RECT 182.200 35.100 182.600 35.200 ;
        RECT 188.600 35.100 189.000 35.200 ;
        RECT 182.200 34.800 189.000 35.100 ;
        RECT 189.400 35.100 189.800 35.200 ;
        RECT 196.600 35.100 197.000 35.200 ;
        RECT 189.400 34.800 197.000 35.100 ;
        RECT 202.200 35.100 202.600 35.200 ;
        RECT 203.000 35.100 203.300 35.800 ;
        RECT 219.800 35.100 220.100 35.800 ;
        RECT 202.200 34.800 220.100 35.100 ;
        RECT 231.000 35.100 231.400 35.200 ;
        RECT 236.600 35.100 237.000 35.200 ;
        RECT 231.000 34.800 237.000 35.100 ;
        RECT 249.400 35.100 249.800 35.200 ;
        RECT 256.600 35.100 257.000 35.200 ;
        RECT 249.400 34.800 257.000 35.100 ;
        RECT 259.800 35.100 260.200 35.200 ;
        RECT 263.000 35.100 263.400 35.200 ;
        RECT 259.800 34.800 263.400 35.100 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 23.000 34.100 23.400 34.200 ;
        RECT 38.200 34.100 38.600 34.200 ;
        RECT 17.400 33.800 38.600 34.100 ;
        RECT 61.400 34.100 61.800 34.200 ;
        RECT 63.800 34.100 64.200 34.200 ;
        RECT 61.400 33.800 64.200 34.100 ;
        RECT 69.400 34.100 69.800 34.200 ;
        RECT 81.400 34.100 81.800 34.200 ;
        RECT 69.400 33.800 81.800 34.100 ;
        RECT 83.800 34.100 84.200 34.200 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 83.800 33.800 89.000 34.100 ;
        RECT 91.800 34.100 92.200 34.200 ;
        RECT 92.600 34.100 93.000 34.200 ;
        RECT 91.800 33.800 93.000 34.100 ;
        RECT 97.400 34.100 97.800 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 97.400 33.800 105.000 34.100 ;
        RECT 117.400 34.100 117.800 34.200 ;
        RECT 123.800 34.100 124.200 34.200 ;
        RECT 133.400 34.100 133.800 34.200 ;
        RECT 144.600 34.100 144.900 34.800 ;
        RECT 117.400 33.800 144.900 34.100 ;
        RECT 154.200 34.100 154.600 34.200 ;
        RECT 175.000 34.100 175.400 34.200 ;
        RECT 154.200 33.800 175.400 34.100 ;
        RECT 175.800 33.800 176.200 34.200 ;
        RECT 177.400 34.100 177.800 34.200 ;
        RECT 188.600 34.100 189.000 34.200 ;
        RECT 177.400 33.800 189.000 34.100 ;
        RECT 189.400 34.100 189.800 34.200 ;
        RECT 190.200 34.100 190.600 34.200 ;
        RECT 189.400 33.800 190.600 34.100 ;
        RECT 195.000 34.100 195.400 34.200 ;
        RECT 201.400 34.100 201.800 34.200 ;
        RECT 195.000 33.800 201.800 34.100 ;
        RECT 207.000 34.100 207.400 34.200 ;
        RECT 222.200 34.100 222.600 34.200 ;
        RECT 225.400 34.100 225.800 34.200 ;
        RECT 207.000 33.800 225.800 34.100 ;
        RECT 4.600 33.100 5.000 33.200 ;
        RECT 7.000 33.100 7.400 33.200 ;
        RECT 9.400 33.100 9.800 33.200 ;
        RECT 4.600 32.800 9.800 33.100 ;
        RECT 11.000 33.100 11.400 33.200 ;
        RECT 12.600 33.100 13.000 33.200 ;
        RECT 11.000 32.800 13.000 33.100 ;
        RECT 19.000 33.100 19.400 33.200 ;
        RECT 22.200 33.100 22.600 33.200 ;
        RECT 19.000 32.800 22.600 33.100 ;
        RECT 27.000 33.100 27.400 33.200 ;
        RECT 32.600 33.100 33.000 33.200 ;
        RECT 27.000 32.800 33.000 33.100 ;
        RECT 59.800 33.100 60.200 33.200 ;
        RECT 61.400 33.100 61.800 33.200 ;
        RECT 59.800 32.800 61.800 33.100 ;
        RECT 103.000 33.100 103.400 33.200 ;
        RECT 134.200 33.100 134.600 33.200 ;
        RECT 103.000 32.800 134.600 33.100 ;
        RECT 153.400 33.100 153.800 33.200 ;
        RECT 160.600 33.100 161.000 33.200 ;
        RECT 153.400 32.800 161.000 33.100 ;
        RECT 161.400 33.100 161.800 33.200 ;
        RECT 175.800 33.100 176.100 33.800 ;
        RECT 161.400 32.800 176.100 33.100 ;
        RECT 187.000 33.100 187.400 33.200 ;
        RECT 193.400 33.100 193.800 33.200 ;
        RECT 199.000 33.100 199.400 33.200 ;
        RECT 187.000 32.800 199.400 33.100 ;
        RECT 202.200 33.100 202.600 33.200 ;
        RECT 207.000 33.100 207.400 33.200 ;
        RECT 202.200 32.800 207.400 33.100 ;
        RECT 210.200 33.100 210.600 33.200 ;
        RECT 215.800 33.100 216.200 33.200 ;
        RECT 210.200 32.800 216.200 33.100 ;
        RECT 219.000 33.100 219.400 33.200 ;
        RECT 255.000 33.100 255.400 33.200 ;
        RECT 219.000 32.800 255.400 33.100 ;
        RECT 25.400 32.100 25.800 32.200 ;
        RECT 31.000 32.100 31.400 32.200 ;
        RECT 34.200 32.100 34.600 32.200 ;
        RECT 25.400 31.800 34.600 32.100 ;
        RECT 44.600 32.100 45.000 32.200 ;
        RECT 53.400 32.100 53.800 32.200 ;
        RECT 44.600 31.800 53.800 32.100 ;
        RECT 58.200 32.100 58.600 32.200 ;
        RECT 64.600 32.100 65.000 32.200 ;
        RECT 58.200 31.800 65.000 32.100 ;
        RECT 70.200 32.100 70.600 32.200 ;
        RECT 124.600 32.100 125.000 32.200 ;
        RECT 70.200 31.800 125.000 32.100 ;
        RECT 159.000 32.100 159.400 32.200 ;
        RECT 179.000 32.100 179.400 32.200 ;
        RECT 159.000 31.800 179.400 32.100 ;
        RECT 214.200 32.100 214.600 32.200 ;
        RECT 232.600 32.100 233.000 32.200 ;
        RECT 214.200 31.800 233.000 32.100 ;
        RECT 26.200 31.100 26.600 31.200 ;
        RECT 63.000 31.100 63.400 31.200 ;
        RECT 26.200 30.800 63.400 31.100 ;
        RECT 91.800 31.100 92.200 31.200 ;
        RECT 95.000 31.100 95.400 31.200 ;
        RECT 91.800 30.800 95.400 31.100 ;
        RECT 130.200 31.100 130.600 31.200 ;
        RECT 170.200 31.100 170.600 31.200 ;
        RECT 130.200 30.800 170.600 31.100 ;
        RECT 184.600 31.100 185.000 31.200 ;
        RECT 191.000 31.100 191.400 31.200 ;
        RECT 201.400 31.100 201.800 31.200 ;
        RECT 203.800 31.100 204.200 31.200 ;
        RECT 184.600 30.800 204.200 31.100 ;
        RECT 219.000 30.800 219.400 31.200 ;
        RECT 235.800 31.100 236.200 31.200 ;
        RECT 246.200 31.100 246.600 31.200 ;
        RECT 247.800 31.100 248.200 31.200 ;
        RECT 261.400 31.100 261.800 31.200 ;
        RECT 235.800 30.800 261.800 31.100 ;
        RECT 219.000 30.200 219.300 30.800 ;
        RECT 35.800 30.100 36.200 30.200 ;
        RECT 39.000 30.100 39.400 30.200 ;
        RECT 35.800 29.800 39.400 30.100 ;
        RECT 41.400 30.100 41.800 30.200 ;
        RECT 45.400 30.100 45.800 30.200 ;
        RECT 41.400 29.800 45.800 30.100 ;
        RECT 141.400 30.100 141.800 30.200 ;
        RECT 144.600 30.100 145.000 30.200 ;
        RECT 141.400 29.800 145.000 30.100 ;
        RECT 219.000 29.800 219.400 30.200 ;
        RECT 222.200 30.100 222.600 30.200 ;
        RECT 226.200 30.100 226.600 30.200 ;
        RECT 222.200 29.800 226.600 30.100 ;
        RECT 237.400 30.100 237.800 30.200 ;
        RECT 248.600 30.100 249.000 30.200 ;
        RECT 237.400 29.800 249.000 30.100 ;
        RECT 20.600 29.100 21.000 29.200 ;
        RECT 27.800 29.100 28.200 29.200 ;
        RECT 20.600 28.800 28.200 29.100 ;
        RECT 31.800 29.100 32.200 29.200 ;
        RECT 35.800 29.100 36.100 29.800 ;
        RECT 31.800 28.800 36.100 29.100 ;
        RECT 37.400 29.100 37.800 29.200 ;
        RECT 42.200 29.100 42.600 29.200 ;
        RECT 37.400 28.800 42.600 29.100 ;
        RECT 43.800 29.100 44.200 29.200 ;
        RECT 46.200 29.100 46.600 29.200 ;
        RECT 43.800 28.800 46.600 29.100 ;
        RECT 73.400 29.100 73.800 29.200 ;
        RECT 97.400 29.100 97.800 29.200 ;
        RECT 114.200 29.100 114.600 29.200 ;
        RECT 73.400 28.800 87.300 29.100 ;
        RECT 97.400 28.800 114.600 29.100 ;
        RECT 155.000 29.100 155.400 29.200 ;
        RECT 163.800 29.100 164.200 29.200 ;
        RECT 172.600 29.100 173.000 29.200 ;
        RECT 182.200 29.100 182.600 29.200 ;
        RECT 184.600 29.100 185.000 29.200 ;
        RECT 155.000 28.800 173.000 29.100 ;
        RECT 181.400 28.800 185.000 29.100 ;
        RECT 191.000 29.100 191.400 29.200 ;
        RECT 195.000 29.100 195.400 29.200 ;
        RECT 191.000 28.800 195.400 29.100 ;
        RECT 195.800 29.100 196.200 29.200 ;
        RECT 203.000 29.100 203.400 29.200 ;
        RECT 195.800 28.800 203.400 29.100 ;
        RECT 205.400 29.100 205.800 29.200 ;
        RECT 210.200 29.100 210.600 29.200 ;
        RECT 205.400 28.800 210.600 29.100 ;
        RECT 220.600 29.100 221.000 29.200 ;
        RECT 221.400 29.100 221.800 29.200 ;
        RECT 220.600 28.800 221.800 29.100 ;
        RECT 223.000 29.100 223.400 29.200 ;
        RECT 223.800 29.100 224.200 29.200 ;
        RECT 223.000 28.800 224.200 29.100 ;
        RECT 227.000 29.100 227.400 29.200 ;
        RECT 234.200 29.100 234.600 29.200 ;
        RECT 243.000 29.100 243.400 29.200 ;
        RECT 227.000 28.800 243.400 29.100 ;
        RECT 87.000 28.200 87.300 28.800 ;
        RECT 29.400 27.800 29.800 28.200 ;
        RECT 32.600 28.100 33.000 28.200 ;
        RECT 47.800 28.100 48.200 28.200 ;
        RECT 32.600 27.800 48.200 28.100 ;
        RECT 48.600 27.800 49.000 28.200 ;
        RECT 79.000 28.100 79.400 28.200 ;
        RECT 85.400 28.100 85.800 28.200 ;
        RECT 86.200 28.100 86.600 28.200 ;
        RECT 79.000 27.800 84.100 28.100 ;
        RECT 85.400 27.800 86.600 28.100 ;
        RECT 87.000 28.100 87.400 28.200 ;
        RECT 94.200 28.100 94.600 28.200 ;
        RECT 87.000 27.800 94.600 28.100 ;
        RECT 116.600 28.100 117.000 28.200 ;
        RECT 156.600 28.100 157.000 28.200 ;
        RECT 116.600 27.800 157.000 28.100 ;
        RECT 160.600 28.100 161.000 28.200 ;
        RECT 205.400 28.100 205.800 28.200 ;
        RECT 160.600 27.800 205.800 28.100 ;
        RECT 213.400 28.100 213.800 28.200 ;
        RECT 239.800 28.100 240.200 28.200 ;
        RECT 213.400 27.800 240.200 28.100 ;
        RECT 253.400 28.100 253.800 28.200 ;
        RECT 263.800 28.100 264.200 28.200 ;
        RECT 253.400 27.800 264.200 28.100 ;
        RECT 6.200 26.800 6.600 27.200 ;
        RECT 29.400 27.100 29.700 27.800 ;
        RECT 16.600 26.800 29.700 27.100 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 42.200 27.100 42.600 27.200 ;
        RECT 48.600 27.100 48.900 27.800 ;
        RECT 54.200 27.100 54.600 27.200 ;
        RECT 42.200 26.800 54.600 27.100 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 66.200 27.100 66.600 27.200 ;
        RECT 61.400 26.800 66.600 27.100 ;
        RECT 71.800 27.100 72.200 27.200 ;
        RECT 83.000 27.100 83.400 27.200 ;
        RECT 71.800 26.800 83.400 27.100 ;
        RECT 83.800 27.100 84.100 27.800 ;
        RECT 89.400 27.100 89.800 27.200 ;
        RECT 83.800 26.800 89.800 27.100 ;
        RECT 117.400 27.100 117.800 27.200 ;
        RECT 118.200 27.100 118.600 27.200 ;
        RECT 117.400 26.800 118.600 27.100 ;
        RECT 142.200 26.800 142.600 27.200 ;
        RECT 149.400 26.800 149.800 27.200 ;
        RECT 167.800 27.100 168.200 27.200 ;
        RECT 200.600 27.100 201.000 27.200 ;
        RECT 167.800 26.800 201.000 27.100 ;
        RECT 201.400 27.100 201.800 27.200 ;
        RECT 203.000 27.100 203.400 27.200 ;
        RECT 201.400 26.800 203.400 27.100 ;
        RECT 207.800 27.100 208.200 27.200 ;
        RECT 218.200 27.100 218.600 27.200 ;
        RECT 207.800 26.800 218.600 27.100 ;
        RECT 238.200 27.100 238.600 27.200 ;
        RECT 239.000 27.100 239.400 27.200 ;
        RECT 238.200 26.800 239.400 27.100 ;
        RECT 239.800 26.800 240.200 27.200 ;
        RECT 6.200 26.100 6.500 26.800 ;
        RECT 16.600 26.200 16.900 26.800 ;
        RECT 10.200 26.100 10.600 26.200 ;
        RECT 6.200 25.800 10.600 26.100 ;
        RECT 12.600 26.100 13.000 26.200 ;
        RECT 16.600 26.100 17.000 26.200 ;
        RECT 12.600 25.800 17.000 26.100 ;
        RECT 21.400 26.100 21.800 26.200 ;
        RECT 24.600 26.100 25.000 26.200 ;
        RECT 21.400 25.800 25.000 26.100 ;
        RECT 35.000 26.100 35.400 26.200 ;
        RECT 39.000 26.100 39.300 26.800 ;
        RECT 35.000 25.800 39.300 26.100 ;
        RECT 47.800 26.100 48.200 26.200 ;
        RECT 60.600 26.100 61.000 26.200 ;
        RECT 47.800 25.800 61.000 26.100 ;
        RECT 73.400 26.100 73.800 26.200 ;
        RECT 104.600 26.100 105.000 26.200 ;
        RECT 113.400 26.100 113.800 26.200 ;
        RECT 73.400 25.800 93.700 26.100 ;
        RECT 104.600 25.800 113.800 26.100 ;
        RECT 116.600 26.100 117.000 26.200 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 134.200 26.100 134.600 26.200 ;
        RECT 116.600 25.800 119.300 26.100 ;
        RECT 127.000 25.800 134.600 26.100 ;
        RECT 137.400 26.100 137.800 26.200 ;
        RECT 142.200 26.100 142.500 26.800 ;
        RECT 137.400 25.800 142.500 26.100 ;
        RECT 147.000 26.100 147.400 26.200 ;
        RECT 149.400 26.100 149.700 26.800 ;
        RECT 151.800 26.100 152.200 26.200 ;
        RECT 165.400 26.100 165.800 26.200 ;
        RECT 168.600 26.100 169.000 26.200 ;
        RECT 147.000 25.800 169.000 26.100 ;
        RECT 175.000 26.100 175.400 26.200 ;
        RECT 203.800 26.100 204.200 26.200 ;
        RECT 175.000 25.800 204.200 26.100 ;
        RECT 207.000 26.100 207.400 26.200 ;
        RECT 216.600 26.100 217.000 26.200 ;
        RECT 207.000 25.800 217.000 26.100 ;
        RECT 239.800 26.100 240.100 26.800 ;
        RECT 244.600 26.100 245.000 26.200 ;
        RECT 239.800 25.800 245.000 26.100 ;
        RECT 250.200 26.100 250.600 26.200 ;
        RECT 251.000 26.100 251.400 26.200 ;
        RECT 250.200 25.800 251.400 26.100 ;
        RECT 93.400 25.200 93.700 25.800 ;
        RECT 119.000 25.200 119.300 25.800 ;
        RECT 47.800 25.100 48.200 25.200 ;
        RECT 50.200 25.100 50.600 25.200 ;
        RECT 47.800 24.800 50.600 25.100 ;
        RECT 52.600 25.100 53.000 25.200 ;
        RECT 67.800 25.100 68.200 25.200 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 52.600 24.800 61.700 25.100 ;
        RECT 67.800 24.800 69.800 25.100 ;
        RECT 83.800 25.100 84.200 25.200 ;
        RECT 84.600 25.100 85.000 25.200 ;
        RECT 83.800 24.800 85.000 25.100 ;
        RECT 93.400 24.800 93.800 25.200 ;
        RECT 102.200 25.100 102.600 25.200 ;
        RECT 103.800 25.100 104.200 25.200 ;
        RECT 102.200 24.800 104.200 25.100 ;
        RECT 119.000 24.800 119.400 25.200 ;
        RECT 151.000 25.100 151.400 25.200 ;
        RECT 158.200 25.100 158.600 25.200 ;
        RECT 151.000 24.800 158.600 25.100 ;
        RECT 166.200 24.800 166.600 25.200 ;
        RECT 168.600 25.100 169.000 25.200 ;
        RECT 243.800 25.100 244.200 25.200 ;
        RECT 247.000 25.100 247.400 25.200 ;
        RECT 168.600 24.800 247.400 25.100 ;
        RECT 61.400 24.200 61.700 24.800 ;
        RECT 61.400 23.800 61.800 24.200 ;
        RECT 104.600 24.100 105.000 24.200 ;
        RECT 109.400 24.100 109.800 24.200 ;
        RECT 123.800 24.100 124.200 24.200 ;
        RECT 104.600 23.800 124.200 24.100 ;
        RECT 124.600 24.100 125.000 24.200 ;
        RECT 139.000 24.100 139.400 24.200 ;
        RECT 159.000 24.100 159.400 24.200 ;
        RECT 124.600 23.800 159.400 24.100 ;
        RECT 166.200 24.100 166.500 24.800 ;
        RECT 175.800 24.100 176.200 24.200 ;
        RECT 166.200 23.800 176.200 24.100 ;
        RECT 196.600 24.100 197.000 24.200 ;
        RECT 256.600 24.100 257.000 24.200 ;
        RECT 196.600 23.800 257.000 24.100 ;
        RECT 25.400 23.100 25.800 23.200 ;
        RECT 42.200 23.100 42.600 23.200 ;
        RECT 50.200 23.100 50.600 23.200 ;
        RECT 25.400 22.800 50.600 23.100 ;
        RECT 88.600 23.100 89.000 23.200 ;
        RECT 175.000 23.100 175.400 23.200 ;
        RECT 88.600 22.800 175.400 23.100 ;
        RECT 67.000 22.100 67.400 22.200 ;
        RECT 75.000 22.100 75.400 22.200 ;
        RECT 67.000 21.800 75.400 22.100 ;
        RECT 171.800 22.100 172.200 22.200 ;
        RECT 181.400 22.100 181.800 22.200 ;
        RECT 171.800 21.800 181.800 22.100 ;
        RECT 183.000 22.100 183.400 22.200 ;
        RECT 222.200 22.100 222.600 22.200 ;
        RECT 183.000 21.800 222.600 22.100 ;
        RECT 63.800 21.100 64.200 21.200 ;
        RECT 106.200 21.100 106.600 21.200 ;
        RECT 63.800 20.800 106.600 21.100 ;
        RECT 108.600 21.100 109.000 21.200 ;
        RECT 119.800 21.100 120.200 21.200 ;
        RECT 108.600 20.800 120.200 21.100 ;
        RECT 193.400 21.100 193.800 21.200 ;
        RECT 227.800 21.100 228.200 21.200 ;
        RECT 193.400 20.800 228.200 21.100 ;
        RECT 101.400 20.100 101.800 20.200 ;
        RECT 108.600 20.100 109.000 20.200 ;
        RECT 114.200 20.100 114.600 20.200 ;
        RECT 101.400 19.800 114.600 20.100 ;
        RECT 165.400 20.100 165.800 20.200 ;
        RECT 237.400 20.100 237.800 20.200 ;
        RECT 165.400 19.800 237.800 20.100 ;
        RECT 255.000 19.800 255.400 20.200 ;
        RECT 255.000 19.200 255.300 19.800 ;
        RECT 1.400 19.100 1.800 19.200 ;
        RECT 7.800 19.100 8.200 19.200 ;
        RECT 18.200 19.100 18.600 19.200 ;
        RECT 1.400 18.800 18.600 19.100 ;
        RECT 67.800 19.100 68.200 19.200 ;
        RECT 80.600 19.100 81.000 19.200 ;
        RECT 67.800 18.800 81.000 19.100 ;
        RECT 83.000 19.100 83.400 19.200 ;
        RECT 86.200 19.100 86.600 19.200 ;
        RECT 83.000 18.800 86.600 19.100 ;
        RECT 96.600 19.100 97.000 19.200 ;
        RECT 97.400 19.100 97.800 19.200 ;
        RECT 96.600 18.800 97.800 19.100 ;
        RECT 106.200 19.100 106.600 19.200 ;
        RECT 130.200 19.100 130.600 19.200 ;
        RECT 106.200 18.800 130.600 19.100 ;
        RECT 186.200 19.100 186.600 19.200 ;
        RECT 195.800 19.100 196.200 19.200 ;
        RECT 186.200 18.800 196.200 19.100 ;
        RECT 254.200 18.800 254.600 19.200 ;
        RECT 255.000 18.800 255.400 19.200 ;
        RECT 254.200 18.200 254.500 18.800 ;
        RECT 41.400 18.100 41.800 18.200 ;
        RECT 52.600 18.100 53.000 18.200 ;
        RECT 57.400 18.100 57.800 18.200 ;
        RECT 100.600 18.100 101.000 18.200 ;
        RECT 41.400 17.800 101.000 18.100 ;
        RECT 118.200 18.100 118.600 18.200 ;
        RECT 132.600 18.100 133.000 18.200 ;
        RECT 118.200 17.800 133.000 18.100 ;
        RECT 159.000 18.100 159.400 18.200 ;
        RECT 159.800 18.100 160.200 18.200 ;
        RECT 159.000 17.800 160.200 18.100 ;
        RECT 250.200 18.100 250.600 18.200 ;
        RECT 251.800 18.100 252.200 18.200 ;
        RECT 250.200 17.800 252.200 18.100 ;
        RECT 254.200 17.800 254.600 18.200 ;
        RECT 19.000 17.100 19.400 17.200 ;
        RECT 19.800 17.100 20.200 17.200 ;
        RECT 19.000 16.800 20.200 17.100 ;
        RECT 63.000 17.100 63.400 17.200 ;
        RECT 73.400 17.100 73.800 17.200 ;
        RECT 74.200 17.100 74.600 17.200 ;
        RECT 63.000 16.800 74.600 17.100 ;
        RECT 85.400 17.100 85.800 17.200 ;
        RECT 87.800 17.100 88.200 17.200 ;
        RECT 93.400 17.100 93.800 17.200 ;
        RECT 85.400 16.800 93.800 17.100 ;
        RECT 100.600 17.100 101.000 17.200 ;
        RECT 183.000 17.100 183.400 17.200 ;
        RECT 100.600 16.800 183.400 17.100 ;
        RECT 208.600 17.100 209.000 17.200 ;
        RECT 211.800 17.100 212.200 17.200 ;
        RECT 208.600 16.800 212.200 17.100 ;
        RECT 227.000 17.100 227.400 17.200 ;
        RECT 232.600 17.100 233.000 17.200 ;
        RECT 227.000 16.800 233.000 17.100 ;
        RECT 251.800 16.800 252.200 17.200 ;
        RECT 8.600 16.100 9.000 16.200 ;
        RECT 11.000 16.100 11.400 16.200 ;
        RECT 8.600 15.800 11.400 16.100 ;
        RECT 11.800 15.800 12.200 16.200 ;
        RECT 14.200 16.100 14.600 16.200 ;
        RECT 17.400 16.100 17.800 16.200 ;
        RECT 62.200 16.100 62.600 16.200 ;
        RECT 14.200 15.800 62.600 16.100 ;
        RECT 73.400 15.800 73.800 16.200 ;
        RECT 83.800 15.800 84.200 16.200 ;
        RECT 91.800 16.100 92.200 16.200 ;
        RECT 92.600 16.100 93.000 16.200 ;
        RECT 91.000 15.800 93.000 16.100 ;
        RECT 93.400 16.100 93.800 16.200 ;
        RECT 94.200 16.100 94.600 16.200 ;
        RECT 93.400 15.800 94.600 16.100 ;
        RECT 123.000 16.100 123.400 16.200 ;
        RECT 125.400 16.100 125.800 16.200 ;
        RECT 165.400 16.100 165.800 16.200 ;
        RECT 123.000 15.800 165.800 16.100 ;
        RECT 175.000 16.100 175.400 16.200 ;
        RECT 176.600 16.100 177.000 16.200 ;
        RECT 175.000 15.800 177.000 16.100 ;
        RECT 183.800 15.800 184.200 16.200 ;
        RECT 187.000 15.800 187.400 16.200 ;
        RECT 211.800 16.100 212.200 16.200 ;
        RECT 218.200 16.100 218.600 16.200 ;
        RECT 211.000 15.800 218.600 16.100 ;
        RECT 228.600 15.800 229.000 16.200 ;
        RECT 251.800 16.100 252.100 16.800 ;
        RECT 252.600 16.100 253.000 16.200 ;
        RECT 251.800 15.800 253.000 16.100 ;
        RECT 11.800 15.200 12.100 15.800 ;
        RECT 73.400 15.200 73.700 15.800 ;
        RECT 10.200 15.100 10.600 15.200 ;
        RECT 7.000 14.800 10.600 15.100 ;
        RECT 11.800 15.100 12.200 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 61.400 15.100 61.800 15.200 ;
        RECT 62.200 15.100 62.600 15.200 ;
        RECT 11.800 14.800 62.600 15.100 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 83.800 15.100 84.100 15.800 ;
        RECT 183.800 15.200 184.100 15.800 ;
        RECT 95.800 15.100 96.200 15.200 ;
        RECT 83.800 14.800 96.200 15.100 ;
        RECT 99.000 15.100 99.400 15.200 ;
        RECT 99.800 15.100 100.200 15.200 ;
        RECT 99.000 14.800 100.200 15.100 ;
        RECT 111.000 15.100 111.400 15.200 ;
        RECT 128.600 15.100 129.000 15.200 ;
        RECT 111.000 14.800 129.000 15.100 ;
        RECT 134.200 15.100 134.600 15.200 ;
        RECT 148.600 15.100 149.000 15.200 ;
        RECT 152.600 15.100 153.000 15.200 ;
        RECT 160.600 15.100 161.000 15.200 ;
        RECT 171.000 15.100 171.400 15.200 ;
        RECT 174.200 15.100 174.600 15.200 ;
        RECT 134.200 14.800 174.600 15.100 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 7.000 14.200 7.300 14.800 ;
        RECT 7.000 13.800 7.400 14.200 ;
        RECT 18.200 14.100 18.600 14.200 ;
        RECT 19.000 14.100 19.400 14.200 ;
        RECT 19.800 14.100 20.200 14.200 ;
        RECT 18.200 13.800 20.200 14.100 ;
        RECT 23.800 14.100 24.200 14.200 ;
        RECT 33.400 14.100 33.800 14.200 ;
        RECT 23.800 13.800 33.800 14.100 ;
        RECT 35.000 14.100 35.400 14.200 ;
        RECT 37.400 14.100 37.800 14.200 ;
        RECT 35.000 13.800 37.800 14.100 ;
        RECT 39.800 13.800 40.200 14.200 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 60.600 14.100 61.000 14.200 ;
        RECT 66.200 14.100 66.600 14.200 ;
        RECT 59.000 13.800 61.000 14.100 ;
        RECT 61.400 13.800 66.600 14.100 ;
        RECT 95.000 14.100 95.400 14.200 ;
        RECT 108.600 14.100 109.000 14.200 ;
        RECT 111.800 14.100 112.200 14.200 ;
        RECT 95.000 13.800 112.200 14.100 ;
        RECT 140.600 14.100 141.000 14.200 ;
        RECT 144.600 14.100 145.000 14.200 ;
        RECT 156.600 14.100 157.000 14.200 ;
        RECT 164.600 14.100 165.000 14.200 ;
        RECT 166.200 14.100 166.600 14.200 ;
        RECT 140.600 13.800 148.900 14.100 ;
        RECT 156.600 13.800 166.600 14.100 ;
        RECT 176.600 14.100 177.000 14.200 ;
        RECT 187.000 14.100 187.300 15.800 ;
        RECT 188.600 15.100 189.000 15.200 ;
        RECT 196.600 15.100 197.000 15.200 ;
        RECT 210.200 15.100 210.600 15.200 ;
        RECT 213.400 15.100 213.800 15.200 ;
        RECT 220.600 15.100 221.000 15.200 ;
        RECT 228.600 15.100 228.900 15.800 ;
        RECT 188.600 14.800 228.900 15.100 ;
        RECT 231.000 15.100 231.400 15.200 ;
        RECT 237.400 15.100 237.800 15.200 ;
        RECT 231.000 14.800 237.800 15.100 ;
        RECT 251.000 15.100 251.400 15.200 ;
        RECT 259.800 15.100 260.200 15.200 ;
        RECT 251.000 14.800 260.200 15.100 ;
        RECT 176.600 13.800 187.300 14.100 ;
        RECT 199.800 14.100 200.200 14.200 ;
        RECT 211.000 14.100 211.400 14.200 ;
        RECT 199.800 13.800 211.400 14.100 ;
        RECT 224.600 14.100 225.000 14.200 ;
        RECT 247.800 14.100 248.200 14.200 ;
        RECT 248.600 14.100 249.000 14.200 ;
        RECT 224.600 13.800 249.000 14.100 ;
        RECT 12.600 13.100 13.000 13.200 ;
        RECT 7.000 12.800 13.000 13.100 ;
        RECT 13.400 13.100 13.800 13.200 ;
        RECT 39.800 13.100 40.100 13.800 ;
        RECT 13.400 12.800 40.100 13.100 ;
        RECT 61.400 13.200 61.700 13.800 ;
        RECT 148.600 13.200 148.900 13.800 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 148.600 12.800 149.000 13.200 ;
        RECT 151.000 13.100 151.400 13.200 ;
        RECT 161.400 13.100 161.800 13.200 ;
        RECT 151.000 12.800 161.800 13.100 ;
        RECT 179.000 13.100 179.400 13.200 ;
        RECT 194.200 13.100 194.600 13.200 ;
        RECT 179.000 12.800 194.600 13.100 ;
        RECT 7.000 12.200 7.300 12.800 ;
        RECT 7.000 11.800 7.400 12.200 ;
        RECT 30.200 12.100 30.600 12.200 ;
        RECT 37.400 12.100 37.800 12.200 ;
        RECT 30.200 11.800 37.800 12.100 ;
        RECT 50.200 12.100 50.600 12.200 ;
        RECT 97.400 12.100 97.800 12.200 ;
        RECT 50.200 11.800 97.800 12.100 ;
        RECT 98.200 12.100 98.600 12.200 ;
        RECT 107.800 12.100 108.200 12.200 ;
        RECT 98.200 11.800 108.200 12.100 ;
        RECT 113.400 12.100 113.800 12.200 ;
        RECT 123.000 12.100 123.400 12.200 ;
        RECT 113.400 11.800 123.400 12.100 ;
        RECT 179.800 12.100 180.200 12.200 ;
        RECT 192.600 12.100 193.000 12.200 ;
        RECT 179.800 11.800 193.000 12.100 ;
        RECT 206.200 12.100 206.600 12.200 ;
        RECT 219.000 12.100 219.400 12.200 ;
        RECT 206.200 11.800 219.400 12.100 ;
        RECT 65.400 11.100 65.800 11.200 ;
        RECT 93.400 11.100 93.800 11.200 ;
        RECT 65.400 10.800 93.800 11.100 ;
        RECT 76.600 10.100 77.000 10.200 ;
        RECT 81.400 10.100 81.800 10.200 ;
        RECT 91.000 10.100 91.400 10.200 ;
        RECT 76.600 9.800 91.400 10.100 ;
        RECT 122.200 10.100 122.600 10.200 ;
        RECT 129.400 10.100 129.800 10.200 ;
        RECT 135.000 10.100 135.400 10.200 ;
        RECT 122.200 9.800 135.400 10.100 ;
        RECT 220.600 10.100 221.000 10.200 ;
        RECT 225.400 10.100 225.800 10.200 ;
        RECT 229.400 10.100 229.800 10.200 ;
        RECT 220.600 9.800 229.800 10.100 ;
        RECT 230.200 10.100 230.600 10.200 ;
        RECT 237.400 10.100 237.800 10.200 ;
        RECT 247.800 10.100 248.200 10.200 ;
        RECT 230.200 9.800 248.200 10.100 ;
        RECT 20.600 9.100 21.000 9.200 ;
        RECT 29.400 9.100 29.800 9.200 ;
        RECT 20.600 8.800 29.800 9.100 ;
        RECT 38.200 9.100 38.600 9.200 ;
        RECT 55.800 9.100 56.200 9.200 ;
        RECT 66.200 9.100 66.600 9.200 ;
        RECT 38.200 8.800 66.600 9.100 ;
        RECT 71.000 9.100 71.400 9.200 ;
        RECT 79.800 9.100 80.200 9.200 ;
        RECT 84.600 9.100 85.000 9.200 ;
        RECT 71.000 8.800 85.000 9.100 ;
        RECT 92.600 9.100 93.000 9.200 ;
        RECT 95.800 9.100 96.200 9.200 ;
        RECT 104.600 9.100 105.000 9.200 ;
        RECT 92.600 8.800 105.000 9.100 ;
        RECT 117.400 9.100 117.800 9.200 ;
        RECT 166.200 9.100 166.600 9.200 ;
        RECT 168.600 9.100 169.000 9.200 ;
        RECT 117.400 8.800 120.100 9.100 ;
        RECT 166.200 8.800 169.000 9.100 ;
        RECT 175.800 9.100 176.200 9.200 ;
        RECT 179.000 9.100 179.400 9.200 ;
        RECT 175.800 8.800 179.400 9.100 ;
        RECT 189.400 9.100 189.800 9.200 ;
        RECT 200.600 9.100 201.000 9.200 ;
        RECT 189.400 8.800 201.000 9.100 ;
        RECT 204.600 9.100 205.000 9.200 ;
        RECT 225.400 9.100 225.800 9.200 ;
        RECT 242.200 9.100 242.600 9.200 ;
        RECT 243.800 9.100 244.200 9.200 ;
        RECT 246.200 9.100 246.600 9.200 ;
        RECT 204.600 8.800 246.600 9.100 ;
        RECT 119.800 8.200 120.100 8.800 ;
        RECT 64.600 8.100 65.000 8.200 ;
        RECT 72.600 8.100 73.000 8.200 ;
        RECT 96.600 8.100 97.000 8.200 ;
        RECT 97.400 8.100 97.800 8.200 ;
        RECT 64.600 7.800 97.800 8.100 ;
        RECT 119.800 7.800 120.200 8.200 ;
        RECT 127.800 8.100 128.200 8.200 ;
        RECT 131.800 8.100 132.200 8.200 ;
        RECT 143.000 8.100 143.400 8.200 ;
        RECT 151.000 8.100 151.400 8.200 ;
        RECT 157.400 8.100 157.800 8.200 ;
        RECT 127.800 7.800 157.800 8.100 ;
        RECT 161.400 8.100 161.800 8.200 ;
        RECT 168.600 8.100 169.000 8.200 ;
        RECT 161.400 7.800 169.000 8.100 ;
        RECT 171.000 8.100 171.400 8.200 ;
        RECT 177.400 8.100 177.800 8.200 ;
        RECT 171.000 7.800 177.800 8.100 ;
        RECT 179.000 8.100 179.400 8.200 ;
        RECT 191.000 8.100 191.400 8.200 ;
        RECT 179.000 7.800 191.400 8.100 ;
        RECT 211.000 8.100 211.400 8.200 ;
        RECT 218.200 8.100 218.600 8.200 ;
        RECT 219.800 8.100 220.200 8.200 ;
        RECT 211.000 7.800 220.200 8.100 ;
        RECT 7.800 7.100 8.200 7.200 ;
        RECT 8.600 7.100 9.000 7.200 ;
        RECT 7.800 6.800 9.000 7.100 ;
        RECT 25.400 7.100 25.800 7.200 ;
        RECT 31.800 7.100 32.200 7.200 ;
        RECT 25.400 6.800 32.200 7.100 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 35.000 7.100 35.400 7.200 ;
        RECT 38.200 7.100 38.600 7.200 ;
        RECT 35.000 6.800 38.600 7.100 ;
        RECT 40.600 7.100 41.000 7.200 ;
        RECT 49.400 7.100 49.800 7.200 ;
        RECT 55.800 7.100 56.200 7.200 ;
        RECT 40.600 6.800 56.200 7.100 ;
        RECT 68.600 7.100 69.000 7.200 ;
        RECT 74.200 7.100 74.600 7.200 ;
        RECT 68.600 6.800 74.600 7.100 ;
        RECT 87.800 7.100 88.200 7.200 ;
        RECT 93.400 7.100 93.800 7.200 ;
        RECT 87.800 6.800 93.800 7.100 ;
        RECT 101.400 7.100 101.800 7.200 ;
        RECT 109.400 7.100 109.800 7.200 ;
        RECT 101.400 6.800 109.800 7.100 ;
        RECT 113.400 7.100 113.800 7.200 ;
        RECT 171.800 7.100 172.200 7.200 ;
        RECT 113.400 6.800 172.200 7.100 ;
        RECT 191.000 7.100 191.300 7.800 ;
        RECT 206.200 7.100 206.600 7.200 ;
        RECT 191.000 6.800 206.600 7.100 ;
        RECT 215.000 6.800 215.400 7.200 ;
        RECT 227.000 6.800 227.400 7.200 ;
        RECT 256.600 6.800 257.000 7.200 ;
        RECT 259.800 6.800 260.200 7.200 ;
        RECT 32.600 6.200 32.900 6.800 ;
        RECT 113.400 6.200 113.700 6.800 ;
        RECT 9.400 5.800 9.800 6.200 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 32.600 6.100 33.000 6.200 ;
        RECT 92.600 6.100 93.000 6.200 ;
        RECT 94.200 6.100 94.600 6.200 ;
        RECT 102.200 6.100 102.600 6.200 ;
        RECT 31.000 5.800 102.600 6.100 ;
        RECT 104.600 6.100 105.000 6.200 ;
        RECT 111.800 6.100 112.200 6.200 ;
        RECT 104.600 5.800 112.200 6.100 ;
        RECT 113.400 5.800 113.800 6.200 ;
        RECT 117.400 6.100 117.800 6.200 ;
        RECT 124.600 6.100 125.000 6.200 ;
        RECT 117.400 5.800 125.000 6.100 ;
        RECT 131.000 6.100 131.400 6.200 ;
        RECT 134.200 6.100 134.600 6.200 ;
        RECT 131.000 5.800 134.600 6.100 ;
        RECT 155.000 6.100 155.400 6.200 ;
        RECT 173.400 6.100 173.800 6.200 ;
        RECT 155.000 5.800 173.800 6.100 ;
        RECT 175.800 6.100 176.200 6.200 ;
        RECT 176.600 6.100 177.000 6.200 ;
        RECT 175.800 5.800 177.000 6.100 ;
        RECT 180.600 6.100 181.000 6.200 ;
        RECT 187.800 6.100 188.200 6.200 ;
        RECT 180.600 5.800 188.200 6.100 ;
        RECT 206.200 6.100 206.600 6.200 ;
        RECT 215.000 6.100 215.300 6.800 ;
        RECT 206.200 5.800 215.300 6.100 ;
        RECT 227.000 6.100 227.300 6.800 ;
        RECT 234.200 6.100 234.600 6.200 ;
        RECT 227.000 5.800 234.600 6.100 ;
        RECT 251.800 6.100 252.200 6.200 ;
        RECT 256.600 6.100 256.900 6.800 ;
        RECT 251.800 5.800 256.900 6.100 ;
        RECT 259.800 6.100 260.100 6.800 ;
        RECT 263.000 6.100 263.400 6.200 ;
        RECT 259.800 5.800 263.400 6.100 ;
        RECT 9.400 5.100 9.700 5.800 ;
        RECT 11.800 5.100 12.200 5.200 ;
        RECT 9.400 4.800 12.200 5.100 ;
        RECT 27.800 5.100 28.200 5.200 ;
        RECT 35.000 5.100 35.400 5.200 ;
        RECT 27.800 4.800 35.400 5.100 ;
        RECT 62.200 5.100 62.600 5.200 ;
        RECT 130.200 5.100 130.600 5.200 ;
        RECT 62.200 4.800 130.600 5.100 ;
        RECT 132.600 5.100 133.000 5.200 ;
        RECT 139.000 5.100 139.400 5.200 ;
        RECT 132.600 4.800 139.400 5.100 ;
        RECT 214.200 5.100 214.600 5.200 ;
        RECT 217.400 5.100 217.800 5.200 ;
        RECT 250.200 5.100 250.600 5.200 ;
        RECT 214.200 4.800 250.600 5.100 ;
        RECT 62.200 4.100 62.600 4.200 ;
        RECT 115.000 4.100 115.400 4.200 ;
        RECT 117.400 4.100 117.800 4.200 ;
        RECT 62.200 3.800 117.800 4.100 ;
      LAYER via3 ;
        RECT 223.000 233.800 223.400 234.200 ;
        RECT 32.600 225.800 33.000 226.200 ;
        RECT 131.800 225.800 132.200 226.200 ;
        RECT 247.000 225.800 247.400 226.200 ;
        RECT 117.400 224.800 117.800 225.200 ;
        RECT 135.000 224.800 135.400 225.200 ;
        RECT 237.400 222.800 237.800 223.200 ;
        RECT 121.400 221.800 121.800 222.200 ;
        RECT 211.800 221.800 212.200 222.200 ;
        RECT 127.800 220.800 128.200 221.200 ;
        RECT 115.000 215.800 115.400 216.200 ;
        RECT 63.800 214.800 64.200 215.200 ;
        RECT 130.200 212.800 130.600 213.200 ;
        RECT 79.800 211.800 80.200 212.200 ;
        RECT 206.200 211.800 206.600 212.200 ;
        RECT 51.800 210.800 52.200 211.200 ;
        RECT 227.800 209.800 228.200 210.200 ;
        RECT 30.200 208.800 30.600 209.200 ;
        RECT 141.400 207.800 141.800 208.200 ;
        RECT 158.200 207.800 158.600 208.200 ;
        RECT 227.800 206.800 228.200 207.200 ;
        RECT 78.200 205.800 78.600 206.200 ;
        RECT 144.600 204.800 145.000 205.200 ;
        RECT 163.000 204.800 163.400 205.200 ;
        RECT 231.000 202.800 231.400 203.200 ;
        RECT 52.600 201.800 53.000 202.200 ;
        RECT 131.800 201.800 132.200 202.200 ;
        RECT 229.400 201.800 229.800 202.200 ;
        RECT 255.800 196.800 256.200 197.200 ;
        RECT 85.400 195.800 85.800 196.200 ;
        RECT 112.600 195.800 113.000 196.200 ;
        RECT 222.200 195.800 222.600 196.200 ;
        RECT 88.600 194.800 89.000 195.200 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 130.200 193.800 130.600 194.200 ;
        RECT 215.800 193.800 216.200 194.200 ;
        RECT 132.600 192.800 133.000 193.200 ;
        RECT 87.800 191.800 88.200 192.200 ;
        RECT 84.600 190.800 85.000 191.200 ;
        RECT 238.200 190.800 238.600 191.200 ;
        RECT 36.600 189.800 37.000 190.200 ;
        RECT 167.000 189.800 167.400 190.200 ;
        RECT 234.200 188.800 234.600 189.200 ;
        RECT 110.200 187.800 110.600 188.200 ;
        RECT 179.800 187.800 180.200 188.200 ;
        RECT 23.000 185.800 23.400 186.200 ;
        RECT 35.800 185.800 36.200 186.200 ;
        RECT 56.600 185.800 57.000 186.200 ;
        RECT 199.800 186.800 200.200 187.200 ;
        RECT 126.200 185.800 126.600 186.200 ;
        RECT 234.200 185.800 234.600 186.200 ;
        RECT 247.000 185.800 247.400 186.200 ;
        RECT 32.600 184.800 33.000 185.200 ;
        RECT 139.800 184.800 140.200 185.200 ;
        RECT 203.800 184.800 204.200 185.200 ;
        RECT 42.200 183.800 42.600 184.200 ;
        RECT 97.400 182.800 97.800 183.200 ;
        RECT 151.800 182.800 152.200 183.200 ;
        RECT 79.000 181.800 79.400 182.200 ;
        RECT 235.000 181.800 235.400 182.200 ;
        RECT 142.200 180.800 142.600 181.200 ;
        RECT 246.200 179.800 246.600 180.200 ;
        RECT 25.400 177.800 25.800 178.200 ;
        RECT 17.400 176.800 17.800 177.200 ;
        RECT 31.000 176.800 31.400 177.200 ;
        RECT 71.000 175.800 71.400 176.200 ;
        RECT 178.200 175.800 178.600 176.200 ;
        RECT 45.400 174.800 45.800 175.200 ;
        RECT 51.800 174.800 52.200 175.200 ;
        RECT 84.600 174.800 85.000 175.200 ;
        RECT 119.000 174.800 119.400 175.200 ;
        RECT 231.000 174.800 231.400 175.200 ;
        RECT 31.000 173.800 31.400 174.200 ;
        RECT 39.000 173.800 39.400 174.200 ;
        RECT 191.800 173.800 192.200 174.200 ;
        RECT 248.600 173.800 249.000 174.200 ;
        RECT 35.800 172.800 36.200 173.200 ;
        RECT 115.800 172.800 116.200 173.200 ;
        RECT 136.600 172.800 137.000 173.200 ;
        RECT 167.800 172.800 168.200 173.200 ;
        RECT 229.400 172.800 229.800 173.200 ;
        RECT 48.600 171.800 49.000 172.200 ;
        RECT 68.600 170.800 69.000 171.200 ;
        RECT 127.000 170.800 127.400 171.200 ;
        RECT 173.400 170.800 173.800 171.200 ;
        RECT 181.400 170.800 181.800 171.200 ;
        RECT 15.800 169.800 16.200 170.200 ;
        RECT 39.000 168.800 39.400 169.200 ;
        RECT 120.600 168.800 121.000 169.200 ;
        RECT 193.400 168.800 193.800 169.200 ;
        RECT 211.000 168.800 211.400 169.200 ;
        RECT 37.400 167.800 37.800 168.200 ;
        RECT 119.000 167.800 119.400 168.200 ;
        RECT 159.800 167.800 160.200 168.200 ;
        RECT 127.000 166.800 127.400 167.200 ;
        RECT 258.200 166.800 258.600 167.200 ;
        RECT 95.000 165.800 95.400 166.200 ;
        RECT 99.800 165.800 100.200 166.200 ;
        RECT 159.000 165.800 159.400 166.200 ;
        RECT 190.200 165.800 190.600 166.200 ;
        RECT 195.800 165.800 196.200 166.200 ;
        RECT 38.200 164.800 38.600 165.200 ;
        RECT 84.600 164.800 85.000 165.200 ;
        RECT 122.200 164.800 122.600 165.200 ;
        RECT 148.600 164.800 149.000 165.200 ;
        RECT 175.000 164.800 175.400 165.200 ;
        RECT 206.200 164.800 206.600 165.200 ;
        RECT 246.200 164.800 246.600 165.200 ;
        RECT 142.200 163.800 142.600 164.200 ;
        RECT 257.400 163.800 257.800 164.200 ;
        RECT 143.000 162.800 143.400 163.200 ;
        RECT 145.400 161.800 145.800 162.200 ;
        RECT 190.200 161.800 190.600 162.200 ;
        RECT 103.800 160.800 104.200 161.200 ;
        RECT 224.600 160.800 225.000 161.200 ;
        RECT 135.000 159.800 135.400 160.200 ;
        RECT 176.600 159.800 177.000 160.200 ;
        RECT 207.000 159.800 207.400 160.200 ;
        RECT 223.000 158.800 223.400 159.200 ;
        RECT 156.600 156.800 157.000 157.200 ;
        RECT 170.200 156.800 170.600 157.200 ;
        RECT 187.000 156.800 187.400 157.200 ;
        RECT 127.800 155.800 128.200 156.200 ;
        RECT 149.400 155.800 149.800 156.200 ;
        RECT 43.800 154.800 44.200 155.200 ;
        RECT 49.400 154.800 49.800 155.200 ;
        RECT 85.400 154.800 85.800 155.200 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 203.800 154.800 204.200 155.200 ;
        RECT 254.200 154.800 254.600 155.200 ;
        RECT 129.400 153.800 129.800 154.200 ;
        RECT 142.200 153.800 142.600 154.200 ;
        RECT 69.400 151.800 69.800 152.200 ;
        RECT 167.000 151.800 167.400 152.200 ;
        RECT 131.800 150.800 132.200 151.200 ;
        RECT 144.600 150.800 145.000 151.200 ;
        RECT 155.000 150.800 155.400 151.200 ;
        RECT 162.200 150.800 162.600 151.200 ;
        RECT 167.000 149.800 167.400 150.200 ;
        RECT 160.600 148.800 161.000 149.200 ;
        RECT 147.000 147.800 147.400 148.200 ;
        RECT 47.000 146.800 47.400 147.200 ;
        RECT 80.600 146.800 81.000 147.200 ;
        RECT 109.400 146.800 109.800 147.200 ;
        RECT 175.000 146.800 175.400 147.200 ;
        RECT 231.800 146.800 232.200 147.200 ;
        RECT 19.000 145.800 19.400 146.200 ;
        RECT 71.800 145.800 72.200 146.200 ;
        RECT 75.000 145.800 75.400 146.200 ;
        RECT 93.400 145.800 93.800 146.200 ;
        RECT 101.400 145.800 101.800 146.200 ;
        RECT 182.200 145.800 182.600 146.200 ;
        RECT 100.600 144.800 101.000 145.200 ;
        RECT 187.800 144.800 188.200 145.200 ;
        RECT 248.600 144.800 249.000 145.200 ;
        RECT 107.800 143.800 108.200 144.200 ;
        RECT 121.400 143.800 121.800 144.200 ;
        RECT 143.000 143.800 143.400 144.200 ;
        RECT 163.000 143.800 163.400 144.200 ;
        RECT 52.600 142.800 53.000 143.200 ;
        RECT 60.600 142.800 61.000 143.200 ;
        RECT 226.200 142.800 226.600 143.200 ;
        RECT 263.000 142.800 263.400 143.200 ;
        RECT 72.600 141.800 73.000 142.200 ;
        RECT 84.600 141.800 85.000 142.200 ;
        RECT 140.600 141.800 141.000 142.200 ;
        RECT 148.600 141.800 149.000 142.200 ;
        RECT 146.200 140.800 146.600 141.200 ;
        RECT 155.000 140.800 155.400 141.200 ;
        RECT 132.600 139.800 133.000 140.200 ;
        RECT 180.600 139.800 181.000 140.200 ;
        RECT 158.200 138.800 158.600 139.200 ;
        RECT 33.400 137.800 33.800 138.200 ;
        RECT 28.600 136.800 29.000 137.200 ;
        RECT 86.200 136.800 86.600 137.200 ;
        RECT 90.200 136.800 90.600 137.200 ;
        RECT 105.400 136.800 105.800 137.200 ;
        RECT 258.200 136.800 258.600 137.200 ;
        RECT 110.200 135.800 110.600 136.200 ;
        RECT 131.000 135.800 131.400 136.200 ;
        RECT 152.600 135.800 153.000 136.200 ;
        RECT 168.600 135.800 169.000 136.200 ;
        RECT 180.600 135.800 181.000 136.200 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 216.600 135.800 217.000 136.200 ;
        RECT 238.200 135.800 238.600 136.200 ;
        RECT 56.600 134.800 57.000 135.200 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 108.600 134.800 109.000 135.200 ;
        RECT 111.800 134.800 112.200 135.200 ;
        RECT 132.600 134.800 133.000 135.200 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 203.800 134.800 204.200 135.200 ;
        RECT 53.400 133.800 53.800 134.200 ;
        RECT 139.000 133.800 139.400 134.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 211.000 133.800 211.400 134.200 ;
        RECT 28.600 132.800 29.000 133.200 ;
        RECT 71.800 132.800 72.200 133.200 ;
        RECT 103.800 132.800 104.200 133.200 ;
        RECT 115.800 132.800 116.200 133.200 ;
        RECT 154.200 132.800 154.600 133.200 ;
        RECT 163.800 132.800 164.200 133.200 ;
        RECT 194.200 132.800 194.600 133.200 ;
        RECT 176.600 130.800 177.000 131.200 ;
        RECT 207.000 130.800 207.400 131.200 ;
        RECT 38.200 129.800 38.600 130.200 ;
        RECT 70.200 129.800 70.600 130.200 ;
        RECT 29.400 128.800 29.800 129.200 ;
        RECT 47.000 128.800 47.400 129.200 ;
        RECT 102.200 128.800 102.600 129.200 ;
        RECT 210.200 128.800 210.600 129.200 ;
        RECT 39.000 126.800 39.400 127.200 ;
        RECT 104.600 126.800 105.000 127.200 ;
        RECT 111.800 126.800 112.200 127.200 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 89.400 125.800 89.800 126.200 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 171.800 125.800 172.200 126.200 ;
        RECT 205.400 125.800 205.800 126.200 ;
        RECT 66.200 124.800 66.600 125.200 ;
        RECT 107.800 124.800 108.200 125.200 ;
        RECT 196.600 124.800 197.000 125.200 ;
        RECT 47.800 123.800 48.200 124.200 ;
        RECT 67.000 123.800 67.400 124.200 ;
        RECT 116.600 123.800 117.000 124.200 ;
        RECT 143.000 123.800 143.400 124.200 ;
        RECT 64.600 122.800 65.000 123.200 ;
        RECT 73.400 122.800 73.800 123.200 ;
        RECT 125.400 122.800 125.800 123.200 ;
        RECT 166.200 122.800 166.600 123.200 ;
        RECT 244.600 122.800 245.000 123.200 ;
        RECT 135.000 121.800 135.400 122.200 ;
        RECT 88.600 120.800 89.000 121.200 ;
        RECT 202.200 120.800 202.600 121.200 ;
        RECT 231.000 119.800 231.400 120.200 ;
        RECT 147.800 118.800 148.200 119.200 ;
        RECT 146.200 117.800 146.600 118.200 ;
        RECT 237.400 117.800 237.800 118.200 ;
        RECT 247.800 117.800 248.200 118.200 ;
        RECT 63.800 115.800 64.200 116.200 ;
        RECT 87.800 115.800 88.200 116.200 ;
        RECT 139.800 115.800 140.200 116.200 ;
        RECT 159.000 115.800 159.400 116.200 ;
        RECT 232.600 115.800 233.000 116.200 ;
        RECT 130.200 114.800 130.600 115.200 ;
        RECT 203.000 114.800 203.400 115.200 ;
        RECT 69.400 113.800 69.800 114.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 79.000 112.800 79.400 113.200 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 91.800 111.800 92.200 112.200 ;
        RECT 257.400 111.800 257.800 112.200 ;
        RECT 42.200 110.800 42.600 111.200 ;
        RECT 51.800 110.800 52.200 111.200 ;
        RECT 92.600 109.800 93.000 110.200 ;
        RECT 173.400 109.800 173.800 110.200 ;
        RECT 25.400 107.800 25.800 108.200 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 144.600 107.800 145.000 108.200 ;
        RECT 160.600 107.800 161.000 108.200 ;
        RECT 167.800 107.800 168.200 108.200 ;
        RECT 141.400 106.800 141.800 107.200 ;
        RECT 165.400 106.800 165.800 107.200 ;
        RECT 239.800 106.800 240.200 107.200 ;
        RECT 88.600 105.800 89.000 106.200 ;
        RECT 153.400 105.800 153.800 106.200 ;
        RECT 167.000 105.800 167.400 106.200 ;
        RECT 212.600 104.800 213.000 105.200 ;
        RECT 164.600 103.800 165.000 104.200 ;
        RECT 187.000 103.800 187.400 104.200 ;
        RECT 94.200 102.800 94.600 103.200 ;
        RECT 200.600 101.800 201.000 102.200 ;
        RECT 199.800 100.800 200.200 101.200 ;
        RECT 47.000 99.800 47.400 100.200 ;
        RECT 80.600 99.800 81.000 100.200 ;
        RECT 41.400 98.800 41.800 99.200 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 161.400 98.800 161.800 99.200 ;
        RECT 58.200 97.800 58.600 98.200 ;
        RECT 71.000 97.800 71.400 98.200 ;
        RECT 195.800 96.800 196.200 97.200 ;
        RECT 42.200 95.800 42.600 96.200 ;
        RECT 248.600 95.800 249.000 96.200 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 32.600 94.800 33.000 95.200 ;
        RECT 131.000 94.800 131.400 95.200 ;
        RECT 181.400 94.800 181.800 95.200 ;
        RECT 71.000 93.800 71.400 94.200 ;
        RECT 142.200 93.800 142.600 94.200 ;
        RECT 24.600 92.800 25.000 93.200 ;
        RECT 89.400 91.800 89.800 92.200 ;
        RECT 103.800 91.800 104.200 92.200 ;
        RECT 184.600 91.800 185.000 92.200 ;
        RECT 187.800 91.800 188.200 92.200 ;
        RECT 121.400 89.800 121.800 90.200 ;
        RECT 174.200 88.800 174.600 89.200 ;
        RECT 257.400 87.800 257.800 88.200 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 147.800 86.800 148.200 87.200 ;
        RECT 189.400 86.800 189.800 87.200 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 172.600 85.800 173.000 86.200 ;
        RECT 216.600 85.800 217.000 86.200 ;
        RECT 160.600 84.800 161.000 85.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 163.000 83.800 163.400 84.200 ;
        RECT 163.800 81.800 164.200 82.200 ;
        RECT 197.400 81.800 197.800 82.200 ;
        RECT 221.400 81.800 221.800 82.200 ;
        RECT 25.400 80.800 25.800 81.200 ;
        RECT 182.200 80.800 182.600 81.200 ;
        RECT 223.800 80.800 224.200 81.200 ;
        RECT 231.800 80.800 232.200 81.200 ;
        RECT 235.000 80.800 235.400 81.200 ;
        RECT 132.600 78.800 133.000 79.200 ;
        RECT 207.000 77.800 207.400 78.200 ;
        RECT 223.000 77.800 223.400 78.200 ;
        RECT 47.000 76.800 47.400 77.200 ;
        RECT 125.400 76.800 125.800 77.200 ;
        RECT 156.600 76.800 157.000 77.200 ;
        RECT 18.200 75.800 18.600 76.200 ;
        RECT 127.800 75.800 128.200 76.200 ;
        RECT 231.000 75.800 231.400 76.200 ;
        RECT 107.000 74.800 107.400 75.200 ;
        RECT 176.600 74.800 177.000 75.200 ;
        RECT 198.200 74.800 198.600 75.200 ;
        RECT 210.200 74.800 210.600 75.200 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 189.400 73.800 189.800 74.200 ;
        RECT 88.600 72.800 89.000 73.200 ;
        RECT 109.400 72.800 109.800 73.200 ;
        RECT 64.600 71.800 65.000 72.200 ;
        RECT 130.200 71.800 130.600 72.200 ;
        RECT 170.200 71.800 170.600 72.200 ;
        RECT 229.400 71.800 229.800 72.200 ;
        RECT 70.200 70.800 70.600 71.200 ;
        RECT 165.400 70.800 165.800 71.200 ;
        RECT 95.000 69.800 95.400 70.200 ;
        RECT 134.200 69.800 134.600 70.200 ;
        RECT 206.200 69.800 206.600 70.200 ;
        RECT 140.600 68.800 141.000 69.200 ;
        RECT 242.200 68.800 242.600 69.200 ;
        RECT 40.600 67.800 41.000 68.200 ;
        RECT 129.400 67.800 129.800 68.200 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 111.800 66.800 112.200 67.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 124.600 65.800 125.000 66.200 ;
        RECT 196.600 65.800 197.000 66.200 ;
        RECT 203.000 65.800 203.400 66.200 ;
        RECT 91.000 64.800 91.400 65.200 ;
        RECT 135.800 64.800 136.200 65.200 ;
        RECT 45.400 63.800 45.800 64.200 ;
        RECT 48.600 63.800 49.000 64.200 ;
        RECT 79.800 61.800 80.200 62.200 ;
        RECT 89.400 61.800 89.800 62.200 ;
        RECT 137.400 61.800 137.800 62.200 ;
        RECT 216.600 61.800 217.000 62.200 ;
        RECT 53.400 60.800 53.800 61.200 ;
        RECT 211.000 60.800 211.400 61.200 ;
        RECT 139.800 59.800 140.200 60.200 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 43.000 56.800 43.400 57.200 ;
        RECT 187.000 56.800 187.400 57.200 ;
        RECT 259.800 55.800 260.200 56.200 ;
        RECT 19.800 54.800 20.200 55.200 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 115.000 54.800 115.400 55.200 ;
        RECT 142.200 54.800 142.600 55.200 ;
        RECT 69.400 51.800 69.800 52.200 ;
        RECT 146.200 51.800 146.600 52.200 ;
        RECT 127.800 50.800 128.200 51.200 ;
        RECT 129.400 49.800 129.800 50.200 ;
        RECT 132.600 48.800 133.000 49.200 ;
        RECT 131.800 47.800 132.200 48.200 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 131.000 46.800 131.400 47.200 ;
        RECT 58.200 45.800 58.600 46.200 ;
        RECT 143.800 45.800 144.200 46.200 ;
        RECT 159.000 45.800 159.400 46.200 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 62.200 44.800 62.600 45.200 ;
        RECT 254.200 44.800 254.600 45.200 ;
        RECT 243.000 43.800 243.400 44.200 ;
        RECT 108.600 42.800 109.000 43.200 ;
        RECT 95.800 41.800 96.200 42.200 ;
        RECT 180.600 41.800 181.000 42.200 ;
        RECT 243.800 41.800 244.200 42.200 ;
        RECT 103.800 40.800 104.200 41.200 ;
        RECT 206.200 39.800 206.600 40.200 ;
        RECT 259.800 39.800 260.200 40.200 ;
        RECT 122.200 38.800 122.600 39.200 ;
        RECT 84.600 37.800 85.000 38.200 ;
        RECT 88.600 37.800 89.000 38.200 ;
        RECT 167.800 37.800 168.200 38.200 ;
        RECT 12.600 36.800 13.000 37.200 ;
        RECT 111.000 36.800 111.400 37.200 ;
        RECT 39.000 35.800 39.400 36.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 63.800 34.800 64.200 35.200 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 102.200 34.800 102.600 35.200 ;
        RECT 188.600 34.800 189.000 35.200 ;
        RECT 23.000 33.800 23.400 34.200 ;
        RECT 175.000 33.800 175.400 34.200 ;
        RECT 201.400 33.800 201.800 34.200 ;
        RECT 160.600 32.800 161.000 33.200 ;
        RECT 255.000 32.800 255.400 33.200 ;
        RECT 124.600 31.800 125.000 32.200 ;
        RECT 63.000 30.800 63.400 31.200 ;
        RECT 172.600 28.800 173.000 29.200 ;
        RECT 221.400 28.800 221.800 29.200 ;
        RECT 54.200 26.800 54.600 27.200 ;
        RECT 247.000 24.800 247.400 25.200 ;
        RECT 237.400 19.800 237.800 20.200 ;
        RECT 7.800 18.800 8.200 19.200 ;
        RECT 97.400 18.800 97.800 19.200 ;
        RECT 159.800 17.800 160.200 18.200 ;
        RECT 251.800 17.800 252.200 18.200 ;
        RECT 19.800 16.800 20.200 17.200 ;
        RECT 232.600 16.800 233.000 17.200 ;
        RECT 92.600 15.800 93.000 16.200 ;
        RECT 94.200 15.800 94.600 16.200 ;
        RECT 252.600 15.800 253.000 16.200 ;
        RECT 62.200 14.800 62.600 15.200 ;
        RECT 99.800 14.800 100.200 15.200 ;
        RECT 220.600 14.800 221.000 15.200 ;
        RECT 84.600 8.800 85.000 9.200 ;
        RECT 179.000 8.800 179.400 9.200 ;
        RECT 96.600 7.800 97.000 8.200 ;
        RECT 219.800 7.800 220.200 8.200 ;
        RECT 176.600 5.800 177.000 6.200 ;
        RECT 11.800 4.800 12.200 5.200 ;
      LAYER metal4 ;
        RECT 32.600 235.800 33.000 236.200 ;
        RECT 32.600 226.200 32.900 235.800 ;
        RECT 223.000 234.100 223.400 234.200 ;
        RECT 222.200 233.800 223.400 234.100 ;
        RECT 129.400 229.800 129.800 230.200 ;
        RECT 32.600 225.800 33.000 226.200 ;
        RECT 51.800 225.800 52.200 226.200 ;
        RECT 125.400 226.100 125.800 226.200 ;
        RECT 126.200 226.100 126.600 226.200 ;
        RECT 125.400 225.800 126.600 226.100 ;
        RECT 31.000 211.800 31.400 212.200 ;
        RECT 30.200 208.800 30.600 209.200 ;
        RECT 30.200 206.200 30.500 208.800 ;
        RECT 30.200 205.800 30.600 206.200 ;
        RECT 17.400 202.800 17.800 203.200 ;
        RECT 17.400 177.200 17.700 202.800 ;
        RECT 19.000 195.800 19.400 196.200 ;
        RECT 17.400 176.800 17.800 177.200 ;
        RECT 15.800 169.800 16.200 170.200 ;
        RECT 11.800 99.800 12.200 100.200 ;
        RECT 7.800 18.800 8.200 19.200 ;
        RECT 7.800 7.200 8.100 18.800 ;
        RECT 11.800 15.200 12.100 99.800 ;
        RECT 15.800 95.200 16.100 169.800 ;
        RECT 19.000 146.200 19.300 195.800 ;
        RECT 23.000 185.800 23.400 186.200 ;
        RECT 19.000 146.100 19.400 146.200 ;
        RECT 19.000 145.800 20.100 146.100 ;
        RECT 16.600 141.800 17.000 142.200 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 16.600 86.100 16.900 141.800 ;
        RECT 18.200 115.800 18.600 116.200 ;
        RECT 17.400 86.100 17.800 86.200 ;
        RECT 16.600 85.800 17.800 86.100 ;
        RECT 12.600 74.800 13.000 75.200 ;
        RECT 12.600 37.200 12.900 74.800 ;
        RECT 16.600 56.200 16.900 85.800 ;
        RECT 18.200 76.200 18.500 115.800 ;
        RECT 19.000 98.800 19.400 99.200 ;
        RECT 18.200 75.800 18.600 76.200 ;
        RECT 16.600 55.800 17.000 56.200 ;
        RECT 16.600 47.200 16.900 55.800 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 12.600 36.800 13.000 37.200 ;
        RECT 19.000 17.100 19.300 98.800 ;
        RECT 19.800 55.200 20.100 145.800 ;
        RECT 23.000 112.200 23.300 185.800 ;
        RECT 25.400 177.800 25.800 178.200 ;
        RECT 23.000 111.800 23.400 112.200 ;
        RECT 19.800 54.800 20.200 55.200 ;
        RECT 19.800 18.200 20.100 54.800 ;
        RECT 23.000 34.200 23.300 111.800 ;
        RECT 25.400 108.200 25.700 177.800 ;
        RECT 31.000 177.200 31.300 211.800 ;
        RECT 31.800 205.800 32.200 206.200 ;
        RECT 31.000 176.800 31.400 177.200 ;
        RECT 31.000 173.800 31.400 174.200 ;
        RECT 27.800 137.100 28.200 137.200 ;
        RECT 28.600 137.100 29.000 137.200 ;
        RECT 27.800 136.800 29.000 137.100 ;
        RECT 30.200 133.800 30.600 134.200 ;
        RECT 28.600 133.100 29.000 133.200 ;
        RECT 29.400 133.100 29.800 133.200 ;
        RECT 28.600 132.800 29.800 133.100 ;
        RECT 30.200 132.200 30.500 133.800 ;
        RECT 30.200 131.800 30.600 132.200 ;
        RECT 29.400 128.800 29.800 129.200 ;
        RECT 29.400 128.200 29.700 128.800 ;
        RECT 30.200 128.200 30.500 131.800 ;
        RECT 31.000 129.200 31.300 173.800 ;
        RECT 31.800 131.200 32.100 205.800 ;
        RECT 32.600 185.200 32.900 225.800 ;
        RECT 51.800 211.200 52.100 225.800 ;
        RECT 117.400 224.800 117.800 225.200 ;
        RECT 111.000 220.800 111.400 221.200 ;
        RECT 63.800 214.800 64.200 215.200 ;
        RECT 51.800 210.800 52.200 211.200 ;
        RECT 35.800 209.800 36.200 210.200 ;
        RECT 33.400 204.800 33.800 205.200 ;
        RECT 32.600 184.800 33.000 185.200 ;
        RECT 33.400 138.200 33.700 204.800 ;
        RECT 35.800 186.200 36.100 209.800 ;
        RECT 44.600 206.100 45.000 206.200 ;
        RECT 45.400 206.100 45.800 206.200 ;
        RECT 44.600 205.800 45.800 206.100 ;
        RECT 42.200 192.800 42.600 193.200 ;
        RECT 43.800 192.800 44.200 193.200 ;
        RECT 36.600 189.800 37.000 190.200 ;
        RECT 35.800 185.800 36.200 186.200 ;
        RECT 35.800 173.800 36.200 174.200 ;
        RECT 35.800 173.200 36.100 173.800 ;
        RECT 35.800 172.800 36.200 173.200 ;
        RECT 36.600 168.100 36.900 189.800 ;
        RECT 41.400 185.800 41.800 186.200 ;
        RECT 39.000 176.800 39.400 177.200 ;
        RECT 39.000 174.200 39.300 176.800 ;
        RECT 39.000 173.800 39.400 174.200 ;
        RECT 39.800 173.800 40.200 174.200 ;
        RECT 39.800 173.200 40.100 173.800 ;
        RECT 39.800 172.800 40.200 173.200 ;
        RECT 39.000 168.800 39.400 169.200 ;
        RECT 37.400 168.100 37.800 168.200 ;
        RECT 36.600 167.800 37.800 168.100 ;
        RECT 39.000 166.200 39.300 168.800 ;
        RECT 39.000 165.800 39.400 166.200 ;
        RECT 38.200 164.800 38.600 165.200 ;
        RECT 33.400 137.800 33.800 138.200 ;
        RECT 35.800 136.800 36.200 137.200 ;
        RECT 31.800 130.800 32.200 131.200 ;
        RECT 31.000 128.800 31.400 129.200 ;
        RECT 29.400 127.800 29.800 128.200 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 31.000 126.200 31.300 128.800 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 31.800 113.200 32.100 130.800 ;
        RECT 35.800 118.200 36.100 136.800 ;
        RECT 38.200 130.200 38.500 164.800 ;
        RECT 38.200 129.800 38.600 130.200 ;
        RECT 38.200 127.100 38.500 129.800 ;
        RECT 39.000 127.100 39.400 127.200 ;
        RECT 38.200 126.800 39.400 127.100 ;
        RECT 35.800 117.800 36.200 118.200 ;
        RECT 31.800 112.800 32.200 113.200 ;
        RECT 25.400 107.800 25.800 108.200 ;
        RECT 24.600 93.100 25.000 93.200 ;
        RECT 23.800 92.800 25.000 93.100 ;
        RECT 23.800 79.200 24.100 92.800 ;
        RECT 25.400 84.200 25.700 107.800 ;
        RECT 25.400 83.800 25.800 84.200 ;
        RECT 25.400 80.800 25.800 81.200 ;
        RECT 23.800 78.800 24.200 79.200 ;
        RECT 23.800 67.200 24.100 78.800 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 23.000 33.800 23.400 34.200 ;
        RECT 25.400 23.200 25.700 80.800 ;
        RECT 31.800 76.200 32.100 112.800 ;
        RECT 32.600 94.800 33.000 95.200 ;
        RECT 31.800 75.800 32.200 76.200 ;
        RECT 31.800 46.200 32.100 75.800 ;
        RECT 31.800 45.800 32.200 46.200 ;
        RECT 25.400 22.800 25.800 23.200 ;
        RECT 19.800 17.800 20.200 18.200 ;
        RECT 19.800 17.100 20.200 17.200 ;
        RECT 19.000 16.800 20.200 17.100 ;
        RECT 11.800 14.800 12.200 15.200 ;
        RECT 7.800 6.800 8.200 7.200 ;
        RECT 11.800 5.200 12.100 14.800 ;
        RECT 32.600 7.200 32.900 94.800 ;
        RECT 39.000 93.200 39.300 126.800 ;
        RECT 41.400 99.200 41.700 185.800 ;
        RECT 42.200 184.200 42.500 192.800 ;
        RECT 42.200 183.800 42.600 184.200 ;
        RECT 42.200 130.200 42.500 183.800 ;
        RECT 43.800 155.200 44.100 192.800 ;
        RECT 51.800 175.200 52.100 210.800 ;
        RECT 52.600 201.800 53.000 202.200 ;
        RECT 44.600 175.100 45.000 175.200 ;
        RECT 45.400 175.100 45.800 175.200 ;
        RECT 44.600 174.800 45.800 175.100 ;
        RECT 47.000 174.800 47.400 175.200 ;
        RECT 51.800 174.800 52.200 175.200 ;
        RECT 47.000 174.200 47.300 174.800 ;
        RECT 47.000 173.800 47.400 174.200 ;
        RECT 48.600 172.800 49.000 173.200 ;
        RECT 48.600 172.200 48.900 172.800 ;
        RECT 48.600 171.800 49.000 172.200 ;
        RECT 51.800 167.200 52.100 174.800 ;
        RECT 52.600 174.200 52.900 201.800 ;
        RECT 56.600 185.800 57.000 186.200 ;
        RECT 56.600 179.200 56.900 185.800 ;
        RECT 56.600 178.800 57.000 179.200 ;
        RECT 52.600 173.800 53.000 174.200 ;
        RECT 51.800 166.800 52.200 167.200 ;
        RECT 43.800 154.800 44.200 155.200 ;
        RECT 49.400 154.800 49.800 155.200 ;
        RECT 47.000 147.100 47.400 147.200 ;
        RECT 47.800 147.100 48.200 147.200 ;
        RECT 47.000 146.800 48.200 147.100 ;
        RECT 42.200 129.800 42.600 130.200 ;
        RECT 47.000 128.800 47.400 129.200 ;
        RECT 44.600 128.100 45.000 128.200 ;
        RECT 45.400 128.100 45.800 128.200 ;
        RECT 44.600 127.800 45.800 128.100 ;
        RECT 47.000 119.200 47.300 128.800 ;
        RECT 47.800 124.800 48.200 125.200 ;
        RECT 47.800 124.200 48.100 124.800 ;
        RECT 47.800 123.800 48.200 124.200 ;
        RECT 47.000 118.800 47.400 119.200 ;
        RECT 47.000 115.800 47.400 116.200 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 42.200 110.800 42.600 111.200 ;
        RECT 41.400 98.800 41.800 99.200 ;
        RECT 42.200 96.200 42.500 110.800 ;
        RECT 42.200 95.800 42.600 96.200 ;
        RECT 39.000 92.800 39.400 93.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 35.000 63.200 35.300 65.800 ;
        RECT 35.000 62.800 35.400 63.200 ;
        RECT 39.000 36.200 39.300 92.800 ;
        RECT 40.600 68.100 41.000 68.200 ;
        RECT 41.400 68.100 41.800 68.200 ;
        RECT 40.600 67.800 41.800 68.100 ;
        RECT 43.000 57.200 43.300 111.800 ;
        RECT 47.000 100.200 47.300 115.800 ;
        RECT 47.000 99.800 47.400 100.200 ;
        RECT 47.000 76.800 47.400 77.200 ;
        RECT 45.400 64.100 45.800 64.200 ;
        RECT 46.200 64.100 46.600 64.200 ;
        RECT 45.400 63.800 46.600 64.100 ;
        RECT 43.000 56.800 43.400 57.200 ;
        RECT 47.000 54.200 47.300 76.800 ;
        RECT 48.600 64.800 49.000 65.200 ;
        RECT 48.600 64.200 48.900 64.800 ;
        RECT 48.600 63.800 49.000 64.200 ;
        RECT 49.400 63.200 49.700 154.800 ;
        RECT 50.200 117.800 50.600 118.200 ;
        RECT 50.200 66.200 50.500 117.800 ;
        RECT 51.800 111.200 52.100 166.800 ;
        RECT 52.600 143.200 52.900 173.800 ;
        RECT 52.600 142.800 53.000 143.200 ;
        RECT 56.600 135.200 56.900 178.800 ;
        RECT 60.600 142.800 61.000 143.200 ;
        RECT 56.600 134.800 57.000 135.200 ;
        RECT 53.400 133.800 53.800 134.200 ;
        RECT 53.400 115.200 53.700 133.800 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 51.800 110.800 52.200 111.200 ;
        RECT 58.200 97.800 58.600 98.200 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 55.800 65.800 57.000 66.100 ;
        RECT 57.400 65.800 57.800 66.200 ;
        RECT 57.400 65.200 57.700 65.800 ;
        RECT 57.400 64.800 57.800 65.200 ;
        RECT 53.400 63.800 53.800 64.200 ;
        RECT 49.400 62.800 49.800 63.200 ;
        RECT 53.400 61.200 53.700 63.800 ;
        RECT 53.400 60.800 53.800 61.200 ;
        RECT 47.000 53.800 47.400 54.200 ;
        RECT 58.200 46.200 58.500 97.800 ;
        RECT 58.200 45.800 58.600 46.200 ;
        RECT 39.000 35.800 39.400 36.200 ;
        RECT 60.600 35.200 60.900 142.800 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 62.200 45.100 62.600 45.200 ;
        RECT 61.400 44.800 62.600 45.100 ;
        RECT 59.800 35.100 60.200 35.200 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 59.800 34.800 61.000 35.100 ;
        RECT 61.400 34.200 61.700 44.800 ;
        RECT 63.000 35.100 63.300 134.800 ;
        RECT 63.800 116.200 64.100 214.800 ;
        RECT 79.800 211.800 80.200 212.200 ;
        RECT 79.800 207.200 80.100 211.800 ;
        RECT 79.800 206.800 80.200 207.200 ;
        RECT 78.200 205.800 78.600 206.200 ;
        RECT 68.600 185.800 69.000 186.200 ;
        RECT 64.600 184.800 65.000 185.200 ;
        RECT 64.600 123.200 64.900 184.800 ;
        RECT 68.600 171.200 68.900 185.800 ;
        RECT 71.800 180.800 72.200 181.200 ;
        RECT 71.000 175.800 71.400 176.200 ;
        RECT 68.600 170.800 69.000 171.200 ;
        RECT 69.400 151.800 69.800 152.200 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 65.400 125.100 65.700 125.800 ;
        RECT 66.200 125.100 66.600 125.200 ;
        RECT 65.400 124.800 66.600 125.100 ;
        RECT 67.000 123.800 67.400 124.200 ;
        RECT 64.600 122.800 65.000 123.200 ;
        RECT 63.800 115.800 64.200 116.200 ;
        RECT 65.400 86.800 65.800 87.200 ;
        RECT 64.600 71.800 65.000 72.200 ;
        RECT 64.600 66.200 64.900 71.800 ;
        RECT 65.400 66.200 65.700 86.800 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 66.200 66.200 66.500 66.800 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 67.000 36.200 67.300 123.800 ;
        RECT 69.400 114.200 69.700 151.800 ;
        RECT 71.000 143.200 71.300 175.800 ;
        RECT 71.800 146.200 72.100 180.800 ;
        RECT 75.800 166.100 76.200 166.200 ;
        RECT 76.600 166.100 77.000 166.200 ;
        RECT 75.800 165.800 77.000 166.100 ;
        RECT 71.800 145.800 72.200 146.200 ;
        RECT 75.000 145.800 75.400 146.200 ;
        RECT 71.000 142.800 71.400 143.200 ;
        RECT 70.200 129.800 70.600 130.200 ;
        RECT 69.400 113.800 69.800 114.200 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 67.800 57.200 68.100 98.800 ;
        RECT 70.200 97.200 70.500 129.800 ;
        RECT 71.000 98.200 71.300 142.800 ;
        RECT 72.600 141.800 73.000 142.200 ;
        RECT 72.600 138.200 72.900 141.800 ;
        RECT 72.600 137.800 73.000 138.200 ;
        RECT 71.800 132.800 72.200 133.200 ;
        RECT 71.800 128.200 72.100 132.800 ;
        RECT 71.800 127.800 72.200 128.200 ;
        RECT 73.400 122.800 73.800 123.200 ;
        RECT 71.000 97.800 71.400 98.200 ;
        RECT 70.200 96.800 70.600 97.200 ;
        RECT 70.200 71.200 70.500 96.800 ;
        RECT 71.000 94.200 71.300 97.800 ;
        RECT 71.000 93.800 71.400 94.200 ;
        RECT 70.200 70.800 70.600 71.200 ;
        RECT 70.200 66.100 70.500 70.800 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 73.400 58.200 73.700 122.800 ;
        RECT 75.000 87.200 75.300 145.800 ;
        RECT 78.200 126.200 78.500 205.800 ;
        RECT 90.200 201.800 90.600 202.200 ;
        RECT 88.600 198.800 89.000 199.200 ;
        RECT 85.400 195.800 85.800 196.200 ;
        RECT 79.800 193.100 80.200 193.200 ;
        RECT 80.600 193.100 81.000 193.200 ;
        RECT 79.800 192.800 81.000 193.100 ;
        RECT 84.600 190.800 85.000 191.200 ;
        RECT 79.000 181.800 79.400 182.200 ;
        RECT 79.000 155.200 79.300 181.800 ;
        RECT 84.600 175.200 84.900 190.800 ;
        RECT 81.400 174.800 81.800 175.200 ;
        RECT 84.600 174.800 85.000 175.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 75.800 125.800 76.200 126.200 ;
        RECT 78.200 125.800 78.600 126.200 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 75.800 86.200 76.100 125.800 ;
        RECT 79.000 113.200 79.300 154.800 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 80.600 147.100 81.000 147.200 ;
        RECT 79.800 146.800 81.000 147.100 ;
        RECT 81.400 144.200 81.700 174.800 ;
        RECT 84.600 164.800 85.000 165.200 ;
        RECT 84.600 149.200 84.900 164.800 ;
        RECT 85.400 155.200 85.700 195.800 ;
        RECT 88.600 195.200 88.900 198.800 ;
        RECT 88.600 194.800 89.000 195.200 ;
        RECT 87.800 191.800 88.200 192.200 ;
        RECT 85.400 154.800 85.800 155.200 ;
        RECT 84.600 148.800 85.000 149.200 ;
        RECT 81.400 143.800 81.800 144.200 ;
        RECT 81.400 126.200 81.700 143.800 ;
        RECT 84.600 141.800 85.000 142.200 ;
        RECT 81.400 125.800 81.800 126.200 ;
        RECT 84.600 118.200 84.900 141.800 ;
        RECT 87.800 140.200 88.100 191.800 ;
        RECT 88.600 157.800 89.000 158.200 ;
        RECT 87.800 139.800 88.200 140.200 ;
        RECT 86.200 136.800 86.600 137.200 ;
        RECT 85.400 126.800 85.800 127.200 ;
        RECT 85.400 126.200 85.700 126.800 ;
        RECT 85.400 125.800 85.800 126.200 ;
        RECT 84.600 117.800 85.000 118.200 ;
        RECT 79.000 112.800 79.400 113.200 ;
        RECT 80.600 100.100 81.000 100.200 ;
        RECT 79.800 99.800 81.000 100.100 ;
        RECT 75.800 85.800 76.200 86.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 74.200 64.200 74.500 65.800 ;
        RECT 74.200 63.800 74.600 64.200 ;
        RECT 79.800 62.200 80.100 99.800 ;
        RECT 80.600 87.800 81.000 88.200 ;
        RECT 79.800 61.800 80.200 62.200 ;
        RECT 68.600 58.100 69.000 58.200 ;
        RECT 68.600 57.800 69.700 58.100 ;
        RECT 73.400 57.800 73.800 58.200 ;
        RECT 67.800 56.800 68.200 57.200 ;
        RECT 69.400 52.200 69.700 57.800 ;
        RECT 69.400 51.800 69.800 52.200 ;
        RECT 80.600 36.200 80.900 87.800 ;
        RECT 84.600 38.200 84.900 117.800 ;
        RECT 84.600 37.800 85.000 38.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 63.800 35.100 64.200 35.200 ;
        RECT 63.000 34.800 64.200 35.100 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 63.000 31.200 63.300 34.800 ;
        RECT 63.000 30.800 63.400 31.200 ;
        RECT 63.000 28.200 63.300 30.800 ;
        RECT 63.000 27.800 63.400 28.200 ;
        RECT 85.400 28.100 85.800 28.200 ;
        RECT 86.200 28.100 86.500 136.800 ;
        RECT 87.000 125.800 87.400 126.200 ;
        RECT 87.000 99.200 87.300 125.800 ;
        RECT 87.800 116.200 88.100 139.800 ;
        RECT 88.600 121.200 88.900 157.800 ;
        RECT 89.400 154.800 89.800 155.200 ;
        RECT 89.400 126.200 89.700 154.800 ;
        RECT 90.200 137.200 90.500 201.800 ;
        RECT 110.200 187.800 110.600 188.200 ;
        RECT 93.400 185.800 93.800 186.200 ;
        RECT 91.800 151.800 92.200 152.200 ;
        RECT 90.200 136.800 90.600 137.200 ;
        RECT 89.400 125.800 89.800 126.200 ;
        RECT 88.600 120.800 89.000 121.200 ;
        RECT 87.800 115.800 88.200 116.200 ;
        RECT 91.800 112.200 92.100 151.800 ;
        RECT 93.400 146.200 93.700 185.800 ;
        RECT 97.400 182.800 97.800 183.200 ;
        RECT 95.000 166.100 95.400 166.200 ;
        RECT 95.800 166.100 96.200 166.200 ;
        RECT 95.000 165.800 96.200 166.100 ;
        RECT 97.400 146.200 97.700 182.800 ;
        RECT 103.000 173.100 103.400 173.200 ;
        RECT 103.800 173.100 104.200 173.200 ;
        RECT 103.000 172.800 104.200 173.100 ;
        RECT 104.600 169.800 105.000 170.200 ;
        RECT 104.600 167.200 104.900 169.800 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 99.800 165.800 100.200 166.200 ;
        RECT 100.600 165.800 101.000 166.200 ;
        RECT 93.400 146.100 93.800 146.200 ;
        RECT 92.600 145.800 93.800 146.100 ;
        RECT 97.400 146.100 97.800 146.200 ;
        RECT 98.200 146.100 98.600 146.200 ;
        RECT 97.400 145.800 98.600 146.100 ;
        RECT 92.600 121.200 92.900 145.800 ;
        RECT 99.800 142.200 100.100 165.800 ;
        RECT 100.600 145.200 100.900 165.800 ;
        RECT 103.800 160.800 104.200 161.200 ;
        RECT 103.800 148.200 104.100 160.800 ;
        RECT 109.400 154.100 109.800 154.200 ;
        RECT 110.200 154.100 110.500 187.800 ;
        RECT 111.000 175.200 111.300 220.800 ;
        RECT 111.800 219.800 112.200 220.200 ;
        RECT 111.000 174.800 111.400 175.200 ;
        RECT 109.400 153.800 110.500 154.100 ;
        RECT 103.800 147.800 104.200 148.200 ;
        RECT 101.400 145.800 101.800 146.200 ;
        RECT 100.600 144.800 101.000 145.200 ;
        RECT 99.800 141.800 100.200 142.200 ;
        RECT 101.400 136.200 101.700 145.800 ;
        RECT 102.200 140.800 102.600 141.200 ;
        RECT 101.400 135.800 101.800 136.200 ;
        RECT 101.400 135.200 101.700 135.800 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 102.200 129.200 102.500 140.800 ;
        RECT 103.800 133.200 104.100 147.800 ;
        RECT 109.400 147.200 109.700 153.800 ;
        RECT 109.400 146.800 109.800 147.200 ;
        RECT 107.800 143.800 108.200 144.200 ;
        RECT 105.400 137.100 105.800 137.200 ;
        RECT 104.600 136.800 105.800 137.100 ;
        RECT 104.600 134.200 104.900 136.800 ;
        RECT 104.600 133.800 105.000 134.200 ;
        RECT 103.800 132.800 104.200 133.200 ;
        RECT 106.200 133.100 106.600 133.200 ;
        RECT 107.000 133.100 107.400 133.200 ;
        RECT 106.200 132.800 107.400 133.100 ;
        RECT 103.000 129.800 103.400 130.200 ;
        RECT 102.200 128.800 102.600 129.200 ;
        RECT 92.600 120.800 93.000 121.200 ;
        RECT 91.800 111.800 92.200 112.200 ;
        RECT 92.600 111.800 93.000 112.200 ;
        RECT 88.600 105.800 89.000 106.200 ;
        RECT 88.600 105.100 88.900 105.800 ;
        RECT 89.400 105.100 89.800 105.200 ;
        RECT 88.600 104.800 89.800 105.100 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 91.800 95.200 92.100 111.800 ;
        RECT 92.600 110.200 92.900 111.800 ;
        RECT 92.600 109.800 93.000 110.200 ;
        RECT 94.200 102.800 94.600 103.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 89.400 91.800 89.800 92.200 ;
        RECT 88.600 73.100 89.000 73.200 ;
        RECT 89.400 73.100 89.700 91.800 ;
        RECT 88.600 72.800 89.700 73.100 ;
        RECT 90.200 80.800 90.600 81.200 ;
        RECT 90.200 66.200 90.500 80.800 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 93.400 65.800 93.800 66.200 ;
        RECT 91.000 64.800 91.400 65.200 ;
        RECT 89.400 61.800 89.800 62.200 ;
        RECT 89.400 55.200 89.700 61.800 ;
        RECT 89.400 55.100 89.800 55.200 ;
        RECT 90.200 55.100 90.600 55.200 ;
        RECT 89.400 54.800 90.600 55.100 ;
        RECT 91.000 47.200 91.300 64.800 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 85.400 27.800 86.500 28.100 ;
        RECT 88.600 37.800 89.000 38.200 ;
        RECT 89.400 37.800 89.800 38.200 ;
        RECT 54.200 27.100 54.600 27.200 ;
        RECT 55.000 27.100 55.400 27.200 ;
        RECT 54.200 26.800 55.400 27.100 ;
        RECT 73.400 25.800 73.800 26.200 ;
        RECT 73.400 18.200 73.700 25.800 ;
        RECT 83.800 25.100 84.200 25.200 ;
        RECT 83.800 24.800 84.900 25.100 ;
        RECT 73.400 17.800 73.800 18.200 ;
        RECT 73.400 15.200 73.700 17.800 ;
        RECT 62.200 14.800 62.600 15.200 ;
        RECT 73.400 14.800 73.800 15.200 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 62.200 5.200 62.500 14.800 ;
        RECT 84.600 9.200 84.900 24.800 ;
        RECT 88.600 23.200 88.900 37.800 ;
        RECT 89.400 35.200 89.700 37.800 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 91.800 34.200 92.100 65.800 ;
        RECT 91.800 33.800 92.200 34.200 ;
        RECT 88.600 22.800 89.000 23.200 ;
        RECT 91.800 18.200 92.100 33.800 ;
        RECT 91.800 17.800 92.200 18.200 ;
        RECT 92.600 15.800 93.000 16.200 ;
        RECT 93.400 16.100 93.700 65.800 ;
        RECT 94.200 55.200 94.500 102.800 ;
        RECT 103.000 86.200 103.300 129.800 ;
        RECT 103.800 102.200 104.100 132.800 ;
        RECT 107.800 131.200 108.100 143.800 ;
        RECT 110.200 135.800 110.600 136.200 ;
        RECT 108.600 134.800 109.000 135.200 ;
        RECT 107.800 130.800 108.200 131.200 ;
        RECT 104.600 126.800 105.000 127.200 ;
        RECT 104.600 125.200 104.900 126.800 ;
        RECT 108.600 125.200 108.900 134.800 ;
        RECT 104.600 124.800 105.000 125.200 ;
        RECT 107.800 124.800 108.200 125.200 ;
        RECT 108.600 125.100 109.000 125.200 ;
        RECT 109.400 125.100 109.800 125.200 ;
        RECT 108.600 124.800 109.800 125.100 ;
        RECT 107.800 124.200 108.100 124.800 ;
        RECT 107.800 123.800 108.200 124.200 ;
        RECT 110.200 123.200 110.500 135.800 ;
        RECT 111.800 135.200 112.100 219.800 ;
        RECT 115.000 216.100 115.400 216.200 ;
        RECT 114.200 215.800 115.400 216.100 ;
        RECT 112.600 195.800 113.000 196.200 ;
        RECT 112.600 149.200 112.900 195.800 ;
        RECT 114.200 185.200 114.500 215.800 ;
        RECT 117.400 206.200 117.700 224.800 ;
        RECT 121.400 221.800 121.800 222.200 ;
        RECT 118.200 211.800 118.600 212.200 ;
        RECT 117.400 205.800 117.800 206.200 ;
        RECT 116.600 204.800 117.000 205.200 ;
        RECT 114.200 184.800 114.600 185.200 ;
        RECT 115.800 172.800 116.200 173.200 ;
        RECT 112.600 148.800 113.000 149.200 ;
        RECT 112.600 145.800 113.000 146.200 ;
        RECT 112.600 145.200 112.900 145.800 ;
        RECT 112.600 144.800 113.000 145.200 ;
        RECT 111.800 134.800 112.200 135.200 ;
        RECT 115.800 133.200 116.100 172.800 ;
        RECT 115.800 132.800 116.200 133.200 ;
        RECT 111.000 127.100 111.400 127.200 ;
        RECT 111.800 127.100 112.200 127.200 ;
        RECT 111.000 126.800 112.200 127.100 ;
        RECT 116.600 124.200 116.900 204.800 ;
        RECT 118.200 175.100 118.500 211.800 ;
        RECT 119.000 175.100 119.400 175.200 ;
        RECT 118.200 174.800 119.400 175.100 ;
        RECT 121.400 174.200 121.700 221.800 ;
        RECT 127.800 221.100 128.200 221.200 ;
        RECT 127.000 220.800 128.200 221.100 ;
        RECT 126.200 185.800 126.600 186.200 ;
        RECT 121.400 173.800 121.800 174.200 ;
        RECT 121.400 169.200 121.700 173.800 ;
        RECT 120.600 168.800 121.000 169.200 ;
        RECT 121.400 168.800 121.800 169.200 ;
        RECT 119.000 168.100 119.400 168.200 ;
        RECT 119.800 168.100 120.200 168.200 ;
        RECT 119.000 167.800 120.200 168.100 ;
        RECT 120.600 143.200 120.900 168.800 ;
        RECT 122.200 164.800 122.600 165.200 ;
        RECT 122.200 144.200 122.500 164.800 ;
        RECT 126.200 148.200 126.500 185.800 ;
        RECT 127.000 171.200 127.300 220.800 ;
        RECT 127.000 170.800 127.400 171.200 ;
        RECT 127.000 166.800 127.400 167.200 ;
        RECT 127.000 156.100 127.300 166.800 ;
        RECT 127.800 156.100 128.200 156.200 ;
        RECT 127.000 155.800 128.200 156.100 ;
        RECT 129.400 154.200 129.700 229.800 ;
        RECT 141.400 226.800 141.800 227.200 ;
        RECT 173.400 226.800 173.800 227.200 ;
        RECT 131.800 225.800 132.200 226.200 ;
        RECT 130.200 212.800 130.600 213.200 ;
        RECT 130.200 194.200 130.500 212.800 ;
        RECT 131.800 202.200 132.100 225.800 ;
        RECT 135.000 224.800 135.400 225.200 ;
        RECT 135.000 215.200 135.300 224.800 ;
        RECT 135.800 223.800 136.200 224.200 ;
        RECT 135.000 214.800 135.400 215.200 ;
        RECT 131.800 201.800 132.200 202.200 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 130.200 193.800 130.600 194.200 ;
        RECT 130.200 188.200 130.500 193.800 ;
        RECT 130.200 187.800 130.600 188.200 ;
        RECT 129.400 153.800 129.800 154.200 ;
        RECT 126.200 147.800 126.600 148.200 ;
        RECT 128.600 147.800 129.000 148.200 ;
        RECT 123.800 145.800 124.200 146.200 ;
        RECT 121.400 143.800 121.800 144.200 ;
        RECT 122.200 143.800 122.600 144.200 ;
        RECT 120.600 142.800 121.000 143.200 ;
        RECT 119.800 136.800 120.200 137.200 ;
        RECT 119.800 135.200 120.100 136.800 ;
        RECT 119.800 134.800 120.200 135.200 ;
        RECT 117.400 126.800 117.800 127.200 ;
        RECT 117.400 126.200 117.700 126.800 ;
        RECT 117.400 125.800 117.800 126.200 ;
        RECT 119.000 125.100 119.400 125.200 ;
        RECT 119.800 125.100 120.200 125.200 ;
        RECT 119.000 124.800 120.200 125.100 ;
        RECT 116.600 123.800 117.000 124.200 ;
        RECT 110.200 122.800 110.600 123.200 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 103.800 101.800 104.200 102.200 ;
        RECT 103.800 92.200 104.100 101.800 ;
        RECT 103.800 91.800 104.200 92.200 ;
        RECT 103.000 85.800 103.400 86.200 ;
        RECT 111.800 84.800 112.200 85.200 ;
        RECT 110.200 80.800 110.600 81.200 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 107.000 75.100 107.400 75.200 ;
        RECT 106.200 74.800 107.400 75.100 ;
        RECT 109.400 72.800 109.800 73.200 ;
        RECT 109.400 71.200 109.700 72.800 ;
        RECT 109.400 70.800 109.800 71.200 ;
        RECT 95.000 69.800 95.400 70.200 ;
        RECT 108.600 69.800 109.000 70.200 ;
        RECT 94.200 54.800 94.600 55.200 ;
        RECT 95.000 27.200 95.300 69.800 ;
        RECT 96.600 67.800 97.000 68.200 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 95.800 42.200 96.100 66.800 ;
        RECT 96.600 66.200 96.900 67.800 ;
        RECT 96.600 65.800 97.000 66.200 ;
        RECT 103.800 64.800 104.200 65.200 ;
        RECT 102.200 56.800 102.600 57.200 ;
        RECT 95.800 41.800 96.200 42.200 ;
        RECT 102.200 35.200 102.500 56.800 ;
        RECT 103.800 41.200 104.100 64.800 ;
        RECT 108.600 43.200 108.900 69.800 ;
        RECT 108.600 42.800 109.000 43.200 ;
        RECT 103.800 40.800 104.200 41.200 ;
        RECT 110.200 37.100 110.500 80.800 ;
        RECT 111.800 67.200 112.100 84.800 ;
        RECT 112.600 74.800 113.000 75.200 ;
        RECT 112.600 74.200 112.900 74.800 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 111.800 66.800 112.200 67.200 ;
        RECT 113.400 63.200 113.700 107.800 ;
        RECT 121.400 90.200 121.700 143.800 ;
        RECT 121.400 89.800 121.800 90.200 ;
        RECT 123.800 86.200 124.100 145.800 ;
        RECT 125.400 122.800 125.800 123.200 ;
        RECT 124.600 116.800 125.000 117.200 ;
        RECT 124.600 111.200 124.900 116.800 ;
        RECT 124.600 110.800 125.000 111.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 120.600 67.100 121.000 67.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 120.600 66.800 121.800 67.100 ;
        RECT 122.200 66.800 122.600 67.200 ;
        RECT 113.400 62.800 113.800 63.200 ;
        RECT 111.000 37.100 111.400 37.200 ;
        RECT 110.200 36.800 111.400 37.100 ;
        RECT 102.200 34.800 102.600 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 106.200 35.100 106.600 35.200 ;
        RECT 105.400 34.800 106.600 35.100 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 94.200 16.100 94.600 16.200 ;
        RECT 93.400 15.800 94.600 16.100 ;
        RECT 92.600 15.200 92.900 15.800 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 84.600 8.800 85.000 9.200 ;
        RECT 94.200 6.200 94.500 15.800 ;
        RECT 95.000 14.200 95.300 26.800 ;
        RECT 97.400 19.100 97.800 19.200 ;
        RECT 96.600 18.800 97.800 19.100 ;
        RECT 95.000 13.800 95.400 14.200 ;
        RECT 96.600 8.200 96.900 18.800 ;
        RECT 99.000 15.100 99.400 15.200 ;
        RECT 99.800 15.100 100.200 15.200 ;
        RECT 99.000 14.800 100.200 15.100 ;
        RECT 96.600 7.800 97.000 8.200 ;
        RECT 113.400 6.200 113.700 62.800 ;
        RECT 115.000 54.800 115.400 55.200 ;
        RECT 115.000 54.200 115.300 54.800 ;
        RECT 115.000 53.800 115.400 54.200 ;
        RECT 122.200 39.200 122.500 66.800 ;
        RECT 123.800 66.200 124.100 85.800 ;
        RECT 125.400 77.200 125.700 122.800 ;
        RECT 128.600 95.200 128.900 147.800 ;
        RECT 131.000 136.200 131.300 194.800 ;
        RECT 132.600 192.800 133.000 193.200 ;
        RECT 131.800 158.800 132.200 159.200 ;
        RECT 131.800 151.200 132.100 158.800 ;
        RECT 131.800 150.800 132.200 151.200 ;
        RECT 131.000 135.800 131.400 136.200 ;
        RECT 130.200 114.800 130.600 115.200 ;
        RECT 128.600 94.800 129.000 95.200 ;
        RECT 125.400 76.800 125.800 77.200 ;
        RECT 125.400 66.200 125.700 76.800 ;
        RECT 127.800 75.800 128.200 76.200 ;
        RECT 127.800 75.200 128.100 75.800 ;
        RECT 127.800 74.800 128.200 75.200 ;
        RECT 130.200 72.200 130.500 114.800 ;
        RECT 131.000 94.800 131.400 95.200 ;
        RECT 130.200 71.800 130.600 72.200 ;
        RECT 127.800 68.800 128.200 69.200 ;
        RECT 123.800 65.800 124.200 66.200 ;
        RECT 124.600 65.800 125.000 66.200 ;
        RECT 125.400 65.800 125.800 66.200 ;
        RECT 124.600 65.200 124.900 65.800 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 127.800 51.200 128.100 68.800 ;
        RECT 128.600 68.100 129.000 68.200 ;
        RECT 129.400 68.100 129.800 68.200 ;
        RECT 128.600 67.800 129.800 68.100 ;
        RECT 130.200 56.200 130.500 71.800 ;
        RECT 130.200 55.800 130.600 56.200 ;
        RECT 127.800 50.800 128.200 51.200 ;
        RECT 129.400 49.800 129.800 50.200 ;
        RECT 129.400 48.200 129.700 49.800 ;
        RECT 129.400 47.800 129.800 48.200 ;
        RECT 131.000 47.200 131.300 94.800 ;
        RECT 131.800 48.200 132.100 150.800 ;
        RECT 132.600 140.200 132.900 192.800 ;
        RECT 135.000 160.200 135.300 214.800 ;
        RECT 135.000 159.800 135.400 160.200 ;
        RECT 135.800 155.200 136.100 223.800 ;
        RECT 141.400 208.200 141.700 226.800 ;
        RECT 173.400 226.200 173.700 226.800 ;
        RECT 173.400 225.800 173.800 226.200 ;
        RECT 211.800 221.800 212.200 222.200 ;
        RECT 179.000 216.800 179.400 217.200 ;
        RECT 170.200 211.800 170.600 212.200 ;
        RECT 141.400 207.800 141.800 208.200 ;
        RECT 158.200 207.800 158.600 208.200 ;
        RECT 144.600 204.800 145.000 205.200 ;
        RECT 144.600 196.200 144.900 204.800 ;
        RECT 154.200 201.800 154.600 202.200 ;
        RECT 144.600 195.800 145.000 196.200 ;
        RECT 139.800 184.800 140.200 185.200 ;
        RECT 136.600 172.800 137.000 173.200 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 132.600 139.800 133.000 140.200 ;
        RECT 132.600 134.800 133.000 135.200 ;
        RECT 132.600 127.200 132.900 134.800 ;
        RECT 132.600 126.800 133.000 127.200 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 135.000 122.200 135.300 124.800 ;
        RECT 135.000 121.800 135.400 122.200 ;
        RECT 134.200 116.800 134.600 117.200 ;
        RECT 134.200 106.200 134.500 116.800 ;
        RECT 136.600 107.200 136.900 172.800 ;
        RECT 139.800 140.200 140.100 184.800 ;
        RECT 141.400 181.800 141.800 182.200 ;
        RECT 142.200 181.800 142.600 182.200 ;
        RECT 140.600 164.800 141.000 165.200 ;
        RECT 140.600 142.200 140.900 164.800 ;
        RECT 141.400 153.200 141.700 181.800 ;
        RECT 142.200 181.200 142.500 181.800 ;
        RECT 142.200 180.800 142.600 181.200 ;
        RECT 142.200 164.200 142.500 180.800 ;
        RECT 142.200 163.800 142.600 164.200 ;
        RECT 142.200 155.200 142.500 163.800 ;
        RECT 143.000 163.100 143.400 163.200 ;
        RECT 143.800 163.100 144.200 163.200 ;
        RECT 143.000 162.800 144.200 163.100 ;
        RECT 142.200 154.800 142.600 155.200 ;
        RECT 142.200 153.800 142.600 154.200 ;
        RECT 141.400 152.800 141.800 153.200 ;
        RECT 140.600 141.800 141.000 142.200 ;
        RECT 139.800 139.800 140.200 140.200 ;
        RECT 137.400 137.800 137.800 138.200 ;
        RECT 136.600 106.800 137.000 107.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 132.600 78.800 133.000 79.200 ;
        RECT 132.600 49.200 132.900 78.800 ;
        RECT 134.200 70.200 134.500 105.800 ;
        RECT 134.200 69.800 134.600 70.200 ;
        RECT 133.400 66.800 133.800 67.200 ;
        RECT 133.400 66.200 133.700 66.800 ;
        RECT 133.400 65.800 133.800 66.200 ;
        RECT 132.600 48.800 133.000 49.200 ;
        RECT 131.800 47.800 132.200 48.200 ;
        RECT 131.000 46.800 131.400 47.200 ;
        RECT 122.200 38.800 122.600 39.200 ;
        RECT 134.200 36.200 134.500 69.800 ;
        RECT 136.600 66.800 137.000 67.200 ;
        RECT 136.600 66.200 136.900 66.800 ;
        RECT 137.400 66.200 137.700 137.800 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 139.000 134.100 139.400 134.200 ;
        RECT 138.200 133.800 139.400 134.100 ;
        RECT 139.800 116.200 140.100 139.800 ;
        RECT 139.800 115.800 140.200 116.200 ;
        RECT 142.200 113.200 142.500 153.800 ;
        RECT 143.800 152.800 144.200 153.200 ;
        RECT 143.000 151.800 143.400 152.200 ;
        RECT 143.000 146.200 143.300 151.800 ;
        RECT 143.000 145.800 143.400 146.200 ;
        RECT 143.000 143.800 143.400 144.200 ;
        RECT 143.000 124.200 143.300 143.800 ;
        RECT 143.800 134.200 144.100 152.800 ;
        RECT 144.600 151.200 144.900 195.800 ;
        RECT 151.800 183.800 152.200 184.200 ;
        RECT 151.800 183.200 152.100 183.800 ;
        RECT 151.800 183.100 152.200 183.200 ;
        RECT 151.000 182.800 152.200 183.100 ;
        RECT 147.800 174.100 148.200 174.200 ;
        RECT 147.800 173.800 148.900 174.100 ;
        RECT 147.000 166.100 147.400 166.200 ;
        RECT 147.800 166.100 148.200 166.200 ;
        RECT 147.000 165.800 148.200 166.100 ;
        RECT 148.600 165.200 148.900 173.800 ;
        RECT 151.000 165.200 151.300 182.800 ;
        RECT 148.600 164.800 149.000 165.200 ;
        RECT 151.000 164.800 151.400 165.200 ;
        RECT 145.400 161.800 145.800 162.200 ;
        RECT 145.400 151.200 145.700 161.800 ;
        RECT 149.400 155.800 149.800 156.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 147.000 153.800 147.400 154.200 ;
        RECT 144.600 150.800 145.000 151.200 ;
        RECT 145.400 150.800 145.800 151.200 ;
        RECT 147.000 148.200 147.300 153.800 ;
        RECT 147.000 147.800 147.400 148.200 ;
        RECT 146.200 143.800 146.600 144.200 ;
        RECT 146.200 141.200 146.500 143.800 ;
        RECT 146.200 140.800 146.600 141.200 ;
        RECT 146.200 139.800 146.600 140.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 144.600 134.100 145.000 134.200 ;
        RECT 145.400 134.100 145.800 134.200 ;
        RECT 144.600 133.800 145.800 134.100 ;
        RECT 144.600 125.800 145.000 126.200 ;
        RECT 144.600 125.200 144.900 125.800 ;
        RECT 144.600 124.800 145.000 125.200 ;
        RECT 143.000 123.800 143.400 124.200 ;
        RECT 144.600 123.800 145.000 124.200 ;
        RECT 143.000 119.200 143.300 123.800 ;
        RECT 143.000 118.800 143.400 119.200 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 141.400 106.800 141.800 107.200 ;
        RECT 140.600 86.800 141.000 87.200 ;
        RECT 140.600 69.200 140.900 86.800 ;
        RECT 141.400 75.200 141.700 106.800 ;
        RECT 142.200 95.800 142.600 96.200 ;
        RECT 142.200 94.200 142.500 95.800 ;
        RECT 142.200 93.800 142.600 94.200 ;
        RECT 142.200 75.800 142.600 76.200 ;
        RECT 142.200 75.200 142.500 75.800 ;
        RECT 141.400 74.800 141.800 75.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 140.600 68.800 141.000 69.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 135.800 64.800 136.200 65.200 ;
        RECT 135.800 54.200 136.100 64.800 ;
        RECT 137.400 64.200 137.700 65.800 ;
        RECT 137.400 63.800 137.800 64.200 ;
        RECT 137.400 62.200 137.700 63.800 ;
        RECT 137.400 61.800 137.800 62.200 ;
        RECT 139.800 59.800 140.200 60.200 ;
        RECT 135.800 53.800 136.200 54.200 ;
        RECT 134.200 35.800 134.600 36.200 ;
        RECT 139.800 35.200 140.100 59.800 ;
        RECT 142.200 55.200 142.500 74.800 ;
        RECT 143.000 58.800 143.400 59.200 ;
        RECT 143.000 55.200 143.300 58.800 ;
        RECT 142.200 54.800 142.600 55.200 ;
        RECT 143.000 54.800 143.400 55.200 ;
        RECT 143.800 46.200 144.100 112.800 ;
        RECT 144.600 108.200 144.900 123.800 ;
        RECT 146.200 118.200 146.500 139.800 ;
        RECT 147.800 126.200 148.100 154.800 ;
        RECT 148.600 141.800 149.000 142.200 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 147.800 118.800 148.200 119.200 ;
        RECT 146.200 117.800 146.600 118.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 144.600 107.800 145.000 108.200 ;
        RECT 146.200 63.800 146.600 64.200 ;
        RECT 146.200 52.200 146.500 63.800 ;
        RECT 146.200 51.800 146.600 52.200 ;
        RECT 143.800 45.800 144.200 46.200 ;
        RECT 139.800 34.800 140.200 35.200 ;
        RECT 124.600 31.800 125.000 32.200 ;
        RECT 118.200 27.800 118.600 28.200 ;
        RECT 117.400 27.100 117.800 27.200 ;
        RECT 118.200 27.100 118.500 27.800 ;
        RECT 117.400 26.800 118.500 27.100 ;
        RECT 124.600 24.200 124.900 31.800 ;
        RECT 147.000 26.200 147.300 113.800 ;
        RECT 147.800 87.200 148.100 118.800 ;
        RECT 148.600 116.200 148.900 141.800 ;
        RECT 148.600 115.800 149.000 116.200 ;
        RECT 148.600 114.800 149.000 115.200 ;
        RECT 148.600 114.200 148.900 114.800 ;
        RECT 148.600 113.800 149.000 114.200 ;
        RECT 147.800 86.800 148.200 87.200 ;
        RECT 149.400 66.200 149.700 155.800 ;
        RECT 152.600 135.800 153.000 136.200 ;
        RECT 152.600 116.200 152.900 135.800 ;
        RECT 154.200 133.200 154.500 201.800 ;
        RECT 155.000 194.800 155.400 195.200 ;
        RECT 155.000 151.200 155.300 194.800 ;
        RECT 156.600 156.800 157.000 157.200 ;
        RECT 156.600 155.200 156.900 156.800 ;
        RECT 156.600 154.800 157.000 155.200 ;
        RECT 155.000 150.800 155.400 151.200 ;
        RECT 155.000 140.800 155.400 141.200 ;
        RECT 155.000 134.200 155.300 140.800 ;
        RECT 158.200 139.200 158.500 207.800 ;
        RECT 163.000 204.800 163.400 205.200 ;
        RECT 159.000 190.800 159.400 191.200 ;
        RECT 159.000 166.200 159.300 190.800 ;
        RECT 159.800 167.800 160.200 168.200 ;
        RECT 159.000 165.800 159.400 166.200 ;
        RECT 158.200 138.800 158.600 139.200 ;
        RECT 155.000 133.800 155.400 134.200 ;
        RECT 154.200 132.800 154.600 133.200 ;
        RECT 152.600 115.800 153.000 116.200 ;
        RECT 150.200 67.800 150.600 68.200 ;
        RECT 150.200 67.200 150.500 67.800 ;
        RECT 150.200 66.800 150.600 67.200 ;
        RECT 149.400 65.800 149.800 66.200 ;
        RECT 152.600 57.200 152.900 115.800 ;
        RECT 155.000 107.200 155.300 133.800 ;
        RECT 159.800 127.200 160.100 167.800 ;
        RECT 162.200 150.800 162.600 151.200 ;
        RECT 160.600 148.800 161.000 149.200 ;
        RECT 160.600 145.200 160.900 148.800 ;
        RECT 160.600 144.800 161.000 145.200 ;
        RECT 161.400 132.800 161.800 133.200 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 159.000 115.800 159.400 116.200 ;
        RECT 155.000 106.800 155.400 107.200 ;
        RECT 153.400 106.100 153.800 106.200 ;
        RECT 154.200 106.100 154.600 106.200 ;
        RECT 153.400 105.800 154.600 106.100 ;
        RECT 155.000 76.200 155.300 106.800 ;
        RECT 156.600 77.100 157.000 77.200 ;
        RECT 157.400 77.100 157.800 77.200 ;
        RECT 156.600 76.800 157.800 77.100 ;
        RECT 155.000 75.800 155.400 76.200 ;
        RECT 152.600 56.800 153.000 57.200 ;
        RECT 159.000 54.200 159.300 115.800 ;
        RECT 159.800 108.100 160.200 108.200 ;
        RECT 160.600 108.100 161.000 108.200 ;
        RECT 159.800 107.800 161.000 108.100 ;
        RECT 161.400 99.200 161.700 132.800 ;
        RECT 161.400 98.800 161.800 99.200 ;
        RECT 162.200 85.200 162.500 150.800 ;
        RECT 163.000 144.200 163.300 204.800 ;
        RECT 166.200 193.800 166.600 194.200 ;
        RECT 166.200 166.200 166.500 193.800 ;
        RECT 167.000 189.800 167.400 190.200 ;
        RECT 167.000 187.200 167.300 189.800 ;
        RECT 167.000 186.800 167.400 187.200 ;
        RECT 169.400 176.800 169.800 177.200 ;
        RECT 167.800 172.800 168.200 173.200 ;
        RECT 167.000 168.800 167.400 169.200 ;
        RECT 163.800 165.800 164.200 166.200 ;
        RECT 166.200 165.800 166.600 166.200 ;
        RECT 163.000 143.800 163.400 144.200 ;
        RECT 163.800 133.200 164.100 165.800 ;
        RECT 165.400 133.800 165.800 134.200 ;
        RECT 163.800 132.800 164.200 133.200 ;
        RECT 164.600 132.800 165.000 133.200 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 160.600 84.800 161.000 85.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 160.600 78.200 160.900 84.800 ;
        RECT 163.000 84.200 163.300 106.800 ;
        RECT 164.600 104.200 164.900 132.800 ;
        RECT 165.400 107.200 165.700 133.800 ;
        RECT 166.200 123.200 166.500 165.800 ;
        RECT 167.000 152.200 167.300 168.800 ;
        RECT 167.000 151.800 167.400 152.200 ;
        RECT 167.000 149.800 167.400 150.200 ;
        RECT 167.000 134.200 167.300 149.800 ;
        RECT 167.000 133.800 167.400 134.200 ;
        RECT 167.800 126.200 168.100 172.800 ;
        RECT 169.400 166.200 169.700 176.800 ;
        RECT 169.400 165.800 169.800 166.200 ;
        RECT 168.600 164.800 169.000 165.200 ;
        RECT 168.600 159.200 168.900 164.800 ;
        RECT 168.600 158.800 169.000 159.200 ;
        RECT 168.600 151.200 168.900 158.800 ;
        RECT 170.200 157.200 170.500 211.800 ;
        RECT 173.400 188.800 173.800 189.200 ;
        RECT 173.400 171.200 173.700 188.800 ;
        RECT 179.000 188.100 179.300 216.800 ;
        RECT 182.200 213.800 182.600 214.200 ;
        RECT 199.800 213.800 200.200 214.200 ;
        RECT 179.800 188.100 180.200 188.200 ;
        RECT 179.000 187.800 180.200 188.100 ;
        RECT 178.200 175.800 178.600 176.200 ;
        RECT 173.400 170.800 173.800 171.200 ;
        RECT 171.800 165.800 172.200 166.200 ;
        RECT 176.600 165.800 177.000 166.200 ;
        RECT 171.800 165.200 172.100 165.800 ;
        RECT 171.800 164.800 172.200 165.200 ;
        RECT 175.000 165.100 175.400 165.200 ;
        RECT 175.800 165.100 176.200 165.200 ;
        RECT 175.000 164.800 176.200 165.100 ;
        RECT 171.800 157.200 172.100 164.800 ;
        RECT 176.600 160.200 176.900 165.800 ;
        RECT 176.600 159.800 177.000 160.200 ;
        RECT 170.200 156.800 170.600 157.200 ;
        RECT 171.800 156.800 172.200 157.200 ;
        RECT 169.400 155.100 169.800 155.200 ;
        RECT 170.200 155.100 170.600 155.200 ;
        RECT 169.400 154.800 170.600 155.100 ;
        RECT 175.000 155.100 175.400 155.200 ;
        RECT 175.800 155.100 176.200 155.200 ;
        RECT 175.000 154.800 176.200 155.100 ;
        RECT 169.400 154.100 169.800 154.200 ;
        RECT 170.200 154.100 170.600 154.200 ;
        RECT 169.400 153.800 170.600 154.100 ;
        RECT 168.600 150.800 169.000 151.200 ;
        RECT 175.000 147.200 175.300 154.800 ;
        RECT 176.600 154.200 176.900 159.800 ;
        RECT 176.600 153.800 177.000 154.200 ;
        RECT 175.000 146.800 175.400 147.200 ;
        RECT 168.600 136.100 169.000 136.200 ;
        RECT 169.400 136.100 169.800 136.200 ;
        RECT 168.600 135.800 169.800 136.100 ;
        RECT 176.600 131.200 176.900 153.800 ;
        RECT 178.200 137.200 178.500 175.800 ;
        RECT 181.400 170.800 181.800 171.200 ;
        RECT 180.600 141.800 181.000 142.200 ;
        RECT 180.600 140.200 180.900 141.800 ;
        RECT 180.600 139.800 181.000 140.200 ;
        RECT 179.000 137.800 179.400 138.200 ;
        RECT 179.000 137.200 179.300 137.800 ;
        RECT 178.200 136.800 178.600 137.200 ;
        RECT 179.000 136.800 179.400 137.200 ;
        RECT 180.600 135.800 181.000 136.200 ;
        RECT 176.600 130.800 177.000 131.200 ;
        RECT 171.800 128.800 172.200 129.200 ;
        RECT 171.800 126.200 172.100 128.800 ;
        RECT 167.800 125.800 168.200 126.200 ;
        RECT 171.800 125.800 172.200 126.200 ;
        RECT 167.800 125.100 168.200 125.200 ;
        RECT 168.600 125.100 169.000 125.200 ;
        RECT 167.800 124.800 169.000 125.100 ;
        RECT 166.200 122.800 166.600 123.200 ;
        RECT 172.600 110.800 173.000 111.200 ;
        RECT 167.800 107.800 168.200 108.200 ;
        RECT 165.400 106.800 165.800 107.200 ;
        RECT 164.600 103.800 165.000 104.200 ;
        RECT 163.000 83.800 163.400 84.200 ;
        RECT 163.800 81.800 164.200 82.200 ;
        RECT 160.600 77.800 161.000 78.200 ;
        RECT 163.000 75.800 163.400 76.200 ;
        RECT 163.000 74.200 163.300 75.800 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 163.800 59.200 164.100 81.800 ;
        RECT 164.600 80.200 164.900 103.800 ;
        RECT 164.600 79.800 165.000 80.200 ;
        RECT 165.400 71.200 165.700 106.800 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 167.000 106.100 167.400 106.200 ;
        RECT 166.200 105.800 167.400 106.100 ;
        RECT 166.200 73.100 166.600 73.200 ;
        RECT 166.200 72.800 167.300 73.100 ;
        RECT 165.400 70.800 165.800 71.200 ;
        RECT 166.200 70.800 166.600 71.200 ;
        RECT 165.400 66.200 165.700 70.800 ;
        RECT 166.200 67.200 166.500 70.800 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 165.400 65.800 165.800 66.200 ;
        RECT 166.200 65.800 166.600 66.200 ;
        RECT 166.200 64.200 166.500 65.800 ;
        RECT 167.000 65.200 167.300 72.800 ;
        RECT 167.800 67.200 168.100 107.800 ;
        RECT 170.200 100.800 170.600 101.200 ;
        RECT 170.200 72.200 170.500 100.800 ;
        RECT 172.600 86.200 172.900 110.800 ;
        RECT 173.400 109.800 173.800 110.200 ;
        RECT 173.400 89.100 173.700 109.800 ;
        RECT 174.200 89.100 174.600 89.200 ;
        RECT 173.400 88.800 174.600 89.100 ;
        RECT 172.600 85.800 173.000 86.200 ;
        RECT 176.600 74.800 177.000 75.200 ;
        RECT 170.200 71.800 170.600 72.200 ;
        RECT 169.400 67.800 169.800 68.200 ;
        RECT 169.400 67.200 169.700 67.800 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 170.200 66.200 170.500 71.800 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 167.000 64.800 167.400 65.200 ;
        RECT 166.200 63.800 166.600 64.200 ;
        RECT 163.800 58.800 164.200 59.200 ;
        RECT 176.600 55.200 176.900 74.800 ;
        RECT 179.000 71.100 179.400 71.200 ;
        RECT 179.800 71.100 180.200 71.200 ;
        RECT 179.000 70.800 180.200 71.100 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 159.000 53.800 159.400 54.200 ;
        RECT 159.000 46.200 159.300 53.800 ;
        RECT 159.000 45.800 159.400 46.200 ;
        RECT 167.800 37.800 168.200 38.200 ;
        RECT 167.000 35.800 167.400 36.200 ;
        RECT 166.200 35.100 166.600 35.200 ;
        RECT 167.000 35.100 167.300 35.800 ;
        RECT 166.200 34.800 167.300 35.100 ;
        RECT 160.600 32.800 161.000 33.200 ;
        RECT 160.600 28.200 160.900 32.800 ;
        RECT 160.600 27.800 161.000 28.200 ;
        RECT 167.800 27.200 168.100 37.800 ;
        RECT 175.000 33.800 175.400 34.200 ;
        RECT 172.600 28.800 173.000 29.200 ;
        RECT 172.600 27.200 172.900 28.800 ;
        RECT 167.800 26.800 168.200 27.200 ;
        RECT 172.600 26.800 173.000 27.200 ;
        RECT 175.000 26.200 175.300 33.800 ;
        RECT 147.000 25.800 147.400 26.200 ;
        RECT 175.000 25.800 175.400 26.200 ;
        RECT 124.600 23.800 125.000 24.200 ;
        RECT 159.000 18.100 159.400 18.200 ;
        RECT 159.800 18.100 160.200 18.200 ;
        RECT 159.000 17.800 160.200 18.100 ;
        RECT 179.000 13.200 179.300 70.800 ;
        RECT 180.600 42.200 180.900 135.800 ;
        RECT 181.400 95.200 181.700 170.800 ;
        RECT 182.200 146.200 182.500 213.800 ;
        RECT 199.800 187.200 200.100 213.800 ;
        RECT 206.200 211.800 206.600 212.200 ;
        RECT 200.600 205.800 201.000 206.200 ;
        RECT 199.800 186.800 200.200 187.200 ;
        RECT 198.200 184.800 198.600 185.200 ;
        RECT 198.200 184.200 198.500 184.800 ;
        RECT 198.200 183.800 198.600 184.200 ;
        RECT 197.400 177.800 197.800 178.200 ;
        RECT 191.800 173.800 192.200 174.200 ;
        RECT 187.000 167.800 187.400 168.200 ;
        RECT 187.000 166.200 187.300 167.800 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 190.200 165.800 190.600 166.200 ;
        RECT 190.200 162.200 190.500 165.800 ;
        RECT 190.200 161.800 190.600 162.200 ;
        RECT 187.000 156.800 187.400 157.200 ;
        RECT 182.200 145.800 182.600 146.200 ;
        RECT 182.200 139.800 182.600 140.200 ;
        RECT 182.200 136.200 182.500 139.800 ;
        RECT 182.200 135.800 182.600 136.200 ;
        RECT 187.000 135.200 187.300 156.800 ;
        RECT 187.800 144.800 188.200 145.200 ;
        RECT 187.000 134.800 187.400 135.200 ;
        RECT 187.000 104.200 187.300 134.800 ;
        RECT 182.200 103.800 182.600 104.200 ;
        RECT 187.000 103.800 187.400 104.200 ;
        RECT 181.400 94.800 181.800 95.200 ;
        RECT 182.200 81.200 182.500 103.800 ;
        RECT 184.600 102.800 185.000 103.200 ;
        RECT 184.600 92.200 184.900 102.800 ;
        RECT 187.800 92.200 188.100 144.800 ;
        RECT 191.800 117.200 192.100 173.800 ;
        RECT 192.600 169.100 193.000 169.200 ;
        RECT 193.400 169.100 193.800 169.200 ;
        RECT 192.600 168.800 193.800 169.100 ;
        RECT 194.200 165.800 194.600 166.200 ;
        RECT 195.800 165.800 196.200 166.200 ;
        RECT 194.200 163.200 194.500 165.800 ;
        RECT 195.800 165.200 196.100 165.800 ;
        RECT 195.800 164.800 196.200 165.200 ;
        RECT 194.200 162.800 194.600 163.200 ;
        RECT 195.800 157.100 196.200 157.200 ;
        RECT 196.600 157.100 197.000 157.200 ;
        RECT 195.800 156.800 197.000 157.100 ;
        RECT 197.400 136.200 197.700 177.800 ;
        RECT 199.800 174.800 200.200 175.200 ;
        RECT 199.000 173.800 199.400 174.200 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 199.000 134.200 199.300 173.800 ;
        RECT 199.800 135.200 200.100 174.800 ;
        RECT 200.600 146.200 200.900 205.800 ;
        RECT 206.200 200.200 206.500 211.800 ;
        RECT 211.800 209.200 212.100 221.800 ;
        RECT 211.800 208.800 212.200 209.200 ;
        RECT 211.800 205.800 212.200 206.200 ;
        RECT 210.200 204.800 210.600 205.200 ;
        RECT 206.200 199.800 206.600 200.200 ;
        RECT 203.800 193.800 204.200 194.200 ;
        RECT 203.800 185.200 204.100 193.800 ;
        RECT 203.800 184.800 204.200 185.200 ;
        RECT 202.200 169.800 202.600 170.200 ;
        RECT 201.400 167.800 201.800 168.200 ;
        RECT 201.400 167.200 201.700 167.800 ;
        RECT 201.400 166.800 201.800 167.200 ;
        RECT 200.600 145.800 201.000 146.200 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 199.000 134.100 199.400 134.200 ;
        RECT 199.800 134.100 200.200 134.200 ;
        RECT 199.000 133.800 200.200 134.100 ;
        RECT 194.200 132.800 194.600 133.200 ;
        RECT 193.400 119.800 193.800 120.200 ;
        RECT 191.800 116.800 192.200 117.200 ;
        RECT 184.600 91.800 185.000 92.200 ;
        RECT 187.000 91.800 187.400 92.200 ;
        RECT 187.800 91.800 188.200 92.200 ;
        RECT 183.800 90.800 184.200 91.200 ;
        RECT 182.200 80.800 182.600 81.200 ;
        RECT 182.200 42.200 182.500 80.800 ;
        RECT 183.000 73.800 183.400 74.200 ;
        RECT 183.000 73.200 183.300 73.800 ;
        RECT 183.000 72.800 183.400 73.200 ;
        RECT 180.600 41.800 181.000 42.200 ;
        RECT 182.200 41.800 182.600 42.200 ;
        RECT 180.600 36.200 180.900 41.800 ;
        RECT 180.600 35.800 181.000 36.200 ;
        RECT 183.800 15.200 184.100 90.800 ;
        RECT 187.000 57.200 187.300 91.800 ;
        RECT 188.600 89.800 189.000 90.200 ;
        RECT 188.600 87.100 188.900 89.800 ;
        RECT 189.400 87.100 189.800 87.200 ;
        RECT 188.600 86.800 189.800 87.100 ;
        RECT 188.600 74.100 189.000 74.200 ;
        RECT 189.400 74.100 189.800 74.200 ;
        RECT 188.600 73.800 189.800 74.100 ;
        RECT 193.400 59.200 193.700 119.800 ;
        RECT 194.200 76.200 194.500 132.800 ;
        RECT 196.600 124.800 197.000 125.200 ;
        RECT 195.800 96.800 196.200 97.200 ;
        RECT 194.200 75.800 194.600 76.200 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 187.000 56.800 187.400 57.200 ;
        RECT 187.000 38.200 187.300 56.800 ;
        RECT 187.000 37.800 187.400 38.200 ;
        RECT 188.600 35.100 189.000 35.200 ;
        RECT 188.600 34.800 189.700 35.100 ;
        RECT 189.400 34.200 189.700 34.800 ;
        RECT 189.400 33.800 189.800 34.200 ;
        RECT 193.400 21.200 193.700 58.800 ;
        RECT 194.200 55.200 194.500 75.800 ;
        RECT 195.800 59.200 196.100 96.800 ;
        RECT 196.600 76.200 196.900 124.800 ;
        RECT 199.800 103.200 200.100 133.800 ;
        RECT 199.800 102.800 200.200 103.200 ;
        RECT 200.600 102.200 200.900 145.800 ;
        RECT 202.200 121.200 202.500 169.800 ;
        RECT 206.200 164.800 206.600 165.200 ;
        RECT 203.000 155.100 203.400 155.200 ;
        RECT 203.800 155.100 204.200 155.200 ;
        RECT 203.000 154.800 204.200 155.100 ;
        RECT 203.000 142.800 203.400 143.200 ;
        RECT 202.200 120.800 202.600 121.200 ;
        RECT 200.600 101.800 201.000 102.200 ;
        RECT 199.800 100.800 200.200 101.200 ;
        RECT 197.400 86.800 197.800 87.200 ;
        RECT 197.400 82.200 197.700 86.800 ;
        RECT 197.400 81.800 197.800 82.200 ;
        RECT 196.600 75.800 197.000 76.200 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 198.200 75.100 198.600 75.200 ;
        RECT 197.400 74.800 198.600 75.100 ;
        RECT 199.800 66.200 200.100 100.800 ;
        RECT 196.600 65.800 197.000 66.200 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 196.600 65.200 196.900 65.800 ;
        RECT 196.600 64.800 197.000 65.200 ;
        RECT 195.800 58.800 196.200 59.200 ;
        RECT 194.200 54.800 194.600 55.200 ;
        RECT 202.200 35.200 202.500 120.800 ;
        RECT 203.000 115.200 203.300 142.800 ;
        RECT 203.800 134.800 204.200 135.200 ;
        RECT 203.000 114.800 203.400 115.200 ;
        RECT 203.800 111.200 204.100 134.800 ;
        RECT 206.200 126.200 206.500 164.800 ;
        RECT 207.000 159.800 207.400 160.200 ;
        RECT 207.000 153.200 207.300 159.800 ;
        RECT 207.000 152.800 207.400 153.200 ;
        RECT 207.000 131.200 207.300 152.800 ;
        RECT 207.800 144.800 208.200 145.200 ;
        RECT 207.800 142.200 208.100 144.800 ;
        RECT 207.800 141.800 208.200 142.200 ;
        RECT 207.000 130.800 207.400 131.200 ;
        RECT 210.200 129.200 210.500 204.800 ;
        RECT 211.000 168.800 211.400 169.200 ;
        RECT 211.000 167.200 211.300 168.800 ;
        RECT 211.000 166.800 211.400 167.200 ;
        RECT 211.000 159.800 211.400 160.200 ;
        RECT 211.000 134.200 211.300 159.800 ;
        RECT 211.000 133.800 211.400 134.200 ;
        RECT 210.200 128.800 210.600 129.200 ;
        RECT 205.400 125.800 205.800 126.200 ;
        RECT 206.200 125.800 206.600 126.200 ;
        RECT 205.400 124.200 205.700 125.800 ;
        RECT 205.400 123.800 205.800 124.200 ;
        RECT 210.200 114.800 210.600 115.200 ;
        RECT 210.200 111.200 210.500 114.800 ;
        RECT 203.800 110.800 204.200 111.200 ;
        RECT 210.200 110.800 210.600 111.200 ;
        RECT 208.600 108.100 209.000 108.200 ;
        RECT 209.400 108.100 209.800 108.200 ;
        RECT 208.600 107.800 209.800 108.100 ;
        RECT 211.000 103.200 211.300 133.800 ;
        RECT 211.800 115.200 212.100 205.800 ;
        RECT 222.200 196.200 222.500 233.800 ;
        RECT 247.000 225.800 247.400 226.200 ;
        RECT 234.200 224.800 234.600 225.200 ;
        RECT 246.200 224.800 246.600 225.200 ;
        RECT 226.200 215.800 226.600 216.200 ;
        RECT 212.600 196.100 213.000 196.200 ;
        RECT 213.400 196.100 213.800 196.200 ;
        RECT 212.600 195.800 213.800 196.100 ;
        RECT 222.200 195.800 222.600 196.200 ;
        RECT 215.800 193.800 216.200 194.200 ;
        RECT 212.600 169.800 213.000 170.200 ;
        RECT 212.600 169.200 212.900 169.800 ;
        RECT 212.600 168.800 213.000 169.200 ;
        RECT 215.800 135.200 216.100 193.800 ;
        RECT 226.200 176.200 226.500 215.800 ;
        RECT 227.800 211.800 228.200 212.200 ;
        RECT 227.800 210.200 228.100 211.800 ;
        RECT 227.800 209.800 228.200 210.200 ;
        RECT 227.800 206.800 228.200 207.200 ;
        RECT 229.400 206.800 229.800 207.200 ;
        RECT 226.200 175.800 226.600 176.200 ;
        RECT 223.000 174.800 223.400 175.200 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 216.600 166.100 217.000 166.200 ;
        RECT 217.400 166.100 217.800 166.200 ;
        RECT 216.600 165.800 217.800 166.100 ;
        RECT 216.600 162.800 217.000 163.200 ;
        RECT 216.600 136.200 216.900 162.800 ;
        RECT 223.000 159.200 223.300 174.800 ;
        RECT 223.800 172.800 224.200 173.200 ;
        RECT 223.000 158.800 223.400 159.200 ;
        RECT 219.800 152.800 220.200 153.200 ;
        RECT 216.600 135.800 217.000 136.200 ;
        RECT 219.800 135.200 220.100 152.800 ;
        RECT 215.800 134.800 216.200 135.200 ;
        RECT 219.000 135.100 219.400 135.200 ;
        RECT 219.800 135.100 220.200 135.200 ;
        RECT 219.000 134.800 220.200 135.100 ;
        RECT 211.800 114.800 212.200 115.200 ;
        RECT 211.000 102.800 211.400 103.200 ;
        RECT 206.200 101.800 206.600 102.200 ;
        RECT 206.200 70.200 206.500 101.800 ;
        RECT 207.000 77.800 207.400 78.200 ;
        RECT 206.200 69.800 206.600 70.200 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 203.000 66.200 203.300 66.800 ;
        RECT 203.000 65.800 203.400 66.200 ;
        RECT 206.200 64.800 206.600 65.200 ;
        RECT 206.200 40.200 206.500 64.800 ;
        RECT 206.200 39.800 206.600 40.200 ;
        RECT 202.200 34.800 202.600 35.200 ;
        RECT 201.400 33.800 201.800 34.200 ;
        RECT 201.400 27.200 201.700 33.800 ;
        RECT 201.400 26.800 201.800 27.200 ;
        RECT 207.000 26.200 207.300 77.800 ;
        RECT 210.200 76.800 210.600 77.200 ;
        RECT 210.200 75.200 210.500 76.800 ;
        RECT 210.200 74.800 210.600 75.200 ;
        RECT 211.000 61.200 211.300 102.800 ;
        RECT 211.000 60.800 211.400 61.200 ;
        RECT 211.800 46.200 212.100 114.800 ;
        RECT 212.600 108.800 213.000 109.200 ;
        RECT 212.600 105.200 212.900 108.800 ;
        RECT 212.600 104.800 213.000 105.200 ;
        RECT 215.800 71.200 216.100 134.800 ;
        RECT 221.400 91.800 221.800 92.200 ;
        RECT 218.200 87.100 218.600 87.200 ;
        RECT 219.000 87.100 219.400 87.200 ;
        RECT 218.200 86.800 219.400 87.100 ;
        RECT 216.600 85.800 217.000 86.200 ;
        RECT 215.800 70.800 216.200 71.200 ;
        RECT 216.600 62.200 216.900 85.800 ;
        RECT 221.400 82.200 221.700 91.800 ;
        RECT 223.000 86.800 223.400 87.200 ;
        RECT 221.400 81.800 221.800 82.200 ;
        RECT 223.000 78.200 223.300 86.800 ;
        RECT 223.800 81.200 224.100 172.800 ;
        RECT 224.600 161.200 224.900 174.800 ;
        RECT 227.800 174.200 228.100 206.800 ;
        RECT 229.400 202.200 229.700 206.800 ;
        RECT 231.000 202.800 231.400 203.200 ;
        RECT 229.400 201.800 229.800 202.200 ;
        RECT 227.800 173.800 228.200 174.200 ;
        RECT 229.400 173.200 229.700 201.800 ;
        RECT 231.000 175.200 231.300 202.800 ;
        RECT 234.200 189.200 234.500 224.800 ;
        RECT 237.400 222.800 237.800 223.200 ;
        RECT 234.200 188.800 234.600 189.200 ;
        RECT 234.200 186.200 234.500 188.800 ;
        RECT 237.400 186.200 237.700 222.800 ;
        RECT 238.200 190.800 238.600 191.200 ;
        RECT 234.200 185.800 234.600 186.200 ;
        RECT 237.400 185.800 237.800 186.200 ;
        RECT 231.000 174.800 231.400 175.200 ;
        RECT 229.400 172.800 229.800 173.200 ;
        RECT 224.600 160.800 225.000 161.200 ;
        RECT 226.200 142.800 226.600 143.200 ;
        RECT 223.800 80.800 224.200 81.200 ;
        RECT 223.000 77.800 223.400 78.200 ;
        RECT 219.000 65.800 219.400 66.200 ;
        RECT 216.600 61.800 217.000 62.200 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 219.000 31.200 219.300 65.800 ;
        RECT 219.800 45.800 220.200 46.200 ;
        RECT 219.000 30.800 219.400 31.200 ;
        RECT 207.800 27.800 208.200 28.200 ;
        RECT 207.800 27.200 208.100 27.800 ;
        RECT 207.800 26.800 208.200 27.200 ;
        RECT 207.000 25.800 207.400 26.200 ;
        RECT 193.400 20.800 193.800 21.200 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 179.000 12.800 179.400 13.200 ;
        RECT 179.000 9.200 179.300 12.800 ;
        RECT 179.000 8.800 179.400 9.200 ;
        RECT 219.800 8.200 220.100 45.800 ;
        RECT 226.200 37.200 226.500 142.800 ;
        RECT 230.200 127.800 230.600 128.200 ;
        RECT 227.000 116.800 227.400 117.200 ;
        RECT 227.000 116.200 227.300 116.800 ;
        RECT 227.000 115.800 227.400 116.200 ;
        RECT 230.200 108.200 230.500 127.800 ;
        RECT 231.000 120.200 231.300 174.800 ;
        RECT 231.800 146.800 232.200 147.200 ;
        RECT 231.800 124.200 232.100 146.800 ;
        RECT 234.200 134.200 234.500 185.800 ;
        RECT 235.000 181.800 235.400 182.200 ;
        RECT 235.000 166.200 235.300 181.800 ;
        RECT 235.000 165.800 235.400 166.200 ;
        RECT 234.200 133.800 234.600 134.200 ;
        RECT 231.800 123.800 232.200 124.200 ;
        RECT 231.000 119.800 231.400 120.200 ;
        RECT 232.600 115.800 233.000 116.200 ;
        RECT 230.200 107.800 230.600 108.200 ;
        RECT 231.800 80.800 232.200 81.200 ;
        RECT 231.000 75.800 231.400 76.200 ;
        RECT 229.400 71.800 229.800 72.200 ;
        RECT 229.400 56.200 229.700 71.800 ;
        RECT 229.400 55.800 229.800 56.200 ;
        RECT 231.000 55.200 231.300 75.800 ;
        RECT 231.800 66.200 232.100 80.800 ;
        RECT 231.800 65.800 232.200 66.200 ;
        RECT 231.000 54.800 231.400 55.200 ;
        RECT 231.000 46.200 231.300 54.800 ;
        RECT 231.000 45.800 231.400 46.200 ;
        RECT 226.200 36.800 226.600 37.200 ;
        RECT 232.600 36.200 232.900 115.800 ;
        RECT 235.000 81.200 235.300 165.800 ;
        RECT 237.400 118.200 237.700 185.800 ;
        RECT 238.200 167.200 238.500 190.800 ;
        RECT 246.200 180.200 246.500 224.800 ;
        RECT 247.000 186.200 247.300 225.800 ;
        RECT 255.000 221.800 255.400 222.200 ;
        RECT 252.600 216.800 253.000 217.200 ;
        RECT 247.000 185.800 247.400 186.200 ;
        RECT 246.200 179.800 246.600 180.200 ;
        RECT 244.600 172.800 245.000 173.200 ;
        RECT 238.200 166.800 238.600 167.200 ;
        RECT 238.200 147.200 238.500 166.800 ;
        RECT 238.200 146.800 238.600 147.200 ;
        RECT 238.200 136.200 238.500 146.800 ;
        RECT 238.200 135.800 238.600 136.200 ;
        RECT 239.800 126.800 240.200 127.200 ;
        RECT 237.400 117.800 237.800 118.200 ;
        RECT 235.000 80.800 235.400 81.200 ;
        RECT 232.600 35.800 233.000 36.200 ;
        RECT 221.400 29.100 221.800 29.200 ;
        RECT 220.600 28.800 221.800 29.100 ;
        RECT 220.600 15.200 220.900 28.800 ;
        RECT 232.600 17.200 232.900 35.800 ;
        RECT 237.400 30.200 237.700 117.800 ;
        RECT 239.800 107.200 240.100 126.800 ;
        RECT 244.600 123.200 244.900 172.800 ;
        RECT 246.200 165.200 246.500 179.800 ;
        RECT 246.200 164.800 246.600 165.200 ;
        RECT 247.000 124.200 247.300 185.800 ;
        RECT 248.600 173.800 249.000 174.200 ;
        RECT 247.800 154.100 248.200 154.200 ;
        RECT 248.600 154.100 248.900 173.800 ;
        RECT 247.800 153.800 248.900 154.100 ;
        RECT 248.600 144.800 249.000 145.200 ;
        RECT 247.000 123.800 247.400 124.200 ;
        RECT 244.600 122.800 245.000 123.200 ;
        RECT 239.800 106.800 240.200 107.200 ;
        RECT 242.200 80.100 242.600 80.200 ;
        RECT 242.200 79.800 243.300 80.100 ;
        RECT 238.200 77.800 238.600 78.200 ;
        RECT 237.400 29.800 237.800 30.200 ;
        RECT 237.400 20.200 237.700 29.800 ;
        RECT 238.200 27.200 238.500 77.800 ;
        RECT 242.200 68.800 242.600 69.200 ;
        RECT 239.800 68.100 240.200 68.200 ;
        RECT 240.600 68.100 241.000 68.200 ;
        RECT 239.800 67.800 241.000 68.100 ;
        RECT 242.200 49.200 242.500 68.800 ;
        RECT 242.200 48.800 242.600 49.200 ;
        RECT 243.000 44.200 243.300 79.800 ;
        RECT 245.400 72.800 245.800 73.200 ;
        RECT 243.800 71.800 244.200 72.200 ;
        RECT 243.000 43.800 243.400 44.200 ;
        RECT 243.800 42.200 244.100 71.800 ;
        RECT 245.400 54.200 245.700 72.800 ;
        RECT 245.400 53.800 245.800 54.200 ;
        RECT 243.800 41.800 244.200 42.200 ;
        RECT 238.200 26.800 238.600 27.200 ;
        RECT 247.000 25.200 247.300 123.800 ;
        RECT 247.800 117.800 248.200 118.200 ;
        RECT 247.800 68.200 248.100 117.800 ;
        RECT 248.600 96.200 248.900 144.800 ;
        RECT 248.600 95.800 249.000 96.200 ;
        RECT 248.600 75.800 249.000 76.200 ;
        RECT 247.800 67.800 248.200 68.200 ;
        RECT 248.600 66.200 248.900 75.800 ;
        RECT 248.600 65.800 249.000 66.200 ;
        RECT 251.800 65.800 252.200 66.200 ;
        RECT 247.000 24.800 247.400 25.200 ;
        RECT 237.400 19.800 237.800 20.200 ;
        RECT 251.800 18.200 252.100 65.800 ;
        RECT 251.800 17.800 252.200 18.200 ;
        RECT 232.600 16.800 233.000 17.200 ;
        RECT 252.600 16.200 252.900 216.800 ;
        RECT 254.200 154.800 254.600 155.200 ;
        RECT 254.200 45.200 254.500 154.800 ;
        RECT 254.200 44.800 254.600 45.200 ;
        RECT 254.200 19.200 254.500 44.800 ;
        RECT 255.000 33.200 255.300 221.800 ;
        RECT 259.000 210.800 259.400 211.200 ;
        RECT 255.800 196.800 256.200 197.200 ;
        RECT 255.800 117.200 256.100 196.800 ;
        RECT 257.400 167.100 257.800 167.200 ;
        RECT 258.200 167.100 258.600 167.200 ;
        RECT 257.400 166.800 258.600 167.100 ;
        RECT 257.400 163.800 257.800 164.200 ;
        RECT 257.400 129.200 257.700 163.800 ;
        RECT 259.000 155.200 259.300 210.800 ;
        RECT 259.000 154.800 259.400 155.200 ;
        RECT 263.000 142.800 263.400 143.200 ;
        RECT 258.200 136.800 258.600 137.200 ;
        RECT 257.400 128.800 257.800 129.200 ;
        RECT 255.800 116.800 256.200 117.200 ;
        RECT 257.400 112.200 257.700 128.800 ;
        RECT 258.200 115.200 258.500 136.800 ;
        RECT 263.000 119.200 263.300 142.800 ;
        RECT 263.000 118.800 263.400 119.200 ;
        RECT 258.200 114.800 258.600 115.200 ;
        RECT 257.400 111.800 257.800 112.200 ;
        RECT 257.400 88.200 257.700 111.800 ;
        RECT 257.400 87.800 257.800 88.200 ;
        RECT 259.800 55.800 260.200 56.200 ;
        RECT 259.800 40.200 260.100 55.800 ;
        RECT 259.800 39.800 260.200 40.200 ;
        RECT 255.000 32.800 255.400 33.200 ;
        RECT 255.000 19.200 255.300 32.800 ;
        RECT 254.200 18.800 254.600 19.200 ;
        RECT 255.000 18.800 255.400 19.200 ;
        RECT 252.600 15.800 253.000 16.200 ;
        RECT 220.600 14.800 221.000 15.200 ;
        RECT 219.800 7.800 220.200 8.200 ;
        RECT 94.200 5.800 94.600 6.200 ;
        RECT 113.400 5.800 113.800 6.200 ;
        RECT 175.800 6.100 176.200 6.200 ;
        RECT 176.600 6.100 177.000 6.200 ;
        RECT 175.800 5.800 177.000 6.100 ;
        RECT 11.800 4.800 12.200 5.200 ;
        RECT 62.200 4.800 62.600 5.200 ;
      LAYER via4 ;
        RECT 126.200 225.800 126.600 226.200 ;
        RECT 29.400 132.800 29.800 133.200 ;
        RECT 47.800 146.800 48.200 147.200 ;
        RECT 45.400 127.800 45.800 128.200 ;
        RECT 41.400 67.800 41.800 68.200 ;
        RECT 46.200 63.800 46.600 64.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 80.600 192.800 81.000 193.200 ;
        RECT 95.800 165.800 96.200 166.200 ;
        RECT 103.800 172.800 104.200 173.200 ;
        RECT 98.200 145.800 98.600 146.200 ;
        RECT 90.200 54.800 90.600 55.200 ;
        RECT 55.000 26.800 55.400 27.200 ;
        RECT 109.400 124.800 109.800 125.200 ;
        RECT 119.800 167.800 120.200 168.200 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 143.800 162.800 144.200 163.200 ;
        RECT 147.800 165.800 148.200 166.200 ;
        RECT 154.200 105.800 154.600 106.200 ;
        RECT 157.400 76.800 157.800 77.200 ;
        RECT 175.800 164.800 176.200 165.200 ;
        RECT 169.400 135.800 169.800 136.200 ;
        RECT 168.600 124.800 169.000 125.200 ;
        RECT 219.800 134.800 220.200 135.200 ;
      LAYER metal5 ;
        RECT 126.200 226.100 126.600 226.200 ;
        RECT 173.400 226.100 173.800 226.200 ;
        RECT 126.200 225.800 173.800 226.100 ;
        RECT 30.200 206.100 30.600 206.200 ;
        RECT 44.600 206.100 45.000 206.200 ;
        RECT 30.200 205.800 45.000 206.100 ;
        RECT 144.600 196.100 145.000 196.200 ;
        RECT 212.600 196.100 213.000 196.200 ;
        RECT 144.600 195.800 213.000 196.100 ;
        RECT 42.200 193.100 42.600 193.200 ;
        RECT 80.600 193.100 81.000 193.200 ;
        RECT 42.200 192.800 81.000 193.100 ;
        RECT 151.800 184.100 152.200 184.200 ;
        RECT 198.200 184.100 198.600 184.200 ;
        RECT 151.800 183.800 198.600 184.100 ;
        RECT 44.600 175.100 45.000 175.200 ;
        RECT 81.400 175.100 81.800 175.200 ;
        RECT 44.600 174.800 81.800 175.100 ;
        RECT 35.800 174.100 36.200 174.200 ;
        RECT 47.000 174.100 47.400 174.200 ;
        RECT 121.400 174.100 121.800 174.200 ;
        RECT 35.800 173.800 40.100 174.100 ;
        RECT 47.000 173.800 121.800 174.100 ;
        RECT 39.800 173.200 40.100 173.800 ;
        RECT 39.800 172.800 40.200 173.200 ;
        RECT 48.600 173.100 49.000 173.200 ;
        RECT 103.800 173.100 104.200 173.200 ;
        RECT 48.600 172.800 104.200 173.100 ;
        RECT 192.600 169.100 193.000 169.200 ;
        RECT 212.600 169.100 213.000 169.200 ;
        RECT 192.600 168.800 213.000 169.100 ;
        RECT 119.800 168.100 120.200 168.200 ;
        RECT 187.000 168.100 187.400 168.200 ;
        RECT 119.800 167.800 187.400 168.100 ;
        RECT 201.400 167.800 201.800 168.200 ;
        RECT 104.600 167.100 105.000 167.200 ;
        RECT 201.400 167.100 201.700 167.800 ;
        RECT 104.600 166.800 201.700 167.100 ;
        RECT 211.000 167.100 211.400 167.200 ;
        RECT 257.400 167.100 257.800 167.200 ;
        RECT 211.000 166.800 257.800 167.100 ;
        RECT 39.000 166.100 39.400 166.200 ;
        RECT 75.800 166.100 76.200 166.200 ;
        RECT 39.000 165.800 76.200 166.100 ;
        RECT 95.800 166.100 96.200 166.200 ;
        RECT 147.800 166.100 148.200 166.200 ;
        RECT 95.800 165.800 148.200 166.100 ;
        RECT 166.200 166.100 166.600 166.200 ;
        RECT 216.600 166.100 217.000 166.200 ;
        RECT 166.200 165.800 217.000 166.100 ;
        RECT 140.600 165.100 141.000 165.200 ;
        RECT 171.800 165.100 172.200 165.200 ;
        RECT 140.600 164.800 172.200 165.100 ;
        RECT 175.800 165.100 176.200 165.200 ;
        RECT 195.800 165.100 196.200 165.200 ;
        RECT 175.800 164.800 196.200 165.100 ;
        RECT 143.800 163.100 144.200 163.200 ;
        RECT 194.200 163.100 194.600 163.200 ;
        RECT 143.800 162.800 194.600 163.100 ;
        RECT 131.800 159.100 132.200 159.200 ;
        RECT 168.600 159.100 169.000 159.200 ;
        RECT 131.800 158.800 169.000 159.100 ;
        RECT 171.800 157.100 172.200 157.200 ;
        RECT 195.800 157.100 196.200 157.200 ;
        RECT 171.800 156.800 196.200 157.100 ;
        RECT 142.200 155.100 142.600 155.200 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 142.200 154.800 148.200 155.100 ;
        RECT 156.600 155.100 157.000 155.200 ;
        RECT 169.400 155.100 169.800 155.200 ;
        RECT 156.600 154.800 169.800 155.100 ;
        RECT 175.000 155.100 175.400 155.200 ;
        RECT 203.000 155.100 203.400 155.200 ;
        RECT 175.000 154.800 203.400 155.100 ;
        RECT 147.000 154.100 147.400 154.200 ;
        RECT 169.400 154.100 169.800 154.200 ;
        RECT 147.000 153.800 169.800 154.100 ;
        RECT 47.800 147.100 48.200 147.200 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 47.800 146.800 80.200 147.100 ;
        RECT 98.200 146.100 98.600 146.200 ;
        RECT 123.800 146.100 124.200 146.200 ;
        RECT 143.000 146.100 143.400 146.200 ;
        RECT 98.200 145.800 143.400 146.100 ;
        RECT 112.600 145.100 113.000 145.200 ;
        RECT 207.800 145.100 208.200 145.200 ;
        RECT 112.600 144.800 208.200 145.100 ;
        RECT 27.800 137.100 28.200 137.200 ;
        RECT 35.800 137.100 36.200 137.200 ;
        RECT 179.000 137.100 179.400 137.200 ;
        RECT 27.800 136.800 179.400 137.100 ;
        RECT 101.400 135.800 101.800 136.200 ;
        RECT 169.400 136.100 169.800 136.200 ;
        RECT 182.200 136.100 182.600 136.200 ;
        RECT 169.400 135.800 182.600 136.100 ;
        RECT 101.400 135.100 101.700 135.800 ;
        RECT 119.800 135.100 120.200 135.200 ;
        RECT 101.400 134.800 120.200 135.100 ;
        RECT 187.000 135.100 187.400 135.200 ;
        RECT 219.800 135.100 220.200 135.200 ;
        RECT 187.000 134.800 220.200 135.100 ;
        RECT 104.600 134.100 105.000 134.200 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 144.600 134.100 145.000 134.200 ;
        RECT 104.600 133.800 145.000 134.100 ;
        RECT 155.000 134.100 155.400 134.200 ;
        RECT 199.000 134.100 199.400 134.200 ;
        RECT 155.000 133.800 199.400 134.100 ;
        RECT 29.400 133.100 29.800 133.200 ;
        RECT 106.200 133.100 106.600 133.200 ;
        RECT 29.400 132.800 106.600 133.100 ;
        RECT 29.400 128.100 29.800 128.200 ;
        RECT 45.400 128.100 45.800 128.200 ;
        RECT 29.400 127.800 45.800 128.100 ;
        RECT 85.400 127.100 85.800 127.200 ;
        RECT 111.000 127.100 111.400 127.200 ;
        RECT 85.400 126.800 111.400 127.100 ;
        RECT 117.400 126.800 117.800 127.200 ;
        RECT 65.400 126.100 65.800 126.200 ;
        RECT 75.800 126.100 76.200 126.200 ;
        RECT 81.400 126.100 81.800 126.200 ;
        RECT 65.400 125.800 81.800 126.100 ;
        RECT 117.400 126.100 117.700 126.800 ;
        RECT 144.600 126.100 145.000 126.200 ;
        RECT 117.400 125.800 145.000 126.100 ;
        RECT 47.800 125.100 48.200 125.200 ;
        RECT 104.600 125.100 105.000 125.200 ;
        RECT 47.800 124.800 105.000 125.100 ;
        RECT 109.400 125.100 109.800 125.200 ;
        RECT 119.000 125.100 119.400 125.200 ;
        RECT 109.400 124.800 119.400 125.100 ;
        RECT 135.000 125.100 135.400 125.200 ;
        RECT 168.600 125.100 169.000 125.200 ;
        RECT 135.000 124.800 169.000 125.100 ;
        RECT 107.800 124.100 108.200 124.200 ;
        RECT 205.400 124.100 205.800 124.200 ;
        RECT 107.800 123.800 205.800 124.100 ;
        RECT 227.000 116.800 227.400 117.200 ;
        RECT 152.600 116.100 153.000 116.200 ;
        RECT 227.000 116.100 227.300 116.800 ;
        RECT 152.600 115.800 227.300 116.100 ;
        RECT 210.200 115.100 210.600 115.200 ;
        RECT 148.600 114.800 210.600 115.100 ;
        RECT 148.600 114.200 148.900 114.800 ;
        RECT 148.600 113.800 149.000 114.200 ;
        RECT 159.800 108.100 160.200 108.200 ;
        RECT 208.600 108.100 209.000 108.200 ;
        RECT 159.800 107.800 209.000 108.100 ;
        RECT 154.200 106.100 154.600 106.200 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 154.200 105.800 166.600 106.100 ;
        RECT 197.400 87.100 197.800 87.200 ;
        RECT 218.200 87.100 218.600 87.200 ;
        RECT 197.400 86.800 218.600 87.100 ;
        RECT 157.400 77.100 157.800 77.200 ;
        RECT 210.200 77.100 210.600 77.200 ;
        RECT 157.400 76.800 210.600 77.100 ;
        RECT 142.200 76.100 142.600 76.200 ;
        RECT 194.200 76.100 194.600 76.200 ;
        RECT 142.200 75.800 194.600 76.100 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 112.600 75.100 113.000 75.200 ;
        RECT 106.200 74.800 113.000 75.100 ;
        RECT 127.800 75.100 128.200 75.200 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 127.800 74.800 197.800 75.100 ;
        RECT 183.000 74.100 183.400 74.200 ;
        RECT 188.600 74.100 189.000 74.200 ;
        RECT 183.000 73.800 189.000 74.100 ;
        RECT 109.400 71.100 109.800 71.200 ;
        RECT 179.000 71.100 179.400 71.200 ;
        RECT 109.400 70.800 179.400 71.100 ;
        RECT 41.400 68.100 41.800 68.200 ;
        RECT 96.600 68.100 97.000 68.200 ;
        RECT 41.400 67.800 97.000 68.100 ;
        RECT 128.600 68.100 129.000 68.200 ;
        RECT 150.200 68.100 150.600 68.200 ;
        RECT 128.600 67.800 150.600 68.100 ;
        RECT 169.400 68.100 169.800 68.200 ;
        RECT 239.800 68.100 240.200 68.200 ;
        RECT 169.400 67.800 240.200 68.100 ;
        RECT 66.200 66.800 66.600 67.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 136.600 67.100 137.000 67.200 ;
        RECT 166.200 67.100 166.600 67.200 ;
        RECT 121.400 66.800 133.700 67.100 ;
        RECT 136.600 66.800 166.600 67.100 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 66.200 66.100 66.500 66.800 ;
        RECT 133.400 66.200 133.700 66.800 ;
        RECT 56.600 65.800 66.500 66.100 ;
        RECT 93.400 66.100 93.800 66.200 ;
        RECT 123.800 66.100 124.200 66.200 ;
        RECT 93.400 65.800 124.200 66.100 ;
        RECT 133.400 65.800 133.800 66.200 ;
        RECT 165.400 66.100 165.800 66.200 ;
        RECT 203.000 66.100 203.300 66.800 ;
        RECT 165.400 65.800 203.300 66.100 ;
        RECT 48.600 65.100 49.000 65.200 ;
        RECT 57.400 65.100 57.800 65.200 ;
        RECT 48.600 64.800 57.800 65.100 ;
        RECT 124.600 65.100 125.000 65.200 ;
        RECT 196.600 65.100 197.000 65.200 ;
        RECT 124.600 64.800 197.000 65.100 ;
        RECT 46.200 64.100 46.600 64.200 ;
        RECT 74.200 64.100 74.600 64.200 ;
        RECT 46.200 63.800 74.600 64.100 ;
        RECT 146.200 64.100 146.600 64.200 ;
        RECT 166.200 64.100 166.600 64.200 ;
        RECT 146.200 63.800 166.600 64.100 ;
        RECT 35.000 63.100 35.400 63.200 ;
        RECT 49.400 63.100 49.800 63.200 ;
        RECT 113.400 63.100 113.800 63.200 ;
        RECT 35.000 62.800 113.800 63.100 ;
        RECT 90.200 55.100 90.600 55.200 ;
        RECT 143.000 55.100 143.400 55.200 ;
        RECT 90.200 54.800 143.400 55.100 ;
        RECT 115.000 54.100 115.400 54.200 ;
        RECT 159.000 54.100 159.400 54.200 ;
        RECT 115.000 53.800 159.400 54.100 ;
        RECT 134.200 36.100 134.600 36.200 ;
        RECT 167.000 36.100 167.400 36.200 ;
        RECT 134.200 35.800 167.400 36.100 ;
        RECT 59.800 35.100 60.200 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 59.800 34.800 105.800 35.100 ;
        RECT 63.000 28.100 63.400 28.200 ;
        RECT 118.200 28.100 118.600 28.200 ;
        RECT 63.000 27.800 118.600 28.100 ;
        RECT 207.800 27.800 208.200 28.200 ;
        RECT 55.000 27.100 55.400 27.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 55.000 26.800 95.400 27.100 ;
        RECT 172.600 27.100 173.000 27.200 ;
        RECT 207.800 27.100 208.100 27.800 ;
        RECT 172.600 26.800 208.100 27.100 ;
        RECT 19.800 18.100 20.200 18.200 ;
        RECT 73.400 18.100 73.800 18.200 ;
        RECT 19.800 17.800 73.800 18.100 ;
        RECT 91.800 18.100 92.200 18.200 ;
        RECT 159.000 18.100 159.400 18.200 ;
        RECT 91.800 17.800 159.400 18.100 ;
        RECT 92.600 15.100 93.000 15.200 ;
        RECT 99.000 15.100 99.400 15.200 ;
        RECT 92.600 14.800 99.400 15.100 ;
        RECT 94.200 6.100 94.600 6.200 ;
        RECT 175.800 6.100 176.200 6.200 ;
        RECT 94.200 5.800 176.200 6.100 ;
  END
END ram32_sdram_2split
END LIBRARY

