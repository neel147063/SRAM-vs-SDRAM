VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram32_sdram_3split
  CLASS BLOCK ;
  FOREIGN ram32_sdram_3split ;
  ORIGIN 2.600 3.000 ;
  SIZE 236.400 BY 216.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.600 200.800 1.000 205.100 ;
        RECT 2.200 200.800 2.600 205.100 ;
        RECT 3.800 200.800 4.200 205.100 ;
        RECT 5.400 200.800 5.800 205.100 ;
        RECT 7.000 200.800 7.400 205.100 ;
        RECT 7.800 200.800 8.200 205.100 ;
        RECT 9.400 200.800 9.800 205.100 ;
        RECT 11.000 200.800 11.400 205.100 ;
        RECT 12.600 200.800 13.000 205.100 ;
        RECT 14.200 200.800 14.600 205.100 ;
        RECT 15.800 200.800 16.200 205.000 ;
        RECT 18.600 200.800 19.000 203.100 ;
        RECT 20.200 200.800 20.600 203.100 ;
        RECT 23.000 200.800 23.400 205.100 ;
        RECT 24.600 200.800 25.000 205.100 ;
        RECT 26.700 200.800 27.100 203.100 ;
        RECT 28.100 200.800 28.500 203.100 ;
        RECT 30.200 200.800 30.600 205.100 ;
        RECT 31.800 200.800 32.200 205.000 ;
        RECT 34.600 200.800 35.000 203.100 ;
        RECT 36.200 200.800 36.600 203.100 ;
        RECT 39.000 200.800 39.400 205.100 ;
        RECT 42.200 200.800 42.600 205.100 ;
        RECT 43.800 200.800 44.200 204.500 ;
        RECT 46.200 200.800 46.600 205.000 ;
        RECT 49.000 200.800 49.400 203.100 ;
        RECT 50.600 200.800 51.000 203.100 ;
        RECT 53.400 200.800 53.800 205.100 ;
        RECT 55.000 200.800 55.400 205.100 ;
        RECT 57.100 200.800 57.500 203.100 ;
        RECT 58.500 200.800 58.900 203.100 ;
        RECT 60.600 200.800 61.000 205.100 ;
        RECT 61.400 200.800 61.800 205.100 ;
        RECT 63.000 200.800 63.400 204.500 ;
        RECT 65.400 200.800 65.800 205.000 ;
        RECT 68.200 200.800 68.600 203.100 ;
        RECT 69.800 200.800 70.200 203.100 ;
        RECT 72.600 200.800 73.000 205.100 ;
        RECT 75.000 200.800 75.400 205.100 ;
        RECT 77.800 200.800 78.200 203.100 ;
        RECT 79.400 200.800 79.800 203.100 ;
        RECT 82.200 200.800 82.600 205.000 ;
        RECT 83.800 200.800 84.200 205.100 ;
        RECT 85.900 200.800 86.300 203.100 ;
        RECT 87.300 200.800 87.700 203.100 ;
        RECT 89.400 200.800 89.800 205.100 ;
        RECT 92.600 200.800 93.000 205.000 ;
        RECT 95.400 200.800 95.800 203.100 ;
        RECT 97.000 200.800 97.400 203.100 ;
        RECT 99.800 200.800 100.200 205.100 ;
        RECT 102.200 200.800 102.600 205.000 ;
        RECT 105.000 200.800 105.400 203.100 ;
        RECT 106.600 200.800 107.000 203.100 ;
        RECT 109.400 200.800 109.800 205.100 ;
        RECT 111.000 200.800 111.400 205.100 ;
        RECT 113.100 200.800 113.500 203.100 ;
        RECT 114.500 200.800 114.900 203.100 ;
        RECT 116.600 200.800 117.000 205.100 ;
        RECT 117.400 200.800 117.800 205.100 ;
        RECT 119.500 200.800 119.900 203.100 ;
        RECT 120.600 200.800 121.000 205.100 ;
        RECT 122.700 200.800 123.100 203.100 ;
        RECT 124.600 200.800 125.000 205.000 ;
        RECT 127.400 200.800 127.800 203.100 ;
        RECT 129.000 200.800 129.400 203.100 ;
        RECT 131.800 200.800 132.200 205.100 ;
        RECT 133.400 200.800 133.800 205.100 ;
        RECT 135.000 200.800 135.400 204.500 ;
        RECT 136.600 200.800 137.000 205.100 ;
        RECT 138.200 200.800 138.600 205.100 ;
        RECT 139.800 200.800 140.200 205.100 ;
        RECT 143.000 200.800 143.400 205.000 ;
        RECT 145.800 200.800 146.200 203.100 ;
        RECT 147.400 200.800 147.800 203.100 ;
        RECT 150.200 200.800 150.600 205.100 ;
        RECT 151.800 200.800 152.200 205.100 ;
        RECT 153.900 200.800 154.300 203.100 ;
        RECT 155.000 200.800 155.400 203.100 ;
        RECT 156.600 200.800 157.000 203.100 ;
        RECT 158.200 200.800 158.600 204.500 ;
        RECT 159.800 200.800 160.200 205.100 ;
        RECT 161.400 200.800 161.800 205.100 ;
        RECT 164.200 200.800 164.600 203.100 ;
        RECT 165.800 200.800 166.200 203.100 ;
        RECT 168.600 200.800 169.000 205.000 ;
        RECT 170.200 200.800 170.600 205.100 ;
        RECT 172.300 200.800 172.700 203.100 ;
        RECT 173.400 200.800 173.800 203.100 ;
        RECT 175.000 200.800 175.400 203.100 ;
        RECT 176.600 200.800 177.000 205.000 ;
        RECT 179.400 200.800 179.800 203.100 ;
        RECT 181.000 200.800 181.400 203.100 ;
        RECT 183.800 200.800 184.200 205.100 ;
        RECT 185.400 200.800 185.800 205.100 ;
        RECT 187.000 200.800 187.400 205.100 ;
        RECT 188.600 200.800 189.000 205.100 ;
        RECT 191.000 200.800 191.400 205.100 ;
        RECT 192.600 200.800 193.000 205.100 ;
        RECT 194.200 200.800 194.600 205.100 ;
        RECT 195.800 200.800 196.200 205.100 ;
        RECT 197.400 200.800 197.800 205.100 ;
        RECT 198.800 200.800 199.200 205.100 ;
        RECT 201.400 200.800 201.800 204.900 ;
        RECT 203.000 200.800 203.400 205.100 ;
        RECT 205.100 200.800 205.500 203.100 ;
        RECT 206.200 200.800 206.600 203.100 ;
        RECT 207.800 200.800 208.200 203.100 ;
        RECT 208.600 200.800 209.000 203.100 ;
        RECT 210.200 200.800 210.600 203.100 ;
        RECT 211.800 200.800 212.200 205.100 ;
        RECT 214.600 200.800 215.000 203.100 ;
        RECT 216.200 200.800 216.600 203.100 ;
        RECT 219.000 200.800 219.400 205.000 ;
        RECT 220.600 200.800 221.000 203.100 ;
        RECT 222.200 200.800 222.600 203.100 ;
        RECT 223.000 200.800 223.400 205.100 ;
        RECT 225.100 200.800 225.500 203.100 ;
        RECT 226.200 200.800 226.600 205.100 ;
        RECT 227.800 200.800 228.200 205.100 ;
        RECT 229.400 200.800 229.800 205.100 ;
        RECT 0.200 200.200 231.000 200.800 ;
        RECT 1.400 195.900 1.800 200.200 ;
        RECT 4.200 197.900 4.600 200.200 ;
        RECT 5.800 197.900 6.200 200.200 ;
        RECT 8.600 196.000 9.000 200.200 ;
        RECT 10.500 197.900 10.900 200.200 ;
        RECT 12.600 195.900 13.000 200.200 ;
        RECT 13.700 197.900 14.100 200.200 ;
        RECT 15.800 195.900 16.200 200.200 ;
        RECT 16.900 197.900 17.300 200.200 ;
        RECT 19.000 195.900 19.400 200.200 ;
        RECT 20.100 197.900 20.500 200.200 ;
        RECT 22.200 195.900 22.600 200.200 ;
        RECT 23.000 195.900 23.400 200.200 ;
        RECT 25.100 197.900 25.500 200.200 ;
        RECT 26.500 197.900 26.900 200.200 ;
        RECT 28.600 195.900 29.000 200.200 ;
        RECT 30.200 196.000 30.600 200.200 ;
        RECT 33.000 197.900 33.400 200.200 ;
        RECT 34.600 197.900 35.000 200.200 ;
        RECT 37.400 195.900 37.800 200.200 ;
        RECT 41.400 196.000 41.800 200.200 ;
        RECT 44.200 197.900 44.600 200.200 ;
        RECT 45.800 197.900 46.200 200.200 ;
        RECT 48.600 195.900 49.000 200.200 ;
        RECT 50.500 197.900 50.900 200.200 ;
        RECT 52.600 195.900 53.000 200.200 ;
        RECT 54.000 195.900 54.400 200.200 ;
        RECT 56.600 196.100 57.000 200.200 ;
        RECT 58.200 195.900 58.600 200.200 ;
        RECT 60.300 197.900 60.700 200.200 ;
        RECT 62.200 196.000 62.600 200.200 ;
        RECT 65.000 197.900 65.400 200.200 ;
        RECT 66.600 197.900 67.000 200.200 ;
        RECT 69.400 195.900 69.800 200.200 ;
        RECT 71.000 195.900 71.400 200.200 ;
        RECT 73.100 197.900 73.500 200.200 ;
        RECT 74.200 195.900 74.600 200.200 ;
        RECT 76.300 197.900 76.700 200.200 ;
        RECT 77.700 197.900 78.100 200.200 ;
        RECT 79.800 195.900 80.200 200.200 ;
        RECT 80.900 197.900 81.300 200.200 ;
        RECT 83.000 195.900 83.400 200.200 ;
        RECT 83.800 195.900 84.200 200.200 ;
        RECT 85.900 197.900 86.300 200.200 ;
        RECT 87.000 195.900 87.400 200.200 ;
        RECT 89.100 197.900 89.500 200.200 ;
        RECT 92.600 196.000 93.000 200.200 ;
        RECT 95.400 197.900 95.800 200.200 ;
        RECT 97.000 197.900 97.400 200.200 ;
        RECT 99.800 195.900 100.200 200.200 ;
        RECT 101.400 195.900 101.800 200.200 ;
        RECT 103.500 197.900 103.900 200.200 ;
        RECT 104.600 195.900 105.000 200.200 ;
        RECT 106.700 197.900 107.100 200.200 ;
        RECT 108.600 196.000 109.000 200.200 ;
        RECT 111.400 197.900 111.800 200.200 ;
        RECT 113.000 197.900 113.400 200.200 ;
        RECT 115.800 195.900 116.200 200.200 ;
        RECT 118.200 196.000 118.600 200.200 ;
        RECT 121.000 197.900 121.400 200.200 ;
        RECT 122.600 197.900 123.000 200.200 ;
        RECT 125.400 195.900 125.800 200.200 ;
        RECT 127.000 195.900 127.400 200.200 ;
        RECT 129.100 197.900 129.500 200.200 ;
        RECT 130.500 197.900 130.900 200.200 ;
        RECT 132.600 195.900 133.000 200.200 ;
        RECT 133.400 195.900 133.800 200.200 ;
        RECT 135.500 197.900 135.900 200.200 ;
        RECT 136.900 197.900 137.300 200.200 ;
        RECT 139.000 195.900 139.400 200.200 ;
        RECT 142.200 195.900 142.600 200.200 ;
        RECT 145.000 197.900 145.400 200.200 ;
        RECT 146.600 197.900 147.000 200.200 ;
        RECT 149.400 196.000 149.800 200.200 ;
        RECT 151.800 195.900 152.200 200.200 ;
        RECT 154.600 197.900 155.000 200.200 ;
        RECT 156.200 197.900 156.600 200.200 ;
        RECT 159.000 196.000 159.400 200.200 ;
        RECT 160.600 195.900 161.000 200.200 ;
        RECT 162.700 197.900 163.100 200.200 ;
        RECT 163.800 197.900 164.200 200.200 ;
        RECT 165.400 197.900 165.800 200.200 ;
        RECT 167.000 195.900 167.400 200.200 ;
        RECT 169.800 197.900 170.200 200.200 ;
        RECT 171.400 197.900 171.800 200.200 ;
        RECT 174.200 196.000 174.600 200.200 ;
        RECT 175.800 195.900 176.200 200.200 ;
        RECT 177.900 197.900 178.300 200.200 ;
        RECT 179.000 197.900 179.400 200.200 ;
        RECT 180.600 197.900 181.000 200.200 ;
        RECT 182.000 195.900 182.400 200.200 ;
        RECT 184.600 196.100 185.000 200.200 ;
        RECT 186.200 195.900 186.600 200.200 ;
        RECT 188.300 197.900 188.700 200.200 ;
        RECT 189.400 197.900 189.800 200.200 ;
        RECT 191.000 197.900 191.400 200.200 ;
        RECT 194.200 195.900 194.600 200.200 ;
        RECT 197.000 197.900 197.400 200.200 ;
        RECT 198.600 197.900 199.000 200.200 ;
        RECT 201.400 196.000 201.800 200.200 ;
        RECT 203.000 195.900 203.400 200.200 ;
        RECT 205.100 197.900 205.500 200.200 ;
        RECT 206.200 197.900 206.600 200.200 ;
        RECT 207.800 197.900 208.200 200.200 ;
        RECT 209.400 195.900 209.800 200.200 ;
        RECT 212.200 197.900 212.600 200.200 ;
        RECT 213.800 197.900 214.200 200.200 ;
        RECT 216.600 196.000 217.000 200.200 ;
        RECT 218.200 195.900 218.600 200.200 ;
        RECT 220.300 197.900 220.700 200.200 ;
        RECT 222.200 195.900 222.600 200.200 ;
        RECT 225.000 197.900 225.400 200.200 ;
        RECT 226.600 197.900 227.000 200.200 ;
        RECT 229.400 196.000 229.800 200.200 ;
        RECT 1.400 180.800 1.800 185.000 ;
        RECT 4.200 180.800 4.600 183.100 ;
        RECT 5.800 180.800 6.200 183.100 ;
        RECT 8.600 180.800 9.000 185.100 ;
        RECT 10.500 180.800 10.900 183.100 ;
        RECT 12.600 180.800 13.000 185.100 ;
        RECT 13.700 180.800 14.100 183.100 ;
        RECT 15.800 180.800 16.200 185.100 ;
        RECT 17.400 180.800 17.800 185.000 ;
        RECT 20.200 180.800 20.600 183.100 ;
        RECT 21.800 180.800 22.200 183.100 ;
        RECT 24.600 180.800 25.000 185.100 ;
        RECT 26.200 180.800 26.600 185.100 ;
        RECT 28.300 180.800 28.700 183.100 ;
        RECT 29.700 180.800 30.100 183.100 ;
        RECT 31.800 180.800 32.200 185.100 ;
        RECT 32.600 180.800 33.000 185.100 ;
        RECT 34.700 180.800 35.100 183.100 ;
        RECT 38.000 180.800 38.400 185.100 ;
        RECT 40.600 180.800 41.000 184.900 ;
        RECT 43.000 180.800 43.400 185.000 ;
        RECT 45.800 180.800 46.200 183.100 ;
        RECT 47.400 180.800 47.800 183.100 ;
        RECT 50.200 180.800 50.600 185.100 ;
        RECT 51.800 180.800 52.200 185.100 ;
        RECT 53.900 180.800 54.300 183.100 ;
        RECT 55.300 180.800 55.700 183.100 ;
        RECT 57.400 180.800 57.800 185.100 ;
        RECT 58.500 180.800 58.900 183.100 ;
        RECT 60.600 180.800 61.000 185.100 ;
        RECT 62.200 180.800 62.600 184.900 ;
        RECT 64.800 180.800 65.200 185.100 ;
        RECT 66.500 180.800 66.900 183.100 ;
        RECT 68.600 180.800 69.000 185.100 ;
        RECT 70.200 180.800 70.600 184.500 ;
        RECT 71.800 180.800 72.200 185.100 ;
        RECT 73.200 180.800 73.600 185.100 ;
        RECT 75.800 180.800 76.200 184.900 ;
        RECT 78.200 180.800 78.600 185.100 ;
        RECT 81.000 180.800 81.400 183.100 ;
        RECT 82.600 180.800 83.000 183.100 ;
        RECT 85.400 180.800 85.800 185.000 ;
        RECT 87.300 180.800 87.700 183.100 ;
        RECT 89.400 180.800 89.800 185.100 ;
        RECT 92.100 180.800 92.500 183.100 ;
        RECT 94.200 180.800 94.600 185.100 ;
        RECT 95.800 180.800 96.200 184.900 ;
        RECT 98.400 180.800 98.800 185.100 ;
        RECT 100.600 180.800 101.000 184.900 ;
        RECT 103.200 180.800 103.600 185.100 ;
        RECT 105.200 180.800 105.600 185.100 ;
        RECT 107.800 180.800 108.200 184.900 ;
        RECT 109.400 180.800 109.800 185.100 ;
        RECT 111.000 180.800 111.400 184.500 ;
        RECT 113.400 180.800 113.800 184.500 ;
        RECT 115.000 180.800 115.400 185.100 ;
        RECT 115.800 180.800 116.200 185.100 ;
        RECT 117.900 180.800 118.300 183.100 ;
        RECT 119.300 180.800 119.700 183.100 ;
        RECT 121.400 180.800 121.800 185.100 ;
        RECT 123.000 180.800 123.400 185.100 ;
        RECT 125.800 180.800 126.200 183.100 ;
        RECT 127.400 180.800 127.800 183.100 ;
        RECT 130.200 180.800 130.600 185.000 ;
        RECT 131.800 180.800 132.200 185.100 ;
        RECT 133.400 180.800 133.800 185.100 ;
        RECT 134.800 180.800 135.200 185.100 ;
        RECT 137.400 180.800 137.800 184.900 ;
        RECT 140.600 180.800 141.000 185.100 ;
        RECT 142.700 180.800 143.100 183.100 ;
        RECT 143.800 180.800 144.200 185.100 ;
        RECT 145.900 180.800 146.300 183.100 ;
        RECT 147.000 180.800 147.400 185.100 ;
        RECT 149.100 180.800 149.500 183.100 ;
        RECT 151.000 180.800 151.400 185.000 ;
        RECT 153.800 180.800 154.200 183.100 ;
        RECT 155.400 180.800 155.800 183.100 ;
        RECT 158.200 180.800 158.600 185.100 ;
        RECT 159.800 180.800 160.200 183.100 ;
        RECT 161.400 180.800 161.800 183.100 ;
        RECT 162.500 180.800 162.900 183.100 ;
        RECT 164.600 180.800 165.000 185.100 ;
        RECT 166.200 180.800 166.600 183.100 ;
        RECT 167.800 180.800 168.200 185.100 ;
        RECT 170.600 180.800 171.000 183.100 ;
        RECT 172.200 180.800 172.600 183.100 ;
        RECT 175.000 180.800 175.400 185.000 ;
        RECT 176.600 180.800 177.000 183.100 ;
        RECT 178.200 180.800 178.600 183.100 ;
        RECT 179.300 180.800 179.700 183.100 ;
        RECT 181.400 180.800 181.800 185.100 ;
        RECT 183.000 180.800 183.400 184.900 ;
        RECT 185.600 180.800 186.000 185.100 ;
        RECT 187.800 180.800 188.200 184.900 ;
        RECT 190.400 180.800 190.800 185.100 ;
        RECT 194.200 180.800 194.600 184.900 ;
        RECT 196.800 180.800 197.200 185.100 ;
        RECT 199.000 180.800 199.400 184.900 ;
        RECT 201.600 180.800 202.000 185.100 ;
        RECT 203.800 180.800 204.200 184.900 ;
        RECT 206.400 180.800 206.800 185.100 ;
        RECT 208.600 180.800 209.000 185.100 ;
        RECT 211.400 180.800 211.800 183.100 ;
        RECT 213.000 180.800 213.400 183.100 ;
        RECT 215.800 180.800 216.200 185.000 ;
        RECT 217.400 180.800 217.800 183.100 ;
        RECT 219.000 180.800 219.400 183.100 ;
        RECT 220.100 180.800 220.500 183.100 ;
        RECT 222.200 180.800 222.600 185.100 ;
        RECT 223.000 180.800 223.400 183.100 ;
        RECT 224.600 180.800 225.000 183.100 ;
        RECT 225.700 180.800 226.100 183.100 ;
        RECT 227.800 180.800 228.200 185.100 ;
        RECT 0.200 180.200 231.000 180.800 ;
        RECT 0.600 175.900 1.000 180.200 ;
        RECT 2.200 175.900 2.600 180.200 ;
        RECT 3.800 175.900 4.200 180.200 ;
        RECT 5.400 175.900 5.800 180.200 ;
        RECT 7.000 175.900 7.400 180.200 ;
        RECT 8.600 175.900 9.000 180.200 ;
        RECT 11.400 177.900 11.800 180.200 ;
        RECT 13.000 177.900 13.400 180.200 ;
        RECT 15.800 176.000 16.200 180.200 ;
        RECT 17.400 175.900 17.800 180.200 ;
        RECT 19.000 175.900 19.400 180.200 ;
        RECT 20.600 175.900 21.000 180.200 ;
        RECT 22.200 175.900 22.600 180.200 ;
        RECT 23.800 175.900 24.200 180.200 ;
        RECT 25.400 176.000 25.800 180.200 ;
        RECT 28.200 177.900 28.600 180.200 ;
        RECT 29.800 177.900 30.200 180.200 ;
        RECT 32.600 175.900 33.000 180.200 ;
        RECT 34.500 177.900 34.900 180.200 ;
        RECT 36.600 175.900 37.000 180.200 ;
        RECT 39.600 175.900 40.000 180.200 ;
        RECT 42.200 176.100 42.600 180.200 ;
        RECT 44.600 176.000 45.000 180.200 ;
        RECT 47.400 177.900 47.800 180.200 ;
        RECT 49.000 177.900 49.400 180.200 ;
        RECT 51.800 175.900 52.200 180.200 ;
        RECT 53.400 175.900 53.800 180.200 ;
        RECT 55.500 177.900 55.900 180.200 ;
        RECT 56.900 177.900 57.300 180.200 ;
        RECT 59.000 175.900 59.400 180.200 ;
        RECT 60.600 176.100 61.000 180.200 ;
        RECT 63.200 175.900 63.600 180.200 ;
        RECT 65.200 175.900 65.600 180.200 ;
        RECT 67.800 176.100 68.200 180.200 ;
        RECT 70.200 176.100 70.600 180.200 ;
        RECT 72.800 175.900 73.200 180.200 ;
        RECT 75.000 176.500 75.400 180.200 ;
        RECT 76.600 175.900 77.000 180.200 ;
        RECT 78.200 176.000 78.600 180.200 ;
        RECT 81.000 177.900 81.400 180.200 ;
        RECT 82.600 177.900 83.000 180.200 ;
        RECT 85.400 175.900 85.800 180.200 ;
        RECT 87.000 175.900 87.400 180.200 ;
        RECT 89.100 177.900 89.500 180.200 ;
        RECT 92.100 177.900 92.500 180.200 ;
        RECT 94.200 175.900 94.600 180.200 ;
        RECT 95.000 175.900 95.400 180.200 ;
        RECT 96.600 175.900 97.000 180.200 ;
        RECT 98.200 175.900 98.600 180.200 ;
        RECT 99.000 177.900 99.400 180.200 ;
        RECT 100.600 177.900 101.000 180.200 ;
        RECT 101.400 175.900 101.800 180.200 ;
        RECT 103.000 175.900 103.400 180.200 ;
        RECT 103.800 175.900 104.200 180.200 ;
        RECT 105.900 177.900 106.300 180.200 ;
        RECT 107.300 177.900 107.700 180.200 ;
        RECT 109.400 175.900 109.800 180.200 ;
        RECT 110.200 175.900 110.600 180.200 ;
        RECT 112.300 177.900 112.700 180.200 ;
        RECT 113.400 175.900 113.800 180.200 ;
        RECT 115.500 177.900 115.900 180.200 ;
        RECT 117.400 176.000 117.800 180.200 ;
        RECT 120.200 177.900 120.600 180.200 ;
        RECT 121.800 177.900 122.200 180.200 ;
        RECT 124.600 175.900 125.000 180.200 ;
        RECT 126.800 175.900 127.200 180.200 ;
        RECT 129.400 176.100 129.800 180.200 ;
        RECT 131.000 177.900 131.400 180.200 ;
        RECT 132.600 177.900 133.000 180.200 ;
        RECT 134.000 175.900 134.400 180.200 ;
        RECT 136.600 176.100 137.000 180.200 ;
        RECT 138.200 175.900 138.600 180.200 ;
        RECT 140.300 177.900 140.700 180.200 ;
        RECT 143.800 175.900 144.200 180.200 ;
        RECT 146.600 177.900 147.000 180.200 ;
        RECT 148.200 177.900 148.600 180.200 ;
        RECT 151.000 176.000 151.400 180.200 ;
        RECT 152.600 175.900 153.000 180.200 ;
        RECT 154.700 177.900 155.100 180.200 ;
        RECT 155.800 177.900 156.200 180.200 ;
        RECT 157.400 177.900 157.800 180.200 ;
        RECT 158.200 175.900 158.600 180.200 ;
        RECT 160.300 177.900 160.700 180.200 ;
        RECT 161.400 177.900 161.800 180.200 ;
        RECT 163.000 177.900 163.400 180.200 ;
        RECT 164.600 176.000 165.000 180.200 ;
        RECT 167.400 177.900 167.800 180.200 ;
        RECT 169.000 177.900 169.400 180.200 ;
        RECT 171.800 175.900 172.200 180.200 ;
        RECT 174.200 176.100 174.600 180.200 ;
        RECT 176.800 175.900 177.200 180.200 ;
        RECT 179.000 176.500 179.400 180.200 ;
        RECT 180.600 175.900 181.000 180.200 ;
        RECT 181.400 177.900 181.800 180.200 ;
        RECT 183.000 177.900 183.400 180.200 ;
        RECT 183.800 177.900 184.200 180.200 ;
        RECT 185.400 177.900 185.800 180.200 ;
        RECT 186.200 177.900 186.600 180.200 ;
        RECT 187.800 177.900 188.200 180.200 ;
        RECT 189.400 176.100 189.800 180.200 ;
        RECT 192.000 175.900 192.400 180.200 ;
        RECT 195.000 177.900 195.400 180.200 ;
        RECT 196.600 177.900 197.000 180.200 ;
        RECT 197.700 177.900 198.100 180.200 ;
        RECT 199.800 175.900 200.200 180.200 ;
        RECT 201.400 175.900 201.800 180.200 ;
        RECT 204.200 177.900 204.600 180.200 ;
        RECT 205.800 177.900 206.200 180.200 ;
        RECT 208.600 176.000 209.000 180.200 ;
        RECT 211.000 176.500 211.400 180.200 ;
        RECT 212.600 175.900 213.000 180.200 ;
        RECT 213.400 177.900 213.800 180.200 ;
        RECT 215.000 177.900 215.400 180.200 ;
        RECT 216.600 175.900 217.000 180.200 ;
        RECT 219.400 177.900 219.800 180.200 ;
        RECT 221.000 177.900 221.400 180.200 ;
        RECT 223.800 176.000 224.200 180.200 ;
        RECT 225.400 177.900 225.800 180.200 ;
        RECT 227.000 177.900 227.400 180.200 ;
        RECT 228.100 177.900 228.500 180.200 ;
        RECT 230.200 175.900 230.600 180.200 ;
        RECT 1.400 160.800 1.800 165.000 ;
        RECT 4.200 160.800 4.600 163.100 ;
        RECT 5.800 160.800 6.200 163.100 ;
        RECT 8.600 160.800 9.000 165.100 ;
        RECT 10.200 160.800 10.600 163.100 ;
        RECT 11.800 160.800 12.200 163.100 ;
        RECT 13.400 160.800 13.800 163.100 ;
        RECT 14.500 160.800 14.900 163.100 ;
        RECT 16.600 160.800 17.000 165.100 ;
        RECT 18.200 160.800 18.600 164.500 ;
        RECT 19.800 160.800 20.200 165.100 ;
        RECT 21.400 160.800 21.800 165.000 ;
        RECT 24.200 160.800 24.600 163.100 ;
        RECT 25.800 160.800 26.200 163.100 ;
        RECT 28.600 160.800 29.000 165.100 ;
        RECT 30.200 160.800 30.600 163.100 ;
        RECT 31.800 160.800 32.200 163.100 ;
        RECT 32.900 160.800 33.300 163.100 ;
        RECT 35.000 160.800 35.400 165.100 ;
        RECT 38.200 160.800 38.600 165.000 ;
        RECT 41.000 160.800 41.400 163.100 ;
        RECT 42.600 160.800 43.000 163.100 ;
        RECT 45.400 160.800 45.800 165.100 ;
        RECT 47.600 160.800 48.000 165.100 ;
        RECT 50.200 160.800 50.600 164.900 ;
        RECT 51.800 160.800 52.200 165.100 ;
        RECT 53.900 160.800 54.300 163.100 ;
        RECT 55.300 160.800 55.700 163.100 ;
        RECT 57.400 160.800 57.800 165.100 ;
        RECT 59.000 160.800 59.400 164.500 ;
        RECT 60.600 160.800 61.000 165.100 ;
        RECT 62.200 160.800 62.600 164.900 ;
        RECT 64.800 160.800 65.200 165.100 ;
        RECT 67.000 160.800 67.400 164.900 ;
        RECT 69.600 160.800 70.000 165.100 ;
        RECT 71.000 160.800 71.400 165.100 ;
        RECT 73.100 160.800 73.500 163.100 ;
        RECT 74.500 160.800 74.900 163.100 ;
        RECT 76.600 160.800 77.000 165.100 ;
        RECT 78.200 160.800 78.600 165.000 ;
        RECT 81.000 160.800 81.400 163.100 ;
        RECT 82.600 160.800 83.000 163.100 ;
        RECT 85.400 160.800 85.800 165.100 ;
        RECT 87.800 160.800 88.200 164.500 ;
        RECT 89.400 160.800 89.800 165.100 ;
        RECT 92.100 160.800 92.500 163.100 ;
        RECT 94.200 160.800 94.600 165.100 ;
        RECT 95.800 160.800 96.200 164.900 ;
        RECT 98.400 160.800 98.800 165.100 ;
        RECT 99.800 160.800 100.200 165.100 ;
        RECT 101.900 160.800 102.300 163.100 ;
        RECT 103.800 160.800 104.200 164.500 ;
        RECT 105.400 160.800 105.800 165.100 ;
        RECT 107.000 160.800 107.400 165.000 ;
        RECT 109.800 160.800 110.200 163.100 ;
        RECT 111.400 160.800 111.800 163.100 ;
        RECT 114.200 160.800 114.600 165.100 ;
        RECT 116.600 160.800 117.000 164.900 ;
        RECT 119.200 160.800 119.600 165.100 ;
        RECT 121.200 160.800 121.600 165.100 ;
        RECT 123.800 160.800 124.200 164.900 ;
        RECT 126.000 160.800 126.400 165.100 ;
        RECT 128.600 160.800 129.000 164.900 ;
        RECT 130.800 160.800 131.200 165.100 ;
        RECT 133.400 160.800 133.800 164.900 ;
        RECT 135.600 160.800 136.000 165.100 ;
        RECT 138.200 160.800 138.600 164.900 ;
        RECT 142.200 160.800 142.600 165.000 ;
        RECT 145.000 160.800 145.400 163.100 ;
        RECT 146.600 160.800 147.000 163.100 ;
        RECT 149.400 160.800 149.800 165.100 ;
        RECT 151.800 160.800 152.200 163.100 ;
        RECT 152.900 160.800 153.300 163.100 ;
        RECT 155.000 160.800 155.400 165.100 ;
        RECT 155.800 160.800 156.200 163.100 ;
        RECT 157.400 160.800 157.800 163.100 ;
        RECT 159.000 160.800 159.400 165.000 ;
        RECT 161.800 160.800 162.200 163.100 ;
        RECT 163.400 160.800 163.800 163.100 ;
        RECT 166.200 160.800 166.600 165.100 ;
        RECT 167.800 160.800 168.200 163.100 ;
        RECT 169.400 160.800 169.800 163.100 ;
        RECT 170.500 160.800 170.900 163.100 ;
        RECT 172.600 160.800 173.000 165.100 ;
        RECT 174.200 160.800 174.600 162.900 ;
        RECT 175.800 160.800 176.200 163.100 ;
        RECT 176.600 160.800 177.000 163.100 ;
        RECT 178.200 160.800 178.600 163.100 ;
        RECT 179.800 160.800 180.200 164.500 ;
        RECT 181.400 160.800 181.800 165.100 ;
        RECT 182.200 160.800 182.600 165.100 ;
        RECT 184.300 160.800 184.700 163.100 ;
        RECT 186.200 160.800 186.600 165.000 ;
        RECT 189.000 160.800 189.400 163.100 ;
        RECT 190.600 160.800 191.000 163.100 ;
        RECT 193.400 160.800 193.800 165.100 ;
        RECT 197.400 160.800 197.800 164.900 ;
        RECT 200.000 160.800 200.400 165.100 ;
        RECT 202.200 160.800 202.600 164.900 ;
        RECT 204.800 160.800 205.200 165.100 ;
        RECT 207.000 160.800 207.400 165.100 ;
        RECT 209.800 160.800 210.200 163.100 ;
        RECT 211.400 160.800 211.800 163.100 ;
        RECT 214.200 160.800 214.600 165.000 ;
        RECT 215.800 160.800 216.200 163.100 ;
        RECT 217.400 160.800 217.800 163.100 ;
        RECT 218.500 160.800 218.900 163.100 ;
        RECT 220.600 160.800 221.000 165.100 ;
        RECT 221.400 160.800 221.800 163.100 ;
        RECT 223.000 160.800 223.400 163.100 ;
        RECT 223.800 160.800 224.200 165.100 ;
        RECT 225.400 160.800 225.800 165.100 ;
        RECT 227.000 160.800 227.400 165.100 ;
        RECT 228.600 160.800 229.000 165.100 ;
        RECT 230.200 160.800 230.600 165.100 ;
        RECT 0.200 160.200 231.000 160.800 ;
        RECT 0.900 157.900 1.300 160.200 ;
        RECT 3.000 155.900 3.400 160.200 ;
        RECT 3.800 157.900 4.200 160.200 ;
        RECT 5.400 157.900 5.800 160.200 ;
        RECT 7.000 156.500 7.400 160.200 ;
        RECT 8.600 155.900 9.000 160.200 ;
        RECT 9.400 155.900 9.800 160.200 ;
        RECT 11.500 157.900 11.900 160.200 ;
        RECT 13.400 156.000 13.800 160.200 ;
        RECT 16.200 157.900 16.600 160.200 ;
        RECT 17.800 157.900 18.200 160.200 ;
        RECT 20.600 155.900 21.000 160.200 ;
        RECT 23.000 156.000 23.400 160.200 ;
        RECT 25.800 157.900 26.200 160.200 ;
        RECT 27.400 157.900 27.800 160.200 ;
        RECT 30.200 155.900 30.600 160.200 ;
        RECT 32.600 156.000 33.000 160.200 ;
        RECT 35.400 157.900 35.800 160.200 ;
        RECT 37.000 157.900 37.400 160.200 ;
        RECT 39.800 155.900 40.200 160.200 ;
        RECT 43.000 155.900 43.400 160.200 ;
        RECT 45.100 157.900 45.500 160.200 ;
        RECT 46.500 157.900 46.900 160.200 ;
        RECT 48.600 155.900 49.000 160.200 ;
        RECT 50.000 155.900 50.400 160.200 ;
        RECT 52.600 156.100 53.000 160.200 ;
        RECT 55.000 156.000 55.400 160.200 ;
        RECT 57.800 157.900 58.200 160.200 ;
        RECT 59.400 157.900 59.800 160.200 ;
        RECT 62.200 155.900 62.600 160.200 ;
        RECT 63.800 155.900 64.200 160.200 ;
        RECT 65.900 157.900 66.300 160.200 ;
        RECT 67.000 157.900 67.400 160.200 ;
        RECT 68.600 157.900 69.000 160.200 ;
        RECT 69.400 157.900 69.800 160.200 ;
        RECT 71.000 155.900 71.400 160.200 ;
        RECT 72.600 156.500 73.000 160.200 ;
        RECT 75.000 156.000 75.400 160.200 ;
        RECT 77.800 157.900 78.200 160.200 ;
        RECT 79.400 157.900 79.800 160.200 ;
        RECT 82.200 155.900 82.600 160.200 ;
        RECT 83.800 155.900 84.200 160.200 ;
        RECT 85.900 157.900 86.300 160.200 ;
        RECT 89.400 156.000 89.800 160.200 ;
        RECT 92.200 157.900 92.600 160.200 ;
        RECT 93.800 157.900 94.200 160.200 ;
        RECT 96.600 155.900 97.000 160.200 ;
        RECT 98.200 157.900 98.600 160.200 ;
        RECT 99.800 157.900 100.200 160.200 ;
        RECT 100.900 157.900 101.300 160.200 ;
        RECT 103.000 155.900 103.400 160.200 ;
        RECT 103.800 157.900 104.200 160.200 ;
        RECT 105.400 157.900 105.800 160.200 ;
        RECT 107.000 156.000 107.400 160.200 ;
        RECT 109.800 157.900 110.200 160.200 ;
        RECT 111.400 157.900 111.800 160.200 ;
        RECT 114.200 155.900 114.600 160.200 ;
        RECT 116.600 156.000 117.000 160.200 ;
        RECT 119.400 157.900 119.800 160.200 ;
        RECT 121.000 157.900 121.400 160.200 ;
        RECT 123.800 155.900 124.200 160.200 ;
        RECT 125.400 155.900 125.800 160.200 ;
        RECT 127.000 156.500 127.400 160.200 ;
        RECT 128.600 157.900 129.000 160.200 ;
        RECT 130.200 157.900 130.600 160.200 ;
        RECT 131.800 156.000 132.200 160.200 ;
        RECT 134.600 157.900 135.000 160.200 ;
        RECT 136.200 157.900 136.600 160.200 ;
        RECT 139.000 155.900 139.400 160.200 ;
        RECT 142.200 157.900 142.600 160.200 ;
        RECT 143.800 157.900 144.200 160.200 ;
        RECT 145.400 157.900 145.800 160.200 ;
        RECT 146.200 155.900 146.600 160.200 ;
        RECT 148.300 157.900 148.700 160.200 ;
        RECT 150.200 156.500 150.600 160.200 ;
        RECT 152.600 155.900 153.000 160.200 ;
        RECT 154.200 156.500 154.600 160.200 ;
        RECT 155.800 157.900 156.200 160.200 ;
        RECT 157.400 157.900 157.800 160.200 ;
        RECT 158.200 157.900 158.600 160.200 ;
        RECT 159.800 157.900 160.200 160.200 ;
        RECT 161.400 155.900 161.800 160.200 ;
        RECT 164.200 157.900 164.600 160.200 ;
        RECT 165.800 157.900 166.200 160.200 ;
        RECT 168.600 156.000 169.000 160.200 ;
        RECT 170.500 157.900 170.900 160.200 ;
        RECT 172.600 155.900 173.000 160.200 ;
        RECT 174.200 156.100 174.600 160.200 ;
        RECT 176.800 155.900 177.200 160.200 ;
        RECT 178.200 157.900 178.600 160.200 ;
        RECT 179.800 157.900 180.200 160.200 ;
        RECT 180.600 155.900 181.000 160.200 ;
        RECT 182.700 157.900 183.100 160.200 ;
        RECT 183.800 157.900 184.200 160.200 ;
        RECT 185.400 157.900 185.800 160.200 ;
        RECT 187.000 155.900 187.400 160.200 ;
        RECT 189.800 157.900 190.200 160.200 ;
        RECT 191.400 157.900 191.800 160.200 ;
        RECT 194.200 156.000 194.600 160.200 ;
        RECT 197.400 157.900 197.800 160.200 ;
        RECT 199.000 157.900 199.400 160.200 ;
        RECT 200.600 156.100 201.000 160.200 ;
        RECT 203.200 155.900 203.600 160.200 ;
        RECT 204.600 155.900 205.000 160.200 ;
        RECT 206.200 156.500 206.600 160.200 ;
        RECT 207.800 155.900 208.200 160.200 ;
        RECT 209.900 157.900 210.300 160.200 ;
        RECT 211.000 157.900 211.400 160.200 ;
        RECT 212.600 157.900 213.000 160.200 ;
        RECT 213.700 157.900 214.100 160.200 ;
        RECT 215.800 155.900 216.200 160.200 ;
        RECT 217.400 155.900 217.800 160.200 ;
        RECT 220.200 157.900 220.600 160.200 ;
        RECT 221.800 157.900 222.200 160.200 ;
        RECT 224.600 156.000 225.000 160.200 ;
        RECT 226.500 157.900 226.900 160.200 ;
        RECT 228.600 155.900 229.000 160.200 ;
        RECT 1.400 140.800 1.800 145.000 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.100 ;
        RECT 10.200 140.800 10.600 145.100 ;
        RECT 12.300 140.800 12.700 143.100 ;
        RECT 13.400 140.800 13.800 143.100 ;
        RECT 15.000 140.800 15.400 143.100 ;
        RECT 15.800 140.800 16.200 143.100 ;
        RECT 17.400 140.800 17.800 143.100 ;
        RECT 18.200 140.800 18.600 143.100 ;
        RECT 19.800 140.800 20.200 143.100 ;
        RECT 20.600 140.800 21.000 145.100 ;
        RECT 22.700 140.800 23.100 143.100 ;
        RECT 23.800 140.800 24.200 143.100 ;
        RECT 25.400 140.800 25.800 143.100 ;
        RECT 27.000 140.800 27.400 145.100 ;
        RECT 30.200 140.800 30.600 145.100 ;
        RECT 31.300 140.800 31.700 143.100 ;
        RECT 33.400 140.800 33.800 145.100 ;
        RECT 35.000 140.800 35.400 144.500 ;
        RECT 36.600 140.800 37.000 145.100 ;
        RECT 39.000 140.800 39.400 145.100 ;
        RECT 41.100 140.800 41.500 143.100 ;
        RECT 42.500 140.800 42.900 143.100 ;
        RECT 44.600 140.800 45.000 145.100 ;
        RECT 45.700 140.800 46.100 143.100 ;
        RECT 47.800 140.800 48.200 145.100 ;
        RECT 48.600 140.800 49.000 145.100 ;
        RECT 50.200 140.800 50.600 144.500 ;
        RECT 52.600 140.800 53.000 144.500 ;
        RECT 54.200 140.800 54.600 145.100 ;
        RECT 55.800 140.800 56.200 145.000 ;
        RECT 58.600 140.800 59.000 143.100 ;
        RECT 60.200 140.800 60.600 143.100 ;
        RECT 63.000 140.800 63.400 145.100 ;
        RECT 64.600 140.800 65.000 145.100 ;
        RECT 66.700 140.800 67.100 143.100 ;
        RECT 68.100 140.800 68.500 143.100 ;
        RECT 70.200 140.800 70.600 145.100 ;
        RECT 71.000 140.800 71.400 145.100 ;
        RECT 73.100 140.800 73.500 143.100 ;
        RECT 75.000 140.800 75.400 144.900 ;
        RECT 77.600 140.800 78.000 145.100 ;
        RECT 79.000 140.800 79.400 145.100 ;
        RECT 80.600 140.800 81.000 145.100 ;
        RECT 82.700 140.800 83.100 145.100 ;
        RECT 84.900 140.800 85.300 143.100 ;
        RECT 87.000 140.800 87.400 145.100 ;
        RECT 90.200 140.800 90.600 142.900 ;
        RECT 91.800 140.800 92.200 143.100 ;
        RECT 92.600 140.800 93.000 143.100 ;
        RECT 94.200 140.800 94.600 142.900 ;
        RECT 95.800 140.800 96.200 145.100 ;
        RECT 97.400 140.800 97.800 145.100 ;
        RECT 98.200 140.800 98.600 143.100 ;
        RECT 99.800 140.800 100.200 142.900 ;
        RECT 103.000 140.800 103.400 145.100 ;
        RECT 103.800 140.800 104.200 143.100 ;
        RECT 105.400 140.800 105.800 142.900 ;
        RECT 107.000 140.800 107.400 145.100 ;
        RECT 108.600 140.800 109.000 144.500 ;
        RECT 110.200 140.800 110.600 145.100 ;
        RECT 114.200 140.800 114.600 145.100 ;
        RECT 116.100 140.800 116.500 145.100 ;
        RECT 118.200 140.800 118.600 145.100 ;
        RECT 120.300 140.800 120.700 143.100 ;
        RECT 121.400 140.800 121.800 143.100 ;
        RECT 123.000 140.800 123.400 143.100 ;
        RECT 123.800 140.800 124.200 143.100 ;
        RECT 125.400 140.800 125.800 143.100 ;
        RECT 126.200 140.800 126.600 143.100 ;
        RECT 127.800 140.800 128.200 143.100 ;
        RECT 128.600 140.800 129.000 145.100 ;
        RECT 130.700 140.800 131.100 143.100 ;
        RECT 131.800 140.800 132.200 143.100 ;
        RECT 133.700 140.800 134.100 143.100 ;
        RECT 135.800 140.800 136.200 145.100 ;
        RECT 136.600 140.800 137.000 143.100 ;
        RECT 138.200 140.800 138.600 143.100 ;
        RECT 140.600 140.800 141.000 145.100 ;
        RECT 142.700 140.800 143.100 143.100 ;
        RECT 143.800 140.800 144.200 143.100 ;
        RECT 145.400 140.800 145.800 143.100 ;
        RECT 147.000 140.800 147.400 144.500 ;
        RECT 150.200 140.800 150.600 143.100 ;
        RECT 151.800 140.800 152.200 142.900 ;
        RECT 154.200 140.800 154.600 143.100 ;
        RECT 155.600 140.800 156.000 145.100 ;
        RECT 158.200 140.800 158.600 144.900 ;
        RECT 160.400 140.800 160.800 145.100 ;
        RECT 163.000 140.800 163.400 144.900 ;
        RECT 165.400 140.800 165.800 145.100 ;
        RECT 168.200 140.800 168.600 143.100 ;
        RECT 169.800 140.800 170.200 143.100 ;
        RECT 172.600 140.800 173.000 145.000 ;
        RECT 174.200 140.800 174.600 145.100 ;
        RECT 176.300 140.800 176.700 143.100 ;
        RECT 177.400 140.800 177.800 143.100 ;
        RECT 179.000 140.800 179.400 143.100 ;
        RECT 180.600 140.800 181.000 145.100 ;
        RECT 183.400 140.800 183.800 143.100 ;
        RECT 185.000 140.800 185.400 143.100 ;
        RECT 187.800 140.800 188.200 145.000 ;
        RECT 189.400 140.800 189.800 145.100 ;
        RECT 191.500 140.800 191.900 143.100 ;
        RECT 194.200 140.800 194.600 143.100 ;
        RECT 195.800 140.800 196.200 143.100 ;
        RECT 197.400 140.800 197.800 145.000 ;
        RECT 200.200 140.800 200.600 143.100 ;
        RECT 201.800 140.800 202.200 143.100 ;
        RECT 204.600 140.800 205.000 145.100 ;
        RECT 207.000 140.800 207.400 143.100 ;
        RECT 208.600 140.800 209.000 145.000 ;
        RECT 211.400 140.800 211.800 143.100 ;
        RECT 213.000 140.800 213.400 143.100 ;
        RECT 215.800 140.800 216.200 145.100 ;
        RECT 217.400 140.800 217.800 145.100 ;
        RECT 219.500 140.800 219.900 143.100 ;
        RECT 221.400 140.800 221.800 145.000 ;
        RECT 224.200 140.800 224.600 143.100 ;
        RECT 225.800 140.800 226.200 143.100 ;
        RECT 228.600 140.800 229.000 145.100 ;
        RECT 0.200 140.200 231.000 140.800 ;
        RECT 1.400 136.000 1.800 140.200 ;
        RECT 4.200 137.900 4.600 140.200 ;
        RECT 5.800 137.900 6.200 140.200 ;
        RECT 8.600 135.900 9.000 140.200 ;
        RECT 10.200 137.900 10.600 140.200 ;
        RECT 11.800 137.900 12.200 140.200 ;
        RECT 12.900 137.900 13.300 140.200 ;
        RECT 15.000 135.900 15.400 140.200 ;
        RECT 16.600 136.000 17.000 140.200 ;
        RECT 19.400 137.900 19.800 140.200 ;
        RECT 21.000 137.900 21.400 140.200 ;
        RECT 23.800 135.900 24.200 140.200 ;
        RECT 25.400 135.900 25.800 140.200 ;
        RECT 27.500 137.900 27.900 140.200 ;
        RECT 29.400 136.000 29.800 140.200 ;
        RECT 32.200 137.900 32.600 140.200 ;
        RECT 33.800 137.900 34.200 140.200 ;
        RECT 36.600 135.900 37.000 140.200 ;
        RECT 39.800 135.900 40.200 140.200 ;
        RECT 41.900 137.900 42.300 140.200 ;
        RECT 43.300 137.900 43.700 140.200 ;
        RECT 45.400 135.900 45.800 140.200 ;
        RECT 46.200 137.900 46.600 140.200 ;
        RECT 47.800 137.900 48.200 140.200 ;
        RECT 48.600 135.900 49.000 140.200 ;
        RECT 50.200 136.500 50.600 140.200 ;
        RECT 52.600 136.000 53.000 140.200 ;
        RECT 55.400 137.900 55.800 140.200 ;
        RECT 57.000 137.900 57.400 140.200 ;
        RECT 59.800 135.900 60.200 140.200 ;
        RECT 61.400 137.900 61.800 140.200 ;
        RECT 63.000 137.900 63.400 140.200 ;
        RECT 64.600 136.000 65.000 140.200 ;
        RECT 67.400 137.900 67.800 140.200 ;
        RECT 69.000 137.900 69.400 140.200 ;
        RECT 71.800 135.900 72.200 140.200 ;
        RECT 73.700 137.900 74.100 140.200 ;
        RECT 75.800 135.900 76.200 140.200 ;
        RECT 76.600 137.900 77.000 140.200 ;
        RECT 78.200 137.900 78.600 140.200 ;
        RECT 79.000 137.900 79.400 140.200 ;
        RECT 80.600 138.100 81.000 140.200 ;
        RECT 82.200 135.900 82.600 140.200 ;
        RECT 84.300 137.900 84.700 140.200 ;
        RECT 87.800 136.000 88.200 140.200 ;
        RECT 90.600 137.900 91.000 140.200 ;
        RECT 92.200 137.900 92.600 140.200 ;
        RECT 95.000 135.900 95.400 140.200 ;
        RECT 96.600 135.900 97.000 140.200 ;
        RECT 99.000 135.900 99.400 140.200 ;
        RECT 100.600 136.500 101.000 140.200 ;
        RECT 102.200 137.900 102.600 140.200 ;
        RECT 103.800 138.100 104.200 140.200 ;
        RECT 105.400 137.900 105.800 140.200 ;
        RECT 107.000 138.100 107.400 140.200 ;
        RECT 108.600 135.900 109.000 140.200 ;
        RECT 110.200 136.500 110.600 140.200 ;
        RECT 112.600 138.100 113.000 140.200 ;
        RECT 114.200 137.900 114.600 140.200 ;
        RECT 115.000 137.900 115.400 140.200 ;
        RECT 116.600 138.100 117.000 140.200 ;
        RECT 118.200 137.900 118.600 140.200 ;
        RECT 119.800 138.100 120.200 140.200 ;
        RECT 122.200 138.100 122.600 140.200 ;
        RECT 123.800 137.900 124.200 140.200 ;
        RECT 125.400 138.100 125.800 140.200 ;
        RECT 127.000 137.900 127.400 140.200 ;
        RECT 127.800 135.900 128.200 140.200 ;
        RECT 130.200 135.900 130.600 140.200 ;
        RECT 131.800 136.500 132.200 140.200 ;
        RECT 133.400 137.900 133.800 140.200 ;
        RECT 135.000 137.900 135.400 140.200 ;
        RECT 135.800 135.900 136.200 140.200 ;
        RECT 139.000 135.900 139.400 140.200 ;
        RECT 141.700 137.900 142.100 140.200 ;
        RECT 143.800 135.900 144.200 140.200 ;
        RECT 144.600 135.900 145.000 140.200 ;
        RECT 146.700 137.900 147.100 140.200 ;
        RECT 148.600 137.900 149.000 140.200 ;
        RECT 149.400 135.900 149.800 140.200 ;
        RECT 151.000 135.900 151.400 140.200 ;
        RECT 152.600 135.900 153.000 140.200 ;
        RECT 155.000 135.900 155.400 140.200 ;
        RECT 156.100 137.900 156.500 140.200 ;
        RECT 158.200 135.900 158.600 140.200 ;
        RECT 159.000 137.900 159.400 140.200 ;
        RECT 160.600 137.900 161.000 140.200 ;
        RECT 161.400 137.900 161.800 140.200 ;
        RECT 163.000 137.900 163.400 140.200 ;
        RECT 163.800 137.900 164.200 140.200 ;
        RECT 165.400 138.100 165.800 140.200 ;
        RECT 167.300 137.900 167.700 140.200 ;
        RECT 169.400 135.900 169.800 140.200 ;
        RECT 170.200 135.900 170.600 140.200 ;
        RECT 172.300 137.900 172.700 140.200 ;
        RECT 173.400 135.900 173.800 140.200 ;
        RECT 175.500 137.900 175.900 140.200 ;
        RECT 176.600 137.900 177.000 140.200 ;
        RECT 178.200 137.900 178.600 140.200 ;
        RECT 179.000 137.900 179.400 140.200 ;
        RECT 180.600 137.900 181.000 140.200 ;
        RECT 181.700 137.900 182.100 140.200 ;
        RECT 183.800 135.900 184.200 140.200 ;
        RECT 184.600 137.900 185.000 140.200 ;
        RECT 186.200 137.900 186.600 140.200 ;
        RECT 189.400 135.900 189.800 140.200 ;
        RECT 192.200 137.900 192.600 140.200 ;
        RECT 193.800 137.900 194.200 140.200 ;
        RECT 196.600 136.000 197.000 140.200 ;
        RECT 198.500 137.900 198.900 140.200 ;
        RECT 200.600 135.900 201.000 140.200 ;
        RECT 202.200 137.900 202.600 140.200 ;
        RECT 203.000 137.900 203.400 140.200 ;
        RECT 204.600 137.900 205.000 140.200 ;
        RECT 205.700 137.900 206.100 140.200 ;
        RECT 207.800 135.900 208.200 140.200 ;
        RECT 209.400 135.900 209.800 140.200 ;
        RECT 212.200 137.900 212.600 140.200 ;
        RECT 213.800 137.900 214.200 140.200 ;
        RECT 216.600 136.000 217.000 140.200 ;
        RECT 219.000 136.000 219.400 140.200 ;
        RECT 221.800 137.900 222.200 140.200 ;
        RECT 223.400 137.900 223.800 140.200 ;
        RECT 226.200 135.900 226.600 140.200 ;
        RECT 228.600 136.500 229.000 140.200 ;
        RECT 0.900 120.800 1.300 123.100 ;
        RECT 3.000 120.800 3.400 125.100 ;
        RECT 4.600 120.800 5.000 125.100 ;
        RECT 7.400 120.800 7.800 123.100 ;
        RECT 9.000 120.800 9.400 123.100 ;
        RECT 11.800 120.800 12.200 125.000 ;
        RECT 13.400 120.800 13.800 123.100 ;
        RECT 15.800 120.800 16.200 125.000 ;
        RECT 18.600 120.800 19.000 123.100 ;
        RECT 20.200 120.800 20.600 123.100 ;
        RECT 23.000 120.800 23.400 125.100 ;
        RECT 24.600 120.800 25.000 123.100 ;
        RECT 26.200 120.800 26.600 125.100 ;
        RECT 28.300 120.800 28.700 123.100 ;
        RECT 29.700 120.800 30.100 123.100 ;
        RECT 31.800 120.800 32.200 125.100 ;
        RECT 33.400 120.800 33.800 125.000 ;
        RECT 36.200 120.800 36.600 123.100 ;
        RECT 37.800 120.800 38.200 123.100 ;
        RECT 40.600 120.800 41.000 125.100 ;
        RECT 44.600 120.800 45.000 123.100 ;
        RECT 45.700 120.800 46.100 123.100 ;
        RECT 47.800 120.800 48.200 125.100 ;
        RECT 48.600 120.800 49.000 125.100 ;
        RECT 50.200 120.800 50.600 125.100 ;
        RECT 51.000 120.800 51.400 125.100 ;
        RECT 53.100 120.800 53.500 123.100 ;
        RECT 54.200 120.800 54.600 123.100 ;
        RECT 55.800 120.800 56.200 123.100 ;
        RECT 56.600 120.800 57.000 123.100 ;
        RECT 58.200 120.800 58.600 125.100 ;
        RECT 60.300 120.800 60.700 123.100 ;
        RECT 61.400 120.800 61.800 123.100 ;
        RECT 63.000 120.800 63.400 123.100 ;
        RECT 63.800 120.800 64.200 123.100 ;
        RECT 66.200 120.800 66.600 125.000 ;
        RECT 69.000 120.800 69.400 123.100 ;
        RECT 70.600 120.800 71.000 123.100 ;
        RECT 73.400 120.800 73.800 125.100 ;
        RECT 75.000 120.800 75.400 123.100 ;
        RECT 76.600 120.800 77.000 123.100 ;
        RECT 78.200 120.800 78.600 125.100 ;
        RECT 80.300 120.800 80.700 123.100 ;
        RECT 81.400 120.800 81.800 123.100 ;
        RECT 83.000 120.800 83.400 123.100 ;
        RECT 84.600 120.800 85.000 125.000 ;
        RECT 87.400 120.800 87.800 123.100 ;
        RECT 89.000 120.800 89.400 123.100 ;
        RECT 91.800 120.800 92.200 125.100 ;
        RECT 95.000 120.800 95.400 123.100 ;
        RECT 96.600 120.800 97.000 123.100 ;
        RECT 99.000 120.800 99.400 125.100 ;
        RECT 100.600 120.800 101.000 122.900 ;
        RECT 102.200 120.800 102.600 123.100 ;
        RECT 103.800 120.800 104.200 122.900 ;
        RECT 105.400 120.800 105.800 123.100 ;
        RECT 106.200 120.800 106.600 125.100 ;
        RECT 109.400 120.800 109.800 125.100 ;
        RECT 111.000 120.800 111.400 122.900 ;
        RECT 112.600 120.800 113.000 123.100 ;
        RECT 114.200 120.800 114.600 122.900 ;
        RECT 115.800 120.800 116.200 123.100 ;
        RECT 116.600 120.800 117.000 125.100 ;
        RECT 119.000 120.800 119.400 123.100 ;
        RECT 120.600 120.800 121.000 122.900 ;
        RECT 122.200 120.800 122.600 125.100 ;
        RECT 123.800 120.800 124.200 124.500 ;
        RECT 126.200 120.800 126.600 125.000 ;
        RECT 129.000 120.800 129.400 123.100 ;
        RECT 130.600 120.800 131.000 123.100 ;
        RECT 133.400 120.800 133.800 125.100 ;
        RECT 135.300 120.800 135.700 123.100 ;
        RECT 137.400 120.800 137.800 125.100 ;
        RECT 138.200 120.800 138.600 123.100 ;
        RECT 139.800 120.800 140.200 123.100 ;
        RECT 142.500 120.800 142.900 123.100 ;
        RECT 144.600 120.800 145.000 125.100 ;
        RECT 145.400 120.800 145.800 123.100 ;
        RECT 147.000 120.800 147.400 123.100 ;
        RECT 148.100 120.800 148.500 123.100 ;
        RECT 150.200 120.800 150.600 125.100 ;
        RECT 151.800 120.800 152.200 123.100 ;
        RECT 153.400 120.800 153.800 125.100 ;
        RECT 156.200 120.800 156.600 123.100 ;
        RECT 157.800 120.800 158.200 123.100 ;
        RECT 160.600 120.800 161.000 125.000 ;
        RECT 162.500 120.800 162.900 123.100 ;
        RECT 164.600 120.800 165.000 125.100 ;
        RECT 166.200 120.800 166.600 122.900 ;
        RECT 167.800 120.800 168.200 123.100 ;
        RECT 168.600 120.800 169.000 123.100 ;
        RECT 170.200 120.800 170.600 123.100 ;
        RECT 171.000 120.800 171.400 125.100 ;
        RECT 172.600 120.800 173.000 124.500 ;
        RECT 174.200 120.800 174.600 125.100 ;
        RECT 176.300 120.800 176.700 123.100 ;
        RECT 177.400 120.800 177.800 123.100 ;
        RECT 179.000 120.800 179.400 123.100 ;
        RECT 180.600 120.800 181.000 125.100 ;
        RECT 183.400 120.800 183.800 123.100 ;
        RECT 185.000 120.800 185.400 123.100 ;
        RECT 187.800 120.800 188.200 125.000 ;
        RECT 189.700 120.800 190.100 123.100 ;
        RECT 191.800 120.800 192.200 125.100 ;
        RECT 195.000 120.800 195.400 124.500 ;
        RECT 196.600 120.800 197.000 125.100 ;
        RECT 198.200 120.800 198.600 124.900 ;
        RECT 200.800 120.800 201.200 125.100 ;
        RECT 203.000 120.800 203.400 124.500 ;
        RECT 205.700 120.800 206.100 123.100 ;
        RECT 207.800 120.800 208.200 125.100 ;
        RECT 209.400 120.800 209.800 124.900 ;
        RECT 212.000 120.800 212.400 125.100 ;
        RECT 213.400 120.800 213.800 123.100 ;
        RECT 215.000 120.800 215.400 123.100 ;
        RECT 216.100 120.800 216.500 123.100 ;
        RECT 218.200 120.800 218.600 125.100 ;
        RECT 219.800 120.800 220.200 125.100 ;
        RECT 222.600 120.800 223.000 123.100 ;
        RECT 224.200 120.800 224.600 123.100 ;
        RECT 227.000 120.800 227.400 125.000 ;
        RECT 229.400 120.800 229.800 124.500 ;
        RECT 0.200 120.200 231.000 120.800 ;
        RECT 0.600 115.900 1.000 120.200 ;
        RECT 2.200 115.900 2.600 120.200 ;
        RECT 3.800 115.900 4.200 120.200 ;
        RECT 5.400 116.000 5.800 120.200 ;
        RECT 8.200 117.900 8.600 120.200 ;
        RECT 9.800 117.900 10.200 120.200 ;
        RECT 12.600 115.900 13.000 120.200 ;
        RECT 14.200 115.900 14.600 120.200 ;
        RECT 16.300 117.900 16.700 120.200 ;
        RECT 17.700 117.900 18.100 120.200 ;
        RECT 19.800 115.900 20.200 120.200 ;
        RECT 20.600 117.900 21.000 120.200 ;
        RECT 22.200 115.900 22.600 120.200 ;
        RECT 25.400 115.900 25.800 120.200 ;
        RECT 26.200 115.900 26.600 120.200 ;
        RECT 29.400 115.900 29.800 120.200 ;
        RECT 31.000 117.900 31.400 120.200 ;
        RECT 31.800 115.900 32.200 120.200 ;
        RECT 33.400 116.500 33.800 120.200 ;
        RECT 35.000 115.900 35.400 120.200 ;
        RECT 37.100 117.900 37.500 120.200 ;
        RECT 39.800 115.900 40.200 120.200 ;
        RECT 41.900 117.900 42.300 120.200 ;
        RECT 43.800 116.500 44.200 120.200 ;
        RECT 45.400 115.900 45.800 120.200 ;
        RECT 46.200 115.900 46.600 120.200 ;
        RECT 48.300 117.900 48.700 120.200 ;
        RECT 49.700 117.900 50.100 120.200 ;
        RECT 51.800 115.900 52.200 120.200 ;
        RECT 53.400 115.900 53.800 120.200 ;
        RECT 56.200 117.900 56.600 120.200 ;
        RECT 57.800 117.900 58.200 120.200 ;
        RECT 60.600 116.000 61.000 120.200 ;
        RECT 63.300 115.900 63.700 120.200 ;
        RECT 66.200 116.500 66.600 120.200 ;
        RECT 67.800 115.900 68.200 120.200 ;
        RECT 68.600 115.900 69.000 120.200 ;
        RECT 70.700 117.900 71.100 120.200 ;
        RECT 72.100 117.900 72.500 120.200 ;
        RECT 74.200 115.900 74.600 120.200 ;
        RECT 75.000 115.900 75.400 120.200 ;
        RECT 78.200 115.900 78.600 120.200 ;
        RECT 79.800 117.900 80.200 120.200 ;
        RECT 80.600 115.900 81.000 120.200 ;
        RECT 82.200 115.900 82.600 120.200 ;
        RECT 83.800 115.900 84.200 120.200 ;
        RECT 86.600 117.900 87.000 120.200 ;
        RECT 88.200 117.900 88.600 120.200 ;
        RECT 91.000 116.000 91.400 120.200 ;
        RECT 94.200 117.900 94.600 120.200 ;
        RECT 95.800 117.900 96.200 120.200 ;
        RECT 96.900 117.900 97.300 120.200 ;
        RECT 99.000 115.900 99.400 120.200 ;
        RECT 99.800 117.900 100.200 120.200 ;
        RECT 101.400 117.900 101.800 120.200 ;
        RECT 102.200 117.900 102.600 120.200 ;
        RECT 103.800 117.900 104.200 120.200 ;
        RECT 104.600 115.900 105.000 120.200 ;
        RECT 106.700 117.900 107.100 120.200 ;
        RECT 107.800 117.900 108.200 120.200 ;
        RECT 109.400 117.900 109.800 120.200 ;
        RECT 111.000 117.900 111.400 120.200 ;
        RECT 111.800 117.900 112.200 120.200 ;
        RECT 113.400 117.900 113.800 120.200 ;
        RECT 115.800 115.900 116.200 120.200 ;
        RECT 117.400 118.100 117.800 120.200 ;
        RECT 119.000 117.900 119.400 120.200 ;
        RECT 119.800 115.900 120.200 120.200 ;
        RECT 122.200 117.900 122.600 120.200 ;
        RECT 123.800 118.100 124.200 120.200 ;
        RECT 125.400 117.900 125.800 120.200 ;
        RECT 127.000 117.900 127.400 120.200 ;
        RECT 128.600 116.500 129.000 120.200 ;
        RECT 130.200 115.900 130.600 120.200 ;
        RECT 131.800 115.900 132.200 120.200 ;
        RECT 134.600 117.900 135.000 120.200 ;
        RECT 136.200 117.900 136.600 120.200 ;
        RECT 139.000 116.000 139.400 120.200 ;
        RECT 142.200 117.900 142.600 120.200 ;
        RECT 143.800 117.900 144.200 120.200 ;
        RECT 144.900 117.900 145.300 120.200 ;
        RECT 147.000 115.900 147.400 120.200 ;
        RECT 147.800 117.900 148.200 120.200 ;
        RECT 149.400 115.900 149.800 120.200 ;
        RECT 152.600 115.900 153.000 120.200 ;
        RECT 153.400 117.900 153.800 120.200 ;
        RECT 155.000 117.900 155.400 120.200 ;
        RECT 156.100 117.900 156.500 120.200 ;
        RECT 158.200 115.900 158.600 120.200 ;
        RECT 159.000 117.900 159.400 120.200 ;
        RECT 160.600 117.900 161.000 120.200 ;
        RECT 161.400 117.900 161.800 120.200 ;
        RECT 163.000 117.900 163.400 120.200 ;
        RECT 164.600 116.500 165.000 120.200 ;
        RECT 167.800 116.500 168.200 120.200 ;
        RECT 170.200 115.900 170.600 120.200 ;
        RECT 171.800 116.500 172.200 120.200 ;
        RECT 173.700 117.900 174.100 120.200 ;
        RECT 175.800 115.900 176.200 120.200 ;
        RECT 178.200 116.500 178.600 120.200 ;
        RECT 179.800 115.900 180.200 120.200 ;
        RECT 181.900 117.900 182.300 120.200 ;
        RECT 183.000 117.900 183.400 120.200 ;
        RECT 184.600 117.900 185.000 120.200 ;
        RECT 186.200 116.500 186.600 120.200 ;
        RECT 188.900 117.900 189.300 120.200 ;
        RECT 191.000 115.900 191.400 120.200 ;
        RECT 194.200 116.000 194.600 120.200 ;
        RECT 197.000 117.900 197.400 120.200 ;
        RECT 198.600 117.900 199.000 120.200 ;
        RECT 201.400 115.900 201.800 120.200 ;
        RECT 203.600 115.900 204.000 120.200 ;
        RECT 206.200 116.100 206.600 120.200 ;
        RECT 207.800 117.900 208.200 120.200 ;
        RECT 209.400 117.900 209.800 120.200 ;
        RECT 211.000 115.900 211.400 120.200 ;
        RECT 213.800 117.900 214.200 120.200 ;
        RECT 215.400 117.900 215.800 120.200 ;
        RECT 218.200 116.000 218.600 120.200 ;
        RECT 220.600 116.000 221.000 120.200 ;
        RECT 223.400 117.900 223.800 120.200 ;
        RECT 225.000 117.900 225.400 120.200 ;
        RECT 227.800 115.900 228.200 120.200 ;
        RECT 0.600 100.800 1.000 103.100 ;
        RECT 2.200 100.800 2.600 103.100 ;
        RECT 3.000 100.800 3.400 103.100 ;
        RECT 4.600 100.800 5.000 103.100 ;
        RECT 6.200 100.800 6.600 103.100 ;
        RECT 7.300 100.800 7.700 103.100 ;
        RECT 9.400 100.800 9.800 105.100 ;
        RECT 11.000 100.800 11.400 105.000 ;
        RECT 13.800 100.800 14.200 103.100 ;
        RECT 15.400 100.800 15.800 103.100 ;
        RECT 18.200 100.800 18.600 105.100 ;
        RECT 19.800 100.800 20.200 105.100 ;
        RECT 21.900 100.800 22.300 103.100 ;
        RECT 23.000 100.800 23.400 103.100 ;
        RECT 24.600 100.800 25.000 103.100 ;
        RECT 25.400 100.800 25.800 105.100 ;
        RECT 27.500 100.800 27.900 103.100 ;
        RECT 28.600 100.800 29.000 105.100 ;
        RECT 30.200 100.800 30.600 104.500 ;
        RECT 31.800 100.800 32.200 103.100 ;
        RECT 35.800 100.800 36.200 105.000 ;
        RECT 38.600 100.800 39.000 103.100 ;
        RECT 40.200 100.800 40.600 103.100 ;
        RECT 43.000 100.800 43.400 105.100 ;
        RECT 45.400 100.800 45.800 104.500 ;
        RECT 47.000 100.800 47.400 105.100 ;
        RECT 48.600 100.800 49.000 105.000 ;
        RECT 51.400 100.800 51.800 103.100 ;
        RECT 53.000 100.800 53.400 103.100 ;
        RECT 55.800 100.800 56.200 105.100 ;
        RECT 57.400 100.800 57.800 103.100 ;
        RECT 59.000 100.800 59.400 103.100 ;
        RECT 60.600 100.800 61.000 103.100 ;
        RECT 61.700 100.800 62.100 103.100 ;
        RECT 63.800 100.800 64.200 105.100 ;
        RECT 65.400 100.800 65.800 105.000 ;
        RECT 68.200 100.800 68.600 103.100 ;
        RECT 69.800 100.800 70.200 103.100 ;
        RECT 72.600 100.800 73.000 105.100 ;
        RECT 75.000 100.800 75.400 104.500 ;
        RECT 76.600 100.800 77.000 105.100 ;
        RECT 77.400 100.800 77.800 105.100 ;
        RECT 79.500 100.800 79.900 103.100 ;
        RECT 80.600 100.800 81.000 105.100 ;
        RECT 82.700 100.800 83.100 103.100 ;
        RECT 84.100 100.800 84.500 103.100 ;
        RECT 86.200 100.800 86.600 105.100 ;
        RECT 89.400 100.800 89.800 105.000 ;
        RECT 92.200 100.800 92.600 103.100 ;
        RECT 93.800 100.800 94.200 103.100 ;
        RECT 96.600 100.800 97.000 105.100 ;
        RECT 98.200 100.800 98.600 105.100 ;
        RECT 100.300 100.800 100.700 103.100 ;
        RECT 101.400 100.800 101.800 103.100 ;
        RECT 103.000 100.800 103.400 103.100 ;
        RECT 104.600 100.800 105.000 105.000 ;
        RECT 107.400 100.800 107.800 103.100 ;
        RECT 109.000 100.800 109.400 103.100 ;
        RECT 111.800 100.800 112.200 105.100 ;
        RECT 113.400 100.800 113.800 105.100 ;
        RECT 115.000 100.800 115.400 105.100 ;
        RECT 117.400 100.800 117.800 105.100 ;
        RECT 118.200 100.800 118.600 105.100 ;
        RECT 119.800 100.800 120.200 104.500 ;
        RECT 122.200 100.800 122.600 104.500 ;
        RECT 123.800 100.800 124.200 105.100 ;
        RECT 124.900 100.800 125.300 103.100 ;
        RECT 127.000 100.800 127.400 105.100 ;
        RECT 128.600 100.800 129.000 105.000 ;
        RECT 131.400 100.800 131.800 103.100 ;
        RECT 133.000 100.800 133.400 103.100 ;
        RECT 135.800 100.800 136.200 105.100 ;
        RECT 137.400 100.800 137.800 105.100 ;
        RECT 139.500 100.800 139.900 103.100 ;
        RECT 142.200 100.800 142.600 103.100 ;
        RECT 143.800 100.800 144.200 103.100 ;
        RECT 144.600 100.800 145.000 103.100 ;
        RECT 146.500 100.800 146.900 103.100 ;
        RECT 148.600 100.800 149.000 105.100 ;
        RECT 149.400 100.800 149.800 105.100 ;
        RECT 151.500 100.800 151.900 103.100 ;
        RECT 152.600 100.800 153.000 103.100 ;
        RECT 154.200 100.800 154.600 103.100 ;
        RECT 156.600 100.800 157.000 105.100 ;
        RECT 157.700 100.800 158.100 103.100 ;
        RECT 159.800 100.800 160.200 105.100 ;
        RECT 161.400 100.800 161.800 104.500 ;
        RECT 164.100 100.800 164.500 103.100 ;
        RECT 166.200 100.800 166.600 105.100 ;
        RECT 167.800 100.800 168.200 103.100 ;
        RECT 169.400 100.800 169.800 105.100 ;
        RECT 172.200 100.800 172.600 103.100 ;
        RECT 173.800 100.800 174.200 103.100 ;
        RECT 176.600 100.800 177.000 105.000 ;
        RECT 178.200 100.800 178.600 103.100 ;
        RECT 179.800 100.800 180.200 103.100 ;
        RECT 180.900 100.800 181.300 103.100 ;
        RECT 183.000 100.800 183.400 105.100 ;
        RECT 183.800 100.800 184.200 103.100 ;
        RECT 185.400 100.800 185.800 103.100 ;
        RECT 186.200 100.800 186.600 105.100 ;
        RECT 188.300 100.800 188.700 103.100 ;
        RECT 189.400 100.800 189.800 103.100 ;
        RECT 191.000 100.800 191.400 103.100 ;
        RECT 194.200 100.800 194.600 105.100 ;
        RECT 197.000 100.800 197.400 103.100 ;
        RECT 198.600 100.800 199.000 103.100 ;
        RECT 201.400 100.800 201.800 105.000 ;
        RECT 203.000 100.800 203.400 105.100 ;
        RECT 204.600 100.800 205.000 105.100 ;
        RECT 206.200 100.800 206.600 105.100 ;
        RECT 207.000 100.800 207.400 105.100 ;
        RECT 209.100 100.800 209.500 103.100 ;
        RECT 211.000 100.800 211.400 105.100 ;
        RECT 213.800 100.800 214.200 103.100 ;
        RECT 215.400 100.800 215.800 103.100 ;
        RECT 218.200 100.800 218.600 105.000 ;
        RECT 220.600 100.800 221.000 105.000 ;
        RECT 223.400 100.800 223.800 103.100 ;
        RECT 225.000 100.800 225.400 103.100 ;
        RECT 227.800 100.800 228.200 105.100 ;
        RECT 0.200 100.200 231.000 100.800 ;
        RECT 1.400 95.900 1.800 100.200 ;
        RECT 4.200 97.900 4.600 100.200 ;
        RECT 5.800 97.900 6.200 100.200 ;
        RECT 8.600 96.000 9.000 100.200 ;
        RECT 10.200 97.900 10.600 100.200 ;
        RECT 11.800 97.900 12.200 100.200 ;
        RECT 12.900 97.900 13.300 100.200 ;
        RECT 15.000 95.900 15.400 100.200 ;
        RECT 15.800 95.900 16.200 100.200 ;
        RECT 17.900 97.900 18.300 100.200 ;
        RECT 19.000 97.900 19.400 100.200 ;
        RECT 20.600 97.900 21.000 100.200 ;
        RECT 22.200 96.000 22.600 100.200 ;
        RECT 25.000 97.900 25.400 100.200 ;
        RECT 26.600 97.900 27.000 100.200 ;
        RECT 29.400 95.900 29.800 100.200 ;
        RECT 31.000 97.900 31.400 100.200 ;
        RECT 32.600 97.900 33.000 100.200 ;
        RECT 34.200 97.900 34.600 100.200 ;
        RECT 35.000 97.900 35.400 100.200 ;
        RECT 38.200 95.900 38.600 100.200 ;
        RECT 40.300 97.900 40.700 100.200 ;
        RECT 41.400 97.900 41.800 100.200 ;
        RECT 43.000 95.900 43.400 100.200 ;
        RECT 46.200 95.900 46.600 100.200 ;
        RECT 47.000 95.900 47.400 100.200 ;
        RECT 49.100 97.900 49.500 100.200 ;
        RECT 50.200 97.900 50.600 100.200 ;
        RECT 51.800 97.900 52.200 100.200 ;
        RECT 52.600 97.900 53.000 100.200 ;
        RECT 54.200 97.900 54.600 100.200 ;
        RECT 55.000 95.900 55.400 100.200 ;
        RECT 57.100 97.900 57.500 100.200 ;
        RECT 59.000 96.000 59.400 100.200 ;
        RECT 61.800 97.900 62.200 100.200 ;
        RECT 63.400 97.900 63.800 100.200 ;
        RECT 66.200 95.900 66.600 100.200 ;
        RECT 67.800 97.900 68.200 100.200 ;
        RECT 69.400 97.900 69.800 100.200 ;
        RECT 70.500 97.900 70.900 100.200 ;
        RECT 72.600 95.900 73.000 100.200 ;
        RECT 73.400 95.900 73.800 100.200 ;
        RECT 75.000 96.500 75.400 100.200 ;
        RECT 76.600 95.900 77.000 100.200 ;
        RECT 78.700 97.900 79.100 100.200 ;
        RECT 80.600 95.900 81.000 100.200 ;
        RECT 83.400 97.900 83.800 100.200 ;
        RECT 85.000 97.900 85.400 100.200 ;
        RECT 87.800 96.000 88.200 100.200 ;
        RECT 91.000 97.900 91.400 100.200 ;
        RECT 92.600 97.900 93.000 100.200 ;
        RECT 94.200 98.100 94.600 100.200 ;
        RECT 95.800 97.900 96.200 100.200 ;
        RECT 96.600 97.900 97.000 100.200 ;
        RECT 98.200 97.900 98.600 100.200 ;
        RECT 99.000 97.900 99.400 100.200 ;
        RECT 100.600 97.900 101.000 100.200 ;
        RECT 101.700 97.900 102.100 100.200 ;
        RECT 103.800 95.900 104.200 100.200 ;
        RECT 104.600 97.900 105.000 100.200 ;
        RECT 106.200 97.900 106.600 100.200 ;
        RECT 107.000 97.900 107.400 100.200 ;
        RECT 108.600 97.900 109.000 100.200 ;
        RECT 110.000 95.900 110.400 100.200 ;
        RECT 112.600 96.100 113.000 100.200 ;
        RECT 114.200 97.900 114.600 100.200 ;
        RECT 115.800 97.900 116.200 100.200 ;
        RECT 116.600 95.900 117.000 100.200 ;
        RECT 118.200 96.500 118.600 100.200 ;
        RECT 119.800 95.900 120.200 100.200 ;
        RECT 121.400 96.500 121.800 100.200 ;
        RECT 123.000 97.900 123.400 100.200 ;
        RECT 124.600 97.900 125.000 100.200 ;
        RECT 127.800 96.500 128.200 100.200 ;
        RECT 130.200 97.900 130.600 100.200 ;
        RECT 131.000 97.900 131.400 100.200 ;
        RECT 132.600 97.900 133.000 100.200 ;
        RECT 133.700 97.900 134.100 100.200 ;
        RECT 135.800 95.900 136.200 100.200 ;
        RECT 139.000 96.000 139.400 100.200 ;
        RECT 141.800 97.900 142.200 100.200 ;
        RECT 143.400 97.900 143.800 100.200 ;
        RECT 146.200 95.900 146.600 100.200 ;
        RECT 148.100 97.900 148.500 100.200 ;
        RECT 150.200 95.900 150.600 100.200 ;
        RECT 151.300 97.900 151.700 100.200 ;
        RECT 153.400 95.900 153.800 100.200 ;
        RECT 154.200 95.900 154.600 100.200 ;
        RECT 155.800 96.500 156.200 100.200 ;
        RECT 158.200 96.500 158.600 100.200 ;
        RECT 159.800 95.900 160.200 100.200 ;
        RECT 161.400 96.000 161.800 100.200 ;
        RECT 164.200 97.900 164.600 100.200 ;
        RECT 165.800 97.900 166.200 100.200 ;
        RECT 168.600 95.900 169.000 100.200 ;
        RECT 171.000 96.000 171.400 100.200 ;
        RECT 173.800 97.900 174.200 100.200 ;
        RECT 175.400 97.900 175.800 100.200 ;
        RECT 178.200 95.900 178.600 100.200 ;
        RECT 179.800 95.900 180.200 100.200 ;
        RECT 181.900 97.900 182.300 100.200 ;
        RECT 183.000 97.900 183.400 100.200 ;
        RECT 184.600 97.900 185.000 100.200 ;
        RECT 185.400 95.900 185.800 100.200 ;
        RECT 187.000 96.500 187.400 100.200 ;
        RECT 188.600 97.900 189.000 100.200 ;
        RECT 190.200 97.900 190.600 100.200 ;
        RECT 193.400 96.500 193.800 100.200 ;
        RECT 196.100 97.900 196.500 100.200 ;
        RECT 198.200 95.900 198.600 100.200 ;
        RECT 199.800 96.500 200.200 100.200 ;
        RECT 202.500 97.900 202.900 100.200 ;
        RECT 204.600 95.900 205.000 100.200 ;
        RECT 206.200 96.000 206.600 100.200 ;
        RECT 209.000 97.900 209.400 100.200 ;
        RECT 210.600 97.900 211.000 100.200 ;
        RECT 213.400 95.900 213.800 100.200 ;
        RECT 215.800 96.000 216.200 100.200 ;
        RECT 218.600 97.900 219.000 100.200 ;
        RECT 220.200 97.900 220.600 100.200 ;
        RECT 223.000 95.900 223.400 100.200 ;
        RECT 225.400 96.500 225.800 100.200 ;
        RECT 227.800 96.500 228.200 100.200 ;
        RECT 1.400 80.800 1.800 85.000 ;
        RECT 4.200 80.800 4.600 83.100 ;
        RECT 5.800 80.800 6.200 83.100 ;
        RECT 8.600 80.800 9.000 85.100 ;
        RECT 10.500 80.800 10.900 83.100 ;
        RECT 12.600 80.800 13.000 85.100 ;
        RECT 13.700 80.800 14.100 83.100 ;
        RECT 15.800 80.800 16.200 85.100 ;
        RECT 16.600 80.800 17.000 85.100 ;
        RECT 18.700 80.800 19.100 83.100 ;
        RECT 20.100 80.800 20.500 83.100 ;
        RECT 22.200 80.800 22.600 85.100 ;
        RECT 23.000 80.800 23.400 85.100 ;
        RECT 25.100 80.800 25.500 83.100 ;
        RECT 26.200 80.800 26.600 85.100 ;
        RECT 28.300 80.800 28.700 83.100 ;
        RECT 30.200 80.800 30.600 85.000 ;
        RECT 33.000 80.800 33.400 83.100 ;
        RECT 34.600 80.800 35.000 83.100 ;
        RECT 37.400 80.800 37.800 85.100 ;
        RECT 40.600 80.800 41.000 83.100 ;
        RECT 42.200 80.800 42.600 83.100 ;
        RECT 43.800 80.800 44.200 85.000 ;
        RECT 46.600 80.800 47.000 83.100 ;
        RECT 48.200 80.800 48.600 83.100 ;
        RECT 51.000 80.800 51.400 85.100 ;
        RECT 52.600 80.800 53.000 85.100 ;
        RECT 54.700 80.800 55.100 83.100 ;
        RECT 55.800 80.800 56.200 83.100 ;
        RECT 57.400 80.800 57.800 83.100 ;
        RECT 58.200 80.800 58.600 83.100 ;
        RECT 59.800 80.800 60.200 85.100 ;
        RECT 63.000 80.800 63.400 85.100 ;
        RECT 64.600 80.800 65.000 83.100 ;
        RECT 65.400 80.800 65.800 85.100 ;
        RECT 67.500 80.800 67.900 83.100 ;
        RECT 68.600 80.800 69.000 85.100 ;
        RECT 70.200 80.800 70.600 85.100 ;
        RECT 71.800 80.800 72.200 85.100 ;
        RECT 73.400 80.800 73.800 85.100 ;
        RECT 75.000 80.800 75.400 85.100 ;
        RECT 75.800 80.800 76.200 83.100 ;
        RECT 77.400 80.800 77.800 82.900 ;
        RECT 79.800 80.800 80.200 85.100 ;
        RECT 82.600 80.800 83.000 83.100 ;
        RECT 84.200 80.800 84.600 83.100 ;
        RECT 87.000 80.800 87.400 85.000 ;
        RECT 90.200 80.800 90.600 85.100 ;
        RECT 92.300 80.800 92.700 83.100 ;
        RECT 93.400 80.800 93.800 83.100 ;
        RECT 95.000 80.800 95.400 83.100 ;
        RECT 95.800 80.800 96.200 85.100 ;
        RECT 97.900 80.800 98.300 83.100 ;
        RECT 99.800 80.800 100.200 85.000 ;
        RECT 102.600 80.800 103.000 83.100 ;
        RECT 104.200 80.800 104.600 83.100 ;
        RECT 107.000 80.800 107.400 85.100 ;
        RECT 108.600 80.800 109.000 85.100 ;
        RECT 110.700 80.800 111.100 83.100 ;
        RECT 112.600 80.800 113.000 84.500 ;
        RECT 115.000 80.800 115.400 85.100 ;
        RECT 117.100 80.800 117.500 83.100 ;
        RECT 118.200 80.800 118.600 85.100 ;
        RECT 120.300 80.800 120.700 83.100 ;
        RECT 122.200 80.800 122.600 85.000 ;
        RECT 125.000 80.800 125.400 83.100 ;
        RECT 126.600 80.800 127.000 83.100 ;
        RECT 129.400 80.800 129.800 85.100 ;
        RECT 131.800 80.800 132.200 85.100 ;
        RECT 134.600 80.800 135.000 83.100 ;
        RECT 136.200 80.800 136.600 83.100 ;
        RECT 139.000 80.800 139.400 85.000 ;
        RECT 142.200 80.800 142.600 83.100 ;
        RECT 143.800 80.800 144.200 83.100 ;
        RECT 144.900 80.800 145.300 83.100 ;
        RECT 147.000 80.800 147.400 85.100 ;
        RECT 147.800 80.800 148.200 83.100 ;
        RECT 149.400 80.800 149.800 83.100 ;
        RECT 150.200 80.800 150.600 83.100 ;
        RECT 151.800 80.800 152.200 83.100 ;
        RECT 153.400 80.800 153.800 84.500 ;
        RECT 156.600 80.800 157.000 84.500 ;
        RECT 159.800 80.800 160.200 84.500 ;
        RECT 163.000 80.800 163.400 84.500 ;
        RECT 165.700 80.800 166.100 83.100 ;
        RECT 167.800 80.800 168.200 85.100 ;
        RECT 168.900 80.800 169.300 83.100 ;
        RECT 171.000 80.800 171.400 85.100 ;
        RECT 172.600 80.800 173.000 84.500 ;
        RECT 174.500 80.800 174.900 83.100 ;
        RECT 176.600 80.800 177.000 85.100 ;
        RECT 179.000 80.800 179.400 84.500 ;
        RECT 180.600 80.800 181.000 85.100 ;
        RECT 182.700 80.800 183.100 83.100 ;
        RECT 183.800 80.800 184.200 83.100 ;
        RECT 185.400 80.800 185.800 83.100 ;
        RECT 186.800 80.800 187.200 85.100 ;
        RECT 189.400 80.800 189.800 84.900 ;
        RECT 192.600 80.800 193.000 85.100 ;
        RECT 194.700 80.800 195.100 83.100 ;
        RECT 195.800 80.800 196.200 83.100 ;
        RECT 197.400 80.800 197.800 83.100 ;
        RECT 199.000 80.800 199.400 85.100 ;
        RECT 201.800 80.800 202.200 83.100 ;
        RECT 203.400 80.800 203.800 83.100 ;
        RECT 206.200 80.800 206.600 85.000 ;
        RECT 208.600 80.800 209.000 84.900 ;
        RECT 211.200 80.800 211.600 85.100 ;
        RECT 213.400 80.800 213.800 85.100 ;
        RECT 216.200 80.800 216.600 83.100 ;
        RECT 217.800 80.800 218.200 83.100 ;
        RECT 220.600 80.800 221.000 85.000 ;
        RECT 222.200 80.800 222.600 83.100 ;
        RECT 223.800 80.800 224.200 83.100 ;
        RECT 224.900 80.800 225.300 83.100 ;
        RECT 227.000 80.800 227.400 85.100 ;
        RECT 227.800 80.800 228.200 83.100 ;
        RECT 229.400 80.800 229.800 83.100 ;
        RECT 0.200 80.200 231.000 80.800 ;
        RECT 1.400 76.000 1.800 80.200 ;
        RECT 4.200 77.900 4.600 80.200 ;
        RECT 5.800 77.900 6.200 80.200 ;
        RECT 8.600 75.900 9.000 80.200 ;
        RECT 10.200 75.900 10.600 80.200 ;
        RECT 12.300 77.900 12.700 80.200 ;
        RECT 13.400 77.900 13.800 80.200 ;
        RECT 15.000 77.900 15.400 80.200 ;
        RECT 15.800 75.900 16.200 80.200 ;
        RECT 17.900 77.900 18.300 80.200 ;
        RECT 19.000 77.900 19.400 80.200 ;
        RECT 20.600 77.900 21.000 80.200 ;
        RECT 22.200 76.000 22.600 80.200 ;
        RECT 25.000 77.900 25.400 80.200 ;
        RECT 26.600 77.900 27.000 80.200 ;
        RECT 29.400 75.900 29.800 80.200 ;
        RECT 31.000 75.900 31.400 80.200 ;
        RECT 34.200 75.900 34.600 80.200 ;
        RECT 35.800 77.900 36.200 80.200 ;
        RECT 36.600 77.900 37.000 80.200 ;
        RECT 39.800 75.900 40.200 80.200 ;
        RECT 43.000 75.900 43.400 80.200 ;
        RECT 43.800 75.900 44.200 80.200 ;
        RECT 45.900 77.900 46.300 80.200 ;
        RECT 47.000 75.900 47.400 80.200 ;
        RECT 49.100 77.900 49.500 80.200 ;
        RECT 51.000 76.500 51.400 80.200 ;
        RECT 52.600 75.900 53.000 80.200 ;
        RECT 53.700 77.900 54.100 80.200 ;
        RECT 55.800 75.900 56.200 80.200 ;
        RECT 56.600 77.900 57.000 80.200 ;
        RECT 58.200 77.900 58.600 80.200 ;
        RECT 59.000 75.900 59.400 80.200 ;
        RECT 61.100 77.900 61.500 80.200 ;
        RECT 62.500 77.900 62.900 80.200 ;
        RECT 64.600 75.900 65.000 80.200 ;
        RECT 65.400 75.900 65.800 80.200 ;
        RECT 67.500 77.900 67.900 80.200 ;
        RECT 68.600 77.900 69.000 80.200 ;
        RECT 70.200 77.900 70.600 80.200 ;
        RECT 71.800 75.900 72.200 80.200 ;
        RECT 74.600 77.900 75.000 80.200 ;
        RECT 76.200 77.900 76.600 80.200 ;
        RECT 79.000 76.000 79.400 80.200 ;
        RECT 80.600 75.900 81.000 80.200 ;
        RECT 83.000 75.900 83.400 80.200 ;
        RECT 85.100 77.900 85.500 80.200 ;
        RECT 86.200 77.900 86.600 80.200 ;
        RECT 87.800 77.900 88.200 80.200 ;
        RECT 91.000 75.900 91.400 80.200 ;
        RECT 93.800 77.900 94.200 80.200 ;
        RECT 95.400 77.900 95.800 80.200 ;
        RECT 98.200 76.000 98.600 80.200 ;
        RECT 100.600 76.100 101.000 80.200 ;
        RECT 103.200 75.900 103.600 80.200 ;
        RECT 104.600 77.900 105.000 80.200 ;
        RECT 106.200 78.100 106.600 80.200 ;
        RECT 107.800 77.900 108.200 80.200 ;
        RECT 109.400 77.900 109.800 80.200 ;
        RECT 110.200 75.900 110.600 80.200 ;
        RECT 112.300 77.900 112.700 80.200 ;
        RECT 113.400 77.900 113.800 80.200 ;
        RECT 115.000 78.100 115.400 80.200 ;
        RECT 116.600 75.900 117.000 80.200 ;
        RECT 118.200 76.500 118.600 80.200 ;
        RECT 119.800 77.900 120.200 80.200 ;
        RECT 121.400 77.900 121.800 80.200 ;
        RECT 122.200 75.900 122.600 80.200 ;
        RECT 123.800 76.500 124.200 80.200 ;
        RECT 126.200 76.000 126.600 80.200 ;
        RECT 129.000 77.900 129.400 80.200 ;
        RECT 130.600 77.900 131.000 80.200 ;
        RECT 133.400 75.900 133.800 80.200 ;
        RECT 135.000 75.900 135.400 80.200 ;
        RECT 137.100 77.900 137.500 80.200 ;
        RECT 138.200 77.900 138.600 80.200 ;
        RECT 139.800 77.900 140.200 80.200 ;
        RECT 142.200 75.900 142.600 80.200 ;
        RECT 144.300 77.900 144.700 80.200 ;
        RECT 145.400 77.900 145.800 80.200 ;
        RECT 147.000 77.900 147.400 80.200 ;
        RECT 148.600 76.000 149.000 80.200 ;
        RECT 151.400 77.900 151.800 80.200 ;
        RECT 153.000 77.900 153.400 80.200 ;
        RECT 155.800 75.900 156.200 80.200 ;
        RECT 157.400 75.900 157.800 80.200 ;
        RECT 159.000 75.900 159.400 80.200 ;
        RECT 160.600 75.900 161.000 80.200 ;
        RECT 162.200 76.000 162.600 80.200 ;
        RECT 165.000 77.900 165.400 80.200 ;
        RECT 166.600 77.900 167.000 80.200 ;
        RECT 169.400 75.900 169.800 80.200 ;
        RECT 171.800 76.500 172.200 80.200 ;
        RECT 173.700 77.900 174.100 80.200 ;
        RECT 175.800 75.900 176.200 80.200 ;
        RECT 177.400 76.500 177.800 80.200 ;
        RECT 179.000 75.900 179.400 80.200 ;
        RECT 180.600 78.100 181.000 80.200 ;
        RECT 182.200 77.900 182.600 80.200 ;
        RECT 183.000 77.900 183.400 80.200 ;
        RECT 184.600 77.900 185.000 80.200 ;
        RECT 186.200 76.100 186.600 80.200 ;
        RECT 188.800 75.900 189.200 80.200 ;
        RECT 192.100 77.900 192.500 80.200 ;
        RECT 194.200 75.900 194.600 80.200 ;
        RECT 195.800 77.900 196.200 80.200 ;
        RECT 197.200 75.900 197.600 80.200 ;
        RECT 199.800 76.100 200.200 80.200 ;
        RECT 202.000 75.900 202.400 80.200 ;
        RECT 204.600 76.100 205.000 80.200 ;
        RECT 207.000 75.900 207.400 80.200 ;
        RECT 209.800 77.900 210.200 80.200 ;
        RECT 211.400 77.900 211.800 80.200 ;
        RECT 214.200 76.000 214.600 80.200 ;
        RECT 215.800 77.900 216.200 80.200 ;
        RECT 217.400 77.900 217.800 80.200 ;
        RECT 218.500 77.900 218.900 80.200 ;
        RECT 220.600 75.900 221.000 80.200 ;
        RECT 221.400 75.900 221.800 80.200 ;
        RECT 223.000 75.900 223.400 80.200 ;
        RECT 224.600 75.900 225.000 80.200 ;
        RECT 226.200 75.900 226.600 80.200 ;
        RECT 227.800 75.900 228.200 80.200 ;
        RECT 229.400 76.500 229.800 80.200 ;
        RECT 0.600 60.800 1.000 65.100 ;
        RECT 2.200 60.800 2.600 65.100 ;
        RECT 3.800 60.800 4.200 65.100 ;
        RECT 5.400 60.800 5.800 65.000 ;
        RECT 8.200 60.800 8.600 63.100 ;
        RECT 9.800 60.800 10.200 63.100 ;
        RECT 12.600 60.800 13.000 65.100 ;
        RECT 14.500 60.800 14.900 63.100 ;
        RECT 16.600 60.800 17.000 65.100 ;
        RECT 17.400 60.800 17.800 63.100 ;
        RECT 19.000 60.800 19.400 65.100 ;
        RECT 21.100 60.800 21.500 63.100 ;
        RECT 23.000 60.800 23.400 65.000 ;
        RECT 25.800 60.800 26.200 63.100 ;
        RECT 27.400 60.800 27.800 63.100 ;
        RECT 30.200 60.800 30.600 65.100 ;
        RECT 31.800 60.800 32.200 65.100 ;
        RECT 33.900 60.800 34.300 63.100 ;
        RECT 35.000 60.800 35.400 65.100 ;
        RECT 36.600 60.800 37.000 64.500 ;
        RECT 40.100 60.800 40.500 63.100 ;
        RECT 42.200 60.800 42.600 65.100 ;
        RECT 43.800 60.800 44.200 64.500 ;
        RECT 45.400 60.800 45.800 65.100 ;
        RECT 46.200 60.800 46.600 63.100 ;
        RECT 47.800 60.800 48.200 63.100 ;
        RECT 48.600 60.800 49.000 63.100 ;
        RECT 50.200 60.800 50.600 63.100 ;
        RECT 51.800 60.800 52.200 65.000 ;
        RECT 54.600 60.800 55.000 63.100 ;
        RECT 56.200 60.800 56.600 63.100 ;
        RECT 59.000 60.800 59.400 65.100 ;
        RECT 60.600 60.800 61.000 63.100 ;
        RECT 62.200 60.800 62.600 63.100 ;
        RECT 63.000 60.800 63.400 63.100 ;
        RECT 64.600 60.800 65.000 63.100 ;
        RECT 65.400 60.800 65.800 63.100 ;
        RECT 67.000 60.800 67.400 63.100 ;
        RECT 68.600 60.800 69.000 64.900 ;
        RECT 71.200 60.800 71.600 65.100 ;
        RECT 72.600 60.800 73.000 65.100 ;
        RECT 74.700 60.800 75.100 63.100 ;
        RECT 75.800 60.800 76.200 63.100 ;
        RECT 77.400 60.800 77.800 63.100 ;
        RECT 79.000 60.800 79.400 65.000 ;
        RECT 81.800 60.800 82.200 63.100 ;
        RECT 83.400 60.800 83.800 63.100 ;
        RECT 86.200 60.800 86.600 65.100 ;
        RECT 90.000 60.800 90.400 65.100 ;
        RECT 92.600 60.800 93.000 64.900 ;
        RECT 94.200 60.800 94.600 63.100 ;
        RECT 95.800 60.800 96.200 63.100 ;
        RECT 96.900 60.800 97.300 63.100 ;
        RECT 99.000 60.800 99.400 65.100 ;
        RECT 100.600 60.800 101.000 64.500 ;
        RECT 103.300 60.800 103.700 63.100 ;
        RECT 105.400 60.800 105.800 65.100 ;
        RECT 106.200 60.800 106.600 65.100 ;
        RECT 108.300 60.800 108.700 63.100 ;
        RECT 109.400 60.800 109.800 63.100 ;
        RECT 111.000 60.800 111.400 63.100 ;
        RECT 111.800 60.800 112.200 63.100 ;
        RECT 113.400 60.800 113.800 63.100 ;
        RECT 114.200 60.800 114.600 63.100 ;
        RECT 115.800 60.800 116.200 63.100 ;
        RECT 116.900 60.800 117.300 63.100 ;
        RECT 119.000 60.800 119.400 65.100 ;
        RECT 119.800 60.800 120.200 65.100 ;
        RECT 121.900 60.800 122.300 63.100 ;
        RECT 123.800 60.800 124.200 64.500 ;
        RECT 126.200 60.800 126.600 65.100 ;
        RECT 128.300 60.800 128.700 63.100 ;
        RECT 130.200 60.800 130.600 65.100 ;
        RECT 133.000 60.800 133.400 63.100 ;
        RECT 134.600 60.800 135.000 63.100 ;
        RECT 137.400 60.800 137.800 65.000 ;
        RECT 141.400 60.800 141.800 64.500 ;
        RECT 143.800 60.800 144.200 63.100 ;
        RECT 145.400 60.800 145.800 62.900 ;
        RECT 147.000 60.800 147.400 65.100 ;
        RECT 149.100 60.800 149.500 63.100 ;
        RECT 151.000 60.800 151.400 64.900 ;
        RECT 153.600 60.800 154.000 65.100 ;
        RECT 155.800 60.800 156.200 64.500 ;
        RECT 159.000 60.800 159.400 64.500 ;
        RECT 162.200 60.800 162.600 64.500 ;
        RECT 164.900 60.800 165.300 63.100 ;
        RECT 167.000 60.800 167.400 65.100 ;
        RECT 168.600 60.800 169.000 64.500 ;
        RECT 171.300 60.800 171.700 63.100 ;
        RECT 173.400 60.800 173.800 65.100 ;
        RECT 175.000 60.800 175.400 65.000 ;
        RECT 177.800 60.800 178.200 63.100 ;
        RECT 179.400 60.800 179.800 63.100 ;
        RECT 182.200 60.800 182.600 65.100 ;
        RECT 183.800 60.800 184.200 63.100 ;
        RECT 185.400 60.800 185.800 63.100 ;
        RECT 186.200 60.800 186.600 63.100 ;
        RECT 187.800 60.800 188.200 63.100 ;
        RECT 189.400 60.800 189.800 64.500 ;
        RECT 191.000 60.800 191.400 65.100 ;
        RECT 194.200 60.800 194.600 65.100 ;
        RECT 197.000 60.800 197.400 63.100 ;
        RECT 198.600 60.800 199.000 63.100 ;
        RECT 201.400 60.800 201.800 65.000 ;
        RECT 203.000 60.800 203.400 65.100 ;
        RECT 205.100 60.800 205.500 63.100 ;
        RECT 206.200 60.800 206.600 63.100 ;
        RECT 207.800 60.800 208.200 63.100 ;
        RECT 208.900 60.800 209.300 63.100 ;
        RECT 211.000 60.800 211.400 65.100 ;
        RECT 212.600 60.800 213.000 65.100 ;
        RECT 215.400 60.800 215.800 63.100 ;
        RECT 217.000 60.800 217.400 63.100 ;
        RECT 219.800 60.800 220.200 65.000 ;
        RECT 222.200 60.800 222.600 65.000 ;
        RECT 225.000 60.800 225.400 63.100 ;
        RECT 226.600 60.800 227.000 63.100 ;
        RECT 229.400 60.800 229.800 65.100 ;
        RECT 0.200 60.200 231.000 60.800 ;
        RECT 1.400 56.500 1.800 60.200 ;
        RECT 3.000 55.900 3.400 60.200 ;
        RECT 4.600 56.000 5.000 60.200 ;
        RECT 7.400 57.900 7.800 60.200 ;
        RECT 9.000 57.900 9.400 60.200 ;
        RECT 11.800 55.900 12.200 60.200 ;
        RECT 13.400 57.900 13.800 60.200 ;
        RECT 15.000 57.900 15.400 60.200 ;
        RECT 15.800 55.900 16.200 60.200 ;
        RECT 17.900 57.900 18.300 60.200 ;
        RECT 19.000 57.900 19.400 60.200 ;
        RECT 20.600 57.900 21.000 60.200 ;
        RECT 21.400 55.900 21.800 60.200 ;
        RECT 23.000 55.900 23.400 60.200 ;
        RECT 24.600 55.900 25.000 60.200 ;
        RECT 26.200 55.900 26.600 60.200 ;
        RECT 27.800 55.900 28.200 60.200 ;
        RECT 28.600 57.900 29.000 60.200 ;
        RECT 30.200 57.900 30.600 60.200 ;
        RECT 31.000 55.900 31.400 60.200 ;
        RECT 33.100 57.900 33.500 60.200 ;
        RECT 36.600 56.000 37.000 60.200 ;
        RECT 39.400 57.900 39.800 60.200 ;
        RECT 41.000 57.900 41.400 60.200 ;
        RECT 43.800 55.900 44.200 60.200 ;
        RECT 45.400 55.900 45.800 60.200 ;
        RECT 47.500 57.900 47.900 60.200 ;
        RECT 48.600 57.900 49.000 60.200 ;
        RECT 50.200 57.900 50.600 60.200 ;
        RECT 51.000 57.900 51.400 60.200 ;
        RECT 52.600 55.900 53.000 60.200 ;
        RECT 54.700 57.900 55.100 60.200 ;
        RECT 55.800 55.900 56.200 60.200 ;
        RECT 57.900 57.900 58.300 60.200 ;
        RECT 59.000 55.900 59.400 60.200 ;
        RECT 61.100 57.900 61.500 60.200 ;
        RECT 63.000 56.000 63.400 60.200 ;
        RECT 65.800 57.900 66.200 60.200 ;
        RECT 67.400 57.900 67.800 60.200 ;
        RECT 70.200 55.900 70.600 60.200 ;
        RECT 72.600 56.500 73.000 60.200 ;
        RECT 74.200 55.900 74.600 60.200 ;
        RECT 75.000 57.900 75.400 60.200 ;
        RECT 76.600 57.900 77.000 60.200 ;
        RECT 78.200 56.100 78.600 60.200 ;
        RECT 80.800 55.900 81.200 60.200 ;
        RECT 82.800 55.900 83.200 60.200 ;
        RECT 85.400 56.100 85.800 60.200 ;
        RECT 89.400 56.100 89.800 60.200 ;
        RECT 92.000 55.900 92.400 60.200 ;
        RECT 94.200 56.000 94.600 60.200 ;
        RECT 97.000 57.900 97.400 60.200 ;
        RECT 98.600 57.900 99.000 60.200 ;
        RECT 101.400 55.900 101.800 60.200 ;
        RECT 103.000 57.900 103.400 60.200 ;
        RECT 104.600 57.900 105.000 60.200 ;
        RECT 105.400 57.900 105.800 60.200 ;
        RECT 107.000 57.900 107.400 60.200 ;
        RECT 107.800 57.900 108.200 60.200 ;
        RECT 109.700 57.900 110.100 60.200 ;
        RECT 111.800 55.900 112.200 60.200 ;
        RECT 113.400 56.500 113.800 60.200 ;
        RECT 115.000 55.900 115.400 60.200 ;
        RECT 116.600 56.100 117.000 60.200 ;
        RECT 119.200 55.900 119.600 60.200 ;
        RECT 121.400 58.100 121.800 60.200 ;
        RECT 123.000 57.900 123.400 60.200 ;
        RECT 123.800 57.900 124.200 60.200 ;
        RECT 125.400 57.900 125.800 60.200 ;
        RECT 127.000 56.500 127.400 60.200 ;
        RECT 128.600 55.900 129.000 60.200 ;
        RECT 129.400 57.900 129.800 60.200 ;
        RECT 131.000 58.100 131.400 60.200 ;
        RECT 132.600 57.900 133.000 60.200 ;
        RECT 134.200 57.900 134.600 60.200 ;
        RECT 135.800 56.100 136.200 60.200 ;
        RECT 138.400 55.900 138.800 60.200 ;
        RECT 142.200 57.900 142.600 60.200 ;
        RECT 144.100 55.900 144.500 60.200 ;
        RECT 146.500 57.900 146.900 60.200 ;
        RECT 148.600 55.900 149.000 60.200 ;
        RECT 149.400 57.900 149.800 60.200 ;
        RECT 151.000 57.900 151.400 60.200 ;
        RECT 152.600 56.000 153.000 60.200 ;
        RECT 155.400 57.900 155.800 60.200 ;
        RECT 157.000 57.900 157.400 60.200 ;
        RECT 159.800 55.900 160.200 60.200 ;
        RECT 161.400 57.900 161.800 60.200 ;
        RECT 163.000 57.900 163.400 60.200 ;
        RECT 164.100 57.900 164.500 60.200 ;
        RECT 166.200 55.900 166.600 60.200 ;
        RECT 167.800 56.100 168.200 60.200 ;
        RECT 170.400 55.900 170.800 60.200 ;
        RECT 172.600 56.000 173.000 60.200 ;
        RECT 175.400 57.900 175.800 60.200 ;
        RECT 177.000 57.900 177.400 60.200 ;
        RECT 179.800 55.900 180.200 60.200 ;
        RECT 181.400 55.900 181.800 60.200 ;
        RECT 183.000 56.500 183.400 60.200 ;
        RECT 185.400 56.100 185.800 60.200 ;
        RECT 188.000 55.900 188.400 60.200 ;
        RECT 189.400 57.900 189.800 60.200 ;
        RECT 191.000 57.900 191.400 60.200 ;
        RECT 193.700 57.900 194.100 60.200 ;
        RECT 195.800 55.900 196.200 60.200 ;
        RECT 197.400 56.500 197.800 60.200 ;
        RECT 199.000 55.900 199.400 60.200 ;
        RECT 200.600 57.900 201.000 60.200 ;
        RECT 202.200 56.100 202.600 60.200 ;
        RECT 204.800 55.900 205.200 60.200 ;
        RECT 207.000 56.100 207.400 60.200 ;
        RECT 209.600 55.900 210.000 60.200 ;
        RECT 211.000 55.900 211.400 60.200 ;
        RECT 212.600 56.500 213.000 60.200 ;
        RECT 214.200 55.900 214.600 60.200 ;
        RECT 216.300 57.900 216.700 60.200 ;
        RECT 218.200 55.900 218.600 60.200 ;
        RECT 221.000 57.900 221.400 60.200 ;
        RECT 222.600 57.900 223.000 60.200 ;
        RECT 225.400 56.000 225.800 60.200 ;
        RECT 227.800 56.500 228.200 60.200 ;
        RECT 229.400 55.900 229.800 60.200 ;
        RECT 1.400 40.800 1.800 45.000 ;
        RECT 4.200 40.800 4.600 43.100 ;
        RECT 5.800 40.800 6.200 43.100 ;
        RECT 8.600 40.800 9.000 45.100 ;
        RECT 10.200 40.800 10.600 43.100 ;
        RECT 11.800 40.800 12.200 43.100 ;
        RECT 12.900 40.800 13.300 43.100 ;
        RECT 15.000 40.800 15.400 45.100 ;
        RECT 15.800 40.800 16.200 43.100 ;
        RECT 17.400 40.800 17.800 43.100 ;
        RECT 19.000 40.800 19.400 45.000 ;
        RECT 21.800 40.800 22.200 43.100 ;
        RECT 23.400 40.800 23.800 43.100 ;
        RECT 26.200 40.800 26.600 45.100 ;
        RECT 27.800 40.800 28.200 43.100 ;
        RECT 29.400 40.800 29.800 43.100 ;
        RECT 30.500 40.800 30.900 43.100 ;
        RECT 32.600 40.800 33.000 45.100 ;
        RECT 33.400 40.800 33.800 43.100 ;
        RECT 35.000 40.800 35.400 43.100 ;
        RECT 38.200 40.800 38.600 45.000 ;
        RECT 41.000 40.800 41.400 43.100 ;
        RECT 42.600 40.800 43.000 43.100 ;
        RECT 45.400 40.800 45.800 45.100 ;
        RECT 47.000 40.800 47.400 45.100 ;
        RECT 49.100 40.800 49.500 43.100 ;
        RECT 50.200 40.800 50.600 43.100 ;
        RECT 51.800 40.800 52.200 43.100 ;
        RECT 53.400 40.800 53.800 45.100 ;
        RECT 56.200 40.800 56.600 43.100 ;
        RECT 57.800 40.800 58.200 43.100 ;
        RECT 60.600 40.800 61.000 45.000 ;
        RECT 62.500 40.800 62.900 43.100 ;
        RECT 64.600 40.800 65.000 45.100 ;
        RECT 66.200 40.800 66.600 45.000 ;
        RECT 69.000 40.800 69.400 43.100 ;
        RECT 70.600 40.800 71.000 43.100 ;
        RECT 73.400 40.800 73.800 45.100 ;
        RECT 75.300 40.800 75.700 43.100 ;
        RECT 77.400 40.800 77.800 45.100 ;
        RECT 78.200 40.800 78.600 45.100 ;
        RECT 80.300 40.800 80.700 43.100 ;
        RECT 81.400 40.800 81.800 43.100 ;
        RECT 83.000 40.800 83.400 43.100 ;
        RECT 84.600 40.800 85.000 45.100 ;
        RECT 87.400 40.800 87.800 43.100 ;
        RECT 89.000 40.800 89.400 43.100 ;
        RECT 91.800 40.800 92.200 45.000 ;
        RECT 95.000 40.800 95.400 45.100 ;
        RECT 97.100 40.800 97.500 43.100 ;
        RECT 98.200 40.800 98.600 43.100 ;
        RECT 99.800 40.800 100.200 43.100 ;
        RECT 101.400 40.800 101.800 45.000 ;
        RECT 104.200 40.800 104.600 43.100 ;
        RECT 105.800 40.800 106.200 43.100 ;
        RECT 108.600 40.800 109.000 45.100 ;
        RECT 110.200 40.800 110.600 43.100 ;
        RECT 112.400 40.800 112.800 45.100 ;
        RECT 115.000 40.800 115.400 44.900 ;
        RECT 117.400 40.800 117.800 44.900 ;
        RECT 120.000 40.800 120.400 45.100 ;
        RECT 121.400 40.800 121.800 43.100 ;
        RECT 123.000 40.800 123.400 43.100 ;
        RECT 123.800 40.800 124.200 43.100 ;
        RECT 125.400 40.800 125.800 43.100 ;
        RECT 127.000 40.800 127.400 45.100 ;
        RECT 129.800 40.800 130.200 43.100 ;
        RECT 131.400 40.800 131.800 43.100 ;
        RECT 134.200 40.800 134.600 45.000 ;
        RECT 135.800 40.800 136.200 43.100 ;
        RECT 137.400 40.800 137.800 43.100 ;
        RECT 138.500 40.800 138.900 43.100 ;
        RECT 140.600 40.800 141.000 45.100 ;
        RECT 143.000 40.800 143.400 45.100 ;
        RECT 144.600 40.800 145.000 45.100 ;
        RECT 145.400 40.800 145.800 43.100 ;
        RECT 147.000 40.800 147.400 43.100 ;
        RECT 147.800 40.800 148.200 45.100 ;
        RECT 149.900 40.800 150.300 43.100 ;
        RECT 151.800 40.800 152.200 45.000 ;
        RECT 154.600 40.800 155.000 43.100 ;
        RECT 156.200 40.800 156.600 43.100 ;
        RECT 159.000 40.800 159.400 45.100 ;
        RECT 161.400 40.800 161.800 44.500 ;
        RECT 163.000 40.800 163.400 45.100 ;
        RECT 165.100 40.800 165.500 43.100 ;
        RECT 166.200 40.800 166.600 43.100 ;
        RECT 167.800 40.800 168.200 43.100 ;
        RECT 169.400 40.800 169.800 45.100 ;
        RECT 172.200 40.800 172.600 43.100 ;
        RECT 173.800 40.800 174.200 43.100 ;
        RECT 176.600 40.800 177.000 45.000 ;
        RECT 178.200 40.800 178.600 45.100 ;
        RECT 179.800 40.800 180.200 44.500 ;
        RECT 182.200 40.800 182.600 44.900 ;
        RECT 184.800 40.800 185.200 45.100 ;
        RECT 187.000 40.800 187.400 45.100 ;
        RECT 189.800 40.800 190.200 43.100 ;
        RECT 191.400 40.800 191.800 43.100 ;
        RECT 194.200 40.800 194.600 45.000 ;
        RECT 198.200 40.800 198.600 44.500 ;
        RECT 199.800 40.800 200.200 45.100 ;
        RECT 200.600 40.800 201.000 45.100 ;
        RECT 202.200 40.800 202.600 44.500 ;
        RECT 204.400 40.800 204.800 45.100 ;
        RECT 207.000 40.800 207.400 44.900 ;
        RECT 208.600 40.800 209.000 43.100 ;
        RECT 210.200 40.800 210.600 43.100 ;
        RECT 211.300 40.800 211.700 43.100 ;
        RECT 213.400 40.800 213.800 45.100 ;
        RECT 214.200 40.800 214.600 43.100 ;
        RECT 215.800 40.800 216.200 43.100 ;
        RECT 216.600 40.800 217.000 45.100 ;
        RECT 218.700 40.800 219.100 43.100 ;
        RECT 220.600 40.800 221.000 45.100 ;
        RECT 223.400 40.800 223.800 43.100 ;
        RECT 225.000 40.800 225.400 43.100 ;
        RECT 227.800 40.800 228.200 45.000 ;
        RECT 0.200 40.200 231.000 40.800 ;
        RECT 0.600 37.900 1.000 40.200 ;
        RECT 2.200 37.900 2.600 40.200 ;
        RECT 3.000 37.900 3.400 40.200 ;
        RECT 4.600 35.900 5.000 40.200 ;
        RECT 6.700 37.900 7.100 40.200 ;
        RECT 7.800 37.900 8.200 40.200 ;
        RECT 9.400 37.900 9.800 40.200 ;
        RECT 10.200 37.900 10.600 40.200 ;
        RECT 11.800 35.900 12.200 40.200 ;
        RECT 15.000 35.900 15.400 40.200 ;
        RECT 16.600 36.000 17.000 40.200 ;
        RECT 19.400 37.900 19.800 40.200 ;
        RECT 21.000 37.900 21.400 40.200 ;
        RECT 23.800 35.900 24.200 40.200 ;
        RECT 25.400 37.900 25.800 40.200 ;
        RECT 27.000 35.900 27.400 40.200 ;
        RECT 30.200 35.900 30.600 40.200 ;
        RECT 31.800 37.900 32.200 40.200 ;
        RECT 33.400 36.000 33.800 40.200 ;
        RECT 36.200 37.900 36.600 40.200 ;
        RECT 37.800 37.900 38.200 40.200 ;
        RECT 40.600 35.900 41.000 40.200 ;
        RECT 44.600 37.900 45.000 40.200 ;
        RECT 45.400 37.900 45.800 40.200 ;
        RECT 47.000 37.900 47.400 40.200 ;
        RECT 48.100 37.900 48.500 40.200 ;
        RECT 50.200 35.900 50.600 40.200 ;
        RECT 51.800 36.500 52.200 40.200 ;
        RECT 53.400 35.900 53.800 40.200 ;
        RECT 54.800 35.900 55.200 40.200 ;
        RECT 57.400 36.100 57.800 40.200 ;
        RECT 59.000 37.900 59.400 40.200 ;
        RECT 60.600 37.900 61.000 40.200 ;
        RECT 61.400 35.900 61.800 40.200 ;
        RECT 63.500 37.900 63.900 40.200 ;
        RECT 64.600 37.900 65.000 40.200 ;
        RECT 66.200 37.900 66.600 40.200 ;
        RECT 67.600 35.900 68.000 40.200 ;
        RECT 70.200 36.100 70.600 40.200 ;
        RECT 71.800 35.900 72.200 40.200 ;
        RECT 73.900 37.900 74.300 40.200 ;
        RECT 75.000 37.900 75.400 40.200 ;
        RECT 76.600 37.900 77.000 40.200 ;
        RECT 77.400 35.900 77.800 40.200 ;
        RECT 79.500 37.900 79.900 40.200 ;
        RECT 80.600 37.900 81.000 40.200 ;
        RECT 82.200 37.900 82.600 40.200 ;
        RECT 83.600 35.900 84.000 40.200 ;
        RECT 86.200 36.100 86.600 40.200 ;
        RECT 90.200 35.900 90.600 40.200 ;
        RECT 93.000 37.900 93.400 40.200 ;
        RECT 94.600 37.900 95.000 40.200 ;
        RECT 97.400 36.000 97.800 40.200 ;
        RECT 99.000 37.900 99.400 40.200 ;
        RECT 100.600 37.900 101.000 40.200 ;
        RECT 101.700 37.900 102.100 40.200 ;
        RECT 103.800 35.900 104.200 40.200 ;
        RECT 104.600 37.900 105.000 40.200 ;
        RECT 106.200 37.900 106.600 40.200 ;
        RECT 107.800 36.100 108.200 40.200 ;
        RECT 110.400 35.900 110.800 40.200 ;
        RECT 111.800 37.900 112.200 40.200 ;
        RECT 113.400 37.900 113.800 40.200 ;
        RECT 114.500 37.900 114.900 40.200 ;
        RECT 116.600 35.900 117.000 40.200 ;
        RECT 117.400 35.900 117.800 40.200 ;
        RECT 119.500 37.900 119.900 40.200 ;
        RECT 121.200 35.900 121.600 40.200 ;
        RECT 123.800 36.100 124.200 40.200 ;
        RECT 126.200 36.100 126.600 40.200 ;
        RECT 128.800 35.900 129.200 40.200 ;
        RECT 131.000 36.100 131.400 40.200 ;
        RECT 133.600 35.900 134.000 40.200 ;
        RECT 135.000 37.900 135.400 40.200 ;
        RECT 136.600 37.900 137.000 40.200 ;
        RECT 137.700 37.900 138.100 40.200 ;
        RECT 139.800 35.900 140.200 40.200 ;
        RECT 143.000 35.900 143.400 40.200 ;
        RECT 145.800 37.900 146.200 40.200 ;
        RECT 147.400 37.900 147.800 40.200 ;
        RECT 150.200 36.000 150.600 40.200 ;
        RECT 151.800 35.900 152.200 40.200 ;
        RECT 155.000 35.900 155.400 40.200 ;
        RECT 156.400 35.900 156.800 40.200 ;
        RECT 159.000 36.100 159.400 40.200 ;
        RECT 160.600 37.900 161.000 40.200 ;
        RECT 162.200 37.900 162.600 40.200 ;
        RECT 163.000 37.900 163.400 40.200 ;
        RECT 164.600 37.900 165.000 40.200 ;
        RECT 165.400 35.900 165.800 40.200 ;
        RECT 167.500 37.900 167.900 40.200 ;
        RECT 169.400 37.900 169.800 40.200 ;
        RECT 170.200 35.900 170.600 40.200 ;
        RECT 171.800 36.500 172.200 40.200 ;
        RECT 173.400 37.900 173.800 40.200 ;
        RECT 175.000 37.900 175.400 40.200 ;
        RECT 176.100 37.900 176.500 40.200 ;
        RECT 178.200 35.900 178.600 40.200 ;
        RECT 179.800 36.100 180.200 40.200 ;
        RECT 182.400 35.900 182.800 40.200 ;
        RECT 184.600 37.900 185.000 40.200 ;
        RECT 186.200 35.900 186.600 40.200 ;
        RECT 189.000 37.900 189.400 40.200 ;
        RECT 190.600 37.900 191.000 40.200 ;
        RECT 193.400 36.000 193.800 40.200 ;
        RECT 196.600 35.900 197.000 40.200 ;
        RECT 198.700 37.900 199.100 40.200 ;
        RECT 199.800 35.900 200.200 40.200 ;
        RECT 201.900 37.900 202.300 40.200 ;
        RECT 203.000 37.900 203.400 40.200 ;
        RECT 204.600 37.900 205.000 40.200 ;
        RECT 206.200 35.900 206.600 40.200 ;
        RECT 209.000 37.900 209.400 40.200 ;
        RECT 210.600 37.900 211.000 40.200 ;
        RECT 213.400 36.000 213.800 40.200 ;
        RECT 215.000 35.900 215.400 40.200 ;
        RECT 217.100 37.900 217.500 40.200 ;
        RECT 218.200 37.900 218.600 40.200 ;
        RECT 219.800 37.900 220.200 40.200 ;
        RECT 221.400 35.900 221.800 40.200 ;
        RECT 224.200 37.900 224.600 40.200 ;
        RECT 225.800 37.900 226.200 40.200 ;
        RECT 228.600 36.000 229.000 40.200 ;
        RECT 0.900 20.800 1.300 23.100 ;
        RECT 3.000 20.800 3.400 25.100 ;
        RECT 4.600 20.800 5.000 25.100 ;
        RECT 7.400 20.800 7.800 23.100 ;
        RECT 9.000 20.800 9.400 23.100 ;
        RECT 11.800 20.800 12.200 25.000 ;
        RECT 14.200 20.800 14.600 25.100 ;
        RECT 17.000 20.800 17.400 23.100 ;
        RECT 18.600 20.800 19.000 23.100 ;
        RECT 21.400 20.800 21.800 25.000 ;
        RECT 23.000 20.800 23.400 23.100 ;
        RECT 24.600 20.800 25.000 23.100 ;
        RECT 26.200 20.800 26.600 23.100 ;
        RECT 27.300 20.800 27.700 23.100 ;
        RECT 29.400 20.800 29.800 25.100 ;
        RECT 30.200 20.800 30.600 25.100 ;
        RECT 31.800 20.800 32.200 25.100 ;
        RECT 33.400 20.800 33.800 25.100 ;
        RECT 35.000 20.800 35.400 25.100 ;
        RECT 36.600 20.800 37.000 25.100 ;
        RECT 39.800 20.800 40.200 25.100 ;
        RECT 42.600 20.800 43.000 23.100 ;
        RECT 44.200 20.800 44.600 23.100 ;
        RECT 47.000 20.800 47.400 25.000 ;
        RECT 48.600 20.800 49.000 25.100 ;
        RECT 50.700 20.800 51.100 23.100 ;
        RECT 51.800 20.800 52.200 23.100 ;
        RECT 53.400 20.800 53.800 23.100 ;
        RECT 54.200 20.800 54.600 23.100 ;
        RECT 55.800 20.800 56.200 23.100 ;
        RECT 56.900 20.800 57.300 23.100 ;
        RECT 59.000 20.800 59.400 25.100 ;
        RECT 60.600 20.800 61.000 25.000 ;
        RECT 63.400 20.800 63.800 23.100 ;
        RECT 65.000 20.800 65.400 23.100 ;
        RECT 67.800 20.800 68.200 25.100 ;
        RECT 70.200 20.800 70.600 25.100 ;
        RECT 73.000 20.800 73.400 23.100 ;
        RECT 74.600 20.800 75.000 23.100 ;
        RECT 77.400 20.800 77.800 25.000 ;
        RECT 79.000 20.800 79.400 23.100 ;
        RECT 80.600 20.800 81.000 23.100 ;
        RECT 81.700 20.800 82.100 23.100 ;
        RECT 83.800 20.800 84.200 25.100 ;
        RECT 87.000 20.800 87.400 25.100 ;
        RECT 89.800 20.800 90.200 23.100 ;
        RECT 91.400 20.800 91.800 23.100 ;
        RECT 94.200 20.800 94.600 25.000 ;
        RECT 95.800 20.800 96.200 23.100 ;
        RECT 97.400 20.800 97.800 23.100 ;
        RECT 98.200 20.800 98.600 23.100 ;
        RECT 99.800 20.800 100.200 23.100 ;
        RECT 100.600 20.800 101.000 23.100 ;
        RECT 102.200 20.800 102.600 23.100 ;
        RECT 103.000 20.800 103.400 25.100 ;
        RECT 105.100 20.800 105.500 23.100 ;
        RECT 107.000 20.800 107.400 25.000 ;
        RECT 109.800 20.800 110.200 23.100 ;
        RECT 111.400 20.800 111.800 23.100 ;
        RECT 114.200 20.800 114.600 25.100 ;
        RECT 116.600 20.800 117.000 25.100 ;
        RECT 119.400 20.800 119.800 23.100 ;
        RECT 121.000 20.800 121.400 23.100 ;
        RECT 123.800 20.800 124.200 25.000 ;
        RECT 125.400 20.800 125.800 23.100 ;
        RECT 127.000 20.800 127.400 23.100 ;
        RECT 127.800 20.800 128.200 25.100 ;
        RECT 129.400 20.800 129.800 25.100 ;
        RECT 131.000 20.800 131.400 25.100 ;
        RECT 132.600 20.800 133.000 25.100 ;
        RECT 134.200 20.800 134.600 25.100 ;
        RECT 135.000 20.800 135.400 25.100 ;
        RECT 136.600 20.800 137.000 25.100 ;
        RECT 138.200 20.800 138.600 25.100 ;
        RECT 139.800 20.800 140.200 25.100 ;
        RECT 141.400 20.800 141.800 25.100 ;
        RECT 143.800 20.800 144.200 23.100 ;
        RECT 145.400 20.800 145.800 23.100 ;
        RECT 146.500 20.800 146.900 23.100 ;
        RECT 148.600 20.800 149.000 25.100 ;
        RECT 150.200 20.800 150.600 25.100 ;
        RECT 153.000 20.800 153.400 23.100 ;
        RECT 154.600 20.800 155.000 23.100 ;
        RECT 157.400 20.800 157.800 25.000 ;
        RECT 159.000 20.800 159.400 25.100 ;
        RECT 161.100 20.800 161.500 23.100 ;
        RECT 162.200 20.800 162.600 25.100 ;
        RECT 164.300 20.800 164.700 23.100 ;
        RECT 165.400 20.800 165.800 23.100 ;
        RECT 167.000 20.800 167.400 23.100 ;
        RECT 168.600 20.800 169.000 25.100 ;
        RECT 171.400 20.800 171.800 23.100 ;
        RECT 173.000 20.800 173.400 23.100 ;
        RECT 175.800 20.800 176.200 25.000 ;
        RECT 178.200 20.800 178.600 25.100 ;
        RECT 181.000 20.800 181.400 23.100 ;
        RECT 182.600 20.800 183.000 23.100 ;
        RECT 185.400 20.800 185.800 25.000 ;
        RECT 189.400 20.800 189.800 25.000 ;
        RECT 192.200 20.800 192.600 23.100 ;
        RECT 193.800 20.800 194.200 23.100 ;
        RECT 196.600 20.800 197.000 25.100 ;
        RECT 198.200 20.800 198.600 23.100 ;
        RECT 199.800 20.800 200.200 23.100 ;
        RECT 201.400 20.800 201.800 24.500 ;
        RECT 203.000 20.800 203.400 25.100 ;
        RECT 203.800 20.800 204.200 25.100 ;
        RECT 205.900 20.800 206.300 23.100 ;
        RECT 207.000 20.800 207.400 23.100 ;
        RECT 208.600 20.800 209.000 23.100 ;
        RECT 210.200 20.800 210.600 25.100 ;
        RECT 213.000 20.800 213.400 23.100 ;
        RECT 214.600 20.800 215.000 23.100 ;
        RECT 217.400 20.800 217.800 25.000 ;
        RECT 219.000 20.800 219.400 23.100 ;
        RECT 220.600 20.800 221.000 23.100 ;
        RECT 222.200 20.800 222.600 25.100 ;
        RECT 225.000 20.800 225.400 23.100 ;
        RECT 226.600 20.800 227.000 23.100 ;
        RECT 229.400 20.800 229.800 25.000 ;
        RECT 0.200 20.200 231.000 20.800 ;
        RECT 1.400 16.000 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 15.900 9.000 20.200 ;
        RECT 10.200 15.900 10.600 20.200 ;
        RECT 12.300 17.900 12.700 20.200 ;
        RECT 14.200 16.000 14.600 20.200 ;
        RECT 17.000 17.900 17.400 20.200 ;
        RECT 18.600 17.900 19.000 20.200 ;
        RECT 21.400 15.900 21.800 20.200 ;
        RECT 23.000 17.900 23.400 20.200 ;
        RECT 25.400 16.000 25.800 20.200 ;
        RECT 28.200 17.900 28.600 20.200 ;
        RECT 29.800 17.900 30.200 20.200 ;
        RECT 32.600 15.900 33.000 20.200 ;
        RECT 34.500 17.900 34.900 20.200 ;
        RECT 36.600 15.900 37.000 20.200 ;
        RECT 39.600 15.900 40.000 20.200 ;
        RECT 42.200 16.100 42.600 20.200 ;
        RECT 44.600 16.500 45.000 20.200 ;
        RECT 46.200 15.900 46.600 20.200 ;
        RECT 47.800 16.000 48.200 20.200 ;
        RECT 50.600 17.900 51.000 20.200 ;
        RECT 52.200 17.900 52.600 20.200 ;
        RECT 55.000 15.900 55.400 20.200 ;
        RECT 56.600 15.900 57.000 20.200 ;
        RECT 58.700 17.900 59.100 20.200 ;
        RECT 59.800 17.900 60.200 20.200 ;
        RECT 61.400 17.900 61.800 20.200 ;
        RECT 62.200 17.900 62.600 20.200 ;
        RECT 63.800 15.900 64.200 20.200 ;
        RECT 65.900 17.900 66.300 20.200 ;
        RECT 67.000 17.900 67.400 20.200 ;
        RECT 68.600 17.900 69.000 20.200 ;
        RECT 70.200 16.000 70.600 20.200 ;
        RECT 73.000 17.900 73.400 20.200 ;
        RECT 74.600 17.900 75.000 20.200 ;
        RECT 77.400 15.900 77.800 20.200 ;
        RECT 79.000 15.900 79.400 20.200 ;
        RECT 80.600 15.900 81.000 20.200 ;
        RECT 82.200 15.900 82.600 20.200 ;
        RECT 84.300 17.900 84.700 20.200 ;
        RECT 85.400 17.900 85.800 20.200 ;
        RECT 87.000 17.900 87.400 20.200 ;
        RECT 90.200 16.000 90.600 20.200 ;
        RECT 93.000 17.900 93.400 20.200 ;
        RECT 94.600 17.900 95.000 20.200 ;
        RECT 97.400 15.900 97.800 20.200 ;
        RECT 99.000 17.900 99.400 20.200 ;
        RECT 101.400 16.000 101.800 20.200 ;
        RECT 104.200 17.900 104.600 20.200 ;
        RECT 105.800 17.900 106.200 20.200 ;
        RECT 108.600 15.900 109.000 20.200 ;
        RECT 110.200 15.900 110.600 20.200 ;
        RECT 112.300 17.900 112.700 20.200 ;
        RECT 113.400 17.900 113.800 20.200 ;
        RECT 115.000 17.900 115.400 20.200 ;
        RECT 116.600 16.100 117.000 20.200 ;
        RECT 119.200 15.900 119.600 20.200 ;
        RECT 120.600 15.900 121.000 20.200 ;
        RECT 122.700 17.900 123.100 20.200 ;
        RECT 123.800 17.900 124.200 20.200 ;
        RECT 125.400 17.900 125.800 20.200 ;
        RECT 127.000 16.500 127.400 20.200 ;
        RECT 128.600 15.900 129.000 20.200 ;
        RECT 129.400 17.900 129.800 20.200 ;
        RECT 131.000 17.900 131.400 20.200 ;
        RECT 132.400 15.900 132.800 20.200 ;
        RECT 135.000 16.100 135.400 20.200 ;
        RECT 136.600 17.900 137.000 20.200 ;
        RECT 138.200 17.900 138.600 20.200 ;
        RECT 140.900 17.900 141.300 20.200 ;
        RECT 143.000 15.900 143.400 20.200 ;
        RECT 144.400 15.900 144.800 20.200 ;
        RECT 147.000 16.100 147.400 20.200 ;
        RECT 149.400 16.000 149.800 20.200 ;
        RECT 152.200 17.900 152.600 20.200 ;
        RECT 153.800 17.900 154.200 20.200 ;
        RECT 156.600 15.900 157.000 20.200 ;
        RECT 159.000 16.000 159.400 20.200 ;
        RECT 161.800 17.900 162.200 20.200 ;
        RECT 163.400 17.900 163.800 20.200 ;
        RECT 166.200 15.900 166.600 20.200 ;
        RECT 167.800 17.900 168.200 20.200 ;
        RECT 169.400 17.900 169.800 20.200 ;
        RECT 170.500 17.900 170.900 20.200 ;
        RECT 172.600 15.900 173.000 20.200 ;
        RECT 174.200 16.000 174.600 20.200 ;
        RECT 177.000 17.900 177.400 20.200 ;
        RECT 178.600 17.900 179.000 20.200 ;
        RECT 181.400 15.900 181.800 20.200 ;
        RECT 183.000 15.900 183.400 20.200 ;
        RECT 184.600 15.900 185.000 20.200 ;
        RECT 185.400 15.900 185.800 20.200 ;
        RECT 187.800 15.900 188.200 20.200 ;
        RECT 189.400 15.900 189.800 20.200 ;
        RECT 192.600 15.900 193.000 20.200 ;
        RECT 195.400 17.900 195.800 20.200 ;
        RECT 197.000 17.900 197.400 20.200 ;
        RECT 199.800 16.000 200.200 20.200 ;
        RECT 202.200 16.100 202.600 20.200 ;
        RECT 204.800 15.900 205.200 20.200 ;
        RECT 206.200 17.900 206.600 20.200 ;
        RECT 207.800 17.900 208.200 20.200 ;
        RECT 208.900 17.900 209.300 20.200 ;
        RECT 211.000 15.900 211.400 20.200 ;
        RECT 211.800 15.900 212.200 20.200 ;
        RECT 213.900 17.900 214.300 20.200 ;
        RECT 215.000 17.900 215.400 20.200 ;
        RECT 216.600 17.900 217.000 20.200 ;
        RECT 217.400 15.900 217.800 20.200 ;
        RECT 219.000 15.900 219.400 20.200 ;
        RECT 220.600 15.900 221.000 20.200 ;
        RECT 222.200 15.900 222.600 20.200 ;
        RECT 223.800 15.900 224.200 20.200 ;
        RECT 224.600 17.900 225.000 20.200 ;
        RECT 226.200 17.900 226.600 20.200 ;
        RECT 227.300 17.900 227.700 20.200 ;
        RECT 229.400 15.900 229.800 20.200 ;
        RECT 0.900 0.800 1.300 3.100 ;
        RECT 3.000 0.800 3.400 5.100 ;
        RECT 3.800 0.800 4.200 3.100 ;
        RECT 5.400 0.800 5.800 3.100 ;
        RECT 6.200 0.800 6.600 5.100 ;
        RECT 7.800 0.800 8.200 4.500 ;
        RECT 9.400 0.800 9.800 5.100 ;
        RECT 11.000 0.800 11.400 5.100 ;
        RECT 12.600 0.800 13.000 5.100 ;
        RECT 13.400 0.800 13.800 3.100 ;
        RECT 15.000 0.800 15.400 3.100 ;
        RECT 15.800 0.800 16.200 5.100 ;
        RECT 17.400 0.800 17.800 5.100 ;
        RECT 19.000 0.800 19.400 5.100 ;
        RECT 20.600 0.800 21.000 4.500 ;
        RECT 22.200 0.800 22.600 5.100 ;
        RECT 23.000 0.800 23.400 5.100 ;
        RECT 24.600 0.800 25.000 5.100 ;
        RECT 26.200 0.800 26.600 5.100 ;
        RECT 27.800 0.800 28.200 5.100 ;
        RECT 29.400 0.800 29.800 5.100 ;
        RECT 31.000 0.800 31.400 5.000 ;
        RECT 33.800 0.800 34.200 3.100 ;
        RECT 35.400 0.800 35.800 3.100 ;
        RECT 38.200 0.800 38.600 5.100 ;
        RECT 41.400 0.800 41.800 3.100 ;
        RECT 43.000 0.800 43.400 3.100 ;
        RECT 43.800 0.800 44.200 3.100 ;
        RECT 45.400 0.800 45.800 3.100 ;
        RECT 46.500 0.800 46.900 3.100 ;
        RECT 48.600 0.800 49.000 5.100 ;
        RECT 50.200 0.800 50.600 5.100 ;
        RECT 53.000 0.800 53.400 3.100 ;
        RECT 54.600 0.800 55.000 3.100 ;
        RECT 57.400 0.800 57.800 5.000 ;
        RECT 59.800 0.800 60.200 5.000 ;
        RECT 62.600 0.800 63.000 3.100 ;
        RECT 64.200 0.800 64.600 3.100 ;
        RECT 67.000 0.800 67.400 5.100 ;
        RECT 69.400 0.800 69.800 5.000 ;
        RECT 72.200 0.800 72.600 3.100 ;
        RECT 73.800 0.800 74.200 3.100 ;
        RECT 76.600 0.800 77.000 5.100 ;
        RECT 79.800 0.800 80.200 4.500 ;
        RECT 82.200 0.800 82.600 4.500 ;
        RECT 86.200 0.800 86.600 5.100 ;
        RECT 87.000 0.800 87.400 5.100 ;
        RECT 91.000 0.800 91.400 5.100 ;
        RECT 93.100 0.800 93.500 3.100 ;
        RECT 94.200 0.800 94.600 3.100 ;
        RECT 95.800 0.800 96.200 3.100 ;
        RECT 97.400 0.800 97.800 5.000 ;
        RECT 100.200 0.800 100.600 3.100 ;
        RECT 101.800 0.800 102.200 3.100 ;
        RECT 104.600 0.800 105.000 5.100 ;
        RECT 106.200 0.800 106.600 5.100 ;
        RECT 107.800 0.800 108.200 5.100 ;
        RECT 109.400 0.800 109.800 5.100 ;
        RECT 111.000 0.800 111.400 5.000 ;
        RECT 113.800 0.800 114.200 3.100 ;
        RECT 115.400 0.800 115.800 3.100 ;
        RECT 118.200 0.800 118.600 5.100 ;
        RECT 120.600 0.800 121.000 5.000 ;
        RECT 123.400 0.800 123.800 3.100 ;
        RECT 125.000 0.800 125.400 3.100 ;
        RECT 127.800 0.800 128.200 5.100 ;
        RECT 129.700 0.800 130.100 3.100 ;
        RECT 131.800 0.800 132.200 5.100 ;
        RECT 133.400 0.800 133.800 5.100 ;
        RECT 136.200 0.800 136.600 3.100 ;
        RECT 137.800 0.800 138.200 3.100 ;
        RECT 140.600 0.800 141.000 5.000 ;
        RECT 144.600 0.800 145.000 5.100 ;
        RECT 147.400 0.800 147.800 3.100 ;
        RECT 149.000 0.800 149.400 3.100 ;
        RECT 151.800 0.800 152.200 5.000 ;
        RECT 153.400 0.800 153.800 3.100 ;
        RECT 155.000 0.800 155.400 3.100 ;
        RECT 156.100 0.800 156.500 3.100 ;
        RECT 158.200 0.800 158.600 5.100 ;
        RECT 159.000 0.800 159.400 5.100 ;
        RECT 161.100 0.800 161.500 3.100 ;
        RECT 162.200 0.800 162.600 3.100 ;
        RECT 163.800 0.800 164.200 3.100 ;
        RECT 165.400 0.800 165.800 5.100 ;
        RECT 168.200 0.800 168.600 3.100 ;
        RECT 169.800 0.800 170.200 3.100 ;
        RECT 172.600 0.800 173.000 5.000 ;
        RECT 174.200 0.800 174.600 3.100 ;
        RECT 175.800 0.800 176.200 3.100 ;
        RECT 176.600 0.800 177.000 5.100 ;
        RECT 179.000 0.800 179.400 3.100 ;
        RECT 180.600 0.800 181.000 3.100 ;
        RECT 182.200 0.800 182.600 4.500 ;
        RECT 184.600 0.800 185.000 5.100 ;
        RECT 187.800 0.800 188.200 4.500 ;
        RECT 190.200 0.800 190.600 5.100 ;
        RECT 195.000 0.800 195.400 4.500 ;
        RECT 197.400 0.800 197.800 5.100 ;
        RECT 200.600 0.800 201.000 5.000 ;
        RECT 203.400 0.800 203.800 3.100 ;
        RECT 205.000 0.800 205.400 3.100 ;
        RECT 207.800 0.800 208.200 5.100 ;
        RECT 210.200 0.800 210.600 5.100 ;
        RECT 213.000 0.800 213.400 3.100 ;
        RECT 214.600 0.800 215.000 3.100 ;
        RECT 217.400 0.800 217.800 5.000 ;
        RECT 219.000 0.800 219.400 3.100 ;
        RECT 220.600 0.800 221.000 3.100 ;
        RECT 222.200 0.800 222.600 5.100 ;
        RECT 225.000 0.800 225.400 3.100 ;
        RECT 226.600 0.800 227.000 3.100 ;
        RECT 229.400 0.800 229.800 5.000 ;
        RECT 0.200 0.200 231.000 0.800 ;
      LAYER via1 ;
        RECT 37.800 200.300 38.200 200.700 ;
        RECT 38.500 200.300 38.900 200.700 ;
        RECT 139.400 200.300 139.800 200.700 ;
        RECT 140.100 200.300 140.500 200.700 ;
        RECT 37.800 180.300 38.200 180.700 ;
        RECT 38.500 180.300 38.900 180.700 ;
        RECT 139.400 180.300 139.800 180.700 ;
        RECT 140.100 180.300 140.500 180.700 ;
        RECT 37.800 160.300 38.200 160.700 ;
        RECT 38.500 160.300 38.900 160.700 ;
        RECT 139.400 160.300 139.800 160.700 ;
        RECT 140.100 160.300 140.500 160.700 ;
        RECT 37.800 140.300 38.200 140.700 ;
        RECT 38.500 140.300 38.900 140.700 ;
        RECT 139.400 140.300 139.800 140.700 ;
        RECT 140.100 140.300 140.500 140.700 ;
        RECT 37.800 120.300 38.200 120.700 ;
        RECT 38.500 120.300 38.900 120.700 ;
        RECT 139.400 120.300 139.800 120.700 ;
        RECT 140.100 120.300 140.500 120.700 ;
        RECT 37.800 100.300 38.200 100.700 ;
        RECT 38.500 100.300 38.900 100.700 ;
        RECT 139.400 100.300 139.800 100.700 ;
        RECT 140.100 100.300 140.500 100.700 ;
        RECT 37.800 80.300 38.200 80.700 ;
        RECT 38.500 80.300 38.900 80.700 ;
        RECT 139.400 80.300 139.800 80.700 ;
        RECT 140.100 80.300 140.500 80.700 ;
        RECT 37.800 60.300 38.200 60.700 ;
        RECT 38.500 60.300 38.900 60.700 ;
        RECT 139.400 60.300 139.800 60.700 ;
        RECT 140.100 60.300 140.500 60.700 ;
        RECT 37.800 40.300 38.200 40.700 ;
        RECT 38.500 40.300 38.900 40.700 ;
        RECT 139.400 40.300 139.800 40.700 ;
        RECT 140.100 40.300 140.500 40.700 ;
        RECT 37.800 20.300 38.200 20.700 ;
        RECT 38.500 20.300 38.900 20.700 ;
        RECT 139.400 20.300 139.800 20.700 ;
        RECT 140.100 20.300 140.500 20.700 ;
        RECT 37.800 0.300 38.200 0.700 ;
        RECT 38.500 0.300 38.900 0.700 ;
        RECT 139.400 0.300 139.800 0.700 ;
        RECT 140.100 0.300 140.500 0.700 ;
      LAYER metal2 ;
        RECT 37.600 200.300 39.200 200.700 ;
        RECT 139.200 200.300 140.800 200.700 ;
        RECT 37.600 180.300 39.200 180.700 ;
        RECT 139.200 180.300 140.800 180.700 ;
        RECT 37.600 160.300 39.200 160.700 ;
        RECT 139.200 160.300 140.800 160.700 ;
        RECT 37.600 140.300 39.200 140.700 ;
        RECT 139.200 140.300 140.800 140.700 ;
        RECT 37.600 120.300 39.200 120.700 ;
        RECT 139.200 120.300 140.800 120.700 ;
        RECT 37.600 100.300 39.200 100.700 ;
        RECT 139.200 100.300 140.800 100.700 ;
        RECT 37.600 80.300 39.200 80.700 ;
        RECT 139.200 80.300 140.800 80.700 ;
        RECT 37.600 60.300 39.200 60.700 ;
        RECT 139.200 60.300 140.800 60.700 ;
        RECT 37.600 40.300 39.200 40.700 ;
        RECT 139.200 40.300 140.800 40.700 ;
        RECT 37.600 20.300 39.200 20.700 ;
        RECT 139.200 20.300 140.800 20.700 ;
        RECT 37.600 0.300 39.200 0.700 ;
        RECT 139.200 0.300 140.800 0.700 ;
      LAYER via2 ;
        RECT 37.800 200.300 38.200 200.700 ;
        RECT 38.500 200.300 38.900 200.700 ;
        RECT 139.400 200.300 139.800 200.700 ;
        RECT 140.100 200.300 140.500 200.700 ;
        RECT 37.800 180.300 38.200 180.700 ;
        RECT 38.500 180.300 38.900 180.700 ;
        RECT 139.400 180.300 139.800 180.700 ;
        RECT 140.100 180.300 140.500 180.700 ;
        RECT 37.800 160.300 38.200 160.700 ;
        RECT 38.500 160.300 38.900 160.700 ;
        RECT 139.400 160.300 139.800 160.700 ;
        RECT 140.100 160.300 140.500 160.700 ;
        RECT 37.800 140.300 38.200 140.700 ;
        RECT 38.500 140.300 38.900 140.700 ;
        RECT 139.400 140.300 139.800 140.700 ;
        RECT 140.100 140.300 140.500 140.700 ;
        RECT 37.800 120.300 38.200 120.700 ;
        RECT 38.500 120.300 38.900 120.700 ;
        RECT 139.400 120.300 139.800 120.700 ;
        RECT 140.100 120.300 140.500 120.700 ;
        RECT 37.800 100.300 38.200 100.700 ;
        RECT 38.500 100.300 38.900 100.700 ;
        RECT 139.400 100.300 139.800 100.700 ;
        RECT 140.100 100.300 140.500 100.700 ;
        RECT 37.800 80.300 38.200 80.700 ;
        RECT 38.500 80.300 38.900 80.700 ;
        RECT 139.400 80.300 139.800 80.700 ;
        RECT 140.100 80.300 140.500 80.700 ;
        RECT 37.800 60.300 38.200 60.700 ;
        RECT 38.500 60.300 38.900 60.700 ;
        RECT 139.400 60.300 139.800 60.700 ;
        RECT 140.100 60.300 140.500 60.700 ;
        RECT 37.800 40.300 38.200 40.700 ;
        RECT 38.500 40.300 38.900 40.700 ;
        RECT 139.400 40.300 139.800 40.700 ;
        RECT 140.100 40.300 140.500 40.700 ;
        RECT 37.800 20.300 38.200 20.700 ;
        RECT 38.500 20.300 38.900 20.700 ;
        RECT 139.400 20.300 139.800 20.700 ;
        RECT 140.100 20.300 140.500 20.700 ;
        RECT 37.800 0.300 38.200 0.700 ;
        RECT 38.500 0.300 38.900 0.700 ;
        RECT 139.400 0.300 139.800 0.700 ;
        RECT 140.100 0.300 140.500 0.700 ;
      LAYER metal3 ;
        RECT 37.600 200.300 39.200 200.700 ;
        RECT 139.200 200.300 140.800 200.700 ;
        RECT 37.600 180.300 39.200 180.700 ;
        RECT 139.200 180.300 140.800 180.700 ;
        RECT 37.600 160.300 39.200 160.700 ;
        RECT 139.200 160.300 140.800 160.700 ;
        RECT 37.600 140.300 39.200 140.700 ;
        RECT 139.200 140.300 140.800 140.700 ;
        RECT 37.600 120.300 39.200 120.700 ;
        RECT 139.200 120.300 140.800 120.700 ;
        RECT 37.600 100.300 39.200 100.700 ;
        RECT 139.200 100.300 140.800 100.700 ;
        RECT 37.600 80.300 39.200 80.700 ;
        RECT 139.200 80.300 140.800 80.700 ;
        RECT 37.600 60.300 39.200 60.700 ;
        RECT 139.200 60.300 140.800 60.700 ;
        RECT 37.600 40.300 39.200 40.700 ;
        RECT 139.200 40.300 140.800 40.700 ;
        RECT 37.600 20.300 39.200 20.700 ;
        RECT 139.200 20.300 140.800 20.700 ;
        RECT 37.600 0.300 39.200 0.700 ;
        RECT 139.200 0.300 140.800 0.700 ;
      LAYER via3 ;
        RECT 37.800 200.300 38.200 200.700 ;
        RECT 38.600 200.300 39.000 200.700 ;
        RECT 139.400 200.300 139.800 200.700 ;
        RECT 140.200 200.300 140.600 200.700 ;
        RECT 37.800 180.300 38.200 180.700 ;
        RECT 38.600 180.300 39.000 180.700 ;
        RECT 139.400 180.300 139.800 180.700 ;
        RECT 140.200 180.300 140.600 180.700 ;
        RECT 37.800 160.300 38.200 160.700 ;
        RECT 38.600 160.300 39.000 160.700 ;
        RECT 139.400 160.300 139.800 160.700 ;
        RECT 140.200 160.300 140.600 160.700 ;
        RECT 37.800 140.300 38.200 140.700 ;
        RECT 38.600 140.300 39.000 140.700 ;
        RECT 139.400 140.300 139.800 140.700 ;
        RECT 140.200 140.300 140.600 140.700 ;
        RECT 37.800 120.300 38.200 120.700 ;
        RECT 38.600 120.300 39.000 120.700 ;
        RECT 139.400 120.300 139.800 120.700 ;
        RECT 140.200 120.300 140.600 120.700 ;
        RECT 37.800 100.300 38.200 100.700 ;
        RECT 38.600 100.300 39.000 100.700 ;
        RECT 139.400 100.300 139.800 100.700 ;
        RECT 140.200 100.300 140.600 100.700 ;
        RECT 37.800 80.300 38.200 80.700 ;
        RECT 38.600 80.300 39.000 80.700 ;
        RECT 139.400 80.300 139.800 80.700 ;
        RECT 140.200 80.300 140.600 80.700 ;
        RECT 37.800 60.300 38.200 60.700 ;
        RECT 38.600 60.300 39.000 60.700 ;
        RECT 139.400 60.300 139.800 60.700 ;
        RECT 140.200 60.300 140.600 60.700 ;
        RECT 37.800 40.300 38.200 40.700 ;
        RECT 38.600 40.300 39.000 40.700 ;
        RECT 139.400 40.300 139.800 40.700 ;
        RECT 140.200 40.300 140.600 40.700 ;
        RECT 37.800 20.300 38.200 20.700 ;
        RECT 38.600 20.300 39.000 20.700 ;
        RECT 139.400 20.300 139.800 20.700 ;
        RECT 140.200 20.300 140.600 20.700 ;
        RECT 37.800 0.300 38.200 0.700 ;
        RECT 38.600 0.300 39.000 0.700 ;
        RECT 139.400 0.300 139.800 0.700 ;
        RECT 140.200 0.300 140.600 0.700 ;
      LAYER metal4 ;
        RECT 37.600 200.300 39.200 200.700 ;
        RECT 139.200 200.300 140.800 200.700 ;
        RECT 37.600 180.300 39.200 180.700 ;
        RECT 139.200 180.300 140.800 180.700 ;
        RECT 37.600 160.300 39.200 160.700 ;
        RECT 139.200 160.300 140.800 160.700 ;
        RECT 37.600 140.300 39.200 140.700 ;
        RECT 139.200 140.300 140.800 140.700 ;
        RECT 37.600 120.300 39.200 120.700 ;
        RECT 139.200 120.300 140.800 120.700 ;
        RECT 37.600 100.300 39.200 100.700 ;
        RECT 139.200 100.300 140.800 100.700 ;
        RECT 37.600 80.300 39.200 80.700 ;
        RECT 139.200 80.300 140.800 80.700 ;
        RECT 37.600 60.300 39.200 60.700 ;
        RECT 139.200 60.300 140.800 60.700 ;
        RECT 37.600 40.300 39.200 40.700 ;
        RECT 139.200 40.300 140.800 40.700 ;
        RECT 37.600 20.300 39.200 20.700 ;
        RECT 139.200 20.300 140.800 20.700 ;
        RECT 37.600 0.300 39.200 0.700 ;
        RECT 139.200 0.300 140.800 0.700 ;
      LAYER via4 ;
        RECT 37.800 200.300 38.200 200.700 ;
        RECT 38.500 200.300 38.900 200.700 ;
        RECT 139.400 200.300 139.800 200.700 ;
        RECT 140.100 200.300 140.500 200.700 ;
        RECT 37.800 180.300 38.200 180.700 ;
        RECT 38.500 180.300 38.900 180.700 ;
        RECT 139.400 180.300 139.800 180.700 ;
        RECT 140.100 180.300 140.500 180.700 ;
        RECT 37.800 160.300 38.200 160.700 ;
        RECT 38.500 160.300 38.900 160.700 ;
        RECT 139.400 160.300 139.800 160.700 ;
        RECT 140.100 160.300 140.500 160.700 ;
        RECT 37.800 140.300 38.200 140.700 ;
        RECT 38.500 140.300 38.900 140.700 ;
        RECT 139.400 140.300 139.800 140.700 ;
        RECT 140.100 140.300 140.500 140.700 ;
        RECT 37.800 120.300 38.200 120.700 ;
        RECT 38.500 120.300 38.900 120.700 ;
        RECT 139.400 120.300 139.800 120.700 ;
        RECT 140.100 120.300 140.500 120.700 ;
        RECT 37.800 100.300 38.200 100.700 ;
        RECT 38.500 100.300 38.900 100.700 ;
        RECT 139.400 100.300 139.800 100.700 ;
        RECT 140.100 100.300 140.500 100.700 ;
        RECT 37.800 80.300 38.200 80.700 ;
        RECT 38.500 80.300 38.900 80.700 ;
        RECT 139.400 80.300 139.800 80.700 ;
        RECT 140.100 80.300 140.500 80.700 ;
        RECT 37.800 60.300 38.200 60.700 ;
        RECT 38.500 60.300 38.900 60.700 ;
        RECT 139.400 60.300 139.800 60.700 ;
        RECT 140.100 60.300 140.500 60.700 ;
        RECT 37.800 40.300 38.200 40.700 ;
        RECT 38.500 40.300 38.900 40.700 ;
        RECT 139.400 40.300 139.800 40.700 ;
        RECT 140.100 40.300 140.500 40.700 ;
        RECT 37.800 20.300 38.200 20.700 ;
        RECT 38.500 20.300 38.900 20.700 ;
        RECT 139.400 20.300 139.800 20.700 ;
        RECT 140.100 20.300 140.500 20.700 ;
        RECT 37.800 0.300 38.200 0.700 ;
        RECT 38.500 0.300 38.900 0.700 ;
        RECT 139.400 0.300 139.800 0.700 ;
        RECT 140.100 0.300 140.500 0.700 ;
      LAYER metal5 ;
        RECT 37.600 200.200 39.200 200.700 ;
        RECT 139.200 200.200 140.800 200.700 ;
        RECT 37.600 180.200 39.200 180.700 ;
        RECT 139.200 180.200 140.800 180.700 ;
        RECT 37.600 160.200 39.200 160.700 ;
        RECT 139.200 160.200 140.800 160.700 ;
        RECT 37.600 140.200 39.200 140.700 ;
        RECT 139.200 140.200 140.800 140.700 ;
        RECT 37.600 120.200 39.200 120.700 ;
        RECT 139.200 120.200 140.800 120.700 ;
        RECT 37.600 100.200 39.200 100.700 ;
        RECT 139.200 100.200 140.800 100.700 ;
        RECT 37.600 80.200 39.200 80.700 ;
        RECT 139.200 80.200 140.800 80.700 ;
        RECT 37.600 60.200 39.200 60.700 ;
        RECT 139.200 60.200 140.800 60.700 ;
        RECT 37.600 40.200 39.200 40.700 ;
        RECT 139.200 40.200 140.800 40.700 ;
        RECT 37.600 20.200 39.200 20.700 ;
        RECT 139.200 20.200 140.800 20.700 ;
        RECT 37.600 0.200 39.200 0.700 ;
        RECT 139.200 0.200 140.800 0.700 ;
      LAYER via5 ;
        RECT 38.600 200.200 39.100 200.700 ;
        RECT 140.200 200.200 140.700 200.700 ;
        RECT 38.600 180.200 39.100 180.700 ;
        RECT 140.200 180.200 140.700 180.700 ;
        RECT 38.600 160.200 39.100 160.700 ;
        RECT 140.200 160.200 140.700 160.700 ;
        RECT 38.600 140.200 39.100 140.700 ;
        RECT 140.200 140.200 140.700 140.700 ;
        RECT 38.600 120.200 39.100 120.700 ;
        RECT 140.200 120.200 140.700 120.700 ;
        RECT 38.600 100.200 39.100 100.700 ;
        RECT 140.200 100.200 140.700 100.700 ;
        RECT 38.600 80.200 39.100 80.700 ;
        RECT 140.200 80.200 140.700 80.700 ;
        RECT 38.600 60.200 39.100 60.700 ;
        RECT 140.200 60.200 140.700 60.700 ;
        RECT 38.600 40.200 39.100 40.700 ;
        RECT 140.200 40.200 140.700 40.700 ;
        RECT 38.600 20.200 39.100 20.700 ;
        RECT 140.200 20.200 140.700 20.700 ;
        RECT 38.600 0.200 39.100 0.700 ;
        RECT 140.200 0.200 140.700 0.700 ;
      LAYER metal6 ;
        RECT 37.600 -3.000 39.200 213.000 ;
        RECT 139.200 -3.000 140.800 213.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 210.200 231.000 210.800 ;
        RECT 0.600 207.900 1.000 210.200 ;
        RECT 2.200 207.900 2.600 210.200 ;
        RECT 3.800 207.900 4.200 210.200 ;
        RECT 5.400 207.900 5.800 210.200 ;
        RECT 7.000 207.900 7.400 210.200 ;
        RECT 7.800 207.900 8.200 210.200 ;
        RECT 9.400 207.900 9.800 210.200 ;
        RECT 11.000 207.900 11.400 210.200 ;
        RECT 12.600 207.900 13.000 210.200 ;
        RECT 14.200 207.900 14.600 210.200 ;
        RECT 15.800 207.900 16.200 210.200 ;
        RECT 18.500 208.900 19.000 210.200 ;
        RECT 20.200 208.900 20.600 210.200 ;
        RECT 23.000 208.000 23.400 210.200 ;
        RECT 25.400 208.300 25.800 210.200 ;
        RECT 29.400 208.300 29.800 210.200 ;
        RECT 31.800 207.900 32.200 210.200 ;
        RECT 34.500 208.900 35.000 210.200 ;
        RECT 36.200 208.900 36.600 210.200 ;
        RECT 39.000 208.000 39.400 210.200 ;
        RECT 42.200 207.900 42.600 210.200 ;
        RECT 43.800 207.900 44.200 210.200 ;
        RECT 46.200 207.900 46.600 210.200 ;
        RECT 48.900 208.900 49.400 210.200 ;
        RECT 50.600 208.900 51.000 210.200 ;
        RECT 53.400 208.000 53.800 210.200 ;
        RECT 55.800 208.300 56.200 210.200 ;
        RECT 59.800 208.300 60.200 210.200 ;
        RECT 61.400 207.900 61.800 210.200 ;
        RECT 63.000 207.900 63.400 210.200 ;
        RECT 65.400 207.900 65.800 210.200 ;
        RECT 68.100 208.900 68.600 210.200 ;
        RECT 69.800 208.900 70.200 210.200 ;
        RECT 72.600 208.000 73.000 210.200 ;
        RECT 75.000 208.000 75.400 210.200 ;
        RECT 77.800 208.900 78.200 210.200 ;
        RECT 79.400 208.900 79.900 210.200 ;
        RECT 82.200 207.900 82.600 210.200 ;
        RECT 84.600 208.300 85.000 210.200 ;
        RECT 88.600 208.300 89.000 210.200 ;
        RECT 92.600 207.900 93.000 210.200 ;
        RECT 95.300 208.900 95.800 210.200 ;
        RECT 97.000 208.900 97.400 210.200 ;
        RECT 99.800 208.000 100.200 210.200 ;
        RECT 102.200 207.900 102.600 210.200 ;
        RECT 104.900 208.900 105.400 210.200 ;
        RECT 106.600 208.900 107.000 210.200 ;
        RECT 109.400 208.000 109.800 210.200 ;
        RECT 111.800 208.300 112.200 210.200 ;
        RECT 115.800 208.300 116.200 210.200 ;
        RECT 118.200 208.300 118.600 210.200 ;
        RECT 121.400 208.300 121.800 210.200 ;
        RECT 124.600 207.900 125.000 210.200 ;
        RECT 127.300 208.900 127.800 210.200 ;
        RECT 129.000 208.900 129.400 210.200 ;
        RECT 131.800 208.000 132.200 210.200 ;
        RECT 133.400 207.900 133.800 210.200 ;
        RECT 135.000 207.900 135.400 210.200 ;
        RECT 136.600 207.900 137.000 210.200 ;
        RECT 138.200 207.900 138.600 210.200 ;
        RECT 139.800 207.900 140.200 210.200 ;
        RECT 143.000 207.900 143.400 210.200 ;
        RECT 145.700 208.900 146.200 210.200 ;
        RECT 147.400 208.900 147.800 210.200 ;
        RECT 150.200 208.000 150.600 210.200 ;
        RECT 152.600 208.300 153.000 210.200 ;
        RECT 156.600 207.900 157.000 210.200 ;
        RECT 158.200 207.900 158.600 210.200 ;
        RECT 159.800 207.900 160.200 210.200 ;
        RECT 161.400 208.000 161.800 210.200 ;
        RECT 164.200 208.900 164.600 210.200 ;
        RECT 165.800 208.900 166.300 210.200 ;
        RECT 168.600 207.900 169.000 210.200 ;
        RECT 171.000 208.300 171.400 210.200 ;
        RECT 175.000 207.900 175.400 210.200 ;
        RECT 176.600 207.900 177.000 210.200 ;
        RECT 179.300 208.900 179.800 210.200 ;
        RECT 181.000 208.900 181.400 210.200 ;
        RECT 183.800 208.000 184.200 210.200 ;
        RECT 185.400 207.900 185.800 210.200 ;
        RECT 187.000 207.900 187.400 210.200 ;
        RECT 188.600 207.900 189.000 210.200 ;
        RECT 191.000 207.900 191.400 210.200 ;
        RECT 192.600 207.900 193.000 210.200 ;
        RECT 194.200 207.900 194.600 210.200 ;
        RECT 195.800 207.900 196.200 210.200 ;
        RECT 197.400 207.900 197.800 210.200 ;
        RECT 198.800 207.500 199.200 210.200 ;
        RECT 201.400 207.700 201.800 210.200 ;
        RECT 203.800 208.300 204.200 210.200 ;
        RECT 207.800 207.900 208.200 210.200 ;
        RECT 208.600 207.900 209.000 210.200 ;
        RECT 211.800 208.000 212.200 210.200 ;
        RECT 214.600 208.900 215.000 210.200 ;
        RECT 216.200 208.900 216.700 210.200 ;
        RECT 219.000 207.900 219.400 210.200 ;
        RECT 222.200 207.900 222.600 210.200 ;
        RECT 223.800 208.300 224.200 210.200 ;
        RECT 226.200 207.900 226.600 210.200 ;
        RECT 227.800 207.900 228.200 210.200 ;
        RECT 229.400 207.900 229.800 210.200 ;
        RECT 1.400 190.800 1.800 193.000 ;
        RECT 4.200 190.800 4.600 192.100 ;
        RECT 5.800 190.800 6.300 192.100 ;
        RECT 8.600 190.800 9.000 193.100 ;
        RECT 11.800 190.800 12.200 192.700 ;
        RECT 15.000 190.800 15.400 192.700 ;
        RECT 18.200 190.800 18.600 192.700 ;
        RECT 21.400 190.800 21.800 192.700 ;
        RECT 23.800 190.800 24.200 192.700 ;
        RECT 27.800 190.800 28.200 192.700 ;
        RECT 30.200 190.800 30.600 193.100 ;
        RECT 32.900 190.800 33.400 192.100 ;
        RECT 34.600 190.800 35.000 192.100 ;
        RECT 37.400 190.800 37.800 193.000 ;
        RECT 41.400 190.800 41.800 193.100 ;
        RECT 44.100 190.800 44.600 192.100 ;
        RECT 45.800 190.800 46.200 192.100 ;
        RECT 48.600 190.800 49.000 193.000 ;
        RECT 51.800 190.800 52.200 192.700 ;
        RECT 54.000 190.800 54.400 193.500 ;
        RECT 56.600 190.800 57.000 193.300 ;
        RECT 59.000 190.800 59.400 192.700 ;
        RECT 62.200 190.800 62.600 193.100 ;
        RECT 64.900 190.800 65.400 192.100 ;
        RECT 66.600 190.800 67.000 192.100 ;
        RECT 69.400 190.800 69.800 193.000 ;
        RECT 71.800 190.800 72.200 192.700 ;
        RECT 75.000 190.800 75.400 192.700 ;
        RECT 79.000 190.800 79.400 192.700 ;
        RECT 82.200 190.800 82.600 192.700 ;
        RECT 84.600 190.800 85.000 192.700 ;
        RECT 87.800 190.800 88.200 192.700 ;
        RECT 92.600 190.800 93.000 193.100 ;
        RECT 95.300 190.800 95.800 192.100 ;
        RECT 97.000 190.800 97.400 192.100 ;
        RECT 99.800 190.800 100.200 193.000 ;
        RECT 102.200 190.800 102.600 192.700 ;
        RECT 105.400 190.800 105.800 192.700 ;
        RECT 108.600 190.800 109.000 193.100 ;
        RECT 111.300 190.800 111.800 192.100 ;
        RECT 113.000 190.800 113.400 192.100 ;
        RECT 115.800 190.800 116.200 193.000 ;
        RECT 118.200 190.800 118.600 193.100 ;
        RECT 120.900 190.800 121.400 192.100 ;
        RECT 122.600 190.800 123.000 192.100 ;
        RECT 125.400 190.800 125.800 193.000 ;
        RECT 127.800 190.800 128.200 192.700 ;
        RECT 131.800 190.800 132.200 192.700 ;
        RECT 134.200 190.800 134.600 192.700 ;
        RECT 138.200 190.800 138.600 192.700 ;
        RECT 142.200 190.800 142.600 193.000 ;
        RECT 145.000 190.800 145.400 192.100 ;
        RECT 146.600 190.800 147.100 192.100 ;
        RECT 149.400 190.800 149.800 193.100 ;
        RECT 151.800 190.800 152.200 193.000 ;
        RECT 154.600 190.800 155.000 192.100 ;
        RECT 156.200 190.800 156.700 192.100 ;
        RECT 159.000 190.800 159.400 193.100 ;
        RECT 161.400 190.800 161.800 192.700 ;
        RECT 165.400 190.800 165.800 193.100 ;
        RECT 167.000 190.800 167.400 193.000 ;
        RECT 169.800 190.800 170.200 192.100 ;
        RECT 171.400 190.800 171.900 192.100 ;
        RECT 174.200 190.800 174.600 193.100 ;
        RECT 176.600 190.800 177.000 192.700 ;
        RECT 180.600 190.800 181.000 193.100 ;
        RECT 182.000 190.800 182.400 193.500 ;
        RECT 184.600 190.800 185.000 193.300 ;
        RECT 187.000 190.800 187.400 192.700 ;
        RECT 191.000 190.800 191.400 193.100 ;
        RECT 194.200 190.800 194.600 193.000 ;
        RECT 197.000 190.800 197.400 192.100 ;
        RECT 198.600 190.800 199.100 192.100 ;
        RECT 201.400 190.800 201.800 193.100 ;
        RECT 203.800 190.800 204.200 192.700 ;
        RECT 207.800 190.800 208.200 193.100 ;
        RECT 209.400 190.800 209.800 193.000 ;
        RECT 212.200 190.800 212.600 192.100 ;
        RECT 213.800 190.800 214.300 192.100 ;
        RECT 216.600 190.800 217.000 193.100 ;
        RECT 219.000 190.800 219.400 192.700 ;
        RECT 222.200 190.800 222.600 193.000 ;
        RECT 225.000 190.800 225.400 192.100 ;
        RECT 226.600 190.800 227.100 192.100 ;
        RECT 229.400 190.800 229.800 193.100 ;
        RECT 0.200 190.200 231.000 190.800 ;
        RECT 1.400 187.900 1.800 190.200 ;
        RECT 4.100 188.900 4.600 190.200 ;
        RECT 5.800 188.900 6.200 190.200 ;
        RECT 8.600 188.000 9.000 190.200 ;
        RECT 11.800 188.300 12.200 190.200 ;
        RECT 15.000 188.300 15.400 190.200 ;
        RECT 17.400 187.900 17.800 190.200 ;
        RECT 20.100 188.900 20.600 190.200 ;
        RECT 21.800 188.900 22.200 190.200 ;
        RECT 24.600 188.000 25.000 190.200 ;
        RECT 27.000 188.300 27.400 190.200 ;
        RECT 31.000 188.300 31.400 190.200 ;
        RECT 33.400 188.300 33.800 190.200 ;
        RECT 38.000 187.500 38.400 190.200 ;
        RECT 40.600 187.700 41.000 190.200 ;
        RECT 43.000 187.900 43.400 190.200 ;
        RECT 45.700 188.900 46.200 190.200 ;
        RECT 47.400 188.900 47.800 190.200 ;
        RECT 50.200 188.000 50.600 190.200 ;
        RECT 52.600 188.300 53.000 190.200 ;
        RECT 56.600 188.300 57.000 190.200 ;
        RECT 59.800 188.300 60.200 190.200 ;
        RECT 62.200 187.700 62.600 190.200 ;
        RECT 64.800 187.500 65.200 190.200 ;
        RECT 67.800 188.300 68.200 190.200 ;
        RECT 70.200 187.900 70.600 190.200 ;
        RECT 71.800 187.900 72.200 190.200 ;
        RECT 73.200 187.500 73.600 190.200 ;
        RECT 75.800 187.700 76.200 190.200 ;
        RECT 78.200 188.000 78.600 190.200 ;
        RECT 81.000 188.900 81.400 190.200 ;
        RECT 82.600 188.900 83.100 190.200 ;
        RECT 85.400 187.900 85.800 190.200 ;
        RECT 88.600 188.300 89.000 190.200 ;
        RECT 93.400 188.300 93.800 190.200 ;
        RECT 95.800 187.700 96.200 190.200 ;
        RECT 98.400 187.500 98.800 190.200 ;
        RECT 100.600 187.700 101.000 190.200 ;
        RECT 103.200 187.500 103.600 190.200 ;
        RECT 105.200 187.500 105.600 190.200 ;
        RECT 107.800 187.700 108.200 190.200 ;
        RECT 109.400 187.900 109.800 190.200 ;
        RECT 111.000 187.900 111.400 190.200 ;
        RECT 113.400 187.900 113.800 190.200 ;
        RECT 115.000 187.900 115.400 190.200 ;
        RECT 116.600 188.300 117.000 190.200 ;
        RECT 120.600 188.300 121.000 190.200 ;
        RECT 123.000 188.000 123.400 190.200 ;
        RECT 125.800 188.900 126.200 190.200 ;
        RECT 127.400 188.900 127.900 190.200 ;
        RECT 130.200 187.900 130.600 190.200 ;
        RECT 131.800 187.900 132.200 190.200 ;
        RECT 133.400 187.900 133.800 190.200 ;
        RECT 134.800 187.500 135.200 190.200 ;
        RECT 137.400 187.700 137.800 190.200 ;
        RECT 141.400 188.300 141.800 190.200 ;
        RECT 144.600 188.300 145.000 190.200 ;
        RECT 147.800 188.300 148.200 190.200 ;
        RECT 151.000 187.900 151.400 190.200 ;
        RECT 153.700 188.900 154.200 190.200 ;
        RECT 155.400 188.900 155.800 190.200 ;
        RECT 158.200 188.000 158.600 190.200 ;
        RECT 159.800 187.900 160.200 190.200 ;
        RECT 163.800 188.300 164.200 190.200 ;
        RECT 166.200 188.900 166.600 190.200 ;
        RECT 167.800 188.000 168.200 190.200 ;
        RECT 170.600 188.900 171.000 190.200 ;
        RECT 172.200 188.900 172.700 190.200 ;
        RECT 175.000 187.900 175.400 190.200 ;
        RECT 176.600 187.900 177.000 190.200 ;
        RECT 180.600 188.300 181.000 190.200 ;
        RECT 183.000 187.700 183.400 190.200 ;
        RECT 185.600 187.500 186.000 190.200 ;
        RECT 187.800 187.700 188.200 190.200 ;
        RECT 190.400 187.500 190.800 190.200 ;
        RECT 194.200 187.700 194.600 190.200 ;
        RECT 196.800 187.500 197.200 190.200 ;
        RECT 199.000 187.700 199.400 190.200 ;
        RECT 201.600 187.500 202.000 190.200 ;
        RECT 203.800 187.700 204.200 190.200 ;
        RECT 206.400 187.500 206.800 190.200 ;
        RECT 208.600 188.000 209.000 190.200 ;
        RECT 211.400 188.900 211.800 190.200 ;
        RECT 213.000 188.900 213.500 190.200 ;
        RECT 215.800 187.900 216.200 190.200 ;
        RECT 217.400 187.900 217.800 190.200 ;
        RECT 221.400 188.300 221.800 190.200 ;
        RECT 223.000 187.900 223.400 190.200 ;
        RECT 227.000 188.300 227.400 190.200 ;
        RECT 0.600 170.800 1.000 173.100 ;
        RECT 2.200 170.800 2.600 173.100 ;
        RECT 3.800 170.800 4.200 173.100 ;
        RECT 5.400 170.800 5.800 173.100 ;
        RECT 7.000 170.800 7.400 173.100 ;
        RECT 8.600 170.800 9.000 173.000 ;
        RECT 11.400 170.800 11.800 172.100 ;
        RECT 13.000 170.800 13.500 172.100 ;
        RECT 15.800 170.800 16.200 173.100 ;
        RECT 17.400 170.800 17.800 173.100 ;
        RECT 19.000 170.800 19.400 173.100 ;
        RECT 20.600 170.800 21.000 173.100 ;
        RECT 22.200 170.800 22.600 173.100 ;
        RECT 23.800 170.800 24.200 173.100 ;
        RECT 25.400 170.800 25.800 173.100 ;
        RECT 28.100 170.800 28.600 172.100 ;
        RECT 29.800 170.800 30.200 172.100 ;
        RECT 32.600 170.800 33.000 173.000 ;
        RECT 35.800 170.800 36.200 172.700 ;
        RECT 39.600 170.800 40.000 173.500 ;
        RECT 42.200 170.800 42.600 173.300 ;
        RECT 44.600 170.800 45.000 173.100 ;
        RECT 47.300 170.800 47.800 172.100 ;
        RECT 49.000 170.800 49.400 172.100 ;
        RECT 51.800 170.800 52.200 173.000 ;
        RECT 54.200 170.800 54.600 172.700 ;
        RECT 58.200 170.800 58.600 172.700 ;
        RECT 60.600 170.800 61.000 173.300 ;
        RECT 63.200 170.800 63.600 173.500 ;
        RECT 65.200 170.800 65.600 173.500 ;
        RECT 67.800 170.800 68.200 173.300 ;
        RECT 70.200 170.800 70.600 173.300 ;
        RECT 72.800 170.800 73.200 173.500 ;
        RECT 75.000 170.800 75.400 173.100 ;
        RECT 76.600 170.800 77.000 173.100 ;
        RECT 78.200 170.800 78.600 173.100 ;
        RECT 80.900 170.800 81.400 172.100 ;
        RECT 82.600 170.800 83.000 172.100 ;
        RECT 85.400 170.800 85.800 173.000 ;
        RECT 87.800 170.800 88.200 172.700 ;
        RECT 93.400 170.800 93.800 172.700 ;
        RECT 95.000 170.800 95.400 173.100 ;
        RECT 96.600 170.800 97.000 173.100 ;
        RECT 98.200 170.800 98.600 173.100 ;
        RECT 99.000 170.800 99.400 173.100 ;
        RECT 101.400 170.800 101.800 173.100 ;
        RECT 103.000 170.800 103.400 173.100 ;
        RECT 104.600 170.800 105.000 172.700 ;
        RECT 108.600 170.800 109.000 172.700 ;
        RECT 111.000 170.800 111.400 172.700 ;
        RECT 114.200 170.800 114.600 172.700 ;
        RECT 117.400 170.800 117.800 173.100 ;
        RECT 120.100 170.800 120.600 172.100 ;
        RECT 121.800 170.800 122.200 172.100 ;
        RECT 124.600 170.800 125.000 173.000 ;
        RECT 126.800 170.800 127.200 173.500 ;
        RECT 129.400 170.800 129.800 173.300 ;
        RECT 132.600 170.800 133.000 173.100 ;
        RECT 134.000 170.800 134.400 173.500 ;
        RECT 136.600 170.800 137.000 173.300 ;
        RECT 139.000 170.800 139.400 172.700 ;
        RECT 143.800 170.800 144.200 173.000 ;
        RECT 146.600 170.800 147.000 172.100 ;
        RECT 148.200 170.800 148.700 172.100 ;
        RECT 151.000 170.800 151.400 173.100 ;
        RECT 153.400 170.800 153.800 172.700 ;
        RECT 157.400 170.800 157.800 173.100 ;
        RECT 159.000 170.800 159.400 172.700 ;
        RECT 163.000 170.800 163.400 173.100 ;
        RECT 164.600 170.800 165.000 173.100 ;
        RECT 167.300 170.800 167.800 172.100 ;
        RECT 169.000 170.800 169.400 172.100 ;
        RECT 171.800 170.800 172.200 173.000 ;
        RECT 174.200 170.800 174.600 173.300 ;
        RECT 176.800 170.800 177.200 173.500 ;
        RECT 179.000 170.800 179.400 173.100 ;
        RECT 180.600 170.800 181.000 173.100 ;
        RECT 181.400 170.800 181.800 173.100 ;
        RECT 183.800 170.800 184.200 173.100 ;
        RECT 187.800 170.800 188.200 173.100 ;
        RECT 189.400 170.800 189.800 173.300 ;
        RECT 192.000 170.800 192.400 173.500 ;
        RECT 196.600 170.800 197.000 173.100 ;
        RECT 199.000 170.800 199.400 172.700 ;
        RECT 201.400 170.800 201.800 173.000 ;
        RECT 204.200 170.800 204.600 172.100 ;
        RECT 205.800 170.800 206.300 172.100 ;
        RECT 208.600 170.800 209.000 173.100 ;
        RECT 211.000 170.800 211.400 173.100 ;
        RECT 212.600 170.800 213.000 173.100 ;
        RECT 213.400 170.800 213.800 173.100 ;
        RECT 216.600 170.800 217.000 173.000 ;
        RECT 219.400 170.800 219.800 172.100 ;
        RECT 221.000 170.800 221.500 172.100 ;
        RECT 223.800 170.800 224.200 173.100 ;
        RECT 225.400 170.800 225.800 173.100 ;
        RECT 229.400 170.800 229.800 172.700 ;
        RECT 0.200 170.200 231.000 170.800 ;
        RECT 1.400 167.900 1.800 170.200 ;
        RECT 4.100 168.900 4.600 170.200 ;
        RECT 5.800 168.900 6.200 170.200 ;
        RECT 8.600 168.000 9.000 170.200 ;
        RECT 10.200 168.900 10.600 170.200 ;
        RECT 11.800 167.900 12.200 170.200 ;
        RECT 15.800 168.300 16.200 170.200 ;
        RECT 18.200 167.900 18.600 170.200 ;
        RECT 19.800 167.900 20.200 170.200 ;
        RECT 21.400 167.900 21.800 170.200 ;
        RECT 24.100 168.900 24.600 170.200 ;
        RECT 25.800 168.900 26.200 170.200 ;
        RECT 28.600 168.000 29.000 170.200 ;
        RECT 30.200 167.900 30.600 170.200 ;
        RECT 34.200 168.300 34.600 170.200 ;
        RECT 38.200 167.900 38.600 170.200 ;
        RECT 40.900 168.900 41.400 170.200 ;
        RECT 42.600 168.900 43.000 170.200 ;
        RECT 45.400 168.000 45.800 170.200 ;
        RECT 47.600 167.500 48.000 170.200 ;
        RECT 50.200 167.700 50.600 170.200 ;
        RECT 52.600 168.300 53.000 170.200 ;
        RECT 56.600 168.300 57.000 170.200 ;
        RECT 59.000 167.900 59.400 170.200 ;
        RECT 60.600 167.900 61.000 170.200 ;
        RECT 62.200 167.700 62.600 170.200 ;
        RECT 64.800 167.500 65.200 170.200 ;
        RECT 67.000 167.700 67.400 170.200 ;
        RECT 69.600 167.500 70.000 170.200 ;
        RECT 71.800 168.300 72.200 170.200 ;
        RECT 75.800 168.300 76.200 170.200 ;
        RECT 78.200 167.900 78.600 170.200 ;
        RECT 80.900 168.900 81.400 170.200 ;
        RECT 82.600 168.900 83.000 170.200 ;
        RECT 85.400 168.000 85.800 170.200 ;
        RECT 87.800 167.900 88.200 170.200 ;
        RECT 89.400 167.900 89.800 170.200 ;
        RECT 93.400 168.300 93.800 170.200 ;
        RECT 95.800 167.700 96.200 170.200 ;
        RECT 98.400 167.500 98.800 170.200 ;
        RECT 100.600 168.300 101.000 170.200 ;
        RECT 103.800 167.900 104.200 170.200 ;
        RECT 105.400 167.900 105.800 170.200 ;
        RECT 107.000 167.900 107.400 170.200 ;
        RECT 109.700 168.900 110.200 170.200 ;
        RECT 111.400 168.900 111.800 170.200 ;
        RECT 114.200 168.000 114.600 170.200 ;
        RECT 116.600 167.700 117.000 170.200 ;
        RECT 119.200 167.500 119.600 170.200 ;
        RECT 121.200 167.500 121.600 170.200 ;
        RECT 123.800 167.700 124.200 170.200 ;
        RECT 126.000 167.500 126.400 170.200 ;
        RECT 128.600 167.700 129.000 170.200 ;
        RECT 130.800 167.500 131.200 170.200 ;
        RECT 133.400 167.700 133.800 170.200 ;
        RECT 135.600 167.500 136.000 170.200 ;
        RECT 138.200 167.700 138.600 170.200 ;
        RECT 142.200 167.900 142.600 170.200 ;
        RECT 144.900 168.900 145.400 170.200 ;
        RECT 146.600 168.900 147.000 170.200 ;
        RECT 149.400 168.000 149.800 170.200 ;
        RECT 151.800 168.900 152.200 170.200 ;
        RECT 154.200 168.300 154.600 170.200 ;
        RECT 155.800 167.900 156.200 170.200 ;
        RECT 159.000 167.900 159.400 170.200 ;
        RECT 161.700 168.900 162.200 170.200 ;
        RECT 163.400 168.900 163.800 170.200 ;
        RECT 166.200 168.000 166.600 170.200 ;
        RECT 167.800 167.900 168.200 170.200 ;
        RECT 171.800 168.300 172.200 170.200 ;
        RECT 175.800 166.900 176.200 170.200 ;
        RECT 176.600 167.900 177.000 170.200 ;
        RECT 179.800 167.900 180.200 170.200 ;
        RECT 181.400 167.900 181.800 170.200 ;
        RECT 183.000 168.300 183.400 170.200 ;
        RECT 186.200 167.900 186.600 170.200 ;
        RECT 188.900 168.900 189.400 170.200 ;
        RECT 190.600 168.900 191.000 170.200 ;
        RECT 193.400 168.000 193.800 170.200 ;
        RECT 197.400 167.700 197.800 170.200 ;
        RECT 200.000 167.500 200.400 170.200 ;
        RECT 202.200 167.700 202.600 170.200 ;
        RECT 204.800 167.500 205.200 170.200 ;
        RECT 207.000 168.000 207.400 170.200 ;
        RECT 209.800 168.900 210.200 170.200 ;
        RECT 211.400 168.900 211.900 170.200 ;
        RECT 214.200 167.900 214.600 170.200 ;
        RECT 215.800 167.900 216.200 170.200 ;
        RECT 219.800 168.300 220.200 170.200 ;
        RECT 221.400 167.900 221.800 170.200 ;
        RECT 223.800 167.900 224.200 170.200 ;
        RECT 225.400 167.900 225.800 170.200 ;
        RECT 227.000 167.900 227.400 170.200 ;
        RECT 228.600 167.900 229.000 170.200 ;
        RECT 230.200 167.900 230.600 170.200 ;
        RECT 2.200 150.800 2.600 152.700 ;
        RECT 5.400 150.800 5.800 153.100 ;
        RECT 7.000 150.800 7.400 153.100 ;
        RECT 8.600 150.800 9.000 153.100 ;
        RECT 10.200 150.800 10.600 152.700 ;
        RECT 13.400 150.800 13.800 153.100 ;
        RECT 16.100 150.800 16.600 152.100 ;
        RECT 17.800 150.800 18.200 152.100 ;
        RECT 20.600 150.800 21.000 153.000 ;
        RECT 23.000 150.800 23.400 153.100 ;
        RECT 25.700 150.800 26.200 152.100 ;
        RECT 27.400 150.800 27.800 152.100 ;
        RECT 30.200 150.800 30.600 153.000 ;
        RECT 32.600 150.800 33.000 153.100 ;
        RECT 35.300 150.800 35.800 152.100 ;
        RECT 37.000 150.800 37.400 152.100 ;
        RECT 39.800 150.800 40.200 153.000 ;
        RECT 43.800 150.800 44.200 152.700 ;
        RECT 47.800 150.800 48.200 152.700 ;
        RECT 50.000 150.800 50.400 153.500 ;
        RECT 52.600 150.800 53.000 153.300 ;
        RECT 55.000 150.800 55.400 153.100 ;
        RECT 57.700 150.800 58.200 152.100 ;
        RECT 59.400 150.800 59.800 152.100 ;
        RECT 62.200 150.800 62.600 153.000 ;
        RECT 64.600 150.800 65.000 152.700 ;
        RECT 68.600 150.800 69.000 153.100 ;
        RECT 69.400 150.800 69.800 152.100 ;
        RECT 71.000 150.800 71.400 153.100 ;
        RECT 72.600 150.800 73.000 153.100 ;
        RECT 75.000 150.800 75.400 153.100 ;
        RECT 77.700 150.800 78.200 152.100 ;
        RECT 79.400 150.800 79.800 152.100 ;
        RECT 82.200 150.800 82.600 153.000 ;
        RECT 84.600 150.800 85.000 152.700 ;
        RECT 89.400 150.800 89.800 153.100 ;
        RECT 92.100 150.800 92.600 152.100 ;
        RECT 93.800 150.800 94.200 152.100 ;
        RECT 96.600 150.800 97.000 153.000 ;
        RECT 99.800 150.800 100.200 153.100 ;
        RECT 102.200 150.800 102.600 152.700 ;
        RECT 105.400 150.800 105.800 153.100 ;
        RECT 107.000 150.800 107.400 153.100 ;
        RECT 109.700 150.800 110.200 152.100 ;
        RECT 111.400 150.800 111.800 152.100 ;
        RECT 114.200 150.800 114.600 153.000 ;
        RECT 116.600 150.800 117.000 153.100 ;
        RECT 119.300 150.800 119.800 152.100 ;
        RECT 121.000 150.800 121.400 152.100 ;
        RECT 123.800 150.800 124.200 153.000 ;
        RECT 125.400 150.800 125.800 153.100 ;
        RECT 127.000 150.800 127.400 153.100 ;
        RECT 130.200 150.800 130.600 153.100 ;
        RECT 131.800 150.800 132.200 153.100 ;
        RECT 134.500 150.800 135.000 152.100 ;
        RECT 136.200 150.800 136.600 152.100 ;
        RECT 139.000 150.800 139.400 153.000 ;
        RECT 142.200 150.800 142.600 152.100 ;
        RECT 145.400 150.800 145.800 153.100 ;
        RECT 147.000 150.800 147.400 152.700 ;
        RECT 149.700 150.800 150.100 153.100 ;
        RECT 151.800 150.800 152.200 152.100 ;
        RECT 152.600 150.800 153.000 153.100 ;
        RECT 154.200 150.800 154.600 153.100 ;
        RECT 155.800 150.800 156.200 153.100 ;
        RECT 158.200 150.800 158.600 153.100 ;
        RECT 161.400 150.800 161.800 153.000 ;
        RECT 164.200 150.800 164.600 152.100 ;
        RECT 165.800 150.800 166.300 152.100 ;
        RECT 168.600 150.800 169.000 153.100 ;
        RECT 171.800 150.800 172.200 152.700 ;
        RECT 174.200 150.800 174.600 153.300 ;
        RECT 176.800 150.800 177.200 153.500 ;
        RECT 178.200 150.800 178.600 153.100 ;
        RECT 181.400 150.800 181.800 152.700 ;
        RECT 185.400 150.800 185.800 153.100 ;
        RECT 187.000 150.800 187.400 153.000 ;
        RECT 189.800 150.800 190.200 152.100 ;
        RECT 191.400 150.800 191.900 152.100 ;
        RECT 194.200 150.800 194.600 153.100 ;
        RECT 197.400 150.800 197.800 153.100 ;
        RECT 200.600 150.800 201.000 153.300 ;
        RECT 203.200 150.800 203.600 153.500 ;
        RECT 204.600 150.800 205.000 153.100 ;
        RECT 206.200 150.800 206.600 153.100 ;
        RECT 208.600 150.800 209.000 152.700 ;
        RECT 212.600 150.800 213.000 153.100 ;
        RECT 215.000 150.800 215.400 152.700 ;
        RECT 217.400 150.800 217.800 153.000 ;
        RECT 220.200 150.800 220.600 152.100 ;
        RECT 221.800 150.800 222.300 152.100 ;
        RECT 224.600 150.800 225.000 153.100 ;
        RECT 227.800 150.800 228.200 152.700 ;
        RECT 0.200 150.200 231.000 150.800 ;
        RECT 1.400 147.900 1.800 150.200 ;
        RECT 4.100 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.200 150.200 ;
        RECT 8.600 148.000 9.000 150.200 ;
        RECT 11.000 148.300 11.400 150.200 ;
        RECT 15.000 147.900 15.400 150.200 ;
        RECT 15.800 147.900 16.200 150.200 ;
        RECT 19.800 147.900 20.200 150.200 ;
        RECT 21.400 148.300 21.800 150.200 ;
        RECT 23.800 148.900 24.200 150.200 ;
        RECT 25.400 148.900 25.800 150.200 ;
        RECT 27.800 148.300 28.200 150.200 ;
        RECT 32.600 148.300 33.000 150.200 ;
        RECT 35.000 147.900 35.400 150.200 ;
        RECT 36.600 147.900 37.000 150.200 ;
        RECT 39.800 148.300 40.200 150.200 ;
        RECT 43.800 148.300 44.200 150.200 ;
        RECT 47.000 148.300 47.400 150.200 ;
        RECT 48.600 147.900 49.000 150.200 ;
        RECT 50.200 147.900 50.600 150.200 ;
        RECT 52.600 147.900 53.000 150.200 ;
        RECT 54.200 147.900 54.600 150.200 ;
        RECT 55.800 147.900 56.200 150.200 ;
        RECT 58.500 148.900 59.000 150.200 ;
        RECT 60.200 148.900 60.600 150.200 ;
        RECT 63.000 148.000 63.400 150.200 ;
        RECT 65.400 148.300 65.800 150.200 ;
        RECT 69.400 148.300 69.800 150.200 ;
        RECT 71.800 148.300 72.200 150.200 ;
        RECT 75.000 147.700 75.400 150.200 ;
        RECT 77.600 147.500 78.000 150.200 ;
        RECT 79.000 147.900 79.400 150.200 ;
        RECT 80.600 147.900 81.000 150.200 ;
        RECT 81.400 148.900 81.800 150.200 ;
        RECT 83.000 148.100 83.400 150.200 ;
        RECT 86.200 148.300 86.600 150.200 ;
        RECT 91.800 146.900 92.200 150.200 ;
        RECT 92.600 146.900 93.000 150.200 ;
        RECT 95.800 147.900 96.200 150.200 ;
        RECT 97.400 147.900 97.800 150.200 ;
        RECT 98.200 146.900 98.600 150.200 ;
        RECT 101.400 148.900 101.800 150.200 ;
        RECT 103.000 148.900 103.400 150.200 ;
        RECT 103.800 146.900 104.200 150.200 ;
        RECT 107.000 147.900 107.400 150.200 ;
        RECT 108.600 147.900 109.000 150.200 ;
        RECT 110.200 148.900 110.600 150.200 ;
        RECT 111.800 148.900 112.200 150.200 ;
        RECT 112.600 148.900 113.000 150.200 ;
        RECT 114.200 148.900 114.600 150.200 ;
        RECT 115.800 148.100 116.200 150.200 ;
        RECT 117.400 148.900 117.800 150.200 ;
        RECT 119.000 148.300 119.400 150.200 ;
        RECT 123.000 147.900 123.400 150.200 ;
        RECT 125.400 147.900 125.800 150.200 ;
        RECT 127.800 147.900 128.200 150.200 ;
        RECT 129.400 148.300 129.800 150.200 ;
        RECT 131.800 148.900 132.200 150.200 ;
        RECT 135.000 148.300 135.400 150.200 ;
        RECT 138.200 147.900 138.600 150.200 ;
        RECT 141.400 148.300 141.800 150.200 ;
        RECT 145.400 147.900 145.800 150.200 ;
        RECT 146.400 147.900 146.800 150.200 ;
        RECT 149.400 147.900 149.800 150.200 ;
        RECT 150.200 146.900 150.600 150.200 ;
        RECT 154.200 148.900 154.600 150.200 ;
        RECT 155.600 147.500 156.000 150.200 ;
        RECT 158.200 147.700 158.600 150.200 ;
        RECT 160.400 147.500 160.800 150.200 ;
        RECT 163.000 147.700 163.400 150.200 ;
        RECT 165.400 148.000 165.800 150.200 ;
        RECT 168.200 148.900 168.600 150.200 ;
        RECT 169.800 148.900 170.300 150.200 ;
        RECT 172.600 147.900 173.000 150.200 ;
        RECT 175.000 148.300 175.400 150.200 ;
        RECT 179.000 147.900 179.400 150.200 ;
        RECT 180.600 148.000 181.000 150.200 ;
        RECT 183.400 148.900 183.800 150.200 ;
        RECT 185.000 148.900 185.500 150.200 ;
        RECT 187.800 147.900 188.200 150.200 ;
        RECT 190.200 148.300 190.600 150.200 ;
        RECT 195.800 147.900 196.200 150.200 ;
        RECT 197.400 147.900 197.800 150.200 ;
        RECT 200.100 148.900 200.600 150.200 ;
        RECT 201.800 148.900 202.200 150.200 ;
        RECT 204.600 148.000 205.000 150.200 ;
        RECT 207.000 148.900 207.400 150.200 ;
        RECT 208.600 147.900 209.000 150.200 ;
        RECT 211.300 148.900 211.800 150.200 ;
        RECT 213.000 148.900 213.400 150.200 ;
        RECT 215.800 148.000 216.200 150.200 ;
        RECT 218.200 148.300 218.600 150.200 ;
        RECT 221.400 147.900 221.800 150.200 ;
        RECT 224.100 148.900 224.600 150.200 ;
        RECT 225.800 148.900 226.200 150.200 ;
        RECT 228.600 148.000 229.000 150.200 ;
        RECT 1.400 130.800 1.800 133.100 ;
        RECT 4.100 130.800 4.600 132.100 ;
        RECT 5.800 130.800 6.200 132.100 ;
        RECT 8.600 130.800 9.000 133.000 ;
        RECT 10.200 130.800 10.600 133.100 ;
        RECT 14.200 130.800 14.600 132.700 ;
        RECT 16.600 130.800 17.000 133.100 ;
        RECT 19.300 130.800 19.800 132.100 ;
        RECT 21.000 130.800 21.400 132.100 ;
        RECT 23.800 130.800 24.200 133.000 ;
        RECT 26.200 130.800 26.600 132.700 ;
        RECT 29.400 130.800 29.800 133.100 ;
        RECT 32.100 130.800 32.600 132.100 ;
        RECT 33.800 130.800 34.200 132.100 ;
        RECT 36.600 130.800 37.000 133.000 ;
        RECT 40.600 130.800 41.000 132.700 ;
        RECT 44.600 130.800 45.000 132.700 ;
        RECT 47.800 130.800 48.200 133.100 ;
        RECT 48.600 130.800 49.000 133.100 ;
        RECT 50.200 130.800 50.600 133.100 ;
        RECT 52.600 130.800 53.000 133.100 ;
        RECT 55.300 130.800 55.800 132.100 ;
        RECT 57.000 130.800 57.400 132.100 ;
        RECT 59.800 130.800 60.200 133.000 ;
        RECT 61.400 130.800 61.800 133.100 ;
        RECT 64.600 130.800 65.000 133.100 ;
        RECT 67.300 130.800 67.800 132.100 ;
        RECT 69.000 130.800 69.400 132.100 ;
        RECT 71.800 130.800 72.200 133.000 ;
        RECT 75.000 130.800 75.400 132.700 ;
        RECT 78.200 130.800 78.600 133.100 ;
        RECT 79.000 130.800 79.400 134.100 ;
        RECT 83.000 130.800 83.400 132.700 ;
        RECT 87.800 130.800 88.200 133.100 ;
        RECT 90.500 130.800 91.000 132.100 ;
        RECT 92.200 130.800 92.600 132.100 ;
        RECT 95.000 130.800 95.400 133.000 ;
        RECT 96.600 130.800 97.000 132.100 ;
        RECT 98.200 130.800 98.600 132.100 ;
        RECT 99.000 130.800 99.400 133.100 ;
        RECT 100.600 130.800 101.000 133.100 ;
        RECT 102.200 130.800 102.600 134.100 ;
        RECT 105.400 130.800 105.800 134.100 ;
        RECT 108.600 130.800 109.000 133.100 ;
        RECT 110.200 130.800 110.600 133.100 ;
        RECT 114.200 130.800 114.600 134.100 ;
        RECT 115.000 130.800 115.400 134.100 ;
        RECT 118.200 130.800 118.600 134.100 ;
        RECT 123.800 130.800 124.200 134.100 ;
        RECT 127.000 130.800 127.400 134.100 ;
        RECT 127.800 130.800 128.200 132.100 ;
        RECT 129.400 130.800 129.800 132.100 ;
        RECT 130.200 130.800 130.600 133.100 ;
        RECT 131.800 130.800 132.200 133.100 ;
        RECT 133.400 130.800 133.800 133.100 ;
        RECT 136.600 130.800 137.000 132.700 ;
        RECT 143.000 130.800 143.400 132.700 ;
        RECT 145.400 130.800 145.800 132.700 ;
        RECT 148.600 130.800 149.000 132.100 ;
        RECT 149.400 130.800 149.800 133.100 ;
        RECT 151.000 130.800 151.400 133.100 ;
        RECT 152.600 130.800 153.000 133.100 ;
        RECT 153.400 130.800 153.800 132.100 ;
        RECT 155.000 130.800 155.400 132.100 ;
        RECT 157.400 130.800 157.800 132.700 ;
        RECT 159.000 130.800 159.400 133.100 ;
        RECT 161.400 130.800 161.800 133.100 ;
        RECT 163.800 130.800 164.200 134.100 ;
        RECT 168.600 130.800 169.000 132.700 ;
        RECT 171.000 130.800 171.400 132.700 ;
        RECT 174.200 130.800 174.600 132.700 ;
        RECT 178.200 130.800 178.600 133.100 ;
        RECT 179.000 130.800 179.400 133.100 ;
        RECT 183.000 130.800 183.400 132.700 ;
        RECT 186.200 130.800 186.600 133.100 ;
        RECT 189.400 130.800 189.800 133.000 ;
        RECT 192.200 130.800 192.600 132.100 ;
        RECT 193.800 130.800 194.300 132.100 ;
        RECT 196.600 130.800 197.000 133.100 ;
        RECT 199.800 130.800 200.200 132.700 ;
        RECT 202.200 130.800 202.600 132.100 ;
        RECT 203.000 130.800 203.400 133.100 ;
        RECT 207.000 130.800 207.400 132.700 ;
        RECT 209.400 130.800 209.800 133.000 ;
        RECT 212.200 130.800 212.600 132.100 ;
        RECT 213.800 130.800 214.300 132.100 ;
        RECT 216.600 130.800 217.000 133.100 ;
        RECT 219.000 130.800 219.400 133.100 ;
        RECT 221.700 130.800 222.200 132.100 ;
        RECT 223.400 130.800 223.800 132.100 ;
        RECT 226.200 130.800 226.600 133.000 ;
        RECT 228.600 130.800 229.000 133.100 ;
        RECT 0.200 130.200 231.000 130.800 ;
        RECT 2.200 128.300 2.600 130.200 ;
        RECT 4.600 128.000 5.000 130.200 ;
        RECT 7.400 128.900 7.800 130.200 ;
        RECT 9.000 128.900 9.500 130.200 ;
        RECT 11.800 127.900 12.200 130.200 ;
        RECT 13.400 128.900 13.800 130.200 ;
        RECT 15.800 127.900 16.200 130.200 ;
        RECT 18.500 128.900 19.000 130.200 ;
        RECT 20.200 128.900 20.600 130.200 ;
        RECT 23.000 128.000 23.400 130.200 ;
        RECT 24.600 128.900 25.000 130.200 ;
        RECT 27.000 128.300 27.400 130.200 ;
        RECT 31.000 128.300 31.400 130.200 ;
        RECT 33.400 127.900 33.800 130.200 ;
        RECT 36.100 128.900 36.600 130.200 ;
        RECT 37.800 128.900 38.200 130.200 ;
        RECT 40.600 128.000 41.000 130.200 ;
        RECT 44.600 128.900 45.000 130.200 ;
        RECT 47.000 128.300 47.400 130.200 ;
        RECT 48.600 127.900 49.000 130.200 ;
        RECT 50.200 127.900 50.600 130.200 ;
        RECT 51.800 128.300 52.200 130.200 ;
        RECT 55.800 127.900 56.200 130.200 ;
        RECT 56.600 128.900 57.000 130.200 ;
        RECT 59.000 128.300 59.400 130.200 ;
        RECT 63.000 127.900 63.400 130.200 ;
        RECT 63.800 128.900 64.200 130.200 ;
        RECT 66.200 127.900 66.600 130.200 ;
        RECT 68.900 128.900 69.400 130.200 ;
        RECT 70.600 128.900 71.000 130.200 ;
        RECT 73.400 128.000 73.800 130.200 ;
        RECT 75.000 128.900 75.400 130.200 ;
        RECT 76.600 128.900 77.000 130.200 ;
        RECT 79.000 128.300 79.400 130.200 ;
        RECT 83.000 127.900 83.400 130.200 ;
        RECT 84.600 127.900 85.000 130.200 ;
        RECT 87.300 128.900 87.800 130.200 ;
        RECT 89.000 128.900 89.400 130.200 ;
        RECT 91.800 128.000 92.200 130.200 ;
        RECT 96.600 127.900 97.000 130.200 ;
        RECT 97.400 128.900 97.800 130.200 ;
        RECT 99.000 128.900 99.400 130.200 ;
        RECT 102.200 126.900 102.600 130.200 ;
        RECT 105.400 126.900 105.800 130.200 ;
        RECT 107.000 128.300 107.400 130.200 ;
        RECT 112.600 126.900 113.000 130.200 ;
        RECT 115.800 126.900 116.200 130.200 ;
        RECT 116.600 128.900 117.000 130.200 ;
        RECT 118.200 128.900 118.600 130.200 ;
        RECT 119.000 126.900 119.400 130.200 ;
        RECT 122.200 127.900 122.600 130.200 ;
        RECT 123.800 127.900 124.200 130.200 ;
        RECT 126.200 127.900 126.600 130.200 ;
        RECT 128.900 128.900 129.400 130.200 ;
        RECT 130.600 128.900 131.000 130.200 ;
        RECT 133.400 128.000 133.800 130.200 ;
        RECT 136.600 128.300 137.000 130.200 ;
        RECT 138.200 127.900 138.600 130.200 ;
        RECT 143.800 128.300 144.200 130.200 ;
        RECT 145.400 127.900 145.800 130.200 ;
        RECT 149.400 128.300 149.800 130.200 ;
        RECT 151.800 128.900 152.200 130.200 ;
        RECT 153.400 128.000 153.800 130.200 ;
        RECT 156.200 128.900 156.600 130.200 ;
        RECT 157.800 128.900 158.300 130.200 ;
        RECT 160.600 127.900 161.000 130.200 ;
        RECT 163.800 128.300 164.200 130.200 ;
        RECT 167.800 126.900 168.200 130.200 ;
        RECT 168.600 127.900 169.000 130.200 ;
        RECT 171.000 127.900 171.400 130.200 ;
        RECT 172.600 127.900 173.000 130.200 ;
        RECT 175.000 128.300 175.400 130.200 ;
        RECT 179.000 127.900 179.400 130.200 ;
        RECT 180.600 128.000 181.000 130.200 ;
        RECT 183.400 128.900 183.800 130.200 ;
        RECT 185.000 128.900 185.500 130.200 ;
        RECT 187.800 127.900 188.200 130.200 ;
        RECT 191.000 128.300 191.400 130.200 ;
        RECT 195.000 127.900 195.400 130.200 ;
        RECT 196.600 127.900 197.000 130.200 ;
        RECT 198.200 127.700 198.600 130.200 ;
        RECT 200.800 127.500 201.200 130.200 ;
        RECT 202.500 127.900 202.900 130.200 ;
        RECT 204.600 128.900 205.000 130.200 ;
        RECT 207.000 128.300 207.400 130.200 ;
        RECT 209.400 127.700 209.800 130.200 ;
        RECT 212.000 127.500 212.400 130.200 ;
        RECT 213.400 127.900 213.800 130.200 ;
        RECT 217.400 128.300 217.800 130.200 ;
        RECT 219.800 128.000 220.200 130.200 ;
        RECT 222.600 128.900 223.000 130.200 ;
        RECT 224.200 128.900 224.700 130.200 ;
        RECT 227.000 127.900 227.400 130.200 ;
        RECT 229.400 127.900 229.800 130.200 ;
        RECT 0.600 110.800 1.000 113.100 ;
        RECT 2.200 110.800 2.600 113.100 ;
        RECT 3.800 110.800 4.200 113.100 ;
        RECT 5.400 110.800 5.800 113.100 ;
        RECT 8.100 110.800 8.600 112.100 ;
        RECT 9.800 110.800 10.200 112.100 ;
        RECT 12.600 110.800 13.000 113.000 ;
        RECT 15.000 110.800 15.400 112.700 ;
        RECT 19.000 110.800 19.400 112.700 ;
        RECT 20.600 110.800 21.000 112.100 ;
        RECT 24.600 110.800 25.000 112.700 ;
        RECT 28.600 110.800 29.000 112.700 ;
        RECT 31.000 110.800 31.400 112.100 ;
        RECT 31.800 110.800 32.200 113.100 ;
        RECT 33.400 110.800 33.800 113.100 ;
        RECT 35.800 110.800 36.200 112.700 ;
        RECT 40.600 110.800 41.000 112.700 ;
        RECT 43.800 110.800 44.200 113.100 ;
        RECT 45.400 110.800 45.800 113.100 ;
        RECT 47.000 110.800 47.400 112.700 ;
        RECT 51.000 110.800 51.400 112.700 ;
        RECT 53.400 110.800 53.800 113.000 ;
        RECT 56.200 110.800 56.600 112.100 ;
        RECT 57.800 110.800 58.300 112.100 ;
        RECT 60.600 110.800 61.000 113.100 ;
        RECT 63.000 110.800 63.400 112.900 ;
        RECT 64.600 110.800 65.000 112.100 ;
        RECT 66.200 110.800 66.600 113.100 ;
        RECT 67.800 110.800 68.200 113.100 ;
        RECT 69.400 110.800 69.800 112.700 ;
        RECT 73.400 110.800 73.800 112.700 ;
        RECT 75.800 110.800 76.200 112.700 ;
        RECT 79.800 110.800 80.200 112.100 ;
        RECT 80.600 110.800 81.000 113.100 ;
        RECT 82.200 110.800 82.600 113.100 ;
        RECT 83.800 110.800 84.200 113.000 ;
        RECT 86.600 110.800 87.000 112.100 ;
        RECT 88.200 110.800 88.700 112.100 ;
        RECT 91.000 110.800 91.400 113.100 ;
        RECT 94.200 110.800 94.600 113.100 ;
        RECT 98.200 110.800 98.600 112.700 ;
        RECT 99.800 110.800 100.200 113.100 ;
        RECT 103.800 110.800 104.200 113.100 ;
        RECT 105.400 110.800 105.800 112.700 ;
        RECT 109.400 110.800 109.800 113.100 ;
        RECT 111.000 110.800 111.400 112.100 ;
        RECT 113.400 110.800 113.800 113.100 ;
        RECT 114.200 110.800 114.600 112.100 ;
        RECT 115.800 110.800 116.200 112.100 ;
        RECT 119.000 110.800 119.400 114.100 ;
        RECT 119.800 110.800 120.200 112.100 ;
        RECT 121.400 110.800 121.800 112.100 ;
        RECT 122.200 110.800 122.600 114.100 ;
        RECT 127.000 110.800 127.400 113.100 ;
        RECT 128.600 110.800 129.000 113.100 ;
        RECT 130.200 110.800 130.600 113.100 ;
        RECT 131.800 110.800 132.200 113.000 ;
        RECT 134.600 110.800 135.000 112.100 ;
        RECT 136.200 110.800 136.700 112.100 ;
        RECT 139.000 110.800 139.400 113.100 ;
        RECT 142.200 110.800 142.600 113.100 ;
        RECT 146.200 110.800 146.600 112.700 ;
        RECT 147.800 110.800 148.200 112.100 ;
        RECT 150.200 110.800 150.600 112.700 ;
        RECT 155.000 110.800 155.400 113.100 ;
        RECT 157.400 110.800 157.800 112.700 ;
        RECT 159.000 110.800 159.400 113.100 ;
        RECT 161.400 110.800 161.800 113.100 ;
        RECT 164.100 110.800 164.500 113.100 ;
        RECT 166.200 110.800 166.600 112.100 ;
        RECT 167.300 110.800 167.700 113.100 ;
        RECT 169.400 110.800 169.800 112.100 ;
        RECT 170.200 110.800 170.600 113.100 ;
        RECT 171.800 110.800 172.200 113.100 ;
        RECT 175.000 110.800 175.400 112.700 ;
        RECT 176.600 110.800 177.000 112.100 ;
        RECT 178.700 110.800 179.100 113.100 ;
        RECT 180.600 110.800 181.000 112.700 ;
        RECT 184.600 110.800 185.000 113.100 ;
        RECT 185.700 110.800 186.100 113.100 ;
        RECT 187.800 110.800 188.200 112.100 ;
        RECT 190.200 110.800 190.600 112.700 ;
        RECT 194.200 110.800 194.600 113.100 ;
        RECT 196.900 110.800 197.400 112.100 ;
        RECT 198.600 110.800 199.000 112.100 ;
        RECT 201.400 110.800 201.800 113.000 ;
        RECT 203.600 110.800 204.000 113.500 ;
        RECT 206.200 110.800 206.600 113.300 ;
        RECT 207.800 110.800 208.200 113.100 ;
        RECT 211.000 110.800 211.400 113.000 ;
        RECT 213.800 110.800 214.200 112.100 ;
        RECT 215.400 110.800 215.900 112.100 ;
        RECT 218.200 110.800 218.600 113.100 ;
        RECT 220.600 110.800 221.000 113.100 ;
        RECT 223.300 110.800 223.800 112.100 ;
        RECT 225.000 110.800 225.400 112.100 ;
        RECT 227.800 110.800 228.200 113.000 ;
        RECT 0.200 110.200 231.000 110.800 ;
        RECT 2.200 107.900 2.600 110.200 ;
        RECT 3.000 108.900 3.400 110.200 ;
        RECT 4.600 107.900 5.000 110.200 ;
        RECT 8.600 108.300 9.000 110.200 ;
        RECT 11.000 107.900 11.400 110.200 ;
        RECT 13.700 108.900 14.200 110.200 ;
        RECT 15.400 108.900 15.800 110.200 ;
        RECT 18.200 108.000 18.600 110.200 ;
        RECT 20.600 108.300 21.000 110.200 ;
        RECT 24.600 107.900 25.000 110.200 ;
        RECT 26.200 108.300 26.600 110.200 ;
        RECT 28.600 107.900 29.000 110.200 ;
        RECT 30.200 107.900 30.600 110.200 ;
        RECT 31.800 108.900 32.200 110.200 ;
        RECT 35.800 107.900 36.200 110.200 ;
        RECT 38.500 108.900 39.000 110.200 ;
        RECT 40.200 108.900 40.600 110.200 ;
        RECT 43.000 108.000 43.400 110.200 ;
        RECT 45.400 107.900 45.800 110.200 ;
        RECT 47.000 107.900 47.400 110.200 ;
        RECT 48.600 107.900 49.000 110.200 ;
        RECT 51.300 108.900 51.800 110.200 ;
        RECT 53.000 108.900 53.400 110.200 ;
        RECT 55.800 108.000 56.200 110.200 ;
        RECT 57.400 108.900 57.800 110.200 ;
        RECT 59.000 107.900 59.400 110.200 ;
        RECT 63.000 108.300 63.400 110.200 ;
        RECT 65.400 107.900 65.800 110.200 ;
        RECT 68.100 108.900 68.600 110.200 ;
        RECT 69.800 108.900 70.200 110.200 ;
        RECT 72.600 108.000 73.000 110.200 ;
        RECT 75.000 107.900 75.400 110.200 ;
        RECT 76.600 107.900 77.000 110.200 ;
        RECT 78.200 108.300 78.600 110.200 ;
        RECT 81.400 108.300 81.800 110.200 ;
        RECT 85.400 108.300 85.800 110.200 ;
        RECT 89.400 107.900 89.800 110.200 ;
        RECT 92.100 108.900 92.600 110.200 ;
        RECT 93.800 108.900 94.200 110.200 ;
        RECT 96.600 108.000 97.000 110.200 ;
        RECT 99.000 108.300 99.400 110.200 ;
        RECT 103.000 107.900 103.400 110.200 ;
        RECT 104.600 107.900 105.000 110.200 ;
        RECT 107.300 108.900 107.800 110.200 ;
        RECT 109.000 108.900 109.400 110.200 ;
        RECT 111.800 108.000 112.200 110.200 ;
        RECT 113.400 107.900 113.800 110.200 ;
        RECT 115.000 107.900 115.400 110.200 ;
        RECT 115.800 108.900 116.200 110.200 ;
        RECT 117.400 108.900 117.800 110.200 ;
        RECT 118.200 107.900 118.600 110.200 ;
        RECT 119.800 107.900 120.200 110.200 ;
        RECT 122.200 107.900 122.600 110.200 ;
        RECT 123.800 107.900 124.200 110.200 ;
        RECT 126.200 108.300 126.600 110.200 ;
        RECT 128.600 107.900 129.000 110.200 ;
        RECT 131.300 108.900 131.800 110.200 ;
        RECT 133.000 108.900 133.400 110.200 ;
        RECT 135.800 108.000 136.200 110.200 ;
        RECT 138.200 108.300 138.600 110.200 ;
        RECT 143.800 107.900 144.200 110.200 ;
        RECT 144.600 108.900 145.000 110.200 ;
        RECT 147.800 108.300 148.200 110.200 ;
        RECT 150.200 108.300 150.600 110.200 ;
        RECT 152.600 107.900 153.000 110.200 ;
        RECT 155.000 108.900 155.400 110.200 ;
        RECT 156.600 108.900 157.000 110.200 ;
        RECT 159.000 108.300 159.400 110.200 ;
        RECT 160.900 107.900 161.300 110.200 ;
        RECT 163.000 108.900 163.400 110.200 ;
        RECT 165.400 108.300 165.800 110.200 ;
        RECT 167.800 108.900 168.200 110.200 ;
        RECT 169.400 108.000 169.800 110.200 ;
        RECT 172.200 108.900 172.600 110.200 ;
        RECT 173.800 108.900 174.300 110.200 ;
        RECT 176.600 107.900 177.000 110.200 ;
        RECT 178.200 107.900 178.600 110.200 ;
        RECT 182.200 108.300 182.600 110.200 ;
        RECT 183.800 107.900 184.200 110.200 ;
        RECT 187.000 108.300 187.400 110.200 ;
        RECT 191.000 107.900 191.400 110.200 ;
        RECT 194.200 108.000 194.600 110.200 ;
        RECT 197.000 108.900 197.400 110.200 ;
        RECT 198.600 108.900 199.100 110.200 ;
        RECT 201.400 107.900 201.800 110.200 ;
        RECT 203.000 107.900 203.400 110.200 ;
        RECT 204.600 107.900 205.000 110.200 ;
        RECT 206.200 107.900 206.600 110.200 ;
        RECT 207.800 108.300 208.200 110.200 ;
        RECT 211.000 108.000 211.400 110.200 ;
        RECT 213.800 108.900 214.200 110.200 ;
        RECT 215.400 108.900 215.900 110.200 ;
        RECT 218.200 107.900 218.600 110.200 ;
        RECT 220.600 107.900 221.000 110.200 ;
        RECT 223.300 108.900 223.800 110.200 ;
        RECT 225.000 108.900 225.400 110.200 ;
        RECT 227.800 108.000 228.200 110.200 ;
        RECT 1.400 90.800 1.800 93.000 ;
        RECT 4.200 90.800 4.600 92.100 ;
        RECT 5.800 90.800 6.300 92.100 ;
        RECT 8.600 90.800 9.000 93.100 ;
        RECT 10.200 90.800 10.600 93.100 ;
        RECT 14.200 90.800 14.600 92.700 ;
        RECT 16.600 90.800 17.000 92.700 ;
        RECT 20.600 90.800 21.000 93.100 ;
        RECT 22.200 90.800 22.600 93.100 ;
        RECT 24.900 90.800 25.400 92.100 ;
        RECT 26.600 90.800 27.000 92.100 ;
        RECT 29.400 90.800 29.800 93.000 ;
        RECT 31.000 90.800 31.400 92.100 ;
        RECT 32.600 90.800 33.000 93.100 ;
        RECT 35.000 90.800 35.400 92.100 ;
        RECT 39.000 90.800 39.400 92.700 ;
        RECT 41.400 90.800 41.800 92.100 ;
        RECT 43.800 90.800 44.200 92.700 ;
        RECT 47.800 90.800 48.200 92.700 ;
        RECT 50.200 90.800 50.600 93.100 ;
        RECT 54.200 90.800 54.600 93.100 ;
        RECT 55.800 90.800 56.200 92.700 ;
        RECT 59.000 90.800 59.400 93.100 ;
        RECT 61.700 90.800 62.200 92.100 ;
        RECT 63.400 90.800 63.800 92.100 ;
        RECT 66.200 90.800 66.600 93.000 ;
        RECT 67.800 90.800 68.200 93.100 ;
        RECT 71.800 90.800 72.200 92.700 ;
        RECT 73.400 90.800 73.800 93.100 ;
        RECT 75.000 90.800 75.400 93.100 ;
        RECT 77.400 90.800 77.800 92.700 ;
        RECT 80.600 90.800 81.000 93.000 ;
        RECT 83.400 90.800 83.800 92.100 ;
        RECT 85.000 90.800 85.500 92.100 ;
        RECT 87.800 90.800 88.200 93.100 ;
        RECT 91.000 90.800 91.400 93.100 ;
        RECT 95.800 90.800 96.200 94.100 ;
        RECT 98.200 90.800 98.600 93.100 ;
        RECT 99.000 90.800 99.400 93.100 ;
        RECT 103.000 90.800 103.400 92.700 ;
        RECT 106.200 90.800 106.600 93.100 ;
        RECT 108.600 90.800 109.000 93.100 ;
        RECT 110.000 90.800 110.400 93.500 ;
        RECT 112.600 90.800 113.000 93.300 ;
        RECT 115.800 90.800 116.200 93.100 ;
        RECT 116.600 90.800 117.000 93.100 ;
        RECT 118.200 90.800 118.600 93.100 ;
        RECT 119.800 90.800 120.200 93.100 ;
        RECT 121.400 90.800 121.800 93.100 ;
        RECT 124.600 90.800 125.000 93.100 ;
        RECT 125.400 90.800 125.800 93.100 ;
        RECT 128.400 90.800 128.800 93.100 ;
        RECT 130.200 90.800 130.600 92.100 ;
        RECT 132.600 90.800 133.000 93.100 ;
        RECT 135.000 90.800 135.400 92.700 ;
        RECT 139.000 90.800 139.400 93.100 ;
        RECT 141.700 90.800 142.200 92.100 ;
        RECT 143.400 90.800 143.800 92.100 ;
        RECT 146.200 90.800 146.600 93.000 ;
        RECT 149.400 90.800 149.800 92.700 ;
        RECT 152.600 90.800 153.000 92.700 ;
        RECT 154.200 90.800 154.600 93.100 ;
        RECT 155.800 90.800 156.200 93.100 ;
        RECT 158.200 90.800 158.600 93.100 ;
        RECT 159.800 90.800 160.200 93.100 ;
        RECT 161.400 90.800 161.800 93.100 ;
        RECT 164.100 90.800 164.600 92.100 ;
        RECT 165.800 90.800 166.200 92.100 ;
        RECT 168.600 90.800 169.000 93.000 ;
        RECT 171.000 90.800 171.400 93.100 ;
        RECT 173.700 90.800 174.200 92.100 ;
        RECT 175.400 90.800 175.800 92.100 ;
        RECT 178.200 90.800 178.600 93.000 ;
        RECT 180.600 90.800 181.000 92.700 ;
        RECT 184.600 90.800 185.000 93.100 ;
        RECT 185.400 90.800 185.800 93.100 ;
        RECT 187.000 90.800 187.400 93.100 ;
        RECT 188.600 90.800 189.000 93.100 ;
        RECT 192.900 90.800 193.300 93.100 ;
        RECT 195.000 90.800 195.400 92.100 ;
        RECT 197.400 90.800 197.800 92.700 ;
        RECT 199.300 90.800 199.700 93.100 ;
        RECT 201.400 90.800 201.800 92.100 ;
        RECT 203.800 90.800 204.200 92.700 ;
        RECT 206.200 90.800 206.600 93.100 ;
        RECT 208.900 90.800 209.400 92.100 ;
        RECT 210.600 90.800 211.000 92.100 ;
        RECT 213.400 90.800 213.800 93.000 ;
        RECT 215.800 90.800 216.200 93.100 ;
        RECT 218.500 90.800 219.000 92.100 ;
        RECT 220.200 90.800 220.600 92.100 ;
        RECT 223.000 90.800 223.400 93.000 ;
        RECT 225.400 90.800 225.800 93.100 ;
        RECT 227.800 90.800 228.200 93.100 ;
        RECT 0.200 90.200 231.000 90.800 ;
        RECT 1.400 87.900 1.800 90.200 ;
        RECT 4.100 88.900 4.600 90.200 ;
        RECT 5.800 88.900 6.200 90.200 ;
        RECT 8.600 88.000 9.000 90.200 ;
        RECT 11.800 88.300 12.200 90.200 ;
        RECT 15.000 88.300 15.400 90.200 ;
        RECT 17.400 88.300 17.800 90.200 ;
        RECT 21.400 88.300 21.800 90.200 ;
        RECT 23.800 88.300 24.200 90.200 ;
        RECT 27.000 88.300 27.400 90.200 ;
        RECT 30.200 87.900 30.600 90.200 ;
        RECT 32.900 88.900 33.400 90.200 ;
        RECT 34.600 88.900 35.000 90.200 ;
        RECT 37.400 88.000 37.800 90.200 ;
        RECT 40.600 87.900 41.000 90.200 ;
        RECT 43.800 87.900 44.200 90.200 ;
        RECT 46.500 88.900 47.000 90.200 ;
        RECT 48.200 88.900 48.600 90.200 ;
        RECT 51.000 88.000 51.400 90.200 ;
        RECT 53.400 88.300 53.800 90.200 ;
        RECT 57.400 87.900 57.800 90.200 ;
        RECT 58.200 88.900 58.600 90.200 ;
        RECT 60.600 88.300 61.000 90.200 ;
        RECT 64.600 88.900 65.000 90.200 ;
        RECT 66.200 88.300 66.600 90.200 ;
        RECT 68.600 87.900 69.000 90.200 ;
        RECT 70.200 87.900 70.600 90.200 ;
        RECT 71.800 87.900 72.200 90.200 ;
        RECT 73.400 87.900 73.800 90.200 ;
        RECT 75.000 87.900 75.400 90.200 ;
        RECT 75.800 86.900 76.200 90.200 ;
        RECT 79.800 88.000 80.200 90.200 ;
        RECT 82.600 88.900 83.000 90.200 ;
        RECT 84.200 88.900 84.700 90.200 ;
        RECT 87.000 87.900 87.400 90.200 ;
        RECT 91.000 88.300 91.400 90.200 ;
        RECT 93.400 87.900 93.800 90.200 ;
        RECT 96.600 88.300 97.000 90.200 ;
        RECT 99.800 87.900 100.200 90.200 ;
        RECT 102.500 88.900 103.000 90.200 ;
        RECT 104.200 88.900 104.600 90.200 ;
        RECT 107.000 88.000 107.400 90.200 ;
        RECT 109.400 88.300 109.800 90.200 ;
        RECT 112.100 87.900 112.500 90.200 ;
        RECT 114.200 88.900 114.600 90.200 ;
        RECT 115.800 88.300 116.200 90.200 ;
        RECT 119.000 88.300 119.400 90.200 ;
        RECT 122.200 87.900 122.600 90.200 ;
        RECT 124.900 88.900 125.400 90.200 ;
        RECT 126.600 88.900 127.000 90.200 ;
        RECT 129.400 88.000 129.800 90.200 ;
        RECT 131.800 88.000 132.200 90.200 ;
        RECT 134.600 88.900 135.000 90.200 ;
        RECT 136.200 88.900 136.700 90.200 ;
        RECT 139.000 87.900 139.400 90.200 ;
        RECT 142.200 87.900 142.600 90.200 ;
        RECT 146.200 88.300 146.600 90.200 ;
        RECT 149.400 87.900 149.800 90.200 ;
        RECT 151.800 87.900 152.200 90.200 ;
        RECT 152.900 87.900 153.300 90.200 ;
        RECT 155.000 88.900 155.400 90.200 ;
        RECT 156.100 87.900 156.500 90.200 ;
        RECT 158.200 88.900 158.600 90.200 ;
        RECT 159.300 87.900 159.700 90.200 ;
        RECT 161.400 88.900 161.800 90.200 ;
        RECT 162.500 87.900 162.900 90.200 ;
        RECT 164.600 88.900 165.000 90.200 ;
        RECT 167.000 88.300 167.400 90.200 ;
        RECT 170.200 88.300 170.600 90.200 ;
        RECT 172.600 87.900 173.000 90.200 ;
        RECT 175.800 88.300 176.200 90.200 ;
        RECT 177.400 88.900 177.800 90.200 ;
        RECT 179.500 87.900 179.900 90.200 ;
        RECT 181.400 88.300 181.800 90.200 ;
        RECT 185.400 87.900 185.800 90.200 ;
        RECT 186.800 87.500 187.200 90.200 ;
        RECT 189.400 87.700 189.800 90.200 ;
        RECT 193.400 88.300 193.800 90.200 ;
        RECT 197.400 87.900 197.800 90.200 ;
        RECT 199.000 88.000 199.400 90.200 ;
        RECT 201.800 88.900 202.200 90.200 ;
        RECT 203.400 88.900 203.900 90.200 ;
        RECT 206.200 87.900 206.600 90.200 ;
        RECT 208.600 87.700 209.000 90.200 ;
        RECT 211.200 87.500 211.600 90.200 ;
        RECT 213.400 88.000 213.800 90.200 ;
        RECT 216.200 88.900 216.600 90.200 ;
        RECT 217.800 88.900 218.300 90.200 ;
        RECT 220.600 87.900 221.000 90.200 ;
        RECT 222.200 87.900 222.600 90.200 ;
        RECT 226.200 88.300 226.600 90.200 ;
        RECT 227.800 87.900 228.200 90.200 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 4.100 70.800 4.600 72.100 ;
        RECT 5.800 70.800 6.200 72.100 ;
        RECT 8.600 70.800 9.000 73.000 ;
        RECT 11.000 70.800 11.400 72.700 ;
        RECT 15.000 70.800 15.400 73.100 ;
        RECT 16.600 70.800 17.000 72.700 ;
        RECT 20.600 70.800 21.000 73.100 ;
        RECT 22.200 70.800 22.600 73.100 ;
        RECT 24.900 70.800 25.400 72.100 ;
        RECT 26.600 70.800 27.000 72.100 ;
        RECT 29.400 70.800 29.800 73.000 ;
        RECT 33.400 70.800 33.800 72.700 ;
        RECT 35.800 70.800 36.200 72.100 ;
        RECT 36.600 70.800 37.000 72.100 ;
        RECT 42.200 70.800 42.600 72.700 ;
        RECT 44.600 70.800 45.000 72.700 ;
        RECT 47.800 70.800 48.200 72.700 ;
        RECT 51.000 70.800 51.400 73.100 ;
        RECT 52.600 70.800 53.000 73.100 ;
        RECT 55.000 70.800 55.400 72.700 ;
        RECT 58.200 70.800 58.600 73.100 ;
        RECT 59.800 70.800 60.200 72.700 ;
        RECT 63.800 70.800 64.200 72.700 ;
        RECT 66.200 70.800 66.600 72.700 ;
        RECT 70.200 70.800 70.600 73.100 ;
        RECT 71.800 70.800 72.200 73.000 ;
        RECT 74.600 70.800 75.000 72.100 ;
        RECT 76.200 70.800 76.700 72.100 ;
        RECT 79.000 70.800 79.400 73.100 ;
        RECT 80.600 70.800 81.000 72.100 ;
        RECT 82.200 70.800 82.600 72.100 ;
        RECT 83.800 70.800 84.200 72.700 ;
        RECT 87.800 70.800 88.200 73.100 ;
        RECT 91.000 70.800 91.400 73.000 ;
        RECT 93.800 70.800 94.200 72.100 ;
        RECT 95.400 70.800 95.900 72.100 ;
        RECT 98.200 70.800 98.600 73.100 ;
        RECT 100.600 70.800 101.000 73.300 ;
        RECT 103.200 70.800 103.600 73.500 ;
        RECT 104.600 70.800 105.000 74.100 ;
        RECT 109.400 70.800 109.800 73.100 ;
        RECT 111.000 70.800 111.400 72.700 ;
        RECT 113.400 70.800 113.800 74.100 ;
        RECT 116.600 70.800 117.000 73.100 ;
        RECT 118.200 70.800 118.600 73.100 ;
        RECT 119.800 70.800 120.200 73.100 ;
        RECT 122.200 70.800 122.600 73.100 ;
        RECT 123.800 70.800 124.200 73.100 ;
        RECT 126.200 70.800 126.600 73.100 ;
        RECT 128.900 70.800 129.400 72.100 ;
        RECT 130.600 70.800 131.000 72.100 ;
        RECT 133.400 70.800 133.800 73.000 ;
        RECT 135.800 70.800 136.200 72.700 ;
        RECT 139.800 70.800 140.200 73.100 ;
        RECT 143.000 70.800 143.400 72.700 ;
        RECT 147.000 70.800 147.400 73.100 ;
        RECT 148.600 70.800 149.000 73.100 ;
        RECT 151.300 70.800 151.800 72.100 ;
        RECT 153.000 70.800 153.400 72.100 ;
        RECT 155.800 70.800 156.200 73.000 ;
        RECT 157.400 70.800 157.800 73.100 ;
        RECT 159.000 70.800 159.400 73.100 ;
        RECT 160.600 70.800 161.000 73.100 ;
        RECT 162.200 70.800 162.600 73.100 ;
        RECT 164.900 70.800 165.400 72.100 ;
        RECT 166.600 70.800 167.000 72.100 ;
        RECT 169.400 70.800 169.800 73.000 ;
        RECT 171.800 70.800 172.200 73.100 ;
        RECT 175.000 70.800 175.400 72.700 ;
        RECT 177.400 70.800 177.800 73.100 ;
        RECT 179.000 70.800 179.400 73.100 ;
        RECT 182.200 70.800 182.600 74.100 ;
        RECT 183.000 70.800 183.400 73.100 ;
        RECT 186.200 70.800 186.600 73.300 ;
        RECT 188.800 70.800 189.200 73.500 ;
        RECT 193.400 70.800 193.800 72.700 ;
        RECT 195.800 70.800 196.200 72.100 ;
        RECT 197.200 70.800 197.600 73.500 ;
        RECT 199.800 70.800 200.200 73.300 ;
        RECT 202.000 70.800 202.400 73.500 ;
        RECT 204.600 70.800 205.000 73.300 ;
        RECT 207.000 70.800 207.400 73.000 ;
        RECT 209.800 70.800 210.200 72.100 ;
        RECT 211.400 70.800 211.900 72.100 ;
        RECT 214.200 70.800 214.600 73.100 ;
        RECT 215.800 70.800 216.200 73.100 ;
        RECT 219.800 70.800 220.200 72.700 ;
        RECT 221.400 70.800 221.800 73.100 ;
        RECT 223.000 70.800 223.400 73.100 ;
        RECT 224.600 70.800 225.000 73.100 ;
        RECT 226.200 70.800 226.600 73.100 ;
        RECT 227.800 70.800 228.200 73.100 ;
        RECT 229.400 70.800 229.800 73.100 ;
        RECT 0.200 70.200 231.000 70.800 ;
        RECT 0.600 67.900 1.000 70.200 ;
        RECT 2.200 67.900 2.600 70.200 ;
        RECT 3.800 67.900 4.200 70.200 ;
        RECT 5.400 67.900 5.800 70.200 ;
        RECT 8.100 68.900 8.600 70.200 ;
        RECT 9.800 68.900 10.200 70.200 ;
        RECT 12.600 68.000 13.000 70.200 ;
        RECT 15.800 68.300 16.200 70.200 ;
        RECT 17.400 68.900 17.800 70.200 ;
        RECT 19.800 68.300 20.200 70.200 ;
        RECT 23.000 67.900 23.400 70.200 ;
        RECT 25.700 68.900 26.200 70.200 ;
        RECT 27.400 68.900 27.800 70.200 ;
        RECT 30.200 68.000 30.600 70.200 ;
        RECT 32.600 68.300 33.000 70.200 ;
        RECT 35.000 67.900 35.400 70.200 ;
        RECT 36.600 67.900 37.000 70.200 ;
        RECT 41.400 68.300 41.800 70.200 ;
        RECT 43.800 67.900 44.200 70.200 ;
        RECT 45.400 67.900 45.800 70.200 ;
        RECT 46.200 67.900 46.600 70.200 ;
        RECT 48.600 67.900 49.000 70.200 ;
        RECT 51.800 67.900 52.200 70.200 ;
        RECT 54.500 68.900 55.000 70.200 ;
        RECT 56.200 68.900 56.600 70.200 ;
        RECT 59.000 68.000 59.400 70.200 ;
        RECT 62.200 67.900 62.600 70.200 ;
        RECT 63.000 67.900 63.400 70.200 ;
        RECT 65.400 67.900 65.800 70.200 ;
        RECT 68.600 67.700 69.000 70.200 ;
        RECT 71.200 67.500 71.600 70.200 ;
        RECT 73.400 68.300 73.800 70.200 ;
        RECT 77.400 67.900 77.800 70.200 ;
        RECT 79.000 67.900 79.400 70.200 ;
        RECT 81.700 68.900 82.200 70.200 ;
        RECT 83.400 68.900 83.800 70.200 ;
        RECT 86.200 68.000 86.600 70.200 ;
        RECT 90.000 67.500 90.400 70.200 ;
        RECT 92.600 67.700 93.000 70.200 ;
        RECT 95.800 67.900 96.200 70.200 ;
        RECT 98.200 68.300 98.600 70.200 ;
        RECT 100.100 67.900 100.500 70.200 ;
        RECT 102.200 68.900 102.600 70.200 ;
        RECT 104.600 68.300 105.000 70.200 ;
        RECT 107.000 68.300 107.400 70.200 ;
        RECT 111.000 67.900 111.400 70.200 ;
        RECT 111.800 67.900 112.200 70.200 ;
        RECT 114.200 67.900 114.600 70.200 ;
        RECT 118.200 68.300 118.600 70.200 ;
        RECT 120.600 68.300 121.000 70.200 ;
        RECT 123.300 67.900 123.700 70.200 ;
        RECT 125.400 68.900 125.800 70.200 ;
        RECT 127.000 68.300 127.400 70.200 ;
        RECT 130.200 68.000 130.600 70.200 ;
        RECT 133.000 68.900 133.400 70.200 ;
        RECT 134.600 68.900 135.100 70.200 ;
        RECT 137.400 67.900 137.800 70.200 ;
        RECT 140.900 67.900 141.300 70.200 ;
        RECT 143.000 68.900 143.400 70.200 ;
        RECT 143.800 66.900 144.200 70.200 ;
        RECT 147.800 68.300 148.200 70.200 ;
        RECT 151.000 67.700 151.400 70.200 ;
        RECT 153.600 67.500 154.000 70.200 ;
        RECT 155.300 67.900 155.700 70.200 ;
        RECT 157.400 68.900 157.800 70.200 ;
        RECT 158.500 67.900 158.900 70.200 ;
        RECT 160.600 68.900 161.000 70.200 ;
        RECT 161.700 67.900 162.100 70.200 ;
        RECT 163.800 68.900 164.200 70.200 ;
        RECT 166.200 68.300 166.600 70.200 ;
        RECT 168.100 67.900 168.500 70.200 ;
        RECT 170.200 68.900 170.600 70.200 ;
        RECT 172.600 68.300 173.000 70.200 ;
        RECT 175.000 67.900 175.400 70.200 ;
        RECT 177.700 68.900 178.200 70.200 ;
        RECT 179.400 68.900 179.800 70.200 ;
        RECT 182.200 68.000 182.600 70.200 ;
        RECT 185.400 67.900 185.800 70.200 ;
        RECT 186.200 67.900 186.600 70.200 ;
        RECT 189.400 67.900 189.800 70.200 ;
        RECT 191.000 67.900 191.400 70.200 ;
        RECT 194.200 68.000 194.600 70.200 ;
        RECT 197.000 68.900 197.400 70.200 ;
        RECT 198.600 68.900 199.100 70.200 ;
        RECT 201.400 67.900 201.800 70.200 ;
        RECT 203.800 68.300 204.200 70.200 ;
        RECT 206.200 67.900 206.600 70.200 ;
        RECT 210.200 68.300 210.600 70.200 ;
        RECT 212.600 68.000 213.000 70.200 ;
        RECT 215.400 68.900 215.800 70.200 ;
        RECT 217.000 68.900 217.500 70.200 ;
        RECT 219.800 67.900 220.200 70.200 ;
        RECT 222.200 67.900 222.600 70.200 ;
        RECT 224.900 68.900 225.400 70.200 ;
        RECT 226.600 68.900 227.000 70.200 ;
        RECT 229.400 68.000 229.800 70.200 ;
        RECT 1.400 50.800 1.800 53.100 ;
        RECT 3.000 50.800 3.400 53.100 ;
        RECT 4.600 50.800 5.000 53.100 ;
        RECT 7.300 50.800 7.800 52.100 ;
        RECT 9.000 50.800 9.400 52.100 ;
        RECT 11.800 50.800 12.200 53.000 ;
        RECT 13.400 50.800 13.800 53.100 ;
        RECT 16.600 50.800 17.000 52.700 ;
        RECT 20.600 50.800 21.000 53.100 ;
        RECT 21.400 50.800 21.800 53.100 ;
        RECT 23.000 50.800 23.400 53.100 ;
        RECT 24.600 50.800 25.000 53.100 ;
        RECT 26.200 50.800 26.600 53.100 ;
        RECT 27.800 50.800 28.200 53.100 ;
        RECT 28.600 50.800 29.000 53.100 ;
        RECT 31.800 50.800 32.200 52.700 ;
        RECT 36.600 50.800 37.000 53.100 ;
        RECT 39.300 50.800 39.800 52.100 ;
        RECT 41.000 50.800 41.400 52.100 ;
        RECT 43.800 50.800 44.200 53.000 ;
        RECT 46.200 50.800 46.600 52.700 ;
        RECT 50.200 50.800 50.600 53.100 ;
        RECT 51.000 50.800 51.400 52.100 ;
        RECT 53.400 50.800 53.800 52.700 ;
        RECT 56.600 50.800 57.000 52.700 ;
        RECT 59.800 50.800 60.200 52.700 ;
        RECT 63.000 50.800 63.400 53.100 ;
        RECT 65.700 50.800 66.200 52.100 ;
        RECT 67.400 50.800 67.800 52.100 ;
        RECT 70.200 50.800 70.600 53.000 ;
        RECT 72.600 50.800 73.000 53.100 ;
        RECT 74.200 50.800 74.600 53.100 ;
        RECT 75.000 50.800 75.400 53.100 ;
        RECT 78.200 50.800 78.600 53.300 ;
        RECT 80.800 50.800 81.200 53.500 ;
        RECT 82.800 50.800 83.200 53.500 ;
        RECT 85.400 50.800 85.800 53.300 ;
        RECT 89.400 50.800 89.800 53.300 ;
        RECT 92.000 50.800 92.400 53.500 ;
        RECT 94.200 50.800 94.600 53.100 ;
        RECT 96.900 50.800 97.400 52.100 ;
        RECT 98.600 50.800 99.000 52.100 ;
        RECT 101.400 50.800 101.800 53.000 ;
        RECT 104.600 50.800 105.000 53.100 ;
        RECT 107.000 50.800 107.400 53.100 ;
        RECT 107.800 50.800 108.200 52.100 ;
        RECT 111.000 50.800 111.400 52.700 ;
        RECT 113.400 50.800 113.800 53.100 ;
        RECT 115.000 50.800 115.400 53.100 ;
        RECT 116.600 50.800 117.000 53.300 ;
        RECT 119.200 50.800 119.600 53.500 ;
        RECT 123.000 50.800 123.400 54.100 ;
        RECT 125.400 50.800 125.800 53.100 ;
        RECT 127.000 50.800 127.400 53.100 ;
        RECT 128.600 50.800 129.000 53.100 ;
        RECT 129.400 50.800 129.800 54.100 ;
        RECT 132.600 50.800 133.000 53.100 ;
        RECT 135.800 50.800 136.200 53.300 ;
        RECT 138.400 50.800 138.800 53.500 ;
        RECT 142.200 50.800 142.600 52.100 ;
        RECT 143.800 50.800 144.200 52.900 ;
        RECT 145.400 50.800 145.800 52.100 ;
        RECT 147.800 50.800 148.200 52.700 ;
        RECT 151.000 50.800 151.400 53.100 ;
        RECT 152.600 50.800 153.000 53.100 ;
        RECT 155.300 50.800 155.800 52.100 ;
        RECT 157.000 50.800 157.400 52.100 ;
        RECT 159.800 50.800 160.200 53.000 ;
        RECT 161.400 50.800 161.800 53.100 ;
        RECT 165.400 50.800 165.800 52.700 ;
        RECT 167.800 50.800 168.200 53.300 ;
        RECT 170.400 50.800 170.800 53.500 ;
        RECT 172.600 50.800 173.000 53.100 ;
        RECT 175.300 50.800 175.800 52.100 ;
        RECT 177.000 50.800 177.400 52.100 ;
        RECT 179.800 50.800 180.200 53.000 ;
        RECT 181.400 50.800 181.800 53.100 ;
        RECT 183.000 50.800 183.400 53.100 ;
        RECT 185.400 50.800 185.800 53.300 ;
        RECT 188.000 50.800 188.400 53.500 ;
        RECT 189.400 50.800 189.800 53.100 ;
        RECT 195.000 50.800 195.400 52.700 ;
        RECT 197.400 50.800 197.800 53.100 ;
        RECT 199.000 50.800 199.400 53.100 ;
        RECT 200.600 50.800 201.000 52.100 ;
        RECT 202.200 50.800 202.600 53.300 ;
        RECT 204.800 50.800 205.200 53.500 ;
        RECT 207.000 50.800 207.400 53.300 ;
        RECT 209.600 50.800 210.000 53.500 ;
        RECT 211.000 50.800 211.400 53.100 ;
        RECT 212.600 50.800 213.000 53.100 ;
        RECT 215.000 50.800 215.400 52.700 ;
        RECT 218.200 50.800 218.600 53.000 ;
        RECT 221.000 50.800 221.400 52.100 ;
        RECT 222.600 50.800 223.100 52.100 ;
        RECT 225.400 50.800 225.800 53.100 ;
        RECT 227.800 50.800 228.200 53.100 ;
        RECT 229.400 50.800 229.800 53.100 ;
        RECT 0.200 50.200 231.000 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 4.100 48.900 4.600 50.200 ;
        RECT 5.800 48.900 6.200 50.200 ;
        RECT 8.600 48.000 9.000 50.200 ;
        RECT 10.200 47.900 10.600 50.200 ;
        RECT 14.200 48.300 14.600 50.200 ;
        RECT 15.800 47.900 16.200 50.200 ;
        RECT 19.000 47.900 19.400 50.200 ;
        RECT 21.700 48.900 22.200 50.200 ;
        RECT 23.400 48.900 23.800 50.200 ;
        RECT 26.200 48.000 26.600 50.200 ;
        RECT 27.800 47.900 28.200 50.200 ;
        RECT 31.800 48.300 32.200 50.200 ;
        RECT 33.400 47.900 33.800 50.200 ;
        RECT 38.200 47.900 38.600 50.200 ;
        RECT 40.900 48.900 41.400 50.200 ;
        RECT 42.600 48.900 43.000 50.200 ;
        RECT 45.400 48.000 45.800 50.200 ;
        RECT 47.800 48.300 48.200 50.200 ;
        RECT 51.800 47.900 52.200 50.200 ;
        RECT 53.400 48.000 53.800 50.200 ;
        RECT 56.200 48.900 56.600 50.200 ;
        RECT 57.800 48.900 58.300 50.200 ;
        RECT 60.600 47.900 61.000 50.200 ;
        RECT 63.800 48.300 64.200 50.200 ;
        RECT 66.200 47.900 66.600 50.200 ;
        RECT 68.900 48.900 69.400 50.200 ;
        RECT 70.600 48.900 71.000 50.200 ;
        RECT 73.400 48.000 73.800 50.200 ;
        RECT 76.600 48.300 77.000 50.200 ;
        RECT 79.000 48.300 79.400 50.200 ;
        RECT 83.000 47.900 83.400 50.200 ;
        RECT 84.600 48.000 85.000 50.200 ;
        RECT 87.400 48.900 87.800 50.200 ;
        RECT 89.000 48.900 89.500 50.200 ;
        RECT 91.800 47.900 92.200 50.200 ;
        RECT 95.800 48.300 96.200 50.200 ;
        RECT 99.800 47.900 100.200 50.200 ;
        RECT 101.400 47.900 101.800 50.200 ;
        RECT 104.100 48.900 104.600 50.200 ;
        RECT 105.800 48.900 106.200 50.200 ;
        RECT 108.600 48.000 109.000 50.200 ;
        RECT 110.200 48.900 110.600 50.200 ;
        RECT 112.400 47.500 112.800 50.200 ;
        RECT 115.000 47.700 115.400 50.200 ;
        RECT 117.400 47.700 117.800 50.200 ;
        RECT 120.000 47.500 120.400 50.200 ;
        RECT 123.000 47.900 123.400 50.200 ;
        RECT 125.400 47.900 125.800 50.200 ;
        RECT 127.000 48.000 127.400 50.200 ;
        RECT 129.800 48.900 130.200 50.200 ;
        RECT 131.400 48.900 131.900 50.200 ;
        RECT 134.200 47.900 134.600 50.200 ;
        RECT 135.800 47.900 136.200 50.200 ;
        RECT 139.800 48.300 140.200 50.200 ;
        RECT 143.000 47.900 143.400 50.200 ;
        RECT 144.600 47.900 145.000 50.200 ;
        RECT 147.000 47.900 147.400 50.200 ;
        RECT 148.600 48.300 149.000 50.200 ;
        RECT 151.800 47.900 152.200 50.200 ;
        RECT 154.500 48.900 155.000 50.200 ;
        RECT 156.200 48.900 156.600 50.200 ;
        RECT 159.000 48.000 159.400 50.200 ;
        RECT 161.400 47.900 161.800 50.200 ;
        RECT 163.800 48.300 164.200 50.200 ;
        RECT 167.800 47.900 168.200 50.200 ;
        RECT 169.400 48.000 169.800 50.200 ;
        RECT 172.200 48.900 172.600 50.200 ;
        RECT 173.800 48.900 174.300 50.200 ;
        RECT 176.600 47.900 177.000 50.200 ;
        RECT 178.200 47.900 178.600 50.200 ;
        RECT 179.800 47.900 180.200 50.200 ;
        RECT 182.200 47.700 182.600 50.200 ;
        RECT 184.800 47.500 185.200 50.200 ;
        RECT 187.000 48.000 187.400 50.200 ;
        RECT 189.800 48.900 190.200 50.200 ;
        RECT 191.400 48.900 191.900 50.200 ;
        RECT 194.200 47.900 194.600 50.200 ;
        RECT 198.200 47.900 198.600 50.200 ;
        RECT 199.800 47.900 200.200 50.200 ;
        RECT 200.600 47.900 201.000 50.200 ;
        RECT 202.200 47.900 202.600 50.200 ;
        RECT 204.400 47.500 204.800 50.200 ;
        RECT 207.000 47.700 207.400 50.200 ;
        RECT 208.600 47.900 209.000 50.200 ;
        RECT 212.600 48.300 213.000 50.200 ;
        RECT 214.200 47.900 214.600 50.200 ;
        RECT 217.400 48.300 217.800 50.200 ;
        RECT 220.600 48.000 221.000 50.200 ;
        RECT 223.400 48.900 223.800 50.200 ;
        RECT 225.000 48.900 225.500 50.200 ;
        RECT 227.800 47.900 228.200 50.200 ;
        RECT 2.200 30.800 2.600 33.100 ;
        RECT 3.000 30.800 3.400 32.100 ;
        RECT 5.400 30.800 5.800 32.700 ;
        RECT 9.400 30.800 9.800 33.100 ;
        RECT 10.200 30.800 10.600 32.100 ;
        RECT 14.200 30.800 14.600 32.700 ;
        RECT 16.600 30.800 17.000 33.100 ;
        RECT 19.300 30.800 19.800 32.100 ;
        RECT 21.000 30.800 21.400 32.100 ;
        RECT 23.800 30.800 24.200 33.000 ;
        RECT 25.400 30.800 25.800 32.100 ;
        RECT 29.400 30.800 29.800 32.700 ;
        RECT 31.800 30.800 32.200 32.100 ;
        RECT 33.400 30.800 33.800 33.100 ;
        RECT 36.100 30.800 36.600 32.100 ;
        RECT 37.800 30.800 38.200 32.100 ;
        RECT 40.600 30.800 41.000 33.000 ;
        RECT 44.600 30.800 45.000 32.100 ;
        RECT 45.400 30.800 45.800 33.100 ;
        RECT 49.400 30.800 49.800 32.700 ;
        RECT 51.800 30.800 52.200 33.100 ;
        RECT 53.400 30.800 53.800 33.100 ;
        RECT 54.800 30.800 55.200 33.500 ;
        RECT 57.400 30.800 57.800 33.300 ;
        RECT 59.000 30.800 59.400 33.100 ;
        RECT 62.200 30.800 62.600 32.700 ;
        RECT 66.200 30.800 66.600 33.100 ;
        RECT 67.600 30.800 68.000 33.500 ;
        RECT 70.200 30.800 70.600 33.300 ;
        RECT 72.600 30.800 73.000 32.700 ;
        RECT 75.000 30.800 75.400 33.100 ;
        RECT 78.200 30.800 78.600 32.700 ;
        RECT 82.200 30.800 82.600 33.100 ;
        RECT 83.600 30.800 84.000 33.500 ;
        RECT 86.200 30.800 86.600 33.300 ;
        RECT 90.200 30.800 90.600 33.000 ;
        RECT 93.000 30.800 93.400 32.100 ;
        RECT 94.600 30.800 95.100 32.100 ;
        RECT 97.400 30.800 97.800 33.100 ;
        RECT 99.000 30.800 99.400 33.100 ;
        RECT 103.000 30.800 103.400 32.700 ;
        RECT 106.200 30.800 106.600 33.100 ;
        RECT 107.800 30.800 108.200 33.300 ;
        RECT 110.400 30.800 110.800 33.500 ;
        RECT 111.800 30.800 112.200 33.100 ;
        RECT 115.800 30.800 116.200 32.700 ;
        RECT 118.200 30.800 118.600 32.700 ;
        RECT 121.200 30.800 121.600 33.500 ;
        RECT 123.800 30.800 124.200 33.300 ;
        RECT 126.200 30.800 126.600 33.300 ;
        RECT 128.800 30.800 129.200 33.500 ;
        RECT 131.000 30.800 131.400 33.300 ;
        RECT 133.600 30.800 134.000 33.500 ;
        RECT 135.000 30.800 135.400 33.100 ;
        RECT 139.000 30.800 139.400 32.700 ;
        RECT 143.000 30.800 143.400 33.000 ;
        RECT 145.800 30.800 146.200 32.100 ;
        RECT 147.400 30.800 147.900 32.100 ;
        RECT 150.200 30.800 150.600 33.100 ;
        RECT 152.600 30.800 153.000 32.700 ;
        RECT 156.400 30.800 156.800 33.500 ;
        RECT 159.000 30.800 159.400 33.300 ;
        RECT 160.600 30.800 161.000 33.100 ;
        RECT 163.000 30.800 163.400 33.100 ;
        RECT 166.200 30.800 166.600 32.700 ;
        RECT 169.400 30.800 169.800 32.100 ;
        RECT 170.200 30.800 170.600 33.100 ;
        RECT 171.800 30.800 172.200 33.100 ;
        RECT 173.400 30.800 173.800 33.100 ;
        RECT 177.400 30.800 177.800 32.700 ;
        RECT 179.800 30.800 180.200 33.300 ;
        RECT 182.400 30.800 182.800 33.500 ;
        RECT 184.600 30.800 185.000 32.100 ;
        RECT 186.200 30.800 186.600 33.000 ;
        RECT 189.000 30.800 189.400 32.100 ;
        RECT 190.600 30.800 191.100 32.100 ;
        RECT 193.400 30.800 193.800 33.100 ;
        RECT 197.400 30.800 197.800 32.700 ;
        RECT 200.600 30.800 201.000 32.700 ;
        RECT 204.600 30.800 205.000 33.100 ;
        RECT 206.200 30.800 206.600 33.000 ;
        RECT 209.000 30.800 209.400 32.100 ;
        RECT 210.600 30.800 211.100 32.100 ;
        RECT 213.400 30.800 213.800 33.100 ;
        RECT 215.800 30.800 216.200 32.700 ;
        RECT 219.800 30.800 220.200 33.100 ;
        RECT 221.400 30.800 221.800 33.000 ;
        RECT 224.200 30.800 224.600 32.100 ;
        RECT 225.800 30.800 226.300 32.100 ;
        RECT 228.600 30.800 229.000 33.100 ;
        RECT 0.200 30.200 231.000 30.800 ;
        RECT 2.200 28.300 2.600 30.200 ;
        RECT 4.600 28.000 5.000 30.200 ;
        RECT 7.400 28.900 7.800 30.200 ;
        RECT 9.000 28.900 9.500 30.200 ;
        RECT 11.800 27.900 12.200 30.200 ;
        RECT 14.200 28.000 14.600 30.200 ;
        RECT 17.000 28.900 17.400 30.200 ;
        RECT 18.600 28.900 19.100 30.200 ;
        RECT 21.400 27.900 21.800 30.200 ;
        RECT 23.000 28.900 23.400 30.200 ;
        RECT 24.600 27.900 25.000 30.200 ;
        RECT 28.600 28.300 29.000 30.200 ;
        RECT 30.200 27.900 30.600 30.200 ;
        RECT 31.800 27.900 32.200 30.200 ;
        RECT 33.400 27.900 33.800 30.200 ;
        RECT 35.000 27.900 35.400 30.200 ;
        RECT 36.600 27.900 37.000 30.200 ;
        RECT 39.800 28.000 40.200 30.200 ;
        RECT 42.600 28.900 43.000 30.200 ;
        RECT 44.200 28.900 44.700 30.200 ;
        RECT 47.000 27.900 47.400 30.200 ;
        RECT 49.400 28.300 49.800 30.200 ;
        RECT 51.800 27.900 52.200 30.200 ;
        RECT 54.200 27.900 54.600 30.200 ;
        RECT 58.200 28.300 58.600 30.200 ;
        RECT 60.600 27.900 61.000 30.200 ;
        RECT 63.300 28.900 63.800 30.200 ;
        RECT 65.000 28.900 65.400 30.200 ;
        RECT 67.800 28.000 68.200 30.200 ;
        RECT 70.200 28.000 70.600 30.200 ;
        RECT 73.000 28.900 73.400 30.200 ;
        RECT 74.600 28.900 75.100 30.200 ;
        RECT 77.400 27.900 77.800 30.200 ;
        RECT 79.000 27.900 79.400 30.200 ;
        RECT 83.000 28.300 83.400 30.200 ;
        RECT 87.000 28.000 87.400 30.200 ;
        RECT 89.800 28.900 90.200 30.200 ;
        RECT 91.400 28.900 91.900 30.200 ;
        RECT 94.200 27.900 94.600 30.200 ;
        RECT 95.800 27.900 96.200 30.200 ;
        RECT 98.200 27.900 98.600 30.200 ;
        RECT 102.200 27.900 102.600 30.200 ;
        RECT 103.800 28.300 104.200 30.200 ;
        RECT 107.000 27.900 107.400 30.200 ;
        RECT 109.700 28.900 110.200 30.200 ;
        RECT 111.400 28.900 111.800 30.200 ;
        RECT 114.200 28.000 114.600 30.200 ;
        RECT 116.600 28.000 117.000 30.200 ;
        RECT 119.400 28.900 119.800 30.200 ;
        RECT 121.000 28.900 121.500 30.200 ;
        RECT 123.800 27.900 124.200 30.200 ;
        RECT 127.000 27.900 127.400 30.200 ;
        RECT 127.800 27.900 128.200 30.200 ;
        RECT 129.400 27.900 129.800 30.200 ;
        RECT 131.000 27.900 131.400 30.200 ;
        RECT 132.600 27.900 133.000 30.200 ;
        RECT 134.200 27.900 134.600 30.200 ;
        RECT 135.000 27.900 135.400 30.200 ;
        RECT 136.600 27.900 137.000 30.200 ;
        RECT 138.200 27.900 138.600 30.200 ;
        RECT 139.800 27.900 140.200 30.200 ;
        RECT 141.400 27.900 141.800 30.200 ;
        RECT 143.800 27.900 144.200 30.200 ;
        RECT 147.800 28.300 148.200 30.200 ;
        RECT 150.200 28.000 150.600 30.200 ;
        RECT 153.000 28.900 153.400 30.200 ;
        RECT 154.600 28.900 155.100 30.200 ;
        RECT 157.400 27.900 157.800 30.200 ;
        RECT 159.800 28.300 160.200 30.200 ;
        RECT 163.000 28.300 163.400 30.200 ;
        RECT 167.000 27.900 167.400 30.200 ;
        RECT 168.600 28.000 169.000 30.200 ;
        RECT 171.400 28.900 171.800 30.200 ;
        RECT 173.000 28.900 173.500 30.200 ;
        RECT 175.800 27.900 176.200 30.200 ;
        RECT 178.200 28.000 178.600 30.200 ;
        RECT 181.000 28.900 181.400 30.200 ;
        RECT 182.600 28.900 183.100 30.200 ;
        RECT 185.400 27.900 185.800 30.200 ;
        RECT 189.400 27.900 189.800 30.200 ;
        RECT 192.100 28.900 192.600 30.200 ;
        RECT 193.800 28.900 194.200 30.200 ;
        RECT 196.600 28.000 197.000 30.200 ;
        RECT 199.800 27.900 200.200 30.200 ;
        RECT 201.400 27.900 201.800 30.200 ;
        RECT 203.000 27.900 203.400 30.200 ;
        RECT 204.600 28.300 205.000 30.200 ;
        RECT 208.600 27.900 209.000 30.200 ;
        RECT 210.200 28.000 210.600 30.200 ;
        RECT 213.000 28.900 213.400 30.200 ;
        RECT 214.600 28.900 215.100 30.200 ;
        RECT 217.400 27.900 217.800 30.200 ;
        RECT 220.600 27.900 221.000 30.200 ;
        RECT 222.200 28.000 222.600 30.200 ;
        RECT 225.000 28.900 225.400 30.200 ;
        RECT 226.600 28.900 227.100 30.200 ;
        RECT 229.400 27.900 229.800 30.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 4.100 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.200 12.100 ;
        RECT 8.600 10.800 9.000 13.000 ;
        RECT 11.000 10.800 11.400 12.700 ;
        RECT 14.200 10.800 14.600 13.100 ;
        RECT 16.900 10.800 17.400 12.100 ;
        RECT 18.600 10.800 19.000 12.100 ;
        RECT 21.400 10.800 21.800 13.000 ;
        RECT 23.000 10.800 23.400 12.100 ;
        RECT 25.400 10.800 25.800 13.100 ;
        RECT 28.100 10.800 28.600 12.100 ;
        RECT 29.800 10.800 30.200 12.100 ;
        RECT 32.600 10.800 33.000 13.000 ;
        RECT 35.800 10.800 36.200 12.700 ;
        RECT 39.600 10.800 40.000 13.500 ;
        RECT 42.200 10.800 42.600 13.300 ;
        RECT 44.600 10.800 45.000 13.100 ;
        RECT 46.200 10.800 46.600 13.100 ;
        RECT 47.800 10.800 48.200 13.100 ;
        RECT 50.500 10.800 51.000 12.100 ;
        RECT 52.200 10.800 52.600 12.100 ;
        RECT 55.000 10.800 55.400 13.000 ;
        RECT 57.400 10.800 57.800 12.700 ;
        RECT 61.400 10.800 61.800 13.100 ;
        RECT 62.200 10.800 62.600 12.100 ;
        RECT 64.600 10.800 65.000 12.700 ;
        RECT 68.600 10.800 69.000 13.100 ;
        RECT 70.200 10.800 70.600 13.100 ;
        RECT 72.900 10.800 73.400 12.100 ;
        RECT 74.600 10.800 75.000 12.100 ;
        RECT 77.400 10.800 77.800 13.000 ;
        RECT 79.000 10.800 79.400 13.100 ;
        RECT 80.600 10.800 81.000 13.100 ;
        RECT 83.000 10.800 83.400 12.700 ;
        RECT 87.000 10.800 87.400 13.100 ;
        RECT 90.200 10.800 90.600 13.100 ;
        RECT 92.900 10.800 93.400 12.100 ;
        RECT 94.600 10.800 95.000 12.100 ;
        RECT 97.400 10.800 97.800 13.000 ;
        RECT 99.000 10.800 99.400 12.100 ;
        RECT 101.400 10.800 101.800 13.100 ;
        RECT 104.100 10.800 104.600 12.100 ;
        RECT 105.800 10.800 106.200 12.100 ;
        RECT 108.600 10.800 109.000 13.000 ;
        RECT 111.000 10.800 111.400 12.700 ;
        RECT 115.000 10.800 115.400 13.100 ;
        RECT 116.600 10.800 117.000 13.300 ;
        RECT 119.200 10.800 119.600 13.500 ;
        RECT 121.400 10.800 121.800 12.700 ;
        RECT 125.400 10.800 125.800 13.100 ;
        RECT 127.000 10.800 127.400 13.100 ;
        RECT 128.600 10.800 129.000 13.100 ;
        RECT 129.400 10.800 129.800 13.100 ;
        RECT 132.400 10.800 132.800 13.500 ;
        RECT 135.000 10.800 135.400 13.300 ;
        RECT 136.600 10.800 137.000 13.100 ;
        RECT 142.200 10.800 142.600 12.700 ;
        RECT 144.400 10.800 144.800 13.500 ;
        RECT 147.000 10.800 147.400 13.300 ;
        RECT 149.400 10.800 149.800 13.100 ;
        RECT 152.100 10.800 152.600 12.100 ;
        RECT 153.800 10.800 154.200 12.100 ;
        RECT 156.600 10.800 157.000 13.000 ;
        RECT 159.000 10.800 159.400 13.100 ;
        RECT 161.700 10.800 162.200 12.100 ;
        RECT 163.400 10.800 163.800 12.100 ;
        RECT 166.200 10.800 166.600 13.000 ;
        RECT 167.800 10.800 168.200 13.100 ;
        RECT 171.800 10.800 172.200 12.700 ;
        RECT 174.200 10.800 174.600 13.100 ;
        RECT 176.900 10.800 177.400 12.100 ;
        RECT 178.600 10.800 179.000 12.100 ;
        RECT 181.400 10.800 181.800 13.000 ;
        RECT 183.000 10.800 183.400 13.100 ;
        RECT 184.600 10.800 185.000 13.100 ;
        RECT 185.400 10.800 185.800 12.100 ;
        RECT 187.000 10.800 187.400 12.100 ;
        RECT 187.800 10.800 188.200 13.100 ;
        RECT 189.400 10.800 189.800 13.100 ;
        RECT 192.600 10.800 193.000 13.000 ;
        RECT 195.400 10.800 195.800 12.100 ;
        RECT 197.000 10.800 197.500 12.100 ;
        RECT 199.800 10.800 200.200 13.100 ;
        RECT 202.200 10.800 202.600 13.300 ;
        RECT 204.800 10.800 205.200 13.500 ;
        RECT 206.200 10.800 206.600 13.100 ;
        RECT 210.200 10.800 210.600 12.700 ;
        RECT 212.600 10.800 213.000 12.700 ;
        RECT 216.600 10.800 217.000 13.100 ;
        RECT 217.400 10.800 217.800 13.100 ;
        RECT 219.000 10.800 219.400 13.100 ;
        RECT 220.600 10.800 221.000 13.100 ;
        RECT 222.200 10.800 222.600 13.100 ;
        RECT 223.800 10.800 224.200 13.100 ;
        RECT 224.600 10.800 225.000 13.100 ;
        RECT 228.600 10.800 229.000 12.700 ;
        RECT 0.200 10.200 231.000 10.800 ;
        RECT 2.200 8.300 2.600 10.200 ;
        RECT 5.400 7.900 5.800 10.200 ;
        RECT 6.200 7.900 6.600 10.200 ;
        RECT 7.800 7.900 8.200 10.200 ;
        RECT 9.400 7.900 9.800 10.200 ;
        RECT 11.000 7.900 11.400 10.200 ;
        RECT 12.600 7.900 13.000 10.200 ;
        RECT 15.000 7.900 15.400 10.200 ;
        RECT 15.800 7.900 16.200 10.200 ;
        RECT 17.400 7.900 17.800 10.200 ;
        RECT 19.000 7.900 19.400 10.200 ;
        RECT 20.600 7.900 21.000 10.200 ;
        RECT 22.200 7.900 22.600 10.200 ;
        RECT 23.000 7.900 23.400 10.200 ;
        RECT 24.600 7.900 25.000 10.200 ;
        RECT 26.200 7.900 26.600 10.200 ;
        RECT 27.800 7.900 28.200 10.200 ;
        RECT 29.400 7.900 29.800 10.200 ;
        RECT 31.000 7.900 31.400 10.200 ;
        RECT 33.700 8.900 34.200 10.200 ;
        RECT 35.400 8.900 35.800 10.200 ;
        RECT 38.200 8.000 38.600 10.200 ;
        RECT 43.000 7.900 43.400 10.200 ;
        RECT 43.800 7.900 44.200 10.200 ;
        RECT 47.800 8.300 48.200 10.200 ;
        RECT 50.200 8.000 50.600 10.200 ;
        RECT 53.000 8.900 53.400 10.200 ;
        RECT 54.600 8.900 55.100 10.200 ;
        RECT 57.400 7.900 57.800 10.200 ;
        RECT 59.800 7.900 60.200 10.200 ;
        RECT 62.500 8.900 63.000 10.200 ;
        RECT 64.200 8.900 64.600 10.200 ;
        RECT 67.000 8.000 67.400 10.200 ;
        RECT 69.400 7.900 69.800 10.200 ;
        RECT 72.100 8.900 72.600 10.200 ;
        RECT 73.800 8.900 74.200 10.200 ;
        RECT 76.600 8.000 77.000 10.200 ;
        RECT 78.200 8.900 78.600 10.200 ;
        RECT 80.300 7.900 80.700 10.200 ;
        RECT 81.700 7.900 82.100 10.200 ;
        RECT 83.800 8.900 84.200 10.200 ;
        RECT 84.600 8.900 85.000 10.200 ;
        RECT 86.200 8.900 86.600 10.200 ;
        RECT 87.000 8.900 87.400 10.200 ;
        RECT 88.600 8.900 89.000 10.200 ;
        RECT 91.800 8.300 92.200 10.200 ;
        RECT 95.800 7.900 96.200 10.200 ;
        RECT 97.400 7.900 97.800 10.200 ;
        RECT 100.100 8.900 100.600 10.200 ;
        RECT 101.800 8.900 102.200 10.200 ;
        RECT 104.600 8.000 105.000 10.200 ;
        RECT 106.200 7.900 106.600 10.200 ;
        RECT 107.800 7.900 108.200 10.200 ;
        RECT 109.400 7.900 109.800 10.200 ;
        RECT 111.000 7.900 111.400 10.200 ;
        RECT 113.700 8.900 114.200 10.200 ;
        RECT 115.400 8.900 115.800 10.200 ;
        RECT 118.200 8.000 118.600 10.200 ;
        RECT 120.600 7.900 121.000 10.200 ;
        RECT 123.300 8.900 123.800 10.200 ;
        RECT 125.000 8.900 125.400 10.200 ;
        RECT 127.800 8.000 128.200 10.200 ;
        RECT 131.000 8.300 131.400 10.200 ;
        RECT 133.400 8.000 133.800 10.200 ;
        RECT 136.200 8.900 136.600 10.200 ;
        RECT 137.800 8.900 138.300 10.200 ;
        RECT 140.600 7.900 141.000 10.200 ;
        RECT 144.600 8.000 145.000 10.200 ;
        RECT 147.400 8.900 147.800 10.200 ;
        RECT 149.000 8.900 149.500 10.200 ;
        RECT 151.800 7.900 152.200 10.200 ;
        RECT 153.400 7.900 153.800 10.200 ;
        RECT 157.400 8.300 157.800 10.200 ;
        RECT 159.800 8.300 160.200 10.200 ;
        RECT 163.800 7.900 164.200 10.200 ;
        RECT 165.400 8.000 165.800 10.200 ;
        RECT 168.200 8.900 168.600 10.200 ;
        RECT 169.800 8.900 170.300 10.200 ;
        RECT 172.600 7.900 173.000 10.200 ;
        RECT 174.200 7.900 174.600 10.200 ;
        RECT 176.600 8.900 177.000 10.200 ;
        RECT 178.200 8.900 178.600 10.200 ;
        RECT 180.600 7.900 181.000 10.200 ;
        RECT 181.700 7.900 182.100 10.200 ;
        RECT 183.800 8.900 184.200 10.200 ;
        RECT 184.600 8.900 185.000 10.200 ;
        RECT 186.200 8.900 186.600 10.200 ;
        RECT 187.300 7.900 187.700 10.200 ;
        RECT 189.400 8.900 189.800 10.200 ;
        RECT 190.200 8.900 190.600 10.200 ;
        RECT 191.800 8.900 192.200 10.200 ;
        RECT 194.500 7.900 194.900 10.200 ;
        RECT 196.600 8.900 197.000 10.200 ;
        RECT 197.400 8.900 197.800 10.200 ;
        RECT 199.000 8.900 199.400 10.200 ;
        RECT 200.600 7.900 201.000 10.200 ;
        RECT 203.300 8.900 203.800 10.200 ;
        RECT 205.000 8.900 205.400 10.200 ;
        RECT 207.800 8.000 208.200 10.200 ;
        RECT 210.200 8.000 210.600 10.200 ;
        RECT 213.000 8.900 213.400 10.200 ;
        RECT 214.600 8.900 215.100 10.200 ;
        RECT 217.400 7.900 217.800 10.200 ;
        RECT 220.600 7.900 221.000 10.200 ;
        RECT 222.200 8.000 222.600 10.200 ;
        RECT 225.000 8.900 225.400 10.200 ;
        RECT 226.600 8.900 227.100 10.200 ;
        RECT 229.400 7.900 229.800 10.200 ;
      LAYER via1 ;
        RECT 88.200 210.300 88.600 210.700 ;
        RECT 88.900 210.300 89.300 210.700 ;
        RECT 191.400 210.300 191.800 210.700 ;
        RECT 192.100 210.300 192.500 210.700 ;
        RECT 88.200 190.300 88.600 190.700 ;
        RECT 88.900 190.300 89.300 190.700 ;
        RECT 191.400 190.300 191.800 190.700 ;
        RECT 192.100 190.300 192.500 190.700 ;
        RECT 88.200 170.300 88.600 170.700 ;
        RECT 88.900 170.300 89.300 170.700 ;
        RECT 191.400 170.300 191.800 170.700 ;
        RECT 192.100 170.300 192.500 170.700 ;
        RECT 88.200 150.300 88.600 150.700 ;
        RECT 88.900 150.300 89.300 150.700 ;
        RECT 191.400 150.300 191.800 150.700 ;
        RECT 192.100 150.300 192.500 150.700 ;
        RECT 88.200 130.300 88.600 130.700 ;
        RECT 88.900 130.300 89.300 130.700 ;
        RECT 191.400 130.300 191.800 130.700 ;
        RECT 192.100 130.300 192.500 130.700 ;
        RECT 88.200 110.300 88.600 110.700 ;
        RECT 88.900 110.300 89.300 110.700 ;
        RECT 191.400 110.300 191.800 110.700 ;
        RECT 192.100 110.300 192.500 110.700 ;
        RECT 88.200 90.300 88.600 90.700 ;
        RECT 88.900 90.300 89.300 90.700 ;
        RECT 191.400 90.300 191.800 90.700 ;
        RECT 192.100 90.300 192.500 90.700 ;
        RECT 88.200 70.300 88.600 70.700 ;
        RECT 88.900 70.300 89.300 70.700 ;
        RECT 191.400 70.300 191.800 70.700 ;
        RECT 192.100 70.300 192.500 70.700 ;
        RECT 88.200 50.300 88.600 50.700 ;
        RECT 88.900 50.300 89.300 50.700 ;
        RECT 191.400 50.300 191.800 50.700 ;
        RECT 192.100 50.300 192.500 50.700 ;
        RECT 88.200 30.300 88.600 30.700 ;
        RECT 88.900 30.300 89.300 30.700 ;
        RECT 191.400 30.300 191.800 30.700 ;
        RECT 192.100 30.300 192.500 30.700 ;
        RECT 88.200 10.300 88.600 10.700 ;
        RECT 88.900 10.300 89.300 10.700 ;
        RECT 191.400 10.300 191.800 10.700 ;
        RECT 192.100 10.300 192.500 10.700 ;
      LAYER metal2 ;
        RECT 88.000 210.300 89.600 210.700 ;
        RECT 191.200 210.300 192.800 210.700 ;
        RECT 88.000 190.300 89.600 190.700 ;
        RECT 191.200 190.300 192.800 190.700 ;
        RECT 88.000 170.300 89.600 170.700 ;
        RECT 191.200 170.300 192.800 170.700 ;
        RECT 88.000 150.300 89.600 150.700 ;
        RECT 191.200 150.300 192.800 150.700 ;
        RECT 88.000 130.300 89.600 130.700 ;
        RECT 191.200 130.300 192.800 130.700 ;
        RECT 88.000 110.300 89.600 110.700 ;
        RECT 191.200 110.300 192.800 110.700 ;
        RECT 88.000 90.300 89.600 90.700 ;
        RECT 191.200 90.300 192.800 90.700 ;
        RECT 88.000 70.300 89.600 70.700 ;
        RECT 191.200 70.300 192.800 70.700 ;
        RECT 88.000 50.300 89.600 50.700 ;
        RECT 191.200 50.300 192.800 50.700 ;
        RECT 88.000 30.300 89.600 30.700 ;
        RECT 191.200 30.300 192.800 30.700 ;
        RECT 88.000 10.300 89.600 10.700 ;
        RECT 191.200 10.300 192.800 10.700 ;
      LAYER via2 ;
        RECT 88.200 210.300 88.600 210.700 ;
        RECT 88.900 210.300 89.300 210.700 ;
        RECT 191.400 210.300 191.800 210.700 ;
        RECT 192.100 210.300 192.500 210.700 ;
        RECT 88.200 190.300 88.600 190.700 ;
        RECT 88.900 190.300 89.300 190.700 ;
        RECT 191.400 190.300 191.800 190.700 ;
        RECT 192.100 190.300 192.500 190.700 ;
        RECT 88.200 170.300 88.600 170.700 ;
        RECT 88.900 170.300 89.300 170.700 ;
        RECT 191.400 170.300 191.800 170.700 ;
        RECT 192.100 170.300 192.500 170.700 ;
        RECT 88.200 150.300 88.600 150.700 ;
        RECT 88.900 150.300 89.300 150.700 ;
        RECT 191.400 150.300 191.800 150.700 ;
        RECT 192.100 150.300 192.500 150.700 ;
        RECT 88.200 130.300 88.600 130.700 ;
        RECT 88.900 130.300 89.300 130.700 ;
        RECT 191.400 130.300 191.800 130.700 ;
        RECT 192.100 130.300 192.500 130.700 ;
        RECT 88.200 110.300 88.600 110.700 ;
        RECT 88.900 110.300 89.300 110.700 ;
        RECT 191.400 110.300 191.800 110.700 ;
        RECT 192.100 110.300 192.500 110.700 ;
        RECT 88.200 90.300 88.600 90.700 ;
        RECT 88.900 90.300 89.300 90.700 ;
        RECT 191.400 90.300 191.800 90.700 ;
        RECT 192.100 90.300 192.500 90.700 ;
        RECT 88.200 70.300 88.600 70.700 ;
        RECT 88.900 70.300 89.300 70.700 ;
        RECT 191.400 70.300 191.800 70.700 ;
        RECT 192.100 70.300 192.500 70.700 ;
        RECT 88.200 50.300 88.600 50.700 ;
        RECT 88.900 50.300 89.300 50.700 ;
        RECT 191.400 50.300 191.800 50.700 ;
        RECT 192.100 50.300 192.500 50.700 ;
        RECT 88.200 30.300 88.600 30.700 ;
        RECT 88.900 30.300 89.300 30.700 ;
        RECT 191.400 30.300 191.800 30.700 ;
        RECT 192.100 30.300 192.500 30.700 ;
        RECT 88.200 10.300 88.600 10.700 ;
        RECT 88.900 10.300 89.300 10.700 ;
        RECT 191.400 10.300 191.800 10.700 ;
        RECT 192.100 10.300 192.500 10.700 ;
      LAYER metal3 ;
        RECT 88.000 210.300 89.600 210.700 ;
        RECT 191.200 210.300 192.800 210.700 ;
        RECT 88.000 190.300 89.600 190.700 ;
        RECT 191.200 190.300 192.800 190.700 ;
        RECT 88.000 170.300 89.600 170.700 ;
        RECT 191.200 170.300 192.800 170.700 ;
        RECT 88.000 150.300 89.600 150.700 ;
        RECT 191.200 150.300 192.800 150.700 ;
        RECT 88.000 130.300 89.600 130.700 ;
        RECT 191.200 130.300 192.800 130.700 ;
        RECT 88.000 110.300 89.600 110.700 ;
        RECT 191.200 110.300 192.800 110.700 ;
        RECT 88.000 90.300 89.600 90.700 ;
        RECT 191.200 90.300 192.800 90.700 ;
        RECT 88.000 70.300 89.600 70.700 ;
        RECT 191.200 70.300 192.800 70.700 ;
        RECT 88.000 50.300 89.600 50.700 ;
        RECT 191.200 50.300 192.800 50.700 ;
        RECT 88.000 30.300 89.600 30.700 ;
        RECT 191.200 30.300 192.800 30.700 ;
        RECT 88.000 10.300 89.600 10.700 ;
        RECT 191.200 10.300 192.800 10.700 ;
      LAYER via3 ;
        RECT 88.200 210.300 88.600 210.700 ;
        RECT 89.000 210.300 89.400 210.700 ;
        RECT 191.400 210.300 191.800 210.700 ;
        RECT 192.200 210.300 192.600 210.700 ;
        RECT 88.200 190.300 88.600 190.700 ;
        RECT 89.000 190.300 89.400 190.700 ;
        RECT 191.400 190.300 191.800 190.700 ;
        RECT 192.200 190.300 192.600 190.700 ;
        RECT 88.200 170.300 88.600 170.700 ;
        RECT 89.000 170.300 89.400 170.700 ;
        RECT 191.400 170.300 191.800 170.700 ;
        RECT 192.200 170.300 192.600 170.700 ;
        RECT 88.200 150.300 88.600 150.700 ;
        RECT 89.000 150.300 89.400 150.700 ;
        RECT 191.400 150.300 191.800 150.700 ;
        RECT 192.200 150.300 192.600 150.700 ;
        RECT 88.200 130.300 88.600 130.700 ;
        RECT 89.000 130.300 89.400 130.700 ;
        RECT 191.400 130.300 191.800 130.700 ;
        RECT 192.200 130.300 192.600 130.700 ;
        RECT 88.200 110.300 88.600 110.700 ;
        RECT 89.000 110.300 89.400 110.700 ;
        RECT 191.400 110.300 191.800 110.700 ;
        RECT 192.200 110.300 192.600 110.700 ;
        RECT 88.200 90.300 88.600 90.700 ;
        RECT 89.000 90.300 89.400 90.700 ;
        RECT 191.400 90.300 191.800 90.700 ;
        RECT 192.200 90.300 192.600 90.700 ;
        RECT 88.200 70.300 88.600 70.700 ;
        RECT 89.000 70.300 89.400 70.700 ;
        RECT 191.400 70.300 191.800 70.700 ;
        RECT 192.200 70.300 192.600 70.700 ;
        RECT 88.200 50.300 88.600 50.700 ;
        RECT 89.000 50.300 89.400 50.700 ;
        RECT 191.400 50.300 191.800 50.700 ;
        RECT 192.200 50.300 192.600 50.700 ;
        RECT 88.200 30.300 88.600 30.700 ;
        RECT 89.000 30.300 89.400 30.700 ;
        RECT 191.400 30.300 191.800 30.700 ;
        RECT 192.200 30.300 192.600 30.700 ;
        RECT 88.200 10.300 88.600 10.700 ;
        RECT 89.000 10.300 89.400 10.700 ;
        RECT 191.400 10.300 191.800 10.700 ;
        RECT 192.200 10.300 192.600 10.700 ;
      LAYER metal4 ;
        RECT 88.000 210.300 89.600 210.700 ;
        RECT 191.200 210.300 192.800 210.700 ;
        RECT 88.000 190.300 89.600 190.700 ;
        RECT 191.200 190.300 192.800 190.700 ;
        RECT 88.000 170.300 89.600 170.700 ;
        RECT 191.200 170.300 192.800 170.700 ;
        RECT 88.000 150.300 89.600 150.700 ;
        RECT 191.200 150.300 192.800 150.700 ;
        RECT 88.000 130.300 89.600 130.700 ;
        RECT 191.200 130.300 192.800 130.700 ;
        RECT 88.000 110.300 89.600 110.700 ;
        RECT 191.200 110.300 192.800 110.700 ;
        RECT 88.000 90.300 89.600 90.700 ;
        RECT 191.200 90.300 192.800 90.700 ;
        RECT 88.000 70.300 89.600 70.700 ;
        RECT 191.200 70.300 192.800 70.700 ;
        RECT 88.000 50.300 89.600 50.700 ;
        RECT 191.200 50.300 192.800 50.700 ;
        RECT 88.000 30.300 89.600 30.700 ;
        RECT 191.200 30.300 192.800 30.700 ;
        RECT 88.000 10.300 89.600 10.700 ;
        RECT 191.200 10.300 192.800 10.700 ;
      LAYER via4 ;
        RECT 88.200 210.300 88.600 210.700 ;
        RECT 88.900 210.300 89.300 210.700 ;
        RECT 191.400 210.300 191.800 210.700 ;
        RECT 192.100 210.300 192.500 210.700 ;
        RECT 88.200 190.300 88.600 190.700 ;
        RECT 88.900 190.300 89.300 190.700 ;
        RECT 191.400 190.300 191.800 190.700 ;
        RECT 192.100 190.300 192.500 190.700 ;
        RECT 88.200 170.300 88.600 170.700 ;
        RECT 88.900 170.300 89.300 170.700 ;
        RECT 191.400 170.300 191.800 170.700 ;
        RECT 192.100 170.300 192.500 170.700 ;
        RECT 88.200 150.300 88.600 150.700 ;
        RECT 88.900 150.300 89.300 150.700 ;
        RECT 191.400 150.300 191.800 150.700 ;
        RECT 192.100 150.300 192.500 150.700 ;
        RECT 88.200 130.300 88.600 130.700 ;
        RECT 88.900 130.300 89.300 130.700 ;
        RECT 191.400 130.300 191.800 130.700 ;
        RECT 192.100 130.300 192.500 130.700 ;
        RECT 88.200 110.300 88.600 110.700 ;
        RECT 88.900 110.300 89.300 110.700 ;
        RECT 191.400 110.300 191.800 110.700 ;
        RECT 192.100 110.300 192.500 110.700 ;
        RECT 88.200 90.300 88.600 90.700 ;
        RECT 88.900 90.300 89.300 90.700 ;
        RECT 191.400 90.300 191.800 90.700 ;
        RECT 192.100 90.300 192.500 90.700 ;
        RECT 88.200 70.300 88.600 70.700 ;
        RECT 88.900 70.300 89.300 70.700 ;
        RECT 191.400 70.300 191.800 70.700 ;
        RECT 192.100 70.300 192.500 70.700 ;
        RECT 88.200 50.300 88.600 50.700 ;
        RECT 88.900 50.300 89.300 50.700 ;
        RECT 191.400 50.300 191.800 50.700 ;
        RECT 192.100 50.300 192.500 50.700 ;
        RECT 88.200 30.300 88.600 30.700 ;
        RECT 88.900 30.300 89.300 30.700 ;
        RECT 191.400 30.300 191.800 30.700 ;
        RECT 192.100 30.300 192.500 30.700 ;
        RECT 88.200 10.300 88.600 10.700 ;
        RECT 88.900 10.300 89.300 10.700 ;
        RECT 191.400 10.300 191.800 10.700 ;
        RECT 192.100 10.300 192.500 10.700 ;
      LAYER metal5 ;
        RECT 88.000 210.200 89.600 210.700 ;
        RECT 191.200 210.200 192.800 210.700 ;
        RECT 88.000 190.200 89.600 190.700 ;
        RECT 191.200 190.200 192.800 190.700 ;
        RECT 88.000 170.200 89.600 170.700 ;
        RECT 191.200 170.200 192.800 170.700 ;
        RECT 88.000 150.200 89.600 150.700 ;
        RECT 191.200 150.200 192.800 150.700 ;
        RECT 88.000 130.200 89.600 130.700 ;
        RECT 191.200 130.200 192.800 130.700 ;
        RECT 88.000 110.200 89.600 110.700 ;
        RECT 191.200 110.200 192.800 110.700 ;
        RECT 88.000 90.200 89.600 90.700 ;
        RECT 191.200 90.200 192.800 90.700 ;
        RECT 88.000 70.200 89.600 70.700 ;
        RECT 191.200 70.200 192.800 70.700 ;
        RECT 88.000 50.200 89.600 50.700 ;
        RECT 191.200 50.200 192.800 50.700 ;
        RECT 88.000 30.200 89.600 30.700 ;
        RECT 191.200 30.200 192.800 30.700 ;
        RECT 88.000 10.200 89.600 10.700 ;
        RECT 191.200 10.200 192.800 10.700 ;
      LAYER via5 ;
        RECT 89.000 210.200 89.500 210.700 ;
        RECT 192.200 210.200 192.700 210.700 ;
        RECT 89.000 190.200 89.500 190.700 ;
        RECT 192.200 190.200 192.700 190.700 ;
        RECT 89.000 170.200 89.500 170.700 ;
        RECT 192.200 170.200 192.700 170.700 ;
        RECT 89.000 150.200 89.500 150.700 ;
        RECT 192.200 150.200 192.700 150.700 ;
        RECT 89.000 130.200 89.500 130.700 ;
        RECT 192.200 130.200 192.700 130.700 ;
        RECT 89.000 110.200 89.500 110.700 ;
        RECT 192.200 110.200 192.700 110.700 ;
        RECT 89.000 90.200 89.500 90.700 ;
        RECT 192.200 90.200 192.700 90.700 ;
        RECT 89.000 70.200 89.500 70.700 ;
        RECT 192.200 70.200 192.700 70.700 ;
        RECT 89.000 50.200 89.500 50.700 ;
        RECT 192.200 50.200 192.700 50.700 ;
        RECT 89.000 30.200 89.500 30.700 ;
        RECT 192.200 30.200 192.700 30.700 ;
        RECT 89.000 10.200 89.500 10.700 ;
        RECT 192.200 10.200 192.700 10.700 ;
      LAYER metal6 ;
        RECT 88.000 -3.000 89.600 213.000 ;
        RECT 191.200 -3.000 192.800 213.000 ;
    END
  END gnd
  PIN en
    PORT
      LAYER metal1 ;
        RECT 175.800 3.800 176.200 5.200 ;
      LAYER metal2 ;
        RECT 175.800 3.800 176.200 4.200 ;
        RECT 175.000 -1.900 175.400 -1.800 ;
        RECT 175.800 -1.900 176.100 3.800 ;
        RECT 175.000 -2.200 176.100 -1.900 ;
    END
  END en
  PIN rw
    PORT
      LAYER metal1 ;
        RECT 161.400 113.400 161.800 114.200 ;
        RECT 166.200 112.800 166.600 113.200 ;
        RECT 169.400 112.800 169.800 113.200 ;
        RECT 166.100 112.400 166.500 112.800 ;
        RECT 169.300 112.400 169.700 112.800 ;
        RECT 203.000 106.800 203.400 107.600 ;
        RECT 154.900 88.200 155.300 88.600 ;
        RECT 158.100 88.200 158.500 88.600 ;
        RECT 155.000 87.800 155.400 88.200 ;
        RECT 158.200 87.800 158.600 88.200 ;
        RECT 155.000 87.200 155.300 87.800 ;
        RECT 155.000 86.800 155.400 87.200 ;
        RECT 157.300 68.200 157.700 68.600 ;
        RECT 163.700 68.200 164.100 68.600 ;
        RECT 157.400 67.800 157.800 68.200 ;
        RECT 163.800 67.800 164.200 68.200 ;
      LAYER via1 ;
        RECT 161.400 113.800 161.800 114.200 ;
      LAYER metal2 ;
        RECT 161.400 113.800 161.800 114.200 ;
        RECT 161.400 113.200 161.700 113.800 ;
        RECT 161.400 112.800 161.800 113.200 ;
        RECT 165.400 113.100 165.800 113.200 ;
        RECT 166.200 113.100 166.600 113.200 ;
        RECT 165.400 112.800 166.600 113.100 ;
        RECT 168.600 113.100 169.000 113.200 ;
        RECT 169.400 113.100 169.800 113.200 ;
        RECT 168.600 112.800 169.800 113.100 ;
        RECT 161.400 101.200 161.700 112.800 ;
        RECT 169.400 109.200 169.700 112.800 ;
        RECT 169.400 108.800 169.800 109.200 ;
        RECT 203.000 108.800 203.400 109.200 ;
        RECT 203.000 108.200 203.300 108.800 ;
        RECT 203.000 107.800 203.400 108.200 ;
        RECT 203.000 107.200 203.300 107.800 ;
        RECT 203.000 106.800 203.400 107.200 ;
        RECT 158.200 100.800 158.600 101.200 ;
        RECT 161.400 100.800 161.800 101.200 ;
        RECT 158.200 88.200 158.500 100.800 ;
        RECT 155.000 87.800 155.400 88.200 ;
        RECT 157.400 88.100 157.800 88.200 ;
        RECT 158.200 88.100 158.600 88.200 ;
        RECT 157.400 87.800 158.600 88.100 ;
        RECT 155.000 87.200 155.300 87.800 ;
        RECT 155.000 86.800 155.400 87.200 ;
        RECT 158.200 73.100 158.500 87.800 ;
        RECT 157.400 72.800 158.500 73.100 ;
        RECT 157.400 68.200 157.700 72.800 ;
        RECT 157.400 67.800 157.800 68.200 ;
        RECT 163.800 67.800 164.200 68.200 ;
        RECT 157.400 67.200 157.700 67.800 ;
        RECT 163.800 67.200 164.100 67.800 ;
        RECT 157.400 66.800 157.800 67.200 ;
        RECT 163.800 66.800 164.200 67.200 ;
      LAYER metal3 ;
        RECT 161.400 113.100 161.800 113.200 ;
        RECT 165.400 113.100 165.800 113.200 ;
        RECT 168.600 113.100 169.000 113.200 ;
        RECT 161.400 112.800 169.000 113.100 ;
        RECT 169.400 109.100 169.800 109.200 ;
        RECT 203.000 109.100 203.400 109.200 ;
        RECT 169.400 108.800 203.400 109.100 ;
        RECT 203.000 108.100 203.400 108.200 ;
        RECT 203.000 107.800 224.100 108.100 ;
        RECT 223.800 107.100 224.100 107.800 ;
        RECT 233.400 107.100 233.800 107.200 ;
        RECT 223.800 106.800 233.800 107.100 ;
        RECT 158.200 101.100 158.600 101.200 ;
        RECT 161.400 101.100 161.800 101.200 ;
        RECT 158.200 100.800 161.800 101.100 ;
        RECT 155.000 88.100 155.400 88.200 ;
        RECT 157.400 88.100 157.800 88.200 ;
        RECT 155.000 87.800 157.800 88.100 ;
        RECT 157.400 67.100 157.800 67.200 ;
        RECT 163.800 67.100 164.200 67.200 ;
        RECT 157.400 66.800 164.200 67.100 ;
    END
  END rw
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 0.600 206.900 1.000 207.200 ;
        RECT 7.800 206.900 8.200 207.200 ;
        RECT 197.400 206.900 197.800 207.200 ;
        RECT 0.600 206.500 1.500 206.900 ;
        RECT 7.800 206.500 8.700 206.900 ;
        RECT 196.900 206.500 197.800 206.900 ;
        RECT 0.600 174.100 1.500 174.500 ;
        RECT 17.400 174.100 18.300 174.500 ;
        RECT 0.600 173.800 1.000 174.100 ;
        RECT 17.400 173.800 17.800 174.100 ;
        RECT 223.800 166.900 224.200 167.200 ;
        RECT 223.800 166.500 224.700 166.900 ;
        RECT 75.000 86.900 75.400 87.200 ;
        RECT 74.500 86.500 75.400 86.900 ;
        RECT 221.400 74.100 222.300 74.500 ;
        RECT 221.400 73.800 221.800 74.100 ;
        RECT 21.400 54.100 22.300 54.500 ;
        RECT 21.400 53.800 21.800 54.100 ;
        RECT 36.600 26.900 37.000 27.200 ;
        RECT 36.100 26.500 37.000 26.900 ;
        RECT 127.800 26.900 128.200 27.200 ;
        RECT 135.000 26.900 135.400 27.200 ;
        RECT 127.800 26.500 128.700 26.900 ;
        RECT 135.000 26.500 135.900 26.900 ;
        RECT 217.400 14.100 218.300 14.500 ;
        RECT 217.400 13.800 217.800 14.100 ;
        RECT 22.200 7.100 22.600 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 22.200 6.900 23.400 7.100 ;
        RECT 22.200 6.800 23.900 6.900 ;
        RECT 23.000 6.500 23.900 6.800 ;
      LAYER via1 ;
        RECT 0.600 206.800 1.000 207.200 ;
        RECT 7.800 206.800 8.200 207.200 ;
        RECT 197.400 206.800 197.800 207.200 ;
        RECT 223.800 166.800 224.200 167.200 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 36.600 26.800 37.000 27.200 ;
        RECT 127.800 26.800 128.200 27.200 ;
        RECT 135.000 26.800 135.400 27.200 ;
      LAYER metal2 ;
        RECT 0.600 206.800 1.000 207.200 ;
        RECT 7.800 206.800 8.200 207.200 ;
        RECT 197.400 206.800 197.800 207.200 ;
        RECT 0.600 205.200 0.900 206.800 ;
        RECT 7.800 205.200 8.100 206.800 ;
        RECT 0.600 204.800 1.000 205.200 ;
        RECT 7.800 204.800 8.200 205.200 ;
        RECT 197.400 183.200 197.700 206.800 ;
        RECT 197.400 182.800 197.800 183.200 ;
        RECT 0.600 173.800 1.000 174.200 ;
        RECT 17.400 173.800 17.800 174.200 ;
        RECT 0.600 171.200 0.900 173.800 ;
        RECT 17.400 171.200 17.700 173.800 ;
        RECT 0.600 170.800 1.000 171.200 ;
        RECT 17.400 170.800 17.800 171.200 ;
        RECT 223.000 167.100 223.400 167.200 ;
        RECT 223.800 167.100 224.200 167.200 ;
        RECT 223.000 166.800 224.200 167.100 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 75.000 83.200 75.300 86.800 ;
        RECT 75.000 82.800 75.400 83.200 ;
        RECT 221.400 73.800 221.800 74.200 ;
        RECT 221.400 73.200 221.700 73.800 ;
        RECT 221.400 72.800 221.800 73.200 ;
        RECT 21.400 53.800 21.800 54.200 ;
        RECT 21.400 50.200 21.700 53.800 ;
        RECT 21.400 49.800 21.800 50.200 ;
        RECT 36.600 49.800 37.000 50.200 ;
        RECT 36.600 27.200 36.900 49.800 ;
        RECT 127.800 27.800 128.200 28.200 ;
        RECT 135.000 27.800 135.400 28.200 ;
        RECT 127.800 27.200 128.100 27.800 ;
        RECT 135.000 27.200 135.300 27.800 ;
        RECT 36.600 26.800 37.000 27.200 ;
        RECT 127.800 26.800 128.200 27.200 ;
        RECT 135.000 26.800 135.400 27.200 ;
        RECT 36.600 20.200 36.900 26.800 ;
        RECT 22.200 19.800 22.600 20.200 ;
        RECT 36.600 19.800 37.000 20.200 ;
        RECT 22.200 7.200 22.500 19.800 ;
        RECT 135.000 18.200 135.300 26.800 ;
        RECT 135.000 17.800 135.400 18.200 ;
        RECT 217.400 17.800 217.800 18.200 ;
        RECT 217.400 14.200 217.700 17.800 ;
        RECT 217.400 13.800 217.800 14.200 ;
        RECT 22.200 6.800 22.600 7.200 ;
      LAYER metal3 ;
        RECT -2.600 205.100 -2.200 205.200 ;
        RECT 0.600 205.100 1.000 205.200 ;
        RECT 7.800 205.100 8.200 205.200 ;
        RECT -2.600 204.800 8.200 205.100 ;
        RECT 197.400 183.100 197.800 183.200 ;
        RECT 219.800 183.100 220.200 183.200 ;
        RECT 197.400 182.800 220.200 183.100 ;
        RECT 0.600 171.100 1.000 171.200 ;
        RECT 17.400 171.100 17.800 171.200 ;
        RECT 46.200 171.100 46.600 171.200 ;
        RECT 0.600 170.800 46.600 171.100 ;
        RECT 219.800 167.100 220.200 167.200 ;
        RECT 223.000 167.100 223.400 167.200 ;
        RECT 219.800 166.800 223.400 167.100 ;
        RECT 44.600 83.100 45.000 83.200 ;
        RECT 46.200 83.100 46.600 83.200 ;
        RECT 75.000 83.100 75.400 83.200 ;
        RECT 107.800 83.100 108.200 83.200 ;
        RECT 44.600 82.800 108.200 83.100 ;
        RECT 219.800 74.100 220.200 74.200 ;
        RECT 219.800 73.800 221.700 74.100 ;
        RECT 221.400 73.200 221.700 73.800 ;
        RECT 221.400 72.800 221.800 73.200 ;
        RECT 21.400 50.100 21.800 50.200 ;
        RECT 36.600 50.100 37.000 50.200 ;
        RECT 44.600 50.100 45.000 50.200 ;
        RECT 21.400 49.800 45.000 50.100 ;
        RECT 107.800 28.100 108.200 28.200 ;
        RECT 127.800 28.100 128.200 28.200 ;
        RECT 135.000 28.100 135.400 28.200 ;
        RECT 107.800 27.800 135.400 28.100 ;
        RECT 22.200 20.100 22.600 20.200 ;
        RECT 36.600 20.100 37.000 20.200 ;
        RECT 22.200 19.800 37.000 20.100 ;
        RECT 135.000 18.100 135.400 18.200 ;
        RECT 217.400 18.100 217.800 18.200 ;
        RECT 219.800 18.100 220.200 18.200 ;
        RECT 135.000 17.800 220.200 18.100 ;
      LAYER via3 ;
        RECT 0.600 204.800 1.000 205.200 ;
        RECT 219.800 182.800 220.200 183.200 ;
        RECT 46.200 170.800 46.600 171.200 ;
        RECT 46.200 82.800 46.600 83.200 ;
        RECT 107.800 82.800 108.200 83.200 ;
        RECT 44.600 49.800 45.000 50.200 ;
        RECT 219.800 17.800 220.200 18.200 ;
      LAYER metal4 ;
        RECT 0.600 204.800 1.000 205.200 ;
        RECT 0.600 171.200 0.900 204.800 ;
        RECT 219.800 182.800 220.200 183.200 ;
        RECT 0.600 170.800 1.000 171.200 ;
        RECT 46.200 170.800 46.600 171.200 ;
        RECT 46.200 83.200 46.500 170.800 ;
        RECT 219.800 167.200 220.100 182.800 ;
        RECT 219.800 166.800 220.200 167.200 ;
        RECT 44.600 82.800 45.000 83.200 ;
        RECT 46.200 82.800 46.600 83.200 ;
        RECT 107.800 82.800 108.200 83.200 ;
        RECT 44.600 50.200 44.900 82.800 ;
        RECT 44.600 49.800 45.000 50.200 ;
        RECT 107.800 28.200 108.100 82.800 ;
        RECT 219.800 74.200 220.100 166.800 ;
        RECT 219.800 73.800 220.200 74.200 ;
        RECT 107.800 27.800 108.200 28.200 ;
        RECT 219.800 18.200 220.100 73.800 ;
        RECT 219.800 17.800 220.200 18.200 ;
    END
  END clk
  PIN ras
    PORT
      LAYER metal1 ;
        RECT 86.200 8.100 86.600 8.600 ;
        RECT 87.000 8.100 87.400 8.600 ;
        RECT 86.200 7.800 87.400 8.100 ;
        RECT 86.200 7.200 86.500 7.800 ;
        RECT 86.200 6.800 86.600 7.200 ;
        RECT 174.200 6.800 174.600 7.600 ;
        RECT 80.600 6.100 81.000 6.200 ;
        RECT 81.400 6.100 81.800 6.200 ;
        RECT 80.200 5.800 82.200 6.100 ;
        RECT 80.200 5.600 80.600 5.800 ;
        RECT 81.800 5.600 82.200 5.800 ;
      LAYER via1 ;
        RECT 81.400 5.800 81.800 6.200 ;
      LAYER metal2 ;
        RECT 81.400 7.800 81.800 8.200 ;
        RECT 86.200 7.800 86.600 8.200 ;
        RECT 81.400 6.200 81.700 7.800 ;
        RECT 86.200 7.200 86.500 7.800 ;
        RECT 86.200 6.800 86.600 7.200 ;
        RECT 174.200 6.800 174.600 7.200 ;
        RECT 174.200 6.200 174.500 6.800 ;
        RECT 81.400 5.800 81.800 6.200 ;
        RECT 174.200 5.800 174.600 6.200 ;
        RECT 81.400 -1.800 81.700 5.800 ;
        RECT 81.400 -2.200 81.800 -1.800 ;
      LAYER metal3 ;
        RECT 81.400 8.100 81.800 8.200 ;
        RECT 86.200 8.100 86.600 8.200 ;
        RECT 81.400 7.800 99.300 8.100 ;
        RECT 99.000 7.100 99.300 7.800 ;
        RECT 99.000 6.800 174.500 7.100 ;
        RECT 174.200 6.200 174.500 6.800 ;
        RECT 174.200 5.800 174.600 6.200 ;
    END
  END ras
  PIN cas
    PORT
      LAYER metal1 ;
        RECT 184.600 7.800 185.000 8.600 ;
        RECT 180.600 7.100 181.000 7.600 ;
        RECT 184.600 7.200 184.900 7.800 ;
        RECT 181.400 7.100 181.800 7.200 ;
        RECT 180.600 6.800 181.800 7.100 ;
        RECT 184.600 6.800 185.000 7.200 ;
        RECT 181.400 6.200 181.700 6.800 ;
        RECT 181.400 6.100 181.800 6.200 ;
        RECT 181.400 5.800 182.200 6.100 ;
        RECT 181.800 5.600 182.200 5.800 ;
      LAYER via1 ;
        RECT 181.400 6.800 181.800 7.200 ;
      LAYER metal2 ;
        RECT 181.400 7.800 181.800 8.200 ;
        RECT 184.600 7.800 185.000 8.200 ;
        RECT 181.400 7.200 181.700 7.800 ;
        RECT 184.600 7.200 184.900 7.800 ;
        RECT 181.400 6.800 181.800 7.200 ;
        RECT 184.600 6.800 185.000 7.200 ;
        RECT 181.400 -1.800 181.700 6.800 ;
        RECT 181.400 -2.200 181.800 -1.800 ;
      LAYER metal3 ;
        RECT 181.400 8.100 181.800 8.200 ;
        RECT 184.600 8.100 185.000 8.200 ;
        RECT 181.400 7.800 185.000 8.100 ;
    END
  END cas
  PIN vas
    PORT
      LAYER metal1 ;
        RECT 190.200 7.800 190.600 8.600 ;
        RECT 197.400 7.800 197.800 8.600 ;
        RECT 187.000 6.100 187.400 6.200 ;
        RECT 194.200 6.100 194.600 6.200 ;
        RECT 187.000 5.800 187.800 6.100 ;
        RECT 194.200 5.800 195.000 6.100 ;
        RECT 187.400 5.600 187.800 5.800 ;
        RECT 194.600 5.600 195.000 5.800 ;
        RECT 179.000 4.400 179.400 5.200 ;
      LAYER via1 ;
        RECT 179.000 4.800 179.400 5.200 ;
      LAYER metal2 ;
        RECT 190.200 7.800 190.600 8.200 ;
        RECT 197.400 7.800 197.800 8.200 ;
        RECT 190.200 6.200 190.500 7.800 ;
        RECT 197.400 6.200 197.700 7.800 ;
        RECT 179.000 5.800 179.400 6.200 ;
        RECT 179.800 5.800 180.200 6.200 ;
        RECT 187.000 6.100 187.400 6.200 ;
        RECT 187.800 6.100 188.200 6.200 ;
        RECT 187.000 5.800 188.200 6.100 ;
        RECT 190.200 5.800 190.600 6.200 ;
        RECT 193.400 6.100 193.800 6.200 ;
        RECT 194.200 6.100 194.600 6.200 ;
        RECT 193.400 5.800 194.600 6.100 ;
        RECT 197.400 5.800 197.800 6.200 ;
        RECT 179.000 5.200 179.300 5.800 ;
        RECT 179.000 4.800 179.400 5.200 ;
        RECT 179.800 -1.800 180.100 5.800 ;
        RECT 179.800 -2.200 180.200 -1.800 ;
      LAYER via2 ;
        RECT 187.800 5.800 188.200 6.200 ;
      LAYER metal3 ;
        RECT 179.000 6.100 179.400 6.200 ;
        RECT 179.800 6.100 180.200 6.200 ;
        RECT 187.800 6.100 188.200 6.200 ;
        RECT 190.200 6.100 190.600 6.200 ;
        RECT 193.400 6.100 193.800 6.200 ;
        RECT 197.400 6.100 197.800 6.200 ;
        RECT 179.000 5.800 197.800 6.100 ;
    END
  END vas
  PIN datain[0]
    PORT
      LAYER metal1 ;
        RECT 0.600 113.400 1.000 114.200 ;
      LAYER via1 ;
        RECT 0.600 113.800 1.000 114.200 ;
      LAYER metal2 ;
        RECT 0.600 114.800 1.000 115.200 ;
        RECT 0.600 114.200 0.900 114.800 ;
        RECT 0.600 113.800 1.000 114.200 ;
      LAYER metal3 ;
        RECT -2.600 115.100 -2.200 115.200 ;
        RECT 0.600 115.100 1.000 115.200 ;
        RECT -2.600 114.800 1.000 115.100 ;
    END
  END datain[0]
  PIN datain[1]
    PORT
      LAYER metal1 ;
        RECT 188.600 206.800 189.000 207.600 ;
      LAYER metal2 ;
        RECT 187.000 212.800 187.400 213.200 ;
        RECT 187.000 208.200 187.300 212.800 ;
        RECT 187.000 207.800 187.400 208.200 ;
        RECT 188.600 207.800 189.000 208.200 ;
        RECT 188.600 207.200 188.900 207.800 ;
        RECT 188.600 206.800 189.000 207.200 ;
      LAYER metal3 ;
        RECT 187.000 208.100 187.400 208.200 ;
        RECT 188.600 208.100 189.000 208.200 ;
        RECT 187.000 207.800 189.000 208.100 ;
    END
  END datain[1]
  PIN datain[2]
    PORT
      LAYER metal1 ;
        RECT 15.800 6.800 16.200 7.600 ;
      LAYER metal2 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 15.800 -1.900 16.100 6.800 ;
        RECT 17.400 -1.900 17.800 -1.800 ;
        RECT 15.800 -2.200 17.800 -1.900 ;
    END
  END datain[2]
  PIN datain[3]
    PORT
      LAYER metal1 ;
        RECT 0.600 66.800 1.000 67.600 ;
      LAYER metal2 ;
        RECT 0.600 66.800 1.000 67.200 ;
        RECT 0.600 65.200 0.900 66.800 ;
        RECT 0.600 64.800 1.000 65.200 ;
      LAYER metal3 ;
        RECT -2.600 65.100 -2.200 65.200 ;
        RECT 0.600 65.100 1.000 65.200 ;
        RECT -2.600 64.800 1.000 65.100 ;
    END
  END datain[3]
  PIN datain[4]
    PORT
      LAYER metal1 ;
        RECT 109.400 6.800 109.800 7.600 ;
      LAYER metal2 ;
        RECT 109.400 6.800 109.800 7.200 ;
        RECT 109.400 1.200 109.700 6.800 ;
        RECT 107.800 0.800 108.200 1.200 ;
        RECT 109.400 0.800 109.800 1.200 ;
        RECT 107.800 -1.800 108.100 0.800 ;
        RECT 107.800 -2.200 108.200 -1.800 ;
      LAYER metal3 ;
        RECT 107.800 1.100 108.200 1.200 ;
        RECT 109.400 1.100 109.800 1.200 ;
        RECT 107.800 0.800 109.800 1.100 ;
    END
  END datain[4]
  PIN datain[5]
    PORT
      LAYER metal1 ;
        RECT 229.400 207.100 229.800 207.600 ;
        RECT 230.200 207.100 230.600 207.200 ;
        RECT 229.400 206.800 230.600 207.100 ;
      LAYER via1 ;
        RECT 230.200 206.800 230.600 207.200 ;
      LAYER metal2 ;
        RECT 230.200 206.800 230.600 207.200 ;
        RECT 230.200 205.200 230.500 206.800 ;
        RECT 230.200 204.800 230.600 205.200 ;
      LAYER metal3 ;
        RECT 230.200 205.100 230.600 205.200 ;
        RECT 233.400 205.100 233.800 205.200 ;
        RECT 230.200 204.800 233.800 205.100 ;
    END
  END datain[5]
  PIN datain[6]
    PORT
      LAYER metal1 ;
        RECT 136.600 206.800 137.000 207.600 ;
      LAYER metal2 ;
        RECT 138.200 212.800 138.600 213.200 ;
        RECT 138.200 208.200 138.500 212.800 ;
        RECT 136.600 207.800 137.000 208.200 ;
        RECT 138.200 207.800 138.600 208.200 ;
        RECT 136.600 207.200 136.900 207.800 ;
        RECT 136.600 206.800 137.000 207.200 ;
      LAYER metal3 ;
        RECT 136.600 208.100 137.000 208.200 ;
        RECT 138.200 208.100 138.600 208.200 ;
        RECT 136.600 207.800 138.600 208.100 ;
    END
  END datain[6]
  PIN datain[7]
    PORT
      LAYER metal1 ;
        RECT 9.400 6.800 9.800 7.600 ;
      LAYER metal2 ;
        RECT 9.400 6.800 9.800 7.200 ;
        RECT 9.400 -1.900 9.700 6.800 ;
        RECT 11.000 -1.900 11.400 -1.800 ;
        RECT 9.400 -2.200 11.400 -1.900 ;
    END
  END datain[7]
  PIN address[0]
    PORT
      LAYER metal1 ;
        RECT 186.200 5.400 186.600 6.200 ;
      LAYER via1 ;
        RECT 186.200 5.800 186.600 6.200 ;
      LAYER metal2 ;
        RECT 186.200 5.800 186.600 6.200 ;
        RECT 185.400 -1.900 185.800 -1.800 ;
        RECT 186.200 -1.900 186.500 5.800 ;
        RECT 185.400 -2.200 186.500 -1.900 ;
    END
  END address[0]
  PIN address[1]
    PORT
      LAYER metal1 ;
        RECT 88.600 6.100 89.000 6.200 ;
        RECT 90.200 6.100 90.600 6.200 ;
        RECT 88.600 5.800 90.600 6.100 ;
        RECT 88.600 5.400 89.000 5.800 ;
      LAYER via1 ;
        RECT 90.200 5.800 90.600 6.200 ;
      LAYER metal2 ;
        RECT 90.200 5.800 90.600 6.200 ;
        RECT 90.200 -1.800 90.500 5.800 ;
        RECT 90.200 -2.200 90.600 -1.800 ;
    END
  END address[1]
  PIN address[2]
    PORT
      LAYER metal1 ;
        RECT 84.600 5.400 85.000 6.200 ;
      LAYER via1 ;
        RECT 84.600 5.800 85.000 6.200 ;
      LAYER metal2 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 84.600 -1.900 84.900 5.800 ;
        RECT 85.400 -1.900 85.800 -1.800 ;
        RECT 84.600 -2.200 85.800 -1.900 ;
    END
  END address[2]
  PIN address[3]
    PORT
      LAYER metal1 ;
        RECT 191.800 6.100 192.200 6.200 ;
        RECT 192.600 6.100 193.000 6.200 ;
        RECT 191.800 5.800 193.000 6.100 ;
        RECT 191.800 5.400 192.200 5.800 ;
      LAYER via1 ;
        RECT 192.600 5.800 193.000 6.200 ;
      LAYER metal2 ;
        RECT 192.600 5.800 193.000 6.200 ;
        RECT 192.600 -1.900 192.900 5.800 ;
        RECT 193.400 -1.900 193.800 -1.800 ;
        RECT 192.600 -2.200 193.800 -1.900 ;
    END
  END address[3]
  PIN address[4]
    PORT
      LAYER metal1 ;
        RECT 199.000 5.400 199.400 6.200 ;
      LAYER via1 ;
        RECT 199.000 5.800 199.400 6.200 ;
      LAYER metal2 ;
        RECT 199.000 5.800 199.400 6.200 ;
        RECT 198.200 -1.900 198.600 -1.800 ;
        RECT 199.000 -1.900 199.300 5.800 ;
        RECT 198.200 -2.200 199.300 -1.900 ;
    END
  END address[4]
  PIN dataout[0]
    PORT
      LAYER metal1 ;
        RECT 172.600 75.900 173.000 79.900 ;
        RECT 172.700 74.800 173.000 75.900 ;
        RECT 172.600 71.100 173.000 74.800 ;
      LAYER via1 ;
        RECT 172.600 76.800 173.000 77.200 ;
      LAYER metal2 ;
        RECT 172.600 77.100 173.000 77.200 ;
        RECT 173.400 77.100 173.800 77.200 ;
        RECT 172.600 76.800 173.800 77.100 ;
      LAYER via2 ;
        RECT 173.400 76.800 173.800 77.200 ;
      LAYER metal3 ;
        RECT 173.400 77.100 173.800 77.200 ;
        RECT 176.600 77.100 177.000 77.200 ;
        RECT 172.600 76.800 177.000 77.100 ;
        RECT 230.200 77.100 230.600 77.200 ;
        RECT 233.400 77.100 233.800 77.200 ;
        RECT 230.200 76.800 233.800 77.100 ;
      LAYER via3 ;
        RECT 176.600 76.800 177.000 77.200 ;
      LAYER metal4 ;
        RECT 176.600 77.100 177.000 77.200 ;
        RECT 177.400 77.100 177.800 77.200 ;
        RECT 176.600 76.800 177.800 77.100 ;
        RECT 229.400 77.100 229.800 77.200 ;
        RECT 230.200 77.100 230.600 77.200 ;
        RECT 229.400 76.800 230.600 77.100 ;
      LAYER via4 ;
        RECT 177.400 76.800 177.800 77.200 ;
      LAYER metal5 ;
        RECT 177.400 77.100 177.800 77.200 ;
        RECT 229.400 77.100 229.800 77.200 ;
        RECT 177.400 76.800 229.800 77.100 ;
    END
  END dataout[0]
  PIN dataout[1]
    PORT
      LAYER metal1 ;
        RECT 230.200 126.200 230.600 129.900 ;
        RECT 230.300 125.100 230.600 126.200 ;
        RECT 230.200 121.100 230.600 125.100 ;
      LAYER via1 ;
        RECT 230.200 123.800 230.600 124.200 ;
      LAYER metal2 ;
        RECT 230.200 124.800 230.600 125.200 ;
        RECT 230.200 124.200 230.500 124.800 ;
        RECT 230.200 123.800 230.600 124.200 ;
      LAYER metal3 ;
        RECT 230.200 125.100 230.600 125.200 ;
        RECT 233.400 125.100 233.800 125.200 ;
        RECT 230.200 124.800 233.800 125.100 ;
    END
  END dataout[1]
  PIN dataout[2]
    PORT
      LAYER metal1 ;
        RECT 230.200 75.900 230.600 79.900 ;
        RECT 230.300 74.800 230.600 75.900 ;
        RECT 230.200 71.100 230.600 74.800 ;
      LAYER via1 ;
        RECT 230.200 73.800 230.600 74.200 ;
      LAYER metal2 ;
        RECT 230.200 74.800 230.600 75.200 ;
        RECT 230.200 74.200 230.500 74.800 ;
        RECT 230.200 73.800 230.600 74.200 ;
      LAYER metal3 ;
        RECT 230.200 75.100 230.600 75.200 ;
        RECT 233.400 75.100 233.800 75.200 ;
        RECT 230.200 74.800 233.800 75.100 ;
    END
  END dataout[2]
  PIN dataout[3]
    PORT
      LAYER metal1 ;
        RECT 173.400 86.200 173.800 89.900 ;
        RECT 173.500 85.100 173.800 86.200 ;
        RECT 173.400 81.100 173.800 85.100 ;
      LAYER via1 ;
        RECT 173.400 83.800 173.800 84.200 ;
      LAYER metal2 ;
        RECT 172.600 84.100 173.000 84.200 ;
        RECT 173.400 84.100 173.800 84.200 ;
        RECT 172.600 83.800 173.800 84.100 ;
      LAYER metal3 ;
        RECT 230.200 85.100 230.600 85.200 ;
        RECT 233.400 85.100 233.800 85.200 ;
        RECT 230.200 84.800 233.800 85.100 ;
        RECT 172.600 84.100 173.000 84.200 ;
        RECT 175.800 84.100 176.200 84.200 ;
        RECT 172.600 83.800 176.200 84.100 ;
      LAYER via3 ;
        RECT 175.800 83.800 176.200 84.200 ;
      LAYER metal4 ;
        RECT 175.800 84.800 176.200 85.200 ;
        RECT 229.400 85.100 229.800 85.200 ;
        RECT 230.200 85.100 230.600 85.200 ;
        RECT 229.400 84.800 230.600 85.100 ;
        RECT 175.800 84.200 176.100 84.800 ;
        RECT 175.800 83.800 176.200 84.200 ;
      LAYER metal5 ;
        RECT 175.800 85.100 176.200 85.200 ;
        RECT 229.400 85.100 229.800 85.200 ;
        RECT 175.800 84.800 229.800 85.100 ;
    END
  END dataout[3]
  PIN dataout[4]
    PORT
      LAYER metal1 ;
        RECT 226.200 95.900 226.600 99.900 ;
        RECT 226.300 94.800 226.600 95.900 ;
        RECT 226.200 91.100 226.600 94.800 ;
      LAYER via1 ;
        RECT 226.200 93.800 226.600 94.200 ;
      LAYER metal2 ;
        RECT 226.200 94.800 226.600 95.200 ;
        RECT 226.200 94.200 226.500 94.800 ;
        RECT 226.200 93.800 226.600 94.200 ;
      LAYER metal3 ;
        RECT 226.200 95.100 226.600 95.200 ;
        RECT 233.400 95.100 233.800 95.200 ;
        RECT 226.200 94.800 233.800 95.100 ;
    END
  END dataout[4]
  PIN dataout[5]
    PORT
      LAYER metal1 ;
        RECT 228.600 97.100 229.000 99.900 ;
        RECT 229.400 97.100 229.800 97.200 ;
        RECT 228.600 96.800 229.800 97.100 ;
        RECT 228.600 95.900 229.000 96.800 ;
        RECT 228.700 94.800 229.000 95.900 ;
        RECT 228.600 91.100 229.000 94.800 ;
      LAYER via1 ;
        RECT 229.400 96.800 229.800 97.200 ;
      LAYER metal2 ;
        RECT 229.400 97.100 229.800 97.200 ;
        RECT 230.200 97.100 230.600 97.200 ;
        RECT 229.400 96.800 230.600 97.100 ;
      LAYER via2 ;
        RECT 230.200 96.800 230.600 97.200 ;
      LAYER metal3 ;
        RECT 230.200 97.100 230.600 97.200 ;
        RECT 233.400 97.100 233.800 97.200 ;
        RECT 230.200 96.800 233.800 97.100 ;
    END
  END dataout[5]
  PIN dataout[6]
    PORT
      LAYER metal1 ;
        RECT 229.400 135.900 229.800 139.900 ;
        RECT 229.500 134.800 229.800 135.900 ;
        RECT 229.400 134.100 229.800 134.800 ;
        RECT 230.200 134.100 230.600 134.200 ;
        RECT 229.400 133.800 230.600 134.100 ;
        RECT 229.400 131.100 229.800 133.800 ;
      LAYER via1 ;
        RECT 230.200 133.800 230.600 134.200 ;
      LAYER metal2 ;
        RECT 230.200 134.800 230.600 135.200 ;
        RECT 230.200 134.200 230.500 134.800 ;
        RECT 230.200 133.800 230.600 134.200 ;
      LAYER metal3 ;
        RECT 230.200 135.100 230.600 135.200 ;
        RECT 233.400 135.100 233.800 135.200 ;
        RECT 230.200 134.800 233.800 135.100 ;
    END
  END dataout[6]
  PIN dataout[7]
    PORT
      LAYER metal1 ;
        RECT 162.200 46.200 162.600 49.900 ;
        RECT 162.300 45.100 162.600 46.200 ;
        RECT 162.200 41.100 162.600 45.100 ;
      LAYER via1 ;
        RECT 162.200 41.800 162.600 42.200 ;
      LAYER metal2 ;
        RECT 162.200 41.800 162.600 42.200 ;
        RECT 162.200 38.200 162.500 41.800 ;
        RECT 162.200 37.800 162.600 38.200 ;
        RECT 161.400 0.800 161.800 1.200 ;
        RECT 161.400 -1.800 161.700 0.800 ;
        RECT 161.400 -2.200 161.800 -1.800 ;
      LAYER metal3 ;
        RECT 162.200 37.800 162.600 38.200 ;
        RECT 162.200 37.200 162.500 37.800 ;
        RECT 162.200 36.800 162.600 37.200 ;
        RECT 161.400 1.100 161.800 1.200 ;
        RECT 162.200 1.100 162.600 1.200 ;
        RECT 161.400 0.800 162.600 1.100 ;
      LAYER via3 ;
        RECT 162.200 0.800 162.600 1.200 ;
      LAYER metal4 ;
        RECT 162.200 36.800 162.600 37.200 ;
        RECT 162.200 1.200 162.500 36.800 ;
        RECT 162.200 0.800 162.600 1.200 ;
    END
  END dataout[7]
  OBS
      LAYER metal1 ;
        RECT 1.400 207.600 1.800 209.900 ;
        RECT 3.000 207.600 3.400 209.900 ;
        RECT 4.600 207.600 5.000 209.900 ;
        RECT 6.200 207.600 6.600 209.900 ;
        RECT 8.600 207.600 9.000 209.900 ;
        RECT 10.200 207.600 10.600 209.900 ;
        RECT 11.800 207.600 12.200 209.900 ;
        RECT 13.400 207.600 13.800 209.900 ;
        RECT 1.400 207.200 2.300 207.600 ;
        RECT 3.000 207.200 4.100 207.600 ;
        RECT 4.600 207.200 5.700 207.600 ;
        RECT 6.200 207.200 7.400 207.600 ;
        RECT 8.600 207.200 9.500 207.600 ;
        RECT 10.200 207.200 11.300 207.600 ;
        RECT 11.800 207.200 12.900 207.600 ;
        RECT 13.400 207.200 14.600 207.600 ;
        RECT 15.000 207.500 15.400 209.900 ;
        RECT 17.200 209.200 17.600 209.900 ;
        RECT 16.600 208.900 17.600 209.200 ;
        RECT 19.400 208.900 19.800 209.900 ;
        RECT 21.500 209.200 22.100 209.900 ;
        RECT 21.400 208.900 22.100 209.200 ;
        RECT 16.600 208.500 17.000 208.900 ;
        RECT 19.400 208.600 19.700 208.900 ;
        RECT 17.400 208.200 17.800 208.600 ;
        RECT 18.300 208.300 19.700 208.600 ;
        RECT 21.400 208.500 21.800 208.900 ;
        RECT 18.300 208.200 18.700 208.300 ;
        RECT 1.900 206.900 2.300 207.200 ;
        RECT 3.700 206.900 4.100 207.200 ;
        RECT 5.300 206.900 5.700 207.200 ;
        RECT 1.900 206.500 3.200 206.900 ;
        RECT 3.700 206.500 4.900 206.900 ;
        RECT 5.300 206.500 6.600 206.900 ;
        RECT 1.900 205.800 2.300 206.500 ;
        RECT 3.700 205.800 4.100 206.500 ;
        RECT 5.300 205.800 5.700 206.500 ;
        RECT 7.000 205.800 7.400 207.200 ;
        RECT 9.100 206.900 9.500 207.200 ;
        RECT 10.900 206.900 11.300 207.200 ;
        RECT 12.500 206.900 12.900 207.200 ;
        RECT 9.100 206.500 10.400 206.900 ;
        RECT 10.900 206.500 12.100 206.900 ;
        RECT 12.500 206.500 13.800 206.900 ;
        RECT 9.100 205.800 9.500 206.500 ;
        RECT 10.900 205.800 11.300 206.500 ;
        RECT 12.500 205.800 12.900 206.500 ;
        RECT 14.200 205.800 14.600 207.200 ;
        RECT 15.400 207.100 16.200 207.200 ;
        RECT 17.500 207.100 17.800 208.200 ;
        RECT 22.300 207.700 22.700 207.800 ;
        RECT 23.800 207.700 24.200 209.900 ;
        RECT 24.600 208.000 25.000 209.900 ;
        RECT 26.200 208.000 26.600 209.900 ;
        RECT 24.600 207.900 26.600 208.000 ;
        RECT 27.000 207.900 27.400 209.900 ;
        RECT 27.800 207.900 28.200 209.900 ;
        RECT 28.600 208.000 29.000 209.900 ;
        RECT 30.200 208.000 30.600 209.900 ;
        RECT 28.600 207.900 30.600 208.000 ;
        RECT 24.700 207.700 26.500 207.900 ;
        RECT 22.300 207.400 24.200 207.700 ;
        RECT 20.300 207.100 20.700 207.200 ;
        RECT 15.400 206.800 20.900 207.100 ;
        RECT 16.900 206.700 17.300 206.800 ;
        RECT 16.100 206.200 16.500 206.300 ;
        RECT 16.100 205.900 18.600 206.200 ;
        RECT 18.200 205.800 18.600 205.900 ;
        RECT 1.400 205.400 2.300 205.800 ;
        RECT 3.000 205.400 4.100 205.800 ;
        RECT 4.600 205.400 5.700 205.800 ;
        RECT 6.200 205.400 7.400 205.800 ;
        RECT 8.600 205.400 9.500 205.800 ;
        RECT 10.200 205.400 11.300 205.800 ;
        RECT 11.800 205.400 12.900 205.800 ;
        RECT 13.400 205.400 14.600 205.800 ;
        RECT 15.000 205.500 17.800 205.600 ;
        RECT 15.000 205.400 17.900 205.500 ;
        RECT 1.400 201.100 1.800 205.400 ;
        RECT 3.000 201.100 3.400 205.400 ;
        RECT 4.600 201.100 5.000 205.400 ;
        RECT 6.200 201.100 6.600 205.400 ;
        RECT 8.600 201.100 9.000 205.400 ;
        RECT 10.200 201.100 10.600 205.400 ;
        RECT 11.800 201.100 12.200 205.400 ;
        RECT 13.400 201.100 13.800 205.400 ;
        RECT 15.000 205.300 19.900 205.400 ;
        RECT 15.000 201.100 15.400 205.300 ;
        RECT 17.500 205.100 19.900 205.300 ;
        RECT 16.600 204.500 19.300 204.800 ;
        RECT 16.600 204.400 17.000 204.500 ;
        RECT 18.900 204.400 19.300 204.500 ;
        RECT 19.600 204.500 19.900 205.100 ;
        RECT 20.600 205.200 20.900 206.800 ;
        RECT 21.400 206.400 21.800 206.500 ;
        RECT 21.400 206.100 23.300 206.400 ;
        RECT 22.900 206.000 23.300 206.100 ;
        RECT 22.100 205.700 22.500 205.800 ;
        RECT 23.800 205.700 24.200 207.400 ;
        RECT 25.000 207.200 25.400 207.400 ;
        RECT 27.000 207.200 27.300 207.900 ;
        RECT 27.900 207.200 28.200 207.900 ;
        RECT 28.700 207.700 30.500 207.900 ;
        RECT 31.000 207.500 31.400 209.900 ;
        RECT 33.200 209.200 33.600 209.900 ;
        RECT 32.600 208.900 33.600 209.200 ;
        RECT 35.400 208.900 35.800 209.900 ;
        RECT 37.500 209.200 38.100 209.900 ;
        RECT 37.400 208.900 38.100 209.200 ;
        RECT 32.600 208.500 33.000 208.900 ;
        RECT 35.400 208.600 35.700 208.900 ;
        RECT 33.400 208.200 33.800 208.600 ;
        RECT 34.300 208.300 35.700 208.600 ;
        RECT 37.400 208.500 37.800 208.900 ;
        RECT 34.300 208.200 34.700 208.300 ;
        RECT 29.800 207.200 30.200 207.400 ;
        RECT 24.600 206.900 25.400 207.200 ;
        RECT 24.600 206.800 25.000 206.900 ;
        RECT 26.100 206.800 27.400 207.200 ;
        RECT 27.800 206.800 29.100 207.200 ;
        RECT 29.800 206.900 30.600 207.200 ;
        RECT 30.200 206.800 30.600 206.900 ;
        RECT 31.400 207.100 32.200 207.200 ;
        RECT 33.500 207.100 33.800 208.200 ;
        RECT 38.300 207.700 38.700 207.800 ;
        RECT 39.800 207.700 40.200 209.900 ;
        RECT 43.000 208.200 43.400 209.900 ;
        RECT 38.300 207.400 40.200 207.700 ;
        RECT 35.000 207.100 35.400 207.200 ;
        RECT 36.300 207.100 36.700 207.200 ;
        RECT 31.400 206.800 36.900 207.100 ;
        RECT 25.400 205.800 25.800 206.600 ;
        RECT 26.100 206.100 26.400 206.800 ;
        RECT 28.800 206.200 29.100 206.800 ;
        RECT 32.900 206.700 33.300 206.800 ;
        RECT 26.100 205.800 28.100 206.100 ;
        RECT 28.600 205.800 29.100 206.200 ;
        RECT 29.400 205.800 29.800 206.600 ;
        RECT 32.100 206.200 32.500 206.300 ;
        RECT 33.400 206.200 33.800 206.300 ;
        RECT 32.100 205.900 34.600 206.200 ;
        RECT 34.200 205.800 34.600 205.900 ;
        RECT 22.100 205.400 24.200 205.700 ;
        RECT 20.600 204.900 21.800 205.200 ;
        RECT 20.300 204.500 20.700 204.600 ;
        RECT 19.600 204.200 20.700 204.500 ;
        RECT 21.500 204.400 21.800 204.900 ;
        RECT 21.500 204.000 22.200 204.400 ;
        RECT 18.300 203.700 18.700 203.800 ;
        RECT 19.700 203.700 20.100 203.800 ;
        RECT 16.600 203.100 17.000 203.500 ;
        RECT 18.300 203.400 20.100 203.700 ;
        RECT 19.400 203.100 19.700 203.400 ;
        RECT 21.400 203.100 21.800 203.500 ;
        RECT 16.600 202.800 17.600 203.100 ;
        RECT 17.200 201.100 17.600 202.800 ;
        RECT 19.400 201.100 19.800 203.100 ;
        RECT 21.500 201.100 22.100 203.100 ;
        RECT 23.800 201.100 24.200 205.400 ;
        RECT 26.100 205.100 26.400 205.800 ;
        RECT 27.800 205.200 28.100 205.800 ;
        RECT 27.000 205.100 27.400 205.200 ;
        RECT 25.900 204.800 26.400 205.100 ;
        RECT 26.700 204.800 27.400 205.100 ;
        RECT 27.800 205.100 28.200 205.200 ;
        RECT 28.800 205.100 29.100 205.800 ;
        RECT 31.000 205.500 33.800 205.600 ;
        RECT 31.000 205.400 33.900 205.500 ;
        RECT 31.000 205.300 35.900 205.400 ;
        RECT 27.800 204.800 28.500 205.100 ;
        RECT 28.800 204.800 29.300 205.100 ;
        RECT 25.900 201.100 26.300 204.800 ;
        RECT 26.700 204.200 27.000 204.800 ;
        RECT 28.200 204.200 28.500 204.800 ;
        RECT 26.600 203.800 27.400 204.200 ;
        RECT 28.200 203.800 28.600 204.200 ;
        RECT 28.900 201.100 29.300 204.800 ;
        RECT 31.000 201.100 31.400 205.300 ;
        RECT 33.500 205.100 35.900 205.300 ;
        RECT 32.600 204.500 35.300 204.800 ;
        RECT 32.600 204.400 33.000 204.500 ;
        RECT 34.900 204.400 35.300 204.500 ;
        RECT 35.600 204.500 35.900 205.100 ;
        RECT 36.600 205.200 36.900 206.800 ;
        RECT 37.400 206.400 37.800 206.500 ;
        RECT 37.400 206.100 39.300 206.400 ;
        RECT 38.900 206.000 39.300 206.100 ;
        RECT 38.100 205.700 38.500 205.800 ;
        RECT 39.800 205.700 40.200 207.400 ;
        RECT 38.100 205.400 40.200 205.700 ;
        RECT 36.600 204.900 37.800 205.200 ;
        RECT 36.300 204.500 36.700 204.600 ;
        RECT 35.600 204.200 36.700 204.500 ;
        RECT 37.500 204.400 37.800 204.900 ;
        RECT 37.500 204.000 38.200 204.400 ;
        RECT 34.300 203.700 34.700 203.800 ;
        RECT 35.700 203.700 36.100 203.800 ;
        RECT 32.600 203.100 33.000 203.500 ;
        RECT 34.300 203.400 36.100 203.700 ;
        RECT 35.400 203.100 35.700 203.400 ;
        RECT 37.400 203.100 37.800 203.500 ;
        RECT 32.600 202.800 33.600 203.100 ;
        RECT 33.200 201.100 33.600 202.800 ;
        RECT 35.400 201.100 35.800 203.100 ;
        RECT 37.500 201.100 38.100 203.100 ;
        RECT 39.800 201.100 40.200 205.400 ;
        RECT 42.900 207.900 43.400 208.200 ;
        RECT 42.900 207.200 43.200 207.900 ;
        RECT 44.600 207.600 45.000 209.900 ;
        RECT 43.700 207.300 45.000 207.600 ;
        RECT 45.400 207.500 45.800 209.900 ;
        RECT 47.600 209.200 48.000 209.900 ;
        RECT 47.000 208.900 48.000 209.200 ;
        RECT 49.800 208.900 50.200 209.900 ;
        RECT 51.900 209.200 52.500 209.900 ;
        RECT 51.800 208.900 52.500 209.200 ;
        RECT 47.000 208.500 47.400 208.900 ;
        RECT 49.800 208.600 50.100 208.900 ;
        RECT 47.800 208.200 48.200 208.600 ;
        RECT 48.700 208.300 50.100 208.600 ;
        RECT 51.800 208.500 52.200 208.900 ;
        RECT 48.700 208.200 49.100 208.300 ;
        RECT 42.900 206.800 43.400 207.200 ;
        RECT 42.900 205.100 43.200 206.800 ;
        RECT 43.700 206.500 44.000 207.300 ;
        RECT 45.800 207.100 46.600 207.200 ;
        RECT 47.900 207.100 48.200 208.200 ;
        RECT 52.700 207.700 53.100 207.800 ;
        RECT 54.200 207.700 54.600 209.900 ;
        RECT 55.000 208.000 55.400 209.900 ;
        RECT 56.600 208.000 57.000 209.900 ;
        RECT 55.000 207.900 57.000 208.000 ;
        RECT 57.400 207.900 57.800 209.900 ;
        RECT 58.200 207.900 58.600 209.900 ;
        RECT 59.000 208.000 59.400 209.900 ;
        RECT 60.600 208.000 61.000 209.900 ;
        RECT 62.200 208.200 62.600 209.900 ;
        RECT 59.000 207.900 61.000 208.000 ;
        RECT 62.100 207.900 62.600 208.200 ;
        RECT 55.100 207.700 56.900 207.900 ;
        RECT 52.700 207.400 54.600 207.700 ;
        RECT 50.700 207.100 51.100 207.200 ;
        RECT 45.800 206.800 51.300 207.100 ;
        RECT 47.300 206.700 47.700 206.800 ;
        RECT 43.500 206.100 44.000 206.500 ;
        RECT 43.700 205.100 44.000 206.100 ;
        RECT 44.500 206.200 44.900 206.600 ;
        RECT 46.500 206.200 46.900 206.300 ;
        RECT 44.500 205.800 45.000 206.200 ;
        RECT 46.500 205.900 49.000 206.200 ;
        RECT 48.600 205.800 49.000 205.900 ;
        RECT 45.400 205.500 48.200 205.600 ;
        RECT 45.400 205.400 48.300 205.500 ;
        RECT 45.400 205.300 50.300 205.400 ;
        RECT 42.900 204.600 43.400 205.100 ;
        RECT 43.700 204.800 45.000 205.100 ;
        RECT 43.000 201.100 43.400 204.600 ;
        RECT 44.600 201.100 45.000 204.800 ;
        RECT 45.400 201.100 45.800 205.300 ;
        RECT 47.900 205.100 50.300 205.300 ;
        RECT 47.000 204.500 49.700 204.800 ;
        RECT 47.000 204.400 47.400 204.500 ;
        RECT 49.300 204.400 49.700 204.500 ;
        RECT 50.000 204.500 50.300 205.100 ;
        RECT 51.000 205.200 51.300 206.800 ;
        RECT 51.800 206.400 52.200 206.500 ;
        RECT 51.800 206.100 53.700 206.400 ;
        RECT 53.300 206.000 53.700 206.100 ;
        RECT 52.500 205.700 52.900 205.800 ;
        RECT 54.200 205.700 54.600 207.400 ;
        RECT 55.400 207.200 55.800 207.400 ;
        RECT 57.400 207.200 57.700 207.900 ;
        RECT 58.300 207.200 58.600 207.900 ;
        RECT 59.100 207.700 60.900 207.900 ;
        RECT 60.200 207.200 60.600 207.400 ;
        RECT 62.100 207.200 62.400 207.900 ;
        RECT 63.800 207.600 64.200 209.900 ;
        RECT 62.900 207.300 64.200 207.600 ;
        RECT 64.600 207.500 65.000 209.900 ;
        RECT 66.800 209.200 67.200 209.900 ;
        RECT 66.200 208.900 67.200 209.200 ;
        RECT 69.000 208.900 69.400 209.900 ;
        RECT 71.100 209.200 71.700 209.900 ;
        RECT 71.000 208.900 71.700 209.200 ;
        RECT 66.200 208.500 66.600 208.900 ;
        RECT 69.000 208.600 69.300 208.900 ;
        RECT 67.000 208.200 67.400 208.600 ;
        RECT 67.900 208.300 69.300 208.600 ;
        RECT 71.000 208.500 71.400 208.900 ;
        RECT 67.900 208.200 68.300 208.300 ;
        RECT 55.000 206.900 55.800 207.200 ;
        RECT 55.000 206.800 55.400 206.900 ;
        RECT 56.500 206.800 57.800 207.200 ;
        RECT 58.200 206.800 59.500 207.200 ;
        RECT 60.200 206.900 61.000 207.200 ;
        RECT 62.100 207.100 62.600 207.200 ;
        RECT 60.600 206.800 61.000 206.900 ;
        RECT 61.400 206.800 62.600 207.100 ;
        RECT 55.800 205.800 56.200 206.600 ;
        RECT 52.500 205.400 54.600 205.700 ;
        RECT 51.000 204.900 52.200 205.200 ;
        RECT 50.700 204.500 51.100 204.600 ;
        RECT 50.000 204.200 51.100 204.500 ;
        RECT 51.900 204.400 52.200 204.900 ;
        RECT 51.900 204.000 52.600 204.400 ;
        RECT 48.700 203.700 49.100 203.800 ;
        RECT 50.100 203.700 50.500 203.800 ;
        RECT 47.000 203.100 47.400 203.500 ;
        RECT 48.700 203.400 50.500 203.700 ;
        RECT 49.800 203.100 50.100 203.400 ;
        RECT 51.800 203.100 52.200 203.500 ;
        RECT 47.000 202.800 48.000 203.100 ;
        RECT 47.600 201.100 48.000 202.800 ;
        RECT 49.800 201.100 50.200 203.100 ;
        RECT 51.900 201.100 52.500 203.100 ;
        RECT 54.200 201.100 54.600 205.400 ;
        RECT 56.500 205.100 56.800 206.800 ;
        RECT 59.200 206.100 59.500 206.800 ;
        RECT 57.400 205.800 59.500 206.100 ;
        RECT 59.800 206.100 60.200 206.600 ;
        RECT 61.400 206.100 61.700 206.800 ;
        RECT 59.800 205.800 61.700 206.100 ;
        RECT 57.400 205.200 57.700 205.800 ;
        RECT 57.400 205.100 57.800 205.200 ;
        RECT 56.300 204.800 56.800 205.100 ;
        RECT 57.100 204.800 57.800 205.100 ;
        RECT 58.200 205.100 58.600 205.200 ;
        RECT 59.200 205.100 59.500 205.800 ;
        RECT 62.100 205.100 62.400 206.800 ;
        RECT 62.900 206.500 63.200 207.300 ;
        RECT 67.100 207.200 67.400 208.200 ;
        RECT 71.900 207.700 72.300 207.800 ;
        RECT 73.400 207.700 73.800 209.900 ;
        RECT 71.900 207.400 73.800 207.700 ;
        RECT 65.000 207.100 65.800 207.200 ;
        RECT 67.000 207.100 67.400 207.200 ;
        RECT 69.900 207.100 70.300 207.200 ;
        RECT 65.000 206.800 70.500 207.100 ;
        RECT 66.500 206.700 66.900 206.800 ;
        RECT 62.700 206.100 63.200 206.500 ;
        RECT 62.900 205.100 63.200 206.100 ;
        RECT 63.700 206.200 64.100 206.600 ;
        RECT 65.700 206.200 66.100 206.300 ;
        RECT 63.700 205.800 64.200 206.200 ;
        RECT 65.700 205.900 68.200 206.200 ;
        RECT 67.800 205.800 68.200 205.900 ;
        RECT 64.600 205.500 67.400 205.600 ;
        RECT 64.600 205.400 67.500 205.500 ;
        RECT 64.600 205.300 69.500 205.400 ;
        RECT 58.200 204.800 58.900 205.100 ;
        RECT 59.200 204.800 59.700 205.100 ;
        RECT 56.300 201.100 56.700 204.800 ;
        RECT 57.100 204.200 57.400 204.800 ;
        RECT 58.600 204.200 58.900 204.800 ;
        RECT 57.000 203.800 57.400 204.200 ;
        RECT 58.200 203.800 59.000 204.200 ;
        RECT 59.300 201.100 59.700 204.800 ;
        RECT 62.100 204.600 62.600 205.100 ;
        RECT 62.900 204.800 64.200 205.100 ;
        RECT 62.200 201.100 62.600 204.600 ;
        RECT 63.800 201.100 64.200 204.800 ;
        RECT 64.600 201.100 65.000 205.300 ;
        RECT 67.100 205.100 69.500 205.300 ;
        RECT 66.200 204.500 68.900 204.800 ;
        RECT 66.200 204.400 66.600 204.500 ;
        RECT 68.500 204.400 68.900 204.500 ;
        RECT 69.200 204.500 69.500 205.100 ;
        RECT 70.200 205.200 70.500 206.800 ;
        RECT 71.000 206.400 71.400 206.500 ;
        RECT 71.000 206.100 72.900 206.400 ;
        RECT 72.500 206.000 72.900 206.100 ;
        RECT 71.700 205.700 72.100 205.800 ;
        RECT 73.400 205.700 73.800 207.400 ;
        RECT 71.700 205.400 73.800 205.700 ;
        RECT 70.200 204.900 71.400 205.200 ;
        RECT 69.900 204.500 70.300 204.600 ;
        RECT 69.200 204.200 70.300 204.500 ;
        RECT 71.100 204.400 71.400 204.900 ;
        RECT 71.100 204.000 71.800 204.400 ;
        RECT 67.900 203.700 68.300 203.800 ;
        RECT 69.300 203.700 69.700 203.800 ;
        RECT 66.200 203.100 66.600 203.500 ;
        RECT 67.900 203.400 69.700 203.700 ;
        RECT 69.000 203.100 69.300 203.400 ;
        RECT 71.000 203.100 71.400 203.500 ;
        RECT 66.200 202.800 67.200 203.100 ;
        RECT 66.800 201.100 67.200 202.800 ;
        RECT 69.000 201.100 69.400 203.100 ;
        RECT 71.100 201.100 71.700 203.100 ;
        RECT 73.400 201.100 73.800 205.400 ;
        RECT 74.200 207.700 74.600 209.900 ;
        RECT 76.300 209.200 76.900 209.900 ;
        RECT 76.300 208.900 77.000 209.200 ;
        RECT 78.600 208.900 79.000 209.900 ;
        RECT 80.800 209.200 81.200 209.900 ;
        RECT 80.800 208.900 81.800 209.200 ;
        RECT 76.600 208.500 77.000 208.900 ;
        RECT 78.700 208.600 79.000 208.900 ;
        RECT 78.700 208.300 80.100 208.600 ;
        RECT 79.700 208.200 80.100 208.300 ;
        RECT 80.600 208.200 81.000 208.600 ;
        RECT 81.400 208.500 81.800 208.900 ;
        RECT 75.700 207.700 76.100 207.800 ;
        RECT 74.200 207.400 76.100 207.700 ;
        RECT 74.200 205.700 74.600 207.400 ;
        RECT 77.700 207.100 78.100 207.200 ;
        RECT 80.600 207.100 80.900 208.200 ;
        RECT 83.000 207.500 83.400 209.900 ;
        RECT 83.800 208.000 84.200 209.900 ;
        RECT 85.400 208.000 85.800 209.900 ;
        RECT 83.800 207.900 85.800 208.000 ;
        RECT 86.200 207.900 86.600 209.900 ;
        RECT 87.000 207.900 87.400 209.900 ;
        RECT 87.800 208.000 88.200 209.900 ;
        RECT 89.400 208.000 89.800 209.900 ;
        RECT 87.800 207.900 89.800 208.000 ;
        RECT 83.900 207.700 85.700 207.900 ;
        RECT 84.200 207.200 84.600 207.400 ;
        RECT 86.200 207.200 86.500 207.900 ;
        RECT 87.100 207.200 87.400 207.900 ;
        RECT 87.900 207.700 89.700 207.900 ;
        RECT 91.800 207.500 92.200 209.900 ;
        RECT 94.000 209.200 94.400 209.900 ;
        RECT 93.400 208.900 94.400 209.200 ;
        RECT 96.200 208.900 96.600 209.900 ;
        RECT 98.300 209.200 98.900 209.900 ;
        RECT 98.200 208.900 98.900 209.200 ;
        RECT 93.400 208.500 93.800 208.900 ;
        RECT 96.200 208.600 96.500 208.900 ;
        RECT 94.200 208.200 94.600 208.600 ;
        RECT 95.100 208.300 96.500 208.600 ;
        RECT 98.200 208.500 98.600 208.900 ;
        RECT 95.100 208.200 95.500 208.300 ;
        RECT 89.000 207.200 89.400 207.400 ;
        RECT 82.200 207.100 83.000 207.200 ;
        RECT 77.500 206.800 83.000 207.100 ;
        RECT 83.800 206.900 84.600 207.200 ;
        RECT 83.800 206.800 84.200 206.900 ;
        RECT 85.300 206.800 86.600 207.200 ;
        RECT 87.000 206.800 88.300 207.200 ;
        RECT 89.000 206.900 89.800 207.200 ;
        RECT 89.400 206.800 89.800 206.900 ;
        RECT 92.200 207.100 93.000 207.200 ;
        RECT 94.300 207.100 94.600 208.200 ;
        RECT 99.100 207.700 99.500 207.800 ;
        RECT 100.600 207.700 101.000 209.900 ;
        RECT 99.100 207.400 101.000 207.700 ;
        RECT 101.400 207.500 101.800 209.900 ;
        RECT 103.600 209.200 104.000 209.900 ;
        RECT 103.000 208.900 104.000 209.200 ;
        RECT 105.800 208.900 106.200 209.900 ;
        RECT 107.900 209.200 108.500 209.900 ;
        RECT 107.800 208.900 108.500 209.200 ;
        RECT 103.000 208.500 103.400 208.900 ;
        RECT 105.800 208.600 106.100 208.900 ;
        RECT 103.800 208.200 104.200 208.600 ;
        RECT 104.700 208.300 106.100 208.600 ;
        RECT 107.800 208.500 108.200 208.900 ;
        RECT 104.700 208.200 105.100 208.300 ;
        RECT 97.100 207.100 97.500 207.200 ;
        RECT 92.200 206.800 97.700 207.100 ;
        RECT 76.600 206.400 77.000 206.500 ;
        RECT 75.100 206.100 77.000 206.400 ;
        RECT 77.500 206.200 77.800 206.800 ;
        RECT 81.100 206.700 81.500 206.800 ;
        RECT 80.600 206.200 81.000 206.300 ;
        RECT 81.900 206.200 82.300 206.300 ;
        RECT 75.100 206.000 75.500 206.100 ;
        RECT 77.400 205.800 77.800 206.200 ;
        RECT 79.800 205.900 82.300 206.200 ;
        RECT 79.800 205.800 80.200 205.900 ;
        RECT 84.600 205.800 85.000 206.600 ;
        RECT 85.300 206.100 85.600 206.800 ;
        RECT 88.000 206.200 88.300 206.800 ;
        RECT 93.700 206.700 94.100 206.800 ;
        RECT 85.300 205.800 87.300 206.100 ;
        RECT 87.800 205.800 88.300 206.200 ;
        RECT 88.600 206.100 89.000 206.600 ;
        RECT 92.900 206.200 93.300 206.300 ;
        RECT 94.200 206.200 94.600 206.300 ;
        RECT 97.400 206.200 97.700 206.800 ;
        RECT 98.200 206.400 98.600 206.500 ;
        RECT 90.200 206.100 90.600 206.200 ;
        RECT 88.600 205.800 90.600 206.100 ;
        RECT 92.900 205.900 95.400 206.200 ;
        RECT 95.000 205.800 95.400 205.900 ;
        RECT 97.400 205.800 97.800 206.200 ;
        RECT 98.200 206.100 100.100 206.400 ;
        RECT 99.700 206.000 100.100 206.100 ;
        RECT 75.900 205.700 76.300 205.800 ;
        RECT 74.200 205.400 76.300 205.700 ;
        RECT 74.200 201.100 74.600 205.400 ;
        RECT 77.500 205.200 77.800 205.800 ;
        RECT 80.600 205.500 83.400 205.600 ;
        RECT 80.500 205.400 83.400 205.500 ;
        RECT 76.600 204.900 77.800 205.200 ;
        RECT 78.500 205.300 83.400 205.400 ;
        RECT 78.500 205.100 80.900 205.300 ;
        RECT 76.600 204.400 76.900 204.900 ;
        RECT 76.200 204.000 76.900 204.400 ;
        RECT 77.700 204.500 78.100 204.600 ;
        RECT 78.500 204.500 78.800 205.100 ;
        RECT 77.700 204.200 78.800 204.500 ;
        RECT 79.100 204.500 81.800 204.800 ;
        RECT 79.100 204.400 79.500 204.500 ;
        RECT 81.400 204.400 81.800 204.500 ;
        RECT 78.300 203.700 78.700 203.800 ;
        RECT 79.700 203.700 80.100 203.800 ;
        RECT 76.600 203.100 77.000 203.500 ;
        RECT 78.300 203.400 80.100 203.700 ;
        RECT 78.700 203.100 79.000 203.400 ;
        RECT 81.400 203.100 81.800 203.500 ;
        RECT 76.300 201.100 76.900 203.100 ;
        RECT 78.600 201.100 79.000 203.100 ;
        RECT 80.800 202.800 81.800 203.100 ;
        RECT 80.800 201.100 81.200 202.800 ;
        RECT 83.000 201.100 83.400 205.300 ;
        RECT 85.300 205.100 85.600 205.800 ;
        RECT 87.000 205.200 87.300 205.800 ;
        RECT 86.200 205.100 86.600 205.200 ;
        RECT 85.100 204.800 85.600 205.100 ;
        RECT 85.900 204.800 86.600 205.100 ;
        RECT 87.000 205.100 87.400 205.200 ;
        RECT 88.000 205.100 88.300 205.800 ;
        RECT 91.800 205.500 94.600 205.600 ;
        RECT 91.800 205.400 94.700 205.500 ;
        RECT 91.800 205.300 96.700 205.400 ;
        RECT 87.000 204.800 87.700 205.100 ;
        RECT 88.000 204.800 88.500 205.100 ;
        RECT 85.100 201.100 85.500 204.800 ;
        RECT 85.900 204.200 86.200 204.800 ;
        RECT 87.400 204.200 87.700 204.800 ;
        RECT 85.800 203.800 86.600 204.200 ;
        RECT 87.400 203.800 87.800 204.200 ;
        RECT 88.100 201.100 88.500 204.800 ;
        RECT 91.800 201.100 92.200 205.300 ;
        RECT 94.300 205.100 96.700 205.300 ;
        RECT 93.400 204.500 96.100 204.800 ;
        RECT 93.400 204.400 93.800 204.500 ;
        RECT 95.700 204.400 96.100 204.500 ;
        RECT 96.400 204.500 96.700 205.100 ;
        RECT 97.400 205.200 97.700 205.800 ;
        RECT 98.900 205.700 99.300 205.800 ;
        RECT 100.600 205.700 101.000 207.400 ;
        RECT 101.800 207.100 102.600 207.200 ;
        RECT 103.900 207.100 104.200 208.200 ;
        RECT 108.700 207.700 109.100 207.800 ;
        RECT 110.200 207.700 110.600 209.900 ;
        RECT 111.000 208.000 111.400 209.900 ;
        RECT 112.600 208.000 113.000 209.900 ;
        RECT 111.000 207.900 113.000 208.000 ;
        RECT 113.400 207.900 113.800 209.900 ;
        RECT 114.200 207.900 114.600 209.900 ;
        RECT 115.000 208.000 115.400 209.900 ;
        RECT 116.600 208.000 117.000 209.900 ;
        RECT 115.000 207.900 117.000 208.000 ;
        RECT 117.400 208.000 117.800 209.900 ;
        RECT 119.000 208.000 119.400 209.900 ;
        RECT 117.400 207.900 119.400 208.000 ;
        RECT 119.800 207.900 120.200 209.900 ;
        RECT 120.600 208.000 121.000 209.900 ;
        RECT 122.200 208.000 122.600 209.900 ;
        RECT 120.600 207.900 122.600 208.000 ;
        RECT 123.000 207.900 123.400 209.900 ;
        RECT 111.100 207.700 112.900 207.900 ;
        RECT 108.700 207.400 110.600 207.700 ;
        RECT 106.700 207.100 107.100 207.200 ;
        RECT 101.800 206.800 107.300 207.100 ;
        RECT 103.300 206.700 103.700 206.800 ;
        RECT 102.500 206.200 102.900 206.300 ;
        RECT 102.500 205.900 105.000 206.200 ;
        RECT 104.600 205.800 105.000 205.900 ;
        RECT 98.900 205.400 101.000 205.700 ;
        RECT 97.400 204.900 98.600 205.200 ;
        RECT 97.100 204.500 97.500 204.600 ;
        RECT 96.400 204.200 97.500 204.500 ;
        RECT 98.300 204.400 98.600 204.900 ;
        RECT 98.300 204.000 99.000 204.400 ;
        RECT 95.100 203.700 95.500 203.800 ;
        RECT 96.500 203.700 96.900 203.800 ;
        RECT 93.400 203.100 93.800 203.500 ;
        RECT 95.100 203.400 96.900 203.700 ;
        RECT 96.200 203.100 96.500 203.400 ;
        RECT 98.200 203.100 98.600 203.500 ;
        RECT 93.400 202.800 94.400 203.100 ;
        RECT 94.000 201.100 94.400 202.800 ;
        RECT 96.200 201.100 96.600 203.100 ;
        RECT 98.300 201.100 98.900 203.100 ;
        RECT 100.600 201.100 101.000 205.400 ;
        RECT 101.400 205.500 104.200 205.600 ;
        RECT 101.400 205.400 104.300 205.500 ;
        RECT 101.400 205.300 106.300 205.400 ;
        RECT 101.400 201.100 101.800 205.300 ;
        RECT 103.900 205.100 106.300 205.300 ;
        RECT 103.000 204.500 105.700 204.800 ;
        RECT 103.000 204.400 103.400 204.500 ;
        RECT 105.300 204.400 105.700 204.500 ;
        RECT 106.000 204.500 106.300 205.100 ;
        RECT 107.000 205.200 107.300 206.800 ;
        RECT 107.800 206.400 108.200 206.500 ;
        RECT 107.800 206.100 109.700 206.400 ;
        RECT 109.300 206.000 109.700 206.100 ;
        RECT 108.500 205.700 108.900 205.800 ;
        RECT 110.200 205.700 110.600 207.400 ;
        RECT 111.400 207.200 111.800 207.400 ;
        RECT 113.400 207.200 113.700 207.900 ;
        RECT 114.300 207.200 114.600 207.900 ;
        RECT 115.100 207.700 116.900 207.900 ;
        RECT 117.500 207.700 119.300 207.900 ;
        RECT 116.200 207.200 116.600 207.400 ;
        RECT 117.800 207.200 118.200 207.400 ;
        RECT 119.800 207.200 120.100 207.900 ;
        RECT 120.700 207.700 122.500 207.900 ;
        RECT 121.000 207.200 121.400 207.400 ;
        RECT 123.000 207.200 123.300 207.900 ;
        RECT 123.800 207.500 124.200 209.900 ;
        RECT 126.000 209.200 126.400 209.900 ;
        RECT 125.400 208.900 126.400 209.200 ;
        RECT 128.200 208.900 128.600 209.900 ;
        RECT 130.300 209.200 130.900 209.900 ;
        RECT 130.200 208.900 130.900 209.200 ;
        RECT 125.400 208.500 125.800 208.900 ;
        RECT 128.200 208.600 128.500 208.900 ;
        RECT 126.200 208.200 126.600 208.600 ;
        RECT 127.100 208.300 128.500 208.600 ;
        RECT 130.200 208.500 130.600 208.900 ;
        RECT 127.100 208.200 127.500 208.300 ;
        RECT 111.000 206.900 111.800 207.200 ;
        RECT 111.000 206.800 111.400 206.900 ;
        RECT 112.500 206.800 113.800 207.200 ;
        RECT 114.200 206.800 115.500 207.200 ;
        RECT 116.200 206.900 117.000 207.200 ;
        RECT 116.600 206.800 117.000 206.900 ;
        RECT 117.400 206.900 118.200 207.200 ;
        RECT 117.400 206.800 117.800 206.900 ;
        RECT 118.900 206.800 120.200 207.200 ;
        RECT 120.600 206.900 121.400 207.200 ;
        RECT 120.600 206.800 121.000 206.900 ;
        RECT 122.100 206.800 123.400 207.200 ;
        RECT 124.200 207.100 125.000 207.200 ;
        RECT 126.300 207.100 126.600 208.200 ;
        RECT 129.400 207.800 129.800 208.200 ;
        RECT 129.400 207.200 129.700 207.800 ;
        RECT 131.100 207.700 131.500 207.800 ;
        RECT 132.600 207.700 133.000 209.900 ;
        RECT 134.200 208.200 134.600 209.900 ;
        RECT 131.100 207.400 133.000 207.700 ;
        RECT 129.100 207.100 129.700 207.200 ;
        RECT 124.200 206.800 129.700 207.100 ;
        RECT 111.800 205.800 112.200 206.600 ;
        RECT 112.500 206.200 112.800 206.800 ;
        RECT 112.500 205.800 113.000 206.200 ;
        RECT 115.200 206.100 115.500 206.800 ;
        RECT 113.400 205.800 115.500 206.100 ;
        RECT 115.800 205.800 116.200 206.600 ;
        RECT 118.200 205.800 118.600 206.600 ;
        RECT 118.900 206.100 119.200 206.800 ;
        RECT 119.800 206.100 120.200 206.200 ;
        RECT 118.900 205.800 120.200 206.100 ;
        RECT 121.400 205.800 121.800 206.600 ;
        RECT 108.500 205.400 110.600 205.700 ;
        RECT 107.000 204.900 108.200 205.200 ;
        RECT 106.700 204.500 107.100 204.600 ;
        RECT 106.000 204.200 107.100 204.500 ;
        RECT 107.900 204.400 108.200 204.900 ;
        RECT 107.900 204.200 108.600 204.400 ;
        RECT 107.900 204.000 109.000 204.200 ;
        RECT 108.300 203.800 109.000 204.000 ;
        RECT 104.700 203.700 105.100 203.800 ;
        RECT 106.100 203.700 106.500 203.800 ;
        RECT 103.000 203.100 103.400 203.500 ;
        RECT 104.700 203.400 106.500 203.700 ;
        RECT 105.800 203.100 106.100 203.400 ;
        RECT 107.800 203.100 108.200 203.500 ;
        RECT 103.000 202.800 104.000 203.100 ;
        RECT 103.600 201.100 104.000 202.800 ;
        RECT 105.800 201.100 106.200 203.100 ;
        RECT 107.900 201.100 108.500 203.100 ;
        RECT 110.200 201.100 110.600 205.400 ;
        RECT 112.500 205.100 112.800 205.800 ;
        RECT 113.400 205.200 113.700 205.800 ;
        RECT 113.400 205.100 113.800 205.200 ;
        RECT 112.300 204.800 112.800 205.100 ;
        RECT 113.100 204.800 113.800 205.100 ;
        RECT 114.200 205.100 114.600 205.200 ;
        RECT 115.200 205.100 115.500 205.800 ;
        RECT 118.900 205.100 119.200 205.800 ;
        RECT 119.800 205.100 120.200 205.200 ;
        RECT 122.100 205.100 122.400 206.800 ;
        RECT 125.700 206.700 126.100 206.800 ;
        RECT 124.900 206.200 125.300 206.300 ;
        RECT 126.200 206.200 126.600 206.300 ;
        RECT 124.900 205.900 127.400 206.200 ;
        RECT 127.000 205.800 127.400 205.900 ;
        RECT 123.800 205.500 126.600 205.600 ;
        RECT 123.800 205.400 126.700 205.500 ;
        RECT 123.800 205.300 128.700 205.400 ;
        RECT 123.000 205.100 123.400 205.200 ;
        RECT 114.200 204.800 114.900 205.100 ;
        RECT 115.200 204.800 115.700 205.100 ;
        RECT 112.300 201.100 112.700 204.800 ;
        RECT 113.100 204.200 113.400 204.800 ;
        RECT 113.000 203.800 113.400 204.200 ;
        RECT 114.600 204.200 114.900 204.800 ;
        RECT 114.600 203.800 115.000 204.200 ;
        RECT 115.300 201.100 115.700 204.800 ;
        RECT 118.700 204.800 119.200 205.100 ;
        RECT 119.500 204.800 120.200 205.100 ;
        RECT 121.900 204.800 122.400 205.100 ;
        RECT 122.700 204.800 123.400 205.100 ;
        RECT 118.700 201.100 119.100 204.800 ;
        RECT 119.500 204.200 119.800 204.800 ;
        RECT 121.900 204.200 122.300 204.800 ;
        RECT 122.700 204.200 123.000 204.800 ;
        RECT 119.400 203.800 119.800 204.200 ;
        RECT 121.400 203.800 122.300 204.200 ;
        RECT 122.600 203.800 123.400 204.200 ;
        RECT 121.900 201.100 122.300 203.800 ;
        RECT 123.800 201.100 124.200 205.300 ;
        RECT 126.300 205.100 128.700 205.300 ;
        RECT 125.400 204.500 128.100 204.800 ;
        RECT 125.400 204.400 125.800 204.500 ;
        RECT 127.700 204.400 128.100 204.500 ;
        RECT 128.400 204.500 128.700 205.100 ;
        RECT 129.400 205.200 129.700 206.800 ;
        RECT 130.200 206.400 130.600 206.500 ;
        RECT 130.200 206.100 132.100 206.400 ;
        RECT 131.700 206.000 132.100 206.100 ;
        RECT 130.900 205.700 131.300 205.800 ;
        RECT 132.600 205.700 133.000 207.400 ;
        RECT 130.900 205.400 133.000 205.700 ;
        RECT 129.400 204.900 130.600 205.200 ;
        RECT 129.100 204.500 129.500 204.600 ;
        RECT 128.400 204.200 129.500 204.500 ;
        RECT 130.300 204.400 130.600 204.900 ;
        RECT 130.300 204.000 131.000 204.400 ;
        RECT 127.100 203.700 127.500 203.800 ;
        RECT 128.500 203.700 128.900 203.800 ;
        RECT 125.400 203.100 125.800 203.500 ;
        RECT 127.100 203.400 128.900 203.700 ;
        RECT 128.200 203.100 128.500 203.400 ;
        RECT 130.200 203.100 130.600 203.500 ;
        RECT 125.400 202.800 126.400 203.100 ;
        RECT 126.000 201.100 126.400 202.800 ;
        RECT 128.200 201.100 128.600 203.100 ;
        RECT 130.300 201.100 130.900 203.100 ;
        RECT 132.600 201.100 133.000 205.400 ;
        RECT 134.100 207.900 134.600 208.200 ;
        RECT 134.100 207.200 134.400 207.900 ;
        RECT 135.800 207.600 136.200 209.900 ;
        RECT 134.900 207.300 136.200 207.600 ;
        RECT 137.400 207.600 137.800 209.900 ;
        RECT 139.000 207.600 139.400 209.900 ;
        RECT 134.100 206.800 134.600 207.200 ;
        RECT 134.100 205.100 134.400 206.800 ;
        RECT 134.900 206.500 135.200 207.300 ;
        RECT 137.400 207.200 139.400 207.600 ;
        RECT 142.200 207.500 142.600 209.900 ;
        RECT 144.400 209.200 144.800 209.900 ;
        RECT 143.800 208.900 144.800 209.200 ;
        RECT 146.600 208.900 147.000 209.900 ;
        RECT 148.700 209.200 149.300 209.900 ;
        RECT 148.600 208.900 149.300 209.200 ;
        RECT 143.800 208.500 144.200 208.900 ;
        RECT 146.600 208.600 146.900 208.900 ;
        RECT 144.600 208.200 145.000 208.600 ;
        RECT 145.500 208.300 146.900 208.600 ;
        RECT 148.600 208.500 149.000 208.900 ;
        RECT 145.500 208.200 145.900 208.300 ;
        RECT 134.700 206.100 135.200 206.500 ;
        RECT 134.900 205.100 135.200 206.100 ;
        RECT 135.700 206.200 136.100 206.600 ;
        RECT 135.700 206.100 136.200 206.200 ;
        RECT 135.700 205.800 137.800 206.100 ;
        RECT 139.000 205.800 139.400 207.200 ;
        RECT 142.600 207.100 143.400 207.200 ;
        RECT 144.700 207.100 145.000 208.200 ;
        RECT 149.500 207.700 149.900 207.800 ;
        RECT 151.000 207.700 151.400 209.900 ;
        RECT 151.800 208.000 152.200 209.900 ;
        RECT 153.400 208.000 153.800 209.900 ;
        RECT 151.800 207.900 153.800 208.000 ;
        RECT 154.200 207.900 154.600 209.900 ;
        RECT 155.300 208.200 155.700 209.900 ;
        RECT 155.300 207.900 156.200 208.200 ;
        RECT 151.900 207.700 153.700 207.900 ;
        RECT 149.500 207.400 151.400 207.700 ;
        RECT 147.500 207.100 147.900 207.200 ;
        RECT 142.600 206.800 148.100 207.100 ;
        RECT 144.100 206.700 144.500 206.800 ;
        RECT 143.300 206.200 143.700 206.300 ;
        RECT 143.300 205.900 145.800 206.200 ;
        RECT 145.400 205.800 145.800 205.900 ;
        RECT 137.400 205.400 139.400 205.800 ;
        RECT 134.100 204.600 134.600 205.100 ;
        RECT 134.900 204.800 136.200 205.100 ;
        RECT 134.200 201.100 134.600 204.600 ;
        RECT 135.800 201.100 136.200 204.800 ;
        RECT 137.400 201.100 137.800 205.400 ;
        RECT 139.000 201.100 139.400 205.400 ;
        RECT 142.200 205.500 145.000 205.600 ;
        RECT 142.200 205.400 145.100 205.500 ;
        RECT 142.200 205.300 147.100 205.400 ;
        RECT 142.200 201.100 142.600 205.300 ;
        RECT 144.700 205.100 147.100 205.300 ;
        RECT 143.800 204.500 146.500 204.800 ;
        RECT 143.800 204.400 144.200 204.500 ;
        RECT 146.100 204.400 146.500 204.500 ;
        RECT 146.800 204.500 147.100 205.100 ;
        RECT 147.800 205.200 148.100 206.800 ;
        RECT 148.600 206.400 149.000 206.500 ;
        RECT 148.600 206.100 150.500 206.400 ;
        RECT 150.100 206.000 150.500 206.100 ;
        RECT 149.300 205.700 149.700 205.800 ;
        RECT 151.000 205.700 151.400 207.400 ;
        RECT 152.200 207.200 152.600 207.400 ;
        RECT 154.200 207.200 154.500 207.900 ;
        RECT 151.800 206.900 152.600 207.200 ;
        RECT 151.800 206.800 152.200 206.900 ;
        RECT 153.300 206.800 154.600 207.200 ;
        RECT 152.600 205.800 153.000 206.600 ;
        RECT 153.300 206.200 153.600 206.800 ;
        RECT 153.300 205.800 153.800 206.200 ;
        RECT 155.800 206.100 156.200 207.900 ;
        RECT 157.400 207.600 157.800 209.900 ;
        RECT 159.000 208.200 159.400 209.900 ;
        RECT 159.000 207.900 159.500 208.200 ;
        RECT 156.600 206.800 157.000 207.600 ;
        RECT 157.400 207.300 158.700 207.600 ;
        RECT 157.500 206.200 157.900 206.600 ;
        RECT 154.200 205.800 156.200 206.100 ;
        RECT 157.400 205.800 157.900 206.200 ;
        RECT 158.400 206.500 158.700 207.300 ;
        RECT 159.200 207.200 159.500 207.900 ;
        RECT 159.000 206.800 159.500 207.200 ;
        RECT 158.400 206.100 158.900 206.500 ;
        RECT 149.300 205.400 151.400 205.700 ;
        RECT 147.800 204.900 149.000 205.200 ;
        RECT 147.500 204.500 147.900 204.600 ;
        RECT 146.800 204.200 147.900 204.500 ;
        RECT 148.700 204.400 149.000 204.900 ;
        RECT 148.700 204.200 149.400 204.400 ;
        RECT 148.700 204.000 149.800 204.200 ;
        RECT 149.100 203.800 149.800 204.000 ;
        RECT 145.500 203.700 145.900 203.800 ;
        RECT 146.900 203.700 147.300 203.800 ;
        RECT 143.800 203.100 144.200 203.500 ;
        RECT 145.500 203.400 147.300 203.700 ;
        RECT 146.600 203.100 146.900 203.400 ;
        RECT 148.600 203.100 149.000 203.500 ;
        RECT 143.800 202.800 144.800 203.100 ;
        RECT 144.400 201.100 144.800 202.800 ;
        RECT 146.600 201.100 147.000 203.100 ;
        RECT 148.700 201.100 149.300 203.100 ;
        RECT 151.000 201.100 151.400 205.400 ;
        RECT 153.300 205.100 153.600 205.800 ;
        RECT 154.200 205.200 154.500 205.800 ;
        RECT 154.200 205.100 154.600 205.200 ;
        RECT 153.100 204.800 153.600 205.100 ;
        RECT 153.900 204.800 154.600 205.100 ;
        RECT 153.100 201.100 153.500 204.800 ;
        RECT 153.900 204.200 154.200 204.800 ;
        RECT 155.000 204.400 155.400 205.200 ;
        RECT 153.800 203.800 154.200 204.200 ;
        RECT 155.800 201.100 156.200 205.800 ;
        RECT 158.400 205.100 158.700 206.100 ;
        RECT 159.200 205.100 159.500 206.800 ;
        RECT 157.400 204.800 158.700 205.100 ;
        RECT 157.400 201.100 157.800 204.800 ;
        RECT 159.000 204.600 159.500 205.100 ;
        RECT 160.600 207.700 161.000 209.900 ;
        RECT 162.700 209.200 163.300 209.900 ;
        RECT 162.700 208.900 163.400 209.200 ;
        RECT 165.000 208.900 165.400 209.900 ;
        RECT 167.200 209.200 167.600 209.900 ;
        RECT 167.200 208.900 168.200 209.200 ;
        RECT 163.000 208.500 163.400 208.900 ;
        RECT 165.100 208.600 165.400 208.900 ;
        RECT 165.100 208.300 166.500 208.600 ;
        RECT 166.100 208.200 166.500 208.300 ;
        RECT 167.000 208.200 167.400 208.600 ;
        RECT 167.800 208.500 168.200 208.900 ;
        RECT 162.100 207.700 162.500 207.800 ;
        RECT 160.600 207.400 162.500 207.700 ;
        RECT 160.600 205.700 161.000 207.400 ;
        RECT 164.100 207.100 164.500 207.200 ;
        RECT 167.000 207.100 167.300 208.200 ;
        RECT 169.400 207.500 169.800 209.900 ;
        RECT 170.200 208.000 170.600 209.900 ;
        RECT 171.800 208.000 172.200 209.900 ;
        RECT 170.200 207.900 172.200 208.000 ;
        RECT 172.600 207.900 173.000 209.900 ;
        RECT 173.700 208.200 174.100 209.900 ;
        RECT 173.700 207.900 174.600 208.200 ;
        RECT 170.300 207.700 172.100 207.900 ;
        RECT 170.600 207.200 171.000 207.400 ;
        RECT 172.600 207.200 172.900 207.900 ;
        RECT 168.600 207.100 169.400 207.200 ;
        RECT 163.900 206.800 169.400 207.100 ;
        RECT 170.200 206.900 171.000 207.200 ;
        RECT 171.700 207.100 173.000 207.200 ;
        RECT 173.400 207.100 173.800 207.200 ;
        RECT 170.200 206.800 170.600 206.900 ;
        RECT 171.700 206.800 173.800 207.100 ;
        RECT 163.000 206.400 163.400 206.500 ;
        RECT 161.500 206.100 163.400 206.400 ;
        RECT 161.500 206.000 161.900 206.100 ;
        RECT 162.300 205.700 162.700 205.800 ;
        RECT 160.600 205.400 162.700 205.700 ;
        RECT 159.000 201.100 159.400 204.600 ;
        RECT 160.600 201.100 161.000 205.400 ;
        RECT 163.900 205.200 164.200 206.800 ;
        RECT 167.500 206.700 167.900 206.800 ;
        RECT 167.000 206.200 167.400 206.300 ;
        RECT 168.300 206.200 168.700 206.300 ;
        RECT 166.200 205.900 168.700 206.200 ;
        RECT 166.200 205.800 166.600 205.900 ;
        RECT 171.000 205.800 171.400 206.600 ;
        RECT 167.000 205.500 169.800 205.600 ;
        RECT 166.900 205.400 169.800 205.500 ;
        RECT 163.000 204.900 164.200 205.200 ;
        RECT 164.900 205.300 169.800 205.400 ;
        RECT 164.900 205.100 167.300 205.300 ;
        RECT 163.000 204.400 163.300 204.900 ;
        RECT 162.600 204.000 163.300 204.400 ;
        RECT 164.100 204.500 164.500 204.600 ;
        RECT 164.900 204.500 165.200 205.100 ;
        RECT 164.100 204.200 165.200 204.500 ;
        RECT 165.500 204.500 168.200 204.800 ;
        RECT 165.500 204.400 165.900 204.500 ;
        RECT 167.800 204.400 168.200 204.500 ;
        RECT 164.700 203.700 165.100 203.800 ;
        RECT 166.100 203.700 166.500 203.800 ;
        RECT 163.000 203.100 163.400 203.500 ;
        RECT 164.700 203.400 166.500 203.700 ;
        RECT 165.100 203.100 165.400 203.400 ;
        RECT 167.800 203.100 168.200 203.500 ;
        RECT 162.700 201.100 163.300 203.100 ;
        RECT 165.000 201.100 165.400 203.100 ;
        RECT 167.200 202.800 168.200 203.100 ;
        RECT 167.200 201.100 167.600 202.800 ;
        RECT 169.400 201.100 169.800 205.300 ;
        RECT 171.700 205.100 172.000 206.800 ;
        RECT 174.200 206.100 174.600 207.900 ;
        RECT 175.000 206.800 175.400 207.600 ;
        RECT 175.800 207.500 176.200 209.900 ;
        RECT 178.000 209.200 178.400 209.900 ;
        RECT 177.400 208.900 178.400 209.200 ;
        RECT 180.200 208.900 180.600 209.900 ;
        RECT 182.300 209.200 182.900 209.900 ;
        RECT 182.200 208.900 182.900 209.200 ;
        RECT 177.400 208.500 177.800 208.900 ;
        RECT 180.200 208.600 180.500 208.900 ;
        RECT 178.200 208.200 178.600 208.600 ;
        RECT 179.100 208.300 180.500 208.600 ;
        RECT 182.200 208.500 182.600 208.900 ;
        RECT 179.100 208.200 179.500 208.300 ;
        RECT 176.200 207.100 177.000 207.200 ;
        RECT 178.300 207.100 178.600 208.200 ;
        RECT 183.100 207.700 183.500 207.800 ;
        RECT 184.600 207.700 185.000 209.900 ;
        RECT 183.100 207.400 185.000 207.700 ;
        RECT 181.100 207.100 181.500 207.200 ;
        RECT 176.200 206.800 181.700 207.100 ;
        RECT 177.700 206.700 178.100 206.800 ;
        RECT 172.600 205.800 174.600 206.100 ;
        RECT 176.900 206.200 177.300 206.300 ;
        RECT 178.200 206.200 178.600 206.300 ;
        RECT 181.400 206.200 181.700 206.800 ;
        RECT 182.200 206.400 182.600 206.500 ;
        RECT 176.900 205.900 179.400 206.200 ;
        RECT 179.000 205.800 179.400 205.900 ;
        RECT 181.400 205.800 181.800 206.200 ;
        RECT 182.200 206.100 184.100 206.400 ;
        RECT 183.700 206.000 184.100 206.100 ;
        RECT 172.600 205.200 172.900 205.800 ;
        RECT 172.600 205.100 173.000 205.200 ;
        RECT 171.500 204.800 172.000 205.100 ;
        RECT 172.300 204.800 173.000 205.100 ;
        RECT 171.500 201.100 171.900 204.800 ;
        RECT 172.300 204.200 172.600 204.800 ;
        RECT 173.400 204.400 173.800 205.200 ;
        RECT 172.200 203.800 172.600 204.200 ;
        RECT 174.200 201.100 174.600 205.800 ;
        RECT 175.800 205.500 178.600 205.600 ;
        RECT 175.800 205.400 178.700 205.500 ;
        RECT 175.800 205.300 180.700 205.400 ;
        RECT 175.800 201.100 176.200 205.300 ;
        RECT 178.300 205.100 180.700 205.300 ;
        RECT 177.400 204.500 180.100 204.800 ;
        RECT 177.400 204.400 177.800 204.500 ;
        RECT 179.700 204.400 180.100 204.500 ;
        RECT 180.400 204.500 180.700 205.100 ;
        RECT 181.400 205.200 181.700 205.800 ;
        RECT 182.900 205.700 183.300 205.800 ;
        RECT 184.600 205.700 185.000 207.400 ;
        RECT 182.900 205.400 185.000 205.700 ;
        RECT 181.400 204.900 182.600 205.200 ;
        RECT 181.100 204.500 181.500 204.600 ;
        RECT 180.400 204.200 181.500 204.500 ;
        RECT 182.300 204.400 182.600 204.900 ;
        RECT 183.000 204.800 183.400 205.400 ;
        RECT 182.300 204.000 183.000 204.400 ;
        RECT 179.100 203.700 179.500 203.800 ;
        RECT 180.500 203.700 180.900 203.800 ;
        RECT 177.400 203.100 177.800 203.500 ;
        RECT 179.100 203.400 180.900 203.700 ;
        RECT 180.200 203.100 180.500 203.400 ;
        RECT 182.200 203.100 182.600 203.500 ;
        RECT 177.400 202.800 178.400 203.100 ;
        RECT 178.000 201.100 178.400 202.800 ;
        RECT 180.200 201.100 180.600 203.100 ;
        RECT 182.300 201.100 182.900 203.100 ;
        RECT 184.600 201.100 185.000 205.400 ;
        RECT 186.200 207.600 186.600 209.900 ;
        RECT 187.800 207.600 188.200 209.900 ;
        RECT 191.800 207.600 192.200 209.900 ;
        RECT 193.400 207.600 193.800 209.900 ;
        RECT 195.000 207.600 195.400 209.900 ;
        RECT 196.600 207.600 197.000 209.900 ;
        RECT 200.100 208.000 200.500 209.500 ;
        RECT 202.200 208.500 202.600 209.500 ;
        RECT 186.200 207.200 188.200 207.600 ;
        RECT 191.000 207.200 192.200 207.600 ;
        RECT 192.700 207.200 193.800 207.600 ;
        RECT 194.300 207.200 195.400 207.600 ;
        RECT 196.100 207.200 197.000 207.600 ;
        RECT 199.700 207.700 200.500 208.000 ;
        RECT 199.700 207.500 200.100 207.700 ;
        RECT 199.700 207.200 200.000 207.500 ;
        RECT 202.300 207.400 202.600 208.500 ;
        RECT 203.000 208.000 203.400 209.900 ;
        RECT 204.600 208.000 205.000 209.900 ;
        RECT 203.000 207.900 205.000 208.000 ;
        RECT 205.400 207.900 205.800 209.900 ;
        RECT 206.500 208.200 206.900 209.900 ;
        RECT 209.900 208.200 210.300 209.900 ;
        RECT 206.500 207.900 207.400 208.200 ;
        RECT 203.100 207.700 204.900 207.900 ;
        RECT 186.200 205.800 186.600 207.200 ;
        RECT 190.200 206.100 190.600 206.200 ;
        RECT 191.000 206.100 191.400 207.200 ;
        RECT 192.700 206.900 193.100 207.200 ;
        RECT 194.300 206.900 194.700 207.200 ;
        RECT 196.100 206.900 196.500 207.200 ;
        RECT 191.800 206.500 193.100 206.900 ;
        RECT 193.500 206.500 194.700 206.900 ;
        RECT 195.200 206.500 196.500 206.900 ;
        RECT 199.000 206.800 200.000 207.200 ;
        RECT 200.500 207.100 202.600 207.400 ;
        RECT 203.400 207.200 203.800 207.400 ;
        RECT 205.400 207.200 205.700 207.900 ;
        RECT 200.500 206.900 201.000 207.100 ;
        RECT 190.200 205.800 191.400 206.100 ;
        RECT 192.700 205.800 193.100 206.500 ;
        RECT 194.300 205.800 194.700 206.500 ;
        RECT 196.100 205.800 196.500 206.500 ;
        RECT 198.200 206.100 198.600 206.200 ;
        RECT 199.000 206.100 199.400 206.200 ;
        RECT 198.200 205.800 199.400 206.100 ;
        RECT 186.200 205.400 188.200 205.800 ;
        RECT 191.000 205.400 192.200 205.800 ;
        RECT 192.700 205.400 193.800 205.800 ;
        RECT 194.300 205.400 195.400 205.800 ;
        RECT 196.100 205.400 197.000 205.800 ;
        RECT 199.000 205.400 199.400 205.800 ;
        RECT 186.200 201.100 186.600 205.400 ;
        RECT 187.800 201.100 188.200 205.400 ;
        RECT 191.800 201.100 192.200 205.400 ;
        RECT 193.400 201.100 193.800 205.400 ;
        RECT 195.000 201.100 195.400 205.400 ;
        RECT 196.600 201.100 197.000 205.400 ;
        RECT 199.700 204.900 200.000 206.800 ;
        RECT 200.300 206.500 201.000 206.900 ;
        RECT 203.000 206.900 203.800 207.200 ;
        RECT 203.000 206.800 203.400 206.900 ;
        RECT 204.500 206.800 205.800 207.200 ;
        RECT 200.700 205.500 201.000 206.500 ;
        RECT 201.400 205.800 201.800 206.600 ;
        RECT 202.200 205.800 202.600 206.600 ;
        RECT 203.800 205.800 204.200 206.600 ;
        RECT 200.700 205.200 202.600 205.500 ;
        RECT 199.700 204.600 200.500 204.900 ;
        RECT 200.100 202.200 200.500 204.600 ;
        RECT 202.300 203.500 202.600 205.200 ;
        RECT 204.500 205.100 204.800 206.800 ;
        RECT 207.000 206.100 207.400 207.900 ;
        RECT 209.400 207.900 210.300 208.200 ;
        RECT 207.800 206.800 208.200 207.600 ;
        RECT 208.600 206.800 209.000 207.600 ;
        RECT 205.400 205.800 207.400 206.100 ;
        RECT 205.400 205.200 205.700 205.800 ;
        RECT 205.400 205.100 205.800 205.200 ;
        RECT 199.800 201.800 200.500 202.200 ;
        RECT 200.100 201.100 200.500 201.800 ;
        RECT 202.200 201.500 202.600 203.500 ;
        RECT 204.300 204.800 204.800 205.100 ;
        RECT 205.100 204.800 205.800 205.100 ;
        RECT 204.300 201.100 204.700 204.800 ;
        RECT 205.100 204.200 205.400 204.800 ;
        RECT 206.200 204.400 206.600 205.200 ;
        RECT 205.000 203.800 205.400 204.200 ;
        RECT 207.000 201.100 207.400 205.800 ;
        RECT 209.400 201.100 209.800 207.900 ;
        RECT 211.000 207.700 211.400 209.900 ;
        RECT 213.100 209.200 213.700 209.900 ;
        RECT 213.100 208.900 213.800 209.200 ;
        RECT 215.400 208.900 215.800 209.900 ;
        RECT 217.600 209.200 218.000 209.900 ;
        RECT 217.600 208.900 218.600 209.200 ;
        RECT 213.400 208.500 213.800 208.900 ;
        RECT 215.500 208.600 215.800 208.900 ;
        RECT 215.500 208.300 216.900 208.600 ;
        RECT 216.500 208.200 216.900 208.300 ;
        RECT 217.400 208.200 217.800 208.600 ;
        RECT 218.200 208.500 218.600 208.900 ;
        RECT 212.500 207.700 212.900 207.800 ;
        RECT 211.000 207.400 212.900 207.700 ;
        RECT 211.000 205.700 211.400 207.400 ;
        RECT 214.500 207.100 214.900 207.200 ;
        RECT 216.600 207.100 217.000 207.200 ;
        RECT 217.400 207.100 217.700 208.200 ;
        RECT 219.800 207.500 220.200 209.900 ;
        RECT 220.900 208.200 221.300 209.900 ;
        RECT 220.900 207.900 221.800 208.200 ;
        RECT 223.000 208.000 223.400 209.900 ;
        RECT 224.600 208.000 225.000 209.900 ;
        RECT 223.000 207.900 225.000 208.000 ;
        RECT 225.400 207.900 225.800 209.900 ;
        RECT 219.000 207.100 219.800 207.200 ;
        RECT 214.300 206.800 219.800 207.100 ;
        RECT 213.400 206.400 213.800 206.500 ;
        RECT 211.900 206.100 213.800 206.400 ;
        RECT 211.900 206.000 212.300 206.100 ;
        RECT 212.700 205.700 213.100 205.800 ;
        RECT 211.000 205.400 213.100 205.700 ;
        RECT 210.200 204.400 210.600 205.200 ;
        RECT 211.000 201.100 211.400 205.400 ;
        RECT 214.300 205.200 214.600 206.800 ;
        RECT 217.900 206.700 218.300 206.800 ;
        RECT 218.700 206.200 219.100 206.300 ;
        RECT 215.000 206.100 215.400 206.200 ;
        RECT 216.600 206.100 219.100 206.200 ;
        RECT 215.000 205.900 219.100 206.100 ;
        RECT 215.000 205.800 217.000 205.900 ;
        RECT 217.400 205.500 220.200 205.600 ;
        RECT 217.300 205.400 220.200 205.500 ;
        RECT 213.400 204.900 214.600 205.200 ;
        RECT 215.300 205.300 220.200 205.400 ;
        RECT 215.300 205.100 217.700 205.300 ;
        RECT 213.400 204.400 213.700 204.900 ;
        RECT 213.000 204.000 213.700 204.400 ;
        RECT 214.500 204.500 214.900 204.600 ;
        RECT 215.300 204.500 215.600 205.100 ;
        RECT 214.500 204.200 215.600 204.500 ;
        RECT 215.900 204.500 218.600 204.800 ;
        RECT 215.900 204.400 216.300 204.500 ;
        RECT 218.200 204.400 218.600 204.500 ;
        RECT 215.100 203.700 215.500 203.800 ;
        RECT 216.500 203.700 216.900 203.800 ;
        RECT 213.400 203.100 213.800 203.500 ;
        RECT 215.100 203.400 216.900 203.700 ;
        RECT 215.500 203.100 215.800 203.400 ;
        RECT 218.200 203.100 218.600 203.500 ;
        RECT 213.100 201.100 213.700 203.100 ;
        RECT 215.400 201.100 215.800 203.100 ;
        RECT 217.600 202.800 218.600 203.100 ;
        RECT 217.600 201.100 218.000 202.800 ;
        RECT 219.800 201.100 220.200 205.300 ;
        RECT 220.600 204.400 221.000 205.200 ;
        RECT 221.400 201.100 221.800 207.900 ;
        RECT 223.100 207.700 224.900 207.900 ;
        RECT 222.200 206.800 222.600 207.600 ;
        RECT 223.400 207.200 223.800 207.400 ;
        RECT 225.400 207.200 225.700 207.900 ;
        RECT 227.000 207.600 227.400 209.900 ;
        RECT 228.600 207.600 229.000 209.900 ;
        RECT 227.000 207.200 229.000 207.600 ;
        RECT 223.000 206.900 223.800 207.200 ;
        RECT 223.000 206.800 223.400 206.900 ;
        RECT 224.500 206.800 225.800 207.200 ;
        RECT 223.800 205.800 224.200 206.600 ;
        RECT 224.500 206.200 224.800 206.800 ;
        RECT 224.500 205.800 225.000 206.200 ;
        RECT 227.000 205.800 227.400 207.200 ;
        RECT 224.500 205.100 224.800 205.800 ;
        RECT 227.000 205.400 229.000 205.800 ;
        RECT 225.400 205.100 225.800 205.200 ;
        RECT 224.300 204.800 224.800 205.100 ;
        RECT 225.100 204.800 225.800 205.100 ;
        RECT 224.300 201.100 224.700 204.800 ;
        RECT 225.100 204.200 225.400 204.800 ;
        RECT 225.000 203.800 225.400 204.200 ;
        RECT 227.000 201.100 227.400 205.400 ;
        RECT 228.600 201.100 229.000 205.400 ;
        RECT 0.600 195.600 1.000 199.900 ;
        RECT 2.700 197.900 3.300 199.900 ;
        RECT 5.000 197.900 5.400 199.900 ;
        RECT 7.200 198.200 7.600 199.900 ;
        RECT 7.200 197.900 8.200 198.200 ;
        RECT 3.000 197.500 3.400 197.900 ;
        RECT 5.100 197.600 5.400 197.900 ;
        RECT 4.700 197.300 6.500 197.600 ;
        RECT 7.800 197.500 8.200 197.900 ;
        RECT 4.700 197.200 5.100 197.300 ;
        RECT 6.100 197.200 6.500 197.300 ;
        RECT 2.600 196.600 3.300 197.000 ;
        RECT 3.000 196.100 3.300 196.600 ;
        RECT 4.100 196.500 5.200 196.800 ;
        RECT 4.100 196.400 4.500 196.500 ;
        RECT 3.000 195.800 4.200 196.100 ;
        RECT 0.600 195.300 2.700 195.600 ;
        RECT 0.600 193.600 1.000 195.300 ;
        RECT 2.300 195.200 2.700 195.300 ;
        RECT 1.500 194.900 1.900 195.000 ;
        RECT 1.500 194.600 3.400 194.900 ;
        RECT 3.000 194.500 3.400 194.600 ;
        RECT 3.900 194.200 4.200 195.800 ;
        RECT 4.900 195.900 5.200 196.500 ;
        RECT 5.500 196.500 5.900 196.600 ;
        RECT 7.800 196.500 8.200 196.600 ;
        RECT 5.500 196.200 8.200 196.500 ;
        RECT 4.900 195.700 7.300 195.900 ;
        RECT 9.400 195.700 9.800 199.900 ;
        RECT 10.600 196.800 11.000 197.200 ;
        RECT 10.600 196.200 10.900 196.800 ;
        RECT 11.300 196.200 11.700 199.900 ;
        RECT 14.500 197.200 14.900 199.900 ;
        RECT 17.700 199.200 18.100 199.900 ;
        RECT 17.700 198.800 18.600 199.200 ;
        RECT 13.400 196.800 14.200 197.200 ;
        RECT 14.500 196.800 15.400 197.200 ;
        RECT 17.000 196.800 17.400 197.200 ;
        RECT 13.800 196.200 14.100 196.800 ;
        RECT 14.500 196.200 14.900 196.800 ;
        RECT 17.000 196.200 17.300 196.800 ;
        RECT 17.700 196.200 18.100 198.800 ;
        RECT 20.900 197.200 21.300 199.900 ;
        RECT 19.800 196.800 20.600 197.200 ;
        RECT 20.900 196.800 21.800 197.200 ;
        RECT 20.200 196.200 20.500 196.800 ;
        RECT 20.900 196.200 21.300 196.800 ;
        RECT 10.200 195.900 10.900 196.200 ;
        RECT 11.200 195.900 11.700 196.200 ;
        RECT 13.400 195.900 14.100 196.200 ;
        RECT 14.400 195.900 14.900 196.200 ;
        RECT 16.600 195.900 17.300 196.200 ;
        RECT 17.600 195.900 18.100 196.200 ;
        RECT 19.800 195.900 20.500 196.200 ;
        RECT 20.800 195.900 21.300 196.200 ;
        RECT 24.300 196.200 24.700 199.900 ;
        RECT 25.000 196.800 25.800 197.200 ;
        RECT 26.600 196.800 27.000 197.200 ;
        RECT 25.100 196.200 25.400 196.800 ;
        RECT 26.600 196.200 26.900 196.800 ;
        RECT 27.300 196.200 27.700 199.900 ;
        RECT 24.300 195.900 24.800 196.200 ;
        RECT 25.100 195.900 25.800 196.200 ;
        RECT 10.200 195.800 10.600 195.900 ;
        RECT 4.900 195.600 9.800 195.700 ;
        RECT 6.900 195.500 9.800 195.600 ;
        RECT 7.000 195.400 9.800 195.500 ;
        RECT 6.200 195.100 6.600 195.200 ;
        RECT 10.200 195.100 10.600 195.200 ;
        RECT 11.200 195.100 11.500 195.900 ;
        RECT 13.400 195.800 13.800 195.900 ;
        RECT 6.200 194.800 8.700 195.100 ;
        RECT 10.200 194.800 11.500 195.100 ;
        RECT 7.000 194.700 7.400 194.800 ;
        RECT 8.300 194.700 8.700 194.800 ;
        RECT 7.500 194.200 7.900 194.300 ;
        RECT 11.200 194.200 11.500 194.800 ;
        RECT 11.800 194.400 12.200 195.200 ;
        RECT 14.400 194.200 14.700 195.900 ;
        RECT 16.600 195.800 17.000 195.900 ;
        RECT 15.000 194.400 15.400 195.200 ;
        RECT 17.600 194.200 17.900 195.900 ;
        RECT 19.800 195.800 20.200 195.900 ;
        RECT 18.200 194.400 18.600 195.200 ;
        RECT 20.800 194.200 21.100 195.900 ;
        RECT 21.400 195.100 21.800 195.200 ;
        RECT 23.000 195.100 23.400 195.200 ;
        RECT 23.800 195.100 24.200 195.200 ;
        RECT 21.400 194.800 24.200 195.100 ;
        RECT 21.400 194.400 21.800 194.800 ;
        RECT 23.800 194.400 24.200 194.800 ;
        RECT 24.500 195.100 24.800 195.900 ;
        RECT 25.400 195.800 25.800 195.900 ;
        RECT 26.200 195.900 26.900 196.200 ;
        RECT 27.200 195.900 27.700 196.200 ;
        RECT 26.200 195.800 26.600 195.900 ;
        RECT 26.200 195.100 26.500 195.800 ;
        RECT 24.500 194.800 26.500 195.100 ;
        RECT 24.500 194.200 24.800 194.800 ;
        RECT 27.200 194.200 27.500 195.900 ;
        RECT 29.400 195.700 29.800 199.900 ;
        RECT 31.600 198.200 32.000 199.900 ;
        RECT 31.000 197.900 32.000 198.200 ;
        RECT 33.800 197.900 34.200 199.900 ;
        RECT 35.900 197.900 36.500 199.900 ;
        RECT 31.000 197.500 31.400 197.900 ;
        RECT 33.800 197.600 34.100 197.900 ;
        RECT 32.700 197.300 34.500 197.600 ;
        RECT 35.800 197.500 36.200 197.900 ;
        RECT 32.700 197.200 33.100 197.300 ;
        RECT 34.100 197.200 34.500 197.300 ;
        RECT 31.000 196.500 31.400 196.600 ;
        RECT 33.300 196.500 33.700 196.600 ;
        RECT 31.000 196.200 33.700 196.500 ;
        RECT 34.000 196.500 35.100 196.800 ;
        RECT 34.000 195.900 34.300 196.500 ;
        RECT 34.700 196.400 35.100 196.500 ;
        RECT 35.900 196.600 36.600 197.000 ;
        RECT 35.900 196.100 36.200 196.600 ;
        RECT 31.900 195.700 34.300 195.900 ;
        RECT 29.400 195.600 34.300 195.700 ;
        RECT 35.000 195.800 36.200 196.100 ;
        RECT 29.400 195.500 32.300 195.600 ;
        RECT 29.400 195.400 32.200 195.500 ;
        RECT 35.000 195.200 35.300 195.800 ;
        RECT 38.200 195.600 38.600 199.900 ;
        RECT 36.500 195.300 38.600 195.600 ;
        RECT 40.600 195.700 41.000 199.900 ;
        RECT 42.800 198.200 43.200 199.900 ;
        RECT 42.200 197.900 43.200 198.200 ;
        RECT 45.000 197.900 45.400 199.900 ;
        RECT 47.100 197.900 47.700 199.900 ;
        RECT 42.200 197.500 42.600 197.900 ;
        RECT 45.000 197.600 45.300 197.900 ;
        RECT 43.900 197.300 45.700 197.600 ;
        RECT 47.000 197.500 47.400 197.900 ;
        RECT 43.900 197.200 44.300 197.300 ;
        RECT 45.300 197.200 45.700 197.300 ;
        RECT 47.500 197.000 48.200 197.200 ;
        RECT 47.100 196.800 48.200 197.000 ;
        RECT 42.200 196.500 42.600 196.600 ;
        RECT 44.500 196.500 44.900 196.600 ;
        RECT 42.200 196.200 44.900 196.500 ;
        RECT 45.200 196.500 46.300 196.800 ;
        RECT 45.200 195.900 45.500 196.500 ;
        RECT 45.900 196.400 46.300 196.500 ;
        RECT 47.100 196.600 47.800 196.800 ;
        RECT 47.100 196.100 47.400 196.600 ;
        RECT 43.100 195.700 45.500 195.900 ;
        RECT 40.600 195.600 45.500 195.700 ;
        RECT 46.200 195.800 47.400 196.100 ;
        RECT 40.600 195.500 43.500 195.600 ;
        RECT 40.600 195.400 43.400 195.500 ;
        RECT 36.500 195.200 36.900 195.300 ;
        RECT 27.800 194.400 28.200 195.200 ;
        RECT 32.600 195.100 33.000 195.200 ;
        RECT 30.500 194.800 33.000 195.100 ;
        RECT 35.000 194.800 35.400 195.200 ;
        RECT 37.300 194.900 37.700 195.000 ;
        RECT 30.500 194.700 30.900 194.800 ;
        RECT 31.800 194.700 32.200 194.800 ;
        RECT 31.300 194.200 31.700 194.300 ;
        RECT 35.000 194.200 35.300 194.800 ;
        RECT 35.800 194.600 37.700 194.900 ;
        RECT 35.800 194.500 36.200 194.600 ;
        RECT 3.900 193.900 9.400 194.200 ;
        RECT 4.100 193.800 4.500 193.900 ;
        RECT 6.200 193.800 6.600 193.900 ;
        RECT 0.600 193.300 2.500 193.600 ;
        RECT 0.600 191.100 1.000 193.300 ;
        RECT 2.100 193.200 2.500 193.300 ;
        RECT 7.000 192.800 7.300 193.900 ;
        RECT 8.600 193.800 9.400 193.900 ;
        RECT 10.200 193.800 11.500 194.200 ;
        RECT 12.600 194.100 13.000 194.200 ;
        RECT 12.200 193.800 13.000 194.100 ;
        RECT 13.400 193.800 14.700 194.200 ;
        RECT 15.800 194.100 16.200 194.200 ;
        RECT 15.400 193.800 16.200 194.100 ;
        RECT 16.600 193.800 17.900 194.200 ;
        RECT 19.000 194.100 19.400 194.200 ;
        RECT 18.600 193.800 19.400 194.100 ;
        RECT 19.800 193.800 21.100 194.200 ;
        RECT 22.200 194.100 22.600 194.200 ;
        RECT 23.000 194.100 23.400 194.200 ;
        RECT 21.800 193.800 23.800 194.100 ;
        RECT 24.500 193.800 25.800 194.200 ;
        RECT 26.200 193.800 27.500 194.200 ;
        RECT 28.600 194.100 29.000 194.200 ;
        RECT 28.200 193.800 29.000 194.100 ;
        RECT 29.800 193.900 35.300 194.200 ;
        RECT 29.800 193.800 30.600 193.900 ;
        RECT 6.100 192.700 6.500 192.800 ;
        RECT 3.000 192.100 3.400 192.500 ;
        RECT 5.100 192.400 6.500 192.700 ;
        RECT 7.000 192.400 7.400 192.800 ;
        RECT 5.100 192.100 5.400 192.400 ;
        RECT 7.800 192.100 8.200 192.500 ;
        RECT 2.700 191.800 3.400 192.100 ;
        RECT 2.700 191.100 3.300 191.800 ;
        RECT 5.000 191.100 5.400 192.100 ;
        RECT 7.200 191.800 8.200 192.100 ;
        RECT 7.200 191.100 7.600 191.800 ;
        RECT 9.400 191.100 9.800 193.500 ;
        RECT 10.300 193.100 10.600 193.800 ;
        RECT 12.200 193.600 12.600 193.800 ;
        RECT 11.100 193.100 12.900 193.300 ;
        RECT 13.500 193.100 13.800 193.800 ;
        RECT 15.400 193.600 15.800 193.800 ;
        RECT 14.300 193.100 16.100 193.300 ;
        RECT 16.700 193.100 17.000 193.800 ;
        RECT 18.600 193.600 19.000 193.800 ;
        RECT 17.500 193.100 19.300 193.300 ;
        RECT 19.900 193.100 20.200 193.800 ;
        RECT 21.800 193.600 22.200 193.800 ;
        RECT 23.400 193.600 23.800 193.800 ;
        RECT 20.700 193.100 22.500 193.300 ;
        RECT 23.100 193.100 24.900 193.300 ;
        RECT 25.400 193.100 25.700 193.800 ;
        RECT 26.300 193.100 26.600 193.800 ;
        RECT 28.200 193.600 28.600 193.800 ;
        RECT 27.100 193.100 28.900 193.300 ;
        RECT 10.200 191.100 10.600 193.100 ;
        RECT 11.000 193.000 13.000 193.100 ;
        RECT 11.000 191.100 11.400 193.000 ;
        RECT 12.600 191.100 13.000 193.000 ;
        RECT 13.400 191.100 13.800 193.100 ;
        RECT 14.200 193.000 16.200 193.100 ;
        RECT 14.200 191.100 14.600 193.000 ;
        RECT 15.800 191.100 16.200 193.000 ;
        RECT 16.600 191.100 17.000 193.100 ;
        RECT 17.400 193.000 19.400 193.100 ;
        RECT 17.400 191.100 17.800 193.000 ;
        RECT 19.000 191.100 19.400 193.000 ;
        RECT 19.800 191.100 20.200 193.100 ;
        RECT 20.600 193.000 22.600 193.100 ;
        RECT 20.600 191.100 21.000 193.000 ;
        RECT 22.200 191.100 22.600 193.000 ;
        RECT 23.000 193.000 25.000 193.100 ;
        RECT 23.000 191.100 23.400 193.000 ;
        RECT 24.600 191.100 25.000 193.000 ;
        RECT 25.400 191.100 25.800 193.100 ;
        RECT 26.200 191.100 26.600 193.100 ;
        RECT 27.000 193.000 29.000 193.100 ;
        RECT 27.000 191.100 27.400 193.000 ;
        RECT 28.600 191.100 29.000 193.000 ;
        RECT 29.400 191.100 29.800 193.500 ;
        RECT 31.900 192.800 32.200 193.900 ;
        RECT 34.700 193.800 35.100 193.900 ;
        RECT 38.200 193.600 38.600 195.300 ;
        RECT 43.800 195.100 44.200 195.200 ;
        RECT 45.400 195.100 45.800 195.200 ;
        RECT 41.700 194.800 45.800 195.100 ;
        RECT 41.700 194.700 42.100 194.800 ;
        RECT 42.500 194.200 42.900 194.300 ;
        RECT 46.200 194.200 46.500 195.800 ;
        RECT 49.400 195.600 49.800 199.900 ;
        RECT 50.600 196.800 51.000 197.200 ;
        RECT 50.600 196.200 50.900 196.800 ;
        RECT 51.300 196.200 51.700 199.900 ;
        RECT 55.300 196.400 55.700 199.900 ;
        RECT 57.400 197.500 57.800 199.500 ;
        RECT 50.200 195.900 50.900 196.200 ;
        RECT 51.200 195.900 51.700 196.200 ;
        RECT 54.900 196.100 55.700 196.400 ;
        RECT 50.200 195.800 50.600 195.900 ;
        RECT 47.700 195.300 49.800 195.600 ;
        RECT 47.700 195.200 48.100 195.300 ;
        RECT 48.500 194.900 48.900 195.000 ;
        RECT 47.000 194.600 48.900 194.900 ;
        RECT 47.000 194.500 47.400 194.600 ;
        RECT 41.000 193.900 46.500 194.200 ;
        RECT 41.000 193.800 41.800 193.900 ;
        RECT 36.700 193.300 38.600 193.600 ;
        RECT 36.700 193.200 37.100 193.300 ;
        RECT 31.000 192.100 31.400 192.500 ;
        RECT 31.800 192.400 32.200 192.800 ;
        RECT 32.700 192.700 33.100 192.800 ;
        RECT 32.700 192.400 34.100 192.700 ;
        RECT 33.800 192.100 34.100 192.400 ;
        RECT 35.800 192.100 36.200 192.500 ;
        RECT 31.000 191.800 32.000 192.100 ;
        RECT 31.600 191.100 32.000 191.800 ;
        RECT 33.800 191.100 34.200 192.100 ;
        RECT 35.800 191.800 36.500 192.100 ;
        RECT 35.900 191.100 36.500 191.800 ;
        RECT 38.200 191.100 38.600 193.300 ;
        RECT 40.600 191.100 41.000 193.500 ;
        RECT 43.100 192.800 43.400 193.900 ;
        RECT 45.900 193.800 46.300 193.900 ;
        RECT 49.400 193.600 49.800 195.300 ;
        RECT 51.200 194.200 51.500 195.900 ;
        RECT 51.800 194.400 52.200 195.200 ;
        RECT 54.200 194.800 54.600 195.600 ;
        RECT 54.900 194.200 55.200 196.100 ;
        RECT 57.500 195.800 57.800 197.500 ;
        RECT 59.500 196.200 59.900 199.900 ;
        RECT 60.200 196.800 60.600 197.200 ;
        RECT 60.300 196.200 60.600 196.800 ;
        RECT 59.500 195.900 60.000 196.200 ;
        RECT 60.300 195.900 61.000 196.200 ;
        RECT 55.900 195.500 57.800 195.800 ;
        RECT 55.900 194.500 56.200 195.500 ;
        RECT 50.200 193.800 51.500 194.200 ;
        RECT 52.600 194.100 53.000 194.200 ;
        RECT 52.200 193.800 53.000 194.100 ;
        RECT 54.200 193.800 55.200 194.200 ;
        RECT 55.500 194.100 56.200 194.500 ;
        RECT 56.600 194.400 57.000 195.200 ;
        RECT 57.400 194.400 57.800 195.200 ;
        RECT 59.000 194.400 59.400 195.200 ;
        RECT 59.700 194.200 60.000 195.900 ;
        RECT 60.600 195.800 61.000 195.900 ;
        RECT 61.400 195.700 61.800 199.900 ;
        RECT 63.600 198.200 64.000 199.900 ;
        RECT 63.000 197.900 64.000 198.200 ;
        RECT 65.800 197.900 66.200 199.900 ;
        RECT 67.900 197.900 68.500 199.900 ;
        RECT 63.000 197.500 63.400 197.900 ;
        RECT 65.800 197.600 66.100 197.900 ;
        RECT 64.700 197.300 66.500 197.600 ;
        RECT 67.800 197.500 68.200 197.900 ;
        RECT 64.700 197.200 65.100 197.300 ;
        RECT 66.100 197.200 66.500 197.300 ;
        RECT 63.000 196.500 63.400 196.600 ;
        RECT 65.300 196.500 65.700 196.600 ;
        RECT 63.000 196.200 65.700 196.500 ;
        RECT 66.000 196.500 67.100 196.800 ;
        RECT 66.000 195.900 66.300 196.500 ;
        RECT 66.700 196.400 67.100 196.500 ;
        RECT 67.900 196.600 68.600 197.000 ;
        RECT 67.900 196.100 68.200 196.600 ;
        RECT 63.900 195.700 66.300 195.900 ;
        RECT 61.400 195.600 66.300 195.700 ;
        RECT 67.000 195.800 68.200 196.100 ;
        RECT 61.400 195.500 64.300 195.600 ;
        RECT 61.400 195.400 64.200 195.500 ;
        RECT 64.600 195.100 65.000 195.200 ;
        RECT 62.500 194.800 65.000 195.100 ;
        RECT 62.500 194.700 62.900 194.800 ;
        RECT 63.800 194.700 64.200 194.800 ;
        RECT 63.300 194.200 63.700 194.300 ;
        RECT 67.000 194.200 67.300 195.800 ;
        RECT 70.200 195.600 70.600 199.900 ;
        RECT 72.300 196.200 72.700 199.900 ;
        RECT 75.500 199.200 75.900 199.900 ;
        RECT 75.000 198.800 75.900 199.200 ;
        RECT 73.000 196.800 73.400 197.200 ;
        RECT 73.100 196.200 73.400 196.800 ;
        RECT 75.500 196.200 75.900 198.800 ;
        RECT 76.200 196.800 76.600 197.200 ;
        RECT 77.400 196.800 78.200 197.200 ;
        RECT 76.300 196.200 76.600 196.800 ;
        RECT 77.800 196.200 78.100 196.800 ;
        RECT 78.500 196.200 78.900 199.900 ;
        RECT 81.000 196.800 81.400 197.200 ;
        RECT 81.000 196.200 81.300 196.800 ;
        RECT 81.700 196.200 82.100 199.900 ;
        RECT 72.300 195.900 72.800 196.200 ;
        RECT 73.100 195.900 73.800 196.200 ;
        RECT 75.500 195.900 76.000 196.200 ;
        RECT 76.300 195.900 77.000 196.200 ;
        RECT 68.500 195.300 70.600 195.600 ;
        RECT 68.500 195.200 68.900 195.300 ;
        RECT 69.300 194.900 69.700 195.000 ;
        RECT 67.800 194.600 69.700 194.900 ;
        RECT 67.800 194.500 68.200 194.600 ;
        RECT 47.900 193.300 49.800 193.600 ;
        RECT 47.900 193.200 48.300 193.300 ;
        RECT 42.200 192.100 42.600 192.500 ;
        RECT 43.000 192.400 43.400 192.800 ;
        RECT 43.900 192.700 44.300 192.800 ;
        RECT 43.900 192.400 45.300 192.700 ;
        RECT 45.000 192.100 45.300 192.400 ;
        RECT 47.000 192.100 47.400 192.500 ;
        RECT 42.200 191.800 43.200 192.100 ;
        RECT 42.800 191.100 43.200 191.800 ;
        RECT 45.000 191.100 45.400 192.100 ;
        RECT 47.000 191.800 47.700 192.100 ;
        RECT 47.100 191.100 47.700 191.800 ;
        RECT 49.400 191.100 49.800 193.300 ;
        RECT 50.300 193.100 50.600 193.800 ;
        RECT 52.200 193.600 52.600 193.800 ;
        RECT 54.900 193.500 55.200 193.800 ;
        RECT 55.700 193.900 56.200 194.100 ;
        RECT 58.200 194.100 58.600 194.200 ;
        RECT 55.700 193.600 57.800 193.900 ;
        RECT 58.200 193.800 59.000 194.100 ;
        RECT 59.700 193.800 61.000 194.200 ;
        RECT 61.800 193.900 67.300 194.200 ;
        RECT 61.800 193.800 62.600 193.900 ;
        RECT 58.600 193.600 59.000 193.800 ;
        RECT 54.900 193.300 55.300 193.500 ;
        RECT 51.100 193.100 52.900 193.300 ;
        RECT 50.200 191.100 50.600 193.100 ;
        RECT 51.000 193.000 53.000 193.100 ;
        RECT 54.900 193.000 55.700 193.300 ;
        RECT 51.000 191.100 51.400 193.000 ;
        RECT 52.600 191.100 53.000 193.000 ;
        RECT 55.300 192.200 55.700 193.000 ;
        RECT 57.500 192.500 57.800 193.600 ;
        RECT 58.300 193.100 60.100 193.300 ;
        RECT 60.600 193.100 60.900 193.800 ;
        RECT 55.300 191.800 56.200 192.200 ;
        RECT 55.300 191.500 55.700 191.800 ;
        RECT 57.400 191.500 57.800 192.500 ;
        RECT 58.200 193.000 60.200 193.100 ;
        RECT 58.200 191.100 58.600 193.000 ;
        RECT 59.800 191.100 60.200 193.000 ;
        RECT 60.600 191.100 61.000 193.100 ;
        RECT 61.400 191.100 61.800 193.500 ;
        RECT 63.900 192.800 64.200 193.900 ;
        RECT 66.700 193.800 67.100 193.900 ;
        RECT 70.200 193.600 70.600 195.300 ;
        RECT 71.800 194.400 72.200 195.200 ;
        RECT 72.500 194.200 72.800 195.900 ;
        RECT 73.400 195.800 73.800 195.900 ;
        RECT 75.000 194.400 75.400 195.200 ;
        RECT 75.700 194.200 76.000 195.900 ;
        RECT 76.600 195.800 77.000 195.900 ;
        RECT 77.400 195.900 78.100 196.200 ;
        RECT 78.400 195.900 78.900 196.200 ;
        RECT 80.600 195.900 81.300 196.200 ;
        RECT 81.600 195.900 82.100 196.200 ;
        RECT 85.100 196.200 85.500 199.900 ;
        RECT 88.300 197.200 88.700 199.900 ;
        RECT 85.800 196.800 86.200 197.200 ;
        RECT 87.800 196.800 88.700 197.200 ;
        RECT 89.000 196.800 89.400 197.200 ;
        RECT 85.900 196.200 86.200 196.800 ;
        RECT 88.300 196.200 88.700 196.800 ;
        RECT 89.100 196.200 89.400 196.800 ;
        RECT 85.100 195.900 85.600 196.200 ;
        RECT 85.900 195.900 86.600 196.200 ;
        RECT 88.300 195.900 88.800 196.200 ;
        RECT 89.100 196.100 89.800 196.200 ;
        RECT 91.000 196.100 91.400 196.200 ;
        RECT 89.100 195.900 91.400 196.100 ;
        RECT 77.400 195.800 77.800 195.900 ;
        RECT 76.600 195.100 76.900 195.800 ;
        RECT 78.400 195.100 78.700 195.900 ;
        RECT 80.600 195.800 81.000 195.900 ;
        RECT 81.600 195.200 81.900 195.900 ;
        RECT 76.600 194.800 78.700 195.100 ;
        RECT 78.400 194.200 78.700 194.800 ;
        RECT 79.000 194.400 79.400 195.200 ;
        RECT 81.400 194.800 81.900 195.200 ;
        RECT 81.600 194.200 81.900 194.800 ;
        RECT 82.200 194.400 82.600 195.200 ;
        RECT 84.600 194.400 85.000 195.200 ;
        RECT 85.300 194.200 85.600 195.900 ;
        RECT 86.200 195.800 86.600 195.900 ;
        RECT 87.800 194.400 88.200 195.200 ;
        RECT 88.500 194.200 88.800 195.900 ;
        RECT 89.400 195.800 91.400 195.900 ;
        RECT 91.800 195.700 92.200 199.900 ;
        RECT 94.000 198.200 94.400 199.900 ;
        RECT 93.400 197.900 94.400 198.200 ;
        RECT 96.200 197.900 96.600 199.900 ;
        RECT 98.300 197.900 98.900 199.900 ;
        RECT 93.400 197.500 93.800 197.900 ;
        RECT 96.200 197.600 96.500 197.900 ;
        RECT 95.100 197.300 96.900 197.600 ;
        RECT 98.200 197.500 98.600 197.900 ;
        RECT 95.100 197.200 95.500 197.300 ;
        RECT 96.500 197.200 96.900 197.300 ;
        RECT 93.400 196.500 93.800 196.600 ;
        RECT 95.700 196.500 96.100 196.600 ;
        RECT 93.400 196.200 96.100 196.500 ;
        RECT 96.400 196.500 97.500 196.800 ;
        RECT 96.400 195.900 96.700 196.500 ;
        RECT 97.100 196.400 97.500 196.500 ;
        RECT 98.300 196.600 99.000 197.000 ;
        RECT 98.300 196.100 98.600 196.600 ;
        RECT 94.300 195.700 96.700 195.900 ;
        RECT 91.800 195.600 96.700 195.700 ;
        RECT 97.400 195.800 98.600 196.100 ;
        RECT 91.800 195.500 94.700 195.600 ;
        RECT 91.800 195.400 94.600 195.500 ;
        RECT 97.400 195.200 97.700 195.800 ;
        RECT 100.600 195.600 101.000 199.900 ;
        RECT 102.700 196.200 103.100 199.900 ;
        RECT 105.900 197.200 106.300 199.900 ;
        RECT 103.400 196.800 103.800 197.200 ;
        RECT 105.400 196.800 106.300 197.200 ;
        RECT 106.600 196.800 107.000 197.200 ;
        RECT 103.500 196.200 103.800 196.800 ;
        RECT 105.900 196.200 106.300 196.800 ;
        RECT 106.700 196.200 107.000 196.800 ;
        RECT 102.700 195.900 103.200 196.200 ;
        RECT 103.500 195.900 104.200 196.200 ;
        RECT 105.900 195.900 106.400 196.200 ;
        RECT 106.700 195.900 107.400 196.200 ;
        RECT 98.900 195.300 101.000 195.600 ;
        RECT 98.900 195.200 99.300 195.300 ;
        RECT 95.000 195.100 95.400 195.200 ;
        RECT 92.900 194.800 95.400 195.100 ;
        RECT 97.400 194.800 97.800 195.200 ;
        RECT 99.700 194.900 100.100 195.000 ;
        RECT 92.900 194.700 93.300 194.800 ;
        RECT 94.200 194.700 94.600 194.800 ;
        RECT 93.700 194.200 94.100 194.300 ;
        RECT 97.400 194.200 97.700 194.800 ;
        RECT 98.200 194.600 100.100 194.900 ;
        RECT 98.200 194.500 98.600 194.600 ;
        RECT 71.000 194.100 71.400 194.200 ;
        RECT 71.000 193.800 71.800 194.100 ;
        RECT 72.500 193.800 73.800 194.200 ;
        RECT 74.200 194.100 74.600 194.200 ;
        RECT 74.200 193.800 75.000 194.100 ;
        RECT 75.700 193.800 77.000 194.200 ;
        RECT 77.400 193.800 78.700 194.200 ;
        RECT 79.800 194.100 80.200 194.200 ;
        RECT 79.400 193.800 80.200 194.100 ;
        RECT 80.600 193.800 81.900 194.200 ;
        RECT 83.000 194.100 83.400 194.200 ;
        RECT 83.800 194.100 84.200 194.200 ;
        RECT 82.600 193.800 84.600 194.100 ;
        RECT 85.300 193.800 86.600 194.200 ;
        RECT 87.000 194.100 87.400 194.200 ;
        RECT 87.000 193.800 87.800 194.100 ;
        RECT 88.500 193.800 89.800 194.200 ;
        RECT 92.200 193.900 97.700 194.200 ;
        RECT 92.200 193.800 93.000 193.900 ;
        RECT 71.400 193.600 71.800 193.800 ;
        RECT 68.700 193.300 70.600 193.600 ;
        RECT 68.700 193.200 69.100 193.300 ;
        RECT 63.000 192.100 63.400 192.500 ;
        RECT 63.800 192.400 64.200 192.800 ;
        RECT 64.700 192.700 65.100 192.800 ;
        RECT 64.700 192.400 66.100 192.700 ;
        RECT 65.800 192.100 66.100 192.400 ;
        RECT 67.800 192.100 68.200 192.500 ;
        RECT 63.000 191.800 64.000 192.100 ;
        RECT 63.600 191.100 64.000 191.800 ;
        RECT 65.800 191.100 66.200 192.100 ;
        RECT 67.800 191.800 68.500 192.100 ;
        RECT 67.900 191.100 68.500 191.800 ;
        RECT 70.200 191.100 70.600 193.300 ;
        RECT 71.100 193.100 72.900 193.300 ;
        RECT 73.400 193.100 73.700 193.800 ;
        RECT 74.600 193.600 75.000 193.800 ;
        RECT 74.300 193.100 76.100 193.300 ;
        RECT 76.600 193.100 76.900 193.800 ;
        RECT 77.500 193.100 77.800 193.800 ;
        RECT 79.400 193.600 79.800 193.800 ;
        RECT 78.300 193.100 80.100 193.300 ;
        RECT 80.700 193.100 81.000 193.800 ;
        RECT 82.600 193.600 83.000 193.800 ;
        RECT 84.200 193.600 84.600 193.800 ;
        RECT 81.500 193.100 83.300 193.300 ;
        RECT 83.900 193.100 85.700 193.300 ;
        RECT 86.200 193.100 86.500 193.800 ;
        RECT 87.400 193.600 87.800 193.800 ;
        RECT 87.100 193.100 88.900 193.300 ;
        RECT 89.400 193.100 89.700 193.800 ;
        RECT 71.000 193.000 73.000 193.100 ;
        RECT 71.000 191.100 71.400 193.000 ;
        RECT 72.600 191.100 73.000 193.000 ;
        RECT 73.400 191.100 73.800 193.100 ;
        RECT 74.200 193.000 76.200 193.100 ;
        RECT 74.200 191.100 74.600 193.000 ;
        RECT 75.800 191.100 76.200 193.000 ;
        RECT 76.600 191.100 77.000 193.100 ;
        RECT 77.400 191.100 77.800 193.100 ;
        RECT 78.200 193.000 80.200 193.100 ;
        RECT 78.200 191.100 78.600 193.000 ;
        RECT 79.800 191.100 80.200 193.000 ;
        RECT 80.600 191.100 81.000 193.100 ;
        RECT 81.400 193.000 83.400 193.100 ;
        RECT 81.400 191.100 81.800 193.000 ;
        RECT 83.000 191.100 83.400 193.000 ;
        RECT 83.800 193.000 85.800 193.100 ;
        RECT 83.800 191.100 84.200 193.000 ;
        RECT 85.400 191.100 85.800 193.000 ;
        RECT 86.200 191.100 86.600 193.100 ;
        RECT 87.000 193.000 89.000 193.100 ;
        RECT 87.000 191.100 87.400 193.000 ;
        RECT 88.600 191.100 89.000 193.000 ;
        RECT 89.400 191.100 89.800 193.100 ;
        RECT 91.800 191.100 92.200 193.500 ;
        RECT 94.300 192.800 94.600 193.900 ;
        RECT 97.100 193.800 97.500 193.900 ;
        RECT 100.600 193.600 101.000 195.300 ;
        RECT 102.200 194.400 102.600 195.200 ;
        RECT 102.900 194.200 103.200 195.900 ;
        RECT 103.800 195.800 104.200 195.900 ;
        RECT 105.400 194.400 105.800 195.200 ;
        RECT 106.100 194.200 106.400 195.900 ;
        RECT 107.000 195.800 107.400 195.900 ;
        RECT 107.800 195.700 108.200 199.900 ;
        RECT 110.000 198.200 110.400 199.900 ;
        RECT 109.400 197.900 110.400 198.200 ;
        RECT 112.200 197.900 112.600 199.900 ;
        RECT 114.300 197.900 114.900 199.900 ;
        RECT 109.400 197.500 109.800 197.900 ;
        RECT 112.200 197.600 112.500 197.900 ;
        RECT 111.100 197.300 112.900 197.600 ;
        RECT 114.200 197.500 114.600 197.900 ;
        RECT 111.100 197.200 111.500 197.300 ;
        RECT 112.500 197.200 112.900 197.300 ;
        RECT 109.400 196.500 109.800 196.600 ;
        RECT 111.700 196.500 112.100 196.600 ;
        RECT 109.400 196.200 112.100 196.500 ;
        RECT 112.400 196.500 113.500 196.800 ;
        RECT 112.400 195.900 112.700 196.500 ;
        RECT 113.100 196.400 113.500 196.500 ;
        RECT 114.300 196.600 115.000 197.000 ;
        RECT 114.300 196.100 114.600 196.600 ;
        RECT 110.300 195.700 112.700 195.900 ;
        RECT 107.800 195.600 112.700 195.700 ;
        RECT 113.400 195.800 114.600 196.100 ;
        RECT 107.800 195.500 110.700 195.600 ;
        RECT 107.800 195.400 110.600 195.500 ;
        RECT 111.000 195.100 111.400 195.200 ;
        RECT 108.900 194.800 111.400 195.100 ;
        RECT 108.900 194.700 109.300 194.800 ;
        RECT 110.200 194.700 110.600 194.800 ;
        RECT 109.700 194.200 110.100 194.300 ;
        RECT 113.400 194.200 113.700 195.800 ;
        RECT 116.600 195.600 117.000 199.900 ;
        RECT 114.900 195.300 117.000 195.600 ;
        RECT 117.400 195.700 117.800 199.900 ;
        RECT 119.600 198.200 120.000 199.900 ;
        RECT 119.000 197.900 120.000 198.200 ;
        RECT 121.800 197.900 122.200 199.900 ;
        RECT 123.900 197.900 124.500 199.900 ;
        RECT 119.000 197.500 119.400 197.900 ;
        RECT 121.800 197.600 122.100 197.900 ;
        RECT 120.700 197.300 122.500 197.600 ;
        RECT 123.800 197.500 124.200 197.900 ;
        RECT 120.700 197.200 121.100 197.300 ;
        RECT 122.100 197.200 122.500 197.300 ;
        RECT 119.000 196.500 119.400 196.600 ;
        RECT 121.300 196.500 121.700 196.600 ;
        RECT 119.000 196.200 121.700 196.500 ;
        RECT 122.000 196.500 123.100 196.800 ;
        RECT 122.000 195.900 122.300 196.500 ;
        RECT 122.700 196.400 123.100 196.500 ;
        RECT 123.900 196.600 124.600 197.000 ;
        RECT 123.900 196.100 124.200 196.600 ;
        RECT 119.900 195.700 122.300 195.900 ;
        RECT 117.400 195.600 122.300 195.700 ;
        RECT 123.000 195.800 124.200 196.100 ;
        RECT 117.400 195.500 120.300 195.600 ;
        RECT 117.400 195.400 120.200 195.500 ;
        RECT 114.900 195.200 115.300 195.300 ;
        RECT 115.700 194.900 116.100 195.000 ;
        RECT 114.200 194.600 116.100 194.900 ;
        RECT 114.200 194.500 114.600 194.600 ;
        RECT 101.400 194.100 101.800 194.200 ;
        RECT 101.400 193.800 102.200 194.100 ;
        RECT 102.900 193.800 104.200 194.200 ;
        RECT 104.600 194.100 105.000 194.200 ;
        RECT 104.600 193.800 105.400 194.100 ;
        RECT 106.100 193.800 107.400 194.200 ;
        RECT 108.200 193.900 113.700 194.200 ;
        RECT 108.200 193.800 109.000 193.900 ;
        RECT 101.800 193.600 102.200 193.800 ;
        RECT 99.100 193.300 101.000 193.600 ;
        RECT 99.100 193.200 99.500 193.300 ;
        RECT 93.400 192.100 93.800 192.500 ;
        RECT 94.200 192.400 94.600 192.800 ;
        RECT 95.100 192.700 95.500 192.800 ;
        RECT 95.100 192.400 96.500 192.700 ;
        RECT 96.200 192.100 96.500 192.400 ;
        RECT 98.200 192.100 98.600 192.500 ;
        RECT 93.400 191.800 94.400 192.100 ;
        RECT 94.000 191.100 94.400 191.800 ;
        RECT 96.200 191.100 96.600 192.100 ;
        RECT 98.200 191.800 98.900 192.100 ;
        RECT 98.300 191.100 98.900 191.800 ;
        RECT 100.600 191.100 101.000 193.300 ;
        RECT 101.500 193.100 103.300 193.300 ;
        RECT 103.800 193.100 104.100 193.800 ;
        RECT 105.000 193.600 105.400 193.800 ;
        RECT 104.700 193.100 106.500 193.300 ;
        RECT 107.000 193.100 107.300 193.800 ;
        RECT 101.400 193.000 103.400 193.100 ;
        RECT 101.400 191.100 101.800 193.000 ;
        RECT 103.000 191.100 103.400 193.000 ;
        RECT 103.800 191.100 104.200 193.100 ;
        RECT 104.600 193.000 106.600 193.100 ;
        RECT 104.600 191.100 105.000 193.000 ;
        RECT 106.200 191.100 106.600 193.000 ;
        RECT 107.000 191.100 107.400 193.100 ;
        RECT 107.800 191.100 108.200 193.500 ;
        RECT 110.300 192.800 110.600 193.900 ;
        RECT 113.100 193.800 113.500 193.900 ;
        RECT 116.600 193.600 117.000 195.300 ;
        RECT 120.600 195.100 121.000 195.200 ;
        RECT 121.400 195.100 121.800 195.200 ;
        RECT 118.500 194.800 121.800 195.100 ;
        RECT 118.500 194.700 118.900 194.800 ;
        RECT 119.300 194.200 119.700 194.300 ;
        RECT 123.000 194.200 123.300 195.800 ;
        RECT 126.200 195.600 126.600 199.900 ;
        RECT 128.300 197.200 128.700 199.900 ;
        RECT 127.800 196.800 128.700 197.200 ;
        RECT 129.000 196.800 129.400 197.200 ;
        RECT 128.300 196.200 128.700 196.800 ;
        RECT 129.100 196.200 129.400 196.800 ;
        RECT 130.600 196.800 131.000 197.200 ;
        RECT 130.600 196.200 130.900 196.800 ;
        RECT 131.300 196.200 131.700 199.900 ;
        RECT 128.300 195.900 128.800 196.200 ;
        RECT 129.100 195.900 129.800 196.200 ;
        RECT 124.500 195.300 126.600 195.600 ;
        RECT 124.500 195.200 124.900 195.300 ;
        RECT 125.300 194.900 125.700 195.000 ;
        RECT 123.800 194.600 125.700 194.900 ;
        RECT 123.800 194.500 124.200 194.600 ;
        RECT 117.800 193.900 123.300 194.200 ;
        RECT 117.800 193.800 118.600 193.900 ;
        RECT 115.100 193.300 117.000 193.600 ;
        RECT 115.100 193.200 115.500 193.300 ;
        RECT 109.400 192.100 109.800 192.500 ;
        RECT 110.200 192.400 110.600 192.800 ;
        RECT 111.100 192.700 111.500 192.800 ;
        RECT 111.100 192.400 112.500 192.700 ;
        RECT 112.200 192.100 112.500 192.400 ;
        RECT 114.200 192.100 114.600 192.500 ;
        RECT 109.400 191.800 110.400 192.100 ;
        RECT 110.000 191.100 110.400 191.800 ;
        RECT 112.200 191.100 112.600 192.100 ;
        RECT 114.200 191.800 114.900 192.100 ;
        RECT 114.300 191.100 114.900 191.800 ;
        RECT 116.600 191.100 117.000 193.300 ;
        RECT 117.400 191.100 117.800 193.500 ;
        RECT 119.900 193.200 120.200 193.900 ;
        RECT 122.700 193.800 123.100 193.900 ;
        RECT 126.200 193.600 126.600 195.300 ;
        RECT 127.800 194.400 128.200 195.200 ;
        RECT 128.500 194.200 128.800 195.900 ;
        RECT 129.400 195.800 129.800 195.900 ;
        RECT 130.200 195.900 130.900 196.200 ;
        RECT 131.200 195.900 131.700 196.200 ;
        RECT 134.700 196.200 135.100 199.900 ;
        RECT 135.400 196.800 136.200 197.200 ;
        RECT 137.000 196.800 137.400 197.200 ;
        RECT 135.500 196.200 135.800 196.800 ;
        RECT 137.000 196.200 137.300 196.800 ;
        RECT 137.700 196.200 138.100 199.900 ;
        RECT 134.700 195.900 135.200 196.200 ;
        RECT 135.500 195.900 136.200 196.200 ;
        RECT 130.200 195.800 130.600 195.900 ;
        RECT 129.400 195.100 129.700 195.800 ;
        RECT 131.200 195.100 131.500 195.900 ;
        RECT 129.400 194.800 131.500 195.100 ;
        RECT 131.200 194.200 131.500 194.800 ;
        RECT 131.800 195.100 132.200 195.200 ;
        RECT 134.200 195.100 134.600 195.200 ;
        RECT 131.800 194.800 134.600 195.100 ;
        RECT 131.800 194.400 132.200 194.800 ;
        RECT 134.200 194.400 134.600 194.800 ;
        RECT 134.900 195.100 135.200 195.900 ;
        RECT 135.800 195.800 136.200 195.900 ;
        RECT 136.600 195.900 137.300 196.200 ;
        RECT 136.600 195.800 137.000 195.900 ;
        RECT 137.600 195.800 138.600 196.200 ;
        RECT 136.600 195.100 136.900 195.800 ;
        RECT 134.900 194.800 136.900 195.100 ;
        RECT 134.900 194.200 135.200 194.800 ;
        RECT 137.600 194.200 137.900 195.800 ;
        RECT 141.400 195.600 141.800 199.900 ;
        RECT 143.500 197.900 144.100 199.900 ;
        RECT 145.800 197.900 146.200 199.900 ;
        RECT 148.000 198.200 148.400 199.900 ;
        RECT 148.000 197.900 149.000 198.200 ;
        RECT 143.800 197.500 144.200 197.900 ;
        RECT 145.900 197.600 146.200 197.900 ;
        RECT 145.500 197.300 147.300 197.600 ;
        RECT 148.600 197.500 149.000 197.900 ;
        RECT 145.500 197.200 145.900 197.300 ;
        RECT 146.900 197.200 147.300 197.300 ;
        RECT 143.400 196.600 144.100 197.000 ;
        RECT 143.800 196.100 144.100 196.600 ;
        RECT 144.900 196.500 146.000 196.800 ;
        RECT 144.900 196.400 145.300 196.500 ;
        RECT 143.800 195.800 145.000 196.100 ;
        RECT 141.400 195.300 143.500 195.600 ;
        RECT 138.200 194.400 138.600 195.200 ;
        RECT 127.000 194.100 127.400 194.200 ;
        RECT 127.000 193.800 127.800 194.100 ;
        RECT 128.500 193.800 129.800 194.200 ;
        RECT 130.200 193.800 131.500 194.200 ;
        RECT 132.600 194.100 133.000 194.200 ;
        RECT 133.400 194.100 133.800 194.200 ;
        RECT 132.200 193.800 134.200 194.100 ;
        RECT 134.900 193.800 136.200 194.200 ;
        RECT 136.600 193.800 137.900 194.200 ;
        RECT 139.000 194.100 139.400 194.200 ;
        RECT 138.600 193.800 139.400 194.100 ;
        RECT 127.400 193.600 127.800 193.800 ;
        RECT 124.700 193.300 126.600 193.600 ;
        RECT 124.700 193.200 125.100 193.300 ;
        RECT 119.000 192.100 119.400 192.500 ;
        RECT 119.800 192.400 120.200 193.200 ;
        RECT 120.700 192.700 121.100 192.800 ;
        RECT 120.700 192.400 122.100 192.700 ;
        RECT 121.800 192.100 122.100 192.400 ;
        RECT 123.800 192.100 124.200 192.500 ;
        RECT 119.000 191.800 120.000 192.100 ;
        RECT 119.600 191.100 120.000 191.800 ;
        RECT 121.800 191.100 122.200 192.100 ;
        RECT 123.800 191.800 124.500 192.100 ;
        RECT 123.900 191.100 124.500 191.800 ;
        RECT 126.200 191.100 126.600 193.300 ;
        RECT 127.100 193.100 128.900 193.300 ;
        RECT 129.400 193.100 129.700 193.800 ;
        RECT 130.300 193.100 130.600 193.800 ;
        RECT 132.200 193.600 132.600 193.800 ;
        RECT 133.800 193.600 134.200 193.800 ;
        RECT 131.100 193.100 132.900 193.300 ;
        RECT 133.500 193.100 135.300 193.300 ;
        RECT 135.800 193.100 136.100 193.800 ;
        RECT 136.700 193.100 137.000 193.800 ;
        RECT 138.600 193.600 139.000 193.800 ;
        RECT 141.400 193.600 141.800 195.300 ;
        RECT 143.100 195.200 143.500 195.300 ;
        RECT 142.300 194.900 142.700 195.000 ;
        RECT 142.300 194.600 144.200 194.900 ;
        RECT 143.800 194.500 144.200 194.600 ;
        RECT 144.700 194.200 145.000 195.800 ;
        RECT 145.700 195.900 146.000 196.500 ;
        RECT 146.300 196.500 146.700 196.600 ;
        RECT 148.600 196.500 149.000 196.600 ;
        RECT 146.300 196.200 149.000 196.500 ;
        RECT 145.700 195.700 148.100 195.900 ;
        RECT 150.200 195.700 150.600 199.900 ;
        RECT 145.700 195.600 150.600 195.700 ;
        RECT 147.700 195.500 150.600 195.600 ;
        RECT 147.800 195.400 150.600 195.500 ;
        RECT 151.000 195.600 151.400 199.900 ;
        RECT 153.100 197.900 153.700 199.900 ;
        RECT 155.400 197.900 155.800 199.900 ;
        RECT 157.600 198.200 158.000 199.900 ;
        RECT 157.600 197.900 158.600 198.200 ;
        RECT 153.400 197.500 153.800 197.900 ;
        RECT 155.500 197.600 155.800 197.900 ;
        RECT 155.100 197.300 156.900 197.600 ;
        RECT 158.200 197.500 158.600 197.900 ;
        RECT 155.100 197.200 155.500 197.300 ;
        RECT 156.500 197.200 156.900 197.300 ;
        RECT 153.000 196.600 153.700 197.000 ;
        RECT 153.400 196.100 153.700 196.600 ;
        RECT 154.500 196.500 155.600 196.800 ;
        RECT 154.500 196.400 154.900 196.500 ;
        RECT 153.400 195.800 154.600 196.100 ;
        RECT 151.000 195.300 153.100 195.600 ;
        RECT 147.000 195.100 147.400 195.200 ;
        RECT 147.000 194.800 149.500 195.100 ;
        RECT 149.100 194.700 149.500 194.800 ;
        RECT 148.300 194.200 148.700 194.300 ;
        RECT 144.700 193.900 150.200 194.200 ;
        RECT 144.900 193.800 145.300 193.900 ;
        RECT 141.400 193.300 143.300 193.600 ;
        RECT 137.500 193.100 139.300 193.300 ;
        RECT 127.000 193.000 129.000 193.100 ;
        RECT 127.000 191.100 127.400 193.000 ;
        RECT 128.600 191.100 129.000 193.000 ;
        RECT 129.400 191.100 129.800 193.100 ;
        RECT 130.200 191.100 130.600 193.100 ;
        RECT 131.000 193.000 133.000 193.100 ;
        RECT 131.000 191.100 131.400 193.000 ;
        RECT 132.600 191.100 133.000 193.000 ;
        RECT 133.400 193.000 135.400 193.100 ;
        RECT 133.400 191.100 133.800 193.000 ;
        RECT 135.000 191.100 135.400 193.000 ;
        RECT 135.800 191.100 136.200 193.100 ;
        RECT 136.600 191.100 137.000 193.100 ;
        RECT 137.400 193.000 139.400 193.100 ;
        RECT 137.400 191.100 137.800 193.000 ;
        RECT 139.000 191.100 139.400 193.000 ;
        RECT 141.400 191.100 141.800 193.300 ;
        RECT 142.900 193.200 143.300 193.300 ;
        RECT 147.800 192.800 148.100 193.900 ;
        RECT 149.400 193.800 150.200 193.900 ;
        RECT 151.000 193.600 151.400 195.300 ;
        RECT 152.700 195.200 153.100 195.300 ;
        RECT 151.900 194.900 152.300 195.000 ;
        RECT 151.900 194.600 153.800 194.900 ;
        RECT 153.400 194.500 153.800 194.600 ;
        RECT 154.300 194.200 154.600 195.800 ;
        RECT 155.300 195.900 155.600 196.500 ;
        RECT 155.900 196.500 156.300 196.600 ;
        RECT 158.200 196.500 158.600 196.600 ;
        RECT 155.900 196.200 158.600 196.500 ;
        RECT 155.300 195.700 157.700 195.900 ;
        RECT 159.800 195.700 160.200 199.900 ;
        RECT 161.900 196.200 162.300 199.900 ;
        RECT 162.600 196.800 163.000 197.200 ;
        RECT 162.700 196.200 163.000 196.800 ;
        RECT 161.900 195.900 162.400 196.200 ;
        RECT 162.700 195.900 163.400 196.200 ;
        RECT 155.300 195.600 160.200 195.700 ;
        RECT 157.300 195.500 160.200 195.600 ;
        RECT 157.400 195.400 160.200 195.500 ;
        RECT 156.600 195.100 157.000 195.200 ;
        RECT 156.600 194.800 159.100 195.100 ;
        RECT 157.400 194.700 157.800 194.800 ;
        RECT 158.700 194.700 159.100 194.800 ;
        RECT 161.400 194.400 161.800 195.200 ;
        RECT 157.900 194.200 158.300 194.300 ;
        RECT 162.100 194.200 162.400 195.900 ;
        RECT 163.000 195.800 163.400 195.900 ;
        RECT 163.800 195.800 164.200 196.600 ;
        RECT 163.000 195.100 163.300 195.800 ;
        RECT 164.600 195.100 165.000 199.900 ;
        RECT 163.000 194.800 165.000 195.100 ;
        RECT 154.300 193.900 159.800 194.200 ;
        RECT 154.500 193.800 154.900 193.900 ;
        RECT 146.900 192.700 147.300 192.800 ;
        RECT 143.800 192.100 144.200 192.500 ;
        RECT 145.900 192.400 147.300 192.700 ;
        RECT 147.800 192.400 148.200 192.800 ;
        RECT 145.900 192.100 146.200 192.400 ;
        RECT 148.600 192.100 149.000 192.500 ;
        RECT 143.500 191.800 144.200 192.100 ;
        RECT 143.500 191.100 144.100 191.800 ;
        RECT 145.800 191.100 146.200 192.100 ;
        RECT 148.000 191.800 149.000 192.100 ;
        RECT 148.000 191.100 148.400 191.800 ;
        RECT 150.200 191.100 150.600 193.500 ;
        RECT 151.000 193.300 152.900 193.600 ;
        RECT 151.000 191.100 151.400 193.300 ;
        RECT 152.500 193.200 152.900 193.300 ;
        RECT 157.400 192.800 157.700 193.900 ;
        RECT 159.000 193.800 159.800 193.900 ;
        RECT 160.600 194.100 161.000 194.200 ;
        RECT 160.600 193.800 161.400 194.100 ;
        RECT 162.100 193.800 163.400 194.200 ;
        RECT 161.000 193.600 161.400 193.800 ;
        RECT 156.500 192.700 156.900 192.800 ;
        RECT 153.400 192.100 153.800 192.500 ;
        RECT 155.500 192.400 156.900 192.700 ;
        RECT 157.400 192.400 157.800 192.800 ;
        RECT 155.500 192.100 155.800 192.400 ;
        RECT 158.200 192.100 158.600 192.500 ;
        RECT 153.100 191.800 153.800 192.100 ;
        RECT 153.100 191.100 153.700 191.800 ;
        RECT 155.400 191.100 155.800 192.100 ;
        RECT 157.600 191.800 158.600 192.100 ;
        RECT 157.600 191.100 158.000 191.800 ;
        RECT 159.800 191.100 160.200 193.500 ;
        RECT 160.700 193.100 162.500 193.300 ;
        RECT 163.000 193.100 163.300 193.800 ;
        RECT 164.600 193.100 165.000 194.800 ;
        RECT 166.200 195.600 166.600 199.900 ;
        RECT 168.300 197.900 168.900 199.900 ;
        RECT 170.600 197.900 171.000 199.900 ;
        RECT 172.800 198.200 173.200 199.900 ;
        RECT 172.800 197.900 173.800 198.200 ;
        RECT 168.600 197.500 169.000 197.900 ;
        RECT 170.700 197.600 171.000 197.900 ;
        RECT 170.300 197.300 172.100 197.600 ;
        RECT 173.400 197.500 173.800 197.900 ;
        RECT 170.300 197.200 170.700 197.300 ;
        RECT 171.700 197.200 172.100 197.300 ;
        RECT 168.200 196.600 168.900 197.000 ;
        RECT 168.600 196.100 168.900 196.600 ;
        RECT 169.700 196.500 170.800 196.800 ;
        RECT 169.700 196.400 170.100 196.500 ;
        RECT 168.600 195.800 169.800 196.100 ;
        RECT 166.200 195.300 168.300 195.600 ;
        RECT 165.400 194.100 165.800 194.200 ;
        RECT 166.200 194.100 166.600 195.300 ;
        RECT 167.900 195.200 168.300 195.300 ;
        RECT 167.100 194.900 167.500 195.000 ;
        RECT 167.100 194.600 169.000 194.900 ;
        RECT 168.600 194.500 169.000 194.600 ;
        RECT 165.400 193.800 166.600 194.100 ;
        RECT 169.500 194.200 169.800 195.800 ;
        RECT 170.500 195.900 170.800 196.500 ;
        RECT 171.100 196.500 171.500 196.600 ;
        RECT 173.400 196.500 173.800 196.600 ;
        RECT 171.100 196.200 173.800 196.500 ;
        RECT 170.500 195.700 172.900 195.900 ;
        RECT 175.000 195.700 175.400 199.900 ;
        RECT 177.100 199.200 177.500 199.900 ;
        RECT 176.600 198.800 177.500 199.200 ;
        RECT 177.100 196.200 177.500 198.800 ;
        RECT 177.800 196.800 178.200 197.200 ;
        RECT 177.900 196.200 178.200 196.800 ;
        RECT 177.100 195.900 177.600 196.200 ;
        RECT 177.900 195.900 178.600 196.200 ;
        RECT 170.500 195.600 175.400 195.700 ;
        RECT 172.500 195.500 175.400 195.600 ;
        RECT 172.600 195.400 175.400 195.500 ;
        RECT 171.000 195.100 171.400 195.200 ;
        RECT 171.800 195.100 172.200 195.200 ;
        RECT 171.000 194.800 174.300 195.100 ;
        RECT 173.900 194.700 174.300 194.800 ;
        RECT 176.600 194.400 177.000 195.200 ;
        RECT 173.100 194.200 173.500 194.300 ;
        RECT 177.300 194.200 177.600 195.900 ;
        RECT 178.200 195.800 178.600 195.900 ;
        RECT 179.000 195.800 179.400 196.600 ;
        RECT 178.200 195.100 178.500 195.800 ;
        RECT 179.800 195.100 180.200 199.900 ;
        RECT 183.300 196.400 183.700 199.900 ;
        RECT 185.400 197.500 185.800 199.500 ;
        RECT 182.900 196.100 183.700 196.400 ;
        RECT 178.200 194.800 180.200 195.100 ;
        RECT 182.200 194.800 182.600 195.600 ;
        RECT 169.500 193.900 175.000 194.200 ;
        RECT 169.700 193.800 170.100 193.900 ;
        RECT 171.000 193.800 171.400 193.900 ;
        RECT 165.400 193.400 165.800 193.800 ;
        RECT 166.200 193.600 166.600 193.800 ;
        RECT 160.600 193.000 162.600 193.100 ;
        RECT 160.600 191.100 161.000 193.000 ;
        RECT 162.200 191.100 162.600 193.000 ;
        RECT 163.000 191.100 163.400 193.100 ;
        RECT 164.100 192.800 165.000 193.100 ;
        RECT 166.200 193.300 168.100 193.600 ;
        RECT 164.100 191.100 164.500 192.800 ;
        RECT 166.200 191.100 166.600 193.300 ;
        RECT 167.700 193.200 168.100 193.300 ;
        RECT 172.600 192.800 172.900 193.900 ;
        RECT 174.200 193.800 175.000 193.900 ;
        RECT 175.800 194.100 176.200 194.200 ;
        RECT 175.800 193.800 176.600 194.100 ;
        RECT 177.300 193.800 178.600 194.200 ;
        RECT 176.200 193.600 176.600 193.800 ;
        RECT 171.700 192.700 172.100 192.800 ;
        RECT 168.600 192.100 169.000 192.500 ;
        RECT 170.700 192.400 172.100 192.700 ;
        RECT 172.600 192.400 173.000 192.800 ;
        RECT 170.700 192.100 171.000 192.400 ;
        RECT 173.400 192.100 173.800 192.500 ;
        RECT 168.300 191.800 169.000 192.100 ;
        RECT 168.300 191.100 168.900 191.800 ;
        RECT 170.600 191.100 171.000 192.100 ;
        RECT 172.800 191.800 173.800 192.100 ;
        RECT 172.800 191.100 173.200 191.800 ;
        RECT 175.000 191.100 175.400 193.500 ;
        RECT 175.900 193.100 177.700 193.300 ;
        RECT 178.200 193.100 178.500 193.800 ;
        RECT 179.800 193.100 180.200 194.800 ;
        RECT 182.900 194.200 183.200 196.100 ;
        RECT 185.500 195.800 185.800 197.500 ;
        RECT 187.500 196.200 187.900 199.900 ;
        RECT 188.200 196.800 188.600 197.200 ;
        RECT 188.300 196.200 188.600 196.800 ;
        RECT 187.500 195.900 188.000 196.200 ;
        RECT 188.300 195.900 189.000 196.200 ;
        RECT 183.900 195.500 185.800 195.800 ;
        RECT 183.900 194.500 184.200 195.500 ;
        RECT 180.600 193.400 181.000 194.200 ;
        RECT 182.200 193.800 183.200 194.200 ;
        RECT 183.500 194.100 184.200 194.500 ;
        RECT 184.600 194.400 185.000 195.200 ;
        RECT 185.400 194.400 185.800 195.200 ;
        RECT 187.000 194.400 187.400 195.200 ;
        RECT 187.700 194.200 188.000 195.900 ;
        RECT 188.600 195.800 189.000 195.900 ;
        RECT 189.400 195.800 189.800 196.600 ;
        RECT 188.600 195.100 188.900 195.800 ;
        RECT 190.200 195.100 190.600 199.900 ;
        RECT 192.600 197.100 193.000 197.200 ;
        RECT 193.400 197.100 193.800 199.900 ;
        RECT 195.500 197.900 196.100 199.900 ;
        RECT 197.800 197.900 198.200 199.900 ;
        RECT 200.000 198.200 200.400 199.900 ;
        RECT 200.000 197.900 201.000 198.200 ;
        RECT 195.800 197.500 196.200 197.900 ;
        RECT 197.900 197.600 198.200 197.900 ;
        RECT 197.500 197.300 199.300 197.600 ;
        RECT 200.600 197.500 201.000 197.900 ;
        RECT 197.500 197.200 197.900 197.300 ;
        RECT 198.900 197.200 199.300 197.300 ;
        RECT 192.600 196.800 193.800 197.100 ;
        RECT 188.600 194.800 190.600 195.100 ;
        RECT 182.900 193.500 183.200 193.800 ;
        RECT 183.700 193.900 184.200 194.100 ;
        RECT 186.200 194.100 186.600 194.200 ;
        RECT 187.700 194.100 189.000 194.200 ;
        RECT 189.400 194.100 189.800 194.200 ;
        RECT 183.700 193.600 185.800 193.900 ;
        RECT 186.200 193.800 187.000 194.100 ;
        RECT 187.700 193.800 189.800 194.100 ;
        RECT 186.600 193.600 187.000 193.800 ;
        RECT 175.800 193.000 177.800 193.100 ;
        RECT 175.800 191.100 176.200 193.000 ;
        RECT 177.400 191.100 177.800 193.000 ;
        RECT 178.200 191.100 178.600 193.100 ;
        RECT 179.300 192.800 180.200 193.100 ;
        RECT 182.900 193.300 183.300 193.500 ;
        RECT 182.900 193.000 183.700 193.300 ;
        RECT 179.300 191.100 179.700 192.800 ;
        RECT 183.300 192.200 183.700 193.000 ;
        RECT 185.500 192.500 185.800 193.600 ;
        RECT 186.300 193.100 188.100 193.300 ;
        RECT 188.600 193.100 188.900 193.800 ;
        RECT 190.200 193.100 190.600 194.800 ;
        RECT 193.400 195.600 193.800 196.800 ;
        RECT 195.400 196.600 196.100 197.000 ;
        RECT 195.800 196.100 196.100 196.600 ;
        RECT 196.900 196.500 198.000 196.800 ;
        RECT 196.900 196.400 197.300 196.500 ;
        RECT 195.800 195.800 197.000 196.100 ;
        RECT 193.400 195.300 195.500 195.600 ;
        RECT 191.000 194.100 191.400 194.200 ;
        RECT 192.600 194.100 193.000 194.200 ;
        RECT 191.000 193.800 193.000 194.100 ;
        RECT 191.000 193.400 191.400 193.800 ;
        RECT 193.400 193.600 193.800 195.300 ;
        RECT 195.100 195.200 195.500 195.300 ;
        RECT 196.700 195.200 197.000 195.800 ;
        RECT 197.700 195.900 198.000 196.500 ;
        RECT 198.300 196.500 198.700 196.600 ;
        RECT 200.600 196.500 201.000 196.600 ;
        RECT 198.300 196.200 201.000 196.500 ;
        RECT 197.700 195.700 200.100 195.900 ;
        RECT 202.200 195.700 202.600 199.900 ;
        RECT 204.300 196.200 204.700 199.900 ;
        RECT 205.000 196.800 205.400 197.200 ;
        RECT 205.100 196.200 205.400 196.800 ;
        RECT 204.300 195.900 204.800 196.200 ;
        RECT 205.100 195.900 205.800 196.200 ;
        RECT 197.700 195.600 202.600 195.700 ;
        RECT 199.700 195.500 202.600 195.600 ;
        RECT 199.800 195.400 202.600 195.500 ;
        RECT 194.300 194.900 194.700 195.000 ;
        RECT 194.300 194.600 196.200 194.900 ;
        RECT 196.600 194.800 197.000 195.200 ;
        RECT 199.000 195.100 199.400 195.200 ;
        RECT 199.000 194.800 201.500 195.100 ;
        RECT 195.800 194.500 196.200 194.600 ;
        RECT 196.700 194.200 197.000 194.800 ;
        RECT 201.100 194.700 201.500 194.800 ;
        RECT 203.800 194.400 204.200 195.200 ;
        RECT 200.300 194.200 200.700 194.300 ;
        RECT 204.500 194.200 204.800 195.900 ;
        RECT 205.400 195.800 205.800 195.900 ;
        RECT 206.200 195.800 206.600 196.600 ;
        RECT 205.400 195.100 205.700 195.800 ;
        RECT 207.000 195.100 207.400 199.900 ;
        RECT 207.800 197.100 208.200 197.200 ;
        RECT 208.600 197.100 209.000 199.900 ;
        RECT 210.700 197.900 211.300 199.900 ;
        RECT 213.000 197.900 213.400 199.900 ;
        RECT 215.200 198.200 215.600 199.900 ;
        RECT 215.200 197.900 216.200 198.200 ;
        RECT 211.000 197.500 211.400 197.900 ;
        RECT 213.100 197.600 213.400 197.900 ;
        RECT 212.700 197.300 214.500 197.600 ;
        RECT 215.800 197.500 216.200 197.900 ;
        RECT 212.700 197.200 213.100 197.300 ;
        RECT 214.100 197.200 214.500 197.300 ;
        RECT 207.800 196.800 209.000 197.100 ;
        RECT 205.400 194.800 207.400 195.100 ;
        RECT 196.700 193.900 202.200 194.200 ;
        RECT 196.900 193.800 197.300 193.900 ;
        RECT 183.300 191.800 184.200 192.200 ;
        RECT 183.300 191.500 183.700 191.800 ;
        RECT 185.400 191.500 185.800 192.500 ;
        RECT 186.200 193.000 188.200 193.100 ;
        RECT 186.200 191.100 186.600 193.000 ;
        RECT 187.800 191.100 188.200 193.000 ;
        RECT 188.600 191.100 189.000 193.100 ;
        RECT 189.700 192.800 190.600 193.100 ;
        RECT 193.400 193.300 195.300 193.600 ;
        RECT 189.700 191.100 190.100 192.800 ;
        RECT 193.400 191.100 193.800 193.300 ;
        RECT 194.900 193.200 195.300 193.300 ;
        RECT 199.800 192.800 200.100 193.900 ;
        RECT 201.400 193.800 202.200 193.900 ;
        RECT 203.000 194.100 203.400 194.200 ;
        RECT 203.000 193.800 203.800 194.100 ;
        RECT 204.500 193.800 205.800 194.200 ;
        RECT 203.400 193.600 203.800 193.800 ;
        RECT 198.900 192.700 199.300 192.800 ;
        RECT 195.800 192.100 196.200 192.500 ;
        RECT 197.900 192.400 199.300 192.700 ;
        RECT 199.800 192.400 200.200 192.800 ;
        RECT 197.900 192.100 198.200 192.400 ;
        RECT 200.600 192.100 201.000 192.500 ;
        RECT 195.500 191.800 196.200 192.100 ;
        RECT 195.500 191.100 196.100 191.800 ;
        RECT 197.800 191.100 198.200 192.100 ;
        RECT 200.000 191.800 201.000 192.100 ;
        RECT 200.000 191.100 200.400 191.800 ;
        RECT 202.200 191.100 202.600 193.500 ;
        RECT 203.100 193.100 204.900 193.300 ;
        RECT 205.400 193.100 205.700 193.800 ;
        RECT 207.000 193.100 207.400 194.800 ;
        RECT 208.600 195.600 209.000 196.800 ;
        RECT 210.600 196.600 211.300 197.000 ;
        RECT 211.000 196.100 211.300 196.600 ;
        RECT 212.100 196.500 213.200 196.800 ;
        RECT 212.100 196.400 212.500 196.500 ;
        RECT 211.000 195.800 212.200 196.100 ;
        RECT 208.600 195.300 210.700 195.600 ;
        RECT 207.800 193.400 208.200 194.200 ;
        RECT 208.600 193.600 209.000 195.300 ;
        RECT 210.300 195.200 210.700 195.300 ;
        RECT 211.900 195.200 212.200 195.800 ;
        RECT 212.900 195.900 213.200 196.500 ;
        RECT 213.500 196.500 213.900 196.600 ;
        RECT 215.800 196.500 216.200 196.600 ;
        RECT 213.500 196.200 216.200 196.500 ;
        RECT 212.900 195.700 215.300 195.900 ;
        RECT 217.400 195.700 217.800 199.900 ;
        RECT 219.500 196.200 219.900 199.900 ;
        RECT 220.200 196.800 220.600 197.200 ;
        RECT 220.300 196.200 220.600 196.800 ;
        RECT 219.500 195.900 220.000 196.200 ;
        RECT 220.300 195.900 221.000 196.200 ;
        RECT 212.900 195.600 217.800 195.700 ;
        RECT 214.900 195.500 217.800 195.600 ;
        RECT 215.000 195.400 217.800 195.500 ;
        RECT 209.500 194.900 209.900 195.000 ;
        RECT 209.500 194.600 211.400 194.900 ;
        RECT 211.800 194.800 212.200 195.200 ;
        RECT 214.200 195.100 214.600 195.200 ;
        RECT 214.200 194.800 216.700 195.100 ;
        RECT 211.000 194.500 211.400 194.600 ;
        RECT 211.900 194.200 212.200 194.800 ;
        RECT 216.300 194.700 216.700 194.800 ;
        RECT 219.000 194.400 219.400 195.200 ;
        RECT 215.500 194.200 215.900 194.300 ;
        RECT 219.700 194.200 220.000 195.900 ;
        RECT 220.600 195.800 221.000 195.900 ;
        RECT 221.400 195.600 221.800 199.900 ;
        RECT 223.500 197.900 224.100 199.900 ;
        RECT 225.800 197.900 226.200 199.900 ;
        RECT 228.000 198.200 228.400 199.900 ;
        RECT 228.000 197.900 229.000 198.200 ;
        RECT 223.800 197.500 224.200 197.900 ;
        RECT 225.900 197.600 226.200 197.900 ;
        RECT 225.500 197.300 227.300 197.600 ;
        RECT 228.600 197.500 229.000 197.900 ;
        RECT 225.500 197.200 225.900 197.300 ;
        RECT 226.900 197.200 227.300 197.300 ;
        RECT 223.400 196.600 224.100 197.000 ;
        RECT 223.800 196.100 224.100 196.600 ;
        RECT 224.900 196.500 226.000 196.800 ;
        RECT 224.900 196.400 225.300 196.500 ;
        RECT 223.800 195.800 225.000 196.100 ;
        RECT 221.400 195.300 223.500 195.600 ;
        RECT 211.900 193.900 217.400 194.200 ;
        RECT 212.100 193.800 212.500 193.900 ;
        RECT 203.000 193.000 205.000 193.100 ;
        RECT 203.000 191.100 203.400 193.000 ;
        RECT 204.600 191.100 205.000 193.000 ;
        RECT 205.400 191.100 205.800 193.100 ;
        RECT 206.500 192.800 207.400 193.100 ;
        RECT 208.600 193.300 210.500 193.600 ;
        RECT 206.500 191.100 206.900 192.800 ;
        RECT 208.600 191.100 209.000 193.300 ;
        RECT 210.100 193.200 210.500 193.300 ;
        RECT 215.000 192.800 215.300 193.900 ;
        RECT 216.600 193.800 217.400 193.900 ;
        RECT 218.200 194.100 218.600 194.200 ;
        RECT 218.200 193.800 219.000 194.100 ;
        RECT 219.700 193.800 221.000 194.200 ;
        RECT 218.600 193.600 219.000 193.800 ;
        RECT 214.100 192.700 214.500 192.800 ;
        RECT 211.000 192.100 211.400 192.500 ;
        RECT 213.100 192.400 214.500 192.700 ;
        RECT 215.000 192.400 215.400 192.800 ;
        RECT 213.100 192.100 213.400 192.400 ;
        RECT 215.800 192.100 216.200 192.500 ;
        RECT 210.700 191.800 211.400 192.100 ;
        RECT 210.700 191.100 211.300 191.800 ;
        RECT 213.000 191.100 213.400 192.100 ;
        RECT 215.200 191.800 216.200 192.100 ;
        RECT 215.200 191.100 215.600 191.800 ;
        RECT 217.400 191.100 217.800 193.500 ;
        RECT 218.300 193.100 220.100 193.300 ;
        RECT 220.600 193.100 220.900 193.800 ;
        RECT 221.400 193.600 221.800 195.300 ;
        RECT 223.100 195.200 223.500 195.300 ;
        RECT 224.700 195.200 225.000 195.800 ;
        RECT 225.700 195.900 226.000 196.500 ;
        RECT 226.300 196.500 226.700 196.600 ;
        RECT 228.600 196.500 229.000 196.600 ;
        RECT 226.300 196.200 229.000 196.500 ;
        RECT 225.700 195.700 228.100 195.900 ;
        RECT 230.200 195.700 230.600 199.900 ;
        RECT 225.700 195.600 230.600 195.700 ;
        RECT 227.700 195.500 230.600 195.600 ;
        RECT 227.800 195.400 230.600 195.500 ;
        RECT 222.300 194.900 222.700 195.000 ;
        RECT 222.300 194.600 224.200 194.900 ;
        RECT 224.600 194.800 225.000 195.200 ;
        RECT 225.400 195.100 225.800 195.200 ;
        RECT 227.000 195.100 227.400 195.200 ;
        RECT 225.400 194.800 229.500 195.100 ;
        RECT 223.800 194.500 224.200 194.600 ;
        RECT 224.700 194.200 225.000 194.800 ;
        RECT 229.100 194.700 229.500 194.800 ;
        RECT 228.300 194.200 228.700 194.300 ;
        RECT 224.700 193.900 230.200 194.200 ;
        RECT 224.900 193.800 225.300 193.900 ;
        RECT 221.400 193.300 223.300 193.600 ;
        RECT 218.200 193.000 220.200 193.100 ;
        RECT 218.200 191.100 218.600 193.000 ;
        RECT 219.800 191.100 220.200 193.000 ;
        RECT 220.600 191.100 221.000 193.100 ;
        RECT 221.400 191.100 221.800 193.300 ;
        RECT 222.900 193.200 223.300 193.300 ;
        RECT 227.800 192.800 228.100 193.900 ;
        RECT 229.400 193.800 230.200 193.900 ;
        RECT 226.900 192.700 227.300 192.800 ;
        RECT 223.800 192.100 224.200 192.500 ;
        RECT 225.900 192.400 227.300 192.700 ;
        RECT 227.800 192.400 228.200 192.800 ;
        RECT 225.900 192.100 226.200 192.400 ;
        RECT 228.600 192.100 229.000 192.500 ;
        RECT 223.500 191.800 224.200 192.100 ;
        RECT 223.500 191.100 224.100 191.800 ;
        RECT 225.800 191.100 226.200 192.100 ;
        RECT 228.000 191.800 229.000 192.100 ;
        RECT 228.000 191.100 228.400 191.800 ;
        RECT 230.200 191.100 230.600 193.500 ;
        RECT 0.600 187.500 1.000 189.900 ;
        RECT 2.800 189.200 3.200 189.900 ;
        RECT 2.200 188.900 3.200 189.200 ;
        RECT 5.000 188.900 5.400 189.900 ;
        RECT 7.100 189.200 7.700 189.900 ;
        RECT 7.000 188.900 7.700 189.200 ;
        RECT 2.200 188.500 2.600 188.900 ;
        RECT 5.000 188.600 5.300 188.900 ;
        RECT 3.000 188.200 3.400 188.600 ;
        RECT 3.900 188.300 5.300 188.600 ;
        RECT 7.000 188.500 7.400 188.900 ;
        RECT 3.900 188.200 4.300 188.300 ;
        RECT 1.000 187.100 1.800 187.200 ;
        RECT 3.100 187.100 3.400 188.200 ;
        RECT 7.900 187.700 8.300 187.800 ;
        RECT 9.400 187.700 9.800 189.900 ;
        RECT 10.200 187.900 10.600 189.900 ;
        RECT 11.000 188.000 11.400 189.900 ;
        RECT 12.600 188.000 13.000 189.900 ;
        RECT 11.000 187.900 13.000 188.000 ;
        RECT 13.400 187.900 13.800 189.900 ;
        RECT 14.200 188.000 14.600 189.900 ;
        RECT 15.800 188.000 16.200 189.900 ;
        RECT 14.200 187.900 16.200 188.000 ;
        RECT 7.900 187.400 9.800 187.700 ;
        RECT 5.900 187.100 6.300 187.200 ;
        RECT 1.000 186.800 6.500 187.100 ;
        RECT 2.500 186.700 2.900 186.800 ;
        RECT 1.700 186.200 2.100 186.300 ;
        RECT 6.200 186.200 6.500 186.800 ;
        RECT 7.000 186.400 7.400 186.500 ;
        RECT 1.700 186.100 4.200 186.200 ;
        RECT 4.600 186.100 5.000 186.200 ;
        RECT 1.700 185.900 5.000 186.100 ;
        RECT 3.800 185.800 5.000 185.900 ;
        RECT 6.200 185.800 6.600 186.200 ;
        RECT 7.000 186.100 8.900 186.400 ;
        RECT 8.500 186.000 8.900 186.100 ;
        RECT 0.600 185.500 3.400 185.600 ;
        RECT 0.600 185.400 3.500 185.500 ;
        RECT 0.600 185.300 5.500 185.400 ;
        RECT 0.600 181.100 1.000 185.300 ;
        RECT 3.100 185.100 5.500 185.300 ;
        RECT 2.200 184.500 4.900 184.800 ;
        RECT 2.200 184.400 2.600 184.500 ;
        RECT 4.500 184.400 4.900 184.500 ;
        RECT 5.200 184.500 5.500 185.100 ;
        RECT 6.200 185.200 6.500 185.800 ;
        RECT 7.700 185.700 8.100 185.800 ;
        RECT 9.400 185.700 9.800 187.400 ;
        RECT 10.300 187.200 10.600 187.900 ;
        RECT 11.100 187.700 12.900 187.900 ;
        RECT 12.200 187.200 12.600 187.400 ;
        RECT 13.500 187.200 13.800 187.900 ;
        RECT 14.300 187.700 16.100 187.900 ;
        RECT 16.600 187.500 17.000 189.900 ;
        RECT 18.800 189.200 19.200 189.900 ;
        RECT 18.200 188.900 19.200 189.200 ;
        RECT 21.000 188.900 21.400 189.900 ;
        RECT 23.100 189.200 23.700 189.900 ;
        RECT 23.000 188.900 23.700 189.200 ;
        RECT 18.200 188.500 18.600 188.900 ;
        RECT 21.000 188.600 21.300 188.900 ;
        RECT 19.000 188.200 19.400 188.600 ;
        RECT 19.900 188.300 21.300 188.600 ;
        RECT 23.000 188.500 23.400 188.900 ;
        RECT 19.900 188.200 20.300 188.300 ;
        RECT 15.400 187.200 15.800 187.400 ;
        RECT 10.200 186.800 11.500 187.200 ;
        RECT 12.200 186.900 13.000 187.200 ;
        RECT 12.600 186.800 13.000 186.900 ;
        RECT 13.400 186.800 14.700 187.200 ;
        RECT 15.400 186.900 16.200 187.200 ;
        RECT 15.800 186.800 16.200 186.900 ;
        RECT 17.000 187.100 17.800 187.200 ;
        RECT 19.100 187.100 19.400 188.200 ;
        RECT 23.900 187.700 24.300 187.800 ;
        RECT 25.400 187.700 25.800 189.900 ;
        RECT 26.200 188.000 26.600 189.900 ;
        RECT 27.800 188.000 28.200 189.900 ;
        RECT 26.200 187.900 28.200 188.000 ;
        RECT 28.600 187.900 29.000 189.900 ;
        RECT 29.400 187.900 29.800 189.900 ;
        RECT 30.200 188.000 30.600 189.900 ;
        RECT 31.800 188.000 32.200 189.900 ;
        RECT 30.200 187.900 32.200 188.000 ;
        RECT 32.600 188.000 33.000 189.900 ;
        RECT 34.200 188.000 34.600 189.900 ;
        RECT 32.600 187.900 34.600 188.000 ;
        RECT 35.000 187.900 35.400 189.900 ;
        RECT 39.300 188.000 39.700 189.500 ;
        RECT 41.400 188.500 41.800 189.500 ;
        RECT 26.300 187.700 28.100 187.900 ;
        RECT 23.900 187.400 25.800 187.700 ;
        RECT 21.900 187.100 22.300 187.200 ;
        RECT 17.000 186.800 22.500 187.100 ;
        RECT 7.700 185.400 9.800 185.700 ;
        RECT 6.200 184.900 7.400 185.200 ;
        RECT 5.900 184.500 6.300 184.600 ;
        RECT 5.200 184.200 6.300 184.500 ;
        RECT 7.100 184.400 7.400 184.900 ;
        RECT 7.100 184.000 7.800 184.400 ;
        RECT 3.900 183.700 4.300 183.800 ;
        RECT 5.300 183.700 5.700 183.800 ;
        RECT 2.200 183.100 2.600 183.500 ;
        RECT 3.900 183.400 5.700 183.700 ;
        RECT 5.000 183.100 5.300 183.400 ;
        RECT 7.000 183.100 7.400 183.500 ;
        RECT 2.200 182.800 3.200 183.100 ;
        RECT 2.800 181.100 3.200 182.800 ;
        RECT 5.000 181.100 5.400 183.100 ;
        RECT 7.100 181.100 7.700 183.100 ;
        RECT 9.400 181.100 9.800 185.400 ;
        RECT 10.200 185.100 10.600 185.200 ;
        RECT 11.200 185.100 11.500 186.800 ;
        RECT 11.800 185.800 12.200 186.600 ;
        RECT 12.600 186.100 13.000 186.200 ;
        RECT 14.400 186.100 14.700 186.800 ;
        RECT 18.500 186.700 18.900 186.800 ;
        RECT 12.600 185.800 14.700 186.100 ;
        RECT 15.000 185.800 15.400 186.600 ;
        RECT 17.700 186.200 18.100 186.300 ;
        RECT 22.200 186.200 22.500 186.800 ;
        RECT 23.000 186.400 23.400 186.500 ;
        RECT 17.700 185.900 20.200 186.200 ;
        RECT 19.800 185.800 20.200 185.900 ;
        RECT 22.200 185.800 22.600 186.200 ;
        RECT 23.000 186.100 24.900 186.400 ;
        RECT 24.500 186.000 24.900 186.100 ;
        RECT 13.400 185.100 13.800 185.200 ;
        RECT 14.400 185.100 14.700 185.800 ;
        RECT 16.600 185.500 19.400 185.600 ;
        RECT 16.600 185.400 19.500 185.500 ;
        RECT 16.600 185.300 21.500 185.400 ;
        RECT 10.200 184.800 10.900 185.100 ;
        RECT 11.200 184.800 11.700 185.100 ;
        RECT 13.400 184.800 14.100 185.100 ;
        RECT 14.400 184.800 14.900 185.100 ;
        RECT 10.600 184.200 10.900 184.800 ;
        RECT 10.600 183.800 11.000 184.200 ;
        RECT 11.300 181.100 11.700 184.800 ;
        RECT 13.800 184.200 14.100 184.800 ;
        RECT 13.400 183.800 14.200 184.200 ;
        RECT 14.500 181.100 14.900 184.800 ;
        RECT 16.600 181.100 17.000 185.300 ;
        RECT 19.100 185.100 21.500 185.300 ;
        RECT 18.200 184.500 20.900 184.800 ;
        RECT 18.200 184.400 18.600 184.500 ;
        RECT 20.500 184.400 20.900 184.500 ;
        RECT 21.200 184.500 21.500 185.100 ;
        RECT 22.200 185.200 22.500 185.800 ;
        RECT 23.700 185.700 24.100 185.800 ;
        RECT 25.400 185.700 25.800 187.400 ;
        RECT 26.600 187.200 27.000 187.400 ;
        RECT 28.600 187.200 28.900 187.900 ;
        RECT 29.500 187.200 29.800 187.900 ;
        RECT 30.300 187.700 32.100 187.900 ;
        RECT 32.700 187.700 34.500 187.900 ;
        RECT 31.400 187.200 31.800 187.400 ;
        RECT 33.000 187.200 33.400 187.400 ;
        RECT 35.000 187.200 35.300 187.900 ;
        RECT 38.900 187.700 39.700 188.000 ;
        RECT 38.900 187.500 39.300 187.700 ;
        RECT 38.900 187.200 39.200 187.500 ;
        RECT 41.500 187.400 41.800 188.500 ;
        RECT 42.200 187.500 42.600 189.900 ;
        RECT 44.400 189.200 44.800 189.900 ;
        RECT 43.800 188.900 44.800 189.200 ;
        RECT 46.600 188.900 47.000 189.900 ;
        RECT 48.700 189.200 49.300 189.900 ;
        RECT 48.600 188.900 49.300 189.200 ;
        RECT 43.800 188.500 44.200 188.900 ;
        RECT 46.600 188.600 46.900 188.900 ;
        RECT 44.600 188.200 45.000 188.600 ;
        RECT 45.500 188.300 46.900 188.600 ;
        RECT 48.600 188.500 49.000 188.900 ;
        RECT 45.500 188.200 45.900 188.300 ;
        RECT 26.200 186.900 27.000 187.200 ;
        RECT 26.200 186.800 26.600 186.900 ;
        RECT 27.700 186.800 29.000 187.200 ;
        RECT 29.400 186.800 30.700 187.200 ;
        RECT 31.400 187.100 32.200 187.200 ;
        RECT 32.600 187.100 33.400 187.200 ;
        RECT 31.400 186.900 33.400 187.100 ;
        RECT 31.800 186.800 33.000 186.900 ;
        RECT 34.100 186.800 35.400 187.200 ;
        RECT 38.200 186.800 39.200 187.200 ;
        RECT 39.700 187.100 41.800 187.400 ;
        RECT 42.600 187.100 43.400 187.200 ;
        RECT 44.700 187.100 45.000 188.200 ;
        RECT 49.500 187.700 49.900 187.800 ;
        RECT 51.000 187.700 51.400 189.900 ;
        RECT 51.800 188.000 52.200 189.900 ;
        RECT 53.400 188.000 53.800 189.900 ;
        RECT 51.800 187.900 53.800 188.000 ;
        RECT 54.200 187.900 54.600 189.900 ;
        RECT 55.000 187.900 55.400 189.900 ;
        RECT 55.800 188.000 56.200 189.900 ;
        RECT 57.400 188.000 57.800 189.900 ;
        RECT 55.800 187.900 57.800 188.000 ;
        RECT 58.200 187.900 58.600 189.900 ;
        RECT 59.000 188.000 59.400 189.900 ;
        RECT 60.600 188.000 61.000 189.900 ;
        RECT 59.000 187.900 61.000 188.000 ;
        RECT 61.400 188.500 61.800 189.500 ;
        RECT 51.900 187.700 53.700 187.900 ;
        RECT 49.500 187.400 51.400 187.700 ;
        RECT 46.200 187.100 46.600 187.200 ;
        RECT 47.500 187.100 47.900 187.200 ;
        RECT 39.700 186.900 40.200 187.100 ;
        RECT 27.000 185.800 27.400 186.600 ;
        RECT 23.700 185.400 25.800 185.700 ;
        RECT 22.200 184.900 23.400 185.200 ;
        RECT 21.900 184.500 22.300 184.600 ;
        RECT 21.200 184.200 22.300 184.500 ;
        RECT 23.100 184.400 23.400 184.900 ;
        RECT 23.100 184.000 23.800 184.400 ;
        RECT 19.900 183.700 20.300 183.800 ;
        RECT 21.300 183.700 21.700 183.800 ;
        RECT 18.200 183.100 18.600 183.500 ;
        RECT 19.900 183.400 21.700 183.700 ;
        RECT 21.000 183.100 21.300 183.400 ;
        RECT 23.000 183.100 23.400 183.500 ;
        RECT 18.200 182.800 19.200 183.100 ;
        RECT 18.800 181.100 19.200 182.800 ;
        RECT 21.000 181.100 21.400 183.100 ;
        RECT 23.100 181.100 23.700 183.100 ;
        RECT 25.400 181.100 25.800 185.400 ;
        RECT 27.700 185.100 28.000 186.800 ;
        RECT 30.400 186.100 30.700 186.800 ;
        RECT 28.600 185.800 30.700 186.100 ;
        RECT 31.000 186.100 31.400 186.600 ;
        RECT 33.400 186.100 33.800 186.600 ;
        RECT 31.000 185.800 33.800 186.100 ;
        RECT 28.600 185.200 28.900 185.800 ;
        RECT 28.600 185.100 29.000 185.200 ;
        RECT 27.500 184.800 28.000 185.100 ;
        RECT 28.300 184.800 29.000 185.100 ;
        RECT 29.400 185.100 29.800 185.200 ;
        RECT 30.400 185.100 30.700 185.800 ;
        RECT 34.100 185.100 34.400 186.800 ;
        RECT 38.200 185.400 38.600 186.200 ;
        RECT 35.000 185.100 35.400 185.200 ;
        RECT 29.400 184.800 30.100 185.100 ;
        RECT 30.400 184.800 30.900 185.100 ;
        RECT 27.500 181.100 27.900 184.800 ;
        RECT 28.300 184.200 28.600 184.800 ;
        RECT 29.800 184.200 30.100 184.800 ;
        RECT 28.200 183.800 28.600 184.200 ;
        RECT 29.400 183.800 30.200 184.200 ;
        RECT 30.500 181.100 30.900 184.800 ;
        RECT 33.900 184.800 34.400 185.100 ;
        RECT 34.700 184.800 35.400 185.100 ;
        RECT 38.900 184.900 39.200 186.800 ;
        RECT 39.500 186.500 40.200 186.900 ;
        RECT 42.600 186.800 48.100 187.100 ;
        RECT 44.100 186.700 44.500 186.800 ;
        RECT 39.900 185.500 40.200 186.500 ;
        RECT 40.600 185.800 41.000 186.600 ;
        RECT 41.400 185.800 41.800 186.600 ;
        RECT 43.300 186.200 43.700 186.300 ;
        RECT 43.300 186.100 45.800 186.200 ;
        RECT 47.000 186.100 47.400 186.200 ;
        RECT 43.300 185.900 47.400 186.100 ;
        RECT 45.400 185.800 47.400 185.900 ;
        RECT 42.200 185.500 45.000 185.600 ;
        RECT 39.900 185.200 41.800 185.500 ;
        RECT 33.900 182.200 34.300 184.800 ;
        RECT 34.700 184.200 35.000 184.800 ;
        RECT 38.900 184.600 39.700 184.900 ;
        RECT 34.600 183.800 35.400 184.200 ;
        RECT 33.400 181.800 34.300 182.200 ;
        RECT 33.900 181.100 34.300 181.800 ;
        RECT 39.300 182.200 39.700 184.600 ;
        RECT 41.500 183.500 41.800 185.200 ;
        RECT 39.300 181.800 40.200 182.200 ;
        RECT 39.300 181.100 39.700 181.800 ;
        RECT 41.400 181.500 41.800 183.500 ;
        RECT 42.200 185.400 45.100 185.500 ;
        RECT 42.200 185.300 47.100 185.400 ;
        RECT 42.200 181.100 42.600 185.300 ;
        RECT 44.700 185.100 47.100 185.300 ;
        RECT 43.800 184.500 46.500 184.800 ;
        RECT 43.800 184.400 44.200 184.500 ;
        RECT 46.100 184.400 46.500 184.500 ;
        RECT 46.800 184.500 47.100 185.100 ;
        RECT 47.800 185.200 48.100 186.800 ;
        RECT 48.600 186.400 49.000 186.500 ;
        RECT 48.600 186.100 50.500 186.400 ;
        RECT 50.100 186.000 50.500 186.100 ;
        RECT 49.300 185.700 49.700 185.800 ;
        RECT 51.000 185.700 51.400 187.400 ;
        RECT 52.200 187.200 52.600 187.400 ;
        RECT 54.200 187.200 54.500 187.900 ;
        RECT 55.100 187.200 55.400 187.900 ;
        RECT 55.900 187.700 57.700 187.900 ;
        RECT 57.000 187.200 57.400 187.400 ;
        RECT 58.300 187.200 58.600 187.900 ;
        RECT 59.100 187.700 60.900 187.900 ;
        RECT 61.400 187.400 61.700 188.500 ;
        RECT 63.500 188.000 63.900 189.500 ;
        RECT 63.500 187.700 64.300 188.000 ;
        RECT 66.200 187.900 66.600 189.900 ;
        RECT 67.000 188.000 67.400 189.900 ;
        RECT 68.600 188.000 69.000 189.900 ;
        RECT 67.000 187.900 69.000 188.000 ;
        RECT 63.900 187.500 64.300 187.700 ;
        RECT 60.200 187.200 60.600 187.400 ;
        RECT 51.800 186.900 52.600 187.200 ;
        RECT 51.800 186.800 52.200 186.900 ;
        RECT 53.300 186.800 54.600 187.200 ;
        RECT 55.000 186.800 56.300 187.200 ;
        RECT 57.000 186.900 57.800 187.200 ;
        RECT 57.400 186.800 57.800 186.900 ;
        RECT 58.200 186.800 59.500 187.200 ;
        RECT 60.200 186.900 61.000 187.200 ;
        RECT 61.400 187.100 63.500 187.400 ;
        RECT 60.600 186.800 61.000 186.900 ;
        RECT 63.000 186.900 63.500 187.100 ;
        RECT 64.000 187.200 64.300 187.500 ;
        RECT 66.300 187.200 66.600 187.900 ;
        RECT 67.100 187.700 68.900 187.900 ;
        RECT 69.400 187.600 69.800 189.900 ;
        RECT 71.000 188.200 71.400 189.900 ;
        RECT 71.000 187.900 71.500 188.200 ;
        RECT 74.500 188.000 74.900 189.500 ;
        RECT 76.600 188.500 77.000 189.500 ;
        RECT 68.200 187.200 68.600 187.400 ;
        RECT 69.400 187.300 70.700 187.600 ;
        RECT 52.600 185.800 53.000 186.600 ;
        RECT 53.300 186.200 53.600 186.800 ;
        RECT 53.300 185.800 53.800 186.200 ;
        RECT 56.000 186.100 56.300 186.800 ;
        RECT 54.200 185.800 56.300 186.100 ;
        RECT 56.600 185.800 57.000 186.600 ;
        RECT 49.300 185.400 51.400 185.700 ;
        RECT 47.800 184.900 49.000 185.200 ;
        RECT 47.500 184.500 47.900 184.600 ;
        RECT 46.800 184.200 47.900 184.500 ;
        RECT 48.700 184.400 49.000 184.900 ;
        RECT 48.700 184.000 49.400 184.400 ;
        RECT 45.500 183.700 45.900 183.800 ;
        RECT 46.900 183.700 47.300 183.800 ;
        RECT 43.800 183.100 44.200 183.500 ;
        RECT 45.500 183.400 47.300 183.700 ;
        RECT 46.600 183.100 46.900 183.400 ;
        RECT 48.600 183.100 49.000 183.500 ;
        RECT 43.800 182.800 44.800 183.100 ;
        RECT 44.400 181.100 44.800 182.800 ;
        RECT 46.600 181.100 47.000 183.100 ;
        RECT 48.700 181.100 49.300 183.100 ;
        RECT 51.000 181.100 51.400 185.400 ;
        RECT 53.300 185.100 53.600 185.800 ;
        RECT 54.200 185.200 54.500 185.800 ;
        RECT 54.200 185.100 54.600 185.200 ;
        RECT 53.100 184.800 53.600 185.100 ;
        RECT 53.900 184.800 54.600 185.100 ;
        RECT 55.000 185.100 55.400 185.200 ;
        RECT 56.000 185.100 56.300 185.800 ;
        RECT 58.200 185.100 58.600 185.200 ;
        RECT 59.200 185.100 59.500 186.800 ;
        RECT 59.800 185.800 60.200 186.600 ;
        RECT 61.400 185.800 61.800 186.600 ;
        RECT 62.200 185.800 62.600 186.600 ;
        RECT 63.000 186.500 63.700 186.900 ;
        RECT 64.000 186.800 65.000 187.200 ;
        RECT 66.200 186.800 67.500 187.200 ;
        RECT 68.200 186.900 69.000 187.200 ;
        RECT 68.600 186.800 69.000 186.900 ;
        RECT 63.000 185.500 63.300 186.500 ;
        RECT 61.400 185.200 63.300 185.500 ;
        RECT 55.000 184.800 55.700 185.100 ;
        RECT 56.000 184.800 56.500 185.100 ;
        RECT 58.200 184.800 58.900 185.100 ;
        RECT 59.200 184.800 59.700 185.100 ;
        RECT 53.100 181.100 53.500 184.800 ;
        RECT 53.900 184.200 54.200 184.800 ;
        RECT 53.800 183.800 54.200 184.200 ;
        RECT 55.400 184.200 55.700 184.800 ;
        RECT 55.400 183.800 55.800 184.200 ;
        RECT 56.100 181.100 56.500 184.800 ;
        RECT 58.600 184.200 58.900 184.800 ;
        RECT 58.600 183.800 59.000 184.200 ;
        RECT 59.300 181.100 59.700 184.800 ;
        RECT 61.400 183.500 61.700 185.200 ;
        RECT 64.000 184.900 64.300 186.800 ;
        RECT 64.600 185.400 65.000 186.200 ;
        RECT 63.500 184.600 64.300 184.900 ;
        RECT 66.200 185.100 66.600 185.200 ;
        RECT 67.200 185.100 67.500 186.800 ;
        RECT 67.800 185.800 68.200 186.600 ;
        RECT 69.500 186.200 69.900 186.600 ;
        RECT 68.600 186.100 69.000 186.200 ;
        RECT 69.400 186.100 69.900 186.200 ;
        RECT 68.600 185.800 69.900 186.100 ;
        RECT 70.400 186.500 70.700 187.300 ;
        RECT 71.200 187.200 71.500 187.900 ;
        RECT 74.100 187.700 74.900 188.000 ;
        RECT 74.100 187.500 74.500 187.700 ;
        RECT 74.100 187.200 74.400 187.500 ;
        RECT 76.700 187.400 77.000 188.500 ;
        RECT 71.000 187.100 71.500 187.200 ;
        RECT 71.800 187.100 72.200 187.200 ;
        RECT 71.000 186.800 72.200 187.100 ;
        RECT 72.600 187.100 73.000 187.200 ;
        RECT 73.400 187.100 74.400 187.200 ;
        RECT 72.600 186.800 74.400 187.100 ;
        RECT 74.900 187.100 77.000 187.400 ;
        RECT 77.400 187.700 77.800 189.900 ;
        RECT 79.500 189.200 80.100 189.900 ;
        RECT 79.500 188.900 80.200 189.200 ;
        RECT 81.800 188.900 82.200 189.900 ;
        RECT 84.000 189.200 84.400 189.900 ;
        RECT 84.000 188.900 85.000 189.200 ;
        RECT 79.800 188.500 80.200 188.900 ;
        RECT 81.900 188.600 82.200 188.900 ;
        RECT 81.900 188.300 83.300 188.600 ;
        RECT 82.900 188.200 83.300 188.300 ;
        RECT 83.800 187.800 84.200 188.600 ;
        RECT 84.600 188.500 85.000 188.900 ;
        RECT 78.900 187.700 79.300 187.800 ;
        RECT 77.400 187.400 79.300 187.700 ;
        RECT 74.900 186.900 75.400 187.100 ;
        RECT 70.400 186.100 70.900 186.500 ;
        RECT 70.400 185.100 70.700 186.100 ;
        RECT 71.200 185.100 71.500 186.800 ;
        RECT 73.400 185.400 73.800 186.200 ;
        RECT 66.200 184.800 66.900 185.100 ;
        RECT 67.200 184.800 67.700 185.100 ;
        RECT 61.400 181.500 61.800 183.500 ;
        RECT 63.500 182.200 63.900 184.600 ;
        RECT 66.600 184.200 66.900 184.800 ;
        RECT 66.600 183.800 67.000 184.200 ;
        RECT 63.500 181.800 64.200 182.200 ;
        RECT 63.500 181.100 63.900 181.800 ;
        RECT 67.300 181.100 67.700 184.800 ;
        RECT 69.400 184.800 70.700 185.100 ;
        RECT 69.400 181.100 69.800 184.800 ;
        RECT 71.000 184.600 71.500 185.100 ;
        RECT 74.100 184.900 74.400 186.800 ;
        RECT 74.700 186.500 75.400 186.900 ;
        RECT 75.100 185.500 75.400 186.500 ;
        RECT 75.800 185.800 76.200 186.600 ;
        RECT 76.600 185.800 77.000 186.600 ;
        RECT 77.400 185.700 77.800 187.400 ;
        RECT 80.900 187.100 81.300 187.200 ;
        RECT 83.800 187.100 84.100 187.800 ;
        RECT 86.200 187.500 86.600 189.900 ;
        RECT 87.000 187.900 87.400 189.900 ;
        RECT 87.800 188.000 88.200 189.900 ;
        RECT 89.400 188.000 89.800 189.900 ;
        RECT 87.800 187.900 89.800 188.000 ;
        RECT 91.800 187.900 92.200 189.900 ;
        RECT 92.600 188.000 93.000 189.900 ;
        RECT 94.200 188.000 94.600 189.900 ;
        RECT 92.600 187.900 94.600 188.000 ;
        RECT 95.000 188.500 95.400 189.500 ;
        RECT 87.100 187.200 87.400 187.900 ;
        RECT 87.900 187.700 89.700 187.900 ;
        RECT 89.000 187.200 89.400 187.400 ;
        RECT 91.900 187.200 92.200 187.900 ;
        RECT 92.700 187.700 94.500 187.900 ;
        RECT 95.000 187.400 95.300 188.500 ;
        RECT 97.100 188.000 97.500 189.500 ;
        RECT 99.800 188.500 100.200 189.500 ;
        RECT 97.100 187.700 97.900 188.000 ;
        RECT 97.500 187.500 97.900 187.700 ;
        RECT 93.800 187.200 94.200 187.400 ;
        RECT 85.400 187.100 86.200 187.200 ;
        RECT 80.700 186.800 86.200 187.100 ;
        RECT 87.000 186.800 88.300 187.200 ;
        RECT 89.000 187.100 89.800 187.200 ;
        RECT 90.200 187.100 90.600 187.200 ;
        RECT 89.000 186.900 90.600 187.100 ;
        RECT 89.400 186.800 90.600 186.900 ;
        RECT 91.800 186.800 93.100 187.200 ;
        RECT 93.800 186.900 94.600 187.200 ;
        RECT 95.000 187.100 97.100 187.400 ;
        RECT 94.200 186.800 94.600 186.900 ;
        RECT 96.600 186.900 97.100 187.100 ;
        RECT 97.600 187.200 97.900 187.500 ;
        RECT 99.800 187.400 100.100 188.500 ;
        RECT 101.900 188.000 102.300 189.500 ;
        RECT 106.500 188.000 106.900 189.500 ;
        RECT 108.600 188.500 109.000 189.500 ;
        RECT 101.900 187.700 102.700 188.000 ;
        RECT 102.300 187.500 102.700 187.700 ;
        RECT 97.600 187.100 98.600 187.200 ;
        RECT 99.000 187.100 99.400 187.200 ;
        RECT 99.800 187.100 101.900 187.400 ;
        RECT 79.800 186.400 80.200 186.500 ;
        RECT 78.300 186.100 80.200 186.400 ;
        RECT 78.300 186.000 78.700 186.100 ;
        RECT 79.100 185.700 79.500 185.800 ;
        RECT 75.100 185.200 77.000 185.500 ;
        RECT 74.100 184.600 74.900 184.900 ;
        RECT 71.000 181.100 71.400 184.600 ;
        RECT 74.500 181.100 74.900 184.600 ;
        RECT 76.700 183.500 77.000 185.200 ;
        RECT 76.600 181.500 77.000 183.500 ;
        RECT 77.400 185.400 79.500 185.700 ;
        RECT 77.400 181.100 77.800 185.400 ;
        RECT 80.700 185.200 81.000 186.800 ;
        RECT 84.300 186.700 84.700 186.800 ;
        RECT 83.800 186.200 84.200 186.300 ;
        RECT 85.100 186.200 85.500 186.300 ;
        RECT 83.000 185.900 85.500 186.200 ;
        RECT 83.000 185.800 83.400 185.900 ;
        RECT 83.800 185.500 86.600 185.600 ;
        RECT 83.700 185.400 86.600 185.500 ;
        RECT 79.800 184.900 81.000 185.200 ;
        RECT 81.700 185.300 86.600 185.400 ;
        RECT 81.700 185.100 84.100 185.300 ;
        RECT 79.800 184.400 80.100 184.900 ;
        RECT 79.400 184.000 80.100 184.400 ;
        RECT 80.900 184.500 81.300 184.600 ;
        RECT 81.700 184.500 82.000 185.100 ;
        RECT 80.900 184.200 82.000 184.500 ;
        RECT 82.300 184.500 85.000 184.800 ;
        RECT 82.300 184.400 82.700 184.500 ;
        RECT 84.600 184.400 85.000 184.500 ;
        RECT 81.500 183.700 81.900 183.800 ;
        RECT 82.900 183.700 83.300 183.800 ;
        RECT 79.800 183.100 80.200 183.500 ;
        RECT 81.500 183.400 83.300 183.700 ;
        RECT 81.900 183.100 82.200 183.400 ;
        RECT 84.600 183.100 85.000 183.500 ;
        RECT 79.500 181.100 80.100 183.100 ;
        RECT 81.800 181.100 82.200 183.100 ;
        RECT 84.000 182.800 85.000 183.100 ;
        RECT 84.000 181.100 84.400 182.800 ;
        RECT 86.200 181.100 86.600 185.300 ;
        RECT 87.000 185.100 87.400 185.200 ;
        RECT 88.000 185.100 88.300 186.800 ;
        RECT 88.600 186.100 89.000 186.600 ;
        RECT 89.400 186.100 89.800 186.200 ;
        RECT 88.600 185.800 89.800 186.100 ;
        RECT 91.800 185.100 92.200 185.200 ;
        RECT 92.800 185.100 93.100 186.800 ;
        RECT 93.400 185.800 93.800 186.600 ;
        RECT 95.000 185.800 95.400 186.600 ;
        RECT 95.800 185.800 96.200 186.600 ;
        RECT 96.600 186.500 97.300 186.900 ;
        RECT 97.600 186.800 99.400 187.100 ;
        RECT 101.400 186.900 101.900 187.100 ;
        RECT 102.400 187.200 102.700 187.500 ;
        RECT 106.100 187.700 106.900 188.000 ;
        RECT 106.100 187.500 106.500 187.700 ;
        RECT 106.100 187.200 106.400 187.500 ;
        RECT 108.700 187.400 109.000 188.500 ;
        RECT 110.200 188.200 110.600 189.900 ;
        RECT 96.600 185.500 96.900 186.500 ;
        RECT 95.000 185.200 96.900 185.500 ;
        RECT 87.000 184.800 87.700 185.100 ;
        RECT 88.000 184.800 88.500 185.100 ;
        RECT 91.800 184.800 92.500 185.100 ;
        RECT 92.800 184.800 93.300 185.100 ;
        RECT 87.400 184.200 87.700 184.800 ;
        RECT 88.100 184.200 88.500 184.800 ;
        RECT 92.200 184.200 92.500 184.800 ;
        RECT 87.400 183.800 87.800 184.200 ;
        RECT 88.100 183.800 89.000 184.200 ;
        RECT 92.200 183.800 92.600 184.200 ;
        RECT 88.100 181.100 88.500 183.800 ;
        RECT 92.900 181.100 93.300 184.800 ;
        RECT 95.000 183.500 95.300 185.200 ;
        RECT 97.600 184.900 97.900 186.800 ;
        RECT 98.200 185.400 98.600 186.200 ;
        RECT 99.800 185.800 100.200 186.600 ;
        RECT 100.600 185.800 101.000 186.600 ;
        RECT 101.400 186.500 102.100 186.900 ;
        RECT 102.400 186.800 103.400 187.200 ;
        RECT 105.400 187.100 106.400 187.200 ;
        RECT 103.800 186.800 106.400 187.100 ;
        RECT 106.900 187.100 109.000 187.400 ;
        RECT 110.100 187.800 110.600 188.200 ;
        RECT 110.100 187.200 110.400 187.800 ;
        RECT 111.800 187.600 112.200 189.900 ;
        RECT 110.900 187.300 112.200 187.600 ;
        RECT 112.600 187.600 113.000 189.900 ;
        RECT 114.200 188.200 114.600 189.900 ;
        RECT 114.200 187.900 114.700 188.200 ;
        RECT 115.800 188.000 116.200 189.900 ;
        RECT 117.400 188.000 117.800 189.900 ;
        RECT 115.800 187.900 117.800 188.000 ;
        RECT 118.200 187.900 118.600 189.900 ;
        RECT 119.000 187.900 119.400 189.900 ;
        RECT 119.800 188.000 120.200 189.900 ;
        RECT 121.400 188.000 121.800 189.900 ;
        RECT 119.800 187.900 121.800 188.000 ;
        RECT 112.600 187.300 113.900 187.600 ;
        RECT 106.900 186.900 107.400 187.100 ;
        RECT 101.400 185.500 101.700 186.500 ;
        RECT 97.100 184.600 97.900 184.900 ;
        RECT 99.800 185.200 101.700 185.500 ;
        RECT 95.000 181.500 95.400 183.500 ;
        RECT 97.100 181.100 97.500 184.600 ;
        RECT 99.800 183.500 100.100 185.200 ;
        RECT 102.400 184.900 102.700 186.800 ;
        RECT 103.000 186.100 103.400 186.200 ;
        RECT 103.800 186.100 104.100 186.800 ;
        RECT 103.000 185.800 104.100 186.100 ;
        RECT 104.600 186.100 105.000 186.200 ;
        RECT 105.400 186.100 105.800 186.200 ;
        RECT 104.600 185.800 105.800 186.100 ;
        RECT 103.000 185.400 103.400 185.800 ;
        RECT 105.400 185.400 105.800 185.800 ;
        RECT 101.900 184.600 102.700 184.900 ;
        RECT 106.100 184.900 106.400 186.800 ;
        RECT 106.700 186.500 107.400 186.900 ;
        RECT 110.100 186.800 110.600 187.200 ;
        RECT 107.100 185.500 107.400 186.500 ;
        RECT 107.800 185.800 108.200 186.600 ;
        RECT 108.600 185.800 109.000 186.600 ;
        RECT 107.100 185.200 109.000 185.500 ;
        RECT 106.100 184.600 106.900 184.900 ;
        RECT 99.800 181.500 100.200 183.500 ;
        RECT 101.900 183.200 102.300 184.600 ;
        RECT 101.900 182.800 102.600 183.200 ;
        RECT 101.900 181.100 102.300 182.800 ;
        RECT 106.500 181.100 106.900 184.600 ;
        RECT 108.700 183.500 109.000 185.200 ;
        RECT 110.100 185.100 110.400 186.800 ;
        RECT 110.900 186.500 111.200 187.300 ;
        RECT 110.700 186.100 111.200 186.500 ;
        RECT 110.900 185.100 111.200 186.100 ;
        RECT 111.700 186.200 112.100 186.600 ;
        RECT 112.700 186.200 113.100 186.600 ;
        RECT 111.700 186.100 112.200 186.200 ;
        RECT 112.600 186.100 113.100 186.200 ;
        RECT 111.700 185.800 113.100 186.100 ;
        RECT 113.600 186.500 113.900 187.300 ;
        RECT 114.400 187.200 114.700 187.900 ;
        RECT 115.900 187.700 117.700 187.900 ;
        RECT 116.200 187.200 116.600 187.400 ;
        RECT 118.200 187.200 118.500 187.900 ;
        RECT 119.100 187.200 119.400 187.900 ;
        RECT 119.900 187.700 121.700 187.900 ;
        RECT 122.200 187.700 122.600 189.900 ;
        RECT 124.300 189.200 124.900 189.900 ;
        RECT 124.300 188.900 125.000 189.200 ;
        RECT 126.600 188.900 127.000 189.900 ;
        RECT 128.800 189.200 129.200 189.900 ;
        RECT 128.800 188.900 129.800 189.200 ;
        RECT 124.600 188.500 125.000 188.900 ;
        RECT 126.700 188.600 127.000 188.900 ;
        RECT 126.700 188.300 128.100 188.600 ;
        RECT 127.700 188.200 128.100 188.300 ;
        RECT 128.600 187.800 129.000 188.600 ;
        RECT 129.400 188.500 129.800 188.900 ;
        RECT 123.700 187.700 124.100 187.800 ;
        RECT 122.200 187.400 124.100 187.700 ;
        RECT 121.000 187.200 121.400 187.400 ;
        RECT 114.200 186.800 114.700 187.200 ;
        RECT 115.800 186.900 116.600 187.200 ;
        RECT 115.800 186.800 116.200 186.900 ;
        RECT 117.300 186.800 118.600 187.200 ;
        RECT 119.000 186.800 120.300 187.200 ;
        RECT 121.000 186.900 121.800 187.200 ;
        RECT 121.400 186.800 121.800 186.900 ;
        RECT 113.600 186.100 114.100 186.500 ;
        RECT 113.600 185.100 113.900 186.100 ;
        RECT 114.400 185.100 114.700 186.800 ;
        RECT 116.600 185.800 117.000 186.600 ;
        RECT 117.300 186.100 117.600 186.800 ;
        RECT 117.300 185.800 119.300 186.100 ;
        RECT 117.300 185.100 117.600 185.800 ;
        RECT 119.000 185.200 119.300 185.800 ;
        RECT 118.200 185.100 118.600 185.200 ;
        RECT 110.100 184.600 110.600 185.100 ;
        RECT 110.900 184.800 112.200 185.100 ;
        RECT 108.600 181.500 109.000 183.500 ;
        RECT 110.200 181.100 110.600 184.600 ;
        RECT 111.800 181.100 112.200 184.800 ;
        RECT 112.600 184.800 113.900 185.100 ;
        RECT 112.600 181.100 113.000 184.800 ;
        RECT 114.200 184.600 114.700 185.100 ;
        RECT 117.100 184.800 117.600 185.100 ;
        RECT 117.900 184.800 118.600 185.100 ;
        RECT 119.000 185.100 119.400 185.200 ;
        RECT 120.000 185.100 120.300 186.800 ;
        RECT 120.600 185.800 121.000 186.600 ;
        RECT 122.200 185.700 122.600 187.400 ;
        RECT 125.700 187.100 126.100 187.200 ;
        RECT 128.600 187.100 128.900 187.800 ;
        RECT 131.000 187.500 131.400 189.900 ;
        RECT 130.200 187.100 131.000 187.200 ;
        RECT 125.500 186.800 131.000 187.100 ;
        RECT 131.800 186.800 132.200 187.600 ;
        RECT 124.600 186.400 125.000 186.500 ;
        RECT 123.100 186.100 125.000 186.400 ;
        RECT 123.100 186.000 123.500 186.100 ;
        RECT 123.900 185.700 124.300 185.800 ;
        RECT 122.200 185.400 124.300 185.700 ;
        RECT 119.000 184.800 119.700 185.100 ;
        RECT 120.000 184.800 120.500 185.100 ;
        RECT 114.200 181.100 114.600 184.600 ;
        RECT 117.100 181.100 117.500 184.800 ;
        RECT 117.900 184.200 118.200 184.800 ;
        RECT 117.800 183.800 118.200 184.200 ;
        RECT 119.400 184.200 119.700 184.800 ;
        RECT 119.400 183.800 119.800 184.200 ;
        RECT 120.100 181.100 120.500 184.800 ;
        RECT 122.200 181.100 122.600 185.400 ;
        RECT 125.500 185.200 125.800 186.800 ;
        RECT 129.100 186.700 129.500 186.800 ;
        RECT 129.900 186.200 130.300 186.300 ;
        RECT 127.000 186.100 127.400 186.200 ;
        RECT 127.800 186.100 130.300 186.200 ;
        RECT 127.000 185.900 130.300 186.100 ;
        RECT 127.000 185.800 128.200 185.900 ;
        RECT 128.600 185.500 131.400 185.600 ;
        RECT 128.500 185.400 131.400 185.500 ;
        RECT 124.600 184.900 125.800 185.200 ;
        RECT 126.500 185.300 131.400 185.400 ;
        RECT 126.500 185.100 128.900 185.300 ;
        RECT 124.600 184.400 124.900 184.900 ;
        RECT 124.200 184.000 124.900 184.400 ;
        RECT 125.700 184.500 126.100 184.600 ;
        RECT 126.500 184.500 126.800 185.100 ;
        RECT 125.700 184.200 126.800 184.500 ;
        RECT 127.100 184.500 129.800 184.800 ;
        RECT 127.100 184.400 127.500 184.500 ;
        RECT 129.400 184.400 129.800 184.500 ;
        RECT 126.300 183.700 126.700 183.800 ;
        RECT 127.700 183.700 128.100 183.800 ;
        RECT 124.600 183.100 125.000 183.500 ;
        RECT 126.300 183.400 128.100 183.700 ;
        RECT 126.700 183.100 127.000 183.400 ;
        RECT 129.400 183.100 129.800 183.500 ;
        RECT 124.300 181.100 124.900 183.100 ;
        RECT 126.600 181.100 127.000 183.100 ;
        RECT 128.800 182.800 129.800 183.100 ;
        RECT 128.800 181.100 129.200 182.800 ;
        RECT 131.000 181.100 131.400 185.300 ;
        RECT 132.600 181.100 133.000 189.900 ;
        RECT 136.100 188.000 136.500 189.500 ;
        RECT 138.200 188.500 138.600 189.500 ;
        RECT 135.700 187.700 136.500 188.000 ;
        RECT 135.700 187.500 136.100 187.700 ;
        RECT 135.700 187.200 136.000 187.500 ;
        RECT 138.300 187.400 138.600 188.500 ;
        RECT 140.600 188.000 141.000 189.900 ;
        RECT 142.200 188.000 142.600 189.900 ;
        RECT 140.600 187.900 142.600 188.000 ;
        RECT 143.000 187.900 143.400 189.900 ;
        RECT 143.800 188.000 144.200 189.900 ;
        RECT 145.400 188.000 145.800 189.900 ;
        RECT 143.800 187.900 145.800 188.000 ;
        RECT 146.200 187.900 146.600 189.900 ;
        RECT 147.000 188.000 147.400 189.900 ;
        RECT 148.600 188.000 149.000 189.900 ;
        RECT 147.000 187.900 149.000 188.000 ;
        RECT 149.400 187.900 149.800 189.900 ;
        RECT 140.700 187.700 142.500 187.900 ;
        RECT 135.000 186.800 136.000 187.200 ;
        RECT 136.500 187.100 138.600 187.400 ;
        RECT 141.000 187.200 141.400 187.400 ;
        RECT 143.000 187.200 143.300 187.900 ;
        RECT 143.900 187.700 145.700 187.900 ;
        RECT 144.200 187.200 144.600 187.400 ;
        RECT 146.200 187.200 146.500 187.900 ;
        RECT 147.100 187.700 148.900 187.900 ;
        RECT 147.400 187.200 147.800 187.400 ;
        RECT 149.400 187.200 149.700 187.900 ;
        RECT 150.200 187.500 150.600 189.900 ;
        RECT 152.400 189.200 152.800 189.900 ;
        RECT 151.800 188.900 152.800 189.200 ;
        RECT 154.600 188.900 155.000 189.900 ;
        RECT 156.700 189.200 157.300 189.900 ;
        RECT 156.600 188.900 157.300 189.200 ;
        RECT 151.800 188.500 152.200 188.900 ;
        RECT 154.600 188.600 154.900 188.900 ;
        RECT 152.600 187.800 153.000 188.600 ;
        RECT 153.500 188.300 154.900 188.600 ;
        RECT 156.600 188.500 157.000 188.900 ;
        RECT 153.500 188.200 153.900 188.300 ;
        RECT 136.500 186.900 137.000 187.100 ;
        RECT 135.000 185.400 135.400 186.200 ;
        RECT 135.700 184.900 136.000 186.800 ;
        RECT 136.300 186.500 137.000 186.900 ;
        RECT 140.600 186.900 141.400 187.200 ;
        RECT 140.600 186.800 141.000 186.900 ;
        RECT 142.100 186.800 143.400 187.200 ;
        RECT 143.800 186.900 144.600 187.200 ;
        RECT 143.800 186.800 144.200 186.900 ;
        RECT 145.300 186.800 146.600 187.200 ;
        RECT 147.000 186.900 147.800 187.200 ;
        RECT 147.000 186.800 147.400 186.900 ;
        RECT 148.500 186.800 149.800 187.200 ;
        RECT 150.600 187.100 151.400 187.200 ;
        RECT 152.700 187.100 153.000 187.800 ;
        RECT 157.500 187.700 157.900 187.800 ;
        RECT 159.000 187.700 159.400 189.900 ;
        RECT 161.100 188.200 161.500 189.900 ;
        RECT 157.500 187.400 159.400 187.700 ;
        RECT 160.600 187.900 161.500 188.200 ;
        RECT 162.200 187.900 162.600 189.900 ;
        RECT 163.000 188.000 163.400 189.900 ;
        RECT 164.600 188.000 165.000 189.900 ;
        RECT 163.000 187.900 165.000 188.000 ;
        RECT 155.500 187.100 155.900 187.200 ;
        RECT 150.600 186.800 156.100 187.100 ;
        RECT 136.700 185.500 137.000 186.500 ;
        RECT 137.400 185.800 137.800 186.600 ;
        RECT 138.200 186.100 138.600 186.600 ;
        RECT 139.000 186.100 139.400 186.200 ;
        RECT 138.200 185.800 139.400 186.100 ;
        RECT 141.400 185.800 141.800 186.600 ;
        RECT 136.700 185.200 138.600 185.500 ;
        RECT 135.700 184.600 136.500 184.900 ;
        RECT 136.100 182.200 136.500 184.600 ;
        RECT 138.300 183.500 138.600 185.200 ;
        RECT 142.100 185.100 142.400 186.800 ;
        RECT 144.600 185.800 145.000 186.600 ;
        RECT 145.300 186.100 145.600 186.800 ;
        RECT 147.000 186.100 147.400 186.200 ;
        RECT 145.300 185.800 147.400 186.100 ;
        RECT 147.800 185.800 148.200 186.600 ;
        RECT 143.000 185.100 143.400 185.200 ;
        RECT 145.300 185.100 145.600 185.800 ;
        RECT 146.200 185.100 146.600 185.200 ;
        RECT 148.500 185.100 148.800 186.800 ;
        RECT 152.100 186.700 152.500 186.800 ;
        RECT 151.300 186.200 151.700 186.300 ;
        RECT 152.600 186.200 153.000 186.300 ;
        RECT 151.300 185.900 153.800 186.200 ;
        RECT 153.400 185.800 153.800 185.900 ;
        RECT 150.200 185.500 153.000 185.600 ;
        RECT 150.200 185.400 153.100 185.500 ;
        RECT 150.200 185.300 155.100 185.400 ;
        RECT 149.400 185.100 149.800 185.200 ;
        RECT 135.800 181.800 136.500 182.200 ;
        RECT 136.100 181.100 136.500 181.800 ;
        RECT 138.200 181.500 138.600 183.500 ;
        RECT 141.900 184.800 142.400 185.100 ;
        RECT 142.700 184.800 143.400 185.100 ;
        RECT 145.100 184.800 145.600 185.100 ;
        RECT 145.900 184.800 146.600 185.100 ;
        RECT 148.300 184.800 148.800 185.100 ;
        RECT 149.100 184.800 149.800 185.100 ;
        RECT 141.900 182.200 142.300 184.800 ;
        RECT 142.700 184.200 143.000 184.800 ;
        RECT 142.600 183.800 143.400 184.200 ;
        RECT 141.400 181.800 142.300 182.200 ;
        RECT 141.900 181.100 142.300 181.800 ;
        RECT 145.100 181.100 145.500 184.800 ;
        RECT 145.900 184.200 146.200 184.800 ;
        RECT 145.800 183.800 146.200 184.200 ;
        RECT 148.300 181.100 148.700 184.800 ;
        RECT 149.100 184.200 149.400 184.800 ;
        RECT 149.000 183.800 149.400 184.200 ;
        RECT 150.200 181.100 150.600 185.300 ;
        RECT 152.700 185.100 155.100 185.300 ;
        RECT 151.800 184.500 154.500 184.800 ;
        RECT 151.800 184.400 152.200 184.500 ;
        RECT 154.100 184.400 154.500 184.500 ;
        RECT 154.800 184.500 155.100 185.100 ;
        RECT 155.800 185.200 156.100 186.800 ;
        RECT 156.600 186.400 157.000 186.500 ;
        RECT 156.600 186.100 158.500 186.400 ;
        RECT 158.100 186.000 158.500 186.100 ;
        RECT 157.300 185.700 157.700 185.800 ;
        RECT 159.000 185.700 159.400 187.400 ;
        RECT 159.800 186.800 160.200 187.600 ;
        RECT 157.300 185.400 159.400 185.700 ;
        RECT 155.800 184.900 157.000 185.200 ;
        RECT 155.500 184.500 155.900 184.600 ;
        RECT 154.800 184.200 155.900 184.500 ;
        RECT 156.700 184.400 157.000 184.900 ;
        RECT 156.700 184.000 157.400 184.400 ;
        RECT 153.500 183.700 153.900 183.800 ;
        RECT 154.900 183.700 155.300 183.800 ;
        RECT 151.800 183.100 152.200 183.500 ;
        RECT 153.500 183.400 155.300 183.700 ;
        RECT 154.600 183.100 154.900 183.400 ;
        RECT 156.600 183.100 157.000 183.500 ;
        RECT 151.800 182.800 152.800 183.100 ;
        RECT 152.400 181.100 152.800 182.800 ;
        RECT 154.600 181.100 155.000 183.100 ;
        RECT 156.700 181.100 157.300 183.100 ;
        RECT 159.000 181.100 159.400 185.400 ;
        RECT 160.600 186.100 161.000 187.900 ;
        RECT 162.300 187.200 162.600 187.900 ;
        RECT 163.100 187.700 164.900 187.900 ;
        RECT 164.200 187.200 164.600 187.400 ;
        RECT 162.200 186.800 163.500 187.200 ;
        RECT 164.200 186.900 165.000 187.200 ;
        RECT 164.600 186.800 165.000 186.900 ;
        RECT 160.600 185.800 162.500 186.100 ;
        RECT 160.600 181.100 161.000 185.800 ;
        RECT 162.200 185.200 162.500 185.800 ;
        RECT 161.400 184.400 161.800 185.200 ;
        RECT 162.200 185.100 162.600 185.200 ;
        RECT 163.200 185.100 163.500 186.800 ;
        RECT 163.800 185.800 164.200 186.600 ;
        RECT 162.200 184.800 162.900 185.100 ;
        RECT 163.200 184.800 163.700 185.100 ;
        RECT 162.600 184.200 162.900 184.800 ;
        RECT 162.600 183.800 163.000 184.200 ;
        RECT 163.300 181.100 163.700 184.800 ;
        RECT 165.400 181.100 165.800 189.900 ;
        RECT 166.200 187.800 166.600 188.600 ;
        RECT 167.000 187.700 167.400 189.900 ;
        RECT 169.100 189.200 169.700 189.900 ;
        RECT 169.100 188.900 169.800 189.200 ;
        RECT 171.400 188.900 171.800 189.900 ;
        RECT 173.600 189.200 174.000 189.900 ;
        RECT 173.600 188.900 174.600 189.200 ;
        RECT 169.400 188.500 169.800 188.900 ;
        RECT 171.500 188.600 171.800 188.900 ;
        RECT 171.500 188.300 172.900 188.600 ;
        RECT 172.500 188.200 172.900 188.300 ;
        RECT 173.400 188.200 173.800 188.600 ;
        RECT 174.200 188.500 174.600 188.900 ;
        RECT 168.500 187.700 168.900 187.800 ;
        RECT 167.000 187.400 169.000 187.700 ;
        RECT 167.000 185.700 167.400 187.400 ;
        RECT 168.600 186.800 169.000 187.400 ;
        RECT 170.500 187.100 170.900 187.200 ;
        RECT 173.400 187.100 173.700 188.200 ;
        RECT 175.800 187.500 176.200 189.900 ;
        RECT 177.900 188.200 178.300 189.900 ;
        RECT 177.400 187.900 178.300 188.200 ;
        RECT 175.000 187.100 175.800 187.200 ;
        RECT 170.300 186.800 175.800 187.100 ;
        RECT 176.600 186.800 177.000 187.600 ;
        RECT 169.400 186.400 169.800 186.500 ;
        RECT 167.900 186.100 169.800 186.400 ;
        RECT 170.300 186.100 170.600 186.800 ;
        RECT 173.900 186.700 174.300 186.800 ;
        RECT 173.400 186.200 173.800 186.300 ;
        RECT 174.700 186.200 175.100 186.300 ;
        RECT 171.000 186.100 171.400 186.200 ;
        RECT 167.900 186.000 168.300 186.100 ;
        RECT 170.200 185.800 171.400 186.100 ;
        RECT 172.600 185.900 175.100 186.200 ;
        RECT 177.400 186.100 177.800 187.900 ;
        RECT 179.000 187.800 179.400 189.900 ;
        RECT 179.800 188.000 180.200 189.900 ;
        RECT 181.400 188.000 181.800 189.900 ;
        RECT 179.800 187.900 181.800 188.000 ;
        RECT 182.200 188.500 182.600 189.500 ;
        RECT 179.100 187.200 179.400 187.800 ;
        RECT 179.900 187.700 181.700 187.900 ;
        RECT 182.200 187.400 182.500 188.500 ;
        RECT 184.300 188.000 184.700 189.500 ;
        RECT 187.000 188.500 187.400 189.500 ;
        RECT 184.300 187.700 185.100 188.000 ;
        RECT 184.700 187.500 185.100 187.700 ;
        RECT 181.000 187.200 181.400 187.400 ;
        RECT 179.000 186.800 180.300 187.200 ;
        RECT 181.000 186.900 181.800 187.200 ;
        RECT 182.200 187.100 184.300 187.400 ;
        RECT 181.400 186.800 181.800 186.900 ;
        RECT 183.800 186.900 184.300 187.100 ;
        RECT 184.800 187.200 185.100 187.500 ;
        RECT 187.000 187.400 187.300 188.500 ;
        RECT 189.100 188.000 189.500 189.500 ;
        RECT 193.400 188.500 193.800 189.500 ;
        RECT 189.100 187.700 189.900 188.000 ;
        RECT 189.500 187.500 189.900 187.700 ;
        RECT 172.600 185.800 173.000 185.900 ;
        RECT 177.400 185.800 179.300 186.100 ;
        RECT 168.700 185.700 169.100 185.800 ;
        RECT 167.000 185.400 169.100 185.700 ;
        RECT 167.000 181.100 167.400 185.400 ;
        RECT 170.300 185.200 170.600 185.800 ;
        RECT 173.400 185.500 176.200 185.600 ;
        RECT 173.300 185.400 176.200 185.500 ;
        RECT 169.400 184.900 170.600 185.200 ;
        RECT 171.300 185.300 176.200 185.400 ;
        RECT 171.300 185.100 173.700 185.300 ;
        RECT 169.400 184.400 169.700 184.900 ;
        RECT 169.000 184.000 169.700 184.400 ;
        RECT 170.500 184.500 170.900 184.600 ;
        RECT 171.300 184.500 171.600 185.100 ;
        RECT 170.500 184.200 171.600 184.500 ;
        RECT 171.900 184.500 174.600 184.800 ;
        RECT 171.900 184.400 172.300 184.500 ;
        RECT 174.200 184.400 174.600 184.500 ;
        RECT 171.100 183.700 171.500 183.800 ;
        RECT 172.500 183.700 172.900 183.800 ;
        RECT 169.400 183.100 169.800 183.500 ;
        RECT 171.100 183.400 172.900 183.700 ;
        RECT 171.500 183.100 171.800 183.400 ;
        RECT 174.200 183.100 174.600 183.500 ;
        RECT 169.100 181.100 169.700 183.100 ;
        RECT 171.400 181.100 171.800 183.100 ;
        RECT 173.600 182.800 174.600 183.100 ;
        RECT 173.600 181.100 174.000 182.800 ;
        RECT 175.800 181.100 176.200 185.300 ;
        RECT 177.400 181.100 177.800 185.800 ;
        RECT 179.000 185.200 179.300 185.800 ;
        RECT 178.200 184.400 178.600 185.200 ;
        RECT 179.000 185.100 179.400 185.200 ;
        RECT 180.000 185.100 180.300 186.800 ;
        RECT 180.600 185.800 181.000 186.600 ;
        RECT 182.200 185.800 182.600 186.600 ;
        RECT 183.000 185.800 183.400 186.600 ;
        RECT 183.800 186.500 184.500 186.900 ;
        RECT 184.800 186.800 185.800 187.200 ;
        RECT 187.000 187.100 189.100 187.400 ;
        RECT 188.600 186.900 189.100 187.100 ;
        RECT 189.600 187.200 189.900 187.500 ;
        RECT 193.400 187.400 193.700 188.500 ;
        RECT 195.500 188.000 195.900 189.500 ;
        RECT 198.200 188.500 198.600 189.500 ;
        RECT 195.500 187.700 196.300 188.000 ;
        RECT 195.900 187.500 196.300 187.700 ;
        RECT 183.800 185.500 184.100 186.500 ;
        RECT 182.200 185.200 184.100 185.500 ;
        RECT 179.000 184.800 179.700 185.100 ;
        RECT 180.000 184.800 180.500 185.100 ;
        RECT 179.400 184.200 179.700 184.800 ;
        RECT 179.400 183.800 179.800 184.200 ;
        RECT 180.100 181.100 180.500 184.800 ;
        RECT 182.200 183.500 182.500 185.200 ;
        RECT 184.800 184.900 185.100 186.800 ;
        RECT 185.400 186.100 185.800 186.200 ;
        RECT 186.200 186.100 186.600 186.200 ;
        RECT 185.400 185.800 186.600 186.100 ;
        RECT 187.000 185.800 187.400 186.600 ;
        RECT 187.800 185.800 188.200 186.600 ;
        RECT 188.600 186.500 189.300 186.900 ;
        RECT 189.600 186.800 190.600 187.200 ;
        RECT 193.400 187.100 195.500 187.400 ;
        RECT 195.000 186.900 195.500 187.100 ;
        RECT 196.000 187.200 196.300 187.500 ;
        RECT 198.200 187.400 198.500 188.500 ;
        RECT 200.300 188.000 200.700 189.500 ;
        RECT 203.000 188.500 203.400 189.500 ;
        RECT 200.300 187.700 201.100 188.000 ;
        RECT 200.700 187.500 201.100 187.700 ;
        RECT 185.400 185.400 185.800 185.800 ;
        RECT 188.600 185.500 188.900 186.500 ;
        RECT 184.300 184.600 185.100 184.900 ;
        RECT 187.000 185.200 188.900 185.500 ;
        RECT 182.200 181.500 182.600 183.500 ;
        RECT 184.300 181.100 184.700 184.600 ;
        RECT 187.000 183.500 187.300 185.200 ;
        RECT 189.600 184.900 189.900 186.800 ;
        RECT 190.200 185.400 190.600 186.200 ;
        RECT 193.400 185.800 193.800 186.600 ;
        RECT 194.200 185.800 194.600 186.600 ;
        RECT 195.000 186.500 195.700 186.900 ;
        RECT 196.000 186.800 197.000 187.200 ;
        RECT 198.200 187.100 200.300 187.400 ;
        RECT 199.800 186.900 200.300 187.100 ;
        RECT 200.800 187.200 201.100 187.500 ;
        RECT 203.000 187.400 203.300 188.500 ;
        RECT 205.100 188.200 205.500 189.500 ;
        RECT 204.600 188.000 205.500 188.200 ;
        RECT 204.600 187.800 205.900 188.000 ;
        RECT 205.100 187.700 205.900 187.800 ;
        RECT 205.500 187.500 205.900 187.700 ;
        RECT 195.000 185.500 195.300 186.500 ;
        RECT 189.100 184.600 189.900 184.900 ;
        RECT 193.400 185.200 195.300 185.500 ;
        RECT 187.000 181.500 187.400 183.500 ;
        RECT 189.100 182.200 189.500 184.600 ;
        RECT 193.400 183.500 193.700 185.200 ;
        RECT 196.000 184.900 196.300 186.800 ;
        RECT 196.600 185.400 197.000 186.200 ;
        RECT 198.200 185.800 198.600 186.600 ;
        RECT 199.000 185.800 199.400 186.600 ;
        RECT 199.800 186.500 200.500 186.900 ;
        RECT 200.800 186.800 201.800 187.200 ;
        RECT 203.000 187.100 205.100 187.400 ;
        RECT 204.600 186.900 205.100 187.100 ;
        RECT 205.600 187.200 205.900 187.500 ;
        RECT 207.800 187.700 208.200 189.900 ;
        RECT 209.900 189.200 210.500 189.900 ;
        RECT 209.900 188.900 210.600 189.200 ;
        RECT 212.200 188.900 212.600 189.900 ;
        RECT 214.400 189.200 214.800 189.900 ;
        RECT 214.400 188.900 215.400 189.200 ;
        RECT 210.200 188.500 210.600 188.900 ;
        RECT 212.300 188.600 212.600 188.900 ;
        RECT 212.300 188.300 213.700 188.600 ;
        RECT 213.300 188.200 213.700 188.300 ;
        RECT 214.200 188.200 214.600 188.600 ;
        RECT 215.000 188.500 215.400 188.900 ;
        RECT 209.300 187.700 209.700 187.800 ;
        RECT 207.800 187.400 209.700 187.700 ;
        RECT 199.800 185.500 200.100 186.500 ;
        RECT 195.500 184.600 196.300 184.900 ;
        RECT 198.200 185.200 200.100 185.500 ;
        RECT 189.100 181.800 189.800 182.200 ;
        RECT 189.100 181.100 189.500 181.800 ;
        RECT 193.400 181.500 193.800 183.500 ;
        RECT 195.500 182.200 195.900 184.600 ;
        RECT 195.000 181.800 195.900 182.200 ;
        RECT 195.500 181.100 195.900 181.800 ;
        RECT 198.200 183.500 198.500 185.200 ;
        RECT 200.800 184.900 201.100 186.800 ;
        RECT 201.400 185.400 201.800 186.200 ;
        RECT 203.000 185.800 203.400 186.600 ;
        RECT 203.800 185.800 204.200 186.600 ;
        RECT 204.600 186.500 205.300 186.900 ;
        RECT 205.600 186.800 206.600 187.200 ;
        RECT 204.600 185.500 204.900 186.500 ;
        RECT 200.300 184.600 201.100 184.900 ;
        RECT 203.000 185.200 204.900 185.500 ;
        RECT 198.200 181.500 198.600 183.500 ;
        RECT 200.300 182.200 200.700 184.600 ;
        RECT 199.800 181.800 200.700 182.200 ;
        RECT 200.300 181.100 200.700 181.800 ;
        RECT 203.000 183.500 203.300 185.200 ;
        RECT 205.600 184.900 205.900 186.800 ;
        RECT 206.200 186.100 206.600 186.200 ;
        RECT 207.000 186.100 207.400 186.200 ;
        RECT 206.200 185.800 207.400 186.100 ;
        RECT 206.200 185.400 206.600 185.800 ;
        RECT 207.800 185.700 208.200 187.400 ;
        RECT 211.300 187.100 211.700 187.200 ;
        RECT 214.200 187.100 214.500 188.200 ;
        RECT 216.600 187.500 217.000 189.900 ;
        RECT 218.700 188.200 219.100 189.900 ;
        RECT 218.200 187.900 219.100 188.200 ;
        RECT 219.800 187.900 220.200 189.900 ;
        RECT 220.600 188.000 221.000 189.900 ;
        RECT 222.200 188.000 222.600 189.900 ;
        RECT 224.300 188.200 224.700 189.900 ;
        RECT 220.600 187.900 222.600 188.000 ;
        RECT 223.800 187.900 224.700 188.200 ;
        RECT 225.400 187.900 225.800 189.900 ;
        RECT 226.200 188.000 226.600 189.900 ;
        RECT 227.800 188.000 228.200 189.900 ;
        RECT 226.200 187.900 228.200 188.000 ;
        RECT 215.800 187.100 216.600 187.200 ;
        RECT 211.100 186.800 216.600 187.100 ;
        RECT 217.400 186.800 217.800 187.600 ;
        RECT 210.200 186.400 210.600 186.500 ;
        RECT 208.700 186.100 210.600 186.400 ;
        RECT 211.100 186.200 211.400 186.800 ;
        RECT 214.700 186.700 215.100 186.800 ;
        RECT 214.200 186.200 214.600 186.300 ;
        RECT 215.500 186.200 215.900 186.300 ;
        RECT 208.700 186.000 209.100 186.100 ;
        RECT 211.000 185.800 211.400 186.200 ;
        RECT 213.400 185.900 215.900 186.200 ;
        RECT 218.200 186.100 218.600 187.900 ;
        RECT 219.900 187.200 220.200 187.900 ;
        RECT 220.700 187.700 222.500 187.900 ;
        RECT 221.800 187.200 222.200 187.400 ;
        RECT 219.000 187.100 219.400 187.200 ;
        RECT 219.800 187.100 221.100 187.200 ;
        RECT 219.000 186.800 221.100 187.100 ;
        RECT 221.800 186.900 222.600 187.200 ;
        RECT 222.200 186.800 222.600 186.900 ;
        RECT 223.000 186.800 223.400 187.600 ;
        RECT 213.400 185.800 213.800 185.900 ;
        RECT 218.200 185.800 220.100 186.100 ;
        RECT 209.500 185.700 209.900 185.800 ;
        RECT 207.800 185.400 209.900 185.700 ;
        RECT 205.100 184.600 205.900 184.900 ;
        RECT 203.000 181.500 203.400 183.500 ;
        RECT 205.100 181.100 205.500 184.600 ;
        RECT 207.800 181.100 208.200 185.400 ;
        RECT 211.100 185.200 211.400 185.800 ;
        RECT 214.200 185.500 217.000 185.600 ;
        RECT 214.100 185.400 217.000 185.500 ;
        RECT 210.200 184.900 211.400 185.200 ;
        RECT 212.100 185.300 217.000 185.400 ;
        RECT 212.100 185.100 214.500 185.300 ;
        RECT 210.200 184.400 210.500 184.900 ;
        RECT 209.800 184.000 210.500 184.400 ;
        RECT 211.300 184.500 211.700 184.600 ;
        RECT 212.100 184.500 212.400 185.100 ;
        RECT 211.300 184.200 212.400 184.500 ;
        RECT 212.700 184.500 215.400 184.800 ;
        RECT 212.700 184.400 213.100 184.500 ;
        RECT 215.000 184.400 215.400 184.500 ;
        RECT 211.900 183.700 212.300 183.800 ;
        RECT 213.300 183.700 213.700 183.800 ;
        RECT 210.200 183.100 210.600 183.500 ;
        RECT 211.900 183.400 213.700 183.700 ;
        RECT 212.300 183.100 212.600 183.400 ;
        RECT 215.000 183.100 215.400 183.500 ;
        RECT 209.900 181.100 210.500 183.100 ;
        RECT 212.200 181.100 212.600 183.100 ;
        RECT 214.400 182.800 215.400 183.100 ;
        RECT 214.400 181.100 214.800 182.800 ;
        RECT 216.600 181.100 217.000 185.300 ;
        RECT 218.200 181.100 218.600 185.800 ;
        RECT 219.800 185.200 220.100 185.800 ;
        RECT 219.000 184.400 219.400 185.200 ;
        RECT 219.800 185.100 220.200 185.200 ;
        RECT 220.800 185.100 221.100 186.800 ;
        RECT 221.400 185.800 221.800 186.600 ;
        RECT 223.800 186.100 224.200 187.900 ;
        RECT 225.500 187.200 225.800 187.900 ;
        RECT 226.300 187.700 228.100 187.900 ;
        RECT 227.400 187.200 227.800 187.400 ;
        RECT 225.400 186.800 226.700 187.200 ;
        RECT 227.400 186.900 228.200 187.200 ;
        RECT 227.800 186.800 228.200 186.900 ;
        RECT 223.800 185.800 225.700 186.100 ;
        RECT 219.800 184.800 220.500 185.100 ;
        RECT 220.800 184.800 221.300 185.100 ;
        RECT 220.200 184.200 220.500 184.800 ;
        RECT 220.200 183.800 220.600 184.200 ;
        RECT 220.900 181.100 221.300 184.800 ;
        RECT 223.800 181.100 224.200 185.800 ;
        RECT 225.400 185.200 225.700 185.800 ;
        RECT 224.600 184.400 225.000 185.200 ;
        RECT 225.400 185.100 225.800 185.200 ;
        RECT 226.400 185.100 226.700 186.800 ;
        RECT 227.000 185.800 227.400 186.600 ;
        RECT 225.400 184.800 226.100 185.100 ;
        RECT 226.400 184.800 226.900 185.100 ;
        RECT 225.800 184.200 226.100 184.800 ;
        RECT 225.800 183.800 226.200 184.200 ;
        RECT 226.500 181.100 226.900 184.800 ;
        RECT 1.400 175.600 1.800 179.900 ;
        RECT 3.000 175.600 3.400 179.900 ;
        RECT 4.600 175.600 5.000 179.900 ;
        RECT 6.200 175.600 6.600 179.900 ;
        RECT 7.800 175.600 8.200 179.900 ;
        RECT 9.900 177.900 10.500 179.900 ;
        RECT 12.200 177.900 12.600 179.900 ;
        RECT 14.400 178.200 14.800 179.900 ;
        RECT 14.400 177.900 15.400 178.200 ;
        RECT 10.200 177.500 10.600 177.900 ;
        RECT 12.300 177.600 12.600 177.900 ;
        RECT 11.900 177.300 13.700 177.600 ;
        RECT 15.000 177.500 15.400 177.900 ;
        RECT 11.900 177.200 12.300 177.300 ;
        RECT 13.300 177.200 13.700 177.300 ;
        RECT 9.800 176.600 10.500 177.000 ;
        RECT 10.200 176.100 10.500 176.600 ;
        RECT 11.300 176.500 12.400 176.800 ;
        RECT 11.300 176.400 11.700 176.500 ;
        RECT 10.200 175.800 11.400 176.100 ;
        RECT 1.400 175.200 2.300 175.600 ;
        RECT 3.000 175.200 4.100 175.600 ;
        RECT 4.600 175.200 5.700 175.600 ;
        RECT 6.200 175.200 7.400 175.600 ;
        RECT 1.900 174.500 2.300 175.200 ;
        RECT 3.700 174.500 4.100 175.200 ;
        RECT 5.300 174.500 5.700 175.200 ;
        RECT 1.900 174.100 3.200 174.500 ;
        RECT 3.700 174.100 4.900 174.500 ;
        RECT 5.300 174.100 6.600 174.500 ;
        RECT 1.900 173.800 2.300 174.100 ;
        RECT 3.700 173.800 4.100 174.100 ;
        RECT 5.300 173.800 5.700 174.100 ;
        RECT 7.000 173.800 7.400 175.200 ;
        RECT 1.400 173.400 2.300 173.800 ;
        RECT 3.000 173.400 4.100 173.800 ;
        RECT 4.600 173.400 5.700 173.800 ;
        RECT 6.200 173.400 7.400 173.800 ;
        RECT 7.800 175.300 9.900 175.600 ;
        RECT 7.800 173.600 8.200 175.300 ;
        RECT 9.500 175.200 9.900 175.300 ;
        RECT 11.100 175.200 11.400 175.800 ;
        RECT 12.100 175.900 12.400 176.500 ;
        RECT 12.700 176.500 13.100 176.600 ;
        RECT 15.000 176.500 15.400 176.600 ;
        RECT 12.700 176.200 15.400 176.500 ;
        RECT 12.100 175.700 14.500 175.900 ;
        RECT 16.600 175.700 17.000 179.900 ;
        RECT 12.100 175.600 17.000 175.700 ;
        RECT 14.100 175.500 17.000 175.600 ;
        RECT 14.200 175.400 17.000 175.500 ;
        RECT 18.200 175.600 18.600 179.900 ;
        RECT 19.800 175.600 20.200 179.900 ;
        RECT 21.400 175.600 21.800 179.900 ;
        RECT 23.000 175.600 23.400 179.900 ;
        RECT 24.600 175.700 25.000 179.900 ;
        RECT 26.800 178.200 27.200 179.900 ;
        RECT 26.200 177.900 27.200 178.200 ;
        RECT 29.000 177.900 29.400 179.900 ;
        RECT 31.100 177.900 31.700 179.900 ;
        RECT 26.200 177.500 26.600 177.900 ;
        RECT 29.000 177.600 29.300 177.900 ;
        RECT 27.900 177.300 29.700 177.600 ;
        RECT 31.000 177.500 31.400 177.900 ;
        RECT 27.900 177.200 28.300 177.300 ;
        RECT 29.300 177.200 29.700 177.300 ;
        RECT 26.200 176.500 26.600 176.600 ;
        RECT 28.500 176.500 28.900 176.600 ;
        RECT 26.200 176.200 28.900 176.500 ;
        RECT 29.200 176.500 30.300 176.800 ;
        RECT 29.200 175.900 29.500 176.500 ;
        RECT 29.900 176.400 30.300 176.500 ;
        RECT 31.100 176.600 31.800 177.000 ;
        RECT 31.100 176.100 31.400 176.600 ;
        RECT 27.100 175.700 29.500 175.900 ;
        RECT 24.600 175.600 29.500 175.700 ;
        RECT 30.200 175.800 31.400 176.100 ;
        RECT 18.200 175.200 19.100 175.600 ;
        RECT 19.800 175.200 20.900 175.600 ;
        RECT 21.400 175.200 22.500 175.600 ;
        RECT 23.000 175.200 24.200 175.600 ;
        RECT 24.600 175.500 27.500 175.600 ;
        RECT 24.600 175.400 27.400 175.500 ;
        RECT 8.700 174.900 9.100 175.000 ;
        RECT 8.700 174.600 10.600 174.900 ;
        RECT 11.000 174.800 11.400 175.200 ;
        RECT 13.400 175.100 13.800 175.200 ;
        RECT 13.400 174.800 15.900 175.100 ;
        RECT 10.200 174.500 10.600 174.600 ;
        RECT 11.100 174.200 11.400 174.800 ;
        RECT 14.200 174.700 14.600 174.800 ;
        RECT 15.500 174.700 15.900 174.800 ;
        RECT 18.700 174.500 19.100 175.200 ;
        RECT 20.500 174.500 20.900 175.200 ;
        RECT 22.100 174.500 22.500 175.200 ;
        RECT 14.700 174.200 15.100 174.300 ;
        RECT 11.100 173.900 16.600 174.200 ;
        RECT 11.300 173.800 11.700 173.900 ;
        RECT 1.400 171.100 1.800 173.400 ;
        RECT 3.000 171.100 3.400 173.400 ;
        RECT 4.600 171.100 5.000 173.400 ;
        RECT 6.200 171.100 6.600 173.400 ;
        RECT 7.800 173.300 9.700 173.600 ;
        RECT 7.800 171.100 8.200 173.300 ;
        RECT 9.300 173.200 9.700 173.300 ;
        RECT 14.200 172.800 14.500 173.900 ;
        RECT 15.800 173.800 16.600 173.900 ;
        RECT 18.700 174.100 20.000 174.500 ;
        RECT 20.500 174.100 21.700 174.500 ;
        RECT 22.100 174.100 23.400 174.500 ;
        RECT 18.700 173.800 19.100 174.100 ;
        RECT 20.500 173.800 20.900 174.100 ;
        RECT 22.100 173.800 22.500 174.100 ;
        RECT 23.800 173.800 24.200 175.200 ;
        RECT 27.800 175.100 28.200 175.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 25.700 174.800 29.000 175.100 ;
        RECT 25.700 174.700 26.100 174.800 ;
        RECT 26.500 174.200 26.900 174.300 ;
        RECT 30.200 174.200 30.500 175.800 ;
        RECT 33.400 175.600 33.800 179.900 ;
        RECT 34.600 176.800 35.000 177.200 ;
        RECT 34.600 176.200 34.900 176.800 ;
        RECT 35.300 176.200 35.700 179.900 ;
        RECT 40.900 176.400 41.300 179.900 ;
        RECT 43.000 177.500 43.400 179.500 ;
        RECT 34.200 175.900 34.900 176.200 ;
        RECT 35.200 175.900 35.700 176.200 ;
        RECT 40.500 176.100 41.300 176.400 ;
        RECT 34.200 175.800 34.600 175.900 ;
        RECT 31.700 175.300 33.800 175.600 ;
        RECT 31.700 175.200 32.100 175.300 ;
        RECT 32.500 174.900 32.900 175.000 ;
        RECT 31.000 174.600 32.900 174.900 ;
        RECT 31.000 174.500 31.400 174.600 ;
        RECT 25.000 173.900 30.500 174.200 ;
        RECT 25.000 173.800 25.800 173.900 ;
        RECT 13.300 172.700 13.700 172.800 ;
        RECT 10.200 172.100 10.600 172.500 ;
        RECT 12.300 172.400 13.700 172.700 ;
        RECT 14.200 172.400 14.600 172.800 ;
        RECT 12.300 172.100 12.600 172.400 ;
        RECT 15.000 172.100 15.400 172.500 ;
        RECT 9.900 171.800 10.600 172.100 ;
        RECT 9.900 171.100 10.500 171.800 ;
        RECT 12.200 171.100 12.600 172.100 ;
        RECT 14.400 171.800 15.400 172.100 ;
        RECT 14.400 171.100 14.800 171.800 ;
        RECT 16.600 171.100 17.000 173.500 ;
        RECT 18.200 173.400 19.100 173.800 ;
        RECT 19.800 173.400 20.900 173.800 ;
        RECT 21.400 173.400 22.500 173.800 ;
        RECT 23.000 173.400 24.200 173.800 ;
        RECT 18.200 171.100 18.600 173.400 ;
        RECT 19.800 171.100 20.200 173.400 ;
        RECT 21.400 171.100 21.800 173.400 ;
        RECT 23.000 171.100 23.400 173.400 ;
        RECT 24.600 171.100 25.000 173.500 ;
        RECT 27.100 172.800 27.400 173.900 ;
        RECT 29.900 173.800 30.300 173.900 ;
        RECT 33.400 173.600 33.800 175.300 ;
        RECT 34.200 175.100 34.600 175.200 ;
        RECT 35.200 175.100 35.500 175.900 ;
        RECT 34.200 174.800 35.500 175.100 ;
        RECT 35.200 174.200 35.500 174.800 ;
        RECT 35.800 174.400 36.200 175.200 ;
        RECT 39.800 174.800 40.200 175.600 ;
        RECT 40.500 174.200 40.800 176.100 ;
        RECT 43.100 175.800 43.400 177.500 ;
        RECT 41.500 175.500 43.400 175.800 ;
        RECT 43.800 175.700 44.200 179.900 ;
        RECT 46.000 178.200 46.400 179.900 ;
        RECT 45.400 177.900 46.400 178.200 ;
        RECT 48.200 177.900 48.600 179.900 ;
        RECT 50.300 177.900 50.900 179.900 ;
        RECT 45.400 177.500 45.800 177.900 ;
        RECT 48.200 177.600 48.500 177.900 ;
        RECT 47.100 177.300 48.900 177.600 ;
        RECT 50.200 177.500 50.600 177.900 ;
        RECT 47.100 177.200 47.500 177.300 ;
        RECT 48.500 177.200 48.900 177.300 ;
        RECT 45.400 176.500 45.800 176.600 ;
        RECT 47.700 176.500 48.100 176.600 ;
        RECT 45.400 176.200 48.100 176.500 ;
        RECT 48.400 176.500 49.500 176.800 ;
        RECT 48.400 175.900 48.700 176.500 ;
        RECT 49.100 176.400 49.500 176.500 ;
        RECT 50.300 176.600 51.000 177.000 ;
        RECT 50.300 176.100 50.600 176.600 ;
        RECT 46.300 175.700 48.700 175.900 ;
        RECT 43.800 175.600 48.700 175.700 ;
        RECT 49.400 175.800 50.600 176.100 ;
        RECT 43.800 175.500 46.700 175.600 ;
        RECT 41.500 174.500 41.800 175.500 ;
        RECT 43.800 175.400 46.600 175.500 ;
        RECT 34.200 173.800 35.500 174.200 ;
        RECT 36.600 174.100 37.000 174.200 ;
        RECT 36.200 173.800 37.000 174.100 ;
        RECT 39.800 173.800 40.800 174.200 ;
        RECT 41.100 174.100 41.800 174.500 ;
        RECT 42.200 174.400 42.600 175.200 ;
        RECT 43.000 174.400 43.400 175.200 ;
        RECT 47.000 175.100 47.400 175.200 ;
        RECT 47.800 175.100 48.200 175.200 ;
        RECT 44.900 174.800 48.200 175.100 ;
        RECT 44.900 174.700 45.300 174.800 ;
        RECT 45.700 174.200 46.100 174.300 ;
        RECT 49.400 174.200 49.700 175.800 ;
        RECT 52.600 175.600 53.000 179.900 ;
        RECT 54.700 176.200 55.100 179.900 ;
        RECT 55.400 176.800 55.800 177.200 ;
        RECT 55.500 176.200 55.800 176.800 ;
        RECT 57.000 176.800 57.400 177.200 ;
        RECT 57.000 176.200 57.300 176.800 ;
        RECT 57.700 176.200 58.100 179.900 ;
        RECT 54.700 175.900 55.200 176.200 ;
        RECT 55.500 175.900 56.200 176.200 ;
        RECT 50.900 175.300 53.000 175.600 ;
        RECT 50.900 175.200 51.300 175.300 ;
        RECT 51.700 174.900 52.100 175.000 ;
        RECT 50.200 174.600 52.100 174.900 ;
        RECT 50.200 174.500 50.600 174.600 ;
        RECT 31.900 173.300 33.800 173.600 ;
        RECT 31.900 173.200 32.300 173.300 ;
        RECT 26.200 172.100 26.600 172.500 ;
        RECT 27.000 172.400 27.400 172.800 ;
        RECT 27.900 172.700 28.300 172.800 ;
        RECT 27.900 172.400 29.300 172.700 ;
        RECT 29.000 172.100 29.300 172.400 ;
        RECT 31.000 172.100 31.400 172.500 ;
        RECT 26.200 171.800 27.200 172.100 ;
        RECT 26.800 171.100 27.200 171.800 ;
        RECT 29.000 171.100 29.400 172.100 ;
        RECT 31.000 171.800 31.700 172.100 ;
        RECT 31.100 171.100 31.700 171.800 ;
        RECT 33.400 171.100 33.800 173.300 ;
        RECT 34.300 173.100 34.600 173.800 ;
        RECT 36.200 173.600 36.600 173.800 ;
        RECT 40.500 173.500 40.800 173.800 ;
        RECT 41.300 173.900 41.800 174.100 ;
        RECT 44.200 173.900 49.700 174.200 ;
        RECT 41.300 173.600 43.400 173.900 ;
        RECT 44.200 173.800 45.000 173.900 ;
        RECT 46.200 173.800 46.600 173.900 ;
        RECT 49.100 173.800 49.500 173.900 ;
        RECT 40.500 173.300 40.900 173.500 ;
        RECT 35.100 173.100 36.900 173.300 ;
        RECT 34.200 171.100 34.600 173.100 ;
        RECT 35.000 173.000 37.000 173.100 ;
        RECT 40.500 173.000 41.300 173.300 ;
        RECT 35.000 171.100 35.400 173.000 ;
        RECT 36.600 171.100 37.000 173.000 ;
        RECT 40.900 172.200 41.300 173.000 ;
        RECT 43.100 172.500 43.400 173.600 ;
        RECT 40.900 171.800 41.800 172.200 ;
        RECT 40.900 171.500 41.300 171.800 ;
        RECT 43.000 171.500 43.400 172.500 ;
        RECT 43.800 171.100 44.200 173.500 ;
        RECT 46.300 172.800 46.600 173.800 ;
        RECT 52.600 173.600 53.000 175.300 ;
        RECT 54.900 175.200 55.200 175.900 ;
        RECT 55.800 175.800 56.200 175.900 ;
        RECT 56.600 175.900 57.300 176.200 ;
        RECT 57.600 175.900 58.100 176.200 ;
        RECT 59.800 177.500 60.200 179.500 ;
        RECT 61.900 179.200 62.300 179.900 ;
        RECT 61.900 178.800 62.600 179.200 ;
        RECT 56.600 175.800 57.000 175.900 ;
        RECT 54.200 174.400 54.600 175.200 ;
        RECT 54.900 174.800 55.400 175.200 ;
        RECT 55.800 175.100 56.100 175.800 ;
        RECT 57.600 175.100 57.900 175.900 ;
        RECT 59.800 175.800 60.100 177.500 ;
        RECT 61.900 176.400 62.300 178.800 ;
        RECT 66.500 176.400 66.900 179.900 ;
        RECT 68.600 177.500 69.000 179.500 ;
        RECT 61.900 176.100 62.700 176.400 ;
        RECT 59.800 175.500 61.700 175.800 ;
        RECT 55.800 174.800 57.900 175.100 ;
        RECT 54.900 174.200 55.200 174.800 ;
        RECT 57.600 174.200 57.900 174.800 ;
        RECT 58.200 174.400 58.600 175.200 ;
        RECT 59.800 174.400 60.200 175.200 ;
        RECT 60.600 174.400 61.000 175.200 ;
        RECT 61.400 174.500 61.700 175.500 ;
        RECT 53.400 174.100 53.800 174.200 ;
        RECT 53.400 173.800 54.200 174.100 ;
        RECT 54.900 173.800 56.200 174.200 ;
        RECT 56.600 173.800 57.900 174.200 ;
        RECT 59.000 174.100 59.400 174.200 ;
        RECT 58.600 173.800 59.400 174.100 ;
        RECT 61.400 174.100 62.100 174.500 ;
        RECT 62.400 174.200 62.700 176.100 ;
        RECT 66.100 176.100 66.900 176.400 ;
        RECT 63.000 174.800 63.400 175.600 ;
        RECT 65.400 174.800 65.800 175.600 ;
        RECT 66.100 175.200 66.400 176.100 ;
        RECT 68.700 175.800 69.000 177.500 ;
        RECT 67.100 175.500 69.000 175.800 ;
        RECT 69.400 177.500 69.800 179.500 ;
        RECT 69.400 175.800 69.700 177.500 ;
        RECT 71.500 176.400 71.900 179.900 ;
        RECT 71.500 176.100 72.300 176.400 ;
        RECT 69.400 175.500 71.300 175.800 ;
        RECT 66.100 174.800 66.600 175.200 ;
        RECT 66.100 174.200 66.400 174.800 ;
        RECT 67.100 174.500 67.400 175.500 ;
        RECT 61.400 173.900 61.900 174.100 ;
        RECT 53.800 173.600 54.200 173.800 ;
        RECT 51.100 173.300 53.000 173.600 ;
        RECT 51.100 173.200 51.500 173.300 ;
        RECT 45.400 172.100 45.800 172.500 ;
        RECT 46.200 172.400 46.600 172.800 ;
        RECT 47.100 172.700 47.500 172.800 ;
        RECT 47.100 172.400 48.500 172.700 ;
        RECT 48.200 172.100 48.500 172.400 ;
        RECT 50.200 172.100 50.600 172.500 ;
        RECT 45.400 171.800 46.400 172.100 ;
        RECT 46.000 171.100 46.400 171.800 ;
        RECT 48.200 171.100 48.600 172.100 ;
        RECT 50.200 171.800 50.900 172.100 ;
        RECT 50.300 171.100 50.900 171.800 ;
        RECT 52.600 171.100 53.000 173.300 ;
        RECT 53.500 173.100 55.300 173.300 ;
        RECT 55.800 173.100 56.100 173.800 ;
        RECT 56.700 173.100 57.000 173.800 ;
        RECT 58.600 173.600 59.000 173.800 ;
        RECT 59.800 173.600 61.900 173.900 ;
        RECT 62.400 173.800 63.400 174.200 ;
        RECT 65.400 173.800 66.400 174.200 ;
        RECT 66.700 174.100 67.400 174.500 ;
        RECT 67.800 174.400 68.200 175.200 ;
        RECT 68.600 174.400 69.000 175.200 ;
        RECT 69.400 174.400 69.800 175.200 ;
        RECT 70.200 174.400 70.600 175.200 ;
        RECT 71.000 174.500 71.300 175.500 ;
        RECT 57.500 173.100 59.300 173.300 ;
        RECT 53.400 173.000 55.400 173.100 ;
        RECT 53.400 171.100 53.800 173.000 ;
        RECT 55.000 171.100 55.400 173.000 ;
        RECT 55.800 171.100 56.200 173.100 ;
        RECT 56.600 171.100 57.000 173.100 ;
        RECT 57.400 173.000 59.400 173.100 ;
        RECT 57.400 171.100 57.800 173.000 ;
        RECT 59.000 171.100 59.400 173.000 ;
        RECT 59.800 172.500 60.100 173.600 ;
        RECT 62.400 173.500 62.700 173.800 ;
        RECT 62.300 173.300 62.700 173.500 ;
        RECT 61.900 173.000 62.700 173.300 ;
        RECT 66.100 173.500 66.400 173.800 ;
        RECT 66.900 173.900 67.400 174.100 ;
        RECT 71.000 174.100 71.700 174.500 ;
        RECT 72.000 174.200 72.300 176.100 ;
        RECT 74.200 176.200 74.600 179.900 ;
        RECT 75.800 176.400 76.200 179.900 ;
        RECT 74.200 175.900 75.500 176.200 ;
        RECT 75.800 175.900 76.300 176.400 ;
        RECT 72.600 174.800 73.000 175.600 ;
        RECT 73.400 175.100 73.800 175.200 ;
        RECT 74.200 175.100 74.700 175.200 ;
        RECT 73.400 174.800 74.700 175.100 ;
        RECT 74.300 174.400 74.700 174.800 ;
        RECT 75.200 174.900 75.500 175.900 ;
        RECT 75.200 174.500 75.700 174.900 ;
        RECT 71.000 173.900 71.500 174.100 ;
        RECT 66.900 173.600 69.000 173.900 ;
        RECT 66.100 173.300 66.500 173.500 ;
        RECT 66.100 173.000 66.900 173.300 ;
        RECT 59.800 171.500 60.200 172.500 ;
        RECT 61.900 171.500 62.300 173.000 ;
        RECT 66.500 171.500 66.900 173.000 ;
        RECT 68.700 172.500 69.000 173.600 ;
        RECT 68.600 171.500 69.000 172.500 ;
        RECT 69.400 173.600 71.500 173.900 ;
        RECT 72.000 173.800 73.000 174.200 ;
        RECT 69.400 172.500 69.700 173.600 ;
        RECT 72.000 173.500 72.300 173.800 ;
        RECT 75.200 173.700 75.500 174.500 ;
        RECT 76.000 174.200 76.300 175.900 ;
        RECT 77.400 175.700 77.800 179.900 ;
        RECT 79.600 178.200 80.000 179.900 ;
        RECT 79.000 177.900 80.000 178.200 ;
        RECT 81.800 177.900 82.200 179.900 ;
        RECT 83.900 177.900 84.500 179.900 ;
        RECT 79.000 177.500 79.400 177.900 ;
        RECT 81.800 177.600 82.100 177.900 ;
        RECT 80.700 177.300 82.500 177.600 ;
        RECT 83.800 177.500 84.200 177.900 ;
        RECT 80.700 177.200 81.100 177.300 ;
        RECT 82.100 177.200 82.500 177.300 ;
        RECT 79.000 176.500 79.400 176.600 ;
        RECT 81.300 176.500 81.700 176.600 ;
        RECT 79.000 176.200 81.700 176.500 ;
        RECT 82.000 176.500 83.100 176.800 ;
        RECT 82.000 175.900 82.300 176.500 ;
        RECT 82.700 176.400 83.100 176.500 ;
        RECT 83.900 176.600 84.600 177.000 ;
        RECT 83.900 176.100 84.200 176.600 ;
        RECT 79.900 175.700 82.300 175.900 ;
        RECT 77.400 175.600 82.300 175.700 ;
        RECT 83.000 175.800 84.200 176.100 ;
        RECT 77.400 175.500 80.300 175.600 ;
        RECT 77.400 175.400 80.200 175.500 ;
        RECT 80.600 175.100 81.000 175.200 ;
        RECT 82.200 175.100 82.600 175.200 ;
        RECT 78.500 174.800 82.600 175.100 ;
        RECT 78.500 174.700 78.900 174.800 ;
        RECT 79.300 174.200 79.700 174.300 ;
        RECT 83.000 174.200 83.300 175.800 ;
        RECT 86.200 175.600 86.600 179.900 ;
        RECT 88.300 176.200 88.700 179.900 ;
        RECT 89.000 176.800 89.400 177.200 ;
        RECT 89.100 176.200 89.400 176.800 ;
        RECT 92.200 176.800 92.600 177.200 ;
        RECT 92.200 176.200 92.500 176.800 ;
        RECT 92.900 176.200 93.300 179.900 ;
        RECT 88.300 175.900 88.800 176.200 ;
        RECT 89.100 175.900 89.800 176.200 ;
        RECT 84.500 175.300 86.600 175.600 ;
        RECT 84.500 175.200 84.900 175.300 ;
        RECT 85.300 174.900 85.700 175.000 ;
        RECT 83.800 174.600 85.700 174.900 ;
        RECT 83.800 174.500 84.200 174.600 ;
        RECT 75.800 173.800 76.300 174.200 ;
        RECT 77.800 173.900 83.300 174.200 ;
        RECT 77.800 173.800 78.600 173.900 ;
        RECT 71.900 173.300 72.300 173.500 ;
        RECT 71.500 173.000 72.300 173.300 ;
        RECT 74.200 173.400 75.500 173.700 ;
        RECT 69.400 171.500 69.800 172.500 ;
        RECT 71.500 172.200 71.900 173.000 ;
        RECT 71.500 171.800 72.200 172.200 ;
        RECT 71.500 171.500 71.900 171.800 ;
        RECT 74.200 171.100 74.600 173.400 ;
        RECT 76.000 173.100 76.300 173.800 ;
        RECT 75.800 172.800 76.300 173.100 ;
        RECT 75.800 171.100 76.200 172.800 ;
        RECT 77.400 171.100 77.800 173.500 ;
        RECT 79.900 172.800 80.200 173.900 ;
        RECT 82.700 173.800 83.100 173.900 ;
        RECT 86.200 173.600 86.600 175.300 ;
        RECT 88.500 175.200 88.800 175.900 ;
        RECT 89.400 175.800 89.800 175.900 ;
        RECT 91.800 175.900 92.500 176.200 ;
        RECT 92.800 175.900 93.300 176.200 ;
        RECT 91.800 175.800 92.200 175.900 ;
        RECT 87.800 174.400 88.200 175.200 ;
        RECT 88.500 174.800 89.000 175.200 ;
        RECT 89.400 175.100 89.700 175.800 ;
        RECT 92.800 175.100 93.100 175.900 ;
        RECT 95.800 175.600 96.200 179.900 ;
        RECT 97.400 175.600 97.800 179.900 ;
        RECT 95.800 175.200 97.800 175.600 ;
        RECT 89.400 174.800 93.100 175.100 ;
        RECT 88.500 174.200 88.800 174.800 ;
        RECT 92.800 174.200 93.100 174.800 ;
        RECT 93.400 174.400 93.800 175.200 ;
        RECT 87.000 174.100 87.400 174.200 ;
        RECT 87.000 173.800 87.800 174.100 ;
        RECT 88.500 173.800 89.800 174.200 ;
        RECT 91.800 173.800 93.100 174.200 ;
        RECT 94.200 174.100 94.600 174.200 ;
        RECT 93.800 173.800 94.600 174.100 ;
        RECT 95.800 173.800 96.200 175.200 ;
        RECT 98.200 174.100 98.600 174.200 ;
        RECT 99.000 174.100 99.400 174.200 ;
        RECT 98.200 173.800 99.400 174.100 ;
        RECT 87.400 173.600 87.800 173.800 ;
        RECT 84.700 173.300 86.600 173.600 ;
        RECT 84.700 173.200 85.100 173.300 ;
        RECT 79.000 172.100 79.400 172.500 ;
        RECT 79.800 172.400 80.200 172.800 ;
        RECT 80.700 172.700 81.100 172.800 ;
        RECT 80.700 172.400 82.100 172.700 ;
        RECT 81.800 172.100 82.100 172.400 ;
        RECT 83.800 172.100 84.200 172.500 ;
        RECT 79.000 171.800 80.000 172.100 ;
        RECT 79.600 171.100 80.000 171.800 ;
        RECT 81.800 171.100 82.200 172.100 ;
        RECT 83.800 171.800 84.500 172.100 ;
        RECT 83.900 171.100 84.500 171.800 ;
        RECT 86.200 171.100 86.600 173.300 ;
        RECT 87.100 173.100 88.900 173.300 ;
        RECT 89.400 173.100 89.700 173.800 ;
        RECT 91.900 173.100 92.200 173.800 ;
        RECT 93.800 173.600 94.200 173.800 ;
        RECT 95.800 173.400 97.800 173.800 ;
        RECT 98.200 173.400 98.600 173.800 ;
        RECT 99.000 173.400 99.400 173.800 ;
        RECT 99.800 174.100 100.200 179.900 ;
        RECT 100.600 175.800 101.000 176.600 ;
        RECT 100.600 174.800 101.000 175.200 ;
        RECT 100.600 174.100 100.900 174.800 ;
        RECT 99.800 173.800 100.900 174.100 ;
        RECT 92.700 173.100 94.500 173.300 ;
        RECT 87.000 173.000 89.000 173.100 ;
        RECT 87.000 171.100 87.400 173.000 ;
        RECT 88.600 171.100 89.000 173.000 ;
        RECT 89.400 171.100 89.800 173.100 ;
        RECT 91.800 171.100 92.200 173.100 ;
        RECT 92.600 173.000 94.600 173.100 ;
        RECT 92.600 171.100 93.000 173.000 ;
        RECT 94.200 171.100 94.600 173.000 ;
        RECT 95.800 171.100 96.200 173.400 ;
        RECT 97.400 171.100 97.800 173.400 ;
        RECT 99.800 173.100 100.200 173.800 ;
        RECT 101.400 173.400 101.800 174.200 ;
        RECT 99.800 172.800 100.700 173.100 ;
        RECT 100.300 171.100 100.700 172.800 ;
        RECT 102.200 171.100 102.600 179.900 ;
        RECT 105.100 176.200 105.500 179.900 ;
        RECT 105.800 176.800 106.200 177.200 ;
        RECT 105.900 176.200 106.200 176.800 ;
        RECT 107.400 176.800 107.800 177.200 ;
        RECT 107.400 176.200 107.700 176.800 ;
        RECT 108.100 176.200 108.500 179.900 ;
        RECT 105.100 175.900 105.600 176.200 ;
        RECT 105.900 175.900 106.600 176.200 ;
        RECT 104.600 174.400 105.000 175.200 ;
        RECT 105.300 175.100 105.600 175.900 ;
        RECT 106.200 175.800 106.600 175.900 ;
        RECT 107.000 175.900 107.700 176.200 ;
        RECT 108.000 175.900 108.500 176.200 ;
        RECT 111.500 176.200 111.900 179.900 ;
        RECT 112.200 176.800 112.600 177.200 ;
        RECT 112.300 176.200 112.600 176.800 ;
        RECT 114.700 176.200 115.100 179.900 ;
        RECT 115.400 176.800 116.200 177.200 ;
        RECT 115.500 176.200 115.800 176.800 ;
        RECT 111.500 175.900 112.000 176.200 ;
        RECT 112.300 175.900 113.000 176.200 ;
        RECT 107.000 175.800 107.400 175.900 ;
        RECT 107.000 175.100 107.300 175.800 ;
        RECT 105.300 174.800 107.300 175.100 ;
        RECT 105.300 174.200 105.600 174.800 ;
        RECT 108.000 174.200 108.300 175.900 ;
        RECT 108.600 174.400 109.000 175.200 ;
        RECT 111.000 174.400 111.400 175.200 ;
        RECT 111.700 174.200 112.000 175.900 ;
        RECT 112.600 175.800 113.000 175.900 ;
        RECT 114.200 175.800 115.200 176.200 ;
        RECT 115.500 175.900 116.200 176.200 ;
        RECT 115.800 175.800 116.200 175.900 ;
        RECT 114.200 174.400 114.600 175.200 ;
        RECT 114.900 174.200 115.200 175.800 ;
        RECT 116.600 175.700 117.000 179.900 ;
        RECT 118.800 178.200 119.200 179.900 ;
        RECT 118.200 177.900 119.200 178.200 ;
        RECT 121.000 177.900 121.400 179.900 ;
        RECT 123.100 177.900 123.700 179.900 ;
        RECT 118.200 177.500 118.600 177.900 ;
        RECT 121.000 177.600 121.300 177.900 ;
        RECT 119.900 177.300 121.700 177.600 ;
        RECT 123.000 177.500 123.400 177.900 ;
        RECT 119.900 177.200 120.300 177.300 ;
        RECT 121.300 177.200 121.700 177.300 ;
        RECT 118.200 176.500 118.600 176.600 ;
        RECT 120.500 176.500 120.900 176.600 ;
        RECT 118.200 176.200 120.900 176.500 ;
        RECT 121.200 176.500 122.300 176.800 ;
        RECT 121.200 175.900 121.500 176.500 ;
        RECT 121.900 176.400 122.300 176.500 ;
        RECT 123.100 176.600 123.800 177.000 ;
        RECT 123.100 176.100 123.400 176.600 ;
        RECT 119.100 175.700 121.500 175.900 ;
        RECT 116.600 175.600 121.500 175.700 ;
        RECT 122.200 175.800 123.400 176.100 ;
        RECT 116.600 175.500 119.500 175.600 ;
        RECT 116.600 175.400 119.400 175.500 ;
        RECT 119.800 175.100 120.200 175.200 ;
        RECT 117.700 174.800 120.200 175.100 ;
        RECT 117.700 174.700 118.100 174.800 ;
        RECT 119.000 174.700 119.400 174.800 ;
        RECT 118.500 174.200 118.900 174.300 ;
        RECT 122.200 174.200 122.500 175.800 ;
        RECT 125.400 175.600 125.800 179.900 ;
        RECT 128.100 176.400 128.500 179.900 ;
        RECT 130.200 177.500 130.600 179.500 ;
        RECT 127.700 176.100 128.500 176.400 ;
        RECT 123.700 175.300 125.800 175.600 ;
        RECT 123.700 175.200 124.100 175.300 ;
        RECT 125.400 175.100 125.800 175.300 ;
        RECT 127.000 175.100 127.400 175.600 ;
        RECT 124.500 174.900 124.900 175.000 ;
        RECT 123.000 174.600 124.900 174.900 ;
        RECT 125.400 174.800 127.400 175.100 ;
        RECT 123.000 174.500 123.400 174.600 ;
        RECT 103.800 174.100 104.200 174.200 ;
        RECT 103.800 173.800 104.600 174.100 ;
        RECT 105.300 173.800 106.600 174.200 ;
        RECT 107.000 173.800 108.300 174.200 ;
        RECT 109.400 174.100 109.800 174.200 ;
        RECT 109.000 173.800 109.800 174.100 ;
        RECT 110.200 174.100 110.600 174.200 ;
        RECT 110.200 173.800 111.000 174.100 ;
        RECT 111.700 173.800 113.000 174.200 ;
        RECT 113.400 174.100 113.800 174.200 ;
        RECT 113.400 173.800 114.200 174.100 ;
        RECT 114.900 173.800 116.200 174.200 ;
        RECT 117.000 173.900 122.500 174.200 ;
        RECT 117.000 173.800 117.800 173.900 ;
        RECT 104.200 173.600 104.600 173.800 ;
        RECT 103.900 173.100 105.700 173.300 ;
        RECT 106.200 173.100 106.500 173.800 ;
        RECT 107.100 173.100 107.400 173.800 ;
        RECT 109.000 173.600 109.400 173.800 ;
        RECT 110.600 173.600 111.000 173.800 ;
        RECT 107.900 173.100 109.700 173.300 ;
        RECT 110.300 173.100 112.100 173.300 ;
        RECT 112.600 173.100 112.900 173.800 ;
        RECT 113.800 173.600 114.200 173.800 ;
        RECT 113.500 173.100 115.300 173.300 ;
        RECT 115.800 173.100 116.100 173.800 ;
        RECT 103.800 173.000 105.800 173.100 ;
        RECT 103.800 171.100 104.200 173.000 ;
        RECT 105.400 171.100 105.800 173.000 ;
        RECT 106.200 171.100 106.600 173.100 ;
        RECT 107.000 171.100 107.400 173.100 ;
        RECT 107.800 173.000 109.800 173.100 ;
        RECT 107.800 171.100 108.200 173.000 ;
        RECT 109.400 171.100 109.800 173.000 ;
        RECT 110.200 173.000 112.200 173.100 ;
        RECT 110.200 171.100 110.600 173.000 ;
        RECT 111.800 171.100 112.200 173.000 ;
        RECT 112.600 171.100 113.000 173.100 ;
        RECT 113.400 173.000 115.400 173.100 ;
        RECT 113.400 171.100 113.800 173.000 ;
        RECT 115.000 171.100 115.400 173.000 ;
        RECT 115.800 171.100 116.200 173.100 ;
        RECT 116.600 171.100 117.000 173.500 ;
        RECT 119.100 172.800 119.400 173.900 ;
        RECT 119.800 173.800 120.200 173.900 ;
        RECT 121.900 173.800 122.300 173.900 ;
        RECT 125.400 173.600 125.800 174.800 ;
        RECT 127.700 174.200 128.000 176.100 ;
        RECT 130.300 175.800 130.600 177.500 ;
        RECT 131.000 175.800 131.400 176.600 ;
        RECT 128.700 175.500 130.600 175.800 ;
        RECT 128.700 174.500 129.000 175.500 ;
        RECT 127.000 173.800 128.000 174.200 ;
        RECT 128.300 174.100 129.000 174.500 ;
        RECT 129.400 174.400 129.800 175.200 ;
        RECT 130.200 174.400 130.600 175.200 ;
        RECT 123.900 173.300 125.800 173.600 ;
        RECT 123.900 173.200 124.300 173.300 ;
        RECT 118.200 172.100 118.600 172.500 ;
        RECT 119.000 172.400 119.400 172.800 ;
        RECT 119.900 172.700 120.300 172.800 ;
        RECT 119.900 172.400 121.300 172.700 ;
        RECT 121.000 172.100 121.300 172.400 ;
        RECT 123.000 172.100 123.400 172.500 ;
        RECT 118.200 171.800 119.200 172.100 ;
        RECT 118.800 171.100 119.200 171.800 ;
        RECT 121.000 171.100 121.400 172.100 ;
        RECT 123.000 171.800 123.700 172.100 ;
        RECT 123.100 171.100 123.700 171.800 ;
        RECT 125.400 171.100 125.800 173.300 ;
        RECT 127.700 173.500 128.000 173.800 ;
        RECT 128.500 173.900 129.000 174.100 ;
        RECT 128.500 173.600 130.600 173.900 ;
        RECT 127.700 173.300 128.100 173.500 ;
        RECT 127.700 173.000 128.500 173.300 ;
        RECT 128.100 172.200 128.500 173.000 ;
        RECT 130.300 172.500 130.600 173.600 ;
        RECT 131.800 173.100 132.200 179.900 ;
        RECT 135.300 176.400 135.700 179.900 ;
        RECT 137.400 177.500 137.800 179.500 ;
        RECT 134.900 176.100 135.700 176.400 ;
        RECT 133.400 175.100 133.800 175.200 ;
        RECT 134.200 175.100 134.600 175.600 ;
        RECT 133.400 174.800 134.600 175.100 ;
        RECT 134.900 174.200 135.200 176.100 ;
        RECT 137.500 175.800 137.800 177.500 ;
        RECT 139.500 176.200 139.900 179.900 ;
        RECT 140.200 176.800 140.600 177.200 ;
        RECT 140.300 176.200 140.600 176.800 ;
        RECT 139.500 175.900 140.000 176.200 ;
        RECT 140.300 176.100 141.000 176.200 ;
        RECT 141.400 176.100 141.800 176.200 ;
        RECT 140.300 175.900 141.800 176.100 ;
        RECT 135.900 175.500 137.800 175.800 ;
        RECT 135.900 174.500 136.200 175.500 ;
        RECT 132.600 173.400 133.000 174.200 ;
        RECT 134.200 173.800 135.200 174.200 ;
        RECT 135.500 174.100 136.200 174.500 ;
        RECT 136.600 174.400 137.000 175.200 ;
        RECT 137.400 174.400 137.800 175.200 ;
        RECT 138.200 174.800 138.600 175.200 ;
        RECT 134.900 173.500 135.200 173.800 ;
        RECT 135.700 173.900 136.200 174.100 ;
        RECT 138.200 174.200 138.500 174.800 ;
        RECT 139.000 174.400 139.400 175.200 ;
        RECT 139.700 175.100 140.000 175.900 ;
        RECT 140.600 175.800 141.800 175.900 ;
        RECT 143.000 175.600 143.400 179.900 ;
        RECT 145.100 177.900 145.700 179.900 ;
        RECT 147.400 177.900 147.800 179.900 ;
        RECT 149.600 178.200 150.000 179.900 ;
        RECT 149.600 177.900 150.600 178.200 ;
        RECT 145.400 177.500 145.800 177.900 ;
        RECT 147.500 177.600 147.800 177.900 ;
        RECT 147.100 177.300 148.900 177.600 ;
        RECT 150.200 177.500 150.600 177.900 ;
        RECT 147.100 177.200 147.500 177.300 ;
        RECT 148.500 177.200 148.900 177.300 ;
        RECT 145.000 176.600 145.700 177.000 ;
        RECT 145.400 176.100 145.700 176.600 ;
        RECT 146.500 176.500 147.600 176.800 ;
        RECT 146.500 176.400 146.900 176.500 ;
        RECT 145.400 175.800 146.600 176.100 ;
        RECT 143.000 175.300 145.100 175.600 ;
        RECT 142.200 175.100 142.600 175.200 ;
        RECT 139.700 174.800 142.600 175.100 ;
        RECT 139.700 174.200 140.000 174.800 ;
        RECT 138.200 174.100 138.600 174.200 ;
        RECT 135.700 173.600 137.800 173.900 ;
        RECT 138.200 173.800 139.000 174.100 ;
        RECT 139.700 173.800 141.000 174.200 ;
        RECT 138.600 173.600 139.000 173.800 ;
        RECT 127.800 171.800 128.500 172.200 ;
        RECT 128.100 171.500 128.500 171.800 ;
        RECT 130.200 171.500 130.600 172.500 ;
        RECT 131.300 172.800 132.200 173.100 ;
        RECT 134.900 173.300 135.300 173.500 ;
        RECT 134.900 173.000 135.700 173.300 ;
        RECT 131.300 171.100 131.700 172.800 ;
        RECT 135.300 172.200 135.700 173.000 ;
        RECT 137.500 172.500 137.800 173.600 ;
        RECT 138.300 173.100 140.100 173.300 ;
        RECT 140.600 173.100 140.900 173.800 ;
        RECT 143.000 173.600 143.400 175.300 ;
        RECT 144.700 175.200 145.100 175.300 ;
        RECT 146.300 175.200 146.600 175.800 ;
        RECT 147.300 175.900 147.600 176.500 ;
        RECT 147.900 176.500 148.300 176.600 ;
        RECT 150.200 176.500 150.600 176.600 ;
        RECT 147.900 176.200 150.600 176.500 ;
        RECT 147.300 175.700 149.700 175.900 ;
        RECT 151.800 175.700 152.200 179.900 ;
        RECT 153.900 176.200 154.300 179.900 ;
        RECT 154.600 176.800 155.000 177.200 ;
        RECT 154.700 176.200 155.000 176.800 ;
        RECT 153.900 175.900 154.400 176.200 ;
        RECT 154.700 175.900 155.400 176.200 ;
        RECT 147.300 175.600 152.200 175.700 ;
        RECT 149.300 175.500 152.200 175.600 ;
        RECT 149.400 175.400 152.200 175.500 ;
        RECT 143.900 174.900 144.300 175.000 ;
        RECT 143.900 174.600 145.800 174.900 ;
        RECT 146.200 174.800 146.600 175.200 ;
        RECT 147.800 175.100 148.200 175.200 ;
        RECT 148.600 175.100 149.000 175.200 ;
        RECT 147.800 174.800 151.100 175.100 ;
        RECT 145.400 174.500 145.800 174.600 ;
        RECT 146.300 174.200 146.600 174.800 ;
        RECT 150.700 174.700 151.100 174.800 ;
        RECT 153.400 174.400 153.800 175.200 ;
        RECT 149.900 174.200 150.300 174.300 ;
        RECT 154.100 174.200 154.400 175.900 ;
        RECT 155.000 175.800 155.400 175.900 ;
        RECT 155.800 175.800 156.200 176.600 ;
        RECT 155.000 175.100 155.300 175.800 ;
        RECT 156.600 175.100 157.000 179.900 ;
        RECT 159.500 176.200 159.900 179.900 ;
        RECT 160.200 176.800 160.600 177.200 ;
        RECT 160.300 176.200 160.600 176.800 ;
        RECT 159.500 175.900 160.000 176.200 ;
        RECT 160.300 175.900 161.000 176.200 ;
        RECT 155.000 174.800 157.000 175.100 ;
        RECT 146.300 173.900 151.800 174.200 ;
        RECT 146.500 173.800 146.900 173.900 ;
        RECT 143.000 173.300 144.900 173.600 ;
        RECT 135.000 171.800 135.700 172.200 ;
        RECT 135.300 171.500 135.700 171.800 ;
        RECT 137.400 171.500 137.800 172.500 ;
        RECT 138.200 173.000 140.200 173.100 ;
        RECT 138.200 171.100 138.600 173.000 ;
        RECT 139.800 171.100 140.200 173.000 ;
        RECT 140.600 171.100 141.000 173.100 ;
        RECT 143.000 171.100 143.400 173.300 ;
        RECT 144.500 173.200 144.900 173.300 ;
        RECT 149.400 172.800 149.700 173.900 ;
        RECT 151.000 173.800 151.800 173.900 ;
        RECT 152.600 174.100 153.000 174.200 ;
        RECT 152.600 173.800 153.400 174.100 ;
        RECT 154.100 173.800 155.400 174.200 ;
        RECT 153.000 173.600 153.400 173.800 ;
        RECT 148.500 172.700 148.900 172.800 ;
        RECT 145.400 172.100 145.800 172.500 ;
        RECT 147.500 172.400 148.900 172.700 ;
        RECT 149.400 172.400 149.800 172.800 ;
        RECT 147.500 172.100 147.800 172.400 ;
        RECT 150.200 172.100 150.600 172.500 ;
        RECT 145.100 171.800 145.800 172.100 ;
        RECT 145.100 171.100 145.700 171.800 ;
        RECT 147.400 171.100 147.800 172.100 ;
        RECT 149.600 171.800 150.600 172.100 ;
        RECT 149.600 171.100 150.000 171.800 ;
        RECT 151.800 171.100 152.200 173.500 ;
        RECT 152.700 173.100 154.500 173.300 ;
        RECT 155.000 173.100 155.300 173.800 ;
        RECT 156.600 173.100 157.000 174.800 ;
        RECT 159.000 174.400 159.400 175.200 ;
        RECT 159.700 174.200 160.000 175.900 ;
        RECT 160.600 175.800 161.000 175.900 ;
        RECT 161.400 175.800 161.800 176.600 ;
        RECT 160.600 175.100 160.900 175.800 ;
        RECT 162.200 175.100 162.600 179.900 ;
        RECT 163.800 175.700 164.200 179.900 ;
        RECT 166.000 178.200 166.400 179.900 ;
        RECT 165.400 177.900 166.400 178.200 ;
        RECT 168.200 177.900 168.600 179.900 ;
        RECT 170.300 177.900 170.900 179.900 ;
        RECT 165.400 177.500 165.800 177.900 ;
        RECT 168.200 177.600 168.500 177.900 ;
        RECT 167.100 177.300 168.900 177.600 ;
        RECT 170.200 177.500 170.600 177.900 ;
        RECT 167.100 177.200 167.500 177.300 ;
        RECT 168.500 177.200 168.900 177.300 ;
        RECT 170.700 177.000 171.400 177.200 ;
        RECT 170.300 176.800 171.400 177.000 ;
        RECT 165.400 176.500 165.800 176.600 ;
        RECT 167.700 176.500 168.100 176.600 ;
        RECT 165.400 176.200 168.100 176.500 ;
        RECT 168.400 176.500 169.500 176.800 ;
        RECT 168.400 175.900 168.700 176.500 ;
        RECT 169.100 176.400 169.500 176.500 ;
        RECT 170.300 176.600 171.000 176.800 ;
        RECT 170.300 176.100 170.600 176.600 ;
        RECT 166.300 175.700 168.700 175.900 ;
        RECT 163.800 175.600 168.700 175.700 ;
        RECT 169.400 175.800 170.600 176.100 ;
        RECT 163.800 175.500 166.700 175.600 ;
        RECT 163.800 175.400 166.600 175.500 ;
        RECT 167.000 175.100 167.400 175.200 ;
        RECT 160.600 174.800 162.600 175.100 ;
        RECT 157.400 173.400 157.800 174.200 ;
        RECT 158.200 174.100 158.600 174.200 ;
        RECT 159.700 174.100 161.000 174.200 ;
        RECT 161.400 174.100 161.800 174.200 ;
        RECT 158.200 173.800 159.000 174.100 ;
        RECT 159.700 173.800 161.800 174.100 ;
        RECT 158.600 173.600 159.000 173.800 ;
        RECT 158.300 173.100 160.100 173.300 ;
        RECT 160.600 173.100 160.900 173.800 ;
        RECT 162.200 173.100 162.600 174.800 ;
        RECT 164.900 174.800 167.400 175.100 ;
        RECT 164.900 174.700 165.300 174.800 ;
        RECT 166.200 174.700 166.600 174.800 ;
        RECT 165.700 174.200 166.100 174.300 ;
        RECT 169.400 174.200 169.700 175.800 ;
        RECT 172.600 175.600 173.000 179.900 ;
        RECT 170.900 175.300 173.000 175.600 ;
        RECT 173.400 177.500 173.800 179.500 ;
        RECT 175.500 179.200 175.900 179.900 ;
        RECT 175.500 178.800 176.200 179.200 ;
        RECT 173.400 175.800 173.700 177.500 ;
        RECT 175.500 176.400 175.900 178.800 ;
        RECT 175.500 176.100 176.300 176.400 ;
        RECT 173.400 175.500 175.300 175.800 ;
        RECT 170.900 175.200 171.300 175.300 ;
        RECT 171.700 174.900 172.100 175.000 ;
        RECT 170.200 174.600 172.100 174.900 ;
        RECT 170.200 174.500 170.600 174.600 ;
        RECT 163.000 173.400 163.400 174.200 ;
        RECT 164.200 173.900 169.700 174.200 ;
        RECT 164.200 173.800 165.000 173.900 ;
        RECT 152.600 173.000 154.600 173.100 ;
        RECT 152.600 171.100 153.000 173.000 ;
        RECT 154.200 171.100 154.600 173.000 ;
        RECT 155.000 171.100 155.400 173.100 ;
        RECT 156.100 172.800 157.000 173.100 ;
        RECT 158.200 173.000 160.200 173.100 ;
        RECT 156.100 171.100 156.500 172.800 ;
        RECT 158.200 171.100 158.600 173.000 ;
        RECT 159.800 171.100 160.200 173.000 ;
        RECT 160.600 171.100 161.000 173.100 ;
        RECT 161.700 172.800 162.600 173.100 ;
        RECT 161.700 171.100 162.100 172.800 ;
        RECT 163.800 171.100 164.200 173.500 ;
        RECT 166.300 173.200 166.600 173.900 ;
        RECT 169.100 173.800 169.500 173.900 ;
        RECT 172.600 173.600 173.000 175.300 ;
        RECT 173.400 174.400 173.800 175.200 ;
        RECT 174.200 174.400 174.600 175.200 ;
        RECT 175.000 174.500 175.300 175.500 ;
        RECT 175.000 174.100 175.700 174.500 ;
        RECT 176.000 174.200 176.300 176.100 ;
        RECT 178.200 176.200 178.600 179.900 ;
        RECT 179.800 176.400 180.200 179.900 ;
        RECT 178.200 175.900 179.500 176.200 ;
        RECT 179.800 175.900 180.300 176.400 ;
        RECT 176.600 174.800 177.000 175.600 ;
        RECT 178.200 174.800 178.700 175.200 ;
        RECT 178.300 174.400 178.700 174.800 ;
        RECT 179.200 174.900 179.500 175.900 ;
        RECT 179.200 174.500 179.700 174.900 ;
        RECT 175.000 173.900 175.500 174.100 ;
        RECT 171.100 173.300 173.000 173.600 ;
        RECT 171.100 173.200 171.500 173.300 ;
        RECT 165.400 172.100 165.800 172.500 ;
        RECT 166.200 172.400 166.600 173.200 ;
        RECT 167.100 172.700 167.500 172.800 ;
        RECT 167.100 172.400 168.500 172.700 ;
        RECT 168.200 172.100 168.500 172.400 ;
        RECT 170.200 172.100 170.600 172.500 ;
        RECT 165.400 171.800 166.400 172.100 ;
        RECT 166.000 171.100 166.400 171.800 ;
        RECT 168.200 171.100 168.600 172.100 ;
        RECT 170.200 171.800 170.900 172.100 ;
        RECT 170.300 171.100 170.900 171.800 ;
        RECT 172.600 171.100 173.000 173.300 ;
        RECT 173.400 173.600 175.500 173.900 ;
        RECT 176.000 173.800 177.000 174.200 ;
        RECT 173.400 172.500 173.700 173.600 ;
        RECT 176.000 173.500 176.300 173.800 ;
        RECT 179.200 173.700 179.500 174.500 ;
        RECT 180.000 174.200 180.300 175.900 ;
        RECT 179.800 173.800 180.300 174.200 ;
        RECT 180.600 174.100 181.000 174.200 ;
        RECT 181.400 174.100 181.800 174.200 ;
        RECT 180.600 173.800 181.800 174.100 ;
        RECT 175.900 173.300 176.300 173.500 ;
        RECT 175.500 173.000 176.300 173.300 ;
        RECT 178.200 173.400 179.500 173.700 ;
        RECT 173.400 171.500 173.800 172.500 ;
        RECT 175.500 171.500 175.900 173.000 ;
        RECT 178.200 171.100 178.600 173.400 ;
        RECT 180.000 173.100 180.300 173.800 ;
        RECT 181.400 173.400 181.800 173.800 ;
        RECT 179.800 172.800 180.300 173.100 ;
        RECT 182.200 173.100 182.600 179.900 ;
        RECT 183.000 175.800 183.400 176.600 ;
        RECT 183.800 173.400 184.200 174.200 ;
        RECT 184.600 173.100 185.000 179.900 ;
        RECT 185.400 175.800 185.800 176.600 ;
        RECT 186.200 175.800 186.600 176.600 ;
        RECT 187.000 173.100 187.400 179.900 ;
        RECT 188.600 177.500 189.000 179.500 ;
        RECT 190.700 179.200 191.100 179.900 ;
        RECT 190.200 178.800 191.100 179.200 ;
        RECT 188.600 175.800 188.900 177.500 ;
        RECT 190.700 176.400 191.100 178.800 ;
        RECT 190.700 176.100 191.500 176.400 ;
        RECT 188.600 175.500 190.500 175.800 ;
        RECT 188.600 174.400 189.000 175.200 ;
        RECT 189.400 174.400 189.800 175.200 ;
        RECT 190.200 174.500 190.500 175.500 ;
        RECT 187.800 173.400 188.200 174.200 ;
        RECT 190.200 174.100 190.900 174.500 ;
        RECT 191.200 174.200 191.500 176.100 ;
        RECT 195.000 175.800 195.400 176.600 ;
        RECT 195.800 176.100 196.200 179.900 ;
        RECT 197.800 176.800 198.200 177.200 ;
        RECT 197.800 176.200 198.100 176.800 ;
        RECT 198.500 176.200 198.900 179.900 ;
        RECT 197.400 176.100 198.100 176.200 ;
        RECT 195.800 175.900 198.100 176.100 ;
        RECT 198.400 175.900 198.900 176.200 ;
        RECT 195.800 175.800 197.800 175.900 ;
        RECT 191.800 175.100 192.200 175.600 ;
        RECT 194.200 175.100 194.600 175.200 ;
        RECT 191.800 174.800 194.600 175.100 ;
        RECT 190.200 173.900 190.700 174.100 ;
        RECT 188.600 173.600 190.700 173.900 ;
        RECT 191.200 173.800 192.200 174.200 ;
        RECT 182.200 172.800 183.100 173.100 ;
        RECT 184.600 172.800 185.500 173.100 ;
        RECT 179.800 171.100 180.200 172.800 ;
        RECT 182.700 172.200 183.100 172.800 ;
        RECT 185.100 172.200 185.500 172.800 ;
        RECT 186.500 172.800 187.400 173.100 ;
        RECT 186.500 172.200 186.900 172.800 ;
        RECT 182.200 171.800 183.100 172.200 ;
        RECT 184.600 171.800 185.500 172.200 ;
        RECT 186.200 171.800 186.900 172.200 ;
        RECT 182.700 171.100 183.100 171.800 ;
        RECT 185.100 171.100 185.500 171.800 ;
        RECT 186.500 171.100 186.900 171.800 ;
        RECT 188.600 172.500 188.900 173.600 ;
        RECT 191.200 173.500 191.500 173.800 ;
        RECT 191.100 173.300 191.500 173.500 ;
        RECT 190.700 173.000 191.500 173.300 ;
        RECT 195.800 173.100 196.200 175.800 ;
        RECT 198.400 175.200 198.700 175.900 ;
        RECT 200.600 175.600 201.000 179.900 ;
        RECT 202.700 177.900 203.300 179.900 ;
        RECT 205.000 177.900 205.400 179.900 ;
        RECT 207.200 178.200 207.600 179.900 ;
        RECT 207.200 177.900 208.200 178.200 ;
        RECT 203.000 177.500 203.400 177.900 ;
        RECT 205.100 177.600 205.400 177.900 ;
        RECT 204.700 177.300 206.500 177.600 ;
        RECT 207.800 177.500 208.200 177.900 ;
        RECT 204.700 177.200 205.100 177.300 ;
        RECT 206.100 177.200 206.500 177.300 ;
        RECT 202.600 176.600 203.300 177.000 ;
        RECT 203.000 176.100 203.300 176.600 ;
        RECT 204.100 176.500 205.200 176.800 ;
        RECT 204.100 176.400 204.500 176.500 ;
        RECT 203.000 175.800 204.200 176.100 ;
        RECT 200.600 175.300 202.700 175.600 ;
        RECT 198.200 174.800 198.700 175.200 ;
        RECT 198.400 174.200 198.700 174.800 ;
        RECT 199.000 174.400 199.400 175.200 ;
        RECT 196.600 173.400 197.000 174.200 ;
        RECT 197.400 173.800 198.700 174.200 ;
        RECT 199.800 174.100 200.200 174.200 ;
        RECT 199.400 173.800 200.200 174.100 ;
        RECT 197.500 173.100 197.800 173.800 ;
        RECT 199.400 173.600 199.800 173.800 ;
        RECT 200.600 173.600 201.000 175.300 ;
        RECT 202.300 175.200 202.700 175.300 ;
        RECT 201.500 174.900 201.900 175.000 ;
        RECT 201.500 174.600 203.400 174.900 ;
        RECT 203.000 174.500 203.400 174.600 ;
        RECT 203.900 174.200 204.200 175.800 ;
        RECT 204.900 175.900 205.200 176.500 ;
        RECT 205.500 176.500 205.900 176.600 ;
        RECT 207.800 176.500 208.200 176.600 ;
        RECT 205.500 176.200 208.200 176.500 ;
        RECT 204.900 175.700 207.300 175.900 ;
        RECT 209.400 175.700 209.800 179.900 ;
        RECT 210.200 176.200 210.600 179.900 ;
        RECT 211.800 176.400 212.200 179.900 ;
        RECT 210.200 175.900 211.500 176.200 ;
        RECT 211.800 175.900 212.300 176.400 ;
        RECT 204.900 175.600 209.800 175.700 ;
        RECT 206.900 175.500 209.800 175.600 ;
        RECT 207.000 175.400 209.800 175.500 ;
        RECT 204.600 175.100 205.000 175.200 ;
        RECT 206.200 175.100 206.600 175.200 ;
        RECT 204.600 174.800 208.700 175.100 ;
        RECT 210.200 174.800 210.700 175.200 ;
        RECT 208.300 174.700 208.700 174.800 ;
        RECT 210.300 174.400 210.700 174.800 ;
        RECT 211.200 174.900 211.500 175.900 ;
        RECT 211.200 174.500 211.700 174.900 ;
        RECT 207.500 174.200 207.900 174.300 ;
        RECT 203.900 173.900 209.400 174.200 ;
        RECT 204.100 173.800 204.500 173.900 ;
        RECT 200.600 173.300 202.500 173.600 ;
        RECT 198.300 173.100 200.100 173.300 ;
        RECT 188.600 171.500 189.000 172.500 ;
        RECT 190.700 171.500 191.100 173.000 ;
        RECT 195.300 172.800 196.200 173.100 ;
        RECT 195.300 171.100 195.700 172.800 ;
        RECT 197.400 171.100 197.800 173.100 ;
        RECT 198.200 173.000 200.200 173.100 ;
        RECT 198.200 171.100 198.600 173.000 ;
        RECT 199.800 171.100 200.200 173.000 ;
        RECT 200.600 171.100 201.000 173.300 ;
        RECT 202.100 173.200 202.500 173.300 ;
        RECT 207.000 172.800 207.300 173.900 ;
        RECT 208.600 173.800 209.400 173.900 ;
        RECT 211.200 173.700 211.500 174.500 ;
        RECT 212.000 174.200 212.300 175.900 ;
        RECT 211.800 174.100 212.300 174.200 ;
        RECT 212.600 174.100 213.000 174.200 ;
        RECT 211.800 173.800 213.000 174.100 ;
        RECT 206.100 172.700 206.500 172.800 ;
        RECT 203.000 172.100 203.400 172.500 ;
        RECT 205.100 172.400 206.500 172.700 ;
        RECT 207.000 172.400 207.400 172.800 ;
        RECT 205.100 172.100 205.400 172.400 ;
        RECT 207.800 172.100 208.200 172.500 ;
        RECT 202.700 171.800 203.400 172.100 ;
        RECT 202.700 171.100 203.300 171.800 ;
        RECT 205.000 171.100 205.400 172.100 ;
        RECT 207.200 171.800 208.200 172.100 ;
        RECT 207.200 171.100 207.600 171.800 ;
        RECT 209.400 171.100 209.800 173.500 ;
        RECT 210.200 173.400 211.500 173.700 ;
        RECT 210.200 171.100 210.600 173.400 ;
        RECT 212.000 173.100 212.300 173.800 ;
        RECT 213.400 173.400 213.800 174.200 ;
        RECT 211.800 172.800 212.300 173.100 ;
        RECT 214.200 173.100 214.600 179.900 ;
        RECT 215.000 175.800 215.400 176.600 ;
        RECT 215.800 175.600 216.200 179.900 ;
        RECT 217.900 177.900 218.500 179.900 ;
        RECT 220.200 177.900 220.600 179.900 ;
        RECT 222.400 178.200 222.800 179.900 ;
        RECT 222.400 177.900 223.400 178.200 ;
        RECT 218.200 177.500 218.600 177.900 ;
        RECT 220.300 177.600 220.600 177.900 ;
        RECT 219.900 177.300 221.700 177.600 ;
        RECT 223.000 177.500 223.400 177.900 ;
        RECT 219.900 177.200 220.300 177.300 ;
        RECT 221.300 177.200 221.700 177.300 ;
        RECT 217.800 176.600 218.500 177.000 ;
        RECT 218.200 176.100 218.500 176.600 ;
        RECT 219.300 176.500 220.400 176.800 ;
        RECT 219.300 176.400 219.700 176.500 ;
        RECT 218.200 175.800 219.400 176.100 ;
        RECT 215.800 175.300 217.900 175.600 ;
        RECT 215.800 173.600 216.200 175.300 ;
        RECT 217.500 175.200 217.900 175.300 ;
        RECT 219.100 175.200 219.400 175.800 ;
        RECT 220.100 175.900 220.400 176.500 ;
        RECT 220.700 176.500 221.100 176.600 ;
        RECT 223.000 176.500 223.400 176.600 ;
        RECT 220.700 176.200 223.400 176.500 ;
        RECT 220.100 175.700 222.500 175.900 ;
        RECT 224.600 175.700 225.000 179.900 ;
        RECT 220.100 175.600 225.000 175.700 ;
        RECT 222.100 175.500 225.000 175.600 ;
        RECT 222.200 175.400 225.000 175.500 ;
        RECT 216.700 174.900 217.100 175.000 ;
        RECT 216.700 174.600 218.600 174.900 ;
        RECT 219.000 174.800 219.400 175.200 ;
        RECT 221.400 175.100 221.800 175.200 ;
        RECT 226.200 175.100 226.600 179.900 ;
        RECT 228.200 176.800 228.600 177.200 ;
        RECT 227.000 175.800 227.400 176.600 ;
        RECT 228.200 176.200 228.500 176.800 ;
        RECT 228.900 176.200 229.300 179.900 ;
        RECT 227.800 175.900 228.500 176.200 ;
        RECT 228.800 175.900 229.300 176.200 ;
        RECT 227.800 175.800 228.200 175.900 ;
        RECT 227.800 175.100 228.100 175.800 ;
        RECT 221.400 174.800 223.900 175.100 ;
        RECT 218.200 174.500 218.600 174.600 ;
        RECT 219.100 174.200 219.400 174.800 ;
        RECT 222.200 174.700 222.600 174.800 ;
        RECT 223.500 174.700 223.900 174.800 ;
        RECT 226.200 174.800 228.100 175.100 ;
        RECT 222.700 174.200 223.100 174.300 ;
        RECT 219.100 173.900 224.600 174.200 ;
        RECT 219.300 173.800 219.700 173.900 ;
        RECT 215.800 173.300 217.700 173.600 ;
        RECT 214.200 172.800 215.100 173.100 ;
        RECT 211.800 171.100 212.200 172.800 ;
        RECT 214.700 172.200 215.100 172.800 ;
        RECT 214.200 171.800 215.100 172.200 ;
        RECT 214.700 171.100 215.100 171.800 ;
        RECT 215.800 171.100 216.200 173.300 ;
        RECT 217.300 173.200 217.700 173.300 ;
        RECT 222.200 172.800 222.500 173.900 ;
        RECT 223.800 173.800 224.600 173.900 ;
        RECT 221.300 172.700 221.700 172.800 ;
        RECT 218.200 172.100 218.600 172.500 ;
        RECT 220.300 172.400 221.700 172.700 ;
        RECT 222.200 172.400 222.600 172.800 ;
        RECT 220.300 172.100 220.600 172.400 ;
        RECT 223.000 172.100 223.400 172.500 ;
        RECT 217.900 171.800 218.600 172.100 ;
        RECT 217.900 171.100 218.500 171.800 ;
        RECT 220.200 171.100 220.600 172.100 ;
        RECT 222.400 171.800 223.400 172.100 ;
        RECT 222.400 171.100 222.800 171.800 ;
        RECT 224.600 171.100 225.000 173.500 ;
        RECT 225.400 173.400 225.800 174.200 ;
        RECT 226.200 173.100 226.600 174.800 ;
        RECT 228.800 174.200 229.100 175.900 ;
        RECT 229.400 174.400 229.800 175.200 ;
        RECT 227.800 173.800 229.100 174.200 ;
        RECT 230.200 174.100 230.600 174.200 ;
        RECT 229.800 173.800 230.600 174.100 ;
        RECT 227.900 173.100 228.200 173.800 ;
        RECT 229.800 173.600 230.200 173.800 ;
        RECT 228.700 173.100 230.500 173.300 ;
        RECT 226.200 172.800 227.100 173.100 ;
        RECT 226.700 171.100 227.100 172.800 ;
        RECT 227.800 171.100 228.200 173.100 ;
        RECT 228.600 173.000 230.600 173.100 ;
        RECT 228.600 171.100 229.000 173.000 ;
        RECT 230.200 171.100 230.600 173.000 ;
        RECT 0.600 167.500 1.000 169.900 ;
        RECT 2.800 169.200 3.200 169.900 ;
        RECT 2.200 168.900 3.200 169.200 ;
        RECT 5.000 168.900 5.400 169.900 ;
        RECT 7.100 169.200 7.700 169.900 ;
        RECT 7.000 168.900 7.700 169.200 ;
        RECT 2.200 168.500 2.600 168.900 ;
        RECT 5.000 168.600 5.300 168.900 ;
        RECT 3.000 168.200 3.400 168.600 ;
        RECT 3.900 168.300 5.300 168.600 ;
        RECT 7.000 168.500 7.400 168.900 ;
        RECT 3.900 168.200 4.300 168.300 ;
        RECT 1.000 167.100 1.800 167.200 ;
        RECT 3.100 167.100 3.400 168.200 ;
        RECT 7.900 167.700 8.300 167.800 ;
        RECT 9.400 167.700 9.800 169.900 ;
        RECT 10.200 167.800 10.600 168.600 ;
        RECT 7.900 167.400 9.800 167.700 ;
        RECT 5.900 167.100 6.300 167.200 ;
        RECT 1.000 166.800 6.500 167.100 ;
        RECT 2.500 166.700 2.900 166.800 ;
        RECT 1.700 166.200 2.100 166.300 ;
        RECT 3.000 166.200 3.400 166.300 ;
        RECT 6.200 166.200 6.500 166.800 ;
        RECT 7.000 166.400 7.400 166.500 ;
        RECT 1.700 165.900 4.200 166.200 ;
        RECT 3.800 165.800 4.200 165.900 ;
        RECT 6.200 165.800 6.600 166.200 ;
        RECT 7.000 166.100 8.900 166.400 ;
        RECT 8.500 166.000 8.900 166.100 ;
        RECT 0.600 165.500 3.400 165.600 ;
        RECT 0.600 165.400 3.500 165.500 ;
        RECT 0.600 165.300 5.500 165.400 ;
        RECT 0.600 161.100 1.000 165.300 ;
        RECT 3.100 165.100 5.500 165.300 ;
        RECT 2.200 164.500 4.900 164.800 ;
        RECT 2.200 164.400 2.600 164.500 ;
        RECT 4.500 164.400 4.900 164.500 ;
        RECT 5.200 164.500 5.500 165.100 ;
        RECT 6.200 165.200 6.500 165.800 ;
        RECT 7.700 165.700 8.100 165.800 ;
        RECT 9.400 165.700 9.800 167.400 ;
        RECT 7.700 165.400 9.800 165.700 ;
        RECT 6.200 164.900 7.400 165.200 ;
        RECT 5.900 164.500 6.300 164.600 ;
        RECT 5.200 164.200 6.300 164.500 ;
        RECT 7.100 164.400 7.400 164.900 ;
        RECT 7.100 164.000 7.800 164.400 ;
        RECT 3.900 163.700 4.300 163.800 ;
        RECT 5.300 163.700 5.700 163.800 ;
        RECT 2.200 163.100 2.600 163.500 ;
        RECT 3.900 163.400 5.700 163.700 ;
        RECT 5.000 163.100 5.300 163.400 ;
        RECT 7.000 163.100 7.400 163.500 ;
        RECT 2.200 162.800 3.200 163.100 ;
        RECT 2.800 161.100 3.200 162.800 ;
        RECT 5.000 161.100 5.400 163.100 ;
        RECT 7.100 161.100 7.700 163.100 ;
        RECT 9.400 161.100 9.800 165.400 ;
        RECT 11.000 161.100 11.400 169.900 ;
        RECT 13.100 168.200 13.500 169.900 ;
        RECT 12.600 167.900 13.500 168.200 ;
        RECT 14.200 167.900 14.600 169.900 ;
        RECT 15.000 168.000 15.400 169.900 ;
        RECT 16.600 168.000 17.000 169.900 ;
        RECT 15.000 167.900 17.000 168.000 ;
        RECT 11.800 166.800 12.200 167.600 ;
        RECT 12.600 166.100 13.000 167.900 ;
        RECT 14.300 167.200 14.600 167.900 ;
        RECT 15.100 167.700 16.900 167.900 ;
        RECT 17.400 167.600 17.800 169.900 ;
        RECT 19.000 168.200 19.400 169.900 ;
        RECT 19.000 167.900 19.500 168.200 ;
        RECT 16.200 167.200 16.600 167.400 ;
        RECT 17.400 167.300 18.700 167.600 ;
        RECT 14.200 166.800 15.500 167.200 ;
        RECT 16.200 166.900 17.000 167.200 ;
        RECT 16.600 166.800 17.000 166.900 ;
        RECT 12.600 165.800 14.500 166.100 ;
        RECT 12.600 161.100 13.000 165.800 ;
        RECT 14.200 165.200 14.500 165.800 ;
        RECT 13.400 164.400 13.800 165.200 ;
        RECT 14.200 165.100 14.600 165.200 ;
        RECT 15.200 165.100 15.500 166.800 ;
        RECT 15.800 165.800 16.200 166.600 ;
        RECT 17.500 166.200 17.900 166.600 ;
        RECT 17.400 165.800 17.900 166.200 ;
        RECT 18.400 166.500 18.700 167.300 ;
        RECT 19.200 167.200 19.500 167.900 ;
        RECT 20.600 167.500 21.000 169.900 ;
        RECT 22.800 169.200 23.200 169.900 ;
        RECT 22.200 168.900 23.200 169.200 ;
        RECT 25.000 168.900 25.400 169.900 ;
        RECT 27.100 169.200 27.700 169.900 ;
        RECT 27.000 168.900 27.700 169.200 ;
        RECT 22.200 168.500 22.600 168.900 ;
        RECT 25.000 168.600 25.300 168.900 ;
        RECT 23.000 168.200 23.400 168.600 ;
        RECT 23.900 168.300 25.300 168.600 ;
        RECT 27.000 168.500 27.400 168.900 ;
        RECT 23.900 168.200 24.300 168.300 ;
        RECT 19.000 167.100 19.500 167.200 ;
        RECT 19.800 167.100 20.200 167.200 ;
        RECT 19.000 166.800 20.200 167.100 ;
        RECT 21.000 167.100 21.800 167.200 ;
        RECT 23.100 167.100 23.400 168.200 ;
        RECT 27.900 167.700 28.300 167.800 ;
        RECT 29.400 167.700 29.800 169.900 ;
        RECT 31.500 168.200 31.900 169.900 ;
        RECT 27.900 167.400 29.800 167.700 ;
        RECT 31.000 167.900 31.900 168.200 ;
        RECT 25.900 167.100 26.300 167.200 ;
        RECT 21.000 166.800 26.500 167.100 ;
        RECT 18.400 166.100 18.900 166.500 ;
        RECT 18.400 165.100 18.700 166.100 ;
        RECT 19.200 165.100 19.500 166.800 ;
        RECT 22.500 166.700 22.900 166.800 ;
        RECT 21.700 166.200 22.100 166.300 ;
        RECT 21.700 165.900 24.200 166.200 ;
        RECT 23.800 165.800 24.200 165.900 ;
        RECT 25.400 166.100 25.800 166.200 ;
        RECT 26.200 166.100 26.500 166.800 ;
        RECT 27.000 166.400 27.400 166.500 ;
        RECT 27.000 166.100 28.900 166.400 ;
        RECT 25.400 165.800 26.500 166.100 ;
        RECT 28.500 166.000 28.900 166.100 ;
        RECT 14.200 164.800 14.900 165.100 ;
        RECT 15.200 164.800 15.700 165.100 ;
        RECT 14.600 164.200 14.900 164.800 ;
        RECT 14.600 163.800 15.000 164.200 ;
        RECT 15.300 161.100 15.700 164.800 ;
        RECT 17.400 164.800 18.700 165.100 ;
        RECT 17.400 161.100 17.800 164.800 ;
        RECT 19.000 164.600 19.500 165.100 ;
        RECT 20.600 165.500 23.400 165.600 ;
        RECT 20.600 165.400 23.500 165.500 ;
        RECT 20.600 165.300 25.500 165.400 ;
        RECT 19.000 161.100 19.400 164.600 ;
        RECT 20.600 161.100 21.000 165.300 ;
        RECT 23.100 165.100 25.500 165.300 ;
        RECT 22.200 164.500 24.900 164.800 ;
        RECT 22.200 164.400 22.600 164.500 ;
        RECT 24.500 164.400 24.900 164.500 ;
        RECT 25.200 164.500 25.500 165.100 ;
        RECT 26.200 165.200 26.500 165.800 ;
        RECT 27.700 165.700 28.100 165.800 ;
        RECT 29.400 165.700 29.800 167.400 ;
        RECT 30.200 166.800 30.600 167.600 ;
        RECT 27.700 165.400 29.800 165.700 ;
        RECT 26.200 164.900 27.400 165.200 ;
        RECT 25.900 164.500 26.300 164.600 ;
        RECT 25.200 164.200 26.300 164.500 ;
        RECT 27.100 164.400 27.400 164.900 ;
        RECT 27.100 164.000 27.800 164.400 ;
        RECT 29.400 164.100 29.800 165.400 ;
        RECT 31.000 166.100 31.400 167.900 ;
        RECT 32.600 167.800 33.000 169.900 ;
        RECT 33.400 168.000 33.800 169.900 ;
        RECT 35.000 168.000 35.400 169.900 ;
        RECT 33.400 167.900 35.400 168.000 ;
        RECT 32.700 167.200 33.000 167.800 ;
        RECT 33.500 167.700 35.300 167.900 ;
        RECT 37.400 167.500 37.800 169.900 ;
        RECT 39.600 169.200 40.000 169.900 ;
        RECT 39.000 168.900 40.000 169.200 ;
        RECT 41.800 168.900 42.200 169.900 ;
        RECT 43.900 169.200 44.500 169.900 ;
        RECT 43.800 168.900 44.500 169.200 ;
        RECT 39.000 168.500 39.400 168.900 ;
        RECT 41.800 168.600 42.100 168.900 ;
        RECT 39.800 168.200 40.200 168.600 ;
        RECT 40.700 168.300 42.100 168.600 ;
        RECT 43.800 168.500 44.200 168.900 ;
        RECT 40.700 168.200 41.100 168.300 ;
        RECT 34.600 167.200 35.000 167.400 ;
        RECT 32.600 166.800 33.900 167.200 ;
        RECT 34.600 166.900 35.400 167.200 ;
        RECT 35.000 166.800 35.400 166.900 ;
        RECT 37.800 167.100 38.600 167.200 ;
        RECT 39.900 167.100 40.200 168.200 ;
        RECT 44.700 167.700 45.100 167.800 ;
        RECT 46.200 167.700 46.600 169.900 ;
        RECT 48.900 168.000 49.300 169.500 ;
        RECT 51.000 168.500 51.400 169.500 ;
        RECT 44.700 167.400 46.600 167.700 ;
        RECT 42.700 167.100 43.100 167.200 ;
        RECT 37.800 166.800 43.300 167.100 ;
        RECT 31.000 165.800 32.900 166.100 ;
        RECT 30.200 164.100 30.600 164.200 ;
        RECT 29.400 163.800 30.600 164.100 ;
        RECT 23.900 163.700 24.300 163.800 ;
        RECT 25.300 163.700 25.700 163.800 ;
        RECT 22.200 163.100 22.600 163.500 ;
        RECT 23.900 163.400 25.700 163.700 ;
        RECT 25.000 163.100 25.300 163.400 ;
        RECT 27.000 163.100 27.400 163.500 ;
        RECT 22.200 162.800 23.200 163.100 ;
        RECT 22.800 161.100 23.200 162.800 ;
        RECT 25.000 161.100 25.400 163.100 ;
        RECT 27.100 161.100 27.700 163.100 ;
        RECT 29.400 161.100 29.800 163.800 ;
        RECT 31.000 161.100 31.400 165.800 ;
        RECT 32.600 165.200 32.900 165.800 ;
        RECT 31.800 164.400 32.200 165.200 ;
        RECT 32.600 165.100 33.000 165.200 ;
        RECT 33.600 165.100 33.900 166.800 ;
        RECT 39.300 166.700 39.700 166.800 ;
        RECT 34.200 166.100 34.600 166.600 ;
        RECT 38.500 166.200 38.900 166.300 ;
        RECT 43.000 166.200 43.300 166.800 ;
        RECT 43.800 166.400 44.200 166.500 ;
        RECT 36.600 166.100 37.000 166.200 ;
        RECT 34.200 165.800 37.000 166.100 ;
        RECT 38.500 166.100 41.000 166.200 ;
        RECT 42.200 166.100 42.600 166.200 ;
        RECT 38.500 165.900 42.600 166.100 ;
        RECT 40.600 165.800 42.600 165.900 ;
        RECT 43.000 165.800 43.400 166.200 ;
        RECT 43.800 166.100 45.700 166.400 ;
        RECT 45.300 166.000 45.700 166.100 ;
        RECT 46.200 166.100 46.600 167.400 ;
        RECT 48.500 167.700 49.300 168.000 ;
        RECT 48.500 167.500 48.900 167.700 ;
        RECT 48.500 167.200 48.800 167.500 ;
        RECT 51.100 167.400 51.400 168.500 ;
        RECT 51.800 168.000 52.200 169.900 ;
        RECT 53.400 168.000 53.800 169.900 ;
        RECT 51.800 167.900 53.800 168.000 ;
        RECT 51.900 167.700 53.700 167.900 ;
        RECT 54.200 167.800 54.600 169.900 ;
        RECT 55.000 167.900 55.400 169.900 ;
        RECT 55.800 168.000 56.200 169.900 ;
        RECT 57.400 168.000 57.800 169.900 ;
        RECT 55.800 167.900 57.800 168.000 ;
        RECT 47.800 166.800 48.800 167.200 ;
        RECT 49.300 167.100 51.400 167.400 ;
        RECT 52.200 167.200 52.600 167.400 ;
        RECT 54.200 167.200 54.500 167.800 ;
        RECT 55.100 167.200 55.400 167.900 ;
        RECT 55.900 167.700 57.700 167.900 ;
        RECT 58.200 167.600 58.600 169.900 ;
        RECT 59.800 168.200 60.200 169.900 ;
        RECT 61.400 168.500 61.800 169.500 ;
        RECT 59.800 167.900 60.300 168.200 ;
        RECT 57.000 167.200 57.400 167.400 ;
        RECT 58.200 167.300 59.500 167.600 ;
        RECT 49.300 166.900 49.800 167.100 ;
        RECT 47.800 166.100 48.200 166.200 ;
        RECT 46.200 165.800 48.200 166.100 ;
        RECT 37.400 165.500 40.200 165.600 ;
        RECT 37.400 165.400 40.300 165.500 ;
        RECT 37.400 165.300 42.300 165.400 ;
        RECT 32.600 164.800 33.300 165.100 ;
        RECT 33.600 164.800 34.100 165.100 ;
        RECT 33.000 164.200 33.300 164.800 ;
        RECT 33.000 163.800 33.400 164.200 ;
        RECT 33.700 161.100 34.100 164.800 ;
        RECT 37.400 161.100 37.800 165.300 ;
        RECT 39.900 165.100 42.300 165.300 ;
        RECT 39.000 164.500 41.700 164.800 ;
        RECT 39.000 164.400 39.400 164.500 ;
        RECT 41.300 164.400 41.700 164.500 ;
        RECT 42.000 164.500 42.300 165.100 ;
        RECT 43.000 165.200 43.300 165.800 ;
        RECT 44.500 165.700 44.900 165.800 ;
        RECT 46.200 165.700 46.600 165.800 ;
        RECT 44.500 165.400 46.600 165.700 ;
        RECT 47.800 165.400 48.200 165.800 ;
        RECT 43.000 164.900 44.200 165.200 ;
        RECT 42.700 164.500 43.100 164.600 ;
        RECT 42.000 164.200 43.100 164.500 ;
        RECT 43.900 164.400 44.200 164.900 ;
        RECT 43.900 164.000 44.600 164.400 ;
        RECT 40.700 163.700 41.100 163.800 ;
        RECT 42.100 163.700 42.500 163.800 ;
        RECT 39.000 163.100 39.400 163.500 ;
        RECT 40.700 163.400 42.500 163.700 ;
        RECT 41.800 163.100 42.100 163.400 ;
        RECT 43.800 163.100 44.200 163.500 ;
        RECT 39.000 162.800 40.000 163.100 ;
        RECT 39.600 161.100 40.000 162.800 ;
        RECT 41.800 161.100 42.200 163.100 ;
        RECT 43.900 161.100 44.500 163.100 ;
        RECT 46.200 161.100 46.600 165.400 ;
        RECT 48.500 164.900 48.800 166.800 ;
        RECT 49.100 166.500 49.800 166.900 ;
        RECT 51.800 166.900 52.600 167.200 ;
        RECT 51.800 166.800 52.200 166.900 ;
        RECT 53.300 166.800 54.600 167.200 ;
        RECT 55.000 166.800 56.300 167.200 ;
        RECT 57.000 166.900 57.800 167.200 ;
        RECT 57.400 166.800 57.800 166.900 ;
        RECT 49.500 165.500 49.800 166.500 ;
        RECT 50.200 165.800 50.600 166.600 ;
        RECT 51.000 165.800 51.400 166.600 ;
        RECT 52.600 165.800 53.000 166.600 ;
        RECT 49.500 165.200 51.400 165.500 ;
        RECT 48.500 164.600 49.300 164.900 ;
        RECT 48.900 162.200 49.300 164.600 ;
        RECT 51.100 163.500 51.400 165.200 ;
        RECT 53.300 165.100 53.600 166.800 ;
        RECT 56.000 166.100 56.300 166.800 ;
        RECT 54.200 165.800 56.300 166.100 ;
        RECT 56.600 165.800 57.000 166.600 ;
        RECT 58.300 166.200 58.700 166.600 ;
        RECT 57.400 166.100 57.800 166.200 ;
        RECT 58.200 166.100 58.700 166.200 ;
        RECT 57.400 165.800 58.700 166.100 ;
        RECT 59.200 166.500 59.500 167.300 ;
        RECT 60.000 167.200 60.300 167.900 ;
        RECT 59.800 166.800 60.300 167.200 ;
        RECT 61.400 167.400 61.700 168.500 ;
        RECT 63.500 168.000 63.900 169.500 ;
        RECT 66.200 168.500 66.600 169.500 ;
        RECT 63.500 167.700 64.300 168.000 ;
        RECT 63.900 167.500 64.300 167.700 ;
        RECT 61.400 167.100 63.500 167.400 ;
        RECT 59.200 166.100 59.700 166.500 ;
        RECT 54.200 165.200 54.500 165.800 ;
        RECT 54.200 165.100 54.600 165.200 ;
        RECT 48.900 161.800 49.800 162.200 ;
        RECT 48.900 161.100 49.300 161.800 ;
        RECT 51.000 161.500 51.400 163.500 ;
        RECT 53.100 164.800 53.600 165.100 ;
        RECT 53.900 164.800 54.600 165.100 ;
        RECT 55.000 165.100 55.400 165.200 ;
        RECT 56.000 165.100 56.300 165.800 ;
        RECT 59.200 165.100 59.500 166.100 ;
        RECT 60.000 165.200 60.300 166.800 ;
        RECT 63.000 166.900 63.500 167.100 ;
        RECT 64.000 167.200 64.300 167.500 ;
        RECT 66.200 167.400 66.500 168.500 ;
        RECT 68.300 168.200 68.700 169.500 ;
        RECT 67.800 168.000 68.700 168.200 ;
        RECT 71.000 168.000 71.400 169.900 ;
        RECT 72.600 168.000 73.000 169.900 ;
        RECT 67.800 167.800 69.100 168.000 ;
        RECT 71.000 167.900 73.000 168.000 ;
        RECT 73.400 167.900 73.800 169.900 ;
        RECT 74.200 167.900 74.600 169.900 ;
        RECT 75.000 168.000 75.400 169.900 ;
        RECT 76.600 168.000 77.000 169.900 ;
        RECT 75.000 167.900 77.000 168.000 ;
        RECT 68.300 167.700 69.100 167.800 ;
        RECT 71.100 167.700 72.900 167.900 ;
        RECT 68.700 167.500 69.100 167.700 ;
        RECT 61.400 165.800 61.800 166.600 ;
        RECT 62.200 165.800 62.600 166.600 ;
        RECT 63.000 166.500 63.700 166.900 ;
        RECT 64.000 166.800 65.000 167.200 ;
        RECT 66.200 167.100 68.300 167.400 ;
        RECT 67.800 166.900 68.300 167.100 ;
        RECT 68.800 167.200 69.100 167.500 ;
        RECT 71.400 167.200 71.800 167.400 ;
        RECT 73.400 167.200 73.700 167.900 ;
        RECT 74.300 167.200 74.600 167.900 ;
        RECT 75.100 167.700 76.900 167.900 ;
        RECT 77.400 167.500 77.800 169.900 ;
        RECT 79.600 169.200 80.000 169.900 ;
        RECT 79.000 168.900 80.000 169.200 ;
        RECT 81.800 168.900 82.200 169.900 ;
        RECT 83.900 169.200 84.500 169.900 ;
        RECT 83.800 168.900 84.500 169.200 ;
        RECT 79.000 168.500 79.400 168.900 ;
        RECT 81.800 168.600 82.100 168.900 ;
        RECT 79.800 168.200 80.200 168.600 ;
        RECT 80.700 168.300 82.100 168.600 ;
        RECT 83.800 168.500 84.200 168.900 ;
        RECT 80.700 168.200 81.100 168.300 ;
        RECT 76.200 167.200 76.600 167.400 ;
        RECT 63.000 165.500 63.300 166.500 ;
        RECT 55.000 164.800 55.700 165.100 ;
        RECT 56.000 164.800 56.500 165.100 ;
        RECT 53.100 161.100 53.500 164.800 ;
        RECT 53.900 164.200 54.200 164.800 ;
        RECT 53.800 163.800 54.200 164.200 ;
        RECT 55.400 164.200 55.700 164.800 ;
        RECT 55.400 163.800 55.800 164.200 ;
        RECT 56.100 161.100 56.500 164.800 ;
        RECT 58.200 164.800 59.500 165.100 ;
        RECT 58.200 161.100 58.600 164.800 ;
        RECT 59.800 164.600 60.300 165.200 ;
        RECT 61.400 165.200 63.300 165.500 ;
        RECT 59.800 161.100 60.200 164.600 ;
        RECT 61.400 163.500 61.700 165.200 ;
        RECT 64.000 164.900 64.300 166.800 ;
        RECT 64.600 165.400 65.000 166.200 ;
        RECT 66.200 165.800 66.600 166.600 ;
        RECT 67.000 165.800 67.400 166.600 ;
        RECT 67.800 166.500 68.500 166.900 ;
        RECT 68.800 166.800 69.800 167.200 ;
        RECT 71.000 166.900 71.800 167.200 ;
        RECT 71.000 166.800 71.400 166.900 ;
        RECT 72.500 166.800 73.800 167.200 ;
        RECT 74.200 166.800 75.500 167.200 ;
        RECT 76.200 166.900 77.000 167.200 ;
        RECT 76.600 166.800 77.000 166.900 ;
        RECT 77.800 167.100 78.600 167.200 ;
        RECT 79.900 167.100 80.200 168.200 ;
        RECT 84.700 167.700 85.100 167.800 ;
        RECT 86.200 167.700 86.600 169.900 ;
        RECT 84.700 167.400 86.600 167.700 ;
        RECT 82.700 167.100 83.100 167.200 ;
        RECT 77.800 166.800 83.300 167.100 ;
        RECT 67.800 165.500 68.100 166.500 ;
        RECT 63.500 164.600 64.300 164.900 ;
        RECT 66.200 165.200 68.100 165.500 ;
        RECT 61.400 161.500 61.800 163.500 ;
        RECT 63.500 162.200 63.900 164.600 ;
        RECT 66.200 163.500 66.500 165.200 ;
        RECT 68.800 164.900 69.100 166.800 ;
        RECT 69.400 165.400 69.800 166.200 ;
        RECT 70.200 166.100 70.600 166.200 ;
        RECT 71.800 166.100 72.200 166.600 ;
        RECT 70.200 165.800 72.200 166.100 ;
        RECT 72.500 166.100 72.800 166.800 ;
        RECT 75.200 166.200 75.500 166.800 ;
        RECT 79.300 166.700 79.700 166.800 ;
        RECT 72.500 165.800 74.500 166.100 ;
        RECT 75.000 165.800 75.500 166.200 ;
        RECT 75.800 165.800 76.200 166.600 ;
        RECT 78.500 166.200 78.900 166.300 ;
        RECT 79.800 166.200 80.200 166.300 ;
        RECT 78.500 165.900 81.000 166.200 ;
        RECT 80.600 165.800 81.000 165.900 ;
        RECT 72.500 165.100 72.800 165.800 ;
        RECT 74.200 165.200 74.500 165.800 ;
        RECT 73.400 165.100 73.800 165.200 ;
        RECT 68.300 164.600 69.100 164.900 ;
        RECT 72.300 164.800 72.800 165.100 ;
        RECT 73.100 164.800 73.800 165.100 ;
        RECT 74.200 165.100 74.600 165.200 ;
        RECT 75.200 165.100 75.500 165.800 ;
        RECT 77.400 165.500 80.200 165.600 ;
        RECT 77.400 165.400 80.300 165.500 ;
        RECT 77.400 165.300 82.300 165.400 ;
        RECT 74.200 164.800 74.900 165.100 ;
        RECT 75.200 164.800 75.700 165.100 ;
        RECT 63.500 161.800 64.200 162.200 ;
        RECT 63.500 161.100 63.900 161.800 ;
        RECT 66.200 161.500 66.600 163.500 ;
        RECT 68.300 161.100 68.700 164.600 ;
        RECT 72.300 161.100 72.700 164.800 ;
        RECT 73.100 164.200 73.400 164.800 ;
        RECT 73.000 163.800 73.400 164.200 ;
        RECT 74.600 164.200 74.900 164.800 ;
        RECT 74.600 163.800 75.000 164.200 ;
        RECT 75.300 161.100 75.700 164.800 ;
        RECT 77.400 161.100 77.800 165.300 ;
        RECT 79.900 165.100 82.300 165.300 ;
        RECT 79.000 164.500 81.700 164.800 ;
        RECT 79.000 164.400 79.400 164.500 ;
        RECT 81.300 164.400 81.700 164.500 ;
        RECT 82.000 164.500 82.300 165.100 ;
        RECT 83.000 165.200 83.300 166.800 ;
        RECT 83.800 166.400 84.200 166.500 ;
        RECT 83.800 166.100 85.700 166.400 ;
        RECT 85.300 166.000 85.700 166.100 ;
        RECT 84.500 165.700 84.900 165.800 ;
        RECT 86.200 165.700 86.600 167.400 ;
        RECT 87.000 167.600 87.400 169.900 ;
        RECT 88.600 168.200 89.000 169.900 ;
        RECT 88.600 167.900 89.100 168.200 ;
        RECT 91.800 167.900 92.200 169.900 ;
        RECT 92.600 168.000 93.000 169.900 ;
        RECT 94.200 168.000 94.600 169.900 ;
        RECT 92.600 167.900 94.600 168.000 ;
        RECT 95.000 168.500 95.400 169.500 ;
        RECT 87.000 167.300 88.300 167.600 ;
        RECT 87.100 166.200 87.500 166.600 ;
        RECT 87.000 165.800 87.500 166.200 ;
        RECT 88.000 166.500 88.300 167.300 ;
        RECT 88.800 167.200 89.100 167.900 ;
        RECT 91.900 167.200 92.200 167.900 ;
        RECT 92.700 167.700 94.500 167.900 ;
        RECT 95.000 167.400 95.300 168.500 ;
        RECT 97.100 168.000 97.500 169.500 ;
        RECT 99.800 168.000 100.200 169.900 ;
        RECT 101.400 168.000 101.800 169.900 ;
        RECT 97.100 167.700 97.900 168.000 ;
        RECT 99.800 167.900 101.800 168.000 ;
        RECT 102.200 167.900 102.600 169.900 ;
        RECT 99.900 167.700 101.700 167.900 ;
        RECT 97.500 167.500 97.900 167.700 ;
        RECT 93.800 167.200 94.200 167.400 ;
        RECT 88.600 167.100 89.100 167.200 ;
        RECT 91.000 167.100 91.400 167.200 ;
        RECT 88.600 166.800 91.400 167.100 ;
        RECT 91.800 166.800 93.100 167.200 ;
        RECT 93.800 166.900 94.600 167.200 ;
        RECT 95.000 167.100 97.100 167.400 ;
        RECT 94.200 166.800 94.600 166.900 ;
        RECT 96.600 166.900 97.100 167.100 ;
        RECT 97.600 167.200 97.900 167.500 ;
        RECT 100.200 167.200 100.600 167.400 ;
        RECT 102.200 167.200 102.500 167.900 ;
        RECT 103.000 167.600 103.400 169.900 ;
        RECT 104.600 168.200 105.000 169.900 ;
        RECT 104.600 167.900 105.100 168.200 ;
        RECT 103.000 167.300 104.300 167.600 ;
        RECT 88.000 166.100 88.500 166.500 ;
        RECT 84.500 165.400 86.600 165.700 ;
        RECT 83.000 164.900 84.200 165.200 ;
        RECT 82.700 164.500 83.100 164.600 ;
        RECT 82.000 164.200 83.100 164.500 ;
        RECT 83.900 164.400 84.200 164.900 ;
        RECT 83.900 164.000 84.600 164.400 ;
        RECT 80.700 163.700 81.100 163.800 ;
        RECT 82.100 163.700 82.500 163.800 ;
        RECT 79.000 163.100 79.400 163.500 ;
        RECT 80.700 163.400 82.500 163.700 ;
        RECT 81.800 163.100 82.100 163.400 ;
        RECT 83.800 163.100 84.200 163.500 ;
        RECT 79.000 162.800 80.000 163.100 ;
        RECT 79.600 161.100 80.000 162.800 ;
        RECT 81.800 161.100 82.200 163.100 ;
        RECT 83.900 161.100 84.500 163.100 ;
        RECT 86.200 161.100 86.600 165.400 ;
        RECT 88.000 165.100 88.300 166.100 ;
        RECT 88.800 165.100 89.100 166.800 ;
        RECT 89.400 166.100 89.800 166.200 ;
        RECT 92.800 166.100 93.100 166.800 ;
        RECT 89.400 165.800 93.100 166.100 ;
        RECT 93.400 165.800 93.800 166.600 ;
        RECT 95.000 165.800 95.400 166.600 ;
        RECT 95.800 165.800 96.200 166.600 ;
        RECT 96.600 166.500 97.300 166.900 ;
        RECT 97.600 166.800 98.600 167.200 ;
        RECT 99.800 166.900 100.600 167.200 ;
        RECT 99.800 166.800 100.200 166.900 ;
        RECT 101.300 166.800 102.600 167.200 ;
        RECT 87.000 164.800 88.300 165.100 ;
        RECT 87.000 161.100 87.400 164.800 ;
        RECT 88.600 164.600 89.100 165.100 ;
        RECT 91.800 165.100 92.200 165.200 ;
        RECT 92.800 165.100 93.100 165.800 ;
        RECT 96.600 165.500 96.900 166.500 ;
        RECT 95.000 165.200 96.900 165.500 ;
        RECT 97.600 165.200 97.900 166.800 ;
        RECT 98.200 165.400 98.600 166.200 ;
        RECT 100.600 165.800 101.000 166.600 ;
        RECT 91.800 164.800 92.500 165.100 ;
        RECT 92.800 164.800 93.300 165.100 ;
        RECT 88.600 161.100 89.000 164.600 ;
        RECT 92.200 164.200 92.500 164.800 ;
        RECT 92.200 163.800 92.600 164.200 ;
        RECT 92.900 161.100 93.300 164.800 ;
        RECT 95.000 163.500 95.300 165.200 ;
        RECT 97.400 164.900 97.900 165.200 ;
        RECT 101.300 165.100 101.600 166.800 ;
        RECT 103.100 166.200 103.500 166.600 ;
        RECT 102.200 166.100 102.600 166.200 ;
        RECT 103.000 166.100 103.500 166.200 ;
        RECT 102.200 165.800 103.500 166.100 ;
        RECT 104.000 166.500 104.300 167.300 ;
        RECT 104.800 167.200 105.100 167.900 ;
        RECT 106.200 167.500 106.600 169.900 ;
        RECT 108.400 169.200 108.800 169.900 ;
        RECT 107.800 168.900 108.800 169.200 ;
        RECT 110.600 168.900 111.000 169.900 ;
        RECT 112.700 169.200 113.300 169.900 ;
        RECT 112.600 168.900 113.300 169.200 ;
        RECT 107.800 168.500 108.200 168.900 ;
        RECT 110.600 168.600 110.900 168.900 ;
        RECT 108.600 168.200 109.000 168.600 ;
        RECT 109.500 168.300 110.900 168.600 ;
        RECT 112.600 168.500 113.000 168.900 ;
        RECT 109.500 168.200 109.900 168.300 ;
        RECT 104.600 166.800 105.100 167.200 ;
        RECT 106.600 167.100 107.400 167.200 ;
        RECT 108.700 167.100 109.000 168.200 ;
        RECT 113.500 167.700 113.900 167.800 ;
        RECT 115.000 167.700 115.400 169.900 ;
        RECT 113.500 167.400 115.400 167.700 ;
        RECT 111.500 167.100 111.900 167.200 ;
        RECT 106.600 166.800 112.100 167.100 ;
        RECT 104.000 166.100 104.500 166.500 ;
        RECT 102.200 165.100 102.600 165.200 ;
        RECT 104.000 165.100 104.300 166.100 ;
        RECT 104.800 165.100 105.100 166.800 ;
        RECT 108.100 166.700 108.500 166.800 ;
        RECT 107.300 166.200 107.700 166.300 ;
        RECT 108.600 166.200 109.000 166.300 ;
        RECT 111.800 166.200 112.100 166.800 ;
        RECT 112.600 166.400 113.000 166.500 ;
        RECT 107.300 165.900 109.800 166.200 ;
        RECT 109.400 165.800 109.800 165.900 ;
        RECT 111.800 165.800 112.200 166.200 ;
        RECT 112.600 166.100 114.500 166.400 ;
        RECT 114.100 166.000 114.500 166.100 ;
        RECT 97.100 164.600 97.900 164.900 ;
        RECT 101.100 164.800 101.600 165.100 ;
        RECT 101.900 164.800 102.600 165.100 ;
        RECT 103.000 164.800 104.300 165.100 ;
        RECT 95.000 161.500 95.400 163.500 ;
        RECT 97.100 161.100 97.500 164.600 ;
        RECT 101.100 162.200 101.500 164.800 ;
        RECT 101.900 164.200 102.200 164.800 ;
        RECT 101.800 163.800 102.200 164.200 ;
        RECT 100.600 161.800 101.500 162.200 ;
        RECT 101.100 161.100 101.500 161.800 ;
        RECT 103.000 161.100 103.400 164.800 ;
        RECT 104.600 164.600 105.100 165.100 ;
        RECT 106.200 165.500 109.000 165.600 ;
        RECT 106.200 165.400 109.100 165.500 ;
        RECT 106.200 165.300 111.100 165.400 ;
        RECT 104.600 161.100 105.000 164.600 ;
        RECT 106.200 161.100 106.600 165.300 ;
        RECT 108.700 165.100 111.100 165.300 ;
        RECT 107.800 164.500 110.500 164.800 ;
        RECT 107.800 164.400 108.200 164.500 ;
        RECT 110.100 164.400 110.500 164.500 ;
        RECT 110.800 164.500 111.100 165.100 ;
        RECT 111.800 165.200 112.100 165.800 ;
        RECT 113.300 165.700 113.700 165.800 ;
        RECT 115.000 165.700 115.400 167.400 ;
        RECT 115.800 168.500 116.200 169.500 ;
        RECT 115.800 167.400 116.100 168.500 ;
        RECT 117.900 168.000 118.300 169.500 ;
        RECT 122.500 168.000 122.900 169.500 ;
        RECT 124.600 168.500 125.000 169.500 ;
        RECT 117.900 167.700 118.700 168.000 ;
        RECT 118.300 167.500 118.700 167.700 ;
        RECT 115.800 167.100 117.900 167.400 ;
        RECT 117.400 166.900 117.900 167.100 ;
        RECT 118.400 167.200 118.700 167.500 ;
        RECT 122.100 167.700 122.900 168.000 ;
        RECT 122.100 167.500 122.500 167.700 ;
        RECT 122.100 167.200 122.400 167.500 ;
        RECT 124.700 167.400 125.000 168.500 ;
        RECT 127.300 168.000 127.700 169.500 ;
        RECT 129.400 168.500 129.800 169.500 ;
        RECT 118.400 167.100 119.400 167.200 ;
        RECT 115.800 165.800 116.200 166.600 ;
        RECT 116.600 165.800 117.000 166.600 ;
        RECT 117.400 166.500 118.100 166.900 ;
        RECT 118.400 166.800 120.900 167.100 ;
        RECT 121.400 166.800 122.400 167.200 ;
        RECT 122.900 167.100 125.000 167.400 ;
        RECT 126.900 167.700 127.700 168.000 ;
        RECT 126.900 167.500 127.300 167.700 ;
        RECT 126.900 167.200 127.200 167.500 ;
        RECT 129.500 167.400 129.800 168.500 ;
        RECT 132.100 168.000 132.500 169.500 ;
        RECT 134.200 168.500 134.600 169.500 ;
        RECT 122.900 166.900 123.400 167.100 ;
        RECT 113.300 165.400 115.400 165.700 ;
        RECT 117.400 165.500 117.700 166.500 ;
        RECT 111.800 164.900 113.000 165.200 ;
        RECT 111.500 164.500 111.900 164.600 ;
        RECT 110.800 164.200 111.900 164.500 ;
        RECT 112.700 164.400 113.000 164.900 ;
        RECT 112.700 164.000 113.400 164.400 ;
        RECT 109.500 163.700 109.900 163.800 ;
        RECT 110.900 163.700 111.300 163.800 ;
        RECT 107.800 163.100 108.200 163.500 ;
        RECT 109.500 163.400 111.300 163.700 ;
        RECT 110.600 163.100 110.900 163.400 ;
        RECT 112.600 163.100 113.000 163.500 ;
        RECT 107.800 162.800 108.800 163.100 ;
        RECT 108.400 161.100 108.800 162.800 ;
        RECT 110.600 161.100 111.000 163.100 ;
        RECT 112.700 161.100 113.300 163.100 ;
        RECT 115.000 161.100 115.400 165.400 ;
        RECT 115.800 165.200 117.700 165.500 ;
        RECT 115.800 163.500 116.100 165.200 ;
        RECT 118.400 164.900 118.700 166.800 ;
        RECT 119.000 165.400 119.400 166.200 ;
        RECT 120.600 166.100 120.900 166.800 ;
        RECT 121.400 166.100 121.800 166.200 ;
        RECT 120.600 165.800 121.800 166.100 ;
        RECT 121.400 165.400 121.800 165.800 ;
        RECT 117.900 164.600 118.700 164.900 ;
        RECT 122.100 164.900 122.400 166.800 ;
        RECT 122.700 166.500 123.400 166.900 ;
        RECT 126.200 166.800 127.200 167.200 ;
        RECT 127.700 167.100 129.800 167.400 ;
        RECT 131.700 167.700 132.500 168.000 ;
        RECT 131.700 167.500 132.100 167.700 ;
        RECT 131.700 167.200 132.000 167.500 ;
        RECT 134.300 167.400 134.600 168.500 ;
        RECT 136.900 168.000 137.300 169.500 ;
        RECT 139.000 168.500 139.400 169.500 ;
        RECT 127.700 166.900 128.200 167.100 ;
        RECT 123.100 165.500 123.400 166.500 ;
        RECT 123.800 165.800 124.200 166.600 ;
        RECT 124.600 165.800 125.000 166.600 ;
        RECT 123.100 165.200 125.000 165.500 ;
        RECT 126.200 165.400 126.600 166.200 ;
        RECT 122.100 164.600 122.900 164.900 ;
        RECT 115.800 161.500 116.200 163.500 ;
        RECT 117.900 161.100 118.300 164.600 ;
        RECT 122.500 162.200 122.900 164.600 ;
        RECT 124.700 163.500 125.000 165.200 ;
        RECT 126.900 164.900 127.200 166.800 ;
        RECT 127.500 166.500 128.200 166.900 ;
        RECT 131.000 166.800 132.000 167.200 ;
        RECT 132.500 167.100 134.600 167.400 ;
        RECT 136.500 167.700 137.300 168.000 ;
        RECT 136.500 167.500 136.900 167.700 ;
        RECT 136.500 167.200 136.800 167.500 ;
        RECT 139.100 167.400 139.400 168.500 ;
        RECT 141.400 167.500 141.800 169.900 ;
        RECT 143.600 169.200 144.000 169.900 ;
        RECT 143.000 168.900 144.000 169.200 ;
        RECT 145.800 168.900 146.200 169.900 ;
        RECT 147.900 169.200 148.500 169.900 ;
        RECT 147.800 168.900 148.500 169.200 ;
        RECT 143.000 168.500 143.400 168.900 ;
        RECT 145.800 168.600 146.100 168.900 ;
        RECT 143.800 168.200 144.200 168.600 ;
        RECT 144.700 168.300 146.100 168.600 ;
        RECT 147.800 168.500 148.200 168.900 ;
        RECT 144.700 168.200 145.100 168.300 ;
        RECT 132.500 166.900 133.000 167.100 ;
        RECT 127.900 165.500 128.200 166.500 ;
        RECT 128.600 165.800 129.000 166.600 ;
        RECT 129.400 165.800 129.800 166.600 ;
        RECT 130.200 166.100 130.600 166.200 ;
        RECT 131.000 166.100 131.400 166.200 ;
        RECT 130.200 165.800 131.400 166.100 ;
        RECT 127.900 165.200 129.800 165.500 ;
        RECT 131.000 165.400 131.400 165.800 ;
        RECT 126.900 164.600 127.700 164.900 ;
        RECT 122.500 161.800 123.400 162.200 ;
        RECT 122.500 161.100 122.900 161.800 ;
        RECT 124.600 161.500 125.000 163.500 ;
        RECT 127.300 162.200 127.700 164.600 ;
        RECT 129.500 163.500 129.800 165.200 ;
        RECT 131.700 165.200 132.000 166.800 ;
        RECT 132.300 166.500 133.000 166.900 ;
        RECT 135.800 166.800 136.800 167.200 ;
        RECT 137.300 167.100 139.400 167.400 ;
        RECT 141.800 167.100 142.600 167.200 ;
        RECT 143.900 167.100 144.200 168.200 ;
        RECT 148.700 167.700 149.100 167.800 ;
        RECT 150.200 167.700 150.600 169.900 ;
        RECT 148.700 167.400 150.600 167.700 ;
        RECT 146.200 167.100 147.100 167.200 ;
        RECT 137.300 166.900 137.800 167.100 ;
        RECT 132.700 165.500 133.000 166.500 ;
        RECT 133.400 165.800 133.800 166.600 ;
        RECT 134.200 165.800 134.600 166.600 ;
        RECT 132.700 165.200 134.600 165.500 ;
        RECT 135.800 165.400 136.200 166.200 ;
        RECT 131.700 164.900 132.200 165.200 ;
        RECT 131.700 164.600 132.500 164.900 ;
        RECT 127.300 161.800 128.200 162.200 ;
        RECT 127.300 161.100 127.700 161.800 ;
        RECT 129.400 161.500 129.800 163.500 ;
        RECT 132.100 161.100 132.500 164.600 ;
        RECT 134.300 163.500 134.600 165.200 ;
        RECT 136.500 164.900 136.800 166.800 ;
        RECT 137.100 166.500 137.800 166.900 ;
        RECT 141.800 166.800 147.300 167.100 ;
        RECT 143.300 166.700 143.700 166.800 ;
        RECT 137.500 165.500 137.800 166.500 ;
        RECT 138.200 165.800 138.600 166.600 ;
        RECT 139.000 165.800 139.400 166.600 ;
        RECT 142.500 166.200 142.900 166.300 ;
        RECT 142.500 165.900 145.000 166.200 ;
        RECT 144.600 165.800 145.000 165.900 ;
        RECT 141.400 165.500 144.200 165.600 ;
        RECT 137.500 165.200 139.400 165.500 ;
        RECT 136.500 164.600 137.300 164.900 ;
        RECT 134.200 161.500 134.600 163.500 ;
        RECT 136.900 162.200 137.300 164.600 ;
        RECT 139.100 163.500 139.400 165.200 ;
        RECT 136.900 161.800 137.800 162.200 ;
        RECT 136.900 161.100 137.300 161.800 ;
        RECT 139.000 161.500 139.400 163.500 ;
        RECT 141.400 165.400 144.300 165.500 ;
        RECT 141.400 165.300 146.300 165.400 ;
        RECT 141.400 161.100 141.800 165.300 ;
        RECT 143.900 165.100 146.300 165.300 ;
        RECT 143.000 164.500 145.700 164.800 ;
        RECT 143.000 164.400 143.400 164.500 ;
        RECT 145.300 164.400 145.700 164.500 ;
        RECT 146.000 164.500 146.300 165.100 ;
        RECT 147.000 165.200 147.300 166.800 ;
        RECT 147.800 166.400 148.200 166.500 ;
        RECT 147.800 166.100 149.700 166.400 ;
        RECT 149.300 166.000 149.700 166.100 ;
        RECT 148.500 165.700 148.900 165.800 ;
        RECT 150.200 165.700 150.600 167.400 ;
        RECT 148.500 165.400 150.600 165.700 ;
        RECT 147.000 164.900 148.200 165.200 ;
        RECT 146.700 164.500 147.100 164.600 ;
        RECT 146.000 164.200 147.100 164.500 ;
        RECT 147.900 164.400 148.200 164.900 ;
        RECT 147.900 164.000 148.600 164.400 ;
        RECT 144.700 163.700 145.100 163.800 ;
        RECT 146.100 163.700 146.500 163.800 ;
        RECT 143.000 163.100 143.400 163.500 ;
        RECT 144.700 163.400 146.500 163.700 ;
        RECT 145.800 163.100 146.100 163.400 ;
        RECT 147.800 163.100 148.200 163.500 ;
        RECT 143.000 162.800 144.000 163.100 ;
        RECT 143.600 161.100 144.000 162.800 ;
        RECT 145.800 161.100 146.200 163.100 ;
        RECT 147.900 161.100 148.500 163.100 ;
        RECT 150.200 161.100 150.600 165.400 ;
        RECT 151.000 161.100 151.400 169.900 ;
        RECT 151.800 167.800 152.200 168.600 ;
        RECT 152.600 167.900 153.000 169.900 ;
        RECT 153.400 168.000 153.800 169.900 ;
        RECT 155.000 168.000 155.400 169.900 ;
        RECT 157.100 168.200 157.500 169.900 ;
        RECT 153.400 167.900 155.400 168.000 ;
        RECT 156.600 167.900 157.500 168.200 ;
        RECT 152.700 167.200 153.000 167.900 ;
        RECT 153.500 167.700 155.300 167.900 ;
        RECT 154.600 167.200 155.000 167.400 ;
        RECT 152.600 166.800 153.900 167.200 ;
        RECT 154.600 166.900 155.400 167.200 ;
        RECT 155.000 166.800 155.400 166.900 ;
        RECT 155.800 166.800 156.200 167.600 ;
        RECT 153.600 166.200 153.900 166.800 ;
        RECT 153.400 165.800 153.900 166.200 ;
        RECT 154.200 165.800 154.600 166.600 ;
        RECT 155.800 166.100 156.200 166.200 ;
        RECT 156.600 166.100 157.000 167.900 ;
        RECT 158.200 167.500 158.600 169.900 ;
        RECT 160.400 169.200 160.800 169.900 ;
        RECT 159.800 168.900 160.800 169.200 ;
        RECT 162.600 168.900 163.000 169.900 ;
        RECT 164.700 169.200 165.300 169.900 ;
        RECT 164.600 168.900 165.300 169.200 ;
        RECT 159.800 168.500 160.200 168.900 ;
        RECT 162.600 168.600 162.900 168.900 ;
        RECT 160.600 168.200 161.000 168.600 ;
        RECT 161.500 168.300 162.900 168.600 ;
        RECT 164.600 168.500 165.000 168.900 ;
        RECT 161.500 168.200 161.900 168.300 ;
        RECT 158.600 167.100 159.400 167.200 ;
        RECT 160.700 167.100 161.000 168.200 ;
        RECT 165.500 167.700 165.900 167.800 ;
        RECT 167.000 167.700 167.400 169.900 ;
        RECT 169.100 168.200 169.500 169.900 ;
        RECT 165.500 167.400 167.400 167.700 ;
        RECT 168.600 167.900 169.500 168.200 ;
        RECT 170.200 167.900 170.600 169.900 ;
        RECT 171.000 168.000 171.400 169.900 ;
        RECT 172.600 168.000 173.000 169.900 ;
        RECT 171.000 167.900 173.000 168.000 ;
        RECT 163.500 167.100 163.900 167.200 ;
        RECT 158.600 166.800 164.100 167.100 ;
        RECT 160.100 166.700 160.500 166.800 ;
        RECT 155.800 165.800 157.000 166.100 ;
        RECT 159.300 166.200 159.700 166.300 ;
        RECT 159.300 165.900 161.800 166.200 ;
        RECT 161.400 165.800 161.800 165.900 ;
        RECT 152.600 165.100 153.000 165.200 ;
        RECT 153.600 165.100 153.900 165.800 ;
        RECT 152.600 164.800 153.300 165.100 ;
        RECT 153.600 164.800 154.100 165.100 ;
        RECT 153.000 164.200 153.300 164.800 ;
        RECT 153.000 163.800 153.400 164.200 ;
        RECT 153.700 161.100 154.100 164.800 ;
        RECT 156.600 161.100 157.000 165.800 ;
        RECT 158.200 165.500 161.000 165.600 ;
        RECT 158.200 165.400 161.100 165.500 ;
        RECT 158.200 165.300 163.100 165.400 ;
        RECT 157.400 164.400 157.800 165.200 ;
        RECT 158.200 161.100 158.600 165.300 ;
        RECT 160.700 165.100 163.100 165.300 ;
        RECT 159.800 164.500 162.500 164.800 ;
        RECT 159.800 164.400 160.200 164.500 ;
        RECT 162.100 164.400 162.500 164.500 ;
        RECT 162.800 164.500 163.100 165.100 ;
        RECT 163.800 165.200 164.100 166.800 ;
        RECT 164.600 166.400 165.000 166.500 ;
        RECT 164.600 166.100 166.500 166.400 ;
        RECT 166.100 166.000 166.500 166.100 ;
        RECT 165.300 165.700 165.700 165.800 ;
        RECT 167.000 165.700 167.400 167.400 ;
        RECT 167.800 166.800 168.200 167.600 ;
        RECT 165.300 165.400 167.400 165.700 ;
        RECT 163.800 164.900 165.000 165.200 ;
        RECT 163.500 164.500 163.900 164.600 ;
        RECT 162.800 164.200 163.900 164.500 ;
        RECT 164.700 164.400 165.000 164.900 ;
        RECT 164.700 164.000 165.400 164.400 ;
        RECT 167.000 164.100 167.400 165.400 ;
        RECT 168.600 166.100 169.000 167.900 ;
        RECT 170.300 167.200 170.600 167.900 ;
        RECT 171.100 167.700 172.900 167.900 ;
        RECT 172.200 167.200 172.600 167.400 ;
        RECT 169.400 167.100 169.800 167.200 ;
        RECT 170.200 167.100 171.500 167.200 ;
        RECT 169.400 166.800 171.500 167.100 ;
        RECT 172.200 166.900 173.000 167.200 ;
        RECT 174.000 167.100 174.400 169.900 ;
        RECT 177.900 168.200 178.300 169.900 ;
        RECT 177.400 167.900 178.300 168.200 ;
        RECT 172.600 166.800 173.000 166.900 ;
        RECT 173.500 166.900 174.400 167.100 ;
        RECT 173.500 166.800 174.300 166.900 ;
        RECT 176.600 166.800 177.000 167.600 ;
        RECT 168.600 165.800 170.500 166.100 ;
        RECT 167.800 164.100 168.200 164.200 ;
        RECT 167.000 163.800 168.200 164.100 ;
        RECT 161.500 163.700 161.900 163.800 ;
        RECT 162.900 163.700 163.300 163.800 ;
        RECT 159.800 163.100 160.200 163.500 ;
        RECT 161.500 163.400 163.300 163.700 ;
        RECT 162.600 163.100 162.900 163.400 ;
        RECT 164.600 163.100 165.000 163.500 ;
        RECT 159.800 162.800 160.800 163.100 ;
        RECT 160.400 161.100 160.800 162.800 ;
        RECT 162.600 161.100 163.000 163.100 ;
        RECT 164.700 161.100 165.300 163.100 ;
        RECT 167.000 161.100 167.400 163.800 ;
        RECT 168.600 161.100 169.000 165.800 ;
        RECT 170.200 165.200 170.500 165.800 ;
        RECT 169.400 164.400 169.800 165.200 ;
        RECT 170.200 165.100 170.600 165.200 ;
        RECT 171.200 165.100 171.500 166.800 ;
        RECT 171.800 165.800 172.200 166.600 ;
        RECT 173.500 165.200 173.800 166.800 ;
        RECT 174.600 165.800 175.400 166.200 ;
        RECT 170.200 164.800 170.900 165.100 ;
        RECT 171.200 164.800 171.700 165.100 ;
        RECT 173.400 164.800 173.800 165.200 ;
        RECT 175.800 164.800 176.200 165.600 ;
        RECT 170.600 164.200 170.900 164.800 ;
        RECT 170.600 163.800 171.000 164.200 ;
        RECT 171.300 161.100 171.700 164.800 ;
        RECT 173.500 163.500 173.800 164.800 ;
        RECT 174.200 163.800 174.600 164.600 ;
        RECT 173.500 163.200 175.300 163.500 ;
        RECT 173.500 163.100 173.800 163.200 ;
        RECT 173.400 161.100 173.800 163.100 ;
        RECT 175.000 163.100 175.300 163.200 ;
        RECT 175.000 161.100 175.400 163.100 ;
        RECT 177.400 161.100 177.800 167.900 ;
        RECT 179.000 167.600 179.400 169.900 ;
        RECT 180.600 168.200 181.000 169.900 ;
        RECT 180.600 167.900 181.100 168.200 ;
        RECT 182.200 168.000 182.600 169.900 ;
        RECT 183.800 168.000 184.200 169.900 ;
        RECT 182.200 167.900 184.200 168.000 ;
        RECT 184.600 167.900 185.000 169.900 ;
        RECT 179.000 167.300 180.300 167.600 ;
        RECT 179.100 166.200 179.500 166.600 ;
        RECT 178.200 166.100 178.600 166.200 ;
        RECT 179.000 166.100 179.500 166.200 ;
        RECT 178.200 165.800 179.500 166.100 ;
        RECT 180.000 166.500 180.300 167.300 ;
        RECT 180.800 167.200 181.100 167.900 ;
        RECT 182.300 167.700 184.100 167.900 ;
        RECT 182.600 167.200 183.000 167.400 ;
        RECT 184.600 167.200 184.900 167.900 ;
        RECT 185.400 167.500 185.800 169.900 ;
        RECT 187.600 169.200 188.000 169.900 ;
        RECT 187.000 168.900 188.000 169.200 ;
        RECT 189.800 168.900 190.200 169.900 ;
        RECT 191.900 169.200 192.500 169.900 ;
        RECT 191.800 168.900 192.500 169.200 ;
        RECT 187.000 168.500 187.400 168.900 ;
        RECT 189.800 168.600 190.100 168.900 ;
        RECT 187.800 168.200 188.200 168.600 ;
        RECT 188.700 168.300 190.100 168.600 ;
        RECT 191.800 168.500 192.200 168.900 ;
        RECT 188.700 168.200 189.100 168.300 ;
        RECT 180.600 166.800 181.100 167.200 ;
        RECT 182.200 166.900 183.000 167.200 ;
        RECT 182.200 166.800 182.600 166.900 ;
        RECT 183.700 166.800 185.000 167.200 ;
        RECT 185.800 167.100 186.600 167.200 ;
        RECT 187.900 167.100 188.200 168.200 ;
        RECT 192.700 167.700 193.100 167.800 ;
        RECT 194.200 167.700 194.600 169.900 ;
        RECT 192.700 167.400 194.600 167.700 ;
        RECT 189.400 167.100 189.800 167.200 ;
        RECT 190.700 167.100 191.100 167.200 ;
        RECT 185.800 166.800 191.300 167.100 ;
        RECT 180.000 166.100 180.500 166.500 ;
        RECT 178.200 164.400 178.600 165.200 ;
        RECT 180.000 165.100 180.300 166.100 ;
        RECT 180.800 165.100 181.100 166.800 ;
        RECT 183.000 165.800 183.400 166.600 ;
        RECT 183.700 165.100 184.000 166.800 ;
        RECT 187.300 166.700 187.700 166.800 ;
        RECT 186.500 166.200 186.900 166.300 ;
        RECT 187.800 166.200 188.200 166.300 ;
        RECT 186.500 165.900 189.000 166.200 ;
        RECT 188.600 165.800 189.000 165.900 ;
        RECT 185.400 165.500 188.200 165.600 ;
        RECT 185.400 165.400 188.300 165.500 ;
        RECT 185.400 165.300 190.300 165.400 ;
        RECT 184.600 165.100 185.000 165.200 ;
        RECT 179.000 164.800 180.300 165.100 ;
        RECT 179.000 161.100 179.400 164.800 ;
        RECT 180.600 164.600 181.100 165.100 ;
        RECT 183.500 164.800 184.000 165.100 ;
        RECT 184.300 164.800 185.000 165.100 ;
        RECT 180.600 161.100 181.000 164.600 ;
        RECT 183.500 161.100 183.900 164.800 ;
        RECT 184.300 164.200 184.600 164.800 ;
        RECT 184.200 163.800 184.600 164.200 ;
        RECT 185.400 161.100 185.800 165.300 ;
        RECT 187.900 165.100 190.300 165.300 ;
        RECT 187.000 164.500 189.700 164.800 ;
        RECT 187.000 164.400 187.400 164.500 ;
        RECT 189.300 164.400 189.700 164.500 ;
        RECT 190.000 164.500 190.300 165.100 ;
        RECT 191.000 165.200 191.300 166.800 ;
        RECT 191.800 166.400 192.200 166.500 ;
        RECT 191.800 166.100 193.700 166.400 ;
        RECT 193.300 166.000 193.700 166.100 ;
        RECT 192.500 165.700 192.900 165.800 ;
        RECT 194.200 165.700 194.600 167.400 ;
        RECT 196.600 168.500 197.000 169.500 ;
        RECT 196.600 167.400 196.900 168.500 ;
        RECT 198.700 168.000 199.100 169.500 ;
        RECT 201.400 168.500 201.800 169.500 ;
        RECT 198.700 167.700 199.500 168.000 ;
        RECT 199.100 167.500 199.500 167.700 ;
        RECT 196.600 167.100 198.700 167.400 ;
        RECT 198.200 166.900 198.700 167.100 ;
        RECT 199.200 167.200 199.500 167.500 ;
        RECT 201.400 167.400 201.700 168.500 ;
        RECT 203.500 168.200 203.900 169.500 ;
        RECT 203.000 168.000 203.900 168.200 ;
        RECT 203.000 167.800 204.300 168.000 ;
        RECT 203.500 167.700 204.300 167.800 ;
        RECT 203.900 167.500 204.300 167.700 ;
        RECT 196.600 165.800 197.000 166.600 ;
        RECT 197.400 165.800 197.800 166.600 ;
        RECT 198.200 166.500 198.900 166.900 ;
        RECT 199.200 166.800 200.200 167.200 ;
        RECT 201.400 167.100 203.500 167.400 ;
        RECT 203.000 166.900 203.500 167.100 ;
        RECT 204.000 167.200 204.300 167.500 ;
        RECT 206.200 167.700 206.600 169.900 ;
        RECT 208.300 169.200 208.900 169.900 ;
        RECT 208.300 168.900 209.000 169.200 ;
        RECT 210.600 168.900 211.000 169.900 ;
        RECT 212.800 169.200 213.200 169.900 ;
        RECT 212.800 168.900 213.800 169.200 ;
        RECT 208.600 168.500 209.000 168.900 ;
        RECT 210.700 168.600 211.000 168.900 ;
        RECT 210.700 168.300 212.100 168.600 ;
        RECT 211.700 168.200 212.100 168.300 ;
        RECT 212.600 168.200 213.000 168.600 ;
        RECT 213.400 168.500 213.800 168.900 ;
        RECT 207.700 167.700 208.100 167.800 ;
        RECT 206.200 167.400 208.200 167.700 ;
        RECT 192.500 165.400 194.600 165.700 ;
        RECT 198.200 165.500 198.500 166.500 ;
        RECT 191.000 164.900 192.200 165.200 ;
        RECT 190.700 164.500 191.100 164.600 ;
        RECT 190.000 164.200 191.100 164.500 ;
        RECT 191.900 164.400 192.200 164.900 ;
        RECT 191.900 164.000 192.600 164.400 ;
        RECT 188.700 163.700 189.100 163.800 ;
        RECT 190.100 163.700 190.500 163.800 ;
        RECT 187.000 163.100 187.400 163.500 ;
        RECT 188.700 163.400 190.500 163.700 ;
        RECT 189.800 163.100 190.100 163.400 ;
        RECT 191.800 163.100 192.200 163.500 ;
        RECT 187.000 162.800 188.000 163.100 ;
        RECT 187.600 161.100 188.000 162.800 ;
        RECT 189.800 161.100 190.200 163.100 ;
        RECT 191.900 161.100 192.500 163.100 ;
        RECT 194.200 161.100 194.600 165.400 ;
        RECT 196.600 165.200 198.500 165.500 ;
        RECT 199.200 165.200 199.500 166.800 ;
        RECT 199.800 165.400 200.200 166.200 ;
        RECT 201.400 165.800 201.800 166.600 ;
        RECT 202.200 165.800 202.600 166.600 ;
        RECT 203.000 166.500 203.700 166.900 ;
        RECT 204.000 166.800 205.000 167.200 ;
        RECT 203.000 165.500 203.300 166.500 ;
        RECT 196.600 163.500 196.900 165.200 ;
        RECT 199.000 164.900 199.500 165.200 ;
        RECT 198.700 164.600 199.500 164.900 ;
        RECT 201.400 165.200 203.300 165.500 ;
        RECT 196.600 161.500 197.000 163.500 ;
        RECT 198.700 161.100 199.100 164.600 ;
        RECT 201.400 163.500 201.700 165.200 ;
        RECT 204.000 164.900 204.300 166.800 ;
        RECT 204.600 166.100 205.000 166.200 ;
        RECT 206.200 166.100 206.600 167.400 ;
        RECT 207.800 166.800 208.200 167.400 ;
        RECT 209.700 167.100 210.100 167.200 ;
        RECT 211.000 167.100 211.400 167.200 ;
        RECT 212.600 167.100 212.900 168.200 ;
        RECT 215.000 167.500 215.400 169.900 ;
        RECT 217.100 168.200 217.500 169.900 ;
        RECT 216.600 167.900 217.500 168.200 ;
        RECT 218.200 167.900 218.600 169.900 ;
        RECT 219.000 168.000 219.400 169.900 ;
        RECT 220.600 168.000 221.000 169.900 ;
        RECT 222.700 168.200 223.100 169.900 ;
        RECT 219.000 167.900 221.000 168.000 ;
        RECT 222.200 167.900 223.100 168.200 ;
        RECT 214.200 167.100 215.000 167.200 ;
        RECT 209.500 166.800 215.000 167.100 ;
        RECT 215.800 166.800 216.200 167.600 ;
        RECT 208.600 166.400 209.000 166.500 ;
        RECT 204.600 165.800 206.600 166.100 ;
        RECT 207.100 166.100 209.000 166.400 ;
        RECT 207.100 166.000 207.500 166.100 ;
        RECT 204.600 165.400 205.000 165.800 ;
        RECT 206.200 165.700 206.600 165.800 ;
        RECT 207.900 165.700 208.300 165.800 ;
        RECT 206.200 165.400 208.300 165.700 ;
        RECT 203.500 164.600 204.300 164.900 ;
        RECT 201.400 161.500 201.800 163.500 ;
        RECT 203.500 161.100 203.900 164.600 ;
        RECT 206.200 161.100 206.600 165.400 ;
        RECT 209.500 165.200 209.800 166.800 ;
        RECT 213.100 166.700 213.500 166.800 ;
        RECT 212.600 166.200 213.000 166.300 ;
        RECT 213.900 166.200 214.300 166.300 ;
        RECT 211.800 165.900 214.300 166.200 ;
        RECT 216.600 166.100 217.000 167.900 ;
        RECT 218.300 167.200 218.600 167.900 ;
        RECT 219.100 167.700 220.900 167.900 ;
        RECT 220.200 167.200 220.600 167.400 ;
        RECT 218.200 166.800 219.500 167.200 ;
        RECT 220.200 166.900 221.000 167.200 ;
        RECT 220.600 166.800 221.000 166.900 ;
        RECT 221.400 166.800 221.800 167.600 ;
        RECT 211.800 165.800 212.200 165.900 ;
        RECT 216.600 165.800 218.500 166.100 ;
        RECT 212.600 165.500 215.400 165.600 ;
        RECT 212.500 165.400 215.400 165.500 ;
        RECT 208.600 164.900 209.800 165.200 ;
        RECT 210.500 165.300 215.400 165.400 ;
        RECT 210.500 165.100 212.900 165.300 ;
        RECT 208.600 164.400 208.900 164.900 ;
        RECT 208.200 164.000 208.900 164.400 ;
        RECT 209.700 164.500 210.100 164.600 ;
        RECT 210.500 164.500 210.800 165.100 ;
        RECT 209.700 164.200 210.800 164.500 ;
        RECT 211.100 164.500 213.800 164.800 ;
        RECT 211.100 164.400 211.500 164.500 ;
        RECT 213.400 164.400 213.800 164.500 ;
        RECT 210.300 163.700 210.700 163.800 ;
        RECT 211.700 163.700 212.100 163.800 ;
        RECT 208.600 163.100 209.000 163.500 ;
        RECT 210.300 163.400 212.100 163.700 ;
        RECT 210.700 163.100 211.000 163.400 ;
        RECT 213.400 163.100 213.800 163.500 ;
        RECT 208.300 161.100 208.900 163.100 ;
        RECT 210.600 161.100 211.000 163.100 ;
        RECT 212.800 162.800 213.800 163.100 ;
        RECT 212.800 161.100 213.200 162.800 ;
        RECT 215.000 161.100 215.400 165.300 ;
        RECT 216.600 161.100 217.000 165.800 ;
        RECT 218.200 165.200 218.500 165.800 ;
        RECT 217.400 164.400 217.800 165.200 ;
        RECT 218.200 165.100 218.600 165.200 ;
        RECT 219.200 165.100 219.500 166.800 ;
        RECT 219.800 165.800 220.200 166.600 ;
        RECT 218.200 164.800 218.900 165.100 ;
        RECT 219.200 164.800 219.700 165.100 ;
        RECT 218.600 164.200 218.900 164.800 ;
        RECT 218.600 163.800 219.000 164.200 ;
        RECT 219.300 161.100 219.700 164.800 ;
        RECT 222.200 161.100 222.600 167.900 ;
        RECT 224.600 167.600 225.000 169.900 ;
        RECT 226.200 167.600 226.600 169.900 ;
        RECT 227.800 167.600 228.200 169.900 ;
        RECT 229.400 167.600 229.800 169.900 ;
        RECT 224.600 167.200 225.500 167.600 ;
        RECT 226.200 167.200 227.300 167.600 ;
        RECT 227.800 167.200 228.900 167.600 ;
        RECT 229.400 167.200 230.600 167.600 ;
        RECT 225.100 166.900 225.500 167.200 ;
        RECT 226.900 166.900 227.300 167.200 ;
        RECT 228.500 166.900 228.900 167.200 ;
        RECT 225.100 166.500 226.400 166.900 ;
        RECT 226.900 166.500 228.100 166.900 ;
        RECT 228.500 166.500 229.800 166.900 ;
        RECT 225.100 165.800 225.500 166.500 ;
        RECT 226.900 165.800 227.300 166.500 ;
        RECT 228.500 165.800 228.900 166.500 ;
        RECT 230.200 165.800 230.600 167.200 ;
        RECT 224.600 165.400 225.500 165.800 ;
        RECT 226.200 165.400 227.300 165.800 ;
        RECT 227.800 165.400 228.900 165.800 ;
        RECT 229.400 165.400 230.600 165.800 ;
        RECT 223.000 164.400 223.400 165.200 ;
        RECT 224.600 161.100 225.000 165.400 ;
        RECT 226.200 161.100 226.600 165.400 ;
        RECT 227.800 161.100 228.200 165.400 ;
        RECT 229.400 161.100 229.800 165.400 ;
        RECT 1.700 159.200 2.100 159.900 ;
        RECT 1.700 158.800 2.600 159.200 ;
        RECT 1.000 156.800 1.400 157.200 ;
        RECT 1.000 156.200 1.300 156.800 ;
        RECT 1.700 156.200 2.100 158.800 ;
        RECT 0.600 155.900 1.300 156.200 ;
        RECT 1.600 155.900 2.100 156.200 ;
        RECT 0.600 155.800 1.000 155.900 ;
        RECT 1.600 154.200 1.900 155.900 ;
        RECT 3.800 155.800 4.200 156.600 ;
        RECT 2.200 155.100 2.600 155.200 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 2.200 154.800 4.200 155.100 ;
        RECT 2.200 154.400 2.600 154.800 ;
        RECT 0.600 153.800 1.900 154.200 ;
        RECT 3.000 154.100 3.400 154.200 ;
        RECT 2.600 153.800 3.400 154.100 ;
        RECT 0.700 153.100 1.000 153.800 ;
        RECT 2.600 153.600 3.000 153.800 ;
        RECT 1.500 153.100 3.300 153.300 ;
        RECT 4.600 153.200 5.000 159.900 ;
        RECT 6.200 156.200 6.600 159.900 ;
        RECT 7.800 156.400 8.200 159.900 ;
        RECT 6.200 155.900 7.500 156.200 ;
        RECT 7.800 155.900 8.300 156.400 ;
        RECT 10.700 156.200 11.100 159.900 ;
        RECT 11.400 156.800 11.800 157.200 ;
        RECT 11.500 156.200 11.800 156.800 ;
        RECT 10.700 155.900 11.200 156.200 ;
        RECT 11.500 155.900 12.200 156.200 ;
        RECT 6.200 154.800 6.700 155.200 ;
        RECT 6.300 154.400 6.700 154.800 ;
        RECT 7.200 154.900 7.500 155.900 ;
        RECT 7.200 154.500 7.700 154.900 ;
        RECT 5.400 153.400 5.800 154.200 ;
        RECT 7.200 153.700 7.500 154.500 ;
        RECT 8.000 154.200 8.300 155.900 ;
        RECT 10.200 154.400 10.600 155.200 ;
        RECT 10.900 154.200 11.200 155.900 ;
        RECT 11.800 155.800 12.200 155.900 ;
        RECT 12.600 155.700 13.000 159.900 ;
        RECT 14.800 158.200 15.200 159.900 ;
        RECT 14.200 157.900 15.200 158.200 ;
        RECT 17.000 157.900 17.400 159.900 ;
        RECT 19.100 157.900 19.700 159.900 ;
        RECT 14.200 157.500 14.600 157.900 ;
        RECT 17.000 157.600 17.300 157.900 ;
        RECT 15.900 157.300 17.700 157.600 ;
        RECT 19.000 157.500 19.400 157.900 ;
        RECT 15.900 157.200 16.300 157.300 ;
        RECT 17.300 157.200 17.700 157.300 ;
        RECT 14.200 156.500 14.600 156.600 ;
        RECT 16.500 156.500 16.900 156.600 ;
        RECT 14.200 156.200 16.900 156.500 ;
        RECT 17.200 156.500 18.300 156.800 ;
        RECT 17.200 155.900 17.500 156.500 ;
        RECT 17.900 156.400 18.300 156.500 ;
        RECT 19.100 156.600 19.800 157.000 ;
        RECT 19.100 156.100 19.400 156.600 ;
        RECT 15.100 155.700 17.500 155.900 ;
        RECT 12.600 155.600 17.500 155.700 ;
        RECT 18.200 155.800 19.400 156.100 ;
        RECT 12.600 155.500 15.500 155.600 ;
        RECT 12.600 155.400 15.400 155.500 ;
        RECT 18.200 155.200 18.500 155.800 ;
        RECT 21.400 155.600 21.800 159.900 ;
        RECT 19.700 155.300 21.800 155.600 ;
        RECT 22.200 155.700 22.600 159.900 ;
        RECT 24.400 158.200 24.800 159.900 ;
        RECT 23.800 157.900 24.800 158.200 ;
        RECT 26.600 157.900 27.000 159.900 ;
        RECT 28.700 157.900 29.300 159.900 ;
        RECT 23.800 157.500 24.200 157.900 ;
        RECT 26.600 157.600 26.900 157.900 ;
        RECT 25.500 157.300 27.300 157.600 ;
        RECT 28.600 157.500 29.000 157.900 ;
        RECT 25.500 157.200 25.900 157.300 ;
        RECT 26.900 157.200 27.300 157.300 ;
        RECT 23.800 156.500 24.200 156.600 ;
        RECT 26.100 156.500 26.500 156.600 ;
        RECT 23.800 156.200 26.500 156.500 ;
        RECT 26.800 156.500 27.900 156.800 ;
        RECT 26.800 155.900 27.100 156.500 ;
        RECT 27.500 156.400 27.900 156.500 ;
        RECT 28.700 156.600 29.400 157.000 ;
        RECT 28.700 156.100 29.000 156.600 ;
        RECT 24.700 155.700 27.100 155.900 ;
        RECT 22.200 155.600 27.100 155.700 ;
        RECT 27.800 155.800 29.000 156.100 ;
        RECT 22.200 155.500 25.100 155.600 ;
        RECT 22.200 155.400 25.000 155.500 ;
        RECT 19.700 155.200 20.100 155.300 ;
        RECT 15.800 155.100 16.200 155.200 ;
        RECT 13.700 154.800 16.200 155.100 ;
        RECT 18.200 154.800 18.600 155.200 ;
        RECT 20.500 154.900 20.900 155.000 ;
        RECT 13.700 154.700 14.100 154.800 ;
        RECT 15.000 154.700 15.400 154.800 ;
        RECT 14.500 154.200 14.900 154.300 ;
        RECT 18.200 154.200 18.500 154.800 ;
        RECT 19.000 154.600 20.900 154.900 ;
        RECT 19.000 154.500 19.400 154.600 ;
        RECT 7.800 154.100 8.300 154.200 ;
        RECT 8.600 154.100 9.000 154.200 ;
        RECT 7.800 153.800 9.000 154.100 ;
        RECT 9.400 154.100 9.800 154.200 ;
        RECT 9.400 153.800 10.200 154.100 ;
        RECT 10.900 153.800 12.200 154.200 ;
        RECT 13.000 153.900 18.500 154.200 ;
        RECT 13.000 153.800 13.800 153.900 ;
        RECT 6.200 153.400 7.500 153.700 ;
        RECT 0.600 151.100 1.000 153.100 ;
        RECT 1.400 153.000 3.400 153.100 ;
        RECT 1.400 151.100 1.800 153.000 ;
        RECT 3.000 151.100 3.400 153.000 ;
        RECT 3.800 152.800 5.000 153.200 ;
        RECT 4.100 151.100 4.500 152.800 ;
        RECT 6.200 151.100 6.600 153.400 ;
        RECT 8.000 153.100 8.300 153.800 ;
        RECT 9.800 153.600 10.200 153.800 ;
        RECT 9.500 153.100 11.300 153.300 ;
        RECT 11.800 153.100 12.100 153.800 ;
        RECT 7.800 152.800 8.300 153.100 ;
        RECT 9.400 153.000 11.400 153.100 ;
        RECT 7.800 151.100 8.200 152.800 ;
        RECT 9.400 151.100 9.800 153.000 ;
        RECT 11.000 151.100 11.400 153.000 ;
        RECT 11.800 151.100 12.200 153.100 ;
        RECT 12.600 151.100 13.000 153.500 ;
        RECT 15.100 152.800 15.400 153.900 ;
        RECT 16.600 153.800 17.000 153.900 ;
        RECT 17.900 153.800 18.300 153.900 ;
        RECT 21.400 153.600 21.800 155.300 ;
        RECT 27.800 155.200 28.100 155.800 ;
        RECT 31.000 155.600 31.400 159.900 ;
        RECT 29.300 155.300 31.400 155.600 ;
        RECT 31.800 155.700 32.200 159.900 ;
        RECT 34.000 158.200 34.400 159.900 ;
        RECT 33.400 157.900 34.400 158.200 ;
        RECT 36.200 157.900 36.600 159.900 ;
        RECT 38.300 157.900 38.900 159.900 ;
        RECT 33.400 157.500 33.800 157.900 ;
        RECT 36.200 157.600 36.500 157.900 ;
        RECT 35.100 157.300 36.900 157.600 ;
        RECT 38.200 157.500 38.600 157.900 ;
        RECT 35.100 157.200 35.500 157.300 ;
        RECT 36.500 157.200 36.900 157.300 ;
        RECT 33.400 156.500 33.800 156.600 ;
        RECT 35.700 156.500 36.100 156.600 ;
        RECT 33.400 156.200 36.100 156.500 ;
        RECT 36.400 156.500 37.500 156.800 ;
        RECT 36.400 155.900 36.700 156.500 ;
        RECT 37.100 156.400 37.500 156.500 ;
        RECT 38.300 156.600 39.000 157.000 ;
        RECT 38.300 156.100 38.600 156.600 ;
        RECT 34.300 155.700 36.700 155.900 ;
        RECT 31.800 155.600 36.700 155.700 ;
        RECT 37.400 155.800 38.600 156.100 ;
        RECT 31.800 155.500 34.700 155.600 ;
        RECT 31.800 155.400 34.600 155.500 ;
        RECT 29.300 155.200 29.700 155.300 ;
        RECT 25.400 155.100 25.800 155.200 ;
        RECT 23.300 154.800 25.800 155.100 ;
        RECT 27.800 154.800 28.200 155.200 ;
        RECT 30.100 154.900 30.500 155.000 ;
        RECT 23.300 154.700 23.700 154.800 ;
        RECT 24.100 154.200 24.500 154.300 ;
        RECT 27.800 154.200 28.100 154.800 ;
        RECT 28.600 154.600 30.500 154.900 ;
        RECT 28.600 154.500 29.000 154.600 ;
        RECT 22.600 153.900 28.100 154.200 ;
        RECT 22.600 153.800 23.400 153.900 ;
        RECT 19.900 153.300 21.800 153.600 ;
        RECT 19.900 153.200 20.300 153.300 ;
        RECT 14.200 152.100 14.600 152.500 ;
        RECT 15.000 152.400 15.400 152.800 ;
        RECT 15.900 152.700 16.300 152.800 ;
        RECT 15.900 152.400 17.300 152.700 ;
        RECT 17.000 152.100 17.300 152.400 ;
        RECT 19.000 152.100 19.400 152.500 ;
        RECT 14.200 151.800 15.200 152.100 ;
        RECT 14.800 151.100 15.200 151.800 ;
        RECT 17.000 151.100 17.400 152.100 ;
        RECT 19.000 151.800 19.700 152.100 ;
        RECT 19.100 151.100 19.700 151.800 ;
        RECT 21.400 151.100 21.800 153.300 ;
        RECT 22.200 151.100 22.600 153.500 ;
        RECT 24.700 152.800 25.000 153.900 ;
        RECT 27.500 153.800 27.900 153.900 ;
        RECT 31.000 153.600 31.400 155.300 ;
        RECT 35.000 155.100 35.400 155.200 ;
        RECT 35.800 155.100 36.200 155.200 ;
        RECT 32.900 154.800 36.200 155.100 ;
        RECT 32.900 154.700 33.300 154.800 ;
        RECT 33.700 154.200 34.100 154.300 ;
        RECT 37.400 154.200 37.700 155.800 ;
        RECT 40.600 155.600 41.000 159.900 ;
        RECT 44.300 157.200 44.700 159.900 ;
        RECT 43.800 156.800 44.700 157.200 ;
        RECT 45.000 156.800 45.400 157.200 ;
        RECT 44.300 156.200 44.700 156.800 ;
        RECT 45.100 156.200 45.400 156.800 ;
        RECT 46.600 156.800 47.000 157.200 ;
        RECT 46.600 156.200 46.900 156.800 ;
        RECT 47.300 156.200 47.700 159.900 ;
        RECT 51.300 156.400 51.700 159.900 ;
        RECT 53.400 157.500 53.800 159.500 ;
        RECT 44.300 155.900 44.800 156.200 ;
        RECT 45.100 155.900 45.800 156.200 ;
        RECT 38.900 155.300 41.000 155.600 ;
        RECT 38.900 155.200 39.300 155.300 ;
        RECT 39.700 154.900 40.100 155.000 ;
        RECT 38.200 154.600 40.100 154.900 ;
        RECT 38.200 154.500 38.600 154.600 ;
        RECT 32.200 153.900 37.700 154.200 ;
        RECT 32.200 153.800 33.000 153.900 ;
        RECT 29.500 153.300 31.400 153.600 ;
        RECT 29.500 153.200 29.900 153.300 ;
        RECT 23.800 152.100 24.200 152.500 ;
        RECT 24.600 152.400 25.000 152.800 ;
        RECT 25.500 152.700 25.900 152.800 ;
        RECT 25.500 152.400 26.900 152.700 ;
        RECT 26.600 152.100 26.900 152.400 ;
        RECT 28.600 152.100 29.000 152.500 ;
        RECT 23.800 151.800 24.800 152.100 ;
        RECT 24.400 151.100 24.800 151.800 ;
        RECT 26.600 151.100 27.000 152.100 ;
        RECT 28.600 151.800 29.300 152.100 ;
        RECT 28.700 151.100 29.300 151.800 ;
        RECT 31.000 151.100 31.400 153.300 ;
        RECT 31.800 151.100 32.200 153.500 ;
        RECT 34.300 152.800 34.600 153.900 ;
        RECT 37.100 153.800 37.500 153.900 ;
        RECT 40.600 153.600 41.000 155.300 ;
        RECT 43.800 154.400 44.200 155.200 ;
        RECT 44.500 154.200 44.800 155.900 ;
        RECT 45.400 155.800 45.800 155.900 ;
        RECT 46.200 155.900 46.900 156.200 ;
        RECT 47.200 155.900 47.700 156.200 ;
        RECT 50.900 156.100 51.700 156.400 ;
        RECT 46.200 155.800 46.600 155.900 ;
        RECT 45.400 155.100 45.700 155.800 ;
        RECT 47.200 155.100 47.500 155.900 ;
        RECT 45.400 154.800 47.500 155.100 ;
        RECT 47.200 154.200 47.500 154.800 ;
        RECT 47.800 154.400 48.200 155.200 ;
        RECT 49.400 155.100 49.800 155.200 ;
        RECT 50.200 155.100 50.600 155.600 ;
        RECT 49.400 154.800 50.600 155.100 ;
        RECT 50.900 154.200 51.200 156.100 ;
        RECT 53.500 155.800 53.800 157.500 ;
        RECT 51.900 155.500 53.800 155.800 ;
        RECT 54.200 155.700 54.600 159.900 ;
        RECT 56.400 158.200 56.800 159.900 ;
        RECT 55.800 157.900 56.800 158.200 ;
        RECT 58.600 157.900 59.000 159.900 ;
        RECT 60.700 157.900 61.300 159.900 ;
        RECT 55.800 157.500 56.200 157.900 ;
        RECT 58.600 157.600 58.900 157.900 ;
        RECT 57.500 157.300 59.300 157.600 ;
        RECT 60.600 157.500 61.000 157.900 ;
        RECT 57.500 157.200 57.900 157.300 ;
        RECT 58.900 157.200 59.300 157.300 ;
        RECT 61.100 157.000 61.800 157.200 ;
        RECT 60.700 156.800 61.800 157.000 ;
        RECT 55.800 156.500 56.200 156.600 ;
        RECT 58.100 156.500 58.500 156.600 ;
        RECT 55.800 156.200 58.500 156.500 ;
        RECT 58.800 156.500 59.900 156.800 ;
        RECT 58.800 155.900 59.100 156.500 ;
        RECT 59.500 156.400 59.900 156.500 ;
        RECT 60.700 156.600 61.400 156.800 ;
        RECT 60.700 156.100 61.000 156.600 ;
        RECT 56.700 155.700 59.100 155.900 ;
        RECT 54.200 155.600 59.100 155.700 ;
        RECT 59.800 155.800 61.000 156.100 ;
        RECT 54.200 155.500 57.100 155.600 ;
        RECT 51.900 154.500 52.200 155.500 ;
        RECT 54.200 155.400 57.000 155.500 ;
        RECT 43.000 154.100 43.400 154.200 ;
        RECT 43.000 153.800 43.800 154.100 ;
        RECT 44.500 153.800 45.800 154.200 ;
        RECT 46.200 153.800 47.500 154.200 ;
        RECT 48.600 154.100 49.000 154.200 ;
        RECT 48.200 153.800 49.000 154.100 ;
        RECT 50.200 153.800 51.200 154.200 ;
        RECT 51.500 154.100 52.200 154.500 ;
        RECT 52.600 154.400 53.000 155.200 ;
        RECT 53.400 154.400 53.800 155.200 ;
        RECT 57.400 155.100 57.800 155.200 ;
        RECT 58.200 155.100 58.600 155.200 ;
        RECT 55.300 154.800 58.600 155.100 ;
        RECT 55.300 154.700 55.700 154.800 ;
        RECT 56.100 154.200 56.500 154.300 ;
        RECT 59.800 154.200 60.100 155.800 ;
        RECT 63.000 155.600 63.400 159.900 ;
        RECT 65.100 156.200 65.500 159.900 ;
        RECT 65.800 156.800 66.200 157.200 ;
        RECT 65.900 156.200 66.200 156.800 ;
        RECT 64.600 155.800 65.600 156.200 ;
        RECT 65.900 155.900 66.600 156.200 ;
        RECT 61.300 155.300 63.400 155.600 ;
        RECT 61.300 155.200 61.700 155.300 ;
        RECT 62.100 154.900 62.500 155.000 ;
        RECT 60.600 154.600 62.500 154.900 ;
        RECT 60.600 154.500 61.000 154.600 ;
        RECT 43.400 153.600 43.800 153.800 ;
        RECT 39.100 153.300 41.000 153.600 ;
        RECT 39.100 153.200 39.500 153.300 ;
        RECT 33.400 152.100 33.800 152.500 ;
        RECT 34.200 152.400 34.600 152.800 ;
        RECT 35.100 152.700 35.500 152.800 ;
        RECT 35.100 152.400 36.500 152.700 ;
        RECT 36.200 152.100 36.500 152.400 ;
        RECT 38.200 152.100 38.600 152.500 ;
        RECT 33.400 151.800 34.400 152.100 ;
        RECT 34.000 151.100 34.400 151.800 ;
        RECT 36.200 151.100 36.600 152.100 ;
        RECT 38.200 151.800 38.900 152.100 ;
        RECT 38.300 151.100 38.900 151.800 ;
        RECT 40.600 151.100 41.000 153.300 ;
        RECT 43.100 153.100 44.900 153.300 ;
        RECT 45.400 153.100 45.700 153.800 ;
        RECT 46.300 153.100 46.600 153.800 ;
        RECT 48.200 153.600 48.600 153.800 ;
        RECT 50.900 153.500 51.200 153.800 ;
        RECT 51.700 153.900 52.200 154.100 ;
        RECT 54.600 153.900 60.100 154.200 ;
        RECT 51.700 153.600 53.800 153.900 ;
        RECT 54.600 153.800 55.400 153.900 ;
        RECT 50.900 153.300 51.300 153.500 ;
        RECT 47.100 153.100 48.900 153.300 ;
        RECT 43.000 153.000 45.000 153.100 ;
        RECT 43.000 151.100 43.400 153.000 ;
        RECT 44.600 151.100 45.000 153.000 ;
        RECT 45.400 151.100 45.800 153.100 ;
        RECT 46.200 151.100 46.600 153.100 ;
        RECT 47.000 153.000 49.000 153.100 ;
        RECT 50.900 153.000 51.700 153.300 ;
        RECT 47.000 151.100 47.400 153.000 ;
        RECT 48.600 151.100 49.000 153.000 ;
        RECT 51.300 152.200 51.700 153.000 ;
        RECT 53.500 152.500 53.800 153.600 ;
        RECT 51.000 151.800 51.700 152.200 ;
        RECT 51.300 151.500 51.700 151.800 ;
        RECT 53.400 151.500 53.800 152.500 ;
        RECT 54.200 151.100 54.600 153.500 ;
        RECT 56.700 152.800 57.000 153.900 ;
        RECT 58.200 153.800 58.600 153.900 ;
        RECT 59.500 153.800 59.900 153.900 ;
        RECT 63.000 153.600 63.400 155.300 ;
        RECT 64.600 154.400 65.000 155.200 ;
        RECT 65.300 154.200 65.600 155.800 ;
        RECT 66.200 155.800 66.600 155.900 ;
        RECT 67.000 155.800 67.400 156.600 ;
        RECT 66.200 155.100 66.500 155.800 ;
        RECT 67.800 155.100 68.200 159.900 ;
        RECT 66.200 154.800 68.200 155.100 ;
        RECT 63.800 154.100 64.200 154.200 ;
        RECT 63.800 153.800 64.600 154.100 ;
        RECT 65.300 153.800 66.600 154.200 ;
        RECT 64.200 153.600 64.600 153.800 ;
        RECT 61.500 153.300 63.400 153.600 ;
        RECT 61.500 153.200 61.900 153.300 ;
        RECT 55.800 152.100 56.200 152.500 ;
        RECT 56.600 152.400 57.000 152.800 ;
        RECT 57.500 152.700 57.900 152.800 ;
        RECT 57.500 152.400 58.900 152.700 ;
        RECT 58.600 152.100 58.900 152.400 ;
        RECT 60.600 152.100 61.000 152.500 ;
        RECT 55.800 151.800 56.800 152.100 ;
        RECT 56.400 151.100 56.800 151.800 ;
        RECT 58.600 151.100 59.000 152.100 ;
        RECT 60.600 151.800 61.300 152.100 ;
        RECT 60.700 151.100 61.300 151.800 ;
        RECT 63.000 151.100 63.400 153.300 ;
        RECT 63.900 153.100 65.700 153.300 ;
        RECT 66.200 153.100 66.500 153.800 ;
        RECT 67.800 153.100 68.200 154.800 ;
        RECT 68.600 154.100 69.000 154.200 ;
        RECT 68.600 153.800 69.700 154.100 ;
        RECT 68.600 153.400 69.000 153.800 ;
        RECT 63.800 153.000 65.800 153.100 ;
        RECT 63.800 151.100 64.200 153.000 ;
        RECT 65.400 151.100 65.800 153.000 ;
        RECT 66.200 151.100 66.600 153.100 ;
        RECT 67.300 152.800 68.200 153.100 ;
        RECT 69.400 153.200 69.700 153.800 ;
        RECT 67.300 151.100 67.700 152.800 ;
        RECT 69.400 152.400 69.800 153.200 ;
        RECT 70.200 151.100 70.600 159.900 ;
        RECT 71.800 156.400 72.200 159.900 ;
        RECT 71.700 155.900 72.200 156.400 ;
        RECT 73.400 156.200 73.800 159.900 ;
        RECT 72.500 155.900 73.800 156.200 ;
        RECT 71.000 154.800 71.400 155.200 ;
        RECT 71.000 154.100 71.300 154.800 ;
        RECT 71.700 154.200 72.000 155.900 ;
        RECT 72.500 154.900 72.800 155.900 ;
        RECT 74.200 155.700 74.600 159.900 ;
        RECT 76.400 158.200 76.800 159.900 ;
        RECT 75.800 157.900 76.800 158.200 ;
        RECT 78.600 157.900 79.000 159.900 ;
        RECT 80.700 157.900 81.300 159.900 ;
        RECT 75.800 157.500 76.200 157.900 ;
        RECT 78.600 157.600 78.900 157.900 ;
        RECT 77.500 157.300 79.300 157.600 ;
        RECT 80.600 157.500 81.000 157.900 ;
        RECT 77.500 157.200 77.900 157.300 ;
        RECT 78.900 157.200 79.300 157.300 ;
        RECT 75.800 156.500 76.200 156.600 ;
        RECT 78.100 156.500 78.500 156.600 ;
        RECT 75.800 156.200 78.500 156.500 ;
        RECT 78.800 156.500 79.900 156.800 ;
        RECT 78.800 155.900 79.100 156.500 ;
        RECT 79.500 156.400 79.900 156.500 ;
        RECT 80.700 156.600 81.400 157.000 ;
        RECT 80.700 156.100 81.000 156.600 ;
        RECT 76.700 155.700 79.100 155.900 ;
        RECT 74.200 155.600 79.100 155.700 ;
        RECT 79.800 155.800 81.000 156.100 ;
        RECT 74.200 155.500 77.100 155.600 ;
        RECT 74.200 155.400 77.000 155.500 ;
        RECT 72.300 154.500 72.800 154.900 ;
        RECT 71.700 154.100 72.200 154.200 ;
        RECT 71.000 153.800 72.200 154.100 ;
        RECT 71.700 153.100 72.000 153.800 ;
        RECT 72.500 153.700 72.800 154.500 ;
        RECT 73.300 154.800 73.800 155.200 ;
        RECT 77.400 155.100 77.800 155.200 ;
        RECT 79.000 155.100 79.400 155.200 ;
        RECT 75.300 154.800 79.400 155.100 ;
        RECT 73.300 154.400 73.700 154.800 ;
        RECT 75.300 154.700 75.700 154.800 ;
        RECT 76.100 154.200 76.500 154.300 ;
        RECT 79.800 154.200 80.100 155.800 ;
        RECT 83.000 155.600 83.400 159.900 ;
        RECT 85.100 156.200 85.500 159.900 ;
        RECT 85.800 156.800 86.200 157.200 ;
        RECT 85.900 156.200 86.200 156.800 ;
        RECT 85.100 155.900 85.600 156.200 ;
        RECT 85.900 155.900 86.600 156.200 ;
        RECT 81.300 155.300 83.400 155.600 ;
        RECT 81.300 155.200 81.700 155.300 ;
        RECT 82.100 154.900 82.500 155.000 ;
        RECT 80.600 154.600 82.500 154.900 ;
        RECT 80.600 154.500 81.000 154.600 ;
        RECT 74.600 153.900 80.200 154.200 ;
        RECT 74.600 153.800 75.400 153.900 ;
        RECT 72.500 153.400 73.800 153.700 ;
        RECT 71.700 152.800 72.200 153.100 ;
        RECT 71.800 151.100 72.200 152.800 ;
        RECT 73.400 151.100 73.800 153.400 ;
        RECT 74.200 151.100 74.600 153.500 ;
        RECT 76.700 152.800 77.000 153.900 ;
        RECT 79.500 153.800 80.200 153.900 ;
        RECT 83.000 153.600 83.400 155.300 ;
        RECT 85.300 155.200 85.600 155.900 ;
        RECT 86.200 155.800 86.600 155.900 ;
        RECT 88.600 155.700 89.000 159.900 ;
        RECT 90.800 158.200 91.200 159.900 ;
        RECT 90.200 157.900 91.200 158.200 ;
        RECT 93.000 157.900 93.400 159.900 ;
        RECT 95.100 157.900 95.700 159.900 ;
        RECT 90.200 157.500 90.600 157.900 ;
        RECT 93.000 157.600 93.300 157.900 ;
        RECT 91.900 157.300 93.700 157.600 ;
        RECT 95.000 157.500 95.400 157.900 ;
        RECT 91.900 157.200 92.300 157.300 ;
        RECT 93.300 157.200 93.700 157.300 ;
        RECT 95.500 157.000 96.200 157.200 ;
        RECT 95.100 156.800 96.200 157.000 ;
        RECT 90.200 156.500 90.600 156.600 ;
        RECT 92.500 156.500 92.900 156.600 ;
        RECT 90.200 156.200 92.900 156.500 ;
        RECT 93.200 156.500 94.300 156.800 ;
        RECT 93.200 155.900 93.500 156.500 ;
        RECT 93.900 156.400 94.300 156.500 ;
        RECT 95.100 156.600 95.800 156.800 ;
        RECT 95.100 156.100 95.400 156.600 ;
        RECT 91.100 155.700 93.500 155.900 ;
        RECT 88.600 155.600 93.500 155.700 ;
        RECT 94.200 155.800 95.400 156.100 ;
        RECT 88.600 155.500 91.500 155.600 ;
        RECT 88.600 155.400 91.400 155.500 ;
        RECT 84.600 154.400 85.000 155.200 ;
        RECT 85.300 154.800 85.800 155.200 ;
        RECT 91.800 155.100 92.200 155.200 ;
        RECT 92.600 155.100 93.000 155.200 ;
        RECT 89.700 154.800 93.000 155.100 ;
        RECT 85.300 154.200 85.600 154.800 ;
        RECT 89.700 154.700 90.100 154.800 ;
        RECT 90.500 154.200 90.900 154.300 ;
        RECT 94.200 154.200 94.500 155.800 ;
        RECT 97.400 155.600 97.800 159.900 ;
        RECT 99.000 157.100 99.400 159.900 ;
        RECT 99.800 157.100 100.200 157.200 ;
        RECT 99.000 156.800 100.200 157.100 ;
        RECT 101.000 156.800 101.400 157.200 ;
        RECT 98.200 155.800 98.600 156.600 ;
        RECT 95.700 155.300 97.800 155.600 ;
        RECT 95.700 155.200 96.100 155.300 ;
        RECT 96.500 154.900 96.900 155.000 ;
        RECT 95.000 154.600 96.900 154.900 ;
        RECT 95.000 154.500 95.400 154.600 ;
        RECT 83.800 154.100 84.200 154.200 ;
        RECT 83.800 153.800 84.600 154.100 ;
        RECT 85.300 153.800 86.600 154.200 ;
        RECT 89.000 153.900 94.500 154.200 ;
        RECT 89.000 153.800 89.800 153.900 ;
        RECT 84.200 153.600 84.600 153.800 ;
        RECT 81.500 153.300 83.400 153.600 ;
        RECT 81.500 153.200 81.900 153.300 ;
        RECT 75.800 152.100 76.200 152.500 ;
        RECT 76.600 152.400 77.000 152.800 ;
        RECT 77.500 152.700 77.900 152.800 ;
        RECT 77.500 152.400 78.900 152.700 ;
        RECT 78.600 152.100 78.900 152.400 ;
        RECT 80.600 152.100 81.000 152.500 ;
        RECT 75.800 151.800 76.800 152.100 ;
        RECT 76.400 151.100 76.800 151.800 ;
        RECT 78.600 151.100 79.000 152.100 ;
        RECT 80.600 151.800 81.300 152.100 ;
        RECT 80.700 151.100 81.300 151.800 ;
        RECT 83.000 151.100 83.400 153.300 ;
        RECT 83.900 153.100 85.700 153.300 ;
        RECT 86.200 153.100 86.500 153.800 ;
        RECT 83.800 153.000 85.800 153.100 ;
        RECT 83.800 151.100 84.200 153.000 ;
        RECT 85.400 151.100 85.800 153.000 ;
        RECT 86.200 151.100 86.600 153.100 ;
        RECT 88.600 151.100 89.000 153.500 ;
        RECT 91.100 152.800 91.400 153.900 ;
        RECT 93.900 153.800 94.300 153.900 ;
        RECT 97.400 153.600 97.800 155.300 ;
        RECT 98.200 154.800 98.600 155.200 ;
        RECT 98.200 154.100 98.500 154.800 ;
        RECT 99.000 154.100 99.400 156.800 ;
        RECT 101.000 156.200 101.300 156.800 ;
        RECT 101.700 156.200 102.100 159.900 ;
        RECT 100.600 155.900 101.300 156.200 ;
        RECT 101.600 155.900 102.100 156.200 ;
        RECT 100.600 155.800 101.000 155.900 ;
        RECT 101.600 155.200 101.900 155.900 ;
        RECT 103.800 155.800 104.200 156.600 ;
        RECT 101.400 154.800 101.900 155.200 ;
        RECT 101.600 154.200 101.900 154.800 ;
        RECT 102.200 154.400 102.600 155.200 ;
        RECT 98.200 153.800 99.400 154.100 ;
        RECT 95.900 153.300 97.800 153.600 ;
        RECT 95.900 153.200 96.300 153.300 ;
        RECT 90.200 152.100 90.600 152.500 ;
        RECT 91.000 152.400 91.400 152.800 ;
        RECT 91.900 152.700 92.300 152.800 ;
        RECT 91.900 152.400 93.300 152.700 ;
        RECT 93.000 152.100 93.300 152.400 ;
        RECT 95.000 152.100 95.400 152.500 ;
        RECT 90.200 151.800 91.200 152.100 ;
        RECT 90.800 151.100 91.200 151.800 ;
        RECT 93.000 151.100 93.400 152.100 ;
        RECT 95.000 151.800 95.700 152.100 ;
        RECT 95.100 151.100 95.700 151.800 ;
        RECT 97.400 151.100 97.800 153.300 ;
        RECT 99.000 153.100 99.400 153.800 ;
        RECT 99.800 153.400 100.200 154.200 ;
        RECT 100.600 153.800 101.900 154.200 ;
        RECT 103.000 154.100 103.400 154.200 ;
        RECT 102.600 153.800 103.400 154.100 ;
        RECT 100.700 153.100 101.000 153.800 ;
        RECT 102.600 153.600 103.000 153.800 ;
        RECT 101.500 153.100 103.300 153.300 ;
        RECT 104.600 153.100 105.000 159.900 ;
        RECT 106.200 155.700 106.600 159.900 ;
        RECT 108.400 158.200 108.800 159.900 ;
        RECT 107.800 157.900 108.800 158.200 ;
        RECT 110.600 157.900 111.000 159.900 ;
        RECT 112.700 157.900 113.300 159.900 ;
        RECT 107.800 157.500 108.200 157.900 ;
        RECT 110.600 157.600 110.900 157.900 ;
        RECT 109.500 157.300 111.300 157.600 ;
        RECT 112.600 157.500 113.000 157.900 ;
        RECT 109.500 157.200 109.900 157.300 ;
        RECT 110.900 157.200 111.300 157.300 ;
        RECT 107.800 156.500 108.200 156.600 ;
        RECT 110.100 156.500 110.500 156.600 ;
        RECT 107.800 156.200 110.500 156.500 ;
        RECT 110.800 156.500 111.900 156.800 ;
        RECT 110.800 155.900 111.100 156.500 ;
        RECT 111.500 156.400 111.900 156.500 ;
        RECT 112.700 156.600 113.400 157.000 ;
        RECT 112.700 156.100 113.000 156.600 ;
        RECT 108.700 155.700 111.100 155.900 ;
        RECT 106.200 155.600 111.100 155.700 ;
        RECT 111.800 155.800 113.000 156.100 ;
        RECT 106.200 155.500 109.100 155.600 ;
        RECT 106.200 155.400 109.000 155.500 ;
        RECT 111.800 155.200 112.100 155.800 ;
        RECT 115.000 155.600 115.400 159.900 ;
        RECT 113.300 155.300 115.400 155.600 ;
        RECT 115.800 155.700 116.200 159.900 ;
        RECT 118.000 158.200 118.400 159.900 ;
        RECT 117.400 157.900 118.400 158.200 ;
        RECT 120.200 157.900 120.600 159.900 ;
        RECT 122.300 157.900 122.900 159.900 ;
        RECT 117.400 157.500 117.800 157.900 ;
        RECT 120.200 157.600 120.500 157.900 ;
        RECT 119.100 157.300 120.900 157.600 ;
        RECT 122.200 157.500 122.600 157.900 ;
        RECT 119.100 157.200 119.500 157.300 ;
        RECT 120.500 157.200 120.900 157.300 ;
        RECT 117.400 156.500 117.800 156.600 ;
        RECT 119.700 156.500 120.100 156.600 ;
        RECT 117.400 156.200 120.100 156.500 ;
        RECT 120.400 156.500 121.500 156.800 ;
        RECT 120.400 155.900 120.700 156.500 ;
        RECT 121.100 156.400 121.500 156.500 ;
        RECT 122.300 156.600 123.000 157.000 ;
        RECT 122.300 156.100 122.600 156.600 ;
        RECT 118.300 155.700 120.700 155.900 ;
        RECT 115.800 155.600 120.700 155.700 ;
        RECT 121.400 155.800 122.600 156.100 ;
        RECT 115.800 155.500 118.700 155.600 ;
        RECT 115.800 155.400 118.600 155.500 ;
        RECT 113.300 155.200 113.700 155.300 ;
        RECT 109.400 155.100 109.800 155.200 ;
        RECT 107.300 154.800 109.800 155.100 ;
        RECT 111.800 154.800 112.200 155.200 ;
        RECT 114.100 154.900 114.500 155.000 ;
        RECT 107.300 154.700 107.700 154.800 ;
        RECT 108.100 154.200 108.500 154.300 ;
        RECT 111.800 154.200 112.100 154.800 ;
        RECT 112.600 154.600 114.500 154.900 ;
        RECT 112.600 154.500 113.000 154.600 ;
        RECT 105.400 153.400 105.800 154.200 ;
        RECT 106.600 153.900 112.100 154.200 ;
        RECT 106.600 153.800 107.400 153.900 ;
        RECT 108.600 153.800 109.000 153.900 ;
        RECT 111.500 153.800 111.900 153.900 ;
        RECT 98.500 152.800 99.400 153.100 ;
        RECT 98.500 151.100 98.900 152.800 ;
        RECT 100.600 151.100 101.000 153.100 ;
        RECT 101.400 153.000 103.400 153.100 ;
        RECT 101.400 151.100 101.800 153.000 ;
        RECT 103.000 151.100 103.400 153.000 ;
        RECT 104.100 152.800 105.000 153.100 ;
        RECT 104.100 152.200 104.500 152.800 ;
        RECT 104.100 151.800 105.000 152.200 ;
        RECT 104.100 151.100 104.500 151.800 ;
        RECT 106.200 151.100 106.600 153.500 ;
        RECT 108.700 152.800 109.000 153.800 ;
        RECT 115.000 153.600 115.400 155.300 ;
        RECT 121.400 155.200 121.700 155.800 ;
        RECT 124.600 155.600 125.000 159.900 ;
        RECT 126.200 156.400 126.600 159.900 ;
        RECT 122.900 155.300 125.000 155.600 ;
        RECT 122.900 155.200 123.300 155.300 ;
        RECT 119.000 155.100 119.400 155.200 ;
        RECT 116.900 154.800 119.400 155.100 ;
        RECT 121.400 154.800 121.800 155.200 ;
        RECT 123.700 154.900 124.100 155.000 ;
        RECT 116.900 154.700 117.300 154.800 ;
        RECT 117.700 154.200 118.100 154.300 ;
        RECT 121.400 154.200 121.700 154.800 ;
        RECT 122.200 154.600 124.100 154.900 ;
        RECT 122.200 154.500 122.600 154.600 ;
        RECT 116.200 153.900 121.700 154.200 ;
        RECT 116.200 153.800 117.000 153.900 ;
        RECT 113.500 153.300 115.400 153.600 ;
        RECT 113.500 153.200 113.900 153.300 ;
        RECT 107.800 152.100 108.200 152.500 ;
        RECT 108.600 152.400 109.000 152.800 ;
        RECT 109.500 152.700 109.900 152.800 ;
        RECT 109.500 152.400 110.900 152.700 ;
        RECT 110.600 152.100 110.900 152.400 ;
        RECT 112.600 152.100 113.000 152.500 ;
        RECT 107.800 151.800 108.800 152.100 ;
        RECT 108.400 151.100 108.800 151.800 ;
        RECT 110.600 151.100 111.000 152.100 ;
        RECT 112.600 151.800 113.300 152.100 ;
        RECT 112.700 151.100 113.300 151.800 ;
        RECT 115.000 151.100 115.400 153.300 ;
        RECT 115.800 151.100 116.200 153.500 ;
        RECT 118.300 152.800 118.600 153.900 ;
        RECT 119.800 153.800 120.200 153.900 ;
        RECT 121.100 153.800 121.500 153.900 ;
        RECT 124.600 153.600 125.000 155.300 ;
        RECT 123.100 153.300 125.000 153.600 ;
        RECT 123.100 153.200 123.500 153.300 ;
        RECT 117.400 152.100 117.800 152.500 ;
        RECT 118.200 152.400 118.600 152.800 ;
        RECT 119.100 152.700 119.500 152.800 ;
        RECT 119.100 152.400 120.500 152.700 ;
        RECT 120.200 152.100 120.500 152.400 ;
        RECT 122.200 152.100 122.600 152.500 ;
        RECT 117.400 151.800 118.400 152.100 ;
        RECT 118.000 151.100 118.400 151.800 ;
        RECT 120.200 151.100 120.600 152.100 ;
        RECT 122.200 151.800 122.900 152.100 ;
        RECT 122.300 151.100 122.900 151.800 ;
        RECT 124.600 151.100 125.000 153.300 ;
        RECT 126.100 155.900 126.600 156.400 ;
        RECT 127.800 156.200 128.200 159.900 ;
        RECT 126.900 155.900 128.200 156.200 ;
        RECT 126.100 154.200 126.400 155.900 ;
        RECT 126.900 154.900 127.200 155.900 ;
        RECT 128.600 155.800 129.000 156.600 ;
        RECT 126.700 154.500 127.200 154.900 ;
        RECT 126.100 153.800 126.600 154.200 ;
        RECT 126.100 153.100 126.400 153.800 ;
        RECT 126.900 153.700 127.200 154.500 ;
        RECT 127.700 154.800 128.200 155.200 ;
        RECT 127.700 154.400 128.100 154.800 ;
        RECT 126.900 153.400 128.200 153.700 ;
        RECT 126.100 152.800 126.600 153.100 ;
        RECT 126.200 151.100 126.600 152.800 ;
        RECT 127.800 151.100 128.200 153.400 ;
        RECT 129.400 153.100 129.800 159.900 ;
        RECT 131.000 155.700 131.400 159.900 ;
        RECT 133.200 158.200 133.600 159.900 ;
        RECT 132.600 157.900 133.600 158.200 ;
        RECT 135.400 157.900 135.800 159.900 ;
        RECT 137.500 157.900 138.100 159.900 ;
        RECT 132.600 157.500 133.000 157.900 ;
        RECT 135.400 157.600 135.700 157.900 ;
        RECT 134.300 157.300 136.100 157.600 ;
        RECT 137.400 157.500 137.800 157.900 ;
        RECT 134.300 157.200 134.700 157.300 ;
        RECT 135.700 157.200 136.100 157.300 ;
        RECT 137.900 157.000 138.600 157.200 ;
        RECT 137.500 156.800 138.600 157.000 ;
        RECT 132.600 156.500 133.000 156.600 ;
        RECT 134.900 156.500 135.300 156.600 ;
        RECT 132.600 156.200 135.300 156.500 ;
        RECT 135.600 156.500 136.700 156.800 ;
        RECT 135.600 155.900 135.900 156.500 ;
        RECT 136.300 156.400 136.700 156.500 ;
        RECT 137.500 156.600 138.200 156.800 ;
        RECT 137.500 156.100 137.800 156.600 ;
        RECT 133.500 155.700 135.900 155.900 ;
        RECT 131.000 155.600 135.900 155.700 ;
        RECT 136.600 155.800 137.800 156.100 ;
        RECT 131.000 155.500 133.900 155.600 ;
        RECT 131.000 155.400 133.800 155.500 ;
        RECT 134.200 155.100 134.600 155.200 ;
        RECT 135.800 155.100 136.200 155.200 ;
        RECT 132.100 154.800 136.200 155.100 ;
        RECT 132.100 154.700 132.500 154.800 ;
        RECT 132.900 154.200 133.300 154.300 ;
        RECT 136.600 154.200 136.900 155.800 ;
        RECT 139.800 155.600 140.200 159.900 ;
        RECT 138.100 155.300 140.200 155.600 ;
        RECT 138.100 155.200 138.500 155.300 ;
        RECT 138.900 154.900 139.300 155.000 ;
        RECT 137.400 154.600 139.300 154.900 ;
        RECT 137.400 154.500 137.800 154.600 ;
        RECT 130.200 153.400 130.600 154.200 ;
        RECT 131.400 153.900 136.900 154.200 ;
        RECT 131.400 153.800 132.200 153.900 ;
        RECT 128.900 152.800 129.800 153.100 ;
        RECT 128.900 151.100 129.300 152.800 ;
        RECT 131.000 151.100 131.400 153.500 ;
        RECT 133.500 152.800 133.800 153.900 ;
        RECT 136.300 153.800 136.700 153.900 ;
        RECT 139.800 153.600 140.200 155.300 ;
        RECT 138.300 153.300 140.200 153.600 ;
        RECT 138.300 153.200 138.700 153.300 ;
        RECT 132.600 152.100 133.000 152.500 ;
        RECT 133.400 152.400 133.800 152.800 ;
        RECT 134.300 152.700 134.700 152.800 ;
        RECT 134.300 152.400 135.700 152.700 ;
        RECT 135.400 152.100 135.700 152.400 ;
        RECT 137.400 152.100 137.800 152.500 ;
        RECT 132.600 151.800 133.600 152.100 ;
        RECT 133.200 151.100 133.600 151.800 ;
        RECT 135.400 151.100 135.800 152.100 ;
        RECT 137.400 151.800 138.100 152.100 ;
        RECT 137.500 151.100 138.100 151.800 ;
        RECT 139.800 151.100 140.200 153.300 ;
        RECT 140.600 153.100 141.000 153.200 ;
        RECT 142.200 153.100 142.600 153.200 ;
        RECT 140.600 152.800 142.600 153.100 ;
        RECT 142.200 152.400 142.600 152.800 ;
        RECT 143.000 151.100 143.400 159.900 ;
        RECT 143.800 155.800 144.200 156.600 ;
        RECT 144.600 156.100 145.000 159.900 ;
        RECT 145.400 156.800 145.800 157.200 ;
        RECT 145.400 156.100 145.700 156.800 ;
        RECT 144.600 155.800 145.700 156.100 ;
        RECT 147.500 156.200 147.900 159.900 ;
        RECT 148.200 156.800 148.600 157.200 ;
        RECT 148.300 156.200 148.600 156.800 ;
        RECT 149.400 156.200 149.800 159.900 ;
        RECT 151.000 156.200 151.400 159.900 ;
        RECT 147.500 155.900 148.000 156.200 ;
        RECT 148.300 155.900 149.000 156.200 ;
        RECT 149.400 155.900 151.400 156.200 ;
        RECT 151.800 155.900 152.200 159.900 ;
        RECT 153.400 156.400 153.800 159.900 ;
        RECT 153.300 155.900 153.800 156.400 ;
        RECT 155.000 156.200 155.400 159.900 ;
        RECT 154.100 155.900 155.400 156.200 ;
        RECT 144.600 153.100 145.000 155.800 ;
        RECT 147.000 154.400 147.400 155.200 ;
        RECT 147.700 154.200 148.000 155.900 ;
        RECT 148.600 155.800 149.000 155.900 ;
        RECT 149.800 155.200 150.200 155.400 ;
        RECT 151.800 155.200 152.100 155.900 ;
        RECT 149.400 154.900 150.200 155.200 ;
        RECT 151.000 154.900 152.200 155.200 ;
        RECT 149.400 154.800 149.800 154.900 ;
        RECT 145.400 153.400 145.800 154.200 ;
        RECT 146.200 154.100 146.600 154.200 ;
        RECT 147.700 154.100 149.000 154.200 ;
        RECT 150.200 154.100 150.600 154.600 ;
        RECT 146.200 153.800 147.000 154.100 ;
        RECT 147.700 153.800 150.600 154.100 ;
        RECT 146.600 153.600 147.000 153.800 ;
        RECT 146.300 153.100 148.100 153.300 ;
        RECT 148.600 153.100 148.900 153.800 ;
        RECT 151.000 153.100 151.300 154.900 ;
        RECT 151.800 154.800 152.200 154.900 ;
        RECT 153.300 154.200 153.600 155.900 ;
        RECT 154.100 154.900 154.400 155.900 ;
        RECT 153.900 154.500 154.400 154.900 ;
        RECT 153.300 153.800 153.800 154.200 ;
        RECT 144.100 152.800 145.000 153.100 ;
        RECT 146.200 153.000 148.200 153.100 ;
        RECT 144.100 151.100 144.500 152.800 ;
        RECT 146.200 151.100 146.600 153.000 ;
        RECT 147.800 151.100 148.200 153.000 ;
        RECT 148.600 151.100 149.000 153.100 ;
        RECT 151.000 151.100 151.400 153.100 ;
        RECT 151.800 152.800 152.200 153.200 ;
        RECT 153.300 153.100 153.600 153.800 ;
        RECT 154.100 153.700 154.400 154.500 ;
        RECT 154.900 154.800 155.400 155.200 ;
        RECT 154.900 154.400 155.300 154.800 ;
        RECT 154.100 153.400 155.400 153.700 ;
        RECT 155.800 153.400 156.200 154.200 ;
        RECT 153.300 152.800 153.800 153.100 ;
        RECT 151.700 152.400 152.100 152.800 ;
        RECT 153.400 151.100 153.800 152.800 ;
        RECT 155.000 151.100 155.400 153.400 ;
        RECT 156.600 153.100 157.000 159.900 ;
        RECT 158.200 157.100 158.600 157.200 ;
        RECT 159.000 157.100 159.400 159.900 ;
        RECT 158.200 156.800 159.400 157.100 ;
        RECT 157.400 155.800 157.800 156.600 ;
        RECT 157.400 154.100 157.800 154.200 ;
        RECT 158.200 154.100 158.600 154.200 ;
        RECT 157.400 153.800 158.600 154.100 ;
        RECT 158.200 153.400 158.600 153.800 ;
        RECT 159.000 153.100 159.400 156.800 ;
        RECT 159.800 155.800 160.200 156.600 ;
        RECT 160.600 155.600 161.000 159.900 ;
        RECT 162.700 157.900 163.300 159.900 ;
        RECT 165.000 157.900 165.400 159.900 ;
        RECT 167.200 158.200 167.600 159.900 ;
        RECT 167.200 157.900 168.200 158.200 ;
        RECT 163.000 157.500 163.400 157.900 ;
        RECT 165.100 157.600 165.400 157.900 ;
        RECT 164.700 157.300 166.500 157.600 ;
        RECT 167.800 157.500 168.200 157.900 ;
        RECT 164.700 157.200 165.100 157.300 ;
        RECT 166.100 157.200 166.500 157.300 ;
        RECT 162.600 156.600 163.300 157.000 ;
        RECT 163.000 156.100 163.300 156.600 ;
        RECT 164.100 156.500 165.200 156.800 ;
        RECT 164.100 156.400 164.500 156.500 ;
        RECT 163.000 155.800 164.200 156.100 ;
        RECT 160.600 155.300 162.700 155.600 ;
        RECT 160.600 153.600 161.000 155.300 ;
        RECT 162.300 155.200 162.700 155.300 ;
        RECT 161.500 154.900 161.900 155.000 ;
        RECT 161.500 154.600 163.400 154.900 ;
        RECT 163.000 154.500 163.400 154.600 ;
        RECT 163.900 154.200 164.200 155.800 ;
        RECT 164.900 155.900 165.200 156.500 ;
        RECT 165.500 156.500 165.900 156.600 ;
        RECT 167.800 156.500 168.200 156.600 ;
        RECT 165.500 156.200 168.200 156.500 ;
        RECT 164.900 155.700 167.300 155.900 ;
        RECT 169.400 155.700 169.800 159.900 ;
        RECT 170.600 156.800 171.000 157.200 ;
        RECT 170.600 156.200 170.900 156.800 ;
        RECT 171.300 156.200 171.700 159.900 ;
        RECT 173.400 157.500 173.800 159.500 ;
        RECT 170.200 155.900 170.900 156.200 ;
        RECT 170.200 155.800 170.600 155.900 ;
        RECT 171.200 155.800 172.200 156.200 ;
        RECT 173.400 155.800 173.700 157.500 ;
        RECT 175.500 156.400 175.900 159.900 ;
        RECT 175.500 156.100 176.300 156.400 ;
        RECT 164.900 155.600 169.800 155.700 ;
        RECT 166.900 155.500 169.800 155.600 ;
        RECT 167.000 155.400 169.800 155.500 ;
        RECT 166.200 155.100 166.600 155.200 ;
        RECT 166.200 154.800 168.700 155.100 ;
        RECT 167.000 154.700 167.400 154.800 ;
        RECT 168.300 154.700 168.700 154.800 ;
        RECT 167.500 154.200 167.900 154.300 ;
        RECT 171.200 154.200 171.500 155.800 ;
        RECT 173.400 155.500 175.300 155.800 ;
        RECT 171.800 154.400 172.200 155.200 ;
        RECT 173.400 154.400 173.800 155.200 ;
        RECT 174.200 154.400 174.600 155.200 ;
        RECT 175.000 154.500 175.300 155.500 ;
        RECT 163.900 153.900 169.400 154.200 ;
        RECT 164.100 153.800 164.500 153.900 ;
        RECT 160.600 153.300 162.500 153.600 ;
        RECT 156.600 152.800 157.500 153.100 ;
        RECT 159.000 152.800 159.900 153.100 ;
        RECT 157.100 151.100 157.500 152.800 ;
        RECT 159.500 151.100 159.900 152.800 ;
        RECT 160.600 151.100 161.000 153.300 ;
        RECT 162.100 153.200 162.500 153.300 ;
        RECT 167.000 152.800 167.300 153.900 ;
        RECT 168.600 153.800 169.400 153.900 ;
        RECT 170.200 153.800 171.500 154.200 ;
        RECT 172.600 154.100 173.000 154.200 ;
        RECT 172.200 153.800 173.000 154.100 ;
        RECT 175.000 154.100 175.700 154.500 ;
        RECT 176.000 154.200 176.300 156.100 ;
        RECT 176.600 155.100 177.000 155.600 ;
        RECT 178.200 155.100 178.600 155.200 ;
        RECT 176.600 154.800 178.600 155.100 ;
        RECT 175.000 153.900 175.500 154.100 ;
        RECT 166.100 152.700 166.500 152.800 ;
        RECT 163.000 152.100 163.400 152.500 ;
        RECT 165.100 152.400 166.500 152.700 ;
        RECT 167.000 152.400 167.400 152.800 ;
        RECT 165.100 152.100 165.400 152.400 ;
        RECT 167.800 152.100 168.200 152.500 ;
        RECT 162.700 151.800 163.400 152.100 ;
        RECT 162.700 151.100 163.300 151.800 ;
        RECT 165.000 151.100 165.400 152.100 ;
        RECT 167.200 151.800 168.200 152.100 ;
        RECT 167.200 151.100 167.600 151.800 ;
        RECT 169.400 151.100 169.800 153.500 ;
        RECT 170.300 153.100 170.600 153.800 ;
        RECT 172.200 153.600 172.600 153.800 ;
        RECT 173.400 153.600 175.500 153.900 ;
        RECT 176.000 153.800 177.000 154.200 ;
        RECT 171.100 153.100 172.900 153.300 ;
        RECT 170.200 151.100 170.600 153.100 ;
        RECT 171.000 153.000 173.000 153.100 ;
        RECT 171.000 151.100 171.400 153.000 ;
        RECT 172.600 151.100 173.000 153.000 ;
        RECT 173.400 152.500 173.700 153.600 ;
        RECT 176.000 153.500 176.300 153.800 ;
        RECT 175.900 153.300 176.300 153.500 ;
        RECT 178.200 153.400 178.600 154.200 ;
        RECT 175.500 153.000 176.300 153.300 ;
        RECT 179.000 153.100 179.400 159.900 ;
        RECT 179.800 155.800 180.200 156.600 ;
        RECT 181.900 156.200 182.300 159.900 ;
        RECT 182.600 156.800 183.000 157.200 ;
        RECT 182.700 156.200 183.000 156.800 ;
        RECT 181.900 155.900 182.400 156.200 ;
        RECT 182.700 155.900 183.400 156.200 ;
        RECT 181.400 154.400 181.800 155.200 ;
        RECT 182.100 154.200 182.400 155.900 ;
        RECT 183.000 155.800 183.400 155.900 ;
        RECT 183.800 155.800 184.200 156.600 ;
        RECT 183.000 155.100 183.300 155.800 ;
        RECT 184.600 155.100 185.000 159.900 ;
        RECT 185.400 157.100 185.800 157.200 ;
        RECT 186.200 157.100 186.600 159.900 ;
        RECT 188.300 157.900 188.900 159.900 ;
        RECT 190.600 157.900 191.000 159.900 ;
        RECT 192.800 158.200 193.200 159.900 ;
        RECT 192.800 157.900 193.800 158.200 ;
        RECT 188.600 157.500 189.000 157.900 ;
        RECT 190.700 157.600 191.000 157.900 ;
        RECT 190.300 157.300 192.100 157.600 ;
        RECT 193.400 157.500 193.800 157.900 ;
        RECT 190.300 157.200 190.700 157.300 ;
        RECT 191.700 157.200 192.100 157.300 ;
        RECT 185.400 156.800 186.600 157.100 ;
        RECT 183.000 154.800 185.000 155.100 ;
        RECT 179.800 154.100 180.200 154.200 ;
        RECT 180.600 154.100 181.000 154.200 ;
        RECT 179.800 153.800 181.400 154.100 ;
        RECT 182.100 153.800 183.400 154.200 ;
        RECT 181.000 153.600 181.400 153.800 ;
        RECT 180.700 153.100 182.500 153.300 ;
        RECT 183.000 153.100 183.300 153.800 ;
        RECT 184.600 153.100 185.000 154.800 ;
        RECT 186.200 155.600 186.600 156.800 ;
        RECT 188.200 156.600 188.900 157.000 ;
        RECT 188.600 156.100 188.900 156.600 ;
        RECT 189.700 156.500 190.800 156.800 ;
        RECT 189.700 156.400 190.100 156.500 ;
        RECT 188.600 155.800 189.800 156.100 ;
        RECT 186.200 155.300 188.300 155.600 ;
        RECT 185.400 154.100 185.800 154.200 ;
        RECT 186.200 154.100 186.600 155.300 ;
        RECT 187.900 155.200 188.300 155.300 ;
        RECT 187.100 154.900 187.500 155.000 ;
        RECT 187.100 154.600 189.000 154.900 ;
        RECT 188.600 154.500 189.000 154.600 ;
        RECT 185.400 153.800 186.600 154.100 ;
        RECT 189.500 154.200 189.800 155.800 ;
        RECT 190.500 155.900 190.800 156.500 ;
        RECT 191.100 156.500 191.500 156.600 ;
        RECT 193.400 156.500 193.800 156.600 ;
        RECT 191.100 156.200 193.800 156.500 ;
        RECT 190.500 155.700 192.900 155.900 ;
        RECT 195.000 155.700 195.400 159.900 ;
        RECT 190.500 155.600 195.400 155.700 ;
        RECT 192.500 155.500 195.400 155.600 ;
        RECT 192.600 155.400 195.400 155.500 ;
        RECT 190.200 155.100 190.600 155.200 ;
        RECT 191.800 155.100 192.200 155.200 ;
        RECT 190.200 154.800 194.300 155.100 ;
        RECT 193.900 154.700 194.300 154.800 ;
        RECT 193.100 154.200 193.500 154.300 ;
        RECT 189.500 153.900 195.000 154.200 ;
        RECT 189.700 153.800 190.100 153.900 ;
        RECT 185.400 153.400 185.800 153.800 ;
        RECT 186.200 153.600 186.600 153.800 ;
        RECT 173.400 151.500 173.800 152.500 ;
        RECT 175.500 152.200 175.900 153.000 ;
        RECT 179.000 152.800 179.900 153.100 ;
        RECT 175.000 151.800 175.900 152.200 ;
        RECT 175.500 151.500 175.900 151.800 ;
        RECT 179.500 152.200 179.900 152.800 ;
        RECT 180.600 153.000 182.600 153.100 ;
        RECT 179.500 151.800 180.200 152.200 ;
        RECT 179.500 151.100 179.900 151.800 ;
        RECT 180.600 151.100 181.000 153.000 ;
        RECT 182.200 151.100 182.600 153.000 ;
        RECT 183.000 151.100 183.400 153.100 ;
        RECT 184.100 152.800 185.000 153.100 ;
        RECT 186.200 153.300 188.100 153.600 ;
        RECT 184.100 151.100 184.500 152.800 ;
        RECT 186.200 151.100 186.600 153.300 ;
        RECT 187.700 153.200 188.100 153.300 ;
        RECT 192.600 152.800 192.900 153.900 ;
        RECT 194.200 153.800 195.000 153.900 ;
        RECT 191.700 152.700 192.100 152.800 ;
        RECT 188.600 152.100 189.000 152.500 ;
        RECT 190.700 152.400 192.100 152.700 ;
        RECT 192.600 152.400 193.000 152.800 ;
        RECT 190.700 152.100 191.000 152.400 ;
        RECT 193.400 152.100 193.800 152.500 ;
        RECT 188.300 151.800 189.000 152.100 ;
        RECT 188.300 151.100 188.900 151.800 ;
        RECT 190.600 151.100 191.000 152.100 ;
        RECT 192.800 151.800 193.800 152.100 ;
        RECT 192.800 151.100 193.200 151.800 ;
        RECT 195.000 151.100 195.400 153.500 ;
        RECT 197.400 153.400 197.800 154.200 ;
        RECT 198.200 153.100 198.600 159.900 ;
        RECT 199.800 157.500 200.200 159.500 ;
        RECT 201.900 159.200 202.300 159.900 ;
        RECT 201.400 158.800 202.300 159.200 ;
        RECT 199.000 155.800 199.400 157.200 ;
        RECT 199.800 155.800 200.100 157.500 ;
        RECT 201.900 156.400 202.300 158.800 ;
        RECT 205.400 156.400 205.800 159.900 ;
        RECT 201.900 156.100 202.700 156.400 ;
        RECT 199.800 155.500 201.700 155.800 ;
        RECT 199.800 154.400 200.200 155.200 ;
        RECT 200.600 154.400 201.000 155.200 ;
        RECT 201.400 154.500 201.700 155.500 ;
        RECT 201.400 154.100 202.100 154.500 ;
        RECT 202.400 154.200 202.700 156.100 ;
        RECT 205.300 155.900 205.800 156.400 ;
        RECT 207.000 156.200 207.400 159.900 ;
        RECT 206.100 155.900 207.400 156.200 ;
        RECT 209.100 156.200 209.500 159.900 ;
        RECT 209.800 156.800 210.200 157.200 ;
        RECT 209.900 156.200 210.200 156.800 ;
        RECT 209.100 155.900 209.600 156.200 ;
        RECT 209.900 155.900 210.600 156.200 ;
        RECT 203.000 154.800 203.400 155.600 ;
        RECT 205.300 154.200 205.600 155.900 ;
        RECT 206.100 154.900 206.400 155.900 ;
        RECT 205.900 154.500 206.400 154.900 ;
        RECT 201.400 153.900 201.900 154.100 ;
        RECT 199.800 153.600 201.900 153.900 ;
        RECT 202.400 153.800 203.400 154.200 ;
        RECT 204.600 154.100 205.000 154.200 ;
        RECT 205.300 154.100 205.800 154.200 ;
        RECT 204.600 153.800 205.800 154.100 ;
        RECT 198.200 152.800 199.100 153.100 ;
        RECT 198.700 152.200 199.100 152.800 ;
        RECT 198.200 151.800 199.100 152.200 ;
        RECT 198.700 151.100 199.100 151.800 ;
        RECT 199.800 152.500 200.100 153.600 ;
        RECT 202.400 153.500 202.700 153.800 ;
        RECT 202.300 153.300 202.700 153.500 ;
        RECT 201.900 153.000 202.700 153.300 ;
        RECT 205.300 153.100 205.600 153.800 ;
        RECT 206.100 153.700 206.400 154.500 ;
        RECT 206.900 154.800 207.400 155.200 ;
        RECT 206.900 154.400 207.300 154.800 ;
        RECT 208.600 154.400 209.000 155.200 ;
        RECT 209.300 154.200 209.600 155.900 ;
        RECT 210.200 155.800 210.600 155.900 ;
        RECT 211.000 155.800 211.400 156.600 ;
        RECT 210.200 155.100 210.500 155.800 ;
        RECT 211.800 155.100 212.200 159.900 ;
        RECT 213.800 156.800 214.200 157.200 ;
        RECT 213.800 156.200 214.100 156.800 ;
        RECT 214.500 156.200 214.900 159.900 ;
        RECT 213.400 155.900 214.100 156.200 ;
        RECT 214.400 155.900 214.900 156.200 ;
        RECT 213.400 155.800 213.800 155.900 ;
        RECT 210.200 154.800 212.200 155.100 ;
        RECT 213.400 155.100 213.800 155.200 ;
        RECT 214.400 155.100 214.700 155.900 ;
        RECT 216.600 155.600 217.000 159.900 ;
        RECT 218.700 157.900 219.300 159.900 ;
        RECT 221.000 157.900 221.400 159.900 ;
        RECT 223.200 158.200 223.600 159.900 ;
        RECT 223.200 157.900 224.200 158.200 ;
        RECT 219.000 157.500 219.400 157.900 ;
        RECT 221.100 157.600 221.400 157.900 ;
        RECT 220.700 157.300 222.500 157.600 ;
        RECT 223.800 157.500 224.200 157.900 ;
        RECT 220.700 157.200 221.100 157.300 ;
        RECT 222.100 157.200 222.500 157.300 ;
        RECT 218.600 156.600 219.300 157.000 ;
        RECT 219.000 156.100 219.300 156.600 ;
        RECT 220.100 156.500 221.200 156.800 ;
        RECT 220.100 156.400 220.500 156.500 ;
        RECT 219.000 155.800 220.200 156.100 ;
        RECT 216.600 155.300 218.700 155.600 ;
        RECT 213.400 154.800 214.700 155.100 ;
        RECT 207.800 154.100 208.200 154.200 ;
        RECT 207.800 153.800 208.600 154.100 ;
        RECT 209.300 153.800 210.600 154.200 ;
        RECT 206.100 153.400 207.400 153.700 ;
        RECT 208.200 153.600 208.600 153.800 ;
        RECT 199.800 151.500 200.200 152.500 ;
        RECT 201.900 151.500 202.300 153.000 ;
        RECT 205.300 152.800 205.800 153.100 ;
        RECT 205.400 151.100 205.800 152.800 ;
        RECT 207.000 151.100 207.400 153.400 ;
        RECT 207.900 153.100 209.700 153.300 ;
        RECT 210.200 153.100 210.500 153.800 ;
        RECT 211.800 153.100 212.200 154.800 ;
        RECT 214.400 154.200 214.700 154.800 ;
        RECT 215.000 154.400 215.400 155.200 ;
        RECT 212.600 153.400 213.000 154.200 ;
        RECT 213.400 153.800 214.700 154.200 ;
        RECT 215.800 154.100 216.200 154.200 ;
        RECT 215.400 153.800 216.200 154.100 ;
        RECT 213.500 153.100 213.800 153.800 ;
        RECT 215.400 153.600 215.800 153.800 ;
        RECT 216.600 153.600 217.000 155.300 ;
        RECT 218.300 155.200 218.700 155.300 ;
        RECT 217.500 154.900 217.900 155.000 ;
        RECT 217.500 154.600 219.400 154.900 ;
        RECT 219.000 154.500 219.400 154.600 ;
        RECT 219.900 154.200 220.200 155.800 ;
        RECT 220.900 155.900 221.200 156.500 ;
        RECT 221.500 156.500 221.900 156.600 ;
        RECT 223.800 156.500 224.200 156.600 ;
        RECT 221.500 156.200 224.200 156.500 ;
        RECT 220.900 155.700 223.300 155.900 ;
        RECT 225.400 155.700 225.800 159.900 ;
        RECT 226.600 156.800 227.000 157.200 ;
        RECT 226.600 156.200 226.900 156.800 ;
        RECT 227.300 156.200 227.700 159.900 ;
        RECT 226.200 155.900 226.900 156.200 ;
        RECT 227.200 155.900 227.700 156.200 ;
        RECT 226.200 155.800 226.600 155.900 ;
        RECT 220.900 155.600 225.800 155.700 ;
        RECT 222.900 155.500 225.800 155.600 ;
        RECT 223.000 155.400 225.800 155.500 ;
        RECT 222.200 155.100 222.600 155.200 ;
        RECT 222.200 154.800 224.700 155.100 ;
        RECT 224.300 154.700 224.700 154.800 ;
        RECT 223.500 154.200 223.900 154.300 ;
        RECT 227.200 154.200 227.500 155.900 ;
        RECT 227.800 154.400 228.200 155.200 ;
        RECT 219.900 153.900 225.400 154.200 ;
        RECT 220.100 153.800 220.500 153.900 ;
        RECT 216.600 153.300 218.500 153.600 ;
        RECT 214.300 153.100 216.100 153.300 ;
        RECT 207.800 153.000 209.800 153.100 ;
        RECT 207.800 151.100 208.200 153.000 ;
        RECT 209.400 151.100 209.800 153.000 ;
        RECT 210.200 151.100 210.600 153.100 ;
        RECT 211.300 152.800 212.200 153.100 ;
        RECT 211.300 151.100 211.700 152.800 ;
        RECT 213.400 151.100 213.800 153.100 ;
        RECT 214.200 153.000 216.200 153.100 ;
        RECT 214.200 151.100 214.600 153.000 ;
        RECT 215.800 151.100 216.200 153.000 ;
        RECT 216.600 151.100 217.000 153.300 ;
        RECT 218.100 153.200 218.500 153.300 ;
        RECT 223.000 152.800 223.300 153.900 ;
        RECT 224.600 153.800 225.400 153.900 ;
        RECT 226.200 153.800 227.500 154.200 ;
        RECT 228.600 154.100 229.000 154.200 ;
        RECT 230.200 154.100 230.600 154.200 ;
        RECT 228.200 153.800 230.600 154.100 ;
        RECT 222.100 152.700 222.500 152.800 ;
        RECT 219.000 152.100 219.400 152.500 ;
        RECT 221.100 152.400 222.500 152.700 ;
        RECT 223.000 152.400 223.400 152.800 ;
        RECT 221.100 152.100 221.400 152.400 ;
        RECT 223.800 152.100 224.200 152.500 ;
        RECT 218.700 151.800 219.400 152.100 ;
        RECT 218.700 151.100 219.300 151.800 ;
        RECT 221.000 151.100 221.400 152.100 ;
        RECT 223.200 151.800 224.200 152.100 ;
        RECT 223.200 151.100 223.600 151.800 ;
        RECT 225.400 151.100 225.800 153.500 ;
        RECT 226.300 153.100 226.600 153.800 ;
        RECT 228.200 153.600 228.600 153.800 ;
        RECT 227.100 153.100 228.900 153.300 ;
        RECT 226.200 151.100 226.600 153.100 ;
        RECT 227.000 153.000 229.000 153.100 ;
        RECT 227.000 151.100 227.400 153.000 ;
        RECT 228.600 151.100 229.000 153.000 ;
        RECT 0.600 147.500 1.000 149.900 ;
        RECT 2.800 149.200 3.200 149.900 ;
        RECT 2.200 148.900 3.200 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.100 149.200 7.700 149.900 ;
        RECT 7.000 148.900 7.700 149.200 ;
        RECT 2.200 148.500 2.600 148.900 ;
        RECT 5.000 148.600 5.300 148.900 ;
        RECT 3.000 148.200 3.400 148.600 ;
        RECT 3.900 148.300 5.300 148.600 ;
        RECT 7.000 148.500 7.400 148.900 ;
        RECT 3.900 148.200 4.300 148.300 ;
        RECT 1.000 147.100 1.800 147.200 ;
        RECT 3.100 147.100 3.400 148.200 ;
        RECT 7.900 147.700 8.300 147.800 ;
        RECT 9.400 147.700 9.800 149.900 ;
        RECT 10.200 148.000 10.600 149.900 ;
        RECT 11.800 148.000 12.200 149.900 ;
        RECT 10.200 147.900 12.200 148.000 ;
        RECT 12.600 147.900 13.000 149.900 ;
        RECT 13.700 148.200 14.100 149.900 ;
        RECT 17.100 148.200 17.500 149.900 ;
        RECT 18.500 149.200 18.900 149.900 ;
        RECT 18.200 148.800 18.900 149.200 ;
        RECT 13.700 147.900 14.600 148.200 ;
        RECT 10.300 147.700 12.100 147.900 ;
        RECT 7.900 147.400 9.800 147.700 ;
        RECT 4.600 147.100 5.000 147.200 ;
        RECT 5.900 147.100 6.300 147.200 ;
        RECT 1.000 146.800 6.500 147.100 ;
        RECT 2.500 146.700 2.900 146.800 ;
        RECT 1.700 146.200 2.100 146.300 ;
        RECT 1.700 145.900 4.200 146.200 ;
        RECT 3.800 145.800 4.200 145.900 ;
        RECT 0.600 145.500 3.400 145.600 ;
        RECT 0.600 145.400 3.500 145.500 ;
        RECT 0.600 145.300 5.500 145.400 ;
        RECT 0.600 141.100 1.000 145.300 ;
        RECT 3.100 145.100 5.500 145.300 ;
        RECT 2.200 144.500 4.900 144.800 ;
        RECT 2.200 144.400 2.600 144.500 ;
        RECT 4.500 144.400 4.900 144.500 ;
        RECT 5.200 144.500 5.500 145.100 ;
        RECT 6.200 145.200 6.500 146.800 ;
        RECT 7.000 146.400 7.400 146.500 ;
        RECT 7.000 146.100 8.900 146.400 ;
        RECT 8.500 146.000 8.900 146.100 ;
        RECT 7.700 145.700 8.100 145.800 ;
        RECT 9.400 145.700 9.800 147.400 ;
        RECT 10.600 147.200 11.000 147.400 ;
        RECT 12.600 147.200 12.900 147.900 ;
        RECT 10.200 146.900 11.000 147.200 ;
        RECT 10.200 146.800 10.600 146.900 ;
        RECT 11.700 146.800 13.000 147.200 ;
        RECT 11.000 145.800 11.400 146.600 ;
        RECT 11.700 146.200 12.000 146.800 ;
        RECT 11.700 145.800 12.200 146.200 ;
        RECT 14.200 146.100 14.600 147.900 ;
        RECT 16.600 147.900 17.500 148.200 ;
        RECT 18.500 148.200 18.900 148.800 ;
        RECT 18.500 147.900 19.400 148.200 ;
        RECT 20.600 148.000 21.000 149.900 ;
        RECT 22.200 148.000 22.600 149.900 ;
        RECT 20.600 147.900 22.600 148.000 ;
        RECT 23.000 147.900 23.400 149.900 ;
        RECT 15.000 147.100 15.400 147.600 ;
        RECT 15.800 147.100 16.200 147.600 ;
        RECT 15.000 146.800 16.200 147.100 ;
        RECT 12.600 145.800 14.600 146.100 ;
        RECT 7.700 145.400 9.800 145.700 ;
        RECT 6.200 144.900 7.400 145.200 ;
        RECT 5.900 144.500 6.300 144.600 ;
        RECT 5.200 144.200 6.300 144.500 ;
        RECT 7.100 144.400 7.400 144.900 ;
        RECT 7.100 144.000 7.800 144.400 ;
        RECT 3.900 143.700 4.300 143.800 ;
        RECT 5.300 143.700 5.700 143.800 ;
        RECT 2.200 143.100 2.600 143.500 ;
        RECT 3.900 143.400 5.700 143.700 ;
        RECT 5.000 143.100 5.300 143.400 ;
        RECT 7.000 143.100 7.400 143.500 ;
        RECT 2.200 142.800 3.200 143.100 ;
        RECT 2.800 141.100 3.200 142.800 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.100 141.100 7.700 143.100 ;
        RECT 9.400 141.100 9.800 145.400 ;
        RECT 11.700 145.100 12.000 145.800 ;
        RECT 12.600 145.200 12.900 145.800 ;
        RECT 12.600 145.100 13.000 145.200 ;
        RECT 11.500 144.800 12.000 145.100 ;
        RECT 12.300 144.800 13.000 145.100 ;
        RECT 11.500 141.100 11.900 144.800 ;
        RECT 12.300 144.200 12.600 144.800 ;
        RECT 13.400 144.400 13.800 145.200 ;
        RECT 12.200 143.800 12.600 144.200 ;
        RECT 14.200 141.100 14.600 145.800 ;
        RECT 16.600 146.100 17.000 147.900 ;
        RECT 17.400 146.100 17.800 146.200 ;
        RECT 16.600 145.800 17.800 146.100 ;
        RECT 16.600 141.100 17.000 145.800 ;
        RECT 17.400 144.400 17.800 145.200 ;
        RECT 18.200 144.400 18.600 145.200 ;
        RECT 19.000 141.100 19.400 147.900 ;
        RECT 20.700 147.700 22.500 147.900 ;
        RECT 19.800 146.800 20.200 147.600 ;
        RECT 21.000 147.200 21.400 147.400 ;
        RECT 23.000 147.200 23.300 147.900 ;
        RECT 23.800 147.800 24.200 148.600 ;
        RECT 20.600 146.900 21.400 147.200 ;
        RECT 20.600 146.800 21.000 146.900 ;
        RECT 22.100 146.800 23.400 147.200 ;
        RECT 21.400 145.800 21.800 146.600 ;
        RECT 22.100 145.100 22.400 146.800 ;
        RECT 24.600 146.100 25.000 149.900 ;
        RECT 25.400 147.800 25.800 148.600 ;
        RECT 26.200 147.100 26.600 149.900 ;
        RECT 27.000 148.000 27.400 149.900 ;
        RECT 28.600 149.600 30.600 149.900 ;
        RECT 28.600 148.000 29.000 149.600 ;
        RECT 27.000 147.900 29.000 148.000 ;
        RECT 29.400 147.900 29.800 149.300 ;
        RECT 30.200 147.900 30.600 149.600 ;
        RECT 31.000 147.900 31.400 149.900 ;
        RECT 31.800 148.000 32.200 149.900 ;
        RECT 33.400 148.000 33.800 149.900 ;
        RECT 31.800 147.900 33.800 148.000 ;
        RECT 27.100 147.700 28.900 147.900 ;
        RECT 27.400 147.200 27.800 147.400 ;
        RECT 29.500 147.200 29.800 147.900 ;
        RECT 31.100 147.200 31.400 147.900 ;
        RECT 31.900 147.700 33.700 147.900 ;
        RECT 34.200 147.600 34.600 149.900 ;
        RECT 35.800 148.200 36.200 149.900 ;
        RECT 35.800 147.900 36.300 148.200 ;
        RECT 39.000 148.000 39.400 149.900 ;
        RECT 40.600 148.000 41.000 149.900 ;
        RECT 39.000 147.900 41.000 148.000 ;
        RECT 41.400 147.900 41.800 149.900 ;
        RECT 42.200 147.900 42.600 149.900 ;
        RECT 43.000 148.000 43.400 149.900 ;
        RECT 44.600 148.000 45.000 149.900 ;
        RECT 43.000 147.900 45.000 148.000 ;
        RECT 45.400 147.900 45.800 149.900 ;
        RECT 46.200 148.000 46.600 149.900 ;
        RECT 47.800 148.000 48.200 149.900 ;
        RECT 49.400 148.200 49.800 149.900 ;
        RECT 46.200 147.900 48.200 148.000 ;
        RECT 49.300 147.900 49.800 148.200 ;
        RECT 33.000 147.200 33.400 147.400 ;
        RECT 34.200 147.300 35.500 147.600 ;
        RECT 27.000 147.100 27.800 147.200 ;
        RECT 26.200 146.900 27.800 147.100 ;
        RECT 28.600 146.900 29.800 147.200 ;
        RECT 26.200 146.800 27.400 146.900 ;
        RECT 28.600 146.800 29.000 146.900 ;
        RECT 24.600 145.800 25.700 146.100 ;
        RECT 23.000 145.100 23.400 145.200 ;
        RECT 21.900 144.800 22.400 145.100 ;
        RECT 22.700 144.800 23.400 145.100 ;
        RECT 21.900 141.100 22.300 144.800 ;
        RECT 22.700 144.200 23.000 144.800 ;
        RECT 22.600 143.800 23.000 144.200 ;
        RECT 24.600 141.100 25.000 145.800 ;
        RECT 25.400 145.200 25.700 145.800 ;
        RECT 25.400 144.800 25.800 145.200 ;
        RECT 26.200 141.100 26.600 146.800 ;
        RECT 27.800 145.800 28.200 146.600 ;
        RECT 28.600 145.100 28.900 146.800 ;
        RECT 29.400 145.800 29.800 146.600 ;
        RECT 30.200 146.400 30.600 147.200 ;
        RECT 31.000 146.800 32.300 147.200 ;
        RECT 33.000 146.900 33.800 147.200 ;
        RECT 33.400 146.800 33.800 146.900 ;
        RECT 32.000 146.200 32.300 146.800 ;
        RECT 31.800 145.800 32.300 146.200 ;
        RECT 32.600 145.800 33.000 146.600 ;
        RECT 34.300 146.200 34.700 146.600 ;
        RECT 34.200 145.800 34.700 146.200 ;
        RECT 35.200 146.500 35.500 147.300 ;
        RECT 36.000 147.200 36.300 147.900 ;
        RECT 39.100 147.700 40.900 147.900 ;
        RECT 39.400 147.200 39.800 147.400 ;
        RECT 41.400 147.200 41.700 147.900 ;
        RECT 42.300 147.200 42.600 147.900 ;
        RECT 43.100 147.700 44.900 147.900 ;
        RECT 44.200 147.200 44.600 147.400 ;
        RECT 45.500 147.200 45.800 147.900 ;
        RECT 46.300 147.700 48.100 147.900 ;
        RECT 47.400 147.200 47.800 147.400 ;
        RECT 49.300 147.200 49.600 147.900 ;
        RECT 51.000 147.600 51.400 149.900 ;
        RECT 50.100 147.300 51.400 147.600 ;
        RECT 51.800 147.600 52.200 149.900 ;
        RECT 53.400 148.200 53.800 149.900 ;
        RECT 53.400 147.900 53.900 148.200 ;
        RECT 51.800 147.300 53.100 147.600 ;
        RECT 35.800 147.100 36.300 147.200 ;
        RECT 36.600 147.100 37.000 147.200 ;
        RECT 35.800 146.800 37.000 147.100 ;
        RECT 39.000 146.900 39.800 147.200 ;
        RECT 39.000 146.800 39.400 146.900 ;
        RECT 40.500 146.800 41.800 147.200 ;
        RECT 42.200 146.800 43.500 147.200 ;
        RECT 44.200 146.900 45.000 147.200 ;
        RECT 44.600 146.800 45.000 146.900 ;
        RECT 45.400 146.800 46.700 147.200 ;
        RECT 47.400 146.900 48.200 147.200 ;
        RECT 47.800 146.800 48.200 146.900 ;
        RECT 49.300 146.800 49.800 147.200 ;
        RECT 35.200 146.100 35.700 146.500 ;
        RECT 31.000 145.100 31.400 145.200 ;
        RECT 32.000 145.100 32.300 145.800 ;
        RECT 35.200 145.100 35.500 146.100 ;
        RECT 36.000 145.100 36.300 146.800 ;
        RECT 39.800 145.800 40.200 146.600 ;
        RECT 40.500 145.100 40.800 146.800 ;
        RECT 41.400 145.100 41.800 145.200 ;
        RECT 28.300 144.200 29.300 145.100 ;
        RECT 31.000 144.800 31.700 145.100 ;
        RECT 32.000 144.800 32.500 145.100 ;
        RECT 31.400 144.200 31.700 144.800 ;
        RECT 28.300 143.800 29.800 144.200 ;
        RECT 31.400 143.800 31.800 144.200 ;
        RECT 28.300 141.100 29.300 143.800 ;
        RECT 32.100 141.100 32.500 144.800 ;
        RECT 34.200 144.800 35.500 145.100 ;
        RECT 34.200 141.100 34.600 144.800 ;
        RECT 35.800 144.600 36.300 145.100 ;
        RECT 40.300 144.800 40.800 145.100 ;
        RECT 41.100 144.800 41.800 145.100 ;
        RECT 42.200 145.100 42.600 145.200 ;
        RECT 43.200 145.100 43.500 146.800 ;
        RECT 43.800 145.800 44.200 146.600 ;
        RECT 44.600 146.100 45.000 146.200 ;
        RECT 45.400 146.100 45.700 146.800 ;
        RECT 44.600 145.800 45.700 146.100 ;
        RECT 45.400 145.100 45.800 145.200 ;
        RECT 46.400 145.100 46.700 146.800 ;
        RECT 47.000 145.800 47.400 146.600 ;
        RECT 49.300 145.100 49.600 146.800 ;
        RECT 50.100 146.500 50.400 147.300 ;
        RECT 49.900 146.100 50.400 146.500 ;
        RECT 50.100 145.100 50.400 146.100 ;
        RECT 50.900 146.200 51.300 146.600 ;
        RECT 51.900 146.200 52.300 146.600 ;
        RECT 50.900 146.100 51.400 146.200 ;
        RECT 51.800 146.100 52.300 146.200 ;
        RECT 50.900 145.800 52.300 146.100 ;
        RECT 52.800 146.500 53.100 147.300 ;
        RECT 53.600 147.200 53.900 147.900 ;
        RECT 55.000 147.500 55.400 149.900 ;
        RECT 57.200 149.200 57.600 149.900 ;
        RECT 56.600 148.900 57.600 149.200 ;
        RECT 59.400 148.900 59.800 149.900 ;
        RECT 61.500 149.200 62.100 149.900 ;
        RECT 61.400 148.900 62.100 149.200 ;
        RECT 56.600 148.500 57.000 148.900 ;
        RECT 59.400 148.600 59.700 148.900 ;
        RECT 57.400 148.200 57.800 148.600 ;
        RECT 58.300 148.300 59.700 148.600 ;
        RECT 61.400 148.500 61.800 148.900 ;
        RECT 58.300 148.200 58.700 148.300 ;
        RECT 57.500 147.200 57.800 148.200 ;
        RECT 62.300 147.700 62.700 147.800 ;
        RECT 63.800 147.700 64.200 149.900 ;
        RECT 64.600 148.000 65.000 149.900 ;
        RECT 66.200 148.000 66.600 149.900 ;
        RECT 64.600 147.900 66.600 148.000 ;
        RECT 67.000 147.900 67.400 149.900 ;
        RECT 67.800 147.900 68.200 149.900 ;
        RECT 68.600 148.000 69.000 149.900 ;
        RECT 70.200 148.000 70.600 149.900 ;
        RECT 68.600 147.900 70.600 148.000 ;
        RECT 71.000 148.000 71.400 149.900 ;
        RECT 72.600 148.000 73.000 149.900 ;
        RECT 71.000 147.900 73.000 148.000 ;
        RECT 73.400 147.900 73.800 149.900 ;
        RECT 74.200 148.500 74.600 149.500 ;
        RECT 64.700 147.700 66.500 147.900 ;
        RECT 62.300 147.400 64.200 147.700 ;
        RECT 53.400 146.800 53.900 147.200 ;
        RECT 55.400 147.100 56.200 147.200 ;
        RECT 57.400 147.100 57.800 147.200 ;
        RECT 58.200 147.100 58.600 147.200 ;
        RECT 60.300 147.100 60.700 147.200 ;
        RECT 55.400 146.800 60.900 147.100 ;
        RECT 52.800 146.100 53.300 146.500 ;
        RECT 52.800 145.100 53.100 146.100 ;
        RECT 53.600 145.100 53.900 146.800 ;
        RECT 56.900 146.700 57.300 146.800 ;
        RECT 56.100 146.200 56.500 146.300 ;
        RECT 56.100 146.100 58.600 146.200 ;
        RECT 59.000 146.100 59.400 146.200 ;
        RECT 56.100 145.900 59.400 146.100 ;
        RECT 58.200 145.800 59.400 145.900 ;
        RECT 42.200 144.800 42.900 145.100 ;
        RECT 43.200 144.800 43.700 145.100 ;
        RECT 45.400 144.800 46.100 145.100 ;
        RECT 46.400 144.800 46.900 145.100 ;
        RECT 35.800 141.100 36.200 144.600 ;
        RECT 40.300 142.200 40.700 144.800 ;
        RECT 41.100 144.200 41.400 144.800 ;
        RECT 41.000 143.800 41.400 144.200 ;
        RECT 42.600 144.200 42.900 144.800 ;
        RECT 42.600 143.800 43.000 144.200 ;
        RECT 39.800 141.800 40.700 142.200 ;
        RECT 40.300 141.100 40.700 141.800 ;
        RECT 43.300 141.100 43.700 144.800 ;
        RECT 45.800 144.200 46.100 144.800 ;
        RECT 45.800 143.800 46.200 144.200 ;
        RECT 46.500 141.100 46.900 144.800 ;
        RECT 49.300 144.600 49.800 145.100 ;
        RECT 50.100 144.800 51.400 145.100 ;
        RECT 49.400 141.100 49.800 144.600 ;
        RECT 51.000 141.100 51.400 144.800 ;
        RECT 51.800 144.800 53.100 145.100 ;
        RECT 51.800 141.100 52.200 144.800 ;
        RECT 53.400 144.600 53.900 145.100 ;
        RECT 55.000 145.500 57.800 145.600 ;
        RECT 55.000 145.400 57.900 145.500 ;
        RECT 55.000 145.300 59.900 145.400 ;
        RECT 53.400 141.100 53.800 144.600 ;
        RECT 55.000 141.100 55.400 145.300 ;
        RECT 57.500 145.100 59.900 145.300 ;
        RECT 56.600 144.500 59.300 144.800 ;
        RECT 56.600 144.400 57.000 144.500 ;
        RECT 58.900 144.400 59.300 144.500 ;
        RECT 59.600 144.500 59.900 145.100 ;
        RECT 60.600 145.200 60.900 146.800 ;
        RECT 61.400 146.400 61.800 146.500 ;
        RECT 61.400 146.100 63.300 146.400 ;
        RECT 62.900 146.000 63.300 146.100 ;
        RECT 62.100 145.700 62.500 145.800 ;
        RECT 63.800 145.700 64.200 147.400 ;
        RECT 65.000 147.200 65.400 147.400 ;
        RECT 67.000 147.200 67.300 147.900 ;
        RECT 67.900 147.200 68.200 147.900 ;
        RECT 68.700 147.700 70.500 147.900 ;
        RECT 71.100 147.700 72.900 147.900 ;
        RECT 69.800 147.200 70.200 147.400 ;
        RECT 71.400 147.200 71.800 147.400 ;
        RECT 73.400 147.200 73.700 147.900 ;
        RECT 74.200 147.400 74.500 148.500 ;
        RECT 76.300 148.000 76.700 149.500 ;
        RECT 76.300 147.700 77.100 148.000 ;
        RECT 76.700 147.500 77.100 147.700 ;
        RECT 64.600 146.900 65.400 147.200 ;
        RECT 64.600 146.800 65.000 146.900 ;
        RECT 66.100 146.800 67.400 147.200 ;
        RECT 67.800 146.800 69.100 147.200 ;
        RECT 69.800 147.100 70.600 147.200 ;
        RECT 71.000 147.100 71.800 147.200 ;
        RECT 69.800 146.900 71.800 147.100 ;
        RECT 70.200 146.800 71.400 146.900 ;
        RECT 72.500 146.800 73.800 147.200 ;
        RECT 74.200 147.100 76.300 147.400 ;
        RECT 75.800 146.900 76.300 147.100 ;
        RECT 76.800 147.200 77.100 147.500 ;
        RECT 65.400 145.800 65.800 146.600 ;
        RECT 66.100 146.200 66.400 146.800 ;
        RECT 66.100 145.800 66.600 146.200 ;
        RECT 68.800 146.100 69.100 146.800 ;
        RECT 67.000 145.800 69.100 146.100 ;
        RECT 69.400 146.100 69.800 146.600 ;
        RECT 71.800 146.100 72.200 146.600 ;
        RECT 69.400 145.800 72.200 146.100 ;
        RECT 62.100 145.400 64.200 145.700 ;
        RECT 60.600 144.900 61.800 145.200 ;
        RECT 60.300 144.500 60.700 144.600 ;
        RECT 59.600 144.200 60.700 144.500 ;
        RECT 61.500 144.400 61.800 144.900 ;
        RECT 61.500 144.000 62.200 144.400 ;
        RECT 58.300 143.700 58.700 143.800 ;
        RECT 59.700 143.700 60.100 143.800 ;
        RECT 56.600 143.100 57.000 143.500 ;
        RECT 58.300 143.400 60.100 143.700 ;
        RECT 59.400 143.100 59.700 143.400 ;
        RECT 61.400 143.100 61.800 143.500 ;
        RECT 56.600 142.800 57.600 143.100 ;
        RECT 57.200 141.100 57.600 142.800 ;
        RECT 59.400 141.100 59.800 143.100 ;
        RECT 61.500 141.100 62.100 143.100 ;
        RECT 63.800 141.100 64.200 145.400 ;
        RECT 66.100 145.100 66.400 145.800 ;
        RECT 67.000 145.200 67.300 145.800 ;
        RECT 67.000 145.100 67.400 145.200 ;
        RECT 65.900 144.800 66.400 145.100 ;
        RECT 66.700 144.800 67.400 145.100 ;
        RECT 67.800 145.100 68.200 145.200 ;
        RECT 68.800 145.100 69.100 145.800 ;
        RECT 72.500 145.100 72.800 146.800 ;
        RECT 74.200 145.800 74.600 146.600 ;
        RECT 75.000 145.800 75.400 146.600 ;
        RECT 75.800 146.500 76.500 146.900 ;
        RECT 76.800 146.800 77.800 147.200 ;
        RECT 79.000 146.800 79.400 147.600 ;
        RECT 75.800 145.500 76.100 146.500 ;
        RECT 74.200 145.200 76.100 145.500 ;
        RECT 73.400 145.100 73.800 145.200 ;
        RECT 67.800 144.800 68.500 145.100 ;
        RECT 68.800 144.800 69.300 145.100 ;
        RECT 65.900 141.100 66.300 144.800 ;
        RECT 66.700 144.200 67.000 144.800 ;
        RECT 66.600 143.800 67.000 144.200 ;
        RECT 68.200 144.200 68.500 144.800 ;
        RECT 68.200 143.800 68.600 144.200 ;
        RECT 68.900 141.100 69.300 144.800 ;
        RECT 72.300 144.800 72.800 145.100 ;
        RECT 73.100 144.800 73.800 145.100 ;
        RECT 72.300 142.200 72.700 144.800 ;
        RECT 73.100 144.200 73.400 144.800 ;
        RECT 73.000 143.800 73.400 144.200 ;
        RECT 71.800 141.800 72.700 142.200 ;
        RECT 72.300 141.100 72.700 141.800 ;
        RECT 74.200 143.500 74.500 145.200 ;
        RECT 76.800 144.900 77.100 146.800 ;
        RECT 77.400 146.100 77.800 146.200 ;
        RECT 78.200 146.100 78.600 146.200 ;
        RECT 77.400 145.800 78.600 146.100 ;
        RECT 79.800 146.100 80.200 149.900 ;
        RECT 82.200 148.900 82.600 149.900 ;
        RECT 81.400 147.800 81.800 148.600 ;
        RECT 82.300 147.800 82.600 148.900 ;
        RECT 83.800 147.900 84.200 149.900 ;
        RECT 84.600 147.900 85.000 149.900 ;
        RECT 85.400 148.000 85.800 149.900 ;
        RECT 87.000 148.000 87.400 149.900 ;
        RECT 85.400 147.900 87.400 148.000 ;
        RECT 90.000 149.100 90.400 149.900 ;
        RECT 91.000 149.100 91.400 149.200 ;
        RECT 90.000 148.800 91.400 149.100 ;
        RECT 82.300 147.500 83.500 147.800 ;
        RECT 82.200 146.800 82.700 147.200 ;
        RECT 82.400 146.400 82.800 146.800 ;
        RECT 80.600 146.100 81.000 146.200 ;
        RECT 79.800 145.800 81.000 146.100 ;
        RECT 83.200 146.000 83.500 147.500 ;
        RECT 83.900 146.200 84.200 147.900 ;
        RECT 84.700 147.200 85.000 147.900 ;
        RECT 85.500 147.700 87.300 147.900 ;
        RECT 86.600 147.200 87.000 147.400 ;
        RECT 84.600 146.800 85.900 147.200 ;
        RECT 86.600 146.900 87.400 147.200 ;
        RECT 90.000 147.100 90.400 148.800 ;
        RECT 87.000 146.800 87.400 146.900 ;
        RECT 89.500 146.900 90.400 147.100 ;
        RECT 94.400 147.100 94.800 149.900 ;
        RECT 94.400 146.900 95.300 147.100 ;
        RECT 89.500 146.800 90.300 146.900 ;
        RECT 94.500 146.800 95.300 146.900 ;
        RECT 95.800 146.800 96.200 147.600 ;
        RECT 77.400 145.400 77.800 145.800 ;
        RECT 76.300 144.600 77.100 144.900 ;
        RECT 74.200 141.500 74.600 143.500 ;
        RECT 76.300 141.100 76.700 144.600 ;
        RECT 79.800 141.100 80.200 145.800 ;
        RECT 83.100 145.700 83.500 146.000 ;
        RECT 83.800 145.800 84.200 146.200 ;
        RECT 81.400 145.600 83.500 145.700 ;
        RECT 81.400 145.400 83.400 145.600 ;
        RECT 81.400 141.100 81.800 145.400 ;
        RECT 83.900 145.100 84.200 145.800 ;
        RECT 83.500 144.800 84.200 145.100 ;
        RECT 84.600 145.100 85.000 145.200 ;
        RECT 85.600 145.100 85.900 146.800 ;
        RECT 86.200 145.800 86.600 146.600 ;
        RECT 89.500 145.200 89.800 146.800 ;
        RECT 90.600 145.800 91.400 146.200 ;
        RECT 93.400 145.800 94.200 146.200 ;
        RECT 84.600 144.800 85.300 145.100 ;
        RECT 85.600 144.800 86.100 145.100 ;
        RECT 89.400 144.800 89.800 145.200 ;
        RECT 91.800 145.100 92.200 145.600 ;
        RECT 92.600 145.100 93.000 145.600 ;
        RECT 91.800 144.800 93.000 145.100 ;
        RECT 95.000 145.200 95.300 146.800 ;
        RECT 95.000 144.800 95.400 145.200 ;
        RECT 83.500 144.200 83.900 144.800 ;
        RECT 85.000 144.200 85.300 144.800 ;
        RECT 83.500 143.800 84.200 144.200 ;
        RECT 85.000 143.800 85.400 144.200 ;
        RECT 83.500 141.100 83.900 143.800 ;
        RECT 85.700 141.100 86.100 144.800 ;
        RECT 89.500 143.500 89.800 144.800 ;
        RECT 90.200 144.100 90.600 144.600 ;
        RECT 91.800 144.100 92.200 144.200 ;
        RECT 90.200 143.800 92.200 144.100 ;
        RECT 94.200 143.800 94.600 144.600 ;
        RECT 95.000 143.500 95.300 144.800 ;
        RECT 89.500 143.200 91.300 143.500 ;
        RECT 89.500 143.100 89.800 143.200 ;
        RECT 89.400 141.100 89.800 143.100 ;
        RECT 91.000 143.100 91.300 143.200 ;
        RECT 93.500 143.200 95.300 143.500 ;
        RECT 93.500 143.100 93.800 143.200 ;
        RECT 91.000 141.100 91.400 143.100 ;
        RECT 93.400 141.100 93.800 143.100 ;
        RECT 95.000 143.100 95.300 143.200 ;
        RECT 95.000 141.100 95.400 143.100 ;
        RECT 96.600 141.100 97.000 149.900 ;
        RECT 100.000 149.200 100.400 149.900 ;
        RECT 100.000 148.800 101.000 149.200 ;
        RECT 102.200 148.900 102.600 149.900 ;
        RECT 105.600 149.200 106.000 149.900 ;
        RECT 100.000 147.100 100.400 148.800 ;
        RECT 102.200 147.200 102.500 148.900 ;
        RECT 105.600 148.800 106.600 149.200 ;
        RECT 103.000 147.800 103.400 148.600 ;
        RECT 100.000 146.900 100.900 147.100 ;
        RECT 100.100 146.800 100.900 146.900 ;
        RECT 99.000 145.800 99.800 146.200 ;
        RECT 98.200 145.100 98.600 145.600 ;
        RECT 100.600 145.200 100.900 146.800 ;
        RECT 102.200 146.800 102.600 147.200 ;
        RECT 105.600 147.100 106.000 148.800 ;
        RECT 107.800 148.200 108.200 149.900 ;
        RECT 107.700 147.900 108.200 148.200 ;
        RECT 107.700 147.200 108.000 147.900 ;
        RECT 109.400 147.600 109.800 149.900 ;
        RECT 111.000 148.900 111.400 149.900 ;
        RECT 110.200 147.800 110.600 148.600 ;
        RECT 108.500 147.300 109.800 147.600 ;
        RECT 107.000 147.100 107.400 147.200 ;
        RECT 107.700 147.100 108.200 147.200 ;
        RECT 105.600 146.900 106.500 147.100 ;
        RECT 105.700 146.800 106.500 146.900 ;
        RECT 107.000 146.800 108.200 147.100 ;
        RECT 101.400 145.400 101.800 146.200 ;
        RECT 102.200 145.200 102.500 146.800 ;
        RECT 104.600 145.800 105.400 146.200 ;
        RECT 99.000 145.100 99.400 145.200 ;
        RECT 98.200 144.800 99.400 145.100 ;
        RECT 100.600 144.800 101.000 145.200 ;
        RECT 102.200 145.100 102.600 145.200 ;
        RECT 99.800 143.800 100.200 144.600 ;
        RECT 100.600 143.500 100.900 144.800 ;
        RECT 99.100 143.200 100.900 143.500 ;
        RECT 99.100 143.100 99.400 143.200 ;
        RECT 99.000 141.100 99.400 143.100 ;
        RECT 100.600 143.100 100.900 143.200 ;
        RECT 101.700 144.700 102.600 145.100 ;
        RECT 103.800 145.100 104.200 145.600 ;
        RECT 106.200 145.200 106.500 146.800 ;
        RECT 104.600 145.100 105.000 145.200 ;
        RECT 103.800 144.800 105.000 145.100 ;
        RECT 106.200 144.800 106.600 145.200 ;
        RECT 107.700 145.100 108.000 146.800 ;
        RECT 108.500 146.500 108.800 147.300 ;
        RECT 111.100 147.200 111.400 148.900 ;
        RECT 111.000 146.800 111.400 147.200 ;
        RECT 108.300 146.100 108.800 146.500 ;
        RECT 108.500 145.100 108.800 146.100 ;
        RECT 109.300 146.200 109.700 146.600 ;
        RECT 109.300 145.800 109.800 146.200 ;
        RECT 111.100 145.100 111.400 146.800 ;
        RECT 113.400 148.800 113.800 149.900 ;
        RECT 113.400 147.200 113.700 148.800 ;
        RECT 114.200 147.800 114.600 148.600 ;
        RECT 115.000 147.900 115.400 149.900 ;
        RECT 116.600 148.900 117.000 149.900 ;
        RECT 113.400 146.800 113.800 147.200 ;
        RECT 111.800 146.100 112.200 146.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 111.800 145.800 113.000 146.100 ;
        RECT 111.800 145.400 112.200 145.800 ;
        RECT 112.600 145.400 113.000 145.800 ;
        RECT 113.400 145.200 113.700 146.800 ;
        RECT 115.000 146.200 115.300 147.900 ;
        RECT 116.600 147.800 116.900 148.900 ;
        RECT 117.400 147.800 117.800 148.600 ;
        RECT 118.200 148.000 118.600 149.900 ;
        RECT 119.800 148.000 120.200 149.900 ;
        RECT 118.200 147.900 120.200 148.000 ;
        RECT 120.600 147.900 121.000 149.900 ;
        RECT 121.700 148.200 122.100 149.900 ;
        RECT 124.100 149.200 124.500 149.900 ;
        RECT 123.800 148.800 124.500 149.200 ;
        RECT 124.100 148.200 124.500 148.800 ;
        RECT 126.500 148.200 126.900 149.900 ;
        RECT 121.700 147.900 122.600 148.200 ;
        RECT 124.100 147.900 125.000 148.200 ;
        RECT 126.500 147.900 127.400 148.200 ;
        RECT 128.600 148.000 129.000 149.900 ;
        RECT 130.200 148.000 130.600 149.900 ;
        RECT 128.600 147.900 130.600 148.000 ;
        RECT 131.000 147.900 131.400 149.900 ;
        RECT 115.700 147.500 116.900 147.800 ;
        RECT 118.300 147.700 120.100 147.900 ;
        RECT 114.200 146.100 114.600 146.200 ;
        RECT 115.000 146.100 115.400 146.200 ;
        RECT 114.200 145.800 115.400 146.100 ;
        RECT 115.700 146.000 116.000 147.500 ;
        RECT 118.600 147.200 119.000 147.400 ;
        RECT 120.600 147.200 120.900 147.900 ;
        RECT 116.500 146.800 117.000 147.200 ;
        RECT 118.200 146.900 119.000 147.200 ;
        RECT 118.200 146.800 118.600 146.900 ;
        RECT 119.700 146.800 121.000 147.200 ;
        RECT 116.400 146.400 116.800 146.800 ;
        RECT 113.400 145.100 113.800 145.200 ;
        RECT 100.600 141.100 101.000 143.100 ;
        RECT 101.700 141.100 102.100 144.700 ;
        RECT 105.400 143.800 105.800 144.600 ;
        RECT 106.200 143.500 106.500 144.800 ;
        RECT 107.700 144.600 108.200 145.100 ;
        RECT 108.500 144.800 109.800 145.100 ;
        RECT 104.700 143.200 106.500 143.500 ;
        RECT 104.700 143.100 105.000 143.200 ;
        RECT 104.600 141.100 105.000 143.100 ;
        RECT 106.200 143.100 106.500 143.200 ;
        RECT 106.200 141.100 106.600 143.100 ;
        RECT 107.800 141.100 108.200 144.600 ;
        RECT 109.400 141.100 109.800 144.800 ;
        RECT 111.000 144.700 111.900 145.100 ;
        RECT 111.500 143.200 111.900 144.700 ;
        RECT 112.900 144.700 113.800 145.100 ;
        RECT 115.000 145.100 115.300 145.800 ;
        RECT 115.700 145.700 116.100 146.000 ;
        RECT 119.000 145.800 119.400 146.600 ;
        RECT 115.700 145.600 117.800 145.700 ;
        RECT 115.800 145.400 117.800 145.600 ;
        RECT 115.000 144.800 115.700 145.100 ;
        RECT 111.500 142.800 112.200 143.200 ;
        RECT 111.500 141.100 111.900 142.800 ;
        RECT 112.900 141.100 113.300 144.700 ;
        RECT 115.300 141.100 115.700 144.800 ;
        RECT 117.400 141.100 117.800 145.400 ;
        RECT 119.700 145.100 120.000 146.800 ;
        RECT 122.200 146.100 122.600 147.900 ;
        RECT 123.000 146.800 123.400 147.600 ;
        RECT 120.600 145.800 122.600 146.100 ;
        RECT 120.600 145.200 120.900 145.800 ;
        RECT 120.600 145.100 121.000 145.200 ;
        RECT 119.500 144.800 120.000 145.100 ;
        RECT 120.300 144.800 121.000 145.100 ;
        RECT 119.500 141.100 119.900 144.800 ;
        RECT 120.300 144.200 120.600 144.800 ;
        RECT 121.400 144.400 121.800 145.200 ;
        RECT 120.200 143.800 120.600 144.200 ;
        RECT 122.200 141.100 122.600 145.800 ;
        RECT 123.800 144.400 124.200 145.200 ;
        RECT 124.600 141.100 125.000 147.900 ;
        RECT 125.400 146.800 125.800 147.600 ;
        RECT 126.200 144.400 126.600 145.200 ;
        RECT 127.000 145.100 127.400 147.900 ;
        RECT 128.700 147.700 130.500 147.900 ;
        RECT 127.800 146.800 128.200 147.600 ;
        RECT 129.000 147.200 129.400 147.400 ;
        RECT 131.000 147.200 131.300 147.900 ;
        RECT 131.800 147.800 132.200 148.600 ;
        RECT 131.800 147.200 132.100 147.800 ;
        RECT 128.600 146.900 129.400 147.200 ;
        RECT 128.600 146.800 129.000 146.900 ;
        RECT 130.100 146.800 131.400 147.200 ;
        RECT 131.800 146.800 132.200 147.200 ;
        RECT 127.800 145.800 128.200 146.200 ;
        RECT 129.400 145.800 129.800 146.600 ;
        RECT 130.100 146.100 130.400 146.800 ;
        RECT 131.800 146.100 132.200 146.200 ;
        RECT 130.100 145.800 132.200 146.100 ;
        RECT 127.800 145.100 128.100 145.800 ;
        RECT 130.100 145.100 130.400 145.800 ;
        RECT 131.000 145.100 131.400 145.200 ;
        RECT 127.000 144.800 128.100 145.100 ;
        RECT 129.900 144.800 130.400 145.100 ;
        RECT 130.700 144.800 131.400 145.100 ;
        RECT 127.000 141.100 127.400 144.800 ;
        RECT 129.900 141.100 130.300 144.800 ;
        RECT 130.700 144.200 131.000 144.800 ;
        RECT 130.600 143.800 131.000 144.200 ;
        RECT 132.600 141.100 133.000 149.900 ;
        RECT 133.400 147.900 133.800 149.900 ;
        RECT 134.200 148.000 134.600 149.900 ;
        RECT 135.800 148.000 136.200 149.900 ;
        RECT 136.900 148.200 137.300 149.900 ;
        RECT 134.200 147.900 136.200 148.000 ;
        RECT 133.500 147.200 133.800 147.900 ;
        RECT 134.300 147.700 136.100 147.900 ;
        RECT 136.600 147.800 137.800 148.200 ;
        RECT 140.600 148.000 141.000 149.900 ;
        RECT 142.200 148.000 142.600 149.900 ;
        RECT 140.600 147.900 142.600 148.000 ;
        RECT 143.000 147.900 143.400 149.900 ;
        RECT 144.100 148.200 144.500 149.900 ;
        RECT 144.100 147.900 145.000 148.200 ;
        RECT 147.700 147.900 148.500 149.900 ;
        RECT 135.400 147.200 135.800 147.400 ;
        RECT 136.600 147.200 136.900 147.800 ;
        RECT 133.400 146.800 134.700 147.200 ;
        RECT 135.400 146.900 136.200 147.200 ;
        RECT 135.800 146.800 136.200 146.900 ;
        RECT 136.600 146.800 137.000 147.200 ;
        RECT 133.400 145.100 133.800 145.200 ;
        RECT 134.400 145.100 134.700 146.800 ;
        RECT 135.000 146.100 135.400 146.600 ;
        RECT 135.800 146.100 136.200 146.200 ;
        RECT 135.000 145.800 136.200 146.100 ;
        RECT 133.400 144.800 134.100 145.100 ;
        RECT 134.400 144.800 134.900 145.100 ;
        RECT 133.800 144.200 134.100 144.800 ;
        RECT 133.800 143.800 134.200 144.200 ;
        RECT 134.500 141.100 134.900 144.800 ;
        RECT 136.600 144.400 137.000 145.200 ;
        RECT 137.400 141.100 137.800 147.800 ;
        RECT 140.700 147.700 142.500 147.900 ;
        RECT 138.200 147.100 138.600 147.600 ;
        RECT 141.000 147.200 141.400 147.400 ;
        RECT 143.000 147.200 143.300 147.900 ;
        RECT 139.000 147.100 139.400 147.200 ;
        RECT 138.200 146.800 139.400 147.100 ;
        RECT 140.600 146.900 141.400 147.200 ;
        RECT 140.600 146.800 141.000 146.900 ;
        RECT 142.100 146.800 143.400 147.200 ;
        RECT 141.400 145.800 141.800 146.600 ;
        RECT 142.100 145.100 142.400 146.800 ;
        RECT 144.600 146.100 145.000 147.900 ;
        RECT 145.400 146.800 145.800 147.600 ;
        RECT 147.900 147.200 148.200 147.900 ;
        RECT 147.000 146.400 147.400 147.200 ;
        RECT 147.800 146.800 148.200 147.200 ;
        RECT 147.900 146.200 148.200 146.800 ;
        RECT 148.600 146.800 149.000 147.200 ;
        RECT 152.000 147.100 152.400 149.900 ;
        RECT 152.000 146.900 152.900 147.100 ;
        RECT 152.100 146.800 152.900 146.900 ;
        RECT 148.600 146.600 148.900 146.800 ;
        RECT 148.500 146.200 148.900 146.600 ;
        RECT 143.000 145.800 145.000 146.100 ;
        RECT 145.400 146.100 145.800 146.200 ;
        RECT 146.200 146.100 146.600 146.200 ;
        RECT 145.400 145.800 147.000 146.100 ;
        RECT 147.800 145.800 148.200 146.200 ;
        RECT 143.000 145.200 143.300 145.800 ;
        RECT 143.000 145.100 143.400 145.200 ;
        RECT 141.900 144.800 142.400 145.100 ;
        RECT 142.700 144.800 143.400 145.100 ;
        RECT 141.900 141.100 142.300 144.800 ;
        RECT 142.700 144.200 143.000 144.800 ;
        RECT 143.800 144.400 144.200 145.200 ;
        RECT 142.600 143.800 143.000 144.200 ;
        RECT 144.600 141.100 145.000 145.800 ;
        RECT 146.600 145.600 147.000 145.800 ;
        RECT 147.900 145.700 148.200 145.800 ;
        RECT 147.900 145.400 148.900 145.700 ;
        RECT 149.400 145.400 149.800 146.200 ;
        RECT 151.000 145.800 151.800 146.200 ;
        RECT 148.600 145.100 148.900 145.400 ;
        RECT 146.200 144.800 148.200 145.100 ;
        RECT 146.200 141.100 146.600 144.800 ;
        RECT 147.800 141.400 148.200 144.800 ;
        RECT 148.600 141.700 149.000 145.100 ;
        RECT 149.400 141.400 149.800 145.100 ;
        RECT 150.200 144.800 150.600 145.600 ;
        RECT 152.600 145.200 152.900 146.800 ;
        RECT 152.600 144.800 153.000 145.200 ;
        RECT 151.800 143.800 152.200 144.600 ;
        RECT 152.600 143.500 152.900 144.800 ;
        RECT 151.100 143.200 152.900 143.500 ;
        RECT 151.100 143.100 151.400 143.200 ;
        RECT 147.800 141.100 149.800 141.400 ;
        RECT 151.000 141.100 151.400 143.100 ;
        RECT 152.600 143.100 152.900 143.200 ;
        RECT 153.400 144.100 153.800 149.900 ;
        RECT 154.200 147.800 154.600 148.600 ;
        RECT 156.900 148.000 157.300 149.500 ;
        RECT 159.000 148.500 159.400 149.500 ;
        RECT 156.500 147.700 157.300 148.000 ;
        RECT 156.500 147.500 156.900 147.700 ;
        RECT 156.500 147.200 156.800 147.500 ;
        RECT 159.100 147.400 159.400 148.500 ;
        RECT 161.700 148.000 162.100 149.500 ;
        RECT 163.800 148.500 164.200 149.500 ;
        RECT 155.800 146.800 156.800 147.200 ;
        RECT 157.300 147.100 159.400 147.400 ;
        RECT 161.300 147.700 162.100 148.000 ;
        RECT 161.300 147.500 161.700 147.700 ;
        RECT 161.300 147.200 161.600 147.500 ;
        RECT 163.900 147.400 164.200 148.500 ;
        RECT 157.300 146.900 157.800 147.100 ;
        RECT 156.500 146.200 156.800 146.800 ;
        RECT 157.100 146.500 157.800 146.900 ;
        RECT 160.600 146.800 161.600 147.200 ;
        RECT 162.100 147.100 164.200 147.400 ;
        RECT 164.600 147.700 165.000 149.900 ;
        RECT 166.700 149.200 167.300 149.900 ;
        RECT 166.700 148.900 167.400 149.200 ;
        RECT 169.000 148.900 169.400 149.900 ;
        RECT 171.200 149.200 171.600 149.900 ;
        RECT 171.200 148.900 172.200 149.200 ;
        RECT 167.000 148.500 167.400 148.900 ;
        RECT 169.100 148.600 169.400 148.900 ;
        RECT 169.100 148.300 170.500 148.600 ;
        RECT 170.100 148.200 170.500 148.300 ;
        RECT 171.000 148.200 171.400 148.600 ;
        RECT 171.800 148.500 172.200 148.900 ;
        RECT 166.100 147.700 166.500 147.800 ;
        RECT 164.600 147.400 166.500 147.700 ;
        RECT 162.100 146.900 162.600 147.100 ;
        RECT 155.000 146.100 155.400 146.200 ;
        RECT 155.800 146.100 156.200 146.200 ;
        RECT 155.000 145.800 156.200 146.100 ;
        RECT 155.800 145.400 156.200 145.800 ;
        RECT 156.500 145.800 157.000 146.200 ;
        RECT 156.500 144.900 156.800 145.800 ;
        RECT 157.500 145.500 157.800 146.500 ;
        RECT 158.200 145.800 158.600 146.600 ;
        RECT 159.000 145.800 159.400 146.600 ;
        RECT 157.500 145.200 159.400 145.500 ;
        RECT 160.600 145.400 161.000 146.200 ;
        RECT 156.500 144.600 157.300 144.900 ;
        RECT 154.200 144.100 154.600 144.200 ;
        RECT 153.400 143.800 154.600 144.100 ;
        RECT 152.600 141.100 153.000 143.100 ;
        RECT 153.400 141.100 153.800 143.800 ;
        RECT 156.900 141.100 157.300 144.600 ;
        RECT 159.100 143.500 159.400 145.200 ;
        RECT 161.300 144.900 161.600 146.800 ;
        RECT 161.900 146.500 162.600 146.900 ;
        RECT 162.300 145.500 162.600 146.500 ;
        RECT 163.000 145.800 163.400 146.600 ;
        RECT 163.800 145.800 164.200 146.600 ;
        RECT 164.600 145.700 165.000 147.400 ;
        RECT 168.100 147.100 169.000 147.200 ;
        RECT 171.000 147.100 171.300 148.200 ;
        RECT 173.400 147.500 173.800 149.900 ;
        RECT 174.200 148.000 174.600 149.900 ;
        RECT 175.800 148.000 176.200 149.900 ;
        RECT 174.200 147.900 176.200 148.000 ;
        RECT 176.600 147.900 177.000 149.900 ;
        RECT 177.700 148.200 178.100 149.900 ;
        RECT 177.700 147.900 178.600 148.200 ;
        RECT 174.300 147.700 176.100 147.900 ;
        RECT 174.600 147.200 175.000 147.400 ;
        RECT 176.600 147.200 176.900 147.900 ;
        RECT 172.600 147.100 173.400 147.200 ;
        RECT 167.900 146.800 173.400 147.100 ;
        RECT 174.200 146.900 175.000 147.200 ;
        RECT 174.200 146.800 174.600 146.900 ;
        RECT 175.700 146.800 177.000 147.200 ;
        RECT 167.000 146.400 167.400 146.500 ;
        RECT 165.500 146.100 167.400 146.400 ;
        RECT 165.500 146.000 165.900 146.100 ;
        RECT 166.300 145.700 166.700 145.800 ;
        RECT 162.300 145.200 164.200 145.500 ;
        RECT 161.300 144.600 162.100 144.900 ;
        RECT 159.000 141.500 159.400 143.500 ;
        RECT 161.700 142.200 162.100 144.600 ;
        RECT 163.900 143.500 164.200 145.200 ;
        RECT 161.700 141.800 162.600 142.200 ;
        RECT 161.700 141.100 162.100 141.800 ;
        RECT 163.800 141.500 164.200 143.500 ;
        RECT 164.600 145.400 166.700 145.700 ;
        RECT 164.600 141.100 165.000 145.400 ;
        RECT 167.900 145.200 168.200 146.800 ;
        RECT 171.500 146.700 171.900 146.800 ;
        RECT 171.000 146.200 171.400 146.300 ;
        RECT 172.300 146.200 172.700 146.300 ;
        RECT 170.200 145.900 172.700 146.200 ;
        RECT 170.200 145.800 170.600 145.900 ;
        RECT 175.000 145.800 175.400 146.600 ;
        RECT 175.700 146.200 176.000 146.800 ;
        RECT 175.700 145.800 176.200 146.200 ;
        RECT 178.200 146.100 178.600 147.900 ;
        RECT 179.800 147.700 180.200 149.900 ;
        RECT 181.900 149.200 182.500 149.900 ;
        RECT 181.900 148.900 182.600 149.200 ;
        RECT 184.200 148.900 184.600 149.900 ;
        RECT 186.400 149.200 186.800 149.900 ;
        RECT 186.400 148.900 187.400 149.200 ;
        RECT 182.200 148.500 182.600 148.900 ;
        RECT 184.300 148.600 184.600 148.900 ;
        RECT 184.300 148.300 185.700 148.600 ;
        RECT 185.300 148.200 185.700 148.300 ;
        RECT 186.200 148.200 186.600 148.600 ;
        RECT 187.000 148.500 187.400 148.900 ;
        RECT 181.300 147.700 181.700 147.800 ;
        RECT 179.000 146.800 179.400 147.600 ;
        RECT 179.800 147.400 181.700 147.700 ;
        RECT 176.600 145.800 178.600 146.100 ;
        RECT 171.000 145.500 173.800 145.600 ;
        RECT 170.900 145.400 173.800 145.500 ;
        RECT 167.000 144.900 168.200 145.200 ;
        RECT 168.900 145.300 173.800 145.400 ;
        RECT 168.900 145.100 171.300 145.300 ;
        RECT 167.000 144.400 167.300 144.900 ;
        RECT 166.600 144.000 167.300 144.400 ;
        RECT 168.100 144.500 168.500 144.600 ;
        RECT 168.900 144.500 169.200 145.100 ;
        RECT 168.100 144.200 169.200 144.500 ;
        RECT 169.500 144.500 172.200 144.800 ;
        RECT 169.500 144.400 169.900 144.500 ;
        RECT 171.800 144.400 172.200 144.500 ;
        RECT 168.700 143.700 169.100 143.800 ;
        RECT 170.100 143.700 170.500 143.800 ;
        RECT 167.000 143.100 167.400 143.500 ;
        RECT 168.700 143.400 170.500 143.700 ;
        RECT 169.100 143.100 169.400 143.400 ;
        RECT 171.800 143.100 172.200 143.500 ;
        RECT 166.700 141.100 167.300 143.100 ;
        RECT 169.000 141.100 169.400 143.100 ;
        RECT 171.200 142.800 172.200 143.100 ;
        RECT 171.200 141.100 171.600 142.800 ;
        RECT 173.400 141.100 173.800 145.300 ;
        RECT 175.700 145.100 176.000 145.800 ;
        RECT 176.600 145.200 176.900 145.800 ;
        RECT 176.600 145.100 177.000 145.200 ;
        RECT 175.500 144.800 176.000 145.100 ;
        RECT 176.300 144.800 177.000 145.100 ;
        RECT 175.500 141.100 175.900 144.800 ;
        RECT 176.300 144.200 176.600 144.800 ;
        RECT 177.400 144.400 177.800 145.200 ;
        RECT 176.200 143.800 176.600 144.200 ;
        RECT 178.200 141.100 178.600 145.800 ;
        RECT 179.800 145.700 180.200 147.400 ;
        RECT 183.300 147.100 183.700 147.200 ;
        RECT 186.200 147.100 186.500 148.200 ;
        RECT 188.600 147.500 189.000 149.900 ;
        RECT 189.400 148.000 189.800 149.900 ;
        RECT 191.000 148.000 191.400 149.900 ;
        RECT 189.400 147.900 191.400 148.000 ;
        RECT 191.800 147.900 192.200 149.900 ;
        RECT 194.500 148.200 194.900 149.900 ;
        RECT 194.500 147.900 195.400 148.200 ;
        RECT 189.500 147.700 191.300 147.900 ;
        RECT 189.800 147.200 190.200 147.400 ;
        RECT 191.800 147.200 192.100 147.900 ;
        RECT 187.800 147.100 188.600 147.200 ;
        RECT 183.100 146.800 188.600 147.100 ;
        RECT 189.400 146.900 190.200 147.200 ;
        RECT 189.400 146.800 189.800 146.900 ;
        RECT 190.900 146.800 192.200 147.200 ;
        RECT 192.600 147.100 193.000 147.200 ;
        RECT 195.000 147.100 195.400 147.900 ;
        RECT 192.600 146.800 195.400 147.100 ;
        RECT 195.800 146.800 196.200 147.600 ;
        RECT 196.600 147.500 197.000 149.900 ;
        RECT 198.800 149.200 199.200 149.900 ;
        RECT 198.200 148.900 199.200 149.200 ;
        RECT 201.000 148.900 201.400 149.900 ;
        RECT 203.100 149.200 203.700 149.900 ;
        RECT 203.000 148.900 203.700 149.200 ;
        RECT 198.200 148.500 198.600 148.900 ;
        RECT 201.000 148.600 201.300 148.900 ;
        RECT 199.000 147.800 199.400 148.600 ;
        RECT 199.900 148.300 201.300 148.600 ;
        RECT 203.000 148.500 203.400 148.900 ;
        RECT 199.900 148.200 200.300 148.300 ;
        RECT 197.000 147.100 197.800 147.200 ;
        RECT 199.100 147.100 199.400 147.800 ;
        RECT 203.900 147.700 204.300 147.800 ;
        RECT 205.400 147.700 205.800 149.900 ;
        RECT 203.900 147.400 205.800 147.700 ;
        RECT 201.900 147.100 202.300 147.200 ;
        RECT 197.000 146.800 202.500 147.100 ;
        RECT 182.200 146.400 182.600 146.500 ;
        RECT 180.700 146.100 182.600 146.400 ;
        RECT 180.700 146.000 181.100 146.100 ;
        RECT 181.500 145.700 181.900 145.800 ;
        RECT 179.800 145.400 181.900 145.700 ;
        RECT 179.000 144.100 179.400 144.200 ;
        RECT 179.800 144.100 180.200 145.400 ;
        RECT 183.100 145.200 183.400 146.800 ;
        RECT 186.700 146.700 187.100 146.800 ;
        RECT 187.500 146.200 187.900 146.300 ;
        RECT 183.800 146.100 184.200 146.200 ;
        RECT 185.400 146.100 187.900 146.200 ;
        RECT 183.800 145.900 187.900 146.100 ;
        RECT 183.800 145.800 185.800 145.900 ;
        RECT 190.200 145.800 190.600 146.600 ;
        RECT 190.900 146.100 191.200 146.800 ;
        RECT 193.400 146.100 193.800 146.200 ;
        RECT 190.900 145.800 193.800 146.100 ;
        RECT 186.200 145.500 189.000 145.600 ;
        RECT 186.100 145.400 189.000 145.500 ;
        RECT 182.200 144.900 183.400 145.200 ;
        RECT 184.100 145.300 189.000 145.400 ;
        RECT 184.100 145.100 186.500 145.300 ;
        RECT 182.200 144.400 182.500 144.900 ;
        RECT 179.000 143.800 180.200 144.100 ;
        RECT 181.800 144.000 182.500 144.400 ;
        RECT 183.300 144.500 183.700 144.600 ;
        RECT 184.100 144.500 184.400 145.100 ;
        RECT 183.300 144.200 184.400 144.500 ;
        RECT 184.700 144.500 187.400 144.800 ;
        RECT 184.700 144.400 185.100 144.500 ;
        RECT 187.000 144.400 187.400 144.500 ;
        RECT 179.800 141.100 180.200 143.800 ;
        RECT 183.900 143.700 184.300 143.800 ;
        RECT 185.300 143.700 185.700 143.800 ;
        RECT 182.200 143.100 182.600 143.500 ;
        RECT 183.900 143.400 185.700 143.700 ;
        RECT 184.300 143.100 184.600 143.400 ;
        RECT 187.000 143.100 187.400 143.500 ;
        RECT 181.900 141.100 182.500 143.100 ;
        RECT 184.200 141.100 184.600 143.100 ;
        RECT 186.400 142.800 187.400 143.100 ;
        RECT 186.400 141.100 186.800 142.800 ;
        RECT 188.600 141.100 189.000 145.300 ;
        RECT 190.900 145.100 191.200 145.800 ;
        RECT 191.800 145.100 192.200 145.200 ;
        RECT 192.600 145.100 193.000 145.200 ;
        RECT 190.700 144.800 191.200 145.100 ;
        RECT 191.500 144.800 193.000 145.100 ;
        RECT 190.700 141.100 191.100 144.800 ;
        RECT 191.500 144.200 191.800 144.800 ;
        RECT 194.200 144.400 194.600 145.200 ;
        RECT 191.400 143.800 191.800 144.200 ;
        RECT 195.000 141.100 195.400 146.800 ;
        RECT 198.500 146.700 198.900 146.800 ;
        RECT 197.700 146.200 198.100 146.300 ;
        RECT 199.000 146.200 199.400 146.300 ;
        RECT 202.200 146.200 202.500 146.800 ;
        RECT 203.000 146.400 203.400 146.500 ;
        RECT 197.700 145.900 200.200 146.200 ;
        RECT 199.800 145.800 200.200 145.900 ;
        RECT 202.200 145.800 202.600 146.200 ;
        RECT 203.000 146.100 204.900 146.400 ;
        RECT 204.500 146.000 204.900 146.100 ;
        RECT 196.600 145.500 199.400 145.600 ;
        RECT 196.600 145.400 199.500 145.500 ;
        RECT 196.600 145.300 201.500 145.400 ;
        RECT 196.600 141.100 197.000 145.300 ;
        RECT 199.100 145.100 201.500 145.300 ;
        RECT 198.200 144.500 200.900 144.800 ;
        RECT 198.200 144.400 198.600 144.500 ;
        RECT 200.500 144.400 200.900 144.500 ;
        RECT 201.200 144.500 201.500 145.100 ;
        RECT 202.200 145.200 202.500 145.800 ;
        RECT 203.700 145.700 204.100 145.800 ;
        RECT 205.400 145.700 205.800 147.400 ;
        RECT 203.700 145.400 205.800 145.700 ;
        RECT 202.200 144.900 203.400 145.200 ;
        RECT 201.900 144.500 202.300 144.600 ;
        RECT 201.200 144.200 202.300 144.500 ;
        RECT 203.100 144.400 203.400 144.900 ;
        RECT 203.100 144.000 203.800 144.400 ;
        RECT 199.900 143.700 200.300 143.800 ;
        RECT 201.300 143.700 201.700 143.800 ;
        RECT 198.200 143.100 198.600 143.500 ;
        RECT 199.900 143.400 201.700 143.700 ;
        RECT 201.000 143.100 201.300 143.400 ;
        RECT 203.000 143.100 203.400 143.500 ;
        RECT 198.200 142.800 199.200 143.100 ;
        RECT 198.800 141.100 199.200 142.800 ;
        RECT 201.000 141.100 201.400 143.100 ;
        RECT 203.100 141.100 203.700 143.100 ;
        RECT 205.400 141.100 205.800 145.400 ;
        RECT 206.200 141.100 206.600 149.900 ;
        RECT 207.000 147.800 207.400 148.600 ;
        RECT 207.800 147.500 208.200 149.900 ;
        RECT 210.000 149.200 210.400 149.900 ;
        RECT 209.400 148.900 210.400 149.200 ;
        RECT 212.200 148.900 212.600 149.900 ;
        RECT 214.300 149.200 214.900 149.900 ;
        RECT 214.200 148.900 214.900 149.200 ;
        RECT 209.400 148.500 209.800 148.900 ;
        RECT 212.200 148.600 212.500 148.900 ;
        RECT 210.200 148.200 210.600 148.600 ;
        RECT 211.100 148.300 212.500 148.600 ;
        RECT 214.200 148.500 214.600 148.900 ;
        RECT 211.100 148.200 211.500 148.300 ;
        RECT 207.000 147.100 207.400 147.200 ;
        RECT 208.200 147.100 209.000 147.200 ;
        RECT 210.300 147.100 210.600 148.200 ;
        RECT 215.100 147.700 215.500 147.800 ;
        RECT 216.600 147.700 217.000 149.900 ;
        RECT 217.400 148.000 217.800 149.900 ;
        RECT 219.000 148.000 219.400 149.900 ;
        RECT 217.400 147.900 219.400 148.000 ;
        RECT 219.800 147.900 220.200 149.900 ;
        RECT 217.500 147.700 219.300 147.900 ;
        RECT 215.100 147.400 217.000 147.700 ;
        RECT 213.100 147.100 213.500 147.200 ;
        RECT 207.000 146.800 213.700 147.100 ;
        RECT 209.700 146.700 210.100 146.800 ;
        RECT 208.900 146.200 209.300 146.300 ;
        RECT 210.200 146.200 210.600 146.300 ;
        RECT 213.400 146.200 213.700 146.800 ;
        RECT 214.200 146.400 214.600 146.500 ;
        RECT 208.900 145.900 211.400 146.200 ;
        RECT 211.000 145.800 211.400 145.900 ;
        RECT 213.400 145.800 213.800 146.200 ;
        RECT 214.200 146.100 216.100 146.400 ;
        RECT 215.700 146.000 216.100 146.100 ;
        RECT 207.800 145.500 210.600 145.600 ;
        RECT 207.800 145.400 210.700 145.500 ;
        RECT 207.800 145.300 212.700 145.400 ;
        RECT 207.800 141.100 208.200 145.300 ;
        RECT 210.300 145.100 212.700 145.300 ;
        RECT 209.400 144.500 212.100 144.800 ;
        RECT 209.400 144.400 209.800 144.500 ;
        RECT 211.700 144.400 212.100 144.500 ;
        RECT 212.400 144.500 212.700 145.100 ;
        RECT 213.400 145.200 213.700 145.800 ;
        RECT 214.900 145.700 215.300 145.800 ;
        RECT 216.600 145.700 217.000 147.400 ;
        RECT 217.800 147.200 218.200 147.400 ;
        RECT 219.800 147.200 220.100 147.900 ;
        RECT 220.600 147.500 221.000 149.900 ;
        RECT 222.800 149.200 223.200 149.900 ;
        RECT 222.200 148.900 223.200 149.200 ;
        RECT 225.000 148.900 225.400 149.900 ;
        RECT 227.100 149.200 227.700 149.900 ;
        RECT 227.000 148.900 227.700 149.200 ;
        RECT 222.200 148.500 222.600 148.900 ;
        RECT 225.000 148.600 225.300 148.900 ;
        RECT 223.000 148.200 223.400 148.600 ;
        RECT 223.900 148.300 225.300 148.600 ;
        RECT 227.000 148.500 227.400 148.900 ;
        RECT 223.900 148.200 224.300 148.300 ;
        RECT 217.400 146.900 218.200 147.200 ;
        RECT 217.400 146.800 217.800 146.900 ;
        RECT 218.900 146.800 220.200 147.200 ;
        RECT 221.000 147.100 221.800 147.200 ;
        RECT 223.100 147.100 223.400 148.200 ;
        RECT 226.200 148.100 226.600 148.200 ;
        RECT 226.200 147.800 228.200 148.100 ;
        RECT 227.800 147.700 228.300 147.800 ;
        RECT 229.400 147.700 229.800 149.900 ;
        RECT 227.800 147.400 229.800 147.700 ;
        RECT 223.800 147.100 224.200 147.200 ;
        RECT 224.600 147.100 225.000 147.200 ;
        RECT 225.900 147.100 226.300 147.200 ;
        RECT 221.000 146.800 226.500 147.100 ;
        RECT 218.200 145.800 218.600 146.600 ;
        RECT 218.900 146.100 219.200 146.800 ;
        RECT 222.500 146.700 222.900 146.800 ;
        RECT 221.700 146.200 222.100 146.300 ;
        RECT 223.000 146.200 223.400 146.300 ;
        RECT 219.800 146.100 220.200 146.200 ;
        RECT 218.900 145.800 220.200 146.100 ;
        RECT 221.700 145.900 224.200 146.200 ;
        RECT 223.800 145.800 224.200 145.900 ;
        RECT 214.900 145.400 217.000 145.700 ;
        RECT 213.400 144.900 214.600 145.200 ;
        RECT 213.100 144.500 213.500 144.600 ;
        RECT 212.400 144.200 213.500 144.500 ;
        RECT 214.300 144.400 214.600 144.900 ;
        RECT 214.300 144.000 215.000 144.400 ;
        RECT 211.100 143.700 211.500 143.800 ;
        RECT 212.500 143.700 212.900 143.800 ;
        RECT 209.400 143.100 209.800 143.500 ;
        RECT 211.100 143.400 212.900 143.700 ;
        RECT 212.200 143.100 212.500 143.400 ;
        RECT 214.200 143.100 214.600 143.500 ;
        RECT 209.400 142.800 210.400 143.100 ;
        RECT 210.000 141.100 210.400 142.800 ;
        RECT 212.200 141.100 212.600 143.100 ;
        RECT 214.300 141.100 214.900 143.100 ;
        RECT 216.600 141.100 217.000 145.400 ;
        RECT 218.900 145.100 219.200 145.800 ;
        RECT 220.600 145.500 223.400 145.600 ;
        RECT 220.600 145.400 223.500 145.500 ;
        RECT 220.600 145.300 225.500 145.400 ;
        RECT 219.800 145.100 220.200 145.200 ;
        RECT 218.700 144.800 219.200 145.100 ;
        RECT 219.500 144.800 220.200 145.100 ;
        RECT 218.700 141.100 219.100 144.800 ;
        RECT 219.500 144.200 219.800 144.800 ;
        RECT 219.400 143.800 219.800 144.200 ;
        RECT 220.600 141.100 221.000 145.300 ;
        RECT 223.100 145.100 225.500 145.300 ;
        RECT 222.200 144.500 224.900 144.800 ;
        RECT 222.200 144.400 222.600 144.500 ;
        RECT 224.500 144.400 224.900 144.500 ;
        RECT 225.200 144.500 225.500 145.100 ;
        RECT 226.200 145.200 226.500 146.800 ;
        RECT 227.000 146.400 227.400 146.500 ;
        RECT 227.000 146.100 228.900 146.400 ;
        RECT 228.500 146.000 228.900 146.100 ;
        RECT 227.700 145.700 228.100 145.800 ;
        RECT 229.400 145.700 229.800 147.400 ;
        RECT 227.700 145.400 229.800 145.700 ;
        RECT 226.200 144.900 227.400 145.200 ;
        RECT 225.900 144.500 226.300 144.600 ;
        RECT 225.200 144.200 226.300 144.500 ;
        RECT 227.100 144.400 227.400 144.900 ;
        RECT 227.100 144.000 227.800 144.400 ;
        RECT 223.900 143.700 224.300 143.800 ;
        RECT 225.300 143.700 225.700 143.800 ;
        RECT 222.200 143.100 222.600 143.500 ;
        RECT 223.900 143.400 225.700 143.700 ;
        RECT 225.000 143.100 225.300 143.400 ;
        RECT 227.000 143.100 227.400 143.500 ;
        RECT 222.200 142.800 223.200 143.100 ;
        RECT 222.800 141.100 223.200 142.800 ;
        RECT 225.000 141.100 225.400 143.100 ;
        RECT 227.100 141.100 227.700 143.100 ;
        RECT 229.400 141.100 229.800 145.400 ;
        RECT 0.600 135.700 1.000 139.900 ;
        RECT 2.800 138.200 3.200 139.900 ;
        RECT 2.200 137.900 3.200 138.200 ;
        RECT 5.000 137.900 5.400 139.900 ;
        RECT 7.100 137.900 7.700 139.900 ;
        RECT 2.200 137.500 2.600 137.900 ;
        RECT 5.000 137.600 5.300 137.900 ;
        RECT 3.900 137.300 5.700 137.600 ;
        RECT 7.000 137.500 7.400 137.900 ;
        RECT 3.900 137.200 4.300 137.300 ;
        RECT 5.300 137.200 5.700 137.300 ;
        RECT 9.400 137.100 9.800 139.900 ;
        RECT 10.200 137.100 10.600 137.200 ;
        RECT 2.200 136.500 2.600 136.600 ;
        RECT 4.500 136.500 4.900 136.600 ;
        RECT 2.200 136.200 4.900 136.500 ;
        RECT 5.200 136.500 6.300 136.800 ;
        RECT 5.200 135.900 5.500 136.500 ;
        RECT 5.900 136.400 6.300 136.500 ;
        RECT 7.100 136.600 7.800 137.000 ;
        RECT 9.400 136.800 10.600 137.100 ;
        RECT 7.100 136.100 7.400 136.600 ;
        RECT 3.100 135.700 5.500 135.900 ;
        RECT 0.600 135.600 5.500 135.700 ;
        RECT 6.200 135.800 7.400 136.100 ;
        RECT 0.600 135.500 3.500 135.600 ;
        RECT 0.600 135.400 3.400 135.500 ;
        RECT 3.800 135.100 4.200 135.200 ;
        RECT 1.700 134.800 4.200 135.100 ;
        RECT 1.700 134.700 2.100 134.800 ;
        RECT 2.500 134.200 2.900 134.300 ;
        RECT 6.200 134.200 6.500 135.800 ;
        RECT 9.400 135.600 9.800 136.800 ;
        RECT 7.700 135.300 9.800 135.600 ;
        RECT 7.700 135.200 8.100 135.300 ;
        RECT 8.500 134.900 8.900 135.000 ;
        RECT 7.000 134.600 8.900 134.900 ;
        RECT 7.000 134.500 7.400 134.600 ;
        RECT 1.000 133.900 6.500 134.200 ;
        RECT 1.000 133.800 1.800 133.900 ;
        RECT 0.600 131.100 1.000 133.500 ;
        RECT 3.100 132.800 3.400 133.900 ;
        RECT 4.600 133.800 5.000 133.900 ;
        RECT 5.900 133.800 6.300 133.900 ;
        RECT 9.400 133.600 9.800 135.300 ;
        RECT 11.000 135.100 11.400 139.900 ;
        RECT 13.000 136.800 13.400 137.200 ;
        RECT 11.800 135.800 12.200 136.600 ;
        RECT 13.000 136.200 13.300 136.800 ;
        RECT 13.700 136.200 14.100 139.900 ;
        RECT 12.600 135.900 13.300 136.200 ;
        RECT 13.600 135.900 14.100 136.200 ;
        RECT 12.600 135.800 13.000 135.900 ;
        RECT 12.600 135.100 12.900 135.800 ;
        RECT 11.000 134.800 12.900 135.100 ;
        RECT 7.900 133.300 9.800 133.600 ;
        RECT 10.200 133.400 10.600 134.200 ;
        RECT 7.900 133.200 8.300 133.300 ;
        RECT 2.200 132.100 2.600 132.500 ;
        RECT 3.000 132.400 3.400 132.800 ;
        RECT 3.900 132.700 4.300 132.800 ;
        RECT 3.900 132.400 5.300 132.700 ;
        RECT 5.000 132.100 5.300 132.400 ;
        RECT 7.000 132.100 7.400 132.500 ;
        RECT 2.200 131.800 3.200 132.100 ;
        RECT 2.800 131.100 3.200 131.800 ;
        RECT 5.000 131.100 5.400 132.100 ;
        RECT 7.000 131.800 7.700 132.100 ;
        RECT 7.100 131.100 7.700 131.800 ;
        RECT 9.400 131.100 9.800 133.300 ;
        RECT 11.000 133.100 11.400 134.800 ;
        RECT 13.600 134.200 13.900 135.900 ;
        RECT 15.800 135.700 16.200 139.900 ;
        RECT 18.000 138.200 18.400 139.900 ;
        RECT 17.400 137.900 18.400 138.200 ;
        RECT 20.200 137.900 20.600 139.900 ;
        RECT 22.300 137.900 22.900 139.900 ;
        RECT 17.400 137.500 17.800 137.900 ;
        RECT 20.200 137.600 20.500 137.900 ;
        RECT 19.100 137.300 20.900 137.600 ;
        RECT 22.200 137.500 22.600 137.900 ;
        RECT 19.100 137.200 19.500 137.300 ;
        RECT 20.500 137.200 20.900 137.300 ;
        RECT 17.400 136.500 17.800 136.600 ;
        RECT 19.700 136.500 20.100 136.600 ;
        RECT 17.400 136.200 20.100 136.500 ;
        RECT 20.400 136.500 21.500 136.800 ;
        RECT 20.400 135.900 20.700 136.500 ;
        RECT 21.100 136.400 21.500 136.500 ;
        RECT 22.300 136.600 23.000 137.000 ;
        RECT 22.300 136.100 22.600 136.600 ;
        RECT 18.300 135.700 20.700 135.900 ;
        RECT 15.800 135.600 20.700 135.700 ;
        RECT 21.400 135.800 22.600 136.100 ;
        RECT 15.800 135.500 18.700 135.600 ;
        RECT 15.800 135.400 18.600 135.500 ;
        RECT 14.200 134.400 14.600 135.200 ;
        RECT 19.000 135.100 19.400 135.200 ;
        RECT 20.600 135.100 21.000 135.200 ;
        RECT 16.900 134.800 21.000 135.100 ;
        RECT 16.900 134.700 17.300 134.800 ;
        RECT 17.700 134.200 18.100 134.300 ;
        RECT 21.400 134.200 21.700 135.800 ;
        RECT 24.600 135.600 25.000 139.900 ;
        RECT 26.700 136.200 27.100 139.900 ;
        RECT 27.400 136.800 27.800 137.200 ;
        RECT 27.500 136.200 27.800 136.800 ;
        RECT 26.700 135.900 27.200 136.200 ;
        RECT 27.500 135.900 28.200 136.200 ;
        RECT 22.900 135.300 25.000 135.600 ;
        RECT 22.900 135.200 23.300 135.300 ;
        RECT 23.700 134.900 24.100 135.000 ;
        RECT 22.200 134.600 24.100 134.900 ;
        RECT 22.200 134.500 22.600 134.600 ;
        RECT 11.800 134.100 12.200 134.200 ;
        RECT 12.600 134.100 13.900 134.200 ;
        RECT 15.000 134.100 15.400 134.200 ;
        RECT 11.800 133.800 13.900 134.100 ;
        RECT 14.600 133.800 15.400 134.100 ;
        RECT 16.200 133.900 21.700 134.200 ;
        RECT 16.200 133.800 17.000 133.900 ;
        RECT 12.700 133.100 13.000 133.800 ;
        RECT 14.600 133.600 15.000 133.800 ;
        RECT 13.500 133.100 15.300 133.300 ;
        RECT 11.000 132.800 11.900 133.100 ;
        RECT 11.500 131.100 11.900 132.800 ;
        RECT 12.600 131.100 13.000 133.100 ;
        RECT 13.400 133.000 15.400 133.100 ;
        RECT 13.400 131.100 13.800 133.000 ;
        RECT 15.000 131.100 15.400 133.000 ;
        RECT 15.800 131.100 16.200 133.500 ;
        RECT 18.300 133.200 18.600 133.900 ;
        RECT 21.100 133.800 21.700 133.900 ;
        RECT 17.400 132.100 17.800 132.500 ;
        RECT 18.200 132.400 18.600 133.200 ;
        RECT 21.400 133.200 21.700 133.800 ;
        RECT 24.600 133.600 25.000 135.300 ;
        RECT 26.900 135.200 27.200 135.900 ;
        RECT 27.800 135.800 28.200 135.900 ;
        RECT 28.600 135.700 29.000 139.900 ;
        RECT 30.800 138.200 31.200 139.900 ;
        RECT 30.200 137.900 31.200 138.200 ;
        RECT 33.000 137.900 33.400 139.900 ;
        RECT 35.100 137.900 35.700 139.900 ;
        RECT 30.200 137.500 30.600 137.900 ;
        RECT 33.000 137.600 33.300 137.900 ;
        RECT 31.900 137.300 33.700 137.600 ;
        RECT 35.000 137.500 35.400 137.900 ;
        RECT 31.900 137.200 32.300 137.300 ;
        RECT 33.300 137.200 33.700 137.300 ;
        RECT 30.200 136.500 30.600 136.600 ;
        RECT 32.500 136.500 32.900 136.600 ;
        RECT 30.200 136.200 32.900 136.500 ;
        RECT 33.200 136.500 34.300 136.800 ;
        RECT 33.200 135.900 33.500 136.500 ;
        RECT 33.900 136.400 34.300 136.500 ;
        RECT 35.100 136.600 35.800 137.000 ;
        RECT 35.100 136.100 35.400 136.600 ;
        RECT 31.100 135.700 33.500 135.900 ;
        RECT 28.600 135.600 33.500 135.700 ;
        RECT 34.200 135.800 35.400 136.100 ;
        RECT 28.600 135.500 31.500 135.600 ;
        RECT 28.600 135.400 31.400 135.500 ;
        RECT 26.200 134.400 26.600 135.200 ;
        RECT 26.900 134.800 27.400 135.200 ;
        RECT 31.800 135.100 32.200 135.200 ;
        RECT 32.600 135.100 33.000 135.200 ;
        RECT 29.700 134.800 33.000 135.100 ;
        RECT 26.900 134.200 27.200 134.800 ;
        RECT 29.700 134.700 30.100 134.800 ;
        RECT 30.500 134.200 30.900 134.300 ;
        RECT 34.200 134.200 34.500 135.800 ;
        RECT 37.400 135.600 37.800 139.900 ;
        RECT 41.100 136.200 41.500 139.900 ;
        RECT 41.800 136.800 42.200 137.200 ;
        RECT 41.900 136.200 42.200 136.800 ;
        RECT 43.400 136.800 43.800 137.200 ;
        RECT 43.400 136.200 43.700 136.800 ;
        RECT 44.100 136.200 44.500 139.900 ;
        RECT 41.100 135.900 41.600 136.200 ;
        RECT 41.900 135.900 42.600 136.200 ;
        RECT 35.700 135.300 37.800 135.600 ;
        RECT 35.700 135.200 36.100 135.300 ;
        RECT 36.500 134.900 36.900 135.000 ;
        RECT 35.000 134.600 36.900 134.900 ;
        RECT 35.000 134.500 35.400 134.600 ;
        RECT 25.400 134.100 25.800 134.200 ;
        RECT 25.400 133.800 26.200 134.100 ;
        RECT 26.900 133.800 28.200 134.200 ;
        RECT 29.000 133.900 34.500 134.200 ;
        RECT 29.000 133.800 29.800 133.900 ;
        RECT 25.800 133.600 26.200 133.800 ;
        RECT 23.100 133.300 25.000 133.600 ;
        RECT 23.100 133.200 23.500 133.300 ;
        RECT 21.400 132.800 21.800 133.200 ;
        RECT 19.100 132.700 19.500 132.800 ;
        RECT 19.100 132.400 20.500 132.700 ;
        RECT 20.200 132.100 20.500 132.400 ;
        RECT 22.200 132.100 22.600 132.500 ;
        RECT 17.400 131.800 18.400 132.100 ;
        RECT 18.000 131.100 18.400 131.800 ;
        RECT 20.200 131.100 20.600 132.100 ;
        RECT 22.200 131.800 22.900 132.100 ;
        RECT 22.300 131.100 22.900 131.800 ;
        RECT 24.600 131.100 25.000 133.300 ;
        RECT 25.500 133.100 27.300 133.300 ;
        RECT 27.800 133.100 28.100 133.800 ;
        RECT 25.400 133.000 27.400 133.100 ;
        RECT 25.400 131.100 25.800 133.000 ;
        RECT 27.000 131.100 27.400 133.000 ;
        RECT 27.800 131.100 28.200 133.100 ;
        RECT 28.600 131.100 29.000 133.500 ;
        RECT 31.100 132.800 31.400 133.900 ;
        RECT 33.400 133.800 34.300 133.900 ;
        RECT 37.400 133.600 37.800 135.300 ;
        RECT 41.300 135.200 41.600 135.900 ;
        RECT 42.200 135.800 42.600 135.900 ;
        RECT 43.000 135.900 43.700 136.200 ;
        RECT 44.000 135.900 44.500 136.200 ;
        RECT 43.000 135.800 43.400 135.900 ;
        RECT 39.800 135.100 40.200 135.200 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 39.800 134.800 41.000 135.100 ;
        RECT 40.600 134.400 41.000 134.800 ;
        RECT 41.300 134.800 41.800 135.200 ;
        RECT 42.200 135.100 42.500 135.800 ;
        RECT 44.000 135.100 44.300 135.900 ;
        RECT 46.200 135.800 46.600 136.600 ;
        RECT 42.200 134.800 44.300 135.100 ;
        RECT 41.300 134.200 41.600 134.800 ;
        RECT 44.000 134.200 44.300 134.800 ;
        RECT 44.600 134.400 45.000 135.200 ;
        RECT 39.800 134.100 40.200 134.200 ;
        RECT 39.800 133.800 40.600 134.100 ;
        RECT 41.300 133.800 42.600 134.200 ;
        RECT 43.000 133.800 44.300 134.200 ;
        RECT 45.400 134.100 45.800 134.200 ;
        RECT 45.000 133.800 45.800 134.100 ;
        RECT 40.200 133.600 40.600 133.800 ;
        RECT 35.900 133.300 37.800 133.600 ;
        RECT 35.900 133.200 36.300 133.300 ;
        RECT 30.200 132.100 30.600 132.500 ;
        RECT 31.000 132.400 31.400 132.800 ;
        RECT 31.900 132.700 32.300 132.800 ;
        RECT 31.900 132.400 33.300 132.700 ;
        RECT 33.000 132.100 33.300 132.400 ;
        RECT 35.000 132.100 35.400 132.500 ;
        RECT 30.200 131.800 31.200 132.100 ;
        RECT 30.800 131.100 31.200 131.800 ;
        RECT 33.000 131.100 33.400 132.100 ;
        RECT 35.000 131.800 35.700 132.100 ;
        RECT 35.100 131.100 35.700 131.800 ;
        RECT 37.400 131.100 37.800 133.300 ;
        RECT 39.900 133.100 41.700 133.300 ;
        RECT 42.200 133.100 42.500 133.800 ;
        RECT 43.100 133.100 43.400 133.800 ;
        RECT 45.000 133.600 45.400 133.800 ;
        RECT 43.900 133.100 45.700 133.300 ;
        RECT 47.000 133.100 47.400 139.900 ;
        RECT 49.400 136.400 49.800 139.900 ;
        RECT 49.300 135.900 49.800 136.400 ;
        RECT 51.000 136.200 51.400 139.900 ;
        RECT 50.100 135.900 51.400 136.200 ;
        RECT 48.600 134.800 49.000 135.200 ;
        RECT 47.800 133.400 48.200 134.200 ;
        RECT 48.600 134.100 48.900 134.800 ;
        RECT 49.300 134.200 49.600 135.900 ;
        RECT 50.100 134.900 50.400 135.900 ;
        RECT 51.800 135.700 52.200 139.900 ;
        RECT 54.000 138.200 54.400 139.900 ;
        RECT 53.400 137.900 54.400 138.200 ;
        RECT 56.200 137.900 56.600 139.900 ;
        RECT 58.300 137.900 58.900 139.900 ;
        RECT 53.400 137.500 53.800 137.900 ;
        RECT 56.200 137.600 56.500 137.900 ;
        RECT 55.100 137.300 56.900 137.600 ;
        RECT 58.200 137.500 58.600 137.900 ;
        RECT 55.100 137.200 55.500 137.300 ;
        RECT 56.500 137.200 56.900 137.300 ;
        RECT 53.400 136.500 53.800 136.600 ;
        RECT 55.700 136.500 56.100 136.600 ;
        RECT 53.400 136.200 56.100 136.500 ;
        RECT 56.400 136.500 57.500 136.800 ;
        RECT 56.400 135.900 56.700 136.500 ;
        RECT 57.100 136.400 57.500 136.500 ;
        RECT 58.300 136.600 59.000 137.000 ;
        RECT 58.300 136.100 58.600 136.600 ;
        RECT 54.300 135.700 56.700 135.900 ;
        RECT 51.800 135.600 56.700 135.700 ;
        RECT 57.400 135.800 58.600 136.100 ;
        RECT 51.800 135.500 54.700 135.600 ;
        RECT 51.800 135.400 54.600 135.500 ;
        RECT 57.400 135.200 57.700 135.800 ;
        RECT 60.600 135.600 61.000 139.900 ;
        RECT 61.400 136.100 61.800 136.200 ;
        RECT 62.200 136.100 62.600 139.900 ;
        RECT 61.400 135.800 62.600 136.100 ;
        RECT 63.000 135.800 63.400 136.600 ;
        RECT 58.900 135.300 61.000 135.600 ;
        RECT 58.900 135.200 59.300 135.300 ;
        RECT 49.900 134.500 50.400 134.900 ;
        RECT 49.300 134.100 49.800 134.200 ;
        RECT 48.600 133.800 49.800 134.100 ;
        RECT 39.800 133.000 41.800 133.100 ;
        RECT 39.800 131.100 40.200 133.000 ;
        RECT 41.400 131.100 41.800 133.000 ;
        RECT 42.200 131.100 42.600 133.100 ;
        RECT 43.000 131.100 43.400 133.100 ;
        RECT 43.800 133.000 45.800 133.100 ;
        RECT 43.800 131.100 44.200 133.000 ;
        RECT 45.400 131.100 45.800 133.000 ;
        RECT 46.500 132.800 47.400 133.100 ;
        RECT 49.300 133.100 49.600 133.800 ;
        RECT 50.100 133.700 50.400 134.500 ;
        RECT 50.900 134.800 51.400 135.200 ;
        RECT 55.000 135.100 55.400 135.200 ;
        RECT 52.900 134.800 55.400 135.100 ;
        RECT 57.400 134.800 57.800 135.200 ;
        RECT 59.700 134.900 60.100 135.000 ;
        RECT 50.900 134.400 51.300 134.800 ;
        RECT 52.900 134.700 53.300 134.800 ;
        RECT 53.700 134.200 54.100 134.300 ;
        RECT 57.400 134.200 57.700 134.800 ;
        RECT 58.200 134.600 60.100 134.900 ;
        RECT 58.200 134.500 58.600 134.600 ;
        RECT 52.200 133.900 57.700 134.200 ;
        RECT 52.200 133.800 53.000 133.900 ;
        RECT 50.100 133.400 51.400 133.700 ;
        RECT 49.300 132.800 49.800 133.100 ;
        RECT 46.500 132.200 46.900 132.800 ;
        RECT 46.200 131.800 46.900 132.200 ;
        RECT 46.500 131.100 46.900 131.800 ;
        RECT 49.400 131.100 49.800 132.800 ;
        RECT 51.000 131.100 51.400 133.400 ;
        RECT 51.800 131.100 52.200 133.500 ;
        RECT 54.300 132.800 54.600 133.900 ;
        RECT 57.100 133.800 57.500 133.900 ;
        RECT 60.600 133.600 61.000 135.300 ;
        RECT 59.100 133.300 61.000 133.600 ;
        RECT 61.400 133.400 61.800 134.200 ;
        RECT 59.100 133.200 59.500 133.300 ;
        RECT 53.400 132.100 53.800 132.500 ;
        RECT 54.200 132.400 54.600 132.800 ;
        RECT 55.100 132.700 55.500 132.800 ;
        RECT 55.100 132.400 56.500 132.700 ;
        RECT 56.200 132.100 56.500 132.400 ;
        RECT 58.200 132.100 58.600 132.500 ;
        RECT 53.400 131.800 54.400 132.100 ;
        RECT 54.000 131.100 54.400 131.800 ;
        RECT 56.200 131.100 56.600 132.100 ;
        RECT 58.200 131.800 58.900 132.100 ;
        RECT 58.300 131.100 58.900 131.800 ;
        RECT 60.600 131.100 61.000 133.300 ;
        RECT 62.200 133.100 62.600 135.800 ;
        RECT 63.800 135.700 64.200 139.900 ;
        RECT 66.000 138.200 66.400 139.900 ;
        RECT 65.400 137.900 66.400 138.200 ;
        RECT 68.200 137.900 68.600 139.900 ;
        RECT 70.300 137.900 70.900 139.900 ;
        RECT 65.400 137.500 65.800 137.900 ;
        RECT 68.200 137.600 68.500 137.900 ;
        RECT 67.100 137.300 68.900 137.600 ;
        RECT 70.200 137.500 70.600 137.900 ;
        RECT 67.100 137.200 67.500 137.300 ;
        RECT 68.500 137.200 68.900 137.300 ;
        RECT 65.400 136.500 65.800 136.600 ;
        RECT 67.700 136.500 68.100 136.600 ;
        RECT 65.400 136.200 68.100 136.500 ;
        RECT 68.400 136.500 69.500 136.800 ;
        RECT 68.400 135.900 68.700 136.500 ;
        RECT 69.100 136.400 69.500 136.500 ;
        RECT 70.300 136.600 71.000 137.000 ;
        RECT 70.300 136.100 70.600 136.600 ;
        RECT 66.300 135.700 68.700 135.900 ;
        RECT 63.800 135.600 68.700 135.700 ;
        RECT 69.400 135.800 70.600 136.100 ;
        RECT 63.800 135.500 66.700 135.600 ;
        RECT 63.800 135.400 66.600 135.500 ;
        RECT 67.000 135.100 67.400 135.200 ;
        RECT 67.800 135.100 68.200 135.200 ;
        RECT 64.900 134.800 68.200 135.100 ;
        RECT 64.900 134.700 65.300 134.800 ;
        RECT 65.700 134.200 66.100 134.300 ;
        RECT 69.400 134.200 69.700 135.800 ;
        RECT 72.600 135.600 73.000 139.900 ;
        RECT 73.800 136.800 74.200 137.200 ;
        RECT 73.800 136.200 74.100 136.800 ;
        RECT 74.500 136.200 74.900 139.900 ;
        RECT 73.400 135.900 74.100 136.200 ;
        RECT 74.400 135.900 74.900 136.200 ;
        RECT 73.400 135.800 73.800 135.900 ;
        RECT 70.900 135.300 73.000 135.600 ;
        RECT 70.900 135.200 71.300 135.300 ;
        RECT 71.700 134.900 72.100 135.000 ;
        RECT 70.200 134.600 72.100 134.900 ;
        RECT 70.200 134.500 70.600 134.600 ;
        RECT 64.200 133.900 69.700 134.200 ;
        RECT 64.200 133.800 65.000 133.900 ;
        RECT 62.200 132.800 63.100 133.100 ;
        RECT 62.700 131.100 63.100 132.800 ;
        RECT 63.800 131.100 64.200 133.500 ;
        RECT 66.300 132.800 66.600 133.900 ;
        RECT 69.100 133.800 69.500 133.900 ;
        RECT 72.600 133.600 73.000 135.300 ;
        RECT 73.400 135.100 73.800 135.200 ;
        RECT 74.400 135.100 74.700 135.900 ;
        RECT 76.600 135.800 77.000 136.600 ;
        RECT 73.400 134.800 74.700 135.100 ;
        RECT 74.400 134.200 74.700 134.800 ;
        RECT 75.000 134.400 75.400 135.200 ;
        RECT 73.400 133.800 74.700 134.200 ;
        RECT 75.800 134.100 76.200 134.200 ;
        RECT 75.400 133.800 76.200 134.100 ;
        RECT 71.100 133.300 73.000 133.600 ;
        RECT 71.100 133.200 71.500 133.300 ;
        RECT 65.400 132.100 65.800 132.500 ;
        RECT 66.200 132.400 66.600 132.800 ;
        RECT 67.100 132.700 67.500 132.800 ;
        RECT 67.100 132.400 68.500 132.700 ;
        RECT 68.200 132.100 68.500 132.400 ;
        RECT 70.200 132.100 70.600 132.500 ;
        RECT 65.400 131.800 66.400 132.100 ;
        RECT 66.000 131.100 66.400 131.800 ;
        RECT 68.200 131.100 68.600 132.100 ;
        RECT 70.200 131.800 70.900 132.100 ;
        RECT 70.300 131.100 70.900 131.800 ;
        RECT 72.600 131.100 73.000 133.300 ;
        RECT 73.500 133.100 73.800 133.800 ;
        RECT 75.400 133.600 75.800 133.800 ;
        RECT 74.300 133.100 76.100 133.300 ;
        RECT 77.400 133.100 77.800 139.900 ;
        RECT 79.800 137.900 80.200 139.900 ;
        RECT 79.900 137.800 80.200 137.900 ;
        RECT 81.400 137.900 81.800 139.900 ;
        RECT 81.400 137.800 81.700 137.900 ;
        RECT 79.900 137.500 81.700 137.800 ;
        RECT 80.600 136.400 81.000 137.200 ;
        RECT 81.400 136.200 81.700 137.500 ;
        RECT 83.500 136.200 83.900 139.900 ;
        RECT 84.200 136.800 84.600 137.200 ;
        RECT 84.300 136.200 84.600 136.800 ;
        RECT 79.000 135.400 79.400 136.200 ;
        RECT 81.400 135.800 81.800 136.200 ;
        RECT 83.500 135.900 84.000 136.200 ;
        RECT 84.300 135.900 85.000 136.200 ;
        RECT 79.800 134.800 80.600 135.200 ;
        RECT 81.400 134.200 81.700 135.800 ;
        RECT 83.700 135.200 84.000 135.900 ;
        RECT 84.600 135.800 85.000 135.900 ;
        RECT 87.000 135.700 87.400 139.900 ;
        RECT 89.200 138.200 89.600 139.900 ;
        RECT 88.600 137.900 89.600 138.200 ;
        RECT 91.400 137.900 91.800 139.900 ;
        RECT 93.500 137.900 94.100 139.900 ;
        RECT 88.600 137.500 89.000 137.900 ;
        RECT 91.400 137.600 91.700 137.900 ;
        RECT 90.300 137.300 92.100 137.600 ;
        RECT 93.400 137.500 93.800 137.900 ;
        RECT 90.300 137.200 90.700 137.300 ;
        RECT 91.700 137.200 92.100 137.300 ;
        RECT 88.600 136.500 89.000 136.600 ;
        RECT 90.900 136.500 91.300 136.600 ;
        RECT 88.600 136.200 91.300 136.500 ;
        RECT 91.600 136.500 92.700 136.800 ;
        RECT 91.600 135.900 91.900 136.500 ;
        RECT 92.300 136.400 92.700 136.500 ;
        RECT 93.500 136.600 94.200 137.000 ;
        RECT 93.500 136.100 93.800 136.600 ;
        RECT 89.500 135.700 91.900 135.900 ;
        RECT 87.000 135.600 91.900 135.700 ;
        RECT 92.600 135.800 93.800 136.100 ;
        RECT 87.000 135.500 89.900 135.600 ;
        RECT 87.000 135.400 89.800 135.500 ;
        RECT 83.000 134.400 83.400 135.200 ;
        RECT 83.700 134.800 84.200 135.200 ;
        RECT 90.200 135.100 90.600 135.200 ;
        RECT 88.100 134.800 90.600 135.100 ;
        RECT 83.700 134.200 84.000 134.800 ;
        RECT 88.100 134.700 88.500 134.800 ;
        RECT 89.400 134.700 89.800 134.800 ;
        RECT 88.900 134.200 89.300 134.300 ;
        RECT 92.600 134.200 92.900 135.800 ;
        RECT 95.800 135.600 96.200 139.900 ;
        RECT 97.900 136.300 98.300 139.900 ;
        RECT 99.800 136.400 100.200 139.900 ;
        RECT 97.400 135.900 98.300 136.300 ;
        RECT 99.700 135.900 100.200 136.400 ;
        RECT 101.400 136.200 101.800 139.900 ;
        RECT 103.000 137.900 103.400 139.900 ;
        RECT 103.100 137.800 103.400 137.900 ;
        RECT 104.600 137.900 105.000 139.900 ;
        RECT 106.200 137.900 106.600 139.900 ;
        RECT 104.600 137.800 104.900 137.900 ;
        RECT 103.100 137.500 104.900 137.800 ;
        RECT 106.300 137.800 106.600 137.900 ;
        RECT 107.800 137.900 108.200 139.900 ;
        RECT 107.800 137.800 108.100 137.900 ;
        RECT 106.300 137.500 108.100 137.800 ;
        RECT 103.800 136.400 104.200 137.200 ;
        RECT 104.600 136.200 104.900 137.500 ;
        RECT 105.400 137.100 105.800 137.200 ;
        RECT 107.000 137.100 107.400 137.200 ;
        RECT 105.400 136.800 107.400 137.100 ;
        RECT 107.000 136.400 107.400 136.800 ;
        RECT 107.800 136.200 108.100 137.500 ;
        RECT 109.400 136.400 109.800 139.900 ;
        RECT 100.500 135.900 101.800 136.200 ;
        RECT 94.100 135.300 96.200 135.600 ;
        RECT 94.100 135.200 94.500 135.300 ;
        RECT 94.900 134.900 95.300 135.000 ;
        RECT 93.400 134.600 95.300 134.900 ;
        RECT 93.400 134.500 93.800 134.600 ;
        RECT 78.200 133.400 78.600 134.200 ;
        RECT 80.900 134.100 81.700 134.200 ;
        RECT 79.800 133.900 81.700 134.100 ;
        RECT 82.200 134.100 82.600 134.200 ;
        RECT 79.800 133.800 81.200 133.900 ;
        RECT 82.200 133.800 83.000 134.100 ;
        RECT 83.700 133.800 85.000 134.200 ;
        RECT 87.400 133.900 92.900 134.200 ;
        RECT 87.400 133.800 88.200 133.900 ;
        RECT 73.400 131.100 73.800 133.100 ;
        RECT 74.200 133.000 76.200 133.100 ;
        RECT 74.200 131.100 74.600 133.000 ;
        RECT 75.800 131.100 76.200 133.000 ;
        RECT 76.900 132.800 77.800 133.100 ;
        RECT 79.800 133.200 80.100 133.800 ;
        RECT 79.800 132.800 80.200 133.200 ;
        RECT 76.900 132.200 77.300 132.800 ;
        RECT 76.600 131.800 77.300 132.200 ;
        RECT 76.900 131.100 77.300 131.800 ;
        RECT 80.800 131.100 81.200 133.800 ;
        RECT 82.600 133.600 83.000 133.800 ;
        RECT 82.300 133.100 84.100 133.300 ;
        RECT 84.600 133.100 84.900 133.800 ;
        RECT 82.200 133.000 84.200 133.100 ;
        RECT 82.200 131.100 82.600 133.000 ;
        RECT 83.800 131.100 84.200 133.000 ;
        RECT 84.600 131.100 85.000 133.100 ;
        RECT 87.000 131.100 87.400 133.500 ;
        RECT 89.500 132.800 89.800 133.900 ;
        RECT 92.300 133.800 92.700 133.900 ;
        RECT 95.800 133.600 96.200 135.300 ;
        RECT 97.500 135.100 97.800 135.900 ;
        RECT 96.600 134.800 97.800 135.100 ;
        RECT 98.200 134.800 98.600 135.600 ;
        RECT 96.600 134.200 96.900 134.800 ;
        RECT 97.500 134.200 97.800 134.800 ;
        RECT 96.600 133.800 97.000 134.200 ;
        RECT 97.400 133.800 97.800 134.200 ;
        RECT 94.300 133.300 96.200 133.600 ;
        RECT 94.300 133.200 94.700 133.300 ;
        RECT 88.600 132.100 89.000 132.500 ;
        RECT 89.400 132.400 89.800 132.800 ;
        RECT 90.300 132.700 90.700 132.800 ;
        RECT 90.300 132.400 91.700 132.700 ;
        RECT 91.400 132.100 91.700 132.400 ;
        RECT 93.400 132.100 93.800 132.500 ;
        RECT 88.600 131.800 89.600 132.100 ;
        RECT 89.200 131.100 89.600 131.800 ;
        RECT 91.400 131.100 91.800 132.100 ;
        RECT 93.400 131.800 94.100 132.100 ;
        RECT 93.500 131.100 94.100 131.800 ;
        RECT 95.800 131.100 96.200 133.300 ;
        RECT 96.600 132.400 97.000 133.200 ;
        RECT 97.500 132.100 97.800 133.800 ;
        RECT 99.700 134.200 100.000 135.900 ;
        RECT 100.500 134.900 100.800 135.900 ;
        RECT 102.200 135.400 102.600 136.200 ;
        RECT 104.600 135.800 105.000 136.200 ;
        RECT 100.300 134.500 100.800 134.900 ;
        RECT 99.700 133.800 100.200 134.200 ;
        RECT 99.700 133.100 100.000 133.800 ;
        RECT 100.500 133.700 100.800 134.500 ;
        RECT 101.300 134.800 101.800 135.200 ;
        RECT 103.000 134.800 103.800 135.200 ;
        RECT 101.300 134.400 101.700 134.800 ;
        RECT 104.600 134.200 104.900 135.800 ;
        RECT 105.400 135.400 105.800 136.200 ;
        RECT 107.800 135.800 108.200 136.200 ;
        RECT 109.300 135.900 109.800 136.400 ;
        RECT 111.000 136.200 111.400 139.900 ;
        RECT 111.800 137.900 112.200 139.900 ;
        RECT 111.900 137.800 112.200 137.900 ;
        RECT 113.400 137.900 113.800 139.900 ;
        RECT 115.800 137.900 116.200 139.900 ;
        RECT 113.400 137.800 113.700 137.900 ;
        RECT 111.900 137.500 113.700 137.800 ;
        RECT 115.900 137.800 116.200 137.900 ;
        RECT 117.400 137.900 117.800 139.900 ;
        RECT 119.000 137.900 119.400 139.900 ;
        RECT 117.400 137.800 117.700 137.900 ;
        RECT 115.900 137.500 117.700 137.800 ;
        RECT 119.100 137.800 119.400 137.900 ;
        RECT 120.600 137.900 121.000 139.900 ;
        RECT 121.400 137.900 121.800 139.900 ;
        RECT 120.600 137.800 120.900 137.900 ;
        RECT 119.100 137.500 120.900 137.800 ;
        RECT 111.900 136.200 112.200 137.500 ;
        RECT 112.600 136.400 113.000 137.200 ;
        RECT 116.600 136.400 117.000 137.200 ;
        RECT 117.400 136.200 117.700 137.500 ;
        RECT 119.800 136.400 120.200 137.200 ;
        RECT 120.600 136.200 120.900 137.500 ;
        RECT 121.500 137.800 121.800 137.900 ;
        RECT 123.000 137.900 123.400 139.900 ;
        RECT 124.600 137.900 125.000 139.900 ;
        RECT 123.000 137.800 123.300 137.900 ;
        RECT 121.500 137.500 123.300 137.800 ;
        RECT 124.700 137.800 125.000 137.900 ;
        RECT 126.200 137.900 126.600 139.900 ;
        RECT 126.200 137.800 126.500 137.900 ;
        RECT 124.700 137.500 126.500 137.800 ;
        RECT 121.500 136.200 121.800 137.500 ;
        RECT 122.200 136.400 122.600 137.200 ;
        RECT 124.700 136.200 125.000 137.500 ;
        RECT 125.400 136.400 125.800 137.200 ;
        RECT 129.100 136.300 129.500 139.900 ;
        RECT 131.000 136.400 131.400 139.900 ;
        RECT 110.100 135.900 111.400 136.200 ;
        RECT 106.200 134.800 107.000 135.200 ;
        RECT 107.800 134.200 108.100 135.800 ;
        RECT 109.300 134.200 109.600 135.900 ;
        RECT 110.100 134.900 110.400 135.900 ;
        RECT 111.800 135.800 112.200 136.200 ;
        RECT 109.900 134.500 110.400 134.900 ;
        RECT 104.100 134.100 104.900 134.200 ;
        RECT 107.300 134.100 108.100 134.200 ;
        RECT 104.000 133.900 104.900 134.100 ;
        RECT 107.200 133.900 108.100 134.100 ;
        RECT 108.600 134.100 109.000 134.200 ;
        RECT 109.300 134.100 109.800 134.200 ;
        RECT 100.500 133.400 101.800 133.700 ;
        RECT 99.700 132.800 100.200 133.100 ;
        RECT 97.400 131.100 97.800 132.100 ;
        RECT 99.800 131.100 100.200 132.800 ;
        RECT 101.400 131.100 101.800 133.400 ;
        RECT 104.000 132.200 104.400 133.900 ;
        RECT 107.200 132.200 107.600 133.900 ;
        RECT 108.600 133.800 109.800 134.100 ;
        RECT 109.300 133.100 109.600 133.800 ;
        RECT 110.100 133.700 110.400 134.500 ;
        RECT 110.900 134.800 111.400 135.200 ;
        RECT 110.900 134.400 111.300 134.800 ;
        RECT 111.900 134.200 112.200 135.800 ;
        RECT 114.200 136.100 114.600 136.200 ;
        RECT 115.000 136.100 115.400 136.200 ;
        RECT 114.200 135.800 115.400 136.100 ;
        RECT 114.200 135.400 114.600 135.800 ;
        RECT 115.000 135.400 115.400 135.800 ;
        RECT 117.400 135.800 117.800 136.200 ;
        RECT 118.200 136.100 118.600 136.200 ;
        RECT 119.000 136.100 119.400 136.200 ;
        RECT 118.200 135.800 119.400 136.100 ;
        RECT 120.600 135.800 121.000 136.200 ;
        RECT 121.400 135.800 121.800 136.200 ;
        RECT 113.000 134.800 113.800 135.200 ;
        RECT 115.800 134.800 116.600 135.200 ;
        RECT 117.400 134.200 117.700 135.800 ;
        RECT 118.200 135.400 118.600 135.800 ;
        RECT 119.000 134.800 119.800 135.200 ;
        RECT 120.600 134.200 120.900 135.800 ;
        RECT 111.900 134.100 112.700 134.200 ;
        RECT 116.900 134.100 117.700 134.200 ;
        RECT 120.100 134.100 120.900 134.200 ;
        RECT 111.900 133.900 112.800 134.100 ;
        RECT 110.100 133.400 111.400 133.700 ;
        RECT 109.300 132.800 109.800 133.100 ;
        RECT 104.000 131.800 105.000 132.200 ;
        RECT 107.200 131.800 108.200 132.200 ;
        RECT 104.000 131.100 104.400 131.800 ;
        RECT 107.200 131.100 107.600 131.800 ;
        RECT 109.400 131.100 109.800 132.800 ;
        RECT 111.000 131.100 111.400 133.400 ;
        RECT 112.400 132.200 112.800 133.900 ;
        RECT 116.800 133.900 117.700 134.100 ;
        RECT 120.000 133.900 120.900 134.100 ;
        RECT 121.500 134.200 121.800 135.800 ;
        RECT 123.800 135.400 124.200 136.200 ;
        RECT 124.600 135.800 125.000 136.200 ;
        RECT 122.600 134.800 123.400 135.200 ;
        RECT 124.700 134.200 125.000 135.800 ;
        RECT 127.000 135.400 127.400 136.200 ;
        RECT 128.600 135.900 129.500 136.300 ;
        RECT 125.800 134.800 126.600 135.200 ;
        RECT 128.700 135.100 129.000 135.900 ;
        RECT 130.900 135.800 131.400 136.400 ;
        RECT 132.600 136.200 133.000 139.900 ;
        RECT 131.700 135.900 133.000 136.200 ;
        RECT 127.800 134.800 129.000 135.100 ;
        RECT 129.400 134.800 129.800 135.600 ;
        RECT 127.800 134.200 128.100 134.800 ;
        RECT 128.700 134.200 129.000 134.800 ;
        RECT 121.500 134.100 122.300 134.200 ;
        RECT 124.700 134.100 125.500 134.200 ;
        RECT 121.500 133.900 122.400 134.100 ;
        RECT 124.700 133.900 125.600 134.100 ;
        RECT 111.800 131.800 112.800 132.200 ;
        RECT 115.800 132.100 116.200 132.200 ;
        RECT 116.800 132.100 117.200 133.900 ;
        RECT 115.800 131.800 117.200 132.100 ;
        RECT 112.400 131.100 112.800 131.800 ;
        RECT 116.800 131.100 117.200 131.800 ;
        RECT 120.000 131.100 120.400 133.900 ;
        RECT 122.000 131.100 122.400 133.900 ;
        RECT 125.200 132.100 125.600 133.900 ;
        RECT 127.800 133.800 128.200 134.200 ;
        RECT 128.600 133.800 129.000 134.200 ;
        RECT 127.800 132.400 128.200 133.200 ;
        RECT 126.200 132.100 126.600 132.200 ;
        RECT 128.700 132.100 129.000 133.800 ;
        RECT 130.900 134.200 131.200 135.800 ;
        RECT 131.700 134.900 132.000 135.900 ;
        RECT 131.500 134.500 132.000 134.900 ;
        RECT 130.900 133.800 131.400 134.200 ;
        RECT 130.900 133.100 131.200 133.800 ;
        RECT 131.700 133.700 132.000 134.500 ;
        RECT 132.500 134.800 133.000 135.200 ;
        RECT 132.500 134.400 132.900 134.800 ;
        RECT 131.700 133.400 133.000 133.700 ;
        RECT 133.400 133.400 133.800 134.200 ;
        RECT 130.900 132.800 131.400 133.100 ;
        RECT 125.200 131.800 126.600 132.100 ;
        RECT 125.200 131.100 125.600 131.800 ;
        RECT 128.600 131.100 129.000 132.100 ;
        RECT 131.000 131.100 131.400 132.800 ;
        RECT 132.600 131.100 133.000 133.400 ;
        RECT 134.200 133.100 134.600 139.900 ;
        RECT 135.000 135.800 135.400 136.600 ;
        RECT 137.100 135.900 138.100 139.900 ;
        RECT 141.800 136.800 142.200 137.200 ;
        RECT 141.800 136.200 142.100 136.800 ;
        RECT 142.500 136.200 142.900 139.900 ;
        RECT 145.900 136.200 146.300 139.900 ;
        RECT 146.600 136.800 147.000 137.200 ;
        RECT 146.700 136.200 147.000 136.800 ;
        RECT 141.400 135.900 142.100 136.200 ;
        RECT 136.600 134.400 137.000 135.200 ;
        RECT 137.400 134.200 137.700 135.900 ;
        RECT 141.400 135.800 141.800 135.900 ;
        RECT 142.400 135.800 143.400 136.200 ;
        RECT 145.900 135.900 146.400 136.200 ;
        RECT 146.700 135.900 147.400 136.200 ;
        RECT 138.200 134.400 138.600 135.200 ;
        RECT 135.800 134.100 136.200 134.200 ;
        RECT 137.400 134.100 137.800 134.200 ;
        RECT 135.800 133.800 136.600 134.100 ;
        RECT 137.400 133.800 138.600 134.100 ;
        RECT 139.000 133.800 139.400 134.600 ;
        RECT 142.400 134.200 142.700 135.800 ;
        RECT 143.000 134.400 143.400 135.200 ;
        RECT 145.400 134.400 145.800 135.200 ;
        RECT 146.100 134.200 146.400 135.900 ;
        RECT 147.000 135.800 147.400 135.900 ;
        RECT 147.800 136.100 148.200 139.900 ;
        RECT 148.600 136.100 149.000 136.200 ;
        RECT 147.800 135.800 149.000 136.100 ;
        RECT 141.400 133.800 142.700 134.200 ;
        RECT 143.800 134.100 144.200 134.200 ;
        RECT 143.400 133.800 144.200 134.100 ;
        RECT 144.600 134.100 145.000 134.200 ;
        RECT 144.600 133.800 145.400 134.100 ;
        RECT 146.100 133.800 147.400 134.200 ;
        RECT 136.200 133.600 136.600 133.800 ;
        RECT 135.900 133.100 137.700 133.300 ;
        RECT 138.300 133.100 138.600 133.800 ;
        RECT 141.500 133.100 141.800 133.800 ;
        RECT 143.400 133.600 143.800 133.800 ;
        RECT 145.000 133.600 145.400 133.800 ;
        RECT 142.300 133.100 144.100 133.300 ;
        RECT 144.700 133.100 146.500 133.300 ;
        RECT 147.000 133.100 147.300 133.800 ;
        RECT 134.200 132.800 135.100 133.100 ;
        RECT 134.700 132.200 135.100 132.800 ;
        RECT 135.800 133.000 137.800 133.100 ;
        RECT 134.700 131.800 135.400 132.200 ;
        RECT 134.700 131.100 135.100 131.800 ;
        RECT 135.800 131.100 136.200 133.000 ;
        RECT 137.400 131.400 137.800 133.000 ;
        RECT 138.200 131.700 138.600 133.100 ;
        RECT 139.000 131.400 139.400 133.100 ;
        RECT 137.400 131.100 139.400 131.400 ;
        RECT 141.400 131.100 141.800 133.100 ;
        RECT 142.200 133.000 144.200 133.100 ;
        RECT 142.200 131.100 142.600 133.000 ;
        RECT 143.800 131.100 144.200 133.000 ;
        RECT 144.600 133.000 146.600 133.100 ;
        RECT 144.600 131.100 145.000 133.000 ;
        RECT 146.200 131.100 146.600 133.000 ;
        RECT 147.000 131.100 147.400 133.100 ;
        RECT 147.800 131.100 148.200 135.800 ;
        RECT 150.200 135.600 150.600 139.900 ;
        RECT 151.800 135.600 152.200 139.900 ;
        RECT 153.700 139.200 154.100 139.900 ;
        RECT 153.400 138.800 154.100 139.200 ;
        RECT 153.700 136.300 154.100 138.800 ;
        RECT 156.200 136.800 156.600 137.200 ;
        RECT 153.700 135.900 154.600 136.300 ;
        RECT 156.200 136.200 156.500 136.800 ;
        RECT 156.900 136.200 157.300 139.900 ;
        RECT 155.800 135.900 156.500 136.200 ;
        RECT 156.800 135.900 157.300 136.200 ;
        RECT 150.200 135.200 152.200 135.600 ;
        RECT 150.200 133.800 150.600 135.200 ;
        RECT 153.400 134.800 153.800 135.600 ;
        RECT 154.200 134.200 154.500 135.900 ;
        RECT 155.800 135.800 156.200 135.900 ;
        RECT 156.800 134.200 157.100 135.900 ;
        RECT 157.400 135.100 157.800 135.200 ;
        RECT 158.200 135.100 158.600 135.200 ;
        RECT 157.400 134.800 158.600 135.100 ;
        RECT 157.400 134.400 157.800 134.800 ;
        RECT 152.600 134.100 153.000 134.200 ;
        RECT 153.400 134.100 153.800 134.200 ;
        RECT 152.600 133.800 153.800 134.100 ;
        RECT 154.200 133.800 154.600 134.200 ;
        RECT 155.800 133.800 157.100 134.200 ;
        RECT 158.200 134.100 158.600 134.200 ;
        RECT 157.800 133.800 158.600 134.100 ;
        RECT 150.200 133.400 152.200 133.800 ;
        RECT 152.600 133.400 153.000 133.800 ;
        RECT 148.600 132.400 149.000 133.200 ;
        RECT 150.200 131.100 150.600 133.400 ;
        RECT 151.800 131.100 152.200 133.400 ;
        RECT 154.200 132.100 154.500 133.800 ;
        RECT 155.000 133.100 155.400 133.200 ;
        RECT 155.900 133.100 156.200 133.800 ;
        RECT 157.800 133.600 158.200 133.800 ;
        RECT 159.000 133.400 159.400 134.200 ;
        RECT 156.700 133.100 158.500 133.300 ;
        RECT 159.800 133.100 160.200 139.900 ;
        RECT 160.600 135.800 161.000 136.600 ;
        RECT 161.400 133.400 161.800 134.200 ;
        RECT 162.200 134.100 162.600 139.900 ;
        RECT 164.600 137.900 165.000 139.900 ;
        RECT 164.700 137.800 165.000 137.900 ;
        RECT 166.200 137.900 166.600 139.900 ;
        RECT 166.200 137.800 166.500 137.900 ;
        RECT 164.700 137.500 166.500 137.800 ;
        RECT 163.000 135.800 163.400 136.600 ;
        RECT 165.400 136.400 165.800 137.200 ;
        RECT 166.200 136.200 166.500 137.500 ;
        RECT 167.400 136.800 167.800 137.200 ;
        RECT 167.400 136.200 167.700 136.800 ;
        RECT 168.100 136.200 168.500 139.900 ;
        RECT 171.500 136.200 171.900 139.900 ;
        RECT 172.200 136.800 172.600 137.200 ;
        RECT 172.300 136.200 172.600 136.800 ;
        RECT 174.700 136.200 175.100 139.900 ;
        RECT 175.400 136.800 175.800 137.200 ;
        RECT 175.500 136.200 175.800 136.800 ;
        RECT 163.800 135.400 164.200 136.200 ;
        RECT 166.200 135.800 166.600 136.200 ;
        RECT 167.000 135.900 167.700 136.200 ;
        RECT 168.000 135.900 168.500 136.200 ;
        RECT 167.000 135.800 167.400 135.900 ;
        RECT 163.000 134.800 163.400 135.200 ;
        RECT 164.600 134.800 165.400 135.200 ;
        RECT 163.000 134.100 163.300 134.800 ;
        RECT 166.200 134.200 166.500 135.800 ;
        RECT 168.000 134.200 168.300 135.900 ;
        RECT 171.000 135.800 172.000 136.200 ;
        RECT 172.300 135.900 173.000 136.200 ;
        RECT 174.700 135.900 175.200 136.200 ;
        RECT 175.500 135.900 176.200 136.200 ;
        RECT 172.600 135.800 173.000 135.900 ;
        RECT 168.600 135.100 169.000 135.200 ;
        RECT 170.200 135.100 170.600 135.200 ;
        RECT 168.600 134.800 170.600 135.100 ;
        RECT 168.600 134.400 169.000 134.800 ;
        RECT 171.000 134.400 171.400 135.200 ;
        RECT 171.700 134.200 172.000 135.800 ;
        RECT 174.200 134.400 174.600 135.200 ;
        RECT 174.900 134.200 175.200 135.900 ;
        RECT 175.800 135.800 176.200 135.900 ;
        RECT 176.600 135.800 177.000 136.600 ;
        RECT 175.800 135.100 176.100 135.800 ;
        RECT 177.400 135.100 177.800 139.900 ;
        RECT 175.800 134.800 177.800 135.100 ;
        RECT 165.700 134.100 166.600 134.200 ;
        RECT 162.200 133.800 163.300 134.100 ;
        RECT 165.600 133.800 166.600 134.100 ;
        RECT 167.000 133.800 168.300 134.200 ;
        RECT 169.400 134.100 169.800 134.200 ;
        RECT 169.000 133.800 169.800 134.100 ;
        RECT 170.200 134.100 170.600 134.200 ;
        RECT 170.200 133.800 171.000 134.100 ;
        RECT 171.700 133.800 173.000 134.200 ;
        RECT 173.400 134.100 173.800 134.200 ;
        RECT 173.400 133.800 174.200 134.100 ;
        RECT 174.900 133.800 176.200 134.200 ;
        RECT 162.200 133.100 162.600 133.800 ;
        RECT 155.000 132.800 156.200 133.100 ;
        RECT 155.000 132.400 155.400 132.800 ;
        RECT 154.200 131.100 154.600 132.100 ;
        RECT 155.800 131.100 156.200 132.800 ;
        RECT 156.600 133.000 158.600 133.100 ;
        RECT 156.600 131.100 157.000 133.000 ;
        RECT 158.200 131.100 158.600 133.000 ;
        RECT 159.800 132.800 160.700 133.100 ;
        RECT 162.200 132.800 163.100 133.100 ;
        RECT 160.300 132.200 160.700 132.800 ;
        RECT 160.300 131.800 161.000 132.200 ;
        RECT 160.300 131.100 160.700 131.800 ;
        RECT 162.700 131.100 163.100 132.800 ;
        RECT 165.600 131.100 166.000 133.800 ;
        RECT 167.100 133.100 167.400 133.800 ;
        RECT 169.000 133.600 169.400 133.800 ;
        RECT 170.600 133.600 171.000 133.800 ;
        RECT 167.900 133.100 169.700 133.300 ;
        RECT 170.300 133.100 172.100 133.300 ;
        RECT 172.600 133.100 172.900 133.800 ;
        RECT 173.800 133.600 174.200 133.800 ;
        RECT 173.500 133.100 175.300 133.300 ;
        RECT 175.800 133.100 176.100 133.800 ;
        RECT 177.400 133.100 177.800 134.800 ;
        RECT 179.800 135.100 180.200 139.900 ;
        RECT 182.500 139.200 182.900 139.900 ;
        RECT 182.500 138.800 183.400 139.200 ;
        RECT 181.800 136.800 182.200 137.200 ;
        RECT 180.600 135.800 181.000 136.600 ;
        RECT 181.800 136.200 182.100 136.800 ;
        RECT 182.500 136.200 182.900 138.800 ;
        RECT 181.400 135.900 182.100 136.200 ;
        RECT 182.400 135.900 182.900 136.200 ;
        RECT 181.400 135.800 181.800 135.900 ;
        RECT 181.400 135.100 181.700 135.800 ;
        RECT 179.800 134.800 181.700 135.100 ;
        RECT 178.200 133.400 178.600 134.200 ;
        RECT 179.000 133.400 179.400 134.200 ;
        RECT 167.000 131.100 167.400 133.100 ;
        RECT 167.800 133.000 169.800 133.100 ;
        RECT 167.800 131.100 168.200 133.000 ;
        RECT 169.400 131.100 169.800 133.000 ;
        RECT 170.200 133.000 172.200 133.100 ;
        RECT 170.200 131.100 170.600 133.000 ;
        RECT 171.800 131.100 172.200 133.000 ;
        RECT 172.600 131.100 173.000 133.100 ;
        RECT 173.400 133.000 175.400 133.100 ;
        RECT 173.400 131.100 173.800 133.000 ;
        RECT 175.000 131.100 175.400 133.000 ;
        RECT 175.800 131.100 176.200 133.100 ;
        RECT 176.900 132.800 177.800 133.100 ;
        RECT 179.800 133.100 180.200 134.800 ;
        RECT 182.400 134.200 182.700 135.900 ;
        RECT 184.600 135.800 185.000 137.200 ;
        RECT 183.000 134.400 183.400 135.200 ;
        RECT 181.400 133.800 182.700 134.200 ;
        RECT 183.800 134.100 184.200 134.200 ;
        RECT 183.400 133.800 184.200 134.100 ;
        RECT 181.500 133.100 181.800 133.800 ;
        RECT 183.400 133.600 183.800 133.800 ;
        RECT 182.300 133.100 184.100 133.300 ;
        RECT 185.400 133.100 185.800 139.900 ;
        RECT 188.600 135.600 189.000 139.900 ;
        RECT 190.700 137.900 191.300 139.900 ;
        RECT 193.000 137.900 193.400 139.900 ;
        RECT 195.200 138.200 195.600 139.900 ;
        RECT 195.200 137.900 196.200 138.200 ;
        RECT 191.000 137.500 191.400 137.900 ;
        RECT 193.100 137.600 193.400 137.900 ;
        RECT 192.700 137.300 194.500 137.600 ;
        RECT 195.800 137.500 196.200 137.900 ;
        RECT 192.700 137.200 193.100 137.300 ;
        RECT 194.100 137.200 194.500 137.300 ;
        RECT 190.600 136.600 191.300 137.000 ;
        RECT 191.000 136.100 191.300 136.600 ;
        RECT 192.100 136.500 193.200 136.800 ;
        RECT 192.100 136.400 192.500 136.500 ;
        RECT 191.000 135.800 192.200 136.100 ;
        RECT 188.600 135.300 190.700 135.600 ;
        RECT 186.200 133.400 186.600 134.200 ;
        RECT 188.600 133.600 189.000 135.300 ;
        RECT 190.300 135.200 190.700 135.300 ;
        RECT 189.500 134.900 189.900 135.000 ;
        RECT 189.500 134.600 191.400 134.900 ;
        RECT 191.000 134.500 191.400 134.600 ;
        RECT 191.900 134.200 192.200 135.800 ;
        RECT 192.900 135.900 193.200 136.500 ;
        RECT 193.500 136.500 193.900 136.600 ;
        RECT 195.800 136.500 196.200 136.600 ;
        RECT 193.500 136.200 196.200 136.500 ;
        RECT 192.900 135.700 195.300 135.900 ;
        RECT 197.400 135.700 197.800 139.900 ;
        RECT 198.600 136.800 199.000 137.200 ;
        RECT 198.600 136.200 198.900 136.800 ;
        RECT 199.300 136.200 199.700 139.900 ;
        RECT 198.200 135.900 198.900 136.200 ;
        RECT 199.200 135.900 199.700 136.200 ;
        RECT 198.200 135.800 198.600 135.900 ;
        RECT 192.900 135.600 197.800 135.700 ;
        RECT 194.900 135.500 197.800 135.600 ;
        RECT 195.000 135.400 197.800 135.500 ;
        RECT 192.600 135.100 193.000 135.200 ;
        RECT 194.200 135.100 194.600 135.200 ;
        RECT 192.600 134.800 196.700 135.100 ;
        RECT 196.300 134.700 196.700 134.800 ;
        RECT 195.500 134.200 195.900 134.300 ;
        RECT 199.200 134.200 199.500 135.900 ;
        RECT 199.800 134.400 200.200 135.200 ;
        RECT 191.900 133.900 197.400 134.200 ;
        RECT 192.100 133.800 192.500 133.900 ;
        RECT 195.000 133.800 195.400 133.900 ;
        RECT 196.600 133.800 197.400 133.900 ;
        RECT 198.200 133.800 199.500 134.200 ;
        RECT 200.600 134.100 201.000 134.200 ;
        RECT 200.200 133.800 201.000 134.100 ;
        RECT 179.800 132.800 180.700 133.100 ;
        RECT 176.900 131.100 177.300 132.800 ;
        RECT 180.300 131.100 180.700 132.800 ;
        RECT 181.400 131.100 181.800 133.100 ;
        RECT 182.200 133.000 184.200 133.100 ;
        RECT 182.200 131.100 182.600 133.000 ;
        RECT 183.800 131.100 184.200 133.000 ;
        RECT 184.900 132.800 185.800 133.100 ;
        RECT 188.600 133.300 190.500 133.600 ;
        RECT 184.900 132.200 185.300 132.800 ;
        RECT 184.900 131.800 185.800 132.200 ;
        RECT 184.900 131.100 185.300 131.800 ;
        RECT 188.600 131.100 189.000 133.300 ;
        RECT 190.100 133.200 190.500 133.300 ;
        RECT 195.000 132.800 195.300 133.800 ;
        RECT 194.100 132.700 194.500 132.800 ;
        RECT 191.000 132.100 191.400 132.500 ;
        RECT 193.100 132.400 194.500 132.700 ;
        RECT 195.000 132.400 195.400 132.800 ;
        RECT 193.100 132.100 193.400 132.400 ;
        RECT 195.800 132.100 196.200 132.500 ;
        RECT 190.700 131.800 191.400 132.100 ;
        RECT 190.700 131.100 191.300 131.800 ;
        RECT 193.000 131.100 193.400 132.100 ;
        RECT 195.200 131.800 196.200 132.100 ;
        RECT 195.200 131.100 195.600 131.800 ;
        RECT 197.400 131.100 197.800 133.500 ;
        RECT 198.300 133.100 198.600 133.800 ;
        RECT 200.200 133.600 200.600 133.800 ;
        RECT 199.100 133.100 200.900 133.300 ;
        RECT 198.200 131.100 198.600 133.100 ;
        RECT 199.000 133.000 201.000 133.100 ;
        RECT 199.000 131.100 199.400 133.000 ;
        RECT 200.600 131.100 201.000 133.000 ;
        RECT 201.400 131.100 201.800 139.900 ;
        RECT 203.800 135.100 204.200 139.900 ;
        RECT 205.800 136.800 206.200 137.200 ;
        RECT 204.600 135.800 205.000 136.600 ;
        RECT 205.800 136.200 206.100 136.800 ;
        RECT 206.500 136.200 206.900 139.900 ;
        RECT 205.400 135.900 206.100 136.200 ;
        RECT 205.400 135.800 205.800 135.900 ;
        RECT 206.400 135.800 207.400 136.200 ;
        RECT 205.400 135.100 205.700 135.800 ;
        RECT 203.800 134.800 205.700 135.100 ;
        RECT 203.000 134.100 203.400 134.200 ;
        RECT 202.200 133.800 203.400 134.100 ;
        RECT 202.200 133.200 202.500 133.800 ;
        RECT 203.000 133.400 203.400 133.800 ;
        RECT 202.200 132.400 202.600 133.200 ;
        RECT 203.800 133.100 204.200 134.800 ;
        RECT 206.400 134.200 206.700 135.800 ;
        RECT 208.600 135.600 209.000 139.900 ;
        RECT 210.700 137.900 211.300 139.900 ;
        RECT 213.000 137.900 213.400 139.900 ;
        RECT 215.200 138.200 215.600 139.900 ;
        RECT 215.200 137.900 216.200 138.200 ;
        RECT 211.000 137.500 211.400 137.900 ;
        RECT 213.100 137.600 213.400 137.900 ;
        RECT 212.700 137.300 214.500 137.600 ;
        RECT 215.800 137.500 216.200 137.900 ;
        RECT 212.700 137.200 213.100 137.300 ;
        RECT 214.100 137.200 214.500 137.300 ;
        RECT 210.600 136.600 211.300 137.000 ;
        RECT 211.000 136.100 211.300 136.600 ;
        RECT 212.100 136.500 213.200 136.800 ;
        RECT 212.100 136.400 212.500 136.500 ;
        RECT 211.000 135.800 212.200 136.100 ;
        RECT 208.600 135.300 210.700 135.600 ;
        RECT 207.000 134.400 207.400 135.200 ;
        RECT 205.400 133.800 206.700 134.200 ;
        RECT 207.800 134.100 208.200 134.200 ;
        RECT 207.400 133.800 208.200 134.100 ;
        RECT 205.500 133.100 205.800 133.800 ;
        RECT 207.400 133.600 207.800 133.800 ;
        RECT 208.600 133.600 209.000 135.300 ;
        RECT 210.300 135.200 210.700 135.300 ;
        RECT 209.500 134.900 209.900 135.000 ;
        RECT 209.500 134.600 211.400 134.900 ;
        RECT 211.000 134.500 211.400 134.600 ;
        RECT 211.900 134.200 212.200 135.800 ;
        RECT 212.900 135.900 213.200 136.500 ;
        RECT 213.500 136.500 213.900 136.600 ;
        RECT 215.800 136.500 216.200 136.600 ;
        RECT 213.500 136.200 216.200 136.500 ;
        RECT 212.900 135.700 215.300 135.900 ;
        RECT 217.400 135.700 217.800 139.900 ;
        RECT 212.900 135.600 217.800 135.700 ;
        RECT 214.900 135.500 217.800 135.600 ;
        RECT 215.000 135.400 217.800 135.500 ;
        RECT 218.200 135.700 218.600 139.900 ;
        RECT 220.400 138.200 220.800 139.900 ;
        RECT 219.800 137.900 220.800 138.200 ;
        RECT 222.600 137.900 223.000 139.900 ;
        RECT 224.700 137.900 225.300 139.900 ;
        RECT 219.800 137.500 220.200 137.900 ;
        RECT 222.600 137.600 222.900 137.900 ;
        RECT 221.500 137.300 223.300 137.600 ;
        RECT 224.600 137.500 225.000 137.900 ;
        RECT 221.500 137.200 221.900 137.300 ;
        RECT 222.900 137.200 223.300 137.300 ;
        RECT 219.800 136.500 220.200 136.600 ;
        RECT 222.100 136.500 222.500 136.600 ;
        RECT 219.800 136.200 222.500 136.500 ;
        RECT 222.800 136.500 223.900 136.800 ;
        RECT 222.800 135.900 223.100 136.500 ;
        RECT 223.500 136.400 223.900 136.500 ;
        RECT 224.700 136.600 225.400 137.000 ;
        RECT 224.700 136.100 225.000 136.600 ;
        RECT 220.700 135.700 223.100 135.900 ;
        RECT 218.200 135.600 223.100 135.700 ;
        RECT 223.800 135.800 225.000 136.100 ;
        RECT 218.200 135.500 221.100 135.600 ;
        RECT 218.200 135.400 221.000 135.500 ;
        RECT 223.800 135.200 224.100 135.800 ;
        RECT 227.000 135.600 227.400 139.900 ;
        RECT 227.800 136.200 228.200 139.900 ;
        RECT 227.800 135.900 228.900 136.200 ;
        RECT 225.300 135.300 227.400 135.600 ;
        RECT 225.300 135.200 225.700 135.300 ;
        RECT 214.200 135.100 214.600 135.200 ;
        RECT 221.400 135.100 221.800 135.200 ;
        RECT 214.200 134.800 216.700 135.100 ;
        RECT 216.300 134.700 216.700 134.800 ;
        RECT 219.300 134.800 221.800 135.100 ;
        RECT 223.800 134.800 224.200 135.200 ;
        RECT 227.000 135.100 227.400 135.300 ;
        RECT 228.600 135.600 228.900 135.900 ;
        RECT 228.600 135.200 229.200 135.600 ;
        RECT 227.800 135.100 228.200 135.200 ;
        RECT 226.100 134.900 226.500 135.000 ;
        RECT 219.300 134.700 219.700 134.800 ;
        RECT 215.500 134.200 215.900 134.300 ;
        RECT 220.100 134.200 220.500 134.300 ;
        RECT 223.800 134.200 224.100 134.800 ;
        RECT 224.600 134.600 226.500 134.900 ;
        RECT 227.000 134.800 228.200 135.100 ;
        RECT 224.600 134.500 225.000 134.600 ;
        RECT 211.900 134.100 217.400 134.200 ;
        RECT 218.600 134.100 224.100 134.200 ;
        RECT 211.900 133.900 224.100 134.100 ;
        RECT 212.100 133.800 212.500 133.900 ;
        RECT 213.400 133.800 213.800 133.900 ;
        RECT 208.600 133.300 210.500 133.600 ;
        RECT 206.300 133.100 208.100 133.300 ;
        RECT 203.800 132.800 204.700 133.100 ;
        RECT 204.300 131.100 204.700 132.800 ;
        RECT 205.400 131.100 205.800 133.100 ;
        RECT 206.200 133.000 208.200 133.100 ;
        RECT 206.200 131.100 206.600 133.000 ;
        RECT 207.800 131.100 208.200 133.000 ;
        RECT 208.600 131.100 209.000 133.300 ;
        RECT 210.100 133.200 210.500 133.300 ;
        RECT 215.000 132.800 215.300 133.900 ;
        RECT 216.600 133.800 219.400 133.900 ;
        RECT 214.100 132.700 214.500 132.800 ;
        RECT 211.000 132.100 211.400 132.500 ;
        RECT 213.100 132.400 214.500 132.700 ;
        RECT 215.000 132.400 215.400 132.800 ;
        RECT 213.100 132.100 213.400 132.400 ;
        RECT 215.800 132.100 216.200 132.500 ;
        RECT 210.700 131.800 211.400 132.100 ;
        RECT 210.700 131.100 211.300 131.800 ;
        RECT 213.000 131.100 213.400 132.100 ;
        RECT 215.200 131.800 216.200 132.100 ;
        RECT 215.200 131.100 215.600 131.800 ;
        RECT 217.400 131.100 217.800 133.500 ;
        RECT 218.200 131.100 218.600 133.500 ;
        RECT 220.700 132.800 221.000 133.900 ;
        RECT 223.500 133.800 223.900 133.900 ;
        RECT 227.000 133.600 227.400 134.800 ;
        RECT 227.800 134.400 228.200 134.800 ;
        RECT 228.600 133.700 228.900 135.200 ;
        RECT 225.500 133.300 227.400 133.600 ;
        RECT 225.500 133.200 225.900 133.300 ;
        RECT 219.800 132.100 220.200 132.500 ;
        RECT 220.600 132.400 221.000 132.800 ;
        RECT 221.500 132.700 221.900 132.800 ;
        RECT 221.500 132.400 222.900 132.700 ;
        RECT 222.600 132.100 222.900 132.400 ;
        RECT 224.600 132.100 225.000 132.500 ;
        RECT 219.800 131.800 220.800 132.100 ;
        RECT 220.400 131.100 220.800 131.800 ;
        RECT 222.600 131.100 223.000 132.100 ;
        RECT 224.600 131.800 225.300 132.100 ;
        RECT 224.700 131.100 225.300 131.800 ;
        RECT 227.000 131.100 227.400 133.300 ;
        RECT 227.800 133.400 228.900 133.700 ;
        RECT 227.800 131.100 228.200 133.400 ;
        RECT 0.600 127.900 1.000 129.900 ;
        RECT 1.400 128.000 1.800 129.900 ;
        RECT 3.000 128.000 3.400 129.900 ;
        RECT 1.400 127.900 3.400 128.000 ;
        RECT 0.700 127.200 1.000 127.900 ;
        RECT 1.500 127.700 3.300 127.900 ;
        RECT 3.800 127.700 4.200 129.900 ;
        RECT 5.900 129.200 6.500 129.900 ;
        RECT 5.900 128.900 6.600 129.200 ;
        RECT 8.200 128.900 8.600 129.900 ;
        RECT 10.400 129.200 10.800 129.900 ;
        RECT 10.400 128.900 11.400 129.200 ;
        RECT 6.200 128.500 6.600 128.900 ;
        RECT 8.300 128.600 8.600 128.900 ;
        RECT 8.300 128.300 9.700 128.600 ;
        RECT 9.300 128.200 9.700 128.300 ;
        RECT 10.200 128.200 10.600 128.600 ;
        RECT 11.000 128.500 11.400 128.900 ;
        RECT 5.300 127.700 5.700 127.800 ;
        RECT 3.800 127.400 5.700 127.700 ;
        RECT 2.600 127.200 3.000 127.400 ;
        RECT 0.600 126.800 1.900 127.200 ;
        RECT 2.600 126.900 3.400 127.200 ;
        RECT 3.000 126.800 3.400 126.900 ;
        RECT 1.600 125.200 1.900 126.800 ;
        RECT 2.200 125.800 2.600 126.600 ;
        RECT 3.800 125.700 4.200 127.400 ;
        RECT 7.300 127.100 7.700 127.200 ;
        RECT 10.200 127.100 10.500 128.200 ;
        RECT 12.600 127.500 13.000 129.900 ;
        RECT 13.400 127.800 13.800 128.600 ;
        RECT 11.800 127.100 12.600 127.200 ;
        RECT 7.100 126.800 12.600 127.100 ;
        RECT 6.200 126.400 6.600 126.500 ;
        RECT 4.700 126.100 6.600 126.400 ;
        RECT 4.700 126.000 5.100 126.100 ;
        RECT 5.500 125.700 5.900 125.800 ;
        RECT 3.800 125.400 5.900 125.700 ;
        RECT 0.600 125.100 1.000 125.200 ;
        RECT 0.600 124.800 1.300 125.100 ;
        RECT 1.600 124.800 2.600 125.200 ;
        RECT 1.000 124.200 1.300 124.800 ;
        RECT 1.000 123.800 1.400 124.200 ;
        RECT 1.700 121.100 2.100 124.800 ;
        RECT 3.800 121.100 4.200 125.400 ;
        RECT 7.100 125.200 7.400 126.800 ;
        RECT 10.700 126.700 11.100 126.800 ;
        RECT 11.500 126.200 11.900 126.300 ;
        RECT 9.400 125.900 11.900 126.200 ;
        RECT 9.400 125.800 9.800 125.900 ;
        RECT 10.200 125.500 13.000 125.600 ;
        RECT 10.100 125.400 13.000 125.500 ;
        RECT 6.200 124.900 7.400 125.200 ;
        RECT 8.100 125.300 13.000 125.400 ;
        RECT 8.100 125.100 10.500 125.300 ;
        RECT 6.200 124.400 6.500 124.900 ;
        RECT 5.800 124.000 6.500 124.400 ;
        RECT 7.300 124.500 7.700 124.600 ;
        RECT 8.100 124.500 8.400 125.100 ;
        RECT 7.300 124.200 8.400 124.500 ;
        RECT 8.700 124.500 11.400 124.800 ;
        RECT 8.700 124.400 9.100 124.500 ;
        RECT 11.000 124.400 11.400 124.500 ;
        RECT 7.900 123.700 8.300 123.800 ;
        RECT 9.300 123.700 9.700 123.800 ;
        RECT 6.200 123.100 6.600 123.500 ;
        RECT 7.900 123.400 9.700 123.700 ;
        RECT 8.300 123.100 8.600 123.400 ;
        RECT 11.000 123.100 11.400 123.500 ;
        RECT 5.900 121.100 6.500 123.100 ;
        RECT 8.200 121.100 8.600 123.100 ;
        RECT 10.400 122.800 11.400 123.100 ;
        RECT 10.400 121.100 10.800 122.800 ;
        RECT 12.600 121.100 13.000 125.300 ;
        RECT 14.200 121.100 14.600 129.900 ;
        RECT 15.000 127.500 15.400 129.900 ;
        RECT 17.200 129.200 17.600 129.900 ;
        RECT 16.600 128.900 17.600 129.200 ;
        RECT 19.400 128.900 19.800 129.900 ;
        RECT 21.500 129.200 22.100 129.900 ;
        RECT 21.400 128.900 22.100 129.200 ;
        RECT 16.600 128.500 17.000 128.900 ;
        RECT 19.400 128.600 19.700 128.900 ;
        RECT 17.400 128.200 17.800 128.600 ;
        RECT 18.300 128.300 19.700 128.600 ;
        RECT 21.400 128.500 21.800 128.900 ;
        RECT 18.300 128.200 18.700 128.300 ;
        RECT 15.400 127.100 16.200 127.200 ;
        RECT 17.500 127.100 17.800 128.200 ;
        RECT 22.300 127.700 22.700 127.800 ;
        RECT 23.800 127.700 24.200 129.900 ;
        RECT 24.600 127.800 25.000 128.600 ;
        RECT 22.300 127.400 24.200 127.700 ;
        RECT 18.200 127.100 18.600 127.200 ;
        RECT 20.300 127.100 20.700 127.200 ;
        RECT 15.400 126.800 20.900 127.100 ;
        RECT 16.900 126.700 17.300 126.800 ;
        RECT 16.100 126.200 16.500 126.300 ;
        RECT 16.100 126.100 18.600 126.200 ;
        RECT 19.000 126.100 19.400 126.200 ;
        RECT 16.100 125.900 19.400 126.100 ;
        RECT 18.200 125.800 19.400 125.900 ;
        RECT 15.000 125.500 17.800 125.600 ;
        RECT 15.000 125.400 17.900 125.500 ;
        RECT 15.000 125.300 19.900 125.400 ;
        RECT 15.000 121.100 15.400 125.300 ;
        RECT 17.500 125.100 19.900 125.300 ;
        RECT 16.600 124.500 19.300 124.800 ;
        RECT 16.600 124.400 17.000 124.500 ;
        RECT 18.900 124.400 19.300 124.500 ;
        RECT 19.600 124.500 19.900 125.100 ;
        RECT 20.600 125.200 20.900 126.800 ;
        RECT 21.400 126.400 21.800 126.500 ;
        RECT 21.400 126.100 23.300 126.400 ;
        RECT 22.900 126.000 23.300 126.100 ;
        RECT 22.100 125.700 22.500 125.800 ;
        RECT 23.800 125.700 24.200 127.400 ;
        RECT 22.100 125.400 24.200 125.700 ;
        RECT 20.600 124.900 21.800 125.200 ;
        RECT 20.300 124.500 20.700 124.600 ;
        RECT 19.600 124.200 20.700 124.500 ;
        RECT 21.500 124.400 21.800 124.900 ;
        RECT 21.500 124.000 22.200 124.400 ;
        RECT 18.300 123.700 18.700 123.800 ;
        RECT 19.700 123.700 20.100 123.800 ;
        RECT 16.600 123.100 17.000 123.500 ;
        RECT 18.300 123.400 20.100 123.700 ;
        RECT 19.400 123.100 19.700 123.400 ;
        RECT 21.400 123.100 21.800 123.500 ;
        RECT 16.600 122.800 17.600 123.100 ;
        RECT 17.200 121.100 17.600 122.800 ;
        RECT 19.400 121.100 19.800 123.100 ;
        RECT 21.500 121.100 22.100 123.100 ;
        RECT 23.800 121.100 24.200 125.400 ;
        RECT 25.400 121.100 25.800 129.900 ;
        RECT 26.200 128.000 26.600 129.900 ;
        RECT 27.800 128.000 28.200 129.900 ;
        RECT 26.200 127.900 28.200 128.000 ;
        RECT 28.600 127.900 29.000 129.900 ;
        RECT 29.400 127.900 29.800 129.900 ;
        RECT 30.200 128.000 30.600 129.900 ;
        RECT 31.800 128.000 32.200 129.900 ;
        RECT 30.200 127.900 32.200 128.000 ;
        RECT 26.300 127.700 28.100 127.900 ;
        RECT 26.600 127.200 27.000 127.400 ;
        RECT 28.600 127.200 28.900 127.900 ;
        RECT 29.500 127.200 29.800 127.900 ;
        RECT 30.300 127.700 32.100 127.900 ;
        RECT 32.600 127.500 33.000 129.900 ;
        RECT 34.800 129.200 35.200 129.900 ;
        RECT 34.200 128.900 35.200 129.200 ;
        RECT 37.000 128.900 37.400 129.900 ;
        RECT 39.100 129.200 39.700 129.900 ;
        RECT 39.000 128.900 39.700 129.200 ;
        RECT 41.400 129.100 41.800 129.900 ;
        RECT 42.200 129.100 42.600 129.200 ;
        RECT 34.200 128.500 34.600 128.900 ;
        RECT 37.000 128.600 37.300 128.900 ;
        RECT 35.000 128.200 35.400 128.600 ;
        RECT 35.900 128.300 37.300 128.600 ;
        RECT 39.000 128.500 39.400 128.900 ;
        RECT 41.400 128.800 42.600 129.100 ;
        RECT 35.900 128.200 36.300 128.300 ;
        RECT 31.400 127.200 31.800 127.400 ;
        RECT 26.200 126.900 27.000 127.200 ;
        RECT 26.200 126.800 26.600 126.900 ;
        RECT 27.700 126.800 29.000 127.200 ;
        RECT 29.400 126.800 30.700 127.200 ;
        RECT 31.400 126.900 32.200 127.200 ;
        RECT 31.800 126.800 32.200 126.900 ;
        RECT 33.000 127.100 33.800 127.200 ;
        RECT 35.100 127.100 35.400 128.200 ;
        RECT 39.900 127.700 40.300 127.800 ;
        RECT 41.400 127.700 41.800 128.800 ;
        RECT 39.900 127.400 41.800 127.700 ;
        RECT 37.900 127.100 38.300 127.200 ;
        RECT 33.000 126.800 38.500 127.100 ;
        RECT 27.000 125.800 27.400 126.600 ;
        RECT 27.700 126.200 28.000 126.800 ;
        RECT 27.700 125.800 28.200 126.200 ;
        RECT 30.400 126.100 30.700 126.800 ;
        RECT 34.500 126.700 34.900 126.800 ;
        RECT 28.600 125.800 30.700 126.100 ;
        RECT 31.000 125.800 31.400 126.600 ;
        RECT 33.700 126.200 34.100 126.300 ;
        RECT 33.700 125.900 36.200 126.200 ;
        RECT 35.800 125.800 36.200 125.900 ;
        RECT 27.700 125.100 28.000 125.800 ;
        RECT 28.600 125.200 28.900 125.800 ;
        RECT 28.600 125.100 29.000 125.200 ;
        RECT 27.500 124.800 28.000 125.100 ;
        RECT 28.300 124.800 29.000 125.100 ;
        RECT 29.400 125.100 29.800 125.200 ;
        RECT 30.400 125.100 30.700 125.800 ;
        RECT 32.600 125.500 35.400 125.600 ;
        RECT 32.600 125.400 35.500 125.500 ;
        RECT 32.600 125.300 37.500 125.400 ;
        RECT 29.400 124.800 30.100 125.100 ;
        RECT 30.400 124.800 30.900 125.100 ;
        RECT 27.500 121.100 27.900 124.800 ;
        RECT 28.300 124.200 28.600 124.800 ;
        RECT 28.200 123.800 28.600 124.200 ;
        RECT 29.800 124.200 30.100 124.800 ;
        RECT 29.800 123.800 30.200 124.200 ;
        RECT 30.500 121.100 30.900 124.800 ;
        RECT 32.600 121.100 33.000 125.300 ;
        RECT 35.100 125.100 37.500 125.300 ;
        RECT 34.200 124.500 36.900 124.800 ;
        RECT 34.200 124.400 34.600 124.500 ;
        RECT 36.500 124.400 36.900 124.500 ;
        RECT 37.200 124.500 37.500 125.100 ;
        RECT 38.200 125.200 38.500 126.800 ;
        RECT 39.000 126.400 39.400 126.500 ;
        RECT 39.000 126.100 40.900 126.400 ;
        RECT 40.500 126.000 40.900 126.100 ;
        RECT 39.700 125.700 40.100 125.800 ;
        RECT 41.400 125.700 41.800 127.400 ;
        RECT 39.700 125.400 41.800 125.700 ;
        RECT 38.200 124.900 39.400 125.200 ;
        RECT 37.900 124.500 38.300 124.600 ;
        RECT 37.200 124.200 38.300 124.500 ;
        RECT 39.100 124.400 39.400 124.900 ;
        RECT 39.100 124.000 39.800 124.400 ;
        RECT 35.900 123.700 36.300 123.800 ;
        RECT 37.300 123.700 37.700 123.800 ;
        RECT 34.200 123.100 34.600 123.500 ;
        RECT 35.900 123.400 37.700 123.700 ;
        RECT 37.000 123.100 37.300 123.400 ;
        RECT 39.000 123.100 39.400 123.500 ;
        RECT 34.200 122.800 35.200 123.100 ;
        RECT 34.800 121.100 35.200 122.800 ;
        RECT 37.000 121.100 37.400 123.100 ;
        RECT 39.100 121.100 39.700 123.100 ;
        RECT 41.400 121.100 41.800 125.400 ;
        RECT 43.800 121.100 44.200 129.900 ;
        RECT 44.600 127.800 45.000 128.600 ;
        RECT 45.400 127.900 45.800 129.900 ;
        RECT 46.200 128.000 46.600 129.900 ;
        RECT 47.800 128.000 48.200 129.900 ;
        RECT 46.200 127.900 48.200 128.000 ;
        RECT 45.500 127.200 45.800 127.900 ;
        RECT 46.300 127.700 48.100 127.900 ;
        RECT 47.400 127.200 47.800 127.400 ;
        RECT 45.400 126.800 46.700 127.200 ;
        RECT 47.400 126.900 48.200 127.200 ;
        RECT 47.800 126.800 48.200 126.900 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 46.400 126.100 46.700 126.800 ;
        RECT 45.400 125.800 46.700 126.100 ;
        RECT 47.000 125.800 47.400 126.600 ;
        RECT 45.400 125.100 45.800 125.200 ;
        RECT 46.400 125.100 46.700 125.800 ;
        RECT 45.400 124.800 46.100 125.100 ;
        RECT 46.400 124.800 46.900 125.100 ;
        RECT 45.800 124.200 46.100 124.800 ;
        RECT 45.800 123.800 46.200 124.200 ;
        RECT 46.500 121.100 46.900 124.800 ;
        RECT 49.400 121.100 49.800 129.900 ;
        RECT 51.000 128.000 51.400 129.900 ;
        RECT 52.600 128.000 53.000 129.900 ;
        RECT 51.000 127.900 53.000 128.000 ;
        RECT 53.400 127.900 53.800 129.900 ;
        RECT 54.500 128.200 54.900 129.900 ;
        RECT 54.500 127.900 55.400 128.200 ;
        RECT 51.100 127.700 52.900 127.900 ;
        RECT 50.200 126.800 50.600 127.600 ;
        RECT 51.400 127.200 51.800 127.400 ;
        RECT 53.400 127.200 53.700 127.900 ;
        RECT 51.000 126.900 51.800 127.200 ;
        RECT 51.000 126.800 51.400 126.900 ;
        RECT 52.500 126.800 53.800 127.200 ;
        RECT 51.800 125.800 52.200 126.600 ;
        RECT 52.500 125.100 52.800 126.800 ;
        RECT 55.000 126.100 55.400 127.900 ;
        RECT 56.600 127.800 57.000 128.600 ;
        RECT 55.800 127.100 56.200 127.600 ;
        RECT 56.600 127.100 56.900 127.800 ;
        RECT 55.800 126.800 56.900 127.100 ;
        RECT 57.400 127.100 57.800 129.900 ;
        RECT 58.200 128.000 58.600 129.900 ;
        RECT 59.800 128.000 60.200 129.900 ;
        RECT 58.200 127.900 60.200 128.000 ;
        RECT 60.600 127.900 61.000 129.900 ;
        RECT 61.700 128.200 62.100 129.900 ;
        RECT 61.700 127.900 62.600 128.200 ;
        RECT 58.300 127.700 60.100 127.900 ;
        RECT 58.600 127.200 59.000 127.400 ;
        RECT 60.600 127.200 60.900 127.900 ;
        RECT 58.200 127.100 59.000 127.200 ;
        RECT 57.400 126.900 59.000 127.100 ;
        RECT 57.400 126.800 58.600 126.900 ;
        RECT 59.700 126.800 61.000 127.200 ;
        RECT 53.400 125.800 55.400 126.100 ;
        RECT 53.400 125.200 53.700 125.800 ;
        RECT 53.400 125.100 53.800 125.200 ;
        RECT 52.300 124.800 52.800 125.100 ;
        RECT 53.100 124.800 53.800 125.100 ;
        RECT 52.300 121.100 52.700 124.800 ;
        RECT 53.100 124.200 53.400 124.800 ;
        RECT 54.200 124.400 54.600 125.200 ;
        RECT 53.000 123.800 53.400 124.200 ;
        RECT 55.000 121.100 55.400 125.800 ;
        RECT 57.400 121.100 57.800 126.800 ;
        RECT 59.000 125.800 59.400 126.600 ;
        RECT 59.700 125.100 60.000 126.800 ;
        RECT 62.200 126.100 62.600 127.900 ;
        RECT 63.800 127.800 64.200 128.600 ;
        RECT 63.000 126.800 63.400 127.600 ;
        RECT 60.600 125.800 62.600 126.100 ;
        RECT 60.600 125.200 60.900 125.800 ;
        RECT 60.600 125.100 61.000 125.200 ;
        RECT 59.500 124.800 60.000 125.100 ;
        RECT 60.300 124.800 61.000 125.100 ;
        RECT 59.500 122.200 59.900 124.800 ;
        RECT 60.300 124.200 60.600 124.800 ;
        RECT 60.200 123.800 60.600 124.200 ;
        RECT 61.400 123.800 61.800 125.200 ;
        RECT 59.000 121.800 59.900 122.200 ;
        RECT 59.500 121.100 59.900 121.800 ;
        RECT 62.200 121.100 62.600 125.800 ;
        RECT 64.600 121.100 65.000 129.900 ;
        RECT 65.400 127.500 65.800 129.900 ;
        RECT 67.600 129.200 68.000 129.900 ;
        RECT 67.000 128.900 68.000 129.200 ;
        RECT 69.800 128.900 70.200 129.900 ;
        RECT 71.900 129.200 72.500 129.900 ;
        RECT 71.800 128.900 72.500 129.200 ;
        RECT 67.000 128.500 67.400 128.900 ;
        RECT 69.800 128.600 70.100 128.900 ;
        RECT 67.800 128.200 68.200 128.600 ;
        RECT 68.700 128.300 70.100 128.600 ;
        RECT 71.800 128.500 72.200 128.900 ;
        RECT 68.700 128.200 69.100 128.300 ;
        RECT 65.800 127.100 66.600 127.200 ;
        RECT 67.900 127.100 68.200 128.200 ;
        RECT 72.700 127.700 73.100 127.800 ;
        RECT 74.200 127.700 74.600 129.900 ;
        RECT 75.000 127.800 75.400 128.600 ;
        RECT 72.700 127.400 74.600 127.700 ;
        RECT 70.700 127.100 71.100 127.200 ;
        RECT 65.800 126.800 71.300 127.100 ;
        RECT 67.300 126.700 67.700 126.800 ;
        RECT 66.500 126.200 66.900 126.300 ;
        RECT 66.500 126.100 69.000 126.200 ;
        RECT 69.400 126.100 69.800 126.200 ;
        RECT 66.500 125.900 69.800 126.100 ;
        RECT 68.600 125.800 69.800 125.900 ;
        RECT 70.200 126.100 70.600 126.200 ;
        RECT 71.000 126.100 71.300 126.800 ;
        RECT 71.800 126.400 72.200 126.500 ;
        RECT 71.800 126.100 73.700 126.400 ;
        RECT 70.200 125.800 71.300 126.100 ;
        RECT 73.300 126.000 73.700 126.100 ;
        RECT 65.400 125.500 68.200 125.600 ;
        RECT 65.400 125.400 68.300 125.500 ;
        RECT 65.400 125.300 70.300 125.400 ;
        RECT 65.400 121.100 65.800 125.300 ;
        RECT 67.900 125.100 70.300 125.300 ;
        RECT 67.000 124.500 69.700 124.800 ;
        RECT 67.000 124.400 67.400 124.500 ;
        RECT 69.300 124.400 69.700 124.500 ;
        RECT 70.000 124.500 70.300 125.100 ;
        RECT 71.000 125.200 71.300 125.800 ;
        RECT 72.500 125.700 72.900 125.800 ;
        RECT 74.200 125.700 74.600 127.400 ;
        RECT 72.500 125.400 74.600 125.700 ;
        RECT 71.000 124.900 72.200 125.200 ;
        RECT 70.700 124.500 71.100 124.600 ;
        RECT 70.000 124.200 71.100 124.500 ;
        RECT 71.900 124.400 72.200 124.900 ;
        RECT 71.900 124.000 72.600 124.400 ;
        RECT 68.700 123.700 69.100 123.800 ;
        RECT 70.100 123.700 70.500 123.800 ;
        RECT 67.000 123.100 67.400 123.500 ;
        RECT 68.700 123.400 70.500 123.700 ;
        RECT 69.800 123.100 70.100 123.400 ;
        RECT 71.800 123.100 72.200 123.500 ;
        RECT 67.000 122.800 68.000 123.100 ;
        RECT 67.600 121.100 68.000 122.800 ;
        RECT 69.800 121.100 70.200 123.100 ;
        RECT 71.900 121.100 72.500 123.100 ;
        RECT 74.200 121.100 74.600 125.400 ;
        RECT 75.000 124.100 75.400 124.200 ;
        RECT 75.800 124.100 76.200 129.900 ;
        RECT 76.600 127.800 77.000 128.600 ;
        RECT 75.000 123.800 76.200 124.100 ;
        RECT 75.800 121.100 76.200 123.800 ;
        RECT 77.400 121.100 77.800 129.900 ;
        RECT 78.200 128.000 78.600 129.900 ;
        RECT 79.800 128.000 80.200 129.900 ;
        RECT 78.200 127.900 80.200 128.000 ;
        RECT 80.600 127.900 81.000 129.900 ;
        RECT 81.700 128.200 82.100 129.900 ;
        RECT 81.700 127.900 82.600 128.200 ;
        RECT 78.300 127.700 80.100 127.900 ;
        RECT 78.600 127.200 79.000 127.400 ;
        RECT 80.600 127.200 80.900 127.900 ;
        RECT 78.200 126.900 79.000 127.200 ;
        RECT 78.200 126.800 78.600 126.900 ;
        RECT 79.700 126.800 81.000 127.200 ;
        RECT 79.000 125.800 79.400 126.600 ;
        RECT 79.700 125.100 80.000 126.800 ;
        RECT 82.200 126.100 82.600 127.900 ;
        RECT 83.000 126.800 83.400 127.600 ;
        RECT 83.800 127.500 84.200 129.900 ;
        RECT 86.000 129.200 86.400 129.900 ;
        RECT 85.400 128.900 86.400 129.200 ;
        RECT 88.200 128.900 88.600 129.900 ;
        RECT 90.300 129.200 90.900 129.900 ;
        RECT 90.200 128.900 90.900 129.200 ;
        RECT 85.400 128.500 85.800 128.900 ;
        RECT 88.200 128.600 88.500 128.900 ;
        RECT 86.200 128.200 86.600 128.600 ;
        RECT 87.100 128.300 88.500 128.600 ;
        RECT 90.200 128.500 90.600 128.900 ;
        RECT 87.100 128.200 87.500 128.300 ;
        RECT 84.200 127.100 85.000 127.200 ;
        RECT 86.300 127.100 86.600 128.200 ;
        RECT 91.100 127.700 91.500 127.800 ;
        RECT 92.600 127.700 93.000 129.900 ;
        RECT 94.200 129.100 94.600 129.200 ;
        RECT 95.300 129.100 95.700 129.900 ;
        RECT 94.200 128.800 95.700 129.100 ;
        RECT 95.300 128.200 95.700 128.800 ;
        RECT 98.200 128.900 98.600 129.900 ;
        RECT 95.300 127.900 96.200 128.200 ;
        RECT 91.100 127.400 93.000 127.700 ;
        RECT 87.000 127.100 87.400 127.200 ;
        RECT 89.100 127.100 89.500 127.200 ;
        RECT 84.200 126.800 89.700 127.100 ;
        RECT 85.700 126.700 86.100 126.800 ;
        RECT 80.600 125.800 82.600 126.100 ;
        RECT 84.900 126.200 85.300 126.300 ;
        RECT 86.200 126.200 86.600 126.300 ;
        RECT 84.900 125.900 87.400 126.200 ;
        RECT 87.000 125.800 87.400 125.900 ;
        RECT 80.600 125.200 80.900 125.800 ;
        RECT 80.600 125.100 81.000 125.200 ;
        RECT 79.500 124.800 80.000 125.100 ;
        RECT 80.300 124.800 81.000 125.100 ;
        RECT 79.500 121.100 79.900 124.800 ;
        RECT 80.300 124.200 80.600 124.800 ;
        RECT 81.400 124.400 81.800 125.200 ;
        RECT 80.200 123.800 80.600 124.200 ;
        RECT 82.200 121.100 82.600 125.800 ;
        RECT 83.800 125.500 86.600 125.600 ;
        RECT 83.800 125.400 86.700 125.500 ;
        RECT 83.800 125.300 88.700 125.400 ;
        RECT 83.800 121.100 84.200 125.300 ;
        RECT 86.300 125.100 88.700 125.300 ;
        RECT 85.400 124.500 88.100 124.800 ;
        RECT 85.400 124.400 85.800 124.500 ;
        RECT 87.700 124.400 88.100 124.500 ;
        RECT 88.400 124.500 88.700 125.100 ;
        RECT 89.400 125.200 89.700 126.800 ;
        RECT 90.200 126.400 90.600 126.500 ;
        RECT 90.200 126.100 92.100 126.400 ;
        RECT 91.700 126.000 92.100 126.100 ;
        RECT 90.900 125.700 91.300 125.800 ;
        RECT 92.600 125.700 93.000 127.400 ;
        RECT 90.900 125.400 93.000 125.700 ;
        RECT 89.400 124.900 90.600 125.200 ;
        RECT 89.100 124.500 89.500 124.600 ;
        RECT 88.400 124.200 89.500 124.500 ;
        RECT 90.300 124.400 90.600 124.900 ;
        RECT 90.300 124.000 91.000 124.400 ;
        RECT 87.100 123.700 87.500 123.800 ;
        RECT 88.500 123.700 88.900 123.800 ;
        RECT 85.400 123.100 85.800 123.500 ;
        RECT 87.100 123.400 88.900 123.700 ;
        RECT 88.200 123.100 88.500 123.400 ;
        RECT 90.200 123.100 90.600 123.500 ;
        RECT 85.400 122.800 86.400 123.100 ;
        RECT 86.000 121.100 86.400 122.800 ;
        RECT 88.200 121.100 88.600 123.100 ;
        RECT 90.300 121.100 90.900 123.100 ;
        RECT 92.600 121.100 93.000 125.400 ;
        RECT 95.000 124.400 95.400 125.200 ;
        RECT 95.800 121.100 96.200 127.900 ;
        RECT 96.600 126.800 97.000 127.600 ;
        RECT 98.200 127.200 98.500 128.900 ;
        RECT 99.000 127.800 99.400 128.600 ;
        RECT 98.200 126.800 98.600 127.200 ;
        RECT 100.400 127.100 100.800 129.900 ;
        RECT 103.600 127.100 104.000 129.900 ;
        RECT 106.200 128.000 106.600 129.900 ;
        RECT 107.800 129.600 109.800 129.900 ;
        RECT 107.800 128.000 108.200 129.600 ;
        RECT 106.200 127.900 108.200 128.000 ;
        RECT 106.300 127.700 108.100 127.900 ;
        RECT 108.600 127.800 109.000 129.300 ;
        RECT 109.400 127.900 109.800 129.600 ;
        RECT 106.600 127.200 107.000 127.400 ;
        RECT 108.700 127.200 109.000 127.800 ;
        RECT 99.900 126.900 100.800 127.100 ;
        RECT 103.100 126.900 104.000 127.100 ;
        RECT 106.200 126.900 107.000 127.200 ;
        RECT 107.800 126.900 109.000 127.200 ;
        RECT 99.900 126.800 100.700 126.900 ;
        RECT 103.100 126.800 103.900 126.900 ;
        RECT 106.200 126.800 106.600 126.900 ;
        RECT 107.800 126.800 108.200 126.900 ;
        RECT 97.400 125.400 97.800 126.200 ;
        RECT 98.200 125.100 98.500 126.800 ;
        RECT 99.900 125.200 100.200 126.800 ;
        RECT 101.000 125.800 101.800 126.200 ;
        RECT 97.700 124.700 98.600 125.100 ;
        RECT 99.800 124.800 100.200 125.200 ;
        RECT 102.200 124.800 102.600 125.600 ;
        RECT 103.100 125.200 103.400 126.800 ;
        RECT 103.800 125.800 105.000 126.200 ;
        RECT 107.000 125.800 107.400 126.600 ;
        RECT 103.000 124.800 103.400 125.200 ;
        RECT 105.400 124.800 105.800 125.600 ;
        RECT 107.800 125.100 108.100 126.800 ;
        RECT 108.600 125.800 109.000 126.600 ;
        RECT 109.400 126.400 109.800 127.200 ;
        RECT 110.800 127.100 111.200 129.900 ;
        RECT 114.000 129.100 114.400 129.900 ;
        RECT 115.000 129.100 115.400 129.200 ;
        RECT 114.000 128.800 115.400 129.100 ;
        RECT 117.400 128.900 117.800 129.900 ;
        RECT 114.000 127.100 114.400 128.800 ;
        RECT 110.300 126.900 111.200 127.100 ;
        RECT 113.500 126.900 114.400 127.100 ;
        RECT 116.600 127.800 117.000 128.600 ;
        RECT 116.600 127.200 116.900 127.800 ;
        RECT 117.500 127.200 117.800 128.900 ;
        RECT 110.300 126.800 111.100 126.900 ;
        RECT 113.500 126.800 114.300 126.900 ;
        RECT 116.600 126.800 117.000 127.200 ;
        RECT 117.400 127.100 117.800 127.200 ;
        RECT 118.200 127.100 118.600 127.200 ;
        RECT 117.400 126.800 118.600 127.100 ;
        RECT 120.800 127.100 121.200 129.900 ;
        RECT 123.000 128.200 123.400 129.900 ;
        RECT 122.900 127.900 123.400 128.200 ;
        RECT 122.900 127.200 123.200 127.900 ;
        RECT 124.600 127.600 125.000 129.900 ;
        RECT 123.700 127.300 125.000 127.600 ;
        RECT 125.400 127.500 125.800 129.900 ;
        RECT 127.600 129.200 128.000 129.900 ;
        RECT 127.000 128.900 128.000 129.200 ;
        RECT 129.800 128.900 130.200 129.900 ;
        RECT 131.900 129.200 132.500 129.900 ;
        RECT 131.800 128.900 132.500 129.200 ;
        RECT 127.000 128.500 127.400 128.900 ;
        RECT 129.800 128.600 130.100 128.900 ;
        RECT 127.800 128.200 128.200 128.600 ;
        RECT 128.700 128.300 130.100 128.600 ;
        RECT 131.800 128.500 132.200 128.900 ;
        RECT 128.700 128.200 129.100 128.300 ;
        RECT 120.800 126.900 121.700 127.100 ;
        RECT 120.900 126.800 121.700 126.900 ;
        RECT 110.300 125.200 110.600 126.800 ;
        RECT 111.400 125.800 112.200 126.200 ;
        RECT 97.700 121.100 98.100 124.700 ;
        RECT 99.900 123.500 100.200 124.800 ;
        RECT 100.600 123.800 101.000 124.600 ;
        RECT 103.100 123.500 103.400 124.800 ;
        RECT 103.800 123.800 104.200 124.600 ;
        RECT 99.900 123.200 101.700 123.500 ;
        RECT 99.900 123.100 100.200 123.200 ;
        RECT 99.800 121.100 100.200 123.100 ;
        RECT 101.400 123.100 101.700 123.200 ;
        RECT 103.100 123.200 104.900 123.500 ;
        RECT 103.100 123.100 103.400 123.200 ;
        RECT 101.400 121.100 101.800 123.100 ;
        RECT 103.000 121.100 103.400 123.100 ;
        RECT 104.600 123.100 104.900 123.200 ;
        RECT 104.600 121.100 105.000 123.100 ;
        RECT 107.500 121.100 108.500 125.100 ;
        RECT 110.200 124.800 110.600 125.200 ;
        RECT 112.600 124.800 113.000 125.600 ;
        RECT 113.500 125.200 113.800 126.800 ;
        RECT 114.600 125.800 115.400 126.200 ;
        RECT 113.400 124.800 113.800 125.200 ;
        RECT 110.300 123.500 110.600 124.800 ;
        RECT 111.000 123.800 111.400 124.600 ;
        RECT 113.500 123.500 113.800 124.800 ;
        RECT 114.200 124.800 115.300 125.100 ;
        RECT 115.800 124.800 116.200 125.600 ;
        RECT 117.500 125.100 117.800 126.800 ;
        RECT 118.200 125.400 118.600 126.200 ;
        RECT 119.800 125.800 120.600 126.200 ;
        RECT 114.200 123.800 114.600 124.800 ;
        RECT 115.000 124.200 115.300 124.800 ;
        RECT 117.400 124.700 118.300 125.100 ;
        RECT 119.000 124.800 119.400 125.600 ;
        RECT 121.400 125.200 121.700 126.800 ;
        RECT 122.900 126.800 123.400 127.200 ;
        RECT 121.400 124.800 121.800 125.200 ;
        RECT 122.900 125.100 123.200 126.800 ;
        RECT 123.700 126.500 124.000 127.300 ;
        RECT 125.800 127.100 126.600 127.200 ;
        RECT 127.900 127.100 128.200 128.200 ;
        RECT 132.700 127.700 133.100 127.800 ;
        RECT 134.200 127.700 134.600 129.900 ;
        RECT 135.000 127.900 135.400 129.900 ;
        RECT 135.800 128.000 136.200 129.900 ;
        RECT 137.400 128.000 137.800 129.900 ;
        RECT 139.500 128.200 139.900 129.900 ;
        RECT 141.400 129.100 141.800 129.200 ;
        RECT 142.200 129.100 142.600 129.900 ;
        RECT 141.400 128.800 142.600 129.100 ;
        RECT 135.800 127.900 137.800 128.000 ;
        RECT 139.000 127.900 139.900 128.200 ;
        RECT 142.200 127.900 142.600 128.800 ;
        RECT 143.000 128.000 143.400 129.900 ;
        RECT 144.600 128.000 145.000 129.900 ;
        RECT 146.700 128.200 147.100 129.900 ;
        RECT 143.000 127.900 145.000 128.000 ;
        RECT 146.200 127.900 147.100 128.200 ;
        RECT 147.800 127.900 148.200 129.900 ;
        RECT 148.600 128.000 149.000 129.900 ;
        RECT 150.200 128.000 150.600 129.900 ;
        RECT 148.600 127.900 150.600 128.000 ;
        RECT 132.700 127.400 134.600 127.700 ;
        RECT 128.600 127.100 129.000 127.200 ;
        RECT 130.700 127.100 131.100 127.200 ;
        RECT 125.800 126.800 131.300 127.100 ;
        RECT 127.300 126.700 127.700 126.800 ;
        RECT 123.500 126.100 124.000 126.500 ;
        RECT 123.700 125.100 124.000 126.100 ;
        RECT 124.500 126.200 124.900 126.600 ;
        RECT 126.500 126.200 126.900 126.300 ;
        RECT 124.500 125.800 125.000 126.200 ;
        RECT 126.500 126.100 129.000 126.200 ;
        RECT 129.400 126.100 129.800 126.200 ;
        RECT 126.500 125.900 129.800 126.100 ;
        RECT 128.600 125.800 129.800 125.900 ;
        RECT 125.400 125.500 128.200 125.600 ;
        RECT 125.400 125.400 128.300 125.500 ;
        RECT 125.400 125.300 130.300 125.400 ;
        RECT 115.000 123.800 115.400 124.200 ;
        RECT 110.300 123.200 112.100 123.500 ;
        RECT 110.300 123.100 110.600 123.200 ;
        RECT 110.200 121.100 110.600 123.100 ;
        RECT 111.800 123.100 112.100 123.200 ;
        RECT 113.500 123.200 115.300 123.500 ;
        RECT 113.500 123.100 113.800 123.200 ;
        RECT 111.800 121.100 112.200 123.100 ;
        RECT 113.400 121.100 113.800 123.100 ;
        RECT 115.000 123.100 115.300 123.200 ;
        RECT 115.000 121.100 115.400 123.100 ;
        RECT 117.900 121.100 118.300 124.700 ;
        RECT 120.600 123.800 121.000 124.600 ;
        RECT 121.400 123.500 121.700 124.800 ;
        RECT 122.900 124.600 123.400 125.100 ;
        RECT 123.700 124.800 125.000 125.100 ;
        RECT 119.900 123.200 121.700 123.500 ;
        RECT 119.900 123.100 120.200 123.200 ;
        RECT 119.800 121.100 120.200 123.100 ;
        RECT 121.400 123.100 121.700 123.200 ;
        RECT 121.400 121.100 121.800 123.100 ;
        RECT 123.000 121.100 123.400 124.600 ;
        RECT 124.600 121.100 125.000 124.800 ;
        RECT 125.400 121.100 125.800 125.300 ;
        RECT 127.900 125.100 130.300 125.300 ;
        RECT 127.000 124.500 129.700 124.800 ;
        RECT 127.000 124.400 127.400 124.500 ;
        RECT 129.300 124.400 129.700 124.500 ;
        RECT 130.000 124.500 130.300 125.100 ;
        RECT 131.000 125.200 131.300 126.800 ;
        RECT 131.800 126.400 132.200 126.500 ;
        RECT 131.800 126.100 133.700 126.400 ;
        RECT 133.300 126.000 133.700 126.100 ;
        RECT 132.500 125.700 132.900 125.800 ;
        RECT 134.200 125.700 134.600 127.400 ;
        RECT 135.100 127.200 135.400 127.900 ;
        RECT 135.900 127.700 137.700 127.900 ;
        RECT 137.000 127.200 137.400 127.400 ;
        RECT 135.000 126.800 136.300 127.200 ;
        RECT 137.000 126.900 137.800 127.200 ;
        RECT 137.400 126.800 137.800 126.900 ;
        RECT 138.200 126.800 138.600 127.600 ;
        RECT 136.000 126.200 136.300 126.800 ;
        RECT 135.800 125.800 136.300 126.200 ;
        RECT 136.600 125.800 137.000 126.600 ;
        RECT 139.000 126.100 139.400 127.900 ;
        RECT 142.300 127.200 142.600 127.900 ;
        RECT 143.100 127.700 144.900 127.900 ;
        RECT 144.200 127.200 144.600 127.400 ;
        RECT 142.200 126.800 143.500 127.200 ;
        RECT 144.200 126.900 145.000 127.200 ;
        RECT 144.600 126.800 145.000 126.900 ;
        RECT 145.400 126.800 145.800 127.600 ;
        RECT 142.200 126.100 142.600 126.200 ;
        RECT 139.000 125.800 142.600 126.100 ;
        RECT 132.500 125.400 134.600 125.700 ;
        RECT 131.000 124.900 132.200 125.200 ;
        RECT 130.700 124.500 131.100 124.600 ;
        RECT 130.000 124.200 131.100 124.500 ;
        RECT 131.900 124.400 132.200 124.900 ;
        RECT 131.900 124.000 132.600 124.400 ;
        RECT 128.700 123.700 129.100 123.800 ;
        RECT 130.100 123.700 130.500 123.800 ;
        RECT 127.000 123.100 127.400 123.500 ;
        RECT 128.700 123.400 130.500 123.700 ;
        RECT 129.800 123.100 130.100 123.400 ;
        RECT 131.800 123.100 132.200 123.500 ;
        RECT 127.000 122.800 128.000 123.100 ;
        RECT 127.600 121.100 128.000 122.800 ;
        RECT 129.800 121.100 130.200 123.100 ;
        RECT 131.900 121.100 132.500 123.100 ;
        RECT 134.200 121.100 134.600 125.400 ;
        RECT 135.000 125.100 135.400 125.200 ;
        RECT 136.000 125.100 136.300 125.800 ;
        RECT 135.000 124.800 135.700 125.100 ;
        RECT 136.000 124.800 136.500 125.100 ;
        RECT 135.400 124.200 135.700 124.800 ;
        RECT 135.400 123.800 135.800 124.200 ;
        RECT 136.100 121.100 136.500 124.800 ;
        RECT 139.000 121.100 139.400 125.800 ;
        RECT 139.800 124.400 140.200 125.200 ;
        RECT 141.400 125.100 141.800 125.200 ;
        RECT 142.200 125.100 142.600 125.200 ;
        RECT 143.200 125.100 143.500 126.800 ;
        RECT 143.800 125.800 144.200 126.600 ;
        RECT 141.400 124.800 142.900 125.100 ;
        RECT 143.200 124.800 143.700 125.100 ;
        RECT 142.600 124.200 142.900 124.800 ;
        RECT 142.600 123.800 143.000 124.200 ;
        RECT 143.300 121.100 143.700 124.800 ;
        RECT 146.200 121.100 146.600 127.900 ;
        RECT 147.900 127.200 148.200 127.900 ;
        RECT 148.700 127.700 150.500 127.900 ;
        RECT 149.800 127.200 150.200 127.400 ;
        RECT 147.800 127.100 149.100 127.200 ;
        RECT 147.000 126.800 149.100 127.100 ;
        RECT 149.800 127.100 150.600 127.200 ;
        RECT 151.000 127.100 151.400 129.900 ;
        RECT 149.800 126.900 151.400 127.100 ;
        RECT 150.200 126.800 151.400 126.900 ;
        RECT 151.800 127.800 152.200 128.600 ;
        RECT 151.800 127.200 152.100 127.800 ;
        RECT 152.600 127.700 153.000 129.900 ;
        RECT 154.700 129.200 155.300 129.900 ;
        RECT 154.700 128.900 155.400 129.200 ;
        RECT 157.000 128.900 157.400 129.900 ;
        RECT 159.200 129.200 159.600 129.900 ;
        RECT 159.200 128.900 160.200 129.200 ;
        RECT 155.000 128.500 155.400 128.900 ;
        RECT 157.100 128.600 157.400 128.900 ;
        RECT 157.100 128.300 158.500 128.600 ;
        RECT 158.100 128.200 158.500 128.300 ;
        RECT 159.000 128.200 159.400 128.600 ;
        RECT 159.800 128.500 160.200 128.900 ;
        RECT 154.100 127.700 154.500 127.800 ;
        RECT 152.600 127.400 154.500 127.700 ;
        RECT 151.800 126.800 152.200 127.200 ;
        RECT 147.000 126.200 147.300 126.800 ;
        RECT 147.000 125.800 147.400 126.200 ;
        RECT 147.000 124.400 147.400 125.200 ;
        RECT 147.800 125.100 148.200 125.200 ;
        RECT 148.800 125.100 149.100 126.800 ;
        RECT 149.400 125.800 149.800 126.600 ;
        RECT 147.800 124.800 148.500 125.100 ;
        RECT 148.800 124.800 149.300 125.100 ;
        RECT 148.200 124.200 148.500 124.800 ;
        RECT 148.200 123.800 148.600 124.200 ;
        RECT 148.900 121.100 149.300 124.800 ;
        RECT 151.000 121.100 151.400 126.800 ;
        RECT 152.600 125.700 153.000 127.400 ;
        RECT 156.100 127.100 156.500 127.200 ;
        RECT 159.000 127.100 159.300 128.200 ;
        RECT 161.400 127.500 161.800 129.900 ;
        RECT 162.200 127.900 162.600 129.900 ;
        RECT 163.000 128.000 163.400 129.900 ;
        RECT 164.600 128.000 165.000 129.900 ;
        RECT 163.000 127.900 165.000 128.000 ;
        RECT 162.300 127.200 162.600 127.900 ;
        RECT 163.100 127.700 164.900 127.900 ;
        RECT 164.200 127.200 164.600 127.400 ;
        RECT 160.600 127.100 161.400 127.200 ;
        RECT 155.900 126.800 161.400 127.100 ;
        RECT 162.200 126.800 163.500 127.200 ;
        RECT 164.200 126.900 165.000 127.200 ;
        RECT 166.000 127.100 166.400 129.900 ;
        RECT 169.900 129.200 170.300 129.900 ;
        RECT 169.400 128.800 170.300 129.200 ;
        RECT 169.900 128.200 170.300 128.800 ;
        RECT 171.800 128.200 172.200 129.900 ;
        RECT 169.400 127.900 170.300 128.200 ;
        RECT 171.700 127.900 172.200 128.200 ;
        RECT 164.600 126.800 165.000 126.900 ;
        RECT 165.500 126.900 166.400 127.100 ;
        RECT 165.500 126.800 166.300 126.900 ;
        RECT 168.600 126.800 169.000 127.600 ;
        RECT 155.000 126.400 155.400 126.500 ;
        RECT 153.500 126.100 155.400 126.400 ;
        RECT 155.900 126.200 156.200 126.800 ;
        RECT 159.500 126.700 159.900 126.800 ;
        RECT 159.000 126.200 159.400 126.300 ;
        RECT 160.300 126.200 160.700 126.300 ;
        RECT 153.500 126.000 153.900 126.100 ;
        RECT 155.800 125.800 156.200 126.200 ;
        RECT 158.200 125.900 160.700 126.200 ;
        RECT 158.200 125.800 158.600 125.900 ;
        RECT 154.300 125.700 154.700 125.800 ;
        RECT 152.600 125.400 154.700 125.700 ;
        RECT 152.600 121.100 153.000 125.400 ;
        RECT 155.900 125.200 156.200 125.800 ;
        RECT 159.000 125.500 161.800 125.600 ;
        RECT 158.900 125.400 161.800 125.500 ;
        RECT 155.000 124.900 156.200 125.200 ;
        RECT 156.900 125.300 161.800 125.400 ;
        RECT 156.900 125.100 159.300 125.300 ;
        RECT 155.000 124.400 155.300 124.900 ;
        RECT 154.600 124.000 155.300 124.400 ;
        RECT 156.100 124.500 156.500 124.600 ;
        RECT 156.900 124.500 157.200 125.100 ;
        RECT 156.100 124.200 157.200 124.500 ;
        RECT 157.500 124.500 160.200 124.800 ;
        RECT 157.500 124.400 157.900 124.500 ;
        RECT 159.800 124.400 160.200 124.500 ;
        RECT 156.700 123.700 157.100 123.800 ;
        RECT 158.100 123.700 158.500 123.800 ;
        RECT 155.000 123.100 155.400 123.500 ;
        RECT 156.700 123.400 158.500 123.700 ;
        RECT 157.100 123.100 157.400 123.400 ;
        RECT 159.800 123.100 160.200 123.500 ;
        RECT 154.700 121.100 155.300 123.100 ;
        RECT 157.000 121.100 157.400 123.100 ;
        RECT 159.200 122.800 160.200 123.100 ;
        RECT 159.200 121.100 159.600 122.800 ;
        RECT 161.400 121.100 161.800 125.300 ;
        RECT 162.200 125.100 162.600 125.200 ;
        RECT 163.200 125.100 163.500 126.800 ;
        RECT 163.800 125.800 164.200 126.600 ;
        RECT 165.500 125.200 165.800 126.800 ;
        RECT 166.600 125.800 167.400 126.200 ;
        RECT 162.200 124.800 162.900 125.100 ;
        RECT 163.200 124.800 163.700 125.100 ;
        RECT 165.400 124.800 165.800 125.200 ;
        RECT 167.800 124.800 168.200 125.600 ;
        RECT 162.600 124.200 162.900 124.800 ;
        RECT 162.600 123.800 163.000 124.200 ;
        RECT 163.300 121.100 163.700 124.800 ;
        RECT 165.500 123.500 165.800 124.800 ;
        RECT 166.200 123.800 166.600 124.600 ;
        RECT 165.500 123.200 167.300 123.500 ;
        RECT 165.500 123.100 165.800 123.200 ;
        RECT 165.400 121.100 165.800 123.100 ;
        RECT 167.000 123.100 167.300 123.200 ;
        RECT 167.000 121.100 167.400 123.100 ;
        RECT 169.400 121.100 169.800 127.900 ;
        RECT 171.700 127.200 172.000 127.900 ;
        RECT 173.400 127.600 173.800 129.900 ;
        RECT 174.200 128.000 174.600 129.900 ;
        RECT 175.800 128.000 176.200 129.900 ;
        RECT 174.200 127.900 176.200 128.000 ;
        RECT 176.600 127.900 177.000 129.900 ;
        RECT 177.700 128.200 178.100 129.900 ;
        RECT 177.700 127.900 178.600 128.200 ;
        RECT 174.300 127.700 176.100 127.900 ;
        RECT 172.500 127.300 173.800 127.600 ;
        RECT 171.700 126.800 172.200 127.200 ;
        RECT 170.200 124.400 170.600 125.200 ;
        RECT 171.700 125.100 172.000 126.800 ;
        RECT 172.500 126.500 172.800 127.300 ;
        RECT 174.600 127.200 175.000 127.400 ;
        RECT 176.600 127.200 176.900 127.900 ;
        RECT 174.200 126.900 175.000 127.200 ;
        RECT 174.200 126.800 174.600 126.900 ;
        RECT 175.700 126.800 177.000 127.200 ;
        RECT 172.300 126.100 172.800 126.500 ;
        RECT 172.500 125.100 172.800 126.100 ;
        RECT 173.300 126.200 173.700 126.600 ;
        RECT 173.300 126.100 173.800 126.200 ;
        RECT 174.200 126.100 174.600 126.200 ;
        RECT 173.300 125.800 174.600 126.100 ;
        RECT 175.000 125.800 175.400 126.600 ;
        RECT 175.700 125.100 176.000 126.800 ;
        RECT 178.200 126.100 178.600 127.900 ;
        RECT 179.800 127.700 180.200 129.900 ;
        RECT 181.900 129.200 182.500 129.900 ;
        RECT 181.900 128.900 182.600 129.200 ;
        RECT 184.200 128.900 184.600 129.900 ;
        RECT 186.400 129.200 186.800 129.900 ;
        RECT 186.400 128.900 187.400 129.200 ;
        RECT 182.200 128.500 182.600 128.900 ;
        RECT 184.300 128.600 184.600 128.900 ;
        RECT 184.300 128.300 185.700 128.600 ;
        RECT 185.300 128.200 185.700 128.300 ;
        RECT 186.200 128.200 186.600 128.600 ;
        RECT 187.000 128.500 187.400 128.900 ;
        RECT 181.300 127.700 181.700 127.800 ;
        RECT 179.000 126.800 179.400 127.600 ;
        RECT 179.800 127.400 181.700 127.700 ;
        RECT 176.600 125.800 178.600 126.100 ;
        RECT 176.600 125.200 176.900 125.800 ;
        RECT 176.600 125.100 177.000 125.200 ;
        RECT 171.700 124.600 172.200 125.100 ;
        RECT 172.500 124.800 173.800 125.100 ;
        RECT 171.800 121.100 172.200 124.600 ;
        RECT 173.400 121.100 173.800 124.800 ;
        RECT 175.500 124.800 176.000 125.100 ;
        RECT 176.300 124.800 177.000 125.100 ;
        RECT 175.500 121.100 175.900 124.800 ;
        RECT 176.300 124.200 176.600 124.800 ;
        RECT 177.400 124.400 177.800 125.200 ;
        RECT 176.200 123.800 176.600 124.200 ;
        RECT 178.200 121.100 178.600 125.800 ;
        RECT 179.800 125.700 180.200 127.400 ;
        RECT 183.300 127.100 183.700 127.200 ;
        RECT 186.200 127.100 186.500 128.200 ;
        RECT 188.600 127.500 189.000 129.900 ;
        RECT 189.400 127.900 189.800 129.900 ;
        RECT 190.200 128.000 190.600 129.900 ;
        RECT 191.800 128.000 192.200 129.900 ;
        RECT 190.200 127.900 192.200 128.000 ;
        RECT 189.500 127.200 189.800 127.900 ;
        RECT 190.300 127.700 192.100 127.900 ;
        RECT 194.200 127.600 194.600 129.900 ;
        RECT 195.800 128.200 196.200 129.900 ;
        RECT 197.400 128.500 197.800 129.500 ;
        RECT 195.800 127.900 196.300 128.200 ;
        RECT 191.400 127.200 191.800 127.400 ;
        RECT 194.200 127.300 195.500 127.600 ;
        RECT 187.800 127.100 188.600 127.200 ;
        RECT 183.100 126.800 188.600 127.100 ;
        RECT 189.400 126.800 190.700 127.200 ;
        RECT 191.400 127.100 192.200 127.200 ;
        RECT 193.400 127.100 193.800 127.200 ;
        RECT 191.400 126.900 193.800 127.100 ;
        RECT 191.800 126.800 193.800 126.900 ;
        RECT 182.200 126.400 182.600 126.500 ;
        RECT 180.700 126.100 182.600 126.400 ;
        RECT 180.700 126.000 181.100 126.100 ;
        RECT 181.500 125.700 181.900 125.800 ;
        RECT 179.800 125.400 181.900 125.700 ;
        RECT 179.800 121.100 180.200 125.400 ;
        RECT 183.100 125.200 183.400 126.800 ;
        RECT 186.700 126.700 187.100 126.800 ;
        RECT 187.500 126.200 187.900 126.300 ;
        RECT 183.800 126.100 184.200 126.200 ;
        RECT 185.400 126.100 187.900 126.200 ;
        RECT 183.800 125.900 187.900 126.100 ;
        RECT 183.800 125.800 185.800 125.900 ;
        RECT 186.200 125.500 189.000 125.600 ;
        RECT 186.100 125.400 189.000 125.500 ;
        RECT 182.200 124.900 183.400 125.200 ;
        RECT 184.100 125.300 189.000 125.400 ;
        RECT 184.100 125.100 186.500 125.300 ;
        RECT 182.200 124.400 182.500 124.900 ;
        RECT 181.800 124.000 182.500 124.400 ;
        RECT 183.300 124.500 183.700 124.600 ;
        RECT 184.100 124.500 184.400 125.100 ;
        RECT 183.300 124.200 184.400 124.500 ;
        RECT 184.700 124.500 187.400 124.800 ;
        RECT 184.700 124.400 185.100 124.500 ;
        RECT 187.000 124.400 187.400 124.500 ;
        RECT 183.900 123.700 184.300 123.800 ;
        RECT 185.300 123.700 185.700 123.800 ;
        RECT 182.200 123.100 182.600 123.500 ;
        RECT 183.900 123.400 185.700 123.700 ;
        RECT 184.300 123.100 184.600 123.400 ;
        RECT 187.000 123.100 187.400 123.500 ;
        RECT 181.900 121.100 182.500 123.100 ;
        RECT 184.200 121.100 184.600 123.100 ;
        RECT 186.400 122.800 187.400 123.100 ;
        RECT 186.400 121.100 186.800 122.800 ;
        RECT 188.600 121.100 189.000 125.300 ;
        RECT 189.400 125.100 189.800 125.200 ;
        RECT 190.400 125.100 190.700 126.800 ;
        RECT 191.000 125.800 191.400 126.600 ;
        RECT 194.300 126.200 194.700 126.600 ;
        RECT 194.200 125.800 194.700 126.200 ;
        RECT 195.200 126.500 195.500 127.300 ;
        RECT 196.000 127.200 196.300 127.900 ;
        RECT 195.800 127.100 196.300 127.200 ;
        RECT 197.400 127.400 197.700 128.500 ;
        RECT 199.500 128.000 199.900 129.500 ;
        RECT 199.500 127.700 200.300 128.000 ;
        RECT 199.900 127.500 200.300 127.700 ;
        RECT 197.400 127.100 199.500 127.400 ;
        RECT 195.800 126.800 196.900 127.100 ;
        RECT 195.200 126.100 195.700 126.500 ;
        RECT 195.200 125.100 195.500 126.100 ;
        RECT 196.000 125.100 196.300 126.800 ;
        RECT 196.600 126.100 196.900 126.800 ;
        RECT 199.000 126.900 199.500 127.100 ;
        RECT 200.000 127.200 200.300 127.500 ;
        RECT 203.800 127.900 204.200 129.900 ;
        RECT 204.500 128.200 204.900 128.600 ;
        RECT 204.600 128.100 205.000 128.200 ;
        RECT 205.400 128.100 205.800 129.900 ;
        RECT 197.400 126.100 197.800 126.600 ;
        RECT 196.600 125.800 197.800 126.100 ;
        RECT 198.200 125.800 198.600 126.600 ;
        RECT 199.000 126.500 199.700 126.900 ;
        RECT 200.000 126.800 201.000 127.200 ;
        RECT 199.000 125.500 199.300 126.500 ;
        RECT 200.000 126.200 200.300 126.800 ;
        RECT 203.000 126.400 203.400 127.200 ;
        RECT 199.800 125.800 200.300 126.200 ;
        RECT 189.400 124.800 190.100 125.100 ;
        RECT 190.400 124.800 190.900 125.100 ;
        RECT 189.800 124.200 190.100 124.800 ;
        RECT 189.800 123.800 190.200 124.200 ;
        RECT 190.500 121.100 190.900 124.800 ;
        RECT 194.200 124.800 195.500 125.100 ;
        RECT 194.200 121.100 194.600 124.800 ;
        RECT 195.800 124.600 196.300 125.100 ;
        RECT 197.400 125.200 199.300 125.500 ;
        RECT 195.800 121.100 196.200 124.600 ;
        RECT 197.400 123.500 197.700 125.200 ;
        RECT 200.000 124.900 200.300 125.800 ;
        RECT 200.600 125.400 201.000 126.200 ;
        RECT 202.200 126.100 202.600 126.200 ;
        RECT 203.800 126.100 204.100 127.900 ;
        RECT 204.600 127.800 205.800 128.100 ;
        RECT 206.200 128.000 206.600 129.900 ;
        RECT 207.800 128.000 208.200 129.900 ;
        RECT 206.200 127.900 208.200 128.000 ;
        RECT 208.600 128.500 209.000 129.500 ;
        RECT 205.500 127.200 205.800 127.800 ;
        RECT 206.300 127.700 208.100 127.900 ;
        RECT 208.600 127.400 208.900 128.500 ;
        RECT 210.700 128.200 211.100 129.500 ;
        RECT 214.700 128.200 215.100 129.900 ;
        RECT 210.200 128.000 211.100 128.200 ;
        RECT 210.200 127.800 211.500 128.000 ;
        RECT 210.700 127.700 211.500 127.800 ;
        RECT 211.100 127.500 211.500 127.700 ;
        RECT 214.200 127.900 215.100 128.200 ;
        RECT 215.800 127.900 216.200 129.900 ;
        RECT 216.600 128.000 217.000 129.900 ;
        RECT 218.200 128.000 218.600 129.900 ;
        RECT 216.600 127.900 218.600 128.000 ;
        RECT 207.400 127.200 207.800 127.400 ;
        RECT 205.400 126.800 206.700 127.200 ;
        RECT 207.400 126.900 208.200 127.200 ;
        RECT 208.600 127.100 210.700 127.400 ;
        RECT 207.800 126.800 208.200 126.900 ;
        RECT 210.200 126.900 210.700 127.100 ;
        RECT 211.200 127.200 211.500 127.500 ;
        RECT 204.600 126.100 205.000 126.200 ;
        RECT 202.200 125.800 203.000 126.100 ;
        RECT 203.800 125.800 205.000 126.100 ;
        RECT 202.600 125.600 203.000 125.800 ;
        RECT 204.600 125.100 204.900 125.800 ;
        RECT 205.400 125.100 205.800 125.200 ;
        RECT 206.400 125.100 206.700 126.800 ;
        RECT 207.000 125.800 207.400 126.600 ;
        RECT 208.600 125.800 209.000 126.600 ;
        RECT 209.400 125.800 209.800 126.600 ;
        RECT 210.200 126.500 210.900 126.900 ;
        RECT 211.200 126.800 212.200 127.200 ;
        RECT 213.400 127.100 213.800 127.600 ;
        RECT 212.600 126.800 213.800 127.100 ;
        RECT 210.200 125.500 210.500 126.500 ;
        RECT 208.600 125.200 210.500 125.500 ;
        RECT 199.500 124.600 200.300 124.900 ;
        RECT 202.200 124.800 204.200 125.100 ;
        RECT 197.400 121.500 197.800 123.500 ;
        RECT 199.500 121.100 199.900 124.600 ;
        RECT 202.200 121.100 202.600 124.800 ;
        RECT 203.800 121.100 204.200 124.800 ;
        RECT 204.600 121.100 205.000 125.100 ;
        RECT 205.400 124.800 206.100 125.100 ;
        RECT 206.400 124.800 206.900 125.100 ;
        RECT 205.800 124.200 206.100 124.800 ;
        RECT 205.800 123.800 206.200 124.200 ;
        RECT 206.500 121.100 206.900 124.800 ;
        RECT 208.600 123.500 208.900 125.200 ;
        RECT 211.200 124.900 211.500 126.800 ;
        RECT 211.800 126.100 212.200 126.200 ;
        RECT 212.600 126.100 212.900 126.800 ;
        RECT 211.800 125.800 212.900 126.100 ;
        RECT 214.200 126.100 214.600 127.900 ;
        RECT 215.900 127.200 216.200 127.900 ;
        RECT 216.700 127.700 218.500 127.900 ;
        RECT 219.000 127.700 219.400 129.900 ;
        RECT 221.100 129.200 221.700 129.900 ;
        RECT 221.100 128.900 221.800 129.200 ;
        RECT 223.400 128.900 223.800 129.900 ;
        RECT 225.600 129.200 226.000 129.900 ;
        RECT 225.600 128.900 226.600 129.200 ;
        RECT 221.400 128.500 221.800 128.900 ;
        RECT 223.500 128.600 223.800 128.900 ;
        RECT 223.500 128.300 224.900 128.600 ;
        RECT 224.500 128.200 224.900 128.300 ;
        RECT 225.400 128.200 225.800 128.600 ;
        RECT 226.200 128.500 226.600 128.900 ;
        RECT 220.500 127.700 220.900 127.800 ;
        RECT 219.000 127.400 220.900 127.700 ;
        RECT 217.800 127.200 218.200 127.400 ;
        RECT 215.800 126.800 217.100 127.200 ;
        RECT 217.800 126.900 218.600 127.200 ;
        RECT 218.200 126.800 218.600 126.900 ;
        RECT 216.800 126.200 217.100 126.800 ;
        RECT 214.200 125.800 216.100 126.100 ;
        RECT 216.600 125.800 217.100 126.200 ;
        RECT 217.400 126.100 217.800 126.600 ;
        RECT 218.200 126.100 218.600 126.200 ;
        RECT 217.400 125.800 218.600 126.100 ;
        RECT 211.800 125.400 212.200 125.800 ;
        RECT 210.700 124.600 211.500 124.900 ;
        RECT 208.600 121.500 209.000 123.500 ;
        RECT 210.700 121.100 211.100 124.600 ;
        RECT 214.200 121.100 214.600 125.800 ;
        RECT 215.800 125.200 216.100 125.800 ;
        RECT 215.000 124.400 215.400 125.200 ;
        RECT 215.800 125.100 216.200 125.200 ;
        RECT 216.800 125.100 217.100 125.800 ;
        RECT 219.000 125.700 219.400 127.400 ;
        RECT 222.500 127.100 222.900 127.200 ;
        RECT 223.800 127.100 224.200 127.200 ;
        RECT 225.400 127.100 225.700 128.200 ;
        RECT 227.800 127.500 228.200 129.900 ;
        RECT 228.600 127.600 229.000 129.900 ;
        RECT 228.600 127.300 229.700 127.600 ;
        RECT 227.000 127.100 227.800 127.200 ;
        RECT 222.300 126.800 227.800 127.100 ;
        RECT 221.400 126.400 221.800 126.500 ;
        RECT 219.900 126.100 221.800 126.400 ;
        RECT 219.900 126.000 220.300 126.100 ;
        RECT 220.700 125.700 221.100 125.800 ;
        RECT 219.000 125.400 221.100 125.700 ;
        RECT 215.800 124.800 216.500 125.100 ;
        RECT 216.800 124.800 217.300 125.100 ;
        RECT 216.200 124.200 216.500 124.800 ;
        RECT 216.200 123.800 216.600 124.200 ;
        RECT 216.900 121.100 217.300 124.800 ;
        RECT 219.000 121.100 219.400 125.400 ;
        RECT 222.300 125.200 222.600 126.800 ;
        RECT 225.900 126.700 226.300 126.800 ;
        RECT 226.700 126.200 227.100 126.300 ;
        RECT 224.600 125.900 227.100 126.200 ;
        RECT 224.600 125.800 225.000 125.900 ;
        RECT 228.600 125.800 229.000 126.600 ;
        RECT 229.400 125.800 229.700 127.300 ;
        RECT 225.400 125.500 228.200 125.600 ;
        RECT 225.300 125.400 228.200 125.500 ;
        RECT 221.400 124.900 222.600 125.200 ;
        RECT 223.300 125.300 228.200 125.400 ;
        RECT 223.300 125.100 225.700 125.300 ;
        RECT 221.400 124.400 221.700 124.900 ;
        RECT 221.000 124.200 221.700 124.400 ;
        RECT 222.500 124.500 222.900 124.600 ;
        RECT 223.300 124.500 223.600 125.100 ;
        RECT 222.500 124.200 223.600 124.500 ;
        RECT 223.900 124.500 226.600 124.800 ;
        RECT 223.900 124.400 224.300 124.500 ;
        RECT 226.200 124.400 226.600 124.500 ;
        RECT 220.600 124.000 221.700 124.200 ;
        RECT 220.600 123.800 221.300 124.000 ;
        RECT 223.100 123.700 223.500 123.800 ;
        RECT 224.500 123.700 224.900 123.800 ;
        RECT 221.400 123.100 221.800 123.500 ;
        RECT 223.100 123.400 224.900 123.700 ;
        RECT 223.500 123.100 223.800 123.400 ;
        RECT 226.200 123.100 226.600 123.500 ;
        RECT 221.100 121.100 221.700 123.100 ;
        RECT 223.400 121.100 223.800 123.100 ;
        RECT 225.600 122.800 226.600 123.100 ;
        RECT 225.600 121.100 226.000 122.800 ;
        RECT 227.800 121.100 228.200 125.300 ;
        RECT 229.400 125.400 230.000 125.800 ;
        RECT 229.400 125.100 229.700 125.400 ;
        RECT 228.600 124.800 229.700 125.100 ;
        RECT 228.600 121.100 229.000 124.800 ;
        RECT 1.400 115.600 1.800 119.900 ;
        RECT 3.000 115.600 3.400 119.900 ;
        RECT 1.400 115.200 3.400 115.600 ;
        RECT 4.600 115.700 5.000 119.900 ;
        RECT 6.800 118.200 7.200 119.900 ;
        RECT 6.200 117.900 7.200 118.200 ;
        RECT 9.000 117.900 9.400 119.900 ;
        RECT 11.100 117.900 11.700 119.900 ;
        RECT 6.200 117.500 6.600 117.900 ;
        RECT 9.000 117.600 9.300 117.900 ;
        RECT 7.900 117.300 9.700 117.600 ;
        RECT 11.000 117.500 11.400 117.900 ;
        RECT 7.900 117.200 8.300 117.300 ;
        RECT 9.300 117.200 9.700 117.300 ;
        RECT 6.200 116.500 6.600 116.600 ;
        RECT 8.500 116.500 8.900 116.600 ;
        RECT 6.200 116.200 8.900 116.500 ;
        RECT 9.200 116.500 10.300 116.800 ;
        RECT 9.200 115.900 9.500 116.500 ;
        RECT 9.900 116.400 10.300 116.500 ;
        RECT 11.100 116.600 11.800 117.000 ;
        RECT 11.100 116.100 11.400 116.600 ;
        RECT 7.100 115.700 9.500 115.900 ;
        RECT 4.600 115.600 9.500 115.700 ;
        RECT 10.200 115.800 11.400 116.100 ;
        RECT 4.600 115.500 7.500 115.600 ;
        RECT 4.600 115.400 7.400 115.500 ;
        RECT 10.200 115.200 10.500 115.800 ;
        RECT 13.400 115.600 13.800 119.900 ;
        RECT 15.500 116.200 15.900 119.900 ;
        RECT 16.200 116.800 16.600 117.200 ;
        RECT 17.400 116.800 18.200 117.200 ;
        RECT 16.300 116.200 16.600 116.800 ;
        RECT 17.800 116.200 18.100 116.800 ;
        RECT 18.500 116.200 18.900 119.900 ;
        RECT 15.500 115.900 16.000 116.200 ;
        RECT 16.300 115.900 17.000 116.200 ;
        RECT 11.700 115.300 13.800 115.600 ;
        RECT 11.700 115.200 12.100 115.300 ;
        RECT 3.000 113.800 3.400 115.200 ;
        RECT 7.800 115.100 8.200 115.200 ;
        RECT 5.700 114.800 8.200 115.100 ;
        RECT 10.200 114.800 10.600 115.200 ;
        RECT 12.500 114.900 12.900 115.000 ;
        RECT 5.700 114.700 6.100 114.800 ;
        RECT 6.500 114.200 6.900 114.300 ;
        RECT 10.200 114.200 10.500 114.800 ;
        RECT 11.000 114.600 12.900 114.900 ;
        RECT 11.000 114.500 11.400 114.600 ;
        RECT 5.000 113.900 10.500 114.200 ;
        RECT 5.000 113.800 5.800 113.900 ;
        RECT 1.400 113.400 3.400 113.800 ;
        RECT 1.400 111.100 1.800 113.400 ;
        RECT 3.000 111.100 3.400 113.400 ;
        RECT 4.600 111.100 5.000 113.500 ;
        RECT 7.100 112.800 7.400 113.900 ;
        RECT 9.900 113.800 10.300 113.900 ;
        RECT 13.400 113.600 13.800 115.300 ;
        RECT 15.700 115.200 16.000 115.900 ;
        RECT 16.600 115.800 17.000 115.900 ;
        RECT 17.400 115.900 18.100 116.200 ;
        RECT 18.400 115.900 18.900 116.200 ;
        RECT 17.400 115.800 17.800 115.900 ;
        RECT 15.000 114.400 15.400 115.200 ;
        RECT 15.700 114.800 16.200 115.200 ;
        RECT 16.600 115.100 16.900 115.800 ;
        RECT 18.400 115.100 18.700 115.900 ;
        RECT 16.600 114.800 18.700 115.100 ;
        RECT 15.700 114.200 16.000 114.800 ;
        RECT 18.400 114.200 18.700 114.800 ;
        RECT 19.000 114.400 19.400 115.200 ;
        RECT 14.200 114.100 14.600 114.200 ;
        RECT 14.200 113.800 15.000 114.100 ;
        RECT 15.700 113.800 17.000 114.200 ;
        RECT 17.400 113.800 18.700 114.200 ;
        RECT 19.800 114.100 20.200 114.200 ;
        RECT 19.400 113.800 20.200 114.100 ;
        RECT 14.600 113.600 15.000 113.800 ;
        RECT 11.900 113.300 13.800 113.600 ;
        RECT 11.900 113.200 12.300 113.300 ;
        RECT 6.200 112.100 6.600 112.500 ;
        RECT 7.000 112.400 7.400 112.800 ;
        RECT 7.900 112.700 8.300 112.800 ;
        RECT 7.900 112.400 9.300 112.700 ;
        RECT 9.000 112.100 9.300 112.400 ;
        RECT 11.000 112.100 11.400 112.500 ;
        RECT 6.200 111.800 7.200 112.100 ;
        RECT 6.800 111.100 7.200 111.800 ;
        RECT 9.000 111.100 9.400 112.100 ;
        RECT 11.000 111.800 11.700 112.100 ;
        RECT 11.100 111.100 11.700 111.800 ;
        RECT 13.400 111.100 13.800 113.300 ;
        RECT 14.300 113.100 16.100 113.300 ;
        RECT 16.600 113.100 16.900 113.800 ;
        RECT 17.500 113.100 17.800 113.800 ;
        RECT 19.400 113.600 19.800 113.800 ;
        RECT 18.300 113.100 20.100 113.300 ;
        RECT 14.200 113.000 16.200 113.100 ;
        RECT 14.200 111.100 14.600 113.000 ;
        RECT 15.800 111.100 16.200 113.000 ;
        RECT 16.600 111.100 17.000 113.100 ;
        RECT 17.400 111.100 17.800 113.100 ;
        RECT 18.200 113.000 20.200 113.100 ;
        RECT 18.200 111.100 18.600 113.000 ;
        RECT 19.800 111.100 20.200 113.000 ;
        RECT 20.600 112.400 21.000 113.200 ;
        RECT 21.400 111.100 21.800 119.900 ;
        RECT 23.500 115.900 24.500 119.900 ;
        RECT 27.500 115.900 28.500 119.900 ;
        RECT 22.200 113.800 22.600 114.600 ;
        RECT 23.000 114.400 23.400 115.200 ;
        RECT 23.900 114.200 24.200 115.900 ;
        RECT 24.600 114.400 25.000 115.200 ;
        RECT 23.800 114.100 24.200 114.200 ;
        RECT 25.400 114.100 25.800 114.200 ;
        RECT 23.000 113.800 24.200 114.100 ;
        RECT 25.000 113.800 25.800 114.100 ;
        RECT 26.200 113.800 26.600 114.600 ;
        RECT 27.000 114.400 27.400 115.200 ;
        RECT 27.900 114.200 28.200 115.900 ;
        RECT 28.600 114.400 29.000 115.200 ;
        RECT 27.800 114.100 28.200 114.200 ;
        RECT 29.400 114.100 29.800 114.200 ;
        RECT 30.200 114.100 30.600 119.900 ;
        RECT 32.600 116.400 33.000 119.900 ;
        RECT 27.000 113.800 28.200 114.100 ;
        RECT 29.000 113.800 30.600 114.100 ;
        RECT 23.000 113.100 23.300 113.800 ;
        RECT 25.000 113.600 25.400 113.800 ;
        RECT 23.900 113.100 25.700 113.300 ;
        RECT 27.000 113.100 27.300 113.800 ;
        RECT 29.000 113.600 29.400 113.800 ;
        RECT 27.900 113.100 29.700 113.300 ;
        RECT 22.200 111.400 22.600 113.100 ;
        RECT 23.000 111.700 23.400 113.100 ;
        RECT 23.800 113.000 25.800 113.100 ;
        RECT 23.800 111.400 24.200 113.000 ;
        RECT 22.200 111.100 24.200 111.400 ;
        RECT 25.400 111.100 25.800 113.000 ;
        RECT 26.200 111.400 26.600 113.100 ;
        RECT 27.000 111.700 27.400 113.100 ;
        RECT 27.800 113.000 29.800 113.100 ;
        RECT 27.800 111.400 28.200 113.000 ;
        RECT 26.200 111.100 28.200 111.400 ;
        RECT 29.400 111.100 29.800 113.000 ;
        RECT 30.200 111.100 30.600 113.800 ;
        RECT 32.500 115.900 33.000 116.400 ;
        RECT 34.200 116.200 34.600 119.900 ;
        RECT 33.300 115.900 34.600 116.200 ;
        RECT 36.300 116.200 36.700 119.900 ;
        RECT 41.100 117.200 41.500 119.900 ;
        RECT 37.000 116.800 37.400 117.200 ;
        RECT 40.600 116.800 41.500 117.200 ;
        RECT 41.800 116.800 42.200 117.200 ;
        RECT 37.100 116.200 37.400 116.800 ;
        RECT 41.100 116.200 41.500 116.800 ;
        RECT 41.900 116.200 42.200 116.800 ;
        RECT 43.000 116.200 43.400 119.900 ;
        RECT 44.600 116.400 45.000 119.900 ;
        RECT 36.300 115.900 36.800 116.200 ;
        RECT 37.100 115.900 37.800 116.200 ;
        RECT 41.100 115.900 41.600 116.200 ;
        RECT 41.900 115.900 42.600 116.200 ;
        RECT 43.000 115.900 44.300 116.200 ;
        RECT 44.600 115.900 45.100 116.400 ;
        RECT 47.500 116.200 47.900 119.900 ;
        RECT 48.200 116.800 48.600 117.200 ;
        RECT 48.300 116.200 48.600 116.800 ;
        RECT 49.800 116.800 50.200 117.200 ;
        RECT 49.800 116.200 50.100 116.800 ;
        RECT 50.500 116.200 50.900 119.900 ;
        RECT 47.500 115.900 48.000 116.200 ;
        RECT 48.300 115.900 49.000 116.200 ;
        RECT 32.500 114.200 32.800 115.900 ;
        RECT 33.300 114.900 33.600 115.900 ;
        RECT 33.100 114.500 33.600 114.900 ;
        RECT 32.500 113.800 33.000 114.200 ;
        RECT 32.500 113.200 32.800 113.800 ;
        RECT 33.300 113.700 33.600 114.500 ;
        RECT 34.100 115.100 34.600 115.200 ;
        RECT 35.000 115.100 35.400 115.200 ;
        RECT 34.100 114.800 35.400 115.100 ;
        RECT 34.100 114.400 34.500 114.800 ;
        RECT 35.800 114.400 36.200 115.200 ;
        RECT 36.500 114.200 36.800 115.900 ;
        RECT 37.400 115.800 37.800 115.900 ;
        RECT 40.600 114.400 41.000 115.200 ;
        RECT 41.300 114.200 41.600 115.900 ;
        RECT 42.200 115.800 42.600 115.900 ;
        RECT 43.000 114.800 43.500 115.200 ;
        RECT 43.100 114.400 43.500 114.800 ;
        RECT 44.000 114.900 44.300 115.900 ;
        RECT 44.000 114.500 44.500 114.900 ;
        RECT 35.000 114.100 35.400 114.200 ;
        RECT 35.000 113.800 35.800 114.100 ;
        RECT 36.500 113.800 37.800 114.200 ;
        RECT 39.800 114.100 40.200 114.200 ;
        RECT 39.800 113.800 40.600 114.100 ;
        RECT 41.300 113.800 42.600 114.200 ;
        RECT 33.300 113.400 34.600 113.700 ;
        RECT 35.400 113.600 35.800 113.800 ;
        RECT 31.000 112.400 31.400 113.200 ;
        RECT 32.500 112.800 33.000 113.200 ;
        RECT 32.600 111.100 33.000 112.800 ;
        RECT 34.200 111.100 34.600 113.400 ;
        RECT 35.100 113.100 36.900 113.300 ;
        RECT 37.400 113.100 37.700 113.800 ;
        RECT 40.200 113.600 40.600 113.800 ;
        RECT 39.900 113.100 41.700 113.300 ;
        RECT 42.200 113.100 42.500 113.800 ;
        RECT 44.000 113.700 44.300 114.500 ;
        RECT 44.800 114.200 45.100 115.900 ;
        RECT 47.000 114.400 47.400 115.200 ;
        RECT 47.700 115.100 48.000 115.900 ;
        RECT 48.600 115.800 49.000 115.900 ;
        RECT 49.400 115.900 50.100 116.200 ;
        RECT 50.400 115.900 50.900 116.200 ;
        RECT 49.400 115.800 49.800 115.900 ;
        RECT 49.400 115.100 49.700 115.800 ;
        RECT 50.400 115.200 50.700 115.900 ;
        RECT 52.600 115.600 53.000 119.900 ;
        RECT 54.700 117.900 55.300 119.900 ;
        RECT 57.000 117.900 57.400 119.900 ;
        RECT 59.200 118.200 59.600 119.900 ;
        RECT 59.200 117.900 60.200 118.200 ;
        RECT 55.000 117.500 55.400 117.900 ;
        RECT 57.100 117.600 57.400 117.900 ;
        RECT 56.700 117.300 58.500 117.600 ;
        RECT 59.800 117.500 60.200 117.900 ;
        RECT 56.700 117.200 57.100 117.300 ;
        RECT 58.100 117.200 58.500 117.300 ;
        RECT 54.600 116.600 55.300 117.000 ;
        RECT 55.000 116.100 55.300 116.600 ;
        RECT 56.100 116.500 57.200 116.800 ;
        RECT 56.100 116.400 56.500 116.500 ;
        RECT 55.000 115.800 56.200 116.100 ;
        RECT 52.600 115.300 54.700 115.600 ;
        RECT 47.700 114.800 49.700 115.100 ;
        RECT 50.200 114.800 50.700 115.200 ;
        RECT 47.700 114.200 48.000 114.800 ;
        RECT 50.400 114.200 50.700 114.800 ;
        RECT 51.000 114.400 51.400 115.200 ;
        RECT 44.600 113.800 45.100 114.200 ;
        RECT 46.200 114.100 46.600 114.200 ;
        RECT 46.200 113.800 47.000 114.100 ;
        RECT 47.700 113.800 49.000 114.200 ;
        RECT 49.400 113.800 50.700 114.200 ;
        RECT 51.800 114.100 52.200 114.200 ;
        RECT 51.400 113.800 52.200 114.100 ;
        RECT 43.000 113.400 44.300 113.700 ;
        RECT 35.000 113.000 37.000 113.100 ;
        RECT 35.000 111.100 35.400 113.000 ;
        RECT 36.600 111.100 37.000 113.000 ;
        RECT 37.400 111.100 37.800 113.100 ;
        RECT 39.800 113.000 41.800 113.100 ;
        RECT 39.800 111.100 40.200 113.000 ;
        RECT 41.400 111.100 41.800 113.000 ;
        RECT 42.200 111.100 42.600 113.100 ;
        RECT 43.000 111.100 43.400 113.400 ;
        RECT 44.800 113.100 45.100 113.800 ;
        RECT 46.600 113.600 47.000 113.800 ;
        RECT 46.300 113.100 48.100 113.300 ;
        RECT 48.600 113.100 48.900 113.800 ;
        RECT 49.500 113.100 49.800 113.800 ;
        RECT 51.400 113.600 51.800 113.800 ;
        RECT 52.600 113.600 53.000 115.300 ;
        RECT 54.300 115.200 54.700 115.300 ;
        RECT 53.500 114.900 53.900 115.000 ;
        RECT 53.500 114.600 55.400 114.900 ;
        RECT 55.000 114.500 55.400 114.600 ;
        RECT 55.900 114.200 56.200 115.800 ;
        RECT 56.900 115.900 57.200 116.500 ;
        RECT 57.500 116.500 57.900 116.600 ;
        RECT 59.800 116.500 60.200 116.600 ;
        RECT 57.500 116.200 60.200 116.500 ;
        RECT 56.900 115.700 59.300 115.900 ;
        RECT 61.400 115.700 61.800 119.900 ;
        RECT 62.500 116.200 62.900 119.900 ;
        RECT 56.900 115.600 61.800 115.700 ;
        RECT 58.900 115.500 61.800 115.600 ;
        RECT 59.000 115.400 61.800 115.500 ;
        RECT 62.200 115.900 62.900 116.200 ;
        RECT 62.200 115.200 62.500 115.900 ;
        RECT 64.600 115.600 65.000 119.900 ;
        RECT 65.400 116.200 65.800 119.900 ;
        RECT 67.000 116.400 67.400 119.900 ;
        RECT 69.900 119.200 70.300 119.900 ;
        RECT 69.400 118.800 70.300 119.200 ;
        RECT 65.400 115.900 66.700 116.200 ;
        RECT 67.000 115.900 67.500 116.400 ;
        RECT 69.900 116.200 70.300 118.800 ;
        RECT 70.600 116.800 71.000 117.200 ;
        RECT 71.800 116.800 72.600 117.200 ;
        RECT 70.700 116.200 71.000 116.800 ;
        RECT 72.200 116.200 72.500 116.800 ;
        RECT 72.900 116.200 73.300 119.900 ;
        RECT 69.900 115.900 70.400 116.200 ;
        RECT 70.700 115.900 71.400 116.200 ;
        RECT 63.000 115.400 65.000 115.600 ;
        RECT 62.900 115.300 65.000 115.400 ;
        RECT 57.400 115.100 57.800 115.200 ;
        RECT 58.200 115.100 58.600 115.200 ;
        RECT 57.400 114.800 60.700 115.100 ;
        RECT 60.300 114.700 60.700 114.800 ;
        RECT 62.200 114.800 62.600 115.200 ;
        RECT 62.900 115.000 63.300 115.300 ;
        RECT 59.500 114.200 59.900 114.300 ;
        RECT 62.200 114.200 62.500 114.800 ;
        RECT 55.900 113.900 61.400 114.200 ;
        RECT 56.100 113.800 56.500 113.900 ;
        RECT 52.600 113.300 54.500 113.600 ;
        RECT 50.300 113.100 52.100 113.300 ;
        RECT 44.600 112.800 45.100 113.100 ;
        RECT 46.200 113.000 48.200 113.100 ;
        RECT 44.600 111.100 45.000 112.800 ;
        RECT 46.200 111.100 46.600 113.000 ;
        RECT 47.800 111.100 48.200 113.000 ;
        RECT 48.600 111.100 49.000 113.100 ;
        RECT 49.400 111.100 49.800 113.100 ;
        RECT 50.200 113.000 52.200 113.100 ;
        RECT 50.200 111.100 50.600 113.000 ;
        RECT 51.800 111.100 52.200 113.000 ;
        RECT 52.600 111.100 53.000 113.300 ;
        RECT 54.100 113.200 54.500 113.300 ;
        RECT 59.000 112.800 59.300 113.900 ;
        RECT 60.600 113.800 61.400 113.900 ;
        RECT 62.200 113.800 62.600 114.200 ;
        RECT 58.100 112.700 58.500 112.800 ;
        RECT 55.000 112.100 55.400 112.500 ;
        RECT 57.100 112.400 58.500 112.700 ;
        RECT 59.000 112.400 59.400 112.800 ;
        RECT 57.100 112.100 57.400 112.400 ;
        RECT 59.800 112.100 60.200 112.500 ;
        RECT 54.700 111.800 55.400 112.100 ;
        RECT 54.700 111.100 55.300 111.800 ;
        RECT 57.000 111.100 57.400 112.100 ;
        RECT 59.200 111.800 60.200 112.100 ;
        RECT 59.200 111.100 59.600 111.800 ;
        RECT 61.400 111.100 61.800 113.500 ;
        RECT 62.200 113.100 62.500 113.800 ;
        RECT 62.900 113.500 63.200 115.000 ;
        RECT 65.400 114.800 65.900 115.200 ;
        RECT 63.600 114.200 64.000 114.600 ;
        RECT 65.500 114.400 65.900 114.800 ;
        RECT 66.400 114.900 66.700 115.900 ;
        RECT 66.400 114.500 66.900 114.900 ;
        RECT 63.700 113.800 64.200 114.200 ;
        RECT 66.400 113.700 66.700 114.500 ;
        RECT 67.200 114.200 67.500 115.900 ;
        RECT 69.400 114.400 69.800 115.200 ;
        RECT 70.100 114.200 70.400 115.900 ;
        RECT 71.000 115.800 71.400 115.900 ;
        RECT 71.800 115.900 72.500 116.200 ;
        RECT 72.800 115.900 73.300 116.200 ;
        RECT 76.300 115.900 77.300 119.900 ;
        RECT 71.800 115.800 72.200 115.900 ;
        RECT 71.000 115.100 71.300 115.800 ;
        RECT 72.800 115.100 73.100 115.900 ;
        RECT 71.000 114.800 73.100 115.100 ;
        RECT 72.800 114.200 73.100 114.800 ;
        RECT 73.400 114.400 73.800 115.200 ;
        RECT 75.800 114.400 76.200 115.200 ;
        RECT 76.600 114.200 76.900 115.900 ;
        RECT 77.400 114.400 77.800 115.200 ;
        RECT 67.000 113.800 67.500 114.200 ;
        RECT 68.600 114.100 69.000 114.200 ;
        RECT 68.600 113.800 69.400 114.100 ;
        RECT 70.100 113.800 71.400 114.200 ;
        RECT 71.800 113.800 73.100 114.200 ;
        RECT 74.200 114.100 74.600 114.200 ;
        RECT 73.800 113.800 74.600 114.100 ;
        RECT 75.000 114.100 75.400 114.200 ;
        RECT 76.600 114.100 77.000 114.200 ;
        RECT 75.000 113.800 75.800 114.100 ;
        RECT 76.600 113.800 77.800 114.100 ;
        RECT 78.200 113.800 78.600 114.600 ;
        RECT 62.900 113.200 64.100 113.500 ;
        RECT 65.400 113.400 66.700 113.700 ;
        RECT 62.200 111.100 62.600 113.100 ;
        RECT 63.800 112.100 64.100 113.200 ;
        RECT 64.600 112.400 65.000 113.200 ;
        RECT 63.800 111.100 64.200 112.100 ;
        RECT 65.400 111.100 65.800 113.400 ;
        RECT 67.200 113.100 67.500 113.800 ;
        RECT 69.000 113.600 69.400 113.800 ;
        RECT 68.700 113.100 70.500 113.300 ;
        RECT 71.000 113.100 71.300 113.800 ;
        RECT 71.900 113.100 72.200 113.800 ;
        RECT 73.800 113.600 74.200 113.800 ;
        RECT 75.400 113.600 75.800 113.800 ;
        RECT 72.700 113.100 74.500 113.300 ;
        RECT 75.100 113.100 76.900 113.300 ;
        RECT 77.500 113.200 77.800 113.800 ;
        RECT 67.000 112.800 67.500 113.100 ;
        RECT 68.600 113.000 70.600 113.100 ;
        RECT 67.000 111.100 67.400 112.800 ;
        RECT 68.600 111.100 69.000 113.000 ;
        RECT 70.200 111.100 70.600 113.000 ;
        RECT 71.000 111.100 71.400 113.100 ;
        RECT 71.800 111.100 72.200 113.100 ;
        RECT 72.600 113.000 74.600 113.100 ;
        RECT 72.600 111.100 73.000 113.000 ;
        RECT 74.200 111.100 74.600 113.000 ;
        RECT 75.000 113.000 77.000 113.100 ;
        RECT 75.000 111.100 75.400 113.000 ;
        RECT 76.600 111.400 77.000 113.000 ;
        RECT 77.400 111.700 77.800 113.200 ;
        RECT 78.200 111.400 78.600 113.100 ;
        RECT 76.600 111.100 78.600 111.400 ;
        RECT 79.000 111.100 79.400 119.900 ;
        RECT 80.600 113.400 81.000 114.200 ;
        RECT 79.800 112.400 80.200 113.200 ;
        RECT 81.400 111.100 81.800 119.900 ;
        RECT 83.000 115.600 83.400 119.900 ;
        RECT 85.100 117.900 85.700 119.900 ;
        RECT 87.400 117.900 87.800 119.900 ;
        RECT 89.600 118.200 90.000 119.900 ;
        RECT 89.600 117.900 90.600 118.200 ;
        RECT 85.400 117.500 85.800 117.900 ;
        RECT 87.500 117.600 87.800 117.900 ;
        RECT 87.100 117.300 88.900 117.600 ;
        RECT 90.200 117.500 90.600 117.900 ;
        RECT 87.100 117.200 87.500 117.300 ;
        RECT 88.500 117.200 88.900 117.300 ;
        RECT 85.000 116.600 85.700 117.000 ;
        RECT 85.400 116.100 85.700 116.600 ;
        RECT 86.500 116.500 87.600 116.800 ;
        RECT 86.500 116.400 86.900 116.500 ;
        RECT 85.400 115.800 86.600 116.100 ;
        RECT 83.000 115.300 85.100 115.600 ;
        RECT 83.000 113.600 83.400 115.300 ;
        RECT 84.700 115.200 85.100 115.300 ;
        RECT 86.300 115.100 86.600 115.800 ;
        RECT 87.300 115.900 87.600 116.500 ;
        RECT 87.900 116.500 88.300 116.600 ;
        RECT 90.200 116.500 90.600 116.600 ;
        RECT 87.900 116.200 90.600 116.500 ;
        RECT 87.300 115.700 89.700 115.900 ;
        RECT 91.800 115.700 92.200 119.900 ;
        RECT 87.300 115.600 92.200 115.700 ;
        RECT 89.300 115.500 92.200 115.600 ;
        RECT 89.400 115.400 92.200 115.500 ;
        RECT 87.000 115.100 87.400 115.200 ;
        RECT 83.900 114.900 84.300 115.000 ;
        RECT 83.900 114.600 85.800 114.900 ;
        RECT 86.200 114.800 87.400 115.100 ;
        RECT 88.600 115.100 89.000 115.200 ;
        RECT 95.000 115.100 95.400 119.900 ;
        RECT 97.000 116.800 97.400 117.200 ;
        RECT 95.800 115.800 96.200 116.600 ;
        RECT 97.000 116.200 97.300 116.800 ;
        RECT 97.700 116.200 98.100 119.900 ;
        RECT 96.600 115.900 97.300 116.200 ;
        RECT 97.600 115.900 98.100 116.200 ;
        RECT 96.600 115.800 97.000 115.900 ;
        RECT 96.600 115.100 96.900 115.800 ;
        RECT 88.600 114.800 91.100 115.100 ;
        RECT 85.400 114.500 85.800 114.600 ;
        RECT 86.300 114.200 86.600 114.800 ;
        RECT 89.400 114.700 89.800 114.800 ;
        RECT 90.700 114.700 91.100 114.800 ;
        RECT 95.000 114.800 96.900 115.100 ;
        RECT 89.900 114.200 90.300 114.300 ;
        RECT 86.300 113.900 91.800 114.200 ;
        RECT 86.500 113.800 86.900 113.900 ;
        RECT 83.000 113.300 84.900 113.600 ;
        RECT 83.000 111.100 83.400 113.300 ;
        RECT 84.500 113.200 84.900 113.300 ;
        RECT 89.400 112.800 89.700 113.900 ;
        RECT 91.000 113.800 91.800 113.900 ;
        RECT 92.600 114.100 93.000 114.200 ;
        RECT 94.200 114.100 94.600 114.200 ;
        RECT 92.600 113.800 94.600 114.100 ;
        RECT 88.500 112.700 88.900 112.800 ;
        RECT 85.400 112.100 85.800 112.500 ;
        RECT 87.500 112.400 88.900 112.700 ;
        RECT 89.400 112.400 89.800 112.800 ;
        RECT 87.500 112.100 87.800 112.400 ;
        RECT 90.200 112.100 90.600 112.500 ;
        RECT 85.100 111.800 85.800 112.100 ;
        RECT 85.100 111.100 85.700 111.800 ;
        RECT 87.400 111.100 87.800 112.100 ;
        RECT 89.600 111.800 90.600 112.100 ;
        RECT 89.600 111.100 90.000 111.800 ;
        RECT 91.800 111.100 92.200 113.500 ;
        RECT 94.200 113.400 94.600 113.800 ;
        RECT 95.000 113.100 95.400 114.800 ;
        RECT 97.600 114.200 97.900 115.900 ;
        RECT 98.200 114.400 98.600 115.200 ;
        RECT 96.600 113.800 97.900 114.200 ;
        RECT 99.000 114.100 99.400 114.200 ;
        RECT 98.600 113.800 99.400 114.100 ;
        RECT 96.700 113.100 97.000 113.800 ;
        RECT 98.600 113.600 99.000 113.800 ;
        RECT 99.800 113.400 100.200 114.200 ;
        RECT 97.500 113.100 99.300 113.300 ;
        RECT 100.600 113.100 101.000 119.900 ;
        RECT 101.400 115.800 101.800 116.600 ;
        RECT 102.200 115.800 102.600 117.200 ;
        RECT 103.000 117.100 103.400 119.900 ;
        RECT 103.000 116.800 104.100 117.100 ;
        RECT 103.000 113.100 103.400 116.800 ;
        RECT 103.800 116.200 104.100 116.800 ;
        RECT 105.900 116.200 106.300 119.900 ;
        RECT 106.600 116.800 107.000 117.200 ;
        RECT 106.700 116.200 107.000 116.800 ;
        RECT 103.800 115.800 104.200 116.200 ;
        RECT 105.900 115.900 106.400 116.200 ;
        RECT 106.700 115.900 107.400 116.200 ;
        RECT 103.800 115.100 104.200 115.200 ;
        RECT 103.800 114.800 104.900 115.100 ;
        RECT 104.600 114.200 104.900 114.800 ;
        RECT 105.400 114.400 105.800 115.200 ;
        RECT 106.100 114.200 106.400 115.900 ;
        RECT 107.000 115.800 107.400 115.900 ;
        RECT 107.800 115.800 108.200 116.600 ;
        RECT 107.000 115.100 107.300 115.800 ;
        RECT 108.600 115.100 109.000 119.900 ;
        RECT 107.000 114.800 109.000 115.100 ;
        RECT 103.800 113.400 104.200 114.200 ;
        RECT 104.600 114.100 105.000 114.200 ;
        RECT 104.600 113.800 105.400 114.100 ;
        RECT 106.100 113.800 107.400 114.200 ;
        RECT 105.000 113.600 105.400 113.800 ;
        RECT 104.700 113.100 106.500 113.300 ;
        RECT 107.000 113.100 107.300 113.800 ;
        RECT 108.600 113.100 109.000 114.800 ;
        RECT 109.400 113.400 109.800 114.200 ;
        RECT 95.000 112.800 95.900 113.100 ;
        RECT 95.500 111.100 95.900 112.800 ;
        RECT 96.600 111.100 97.000 113.100 ;
        RECT 97.400 113.000 99.400 113.100 ;
        RECT 97.400 111.100 97.800 113.000 ;
        RECT 99.000 111.100 99.400 113.000 ;
        RECT 100.600 112.800 101.500 113.100 ;
        RECT 101.100 112.200 101.500 112.800 ;
        RECT 102.500 112.800 103.400 113.100 ;
        RECT 104.600 113.000 106.600 113.100 ;
        RECT 101.100 111.800 101.800 112.200 ;
        RECT 101.100 111.100 101.500 111.800 ;
        RECT 102.500 111.100 102.900 112.800 ;
        RECT 104.600 111.100 105.000 113.000 ;
        RECT 106.200 111.100 106.600 113.000 ;
        RECT 107.000 111.100 107.400 113.100 ;
        RECT 108.100 112.800 109.000 113.100 ;
        RECT 108.100 111.100 108.500 112.800 ;
        RECT 110.200 111.100 110.600 119.900 ;
        RECT 111.800 115.800 112.200 116.600 ;
        RECT 111.000 112.400 111.400 113.200 ;
        RECT 112.600 113.100 113.000 119.900 ;
        RECT 114.500 119.200 114.900 119.900 ;
        RECT 114.200 118.800 114.900 119.200 ;
        RECT 114.500 116.300 114.900 118.800 ;
        RECT 116.600 117.900 117.000 119.900 ;
        RECT 116.700 117.800 117.000 117.900 ;
        RECT 118.200 117.900 118.600 119.900 ;
        RECT 118.200 117.800 118.500 117.900 ;
        RECT 116.700 117.500 118.500 117.800 ;
        RECT 114.500 115.900 115.400 116.300 ;
        RECT 116.700 116.200 117.000 117.500 ;
        RECT 117.400 116.400 117.800 117.200 ;
        RECT 121.100 116.300 121.500 119.900 ;
        RECT 123.000 117.900 123.400 119.900 ;
        RECT 123.100 117.800 123.400 117.900 ;
        RECT 124.600 117.900 125.000 119.900 ;
        RECT 124.600 117.800 124.900 117.900 ;
        RECT 123.100 117.500 124.900 117.800 ;
        RECT 123.800 116.400 124.200 117.200 ;
        RECT 114.200 114.800 114.600 115.600 ;
        RECT 115.000 114.200 115.300 115.900 ;
        RECT 116.600 115.800 117.000 116.200 ;
        RECT 116.700 114.200 117.000 115.800 ;
        RECT 119.000 115.400 119.400 116.200 ;
        RECT 120.600 115.900 121.500 116.300 ;
        RECT 124.600 116.200 124.900 117.500 ;
        RECT 122.200 116.100 122.600 116.200 ;
        RECT 123.000 116.100 123.400 116.200 ;
        RECT 117.800 114.800 118.600 115.200 ;
        RECT 120.700 114.200 121.000 115.900 ;
        RECT 122.200 115.800 123.400 116.100 ;
        RECT 124.600 115.800 125.000 116.200 ;
        RECT 125.400 115.800 125.800 116.600 ;
        RECT 121.400 114.800 121.800 115.600 ;
        RECT 122.200 115.400 122.600 115.800 ;
        RECT 123.000 114.800 123.800 115.200 ;
        RECT 124.600 114.200 124.900 115.800 ;
        RECT 113.400 113.400 113.800 114.200 ;
        RECT 115.000 113.800 115.400 114.200 ;
        RECT 116.700 114.100 117.500 114.200 ;
        RECT 116.700 113.900 117.600 114.100 ;
        RECT 112.100 112.800 113.000 113.100 ;
        RECT 112.100 112.200 112.500 112.800 ;
        RECT 111.800 111.800 112.500 112.200 ;
        RECT 112.100 111.100 112.500 111.800 ;
        RECT 115.000 112.100 115.300 113.800 ;
        RECT 115.800 112.400 116.200 113.200 ;
        RECT 117.200 112.100 117.600 113.900 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 120.600 114.100 121.000 114.200 ;
        RECT 124.100 114.100 124.900 114.200 ;
        RECT 120.600 113.800 121.700 114.100 ;
        RECT 119.800 113.200 120.100 113.800 ;
        RECT 119.800 112.400 120.200 113.200 ;
        RECT 118.200 112.100 118.600 112.200 ;
        RECT 120.700 112.100 121.000 113.800 ;
        RECT 121.400 113.200 121.700 113.800 ;
        RECT 124.000 113.900 124.900 114.100 ;
        RECT 121.400 112.800 121.800 113.200 ;
        RECT 115.000 111.100 115.400 112.100 ;
        RECT 117.200 111.800 118.600 112.100 ;
        RECT 117.200 111.100 117.600 111.800 ;
        RECT 120.600 111.100 121.000 112.100 ;
        RECT 124.000 111.100 124.400 113.900 ;
        RECT 126.200 113.100 126.600 119.900 ;
        RECT 127.800 116.200 128.200 119.900 ;
        RECT 129.400 116.400 129.800 119.900 ;
        RECT 127.800 115.900 129.100 116.200 ;
        RECT 129.400 115.900 129.900 116.400 ;
        RECT 127.800 114.800 128.300 115.200 ;
        RECT 127.900 114.400 128.300 114.800 ;
        RECT 128.800 114.900 129.100 115.900 ;
        RECT 128.800 114.500 129.300 114.900 ;
        RECT 127.000 113.400 127.400 114.200 ;
        RECT 128.800 113.700 129.100 114.500 ;
        RECT 129.600 114.200 129.900 115.900 ;
        RECT 129.400 113.800 129.900 114.200 ;
        RECT 127.800 113.400 129.100 113.700 ;
        RECT 125.700 112.800 126.600 113.100 ;
        RECT 125.700 112.200 126.100 112.800 ;
        RECT 125.700 111.800 126.600 112.200 ;
        RECT 125.700 111.100 126.100 111.800 ;
        RECT 127.800 111.100 128.200 113.400 ;
        RECT 129.600 113.100 129.900 113.800 ;
        RECT 129.400 112.800 129.900 113.100 ;
        RECT 131.000 115.600 131.400 119.900 ;
        RECT 133.100 117.900 133.700 119.900 ;
        RECT 135.400 117.900 135.800 119.900 ;
        RECT 137.600 118.200 138.000 119.900 ;
        RECT 137.600 117.900 138.600 118.200 ;
        RECT 133.400 117.500 133.800 117.900 ;
        RECT 135.500 117.600 135.800 117.900 ;
        RECT 135.100 117.300 136.900 117.600 ;
        RECT 138.200 117.500 138.600 117.900 ;
        RECT 135.100 117.200 135.500 117.300 ;
        RECT 136.500 117.200 136.900 117.300 ;
        RECT 133.000 116.600 133.700 117.000 ;
        RECT 133.400 116.100 133.700 116.600 ;
        RECT 134.500 116.500 135.600 116.800 ;
        RECT 134.500 116.400 134.900 116.500 ;
        RECT 133.400 115.800 134.600 116.100 ;
        RECT 131.000 115.300 133.100 115.600 ;
        RECT 131.000 113.600 131.400 115.300 ;
        RECT 132.700 115.200 133.100 115.300 ;
        RECT 131.900 114.900 132.300 115.000 ;
        RECT 131.900 114.600 133.800 114.900 ;
        RECT 133.400 114.500 133.800 114.600 ;
        RECT 134.300 114.200 134.600 115.800 ;
        RECT 135.300 115.900 135.600 116.500 ;
        RECT 135.900 116.500 136.300 116.600 ;
        RECT 138.200 116.500 138.600 116.600 ;
        RECT 135.900 116.200 138.600 116.500 ;
        RECT 135.300 115.700 137.700 115.900 ;
        RECT 139.800 115.700 140.200 119.900 ;
        RECT 135.300 115.600 140.200 115.700 ;
        RECT 137.300 115.500 140.200 115.600 ;
        RECT 137.400 115.400 140.200 115.500 ;
        RECT 136.600 115.100 137.000 115.200 ;
        RECT 143.000 115.100 143.400 119.900 ;
        RECT 145.000 116.800 145.400 117.200 ;
        RECT 143.800 115.800 144.200 116.600 ;
        RECT 145.000 116.200 145.300 116.800 ;
        RECT 145.700 116.200 146.100 119.900 ;
        RECT 144.600 115.900 145.300 116.200 ;
        RECT 145.600 115.900 146.100 116.200 ;
        RECT 144.600 115.800 145.000 115.900 ;
        RECT 144.600 115.100 144.900 115.800 ;
        RECT 136.600 114.800 139.100 115.100 ;
        RECT 137.400 114.700 137.800 114.800 ;
        RECT 138.700 114.700 139.100 114.800 ;
        RECT 143.000 114.800 144.900 115.100 ;
        RECT 137.900 114.200 138.300 114.300 ;
        RECT 134.300 113.900 139.800 114.200 ;
        RECT 134.500 113.800 134.900 113.900 ;
        RECT 131.000 113.300 132.900 113.600 ;
        RECT 129.400 111.100 129.800 112.800 ;
        RECT 131.000 111.100 131.400 113.300 ;
        RECT 132.500 113.200 132.900 113.300 ;
        RECT 137.400 112.800 137.700 113.900 ;
        RECT 139.000 113.800 139.800 113.900 ;
        RECT 136.500 112.700 136.900 112.800 ;
        RECT 133.400 112.100 133.800 112.500 ;
        RECT 135.500 112.400 136.900 112.700 ;
        RECT 137.400 112.400 137.800 112.800 ;
        RECT 135.500 112.100 135.800 112.400 ;
        RECT 138.200 112.100 138.600 112.500 ;
        RECT 133.100 111.800 133.800 112.100 ;
        RECT 133.100 111.100 133.700 111.800 ;
        RECT 135.400 111.100 135.800 112.100 ;
        RECT 137.600 111.800 138.600 112.100 ;
        RECT 137.600 111.100 138.000 111.800 ;
        RECT 139.800 111.100 140.200 113.500 ;
        RECT 142.200 113.400 142.600 114.200 ;
        RECT 143.000 113.100 143.400 114.800 ;
        RECT 145.600 114.200 145.900 115.900 ;
        RECT 146.200 114.400 146.600 115.200 ;
        RECT 148.600 115.100 149.000 119.900 ;
        RECT 150.700 115.900 151.700 119.900 ;
        RECT 150.200 115.100 150.600 115.200 ;
        RECT 148.600 114.800 150.600 115.100 ;
        RECT 144.600 113.800 145.900 114.200 ;
        RECT 147.000 114.100 147.400 114.200 ;
        RECT 146.600 113.800 147.400 114.100 ;
        RECT 144.700 113.100 145.000 113.800 ;
        RECT 146.600 113.600 147.000 113.800 ;
        RECT 145.500 113.100 147.300 113.300 ;
        RECT 143.000 112.800 143.900 113.100 ;
        RECT 143.500 111.100 143.900 112.800 ;
        RECT 144.600 111.100 145.000 113.100 ;
        RECT 145.400 113.000 147.400 113.100 ;
        RECT 145.400 111.100 145.800 113.000 ;
        RECT 147.000 111.100 147.400 113.000 ;
        RECT 147.800 112.400 148.200 113.200 ;
        RECT 148.600 111.100 149.000 114.800 ;
        RECT 150.200 114.400 150.600 114.800 ;
        RECT 151.000 114.200 151.300 115.900 ;
        RECT 153.400 115.800 153.800 116.600 ;
        RECT 151.800 114.400 152.200 115.200 ;
        RECT 149.400 114.100 149.800 114.200 ;
        RECT 151.000 114.100 151.400 114.200 ;
        RECT 152.600 114.100 153.000 114.600 ;
        RECT 153.400 114.100 153.800 114.200 ;
        RECT 149.400 113.800 150.200 114.100 ;
        RECT 151.000 113.800 152.200 114.100 ;
        RECT 152.600 113.800 153.800 114.100 ;
        RECT 149.800 113.600 150.200 113.800 ;
        RECT 149.500 113.100 151.300 113.300 ;
        RECT 151.900 113.100 152.200 113.800 ;
        RECT 154.200 113.100 154.600 119.900 ;
        RECT 156.200 116.800 156.600 117.200 ;
        RECT 156.200 116.200 156.500 116.800 ;
        RECT 156.900 116.200 157.300 119.900 ;
        RECT 155.800 115.900 156.500 116.200 ;
        RECT 156.800 115.900 157.300 116.200 ;
        RECT 155.800 115.800 156.200 115.900 ;
        RECT 156.800 114.200 157.100 115.900 ;
        RECT 157.400 114.400 157.800 115.200 ;
        RECT 155.000 113.400 155.400 114.200 ;
        RECT 155.800 113.800 157.100 114.200 ;
        RECT 158.200 114.100 158.600 114.200 ;
        RECT 157.800 113.800 158.600 114.100 ;
        RECT 155.900 113.100 156.200 113.800 ;
        RECT 157.800 113.600 158.200 113.800 ;
        RECT 159.000 113.400 159.400 114.200 ;
        RECT 156.700 113.100 158.500 113.300 ;
        RECT 159.800 113.100 160.200 119.900 ;
        RECT 160.600 115.800 161.000 116.600 ;
        RECT 162.200 113.100 162.600 119.900 ;
        RECT 163.000 115.800 163.400 116.600 ;
        RECT 163.800 116.200 164.200 119.900 ;
        RECT 165.400 116.200 165.800 119.900 ;
        RECT 163.800 115.900 165.800 116.200 ;
        RECT 166.200 115.800 166.600 119.900 ;
        RECT 167.000 116.200 167.400 119.900 ;
        RECT 168.600 116.200 169.000 119.900 ;
        RECT 167.000 115.900 169.000 116.200 ;
        RECT 169.400 115.900 169.800 119.900 ;
        RECT 171.000 116.400 171.400 119.900 ;
        RECT 170.900 115.900 171.400 116.400 ;
        RECT 172.600 116.200 173.000 119.900 ;
        RECT 173.800 116.800 174.200 117.200 ;
        RECT 173.800 116.200 174.100 116.800 ;
        RECT 174.500 116.200 174.900 119.900 ;
        RECT 171.700 115.900 173.000 116.200 ;
        RECT 173.400 115.900 174.100 116.200 ;
        RECT 164.200 115.200 164.600 115.400 ;
        RECT 166.200 115.200 166.500 115.800 ;
        RECT 167.400 115.200 167.800 115.400 ;
        RECT 169.400 115.200 169.700 115.900 ;
        RECT 163.800 114.900 164.600 115.200 ;
        RECT 165.400 114.900 166.600 115.200 ;
        RECT 163.800 114.800 164.200 114.900 ;
        RECT 164.600 113.800 165.000 114.600 ;
        RECT 165.400 113.100 165.700 114.900 ;
        RECT 166.200 114.800 166.600 114.900 ;
        RECT 167.000 114.900 167.800 115.200 ;
        RECT 168.600 114.900 169.800 115.200 ;
        RECT 167.000 114.800 167.400 114.900 ;
        RECT 167.800 113.800 168.200 114.600 ;
        RECT 168.600 113.100 168.900 114.900 ;
        RECT 169.400 114.800 169.800 114.900 ;
        RECT 170.900 114.200 171.200 115.900 ;
        RECT 171.700 114.900 172.000 115.900 ;
        RECT 173.400 115.800 173.800 115.900 ;
        RECT 174.400 115.800 175.400 116.200 ;
        RECT 176.600 115.900 177.000 119.900 ;
        RECT 177.400 116.200 177.800 119.900 ;
        RECT 179.000 116.200 179.400 119.900 ;
        RECT 181.100 116.200 181.500 119.900 ;
        RECT 181.800 116.800 182.200 117.200 ;
        RECT 181.900 116.200 182.200 116.800 ;
        RECT 177.400 115.900 179.400 116.200 ;
        RECT 171.500 114.500 172.000 114.900 ;
        RECT 170.900 113.800 171.400 114.200 ;
        RECT 170.900 113.100 171.200 113.800 ;
        RECT 171.700 113.700 172.000 114.500 ;
        RECT 172.500 115.100 173.000 115.200 ;
        RECT 173.400 115.100 173.800 115.200 ;
        RECT 172.500 114.800 173.800 115.100 ;
        RECT 172.500 114.400 172.900 114.800 ;
        RECT 174.400 114.200 174.700 115.800 ;
        RECT 176.700 115.200 177.000 115.900 ;
        RECT 180.600 115.800 181.600 116.200 ;
        RECT 181.900 115.900 182.600 116.200 ;
        RECT 182.200 115.800 182.600 115.900 ;
        RECT 183.000 115.800 183.400 116.600 ;
        RECT 178.600 115.200 179.000 115.400 ;
        RECT 175.000 115.100 175.400 115.200 ;
        RECT 176.600 115.100 177.800 115.200 ;
        RECT 175.000 114.900 177.800 115.100 ;
        RECT 178.600 115.100 179.400 115.200 ;
        RECT 179.800 115.100 180.200 115.200 ;
        RECT 178.600 114.900 180.200 115.100 ;
        RECT 175.000 114.800 177.000 114.900 ;
        RECT 175.000 114.400 175.400 114.800 ;
        RECT 173.400 113.800 174.700 114.200 ;
        RECT 175.800 114.100 176.200 114.200 ;
        RECT 175.400 113.800 176.200 114.100 ;
        RECT 171.700 113.400 173.000 113.700 ;
        RECT 149.400 113.000 151.400 113.100 ;
        RECT 149.400 111.100 149.800 113.000 ;
        RECT 151.000 111.400 151.400 113.000 ;
        RECT 151.800 111.700 152.200 113.100 ;
        RECT 152.600 111.400 153.000 113.100 ;
        RECT 151.000 111.100 153.000 111.400 ;
        RECT 153.700 112.800 154.600 113.100 ;
        RECT 153.700 112.200 154.100 112.800 ;
        RECT 153.700 111.800 154.600 112.200 ;
        RECT 153.700 111.100 154.100 111.800 ;
        RECT 155.800 111.100 156.200 113.100 ;
        RECT 156.600 113.000 158.600 113.100 ;
        RECT 156.600 111.100 157.000 113.000 ;
        RECT 158.200 111.100 158.600 113.000 ;
        RECT 159.800 112.800 160.700 113.100 ;
        RECT 162.200 112.800 163.100 113.100 ;
        RECT 160.300 112.200 160.700 112.800 ;
        RECT 160.300 111.800 161.000 112.200 ;
        RECT 160.300 111.100 160.700 111.800 ;
        RECT 162.700 111.100 163.100 112.800 ;
        RECT 165.400 111.100 165.800 113.100 ;
        RECT 168.600 111.100 169.000 113.100 ;
        RECT 170.900 112.800 171.400 113.100 ;
        RECT 171.000 111.100 171.400 112.800 ;
        RECT 172.600 111.100 173.000 113.400 ;
        RECT 173.500 113.100 173.800 113.800 ;
        RECT 175.400 113.600 175.800 113.800 ;
        RECT 174.300 113.100 176.100 113.300 ;
        RECT 173.400 111.100 173.800 113.100 ;
        RECT 174.200 113.000 176.200 113.100 ;
        RECT 174.200 111.100 174.600 113.000 ;
        RECT 175.800 111.100 176.200 113.000 ;
        RECT 176.600 112.800 177.000 113.200 ;
        RECT 177.500 113.100 177.800 114.900 ;
        RECT 179.000 114.800 180.200 114.900 ;
        RECT 178.200 113.800 178.600 114.600 ;
        RECT 180.600 114.400 181.000 115.200 ;
        RECT 181.300 114.200 181.600 115.800 ;
        RECT 179.800 114.100 180.200 114.200 ;
        RECT 179.800 113.800 180.600 114.100 ;
        RECT 181.300 113.800 182.600 114.200 ;
        RECT 180.200 113.600 180.600 113.800 ;
        RECT 179.900 113.100 181.700 113.300 ;
        RECT 182.200 113.100 182.500 113.800 ;
        RECT 183.800 113.100 184.200 119.900 ;
        RECT 185.400 116.200 185.800 119.900 ;
        RECT 187.000 116.200 187.400 119.900 ;
        RECT 185.400 115.900 187.400 116.200 ;
        RECT 187.800 115.900 188.200 119.900 ;
        RECT 189.000 116.800 189.400 117.200 ;
        RECT 189.000 116.200 189.300 116.800 ;
        RECT 189.700 116.200 190.100 119.900 ;
        RECT 188.600 115.900 189.300 116.200 ;
        RECT 189.600 115.900 190.100 116.200 ;
        RECT 185.800 115.200 186.200 115.400 ;
        RECT 187.800 115.200 188.100 115.900 ;
        RECT 188.600 115.800 189.000 115.900 ;
        RECT 185.400 114.900 186.200 115.200 ;
        RECT 187.000 115.100 188.200 115.200 ;
        RECT 188.600 115.100 189.000 115.200 ;
        RECT 187.000 114.900 189.000 115.100 ;
        RECT 185.400 114.800 185.800 114.900 ;
        RECT 184.600 113.400 185.000 114.200 ;
        RECT 186.200 113.800 186.600 114.600 ;
        RECT 176.700 112.400 177.100 112.800 ;
        RECT 177.400 111.100 177.800 113.100 ;
        RECT 179.800 113.000 181.800 113.100 ;
        RECT 179.800 111.100 180.200 113.000 ;
        RECT 181.400 111.100 181.800 113.000 ;
        RECT 182.200 111.100 182.600 113.100 ;
        RECT 183.300 112.800 184.200 113.100 ;
        RECT 187.000 113.100 187.300 114.900 ;
        RECT 187.800 114.800 189.000 114.900 ;
        RECT 189.600 114.200 189.900 115.900 ;
        RECT 193.400 115.700 193.800 119.900 ;
        RECT 195.600 118.200 196.000 119.900 ;
        RECT 195.000 117.900 196.000 118.200 ;
        RECT 197.800 117.900 198.200 119.900 ;
        RECT 199.900 117.900 200.500 119.900 ;
        RECT 195.000 117.500 195.400 117.900 ;
        RECT 197.800 117.600 198.100 117.900 ;
        RECT 196.700 117.300 198.500 117.600 ;
        RECT 199.800 117.500 200.200 117.900 ;
        RECT 196.700 117.200 197.100 117.300 ;
        RECT 198.100 117.200 198.500 117.300 ;
        RECT 195.000 116.500 195.400 116.600 ;
        RECT 197.300 116.500 197.700 116.600 ;
        RECT 195.000 116.200 197.700 116.500 ;
        RECT 198.000 116.500 199.100 116.800 ;
        RECT 198.000 115.900 198.300 116.500 ;
        RECT 198.700 116.400 199.100 116.500 ;
        RECT 199.900 116.600 200.600 117.000 ;
        RECT 199.900 116.100 200.200 116.600 ;
        RECT 195.900 115.700 198.300 115.900 ;
        RECT 193.400 115.600 198.300 115.700 ;
        RECT 199.000 115.800 200.200 116.100 ;
        RECT 193.400 115.500 196.300 115.600 ;
        RECT 193.400 115.400 196.200 115.500 ;
        RECT 190.200 115.100 190.600 115.200 ;
        RECT 192.600 115.100 193.000 115.200 ;
        RECT 196.600 115.100 197.000 115.200 ;
        RECT 190.200 114.800 193.000 115.100 ;
        RECT 194.500 114.800 197.000 115.100 ;
        RECT 190.200 114.400 190.600 114.800 ;
        RECT 194.500 114.700 194.900 114.800 ;
        RECT 195.800 114.700 196.200 114.800 ;
        RECT 195.300 114.200 195.700 114.300 ;
        RECT 199.000 114.200 199.300 115.800 ;
        RECT 202.200 115.600 202.600 119.900 ;
        RECT 204.900 116.400 205.300 119.900 ;
        RECT 207.000 117.500 207.400 119.500 ;
        RECT 204.500 116.100 205.300 116.400 ;
        RECT 200.500 115.300 202.600 115.600 ;
        RECT 200.500 115.200 200.900 115.300 ;
        RECT 201.300 114.900 201.700 115.000 ;
        RECT 199.800 114.600 201.700 114.900 ;
        RECT 199.800 114.500 200.200 114.600 ;
        RECT 188.600 113.800 189.900 114.200 ;
        RECT 191.000 114.100 191.400 114.200 ;
        RECT 191.800 114.100 192.200 114.200 ;
        RECT 190.600 113.800 192.200 114.100 ;
        RECT 193.800 113.900 199.300 114.200 ;
        RECT 193.800 113.800 194.600 113.900 ;
        RECT 187.800 113.100 188.200 113.200 ;
        RECT 188.700 113.100 189.000 113.800 ;
        RECT 190.600 113.600 191.000 113.800 ;
        RECT 189.500 113.100 191.300 113.300 ;
        RECT 183.300 112.200 183.700 112.800 ;
        RECT 183.000 111.800 183.700 112.200 ;
        RECT 183.300 111.100 183.700 111.800 ;
        RECT 187.000 111.100 187.400 113.100 ;
        RECT 187.800 112.800 189.000 113.100 ;
        RECT 187.700 112.400 188.100 112.800 ;
        RECT 188.600 111.100 189.000 112.800 ;
        RECT 189.400 113.000 191.400 113.100 ;
        RECT 189.400 111.100 189.800 113.000 ;
        RECT 191.000 111.100 191.400 113.000 ;
        RECT 193.400 111.100 193.800 113.500 ;
        RECT 195.900 112.800 196.200 113.900 ;
        RECT 196.600 113.800 197.000 113.900 ;
        RECT 198.700 113.800 199.100 113.900 ;
        RECT 202.200 113.600 202.600 115.300 ;
        RECT 203.800 114.800 204.200 115.600 ;
        RECT 204.500 114.200 204.800 116.100 ;
        RECT 207.100 115.800 207.400 117.500 ;
        RECT 205.500 115.500 207.400 115.800 ;
        RECT 205.500 114.500 205.800 115.500 ;
        RECT 203.000 114.100 203.400 114.200 ;
        RECT 203.800 114.100 204.800 114.200 ;
        RECT 205.100 114.100 205.800 114.500 ;
        RECT 206.200 114.400 206.600 115.200 ;
        RECT 207.000 114.400 207.400 115.200 ;
        RECT 203.000 113.800 204.800 114.100 ;
        RECT 200.700 113.300 202.600 113.600 ;
        RECT 200.700 113.200 201.100 113.300 ;
        RECT 195.000 112.100 195.400 112.500 ;
        RECT 195.800 112.400 196.200 112.800 ;
        RECT 196.700 112.700 197.100 112.800 ;
        RECT 196.700 112.400 198.100 112.700 ;
        RECT 197.800 112.100 198.100 112.400 ;
        RECT 199.800 112.100 200.200 112.500 ;
        RECT 195.000 111.800 196.000 112.100 ;
        RECT 195.600 111.100 196.000 111.800 ;
        RECT 197.800 111.100 198.200 112.100 ;
        RECT 199.800 111.800 200.500 112.100 ;
        RECT 199.900 111.100 200.500 111.800 ;
        RECT 202.200 111.100 202.600 113.300 ;
        RECT 204.500 113.500 204.800 113.800 ;
        RECT 205.300 113.900 205.800 114.100 ;
        RECT 205.300 113.600 207.400 113.900 ;
        RECT 204.500 113.300 204.900 113.500 ;
        RECT 204.500 113.000 205.300 113.300 ;
        RECT 204.900 111.500 205.300 113.000 ;
        RECT 207.100 112.500 207.400 113.600 ;
        RECT 207.800 113.400 208.200 114.200 ;
        RECT 208.600 113.100 209.000 119.900 ;
        RECT 209.400 115.800 209.800 116.600 ;
        RECT 210.200 115.600 210.600 119.900 ;
        RECT 212.300 117.900 212.900 119.900 ;
        RECT 214.600 117.900 215.000 119.900 ;
        RECT 216.800 118.200 217.200 119.900 ;
        RECT 216.800 117.900 217.800 118.200 ;
        RECT 212.600 117.500 213.000 117.900 ;
        RECT 214.700 117.600 215.000 117.900 ;
        RECT 214.300 117.300 216.100 117.600 ;
        RECT 217.400 117.500 217.800 117.900 ;
        RECT 214.300 117.200 214.700 117.300 ;
        RECT 215.700 117.200 216.100 117.300 ;
        RECT 212.200 116.600 212.900 117.000 ;
        RECT 212.600 116.100 212.900 116.600 ;
        RECT 213.700 116.500 214.800 116.800 ;
        RECT 213.700 116.400 214.100 116.500 ;
        RECT 212.600 115.800 213.800 116.100 ;
        RECT 210.200 115.300 212.300 115.600 ;
        RECT 210.200 113.600 210.600 115.300 ;
        RECT 211.900 115.200 212.300 115.300 ;
        RECT 211.100 114.900 211.500 115.000 ;
        RECT 211.100 114.600 213.000 114.900 ;
        RECT 212.600 114.500 213.000 114.600 ;
        RECT 213.500 114.200 213.800 115.800 ;
        RECT 214.500 115.900 214.800 116.500 ;
        RECT 215.100 116.500 215.500 116.600 ;
        RECT 217.400 116.500 217.800 116.600 ;
        RECT 215.100 116.200 217.800 116.500 ;
        RECT 214.500 115.700 216.900 115.900 ;
        RECT 219.000 115.700 219.400 119.900 ;
        RECT 214.500 115.600 219.400 115.700 ;
        RECT 216.500 115.500 219.400 115.600 ;
        RECT 216.600 115.400 219.400 115.500 ;
        RECT 219.800 115.700 220.200 119.900 ;
        RECT 222.000 118.200 222.400 119.900 ;
        RECT 221.400 117.900 222.400 118.200 ;
        RECT 224.200 117.900 224.600 119.900 ;
        RECT 226.300 117.900 226.900 119.900 ;
        RECT 221.400 117.500 221.800 117.900 ;
        RECT 224.200 117.600 224.500 117.900 ;
        RECT 223.100 117.300 224.900 117.600 ;
        RECT 226.200 117.500 226.600 117.900 ;
        RECT 223.100 117.200 223.500 117.300 ;
        RECT 224.500 117.200 224.900 117.300 ;
        RECT 221.400 116.500 221.800 116.600 ;
        RECT 223.700 116.500 224.100 116.600 ;
        RECT 221.400 116.200 224.100 116.500 ;
        RECT 224.400 116.500 225.500 116.800 ;
        RECT 224.400 115.900 224.700 116.500 ;
        RECT 225.100 116.400 225.500 116.500 ;
        RECT 226.300 116.600 227.000 117.000 ;
        RECT 226.300 116.100 226.600 116.600 ;
        RECT 222.300 115.700 224.700 115.900 ;
        RECT 219.800 115.600 224.700 115.700 ;
        RECT 225.400 115.800 226.600 116.100 ;
        RECT 219.800 115.500 222.700 115.600 ;
        RECT 219.800 115.400 222.600 115.500 ;
        RECT 215.800 115.100 216.200 115.200 ;
        RECT 223.000 115.100 223.400 115.200 ;
        RECT 215.800 114.800 218.300 115.100 ;
        RECT 216.600 114.700 217.000 114.800 ;
        RECT 217.900 114.700 218.300 114.800 ;
        RECT 220.900 114.800 223.400 115.100 ;
        RECT 220.900 114.700 221.300 114.800 ;
        RECT 217.100 114.200 217.500 114.300 ;
        RECT 221.700 114.200 222.100 114.300 ;
        RECT 225.400 114.200 225.700 115.800 ;
        RECT 228.600 115.600 229.000 119.900 ;
        RECT 226.900 115.300 229.000 115.600 ;
        RECT 226.900 115.200 227.300 115.300 ;
        RECT 227.700 114.900 228.100 115.000 ;
        RECT 226.200 114.600 228.100 114.900 ;
        RECT 226.200 114.500 226.600 114.600 ;
        RECT 213.500 113.900 219.000 114.200 ;
        RECT 213.700 113.800 214.100 113.900 ;
        RECT 210.200 113.300 212.100 113.600 ;
        RECT 208.600 112.800 209.500 113.100 ;
        RECT 207.000 111.500 207.400 112.500 ;
        RECT 209.100 112.200 209.500 112.800 ;
        RECT 208.600 111.800 209.500 112.200 ;
        RECT 209.100 111.100 209.500 111.800 ;
        RECT 210.200 111.100 210.600 113.300 ;
        RECT 211.700 113.200 212.100 113.300 ;
        RECT 216.600 113.200 216.900 113.900 ;
        RECT 218.200 113.800 219.000 113.900 ;
        RECT 220.200 113.900 225.700 114.200 ;
        RECT 220.200 113.800 221.000 113.900 ;
        RECT 215.700 112.700 216.100 112.800 ;
        RECT 212.600 112.100 213.000 112.500 ;
        RECT 214.700 112.400 216.100 112.700 ;
        RECT 216.600 112.400 217.000 113.200 ;
        RECT 214.700 112.100 215.000 112.400 ;
        RECT 217.400 112.100 217.800 112.500 ;
        RECT 212.300 111.800 213.000 112.100 ;
        RECT 212.300 111.100 212.900 111.800 ;
        RECT 214.600 111.100 215.000 112.100 ;
        RECT 216.800 111.800 217.800 112.100 ;
        RECT 216.800 111.100 217.200 111.800 ;
        RECT 219.000 111.100 219.400 113.500 ;
        RECT 219.800 111.100 220.200 113.500 ;
        RECT 222.300 113.200 222.600 113.900 ;
        RECT 225.100 113.800 225.500 113.900 ;
        RECT 228.600 113.600 229.000 115.300 ;
        RECT 227.100 113.300 229.000 113.600 ;
        RECT 227.100 113.200 227.500 113.300 ;
        RECT 221.400 112.100 221.800 112.500 ;
        RECT 222.200 112.400 222.600 113.200 ;
        RECT 223.100 112.700 223.500 112.800 ;
        RECT 223.100 112.400 224.500 112.700 ;
        RECT 224.200 112.100 224.500 112.400 ;
        RECT 226.200 112.100 226.600 112.500 ;
        RECT 221.400 111.800 222.400 112.100 ;
        RECT 222.000 111.100 222.400 111.800 ;
        RECT 224.200 111.100 224.600 112.100 ;
        RECT 226.200 111.800 226.900 112.100 ;
        RECT 226.300 111.100 226.900 111.800 ;
        RECT 228.600 111.100 229.000 113.300 ;
        RECT 0.900 109.200 1.300 109.900 ;
        RECT 0.900 108.800 1.800 109.200 ;
        RECT 0.900 108.200 1.300 108.800 ;
        RECT 0.900 107.900 1.800 108.200 ;
        RECT 0.600 104.400 1.000 105.200 ;
        RECT 1.400 101.100 1.800 107.900 ;
        RECT 3.000 107.800 3.400 108.600 ;
        RECT 2.200 107.100 2.600 107.600 ;
        RECT 2.200 106.800 3.300 107.100 ;
        RECT 3.000 106.200 3.300 106.800 ;
        RECT 3.000 105.800 3.400 106.200 ;
        RECT 3.800 106.100 4.200 109.900 ;
        RECT 5.900 108.200 6.300 109.900 ;
        RECT 5.400 107.900 6.300 108.200 ;
        RECT 7.000 107.900 7.400 109.900 ;
        RECT 7.800 108.000 8.200 109.900 ;
        RECT 9.400 108.000 9.800 109.900 ;
        RECT 7.800 107.900 9.800 108.000 ;
        RECT 4.600 106.800 5.000 107.600 ;
        RECT 5.400 106.100 5.800 107.900 ;
        RECT 7.100 107.200 7.400 107.900 ;
        RECT 7.900 107.700 9.700 107.900 ;
        RECT 10.200 107.500 10.600 109.900 ;
        RECT 12.400 109.200 12.800 109.900 ;
        RECT 11.800 108.900 12.800 109.200 ;
        RECT 14.600 108.900 15.000 109.900 ;
        RECT 16.700 109.200 17.300 109.900 ;
        RECT 16.600 108.900 17.300 109.200 ;
        RECT 11.800 108.500 12.200 108.900 ;
        RECT 14.600 108.600 14.900 108.900 ;
        RECT 12.600 108.200 13.000 108.600 ;
        RECT 13.500 108.300 14.900 108.600 ;
        RECT 16.600 108.500 17.000 108.900 ;
        RECT 13.500 108.200 13.900 108.300 ;
        RECT 9.000 107.200 9.400 107.400 ;
        RECT 7.000 106.800 8.300 107.200 ;
        RECT 9.000 106.900 9.800 107.200 ;
        RECT 9.400 106.800 9.800 106.900 ;
        RECT 10.600 107.100 11.400 107.200 ;
        RECT 12.700 107.100 13.000 108.200 ;
        RECT 17.500 107.700 17.900 107.800 ;
        RECT 19.000 107.700 19.400 109.900 ;
        RECT 19.800 108.000 20.200 109.900 ;
        RECT 21.400 108.000 21.800 109.900 ;
        RECT 19.800 107.900 21.800 108.000 ;
        RECT 22.200 107.900 22.600 109.900 ;
        RECT 23.300 108.200 23.700 109.900 ;
        RECT 23.300 107.900 24.200 108.200 ;
        RECT 25.400 108.000 25.800 109.900 ;
        RECT 27.000 108.000 27.400 109.900 ;
        RECT 25.400 107.900 27.400 108.000 ;
        RECT 27.800 107.900 28.200 109.900 ;
        RECT 29.400 108.200 29.800 109.900 ;
        RECT 29.300 107.900 29.800 108.200 ;
        RECT 19.900 107.700 21.700 107.900 ;
        RECT 17.500 107.400 19.400 107.700 ;
        RECT 15.500 107.100 15.900 107.200 ;
        RECT 10.600 106.800 16.100 107.100 ;
        RECT 3.800 105.800 4.900 106.100 ;
        RECT 3.800 101.100 4.200 105.800 ;
        RECT 4.600 105.200 4.900 105.800 ;
        RECT 5.400 105.800 7.300 106.100 ;
        RECT 4.600 104.800 5.000 105.200 ;
        RECT 5.400 101.100 5.800 105.800 ;
        RECT 7.000 105.200 7.300 105.800 ;
        RECT 8.000 105.200 8.300 106.800 ;
        RECT 12.100 106.700 12.500 106.800 ;
        RECT 8.600 106.100 9.000 106.600 ;
        RECT 11.300 106.200 11.700 106.300 ;
        RECT 9.400 106.100 9.800 106.200 ;
        RECT 8.600 105.800 9.800 106.100 ;
        RECT 11.300 106.100 13.800 106.200 ;
        RECT 15.000 106.100 15.400 106.200 ;
        RECT 11.300 105.900 15.400 106.100 ;
        RECT 13.400 105.800 15.400 105.900 ;
        RECT 10.200 105.500 13.000 105.600 ;
        RECT 10.200 105.400 13.100 105.500 ;
        RECT 10.200 105.300 15.100 105.400 ;
        RECT 6.200 104.400 6.600 105.200 ;
        RECT 7.000 105.100 7.400 105.200 ;
        RECT 7.000 104.800 7.700 105.100 ;
        RECT 8.000 104.800 9.000 105.200 ;
        RECT 7.400 104.200 7.700 104.800 ;
        RECT 7.400 103.800 7.800 104.200 ;
        RECT 8.100 101.100 8.500 104.800 ;
        RECT 10.200 101.100 10.600 105.300 ;
        RECT 12.700 105.100 15.100 105.300 ;
        RECT 11.800 104.500 14.500 104.800 ;
        RECT 11.800 104.400 12.200 104.500 ;
        RECT 14.100 104.400 14.500 104.500 ;
        RECT 14.800 104.500 15.100 105.100 ;
        RECT 15.800 105.200 16.100 106.800 ;
        RECT 16.600 106.400 17.000 106.500 ;
        RECT 16.600 106.100 18.500 106.400 ;
        RECT 18.100 106.000 18.500 106.100 ;
        RECT 17.300 105.700 17.700 105.800 ;
        RECT 19.000 105.700 19.400 107.400 ;
        RECT 20.200 107.200 20.600 107.400 ;
        RECT 22.200 107.200 22.500 107.900 ;
        RECT 19.800 106.900 20.600 107.200 ;
        RECT 19.800 106.800 20.200 106.900 ;
        RECT 21.300 106.800 22.600 107.200 ;
        RECT 20.600 105.800 21.000 106.600 ;
        RECT 21.300 106.200 21.600 106.800 ;
        RECT 21.300 105.800 21.800 106.200 ;
        RECT 23.800 106.100 24.200 107.900 ;
        RECT 25.500 107.700 27.300 107.900 ;
        RECT 24.600 106.800 25.000 107.600 ;
        RECT 25.800 107.200 26.200 107.400 ;
        RECT 27.800 107.200 28.100 107.900 ;
        RECT 29.300 107.200 29.600 107.900 ;
        RECT 31.000 107.600 31.400 109.900 ;
        RECT 31.800 107.800 32.200 108.600 ;
        RECT 30.100 107.300 31.400 107.600 ;
        RECT 25.400 106.900 26.200 107.200 ;
        RECT 25.400 106.800 25.800 106.900 ;
        RECT 26.900 106.800 28.200 107.200 ;
        RECT 29.300 106.800 29.800 107.200 ;
        RECT 22.200 105.800 24.200 106.100 ;
        RECT 26.200 105.800 26.600 106.600 ;
        RECT 17.300 105.400 19.400 105.700 ;
        RECT 15.800 104.900 17.000 105.200 ;
        RECT 15.500 104.500 15.900 104.600 ;
        RECT 14.800 104.200 15.900 104.500 ;
        RECT 16.700 104.400 17.000 104.900 ;
        RECT 16.700 104.000 17.400 104.400 ;
        RECT 13.500 103.700 13.900 103.800 ;
        RECT 14.900 103.700 15.300 103.800 ;
        RECT 11.800 103.100 12.200 103.500 ;
        RECT 13.500 103.400 15.300 103.700 ;
        RECT 14.600 103.100 14.900 103.400 ;
        RECT 16.600 103.100 17.000 103.500 ;
        RECT 11.800 102.800 12.800 103.100 ;
        RECT 12.400 101.100 12.800 102.800 ;
        RECT 14.600 101.100 15.000 103.100 ;
        RECT 16.700 101.100 17.300 103.100 ;
        RECT 19.000 101.100 19.400 105.400 ;
        RECT 21.300 105.100 21.600 105.800 ;
        RECT 22.200 105.200 22.500 105.800 ;
        RECT 22.200 105.100 22.600 105.200 ;
        RECT 21.100 104.800 21.600 105.100 ;
        RECT 21.900 104.800 22.600 105.100 ;
        RECT 21.100 101.100 21.500 104.800 ;
        RECT 21.900 104.200 22.200 104.800 ;
        RECT 23.000 104.400 23.400 105.200 ;
        RECT 21.800 103.800 22.200 104.200 ;
        RECT 23.800 101.100 24.200 105.800 ;
        RECT 26.900 105.100 27.200 106.800 ;
        RECT 27.800 105.100 28.200 105.200 ;
        RECT 26.700 104.800 27.200 105.100 ;
        RECT 27.500 104.800 28.200 105.100 ;
        RECT 29.300 105.100 29.600 106.800 ;
        RECT 30.100 106.500 30.400 107.300 ;
        RECT 31.800 106.800 32.200 107.200 ;
        RECT 29.900 106.100 30.400 106.500 ;
        RECT 30.100 105.100 30.400 106.100 ;
        RECT 30.900 106.200 31.300 106.600 ;
        RECT 30.900 106.100 31.400 106.200 ;
        RECT 31.800 106.100 32.100 106.800 ;
        RECT 30.900 105.800 32.100 106.100 ;
        RECT 26.700 102.200 27.100 104.800 ;
        RECT 27.500 104.200 27.800 104.800 ;
        RECT 29.300 104.600 29.800 105.100 ;
        RECT 30.100 104.800 31.400 105.100 ;
        RECT 27.400 103.800 27.800 104.200 ;
        RECT 26.200 101.800 27.100 102.200 ;
        RECT 26.700 101.100 27.100 101.800 ;
        RECT 29.400 101.100 29.800 104.600 ;
        RECT 31.000 101.100 31.400 104.800 ;
        RECT 32.600 102.100 33.000 109.900 ;
        RECT 35.000 107.500 35.400 109.900 ;
        RECT 37.200 109.200 37.600 109.900 ;
        RECT 36.600 108.900 37.600 109.200 ;
        RECT 39.400 108.900 39.800 109.900 ;
        RECT 41.500 109.200 42.100 109.900 ;
        RECT 41.400 108.900 42.100 109.200 ;
        RECT 36.600 108.500 37.000 108.900 ;
        RECT 39.400 108.600 39.700 108.900 ;
        RECT 37.400 108.200 37.800 108.600 ;
        RECT 38.300 108.300 39.700 108.600 ;
        RECT 41.400 108.500 41.800 108.900 ;
        RECT 38.300 108.200 38.700 108.300 ;
        RECT 35.400 107.100 36.200 107.200 ;
        RECT 37.500 107.100 37.800 108.200 ;
        RECT 42.200 107.800 42.600 108.200 ;
        RECT 42.200 107.700 42.700 107.800 ;
        RECT 43.800 107.700 44.200 109.900 ;
        RECT 42.200 107.400 44.200 107.700 ;
        RECT 40.300 107.100 40.700 107.200 ;
        RECT 35.400 106.800 40.900 107.100 ;
        RECT 36.900 106.700 37.300 106.800 ;
        RECT 36.100 106.200 36.500 106.300 ;
        RECT 37.400 106.200 37.800 106.300 ;
        RECT 40.600 106.200 40.900 106.800 ;
        RECT 41.400 106.400 41.800 106.500 ;
        RECT 36.100 105.900 38.600 106.200 ;
        RECT 38.200 105.800 38.600 105.900 ;
        RECT 40.600 105.800 41.000 106.200 ;
        RECT 41.400 106.100 43.300 106.400 ;
        RECT 42.900 106.000 43.300 106.100 ;
        RECT 35.000 105.500 37.800 105.600 ;
        RECT 35.000 105.400 37.900 105.500 ;
        RECT 35.000 105.300 39.900 105.400 ;
        RECT 33.400 102.100 33.800 102.200 ;
        RECT 32.600 101.800 33.800 102.100 ;
        RECT 32.600 101.100 33.000 101.800 ;
        RECT 35.000 101.100 35.400 105.300 ;
        RECT 37.500 105.100 39.900 105.300 ;
        RECT 36.600 104.500 39.300 104.800 ;
        RECT 36.600 104.400 37.000 104.500 ;
        RECT 38.900 104.400 39.300 104.500 ;
        RECT 39.600 104.500 39.900 105.100 ;
        RECT 40.600 105.200 40.900 105.800 ;
        RECT 42.100 105.700 42.500 105.800 ;
        RECT 43.800 105.700 44.200 107.400 ;
        RECT 44.600 107.600 45.000 109.900 ;
        RECT 46.200 108.200 46.600 109.900 ;
        RECT 46.200 107.900 46.700 108.200 ;
        RECT 44.600 107.300 45.900 107.600 ;
        RECT 44.700 106.200 45.100 106.600 ;
        RECT 44.600 105.800 45.100 106.200 ;
        RECT 45.600 106.500 45.900 107.300 ;
        RECT 46.400 107.200 46.700 107.900 ;
        RECT 47.800 107.500 48.200 109.900 ;
        RECT 50.000 109.200 50.400 109.900 ;
        RECT 49.400 108.900 50.400 109.200 ;
        RECT 52.200 108.900 52.600 109.900 ;
        RECT 54.300 109.200 54.900 109.900 ;
        RECT 54.200 108.900 54.900 109.200 ;
        RECT 49.400 108.500 49.800 108.900 ;
        RECT 52.200 108.600 52.500 108.900 ;
        RECT 50.200 108.200 50.600 108.600 ;
        RECT 51.100 108.300 52.500 108.600 ;
        RECT 54.200 108.500 54.600 108.900 ;
        RECT 51.100 108.200 51.500 108.300 ;
        RECT 46.200 106.800 46.700 107.200 ;
        RECT 48.200 107.100 49.000 107.200 ;
        RECT 50.300 107.100 50.600 108.200 ;
        RECT 55.100 107.700 55.500 107.800 ;
        RECT 56.600 107.700 57.000 109.900 ;
        RECT 57.400 107.800 57.800 108.600 ;
        RECT 55.100 107.400 57.000 107.700 ;
        RECT 53.100 107.100 53.500 107.200 ;
        RECT 48.200 106.800 53.700 107.100 ;
        RECT 45.600 106.100 46.100 106.500 ;
        RECT 42.100 105.400 44.200 105.700 ;
        RECT 40.600 104.900 41.800 105.200 ;
        RECT 40.300 104.500 40.700 104.600 ;
        RECT 39.600 104.200 40.700 104.500 ;
        RECT 41.500 104.400 41.800 104.900 ;
        RECT 41.500 104.000 42.200 104.400 ;
        RECT 38.300 103.700 38.700 103.800 ;
        RECT 39.700 103.700 40.100 103.800 ;
        RECT 36.600 103.100 37.000 103.500 ;
        RECT 38.300 103.400 40.100 103.700 ;
        RECT 39.400 103.100 39.700 103.400 ;
        RECT 41.400 103.100 41.800 103.500 ;
        RECT 36.600 102.800 37.600 103.100 ;
        RECT 37.200 101.100 37.600 102.800 ;
        RECT 39.400 101.100 39.800 103.100 ;
        RECT 41.500 101.100 42.100 103.100 ;
        RECT 43.800 101.100 44.200 105.400 ;
        RECT 45.600 105.100 45.900 106.100 ;
        RECT 46.400 105.100 46.700 106.800 ;
        RECT 49.700 106.700 50.100 106.800 ;
        RECT 48.900 106.200 49.300 106.300 ;
        RECT 48.900 106.100 51.400 106.200 ;
        RECT 52.600 106.100 53.000 106.200 ;
        RECT 48.900 105.900 53.000 106.100 ;
        RECT 51.000 105.800 53.000 105.900 ;
        RECT 44.600 104.800 45.900 105.100 ;
        RECT 44.600 101.100 45.000 104.800 ;
        RECT 46.200 104.600 46.700 105.100 ;
        RECT 47.800 105.500 50.600 105.600 ;
        RECT 47.800 105.400 50.700 105.500 ;
        RECT 47.800 105.300 52.700 105.400 ;
        RECT 46.200 101.100 46.600 104.600 ;
        RECT 47.800 101.100 48.200 105.300 ;
        RECT 50.300 105.100 52.700 105.300 ;
        RECT 49.400 104.500 52.100 104.800 ;
        RECT 49.400 104.400 49.800 104.500 ;
        RECT 51.700 104.400 52.100 104.500 ;
        RECT 52.400 104.500 52.700 105.100 ;
        RECT 53.400 105.200 53.700 106.800 ;
        RECT 54.200 106.400 54.600 106.500 ;
        RECT 54.200 106.100 56.100 106.400 ;
        RECT 55.700 106.000 56.100 106.100 ;
        RECT 54.900 105.700 55.300 105.800 ;
        RECT 56.600 105.700 57.000 107.400 ;
        RECT 54.900 105.400 57.000 105.700 ;
        RECT 53.400 104.900 54.600 105.200 ;
        RECT 53.100 104.500 53.500 104.600 ;
        RECT 52.400 104.200 53.500 104.500 ;
        RECT 54.300 104.400 54.600 104.900 ;
        RECT 54.300 104.000 55.000 104.400 ;
        RECT 51.100 103.700 51.500 103.800 ;
        RECT 52.500 103.700 52.900 103.800 ;
        RECT 49.400 103.100 49.800 103.500 ;
        RECT 51.100 103.400 52.900 103.700 ;
        RECT 52.200 103.100 52.500 103.400 ;
        RECT 54.200 103.100 54.600 103.500 ;
        RECT 49.400 102.800 50.400 103.100 ;
        RECT 50.000 101.100 50.400 102.800 ;
        RECT 52.200 101.100 52.600 103.100 ;
        RECT 54.300 101.100 54.900 103.100 ;
        RECT 56.600 101.100 57.000 105.400 ;
        RECT 58.200 104.100 58.600 109.900 ;
        RECT 60.300 108.200 60.700 109.900 ;
        RECT 59.800 107.900 60.700 108.200 ;
        RECT 61.400 107.900 61.800 109.900 ;
        RECT 62.200 108.000 62.600 109.900 ;
        RECT 63.800 108.000 64.200 109.900 ;
        RECT 62.200 107.900 64.200 108.000 ;
        RECT 59.000 106.800 59.400 107.600 ;
        RECT 59.800 106.100 60.200 107.900 ;
        RECT 61.500 107.200 61.800 107.900 ;
        RECT 62.300 107.700 64.100 107.900 ;
        RECT 64.600 107.500 65.000 109.900 ;
        RECT 66.800 109.200 67.200 109.900 ;
        RECT 66.200 108.900 67.200 109.200 ;
        RECT 69.000 108.900 69.400 109.900 ;
        RECT 71.100 109.200 71.700 109.900 ;
        RECT 71.000 108.900 71.700 109.200 ;
        RECT 66.200 108.500 66.600 108.900 ;
        RECT 69.000 108.600 69.300 108.900 ;
        RECT 67.000 108.200 67.400 108.600 ;
        RECT 67.900 108.300 69.300 108.600 ;
        RECT 71.000 108.500 71.400 108.900 ;
        RECT 67.900 108.200 68.300 108.300 ;
        RECT 63.400 107.200 63.800 107.400 ;
        RECT 61.400 106.800 62.700 107.200 ;
        RECT 63.400 106.900 64.200 107.200 ;
        RECT 63.800 106.800 64.200 106.900 ;
        RECT 65.000 107.100 65.800 107.200 ;
        RECT 67.100 107.100 67.400 108.200 ;
        RECT 71.900 107.700 72.300 107.800 ;
        RECT 73.400 107.700 73.800 109.900 ;
        RECT 71.900 107.400 73.800 107.700 ;
        RECT 69.900 107.100 70.600 107.200 ;
        RECT 65.000 106.800 70.600 107.100 ;
        RECT 59.800 105.800 61.700 106.100 ;
        RECT 59.000 104.100 59.400 104.200 ;
        RECT 58.200 103.800 59.400 104.100 ;
        RECT 58.200 101.100 58.600 103.800 ;
        RECT 59.800 101.100 60.200 105.800 ;
        RECT 61.400 105.200 61.700 105.800 ;
        RECT 60.600 104.400 61.000 105.200 ;
        RECT 61.400 105.100 61.800 105.200 ;
        RECT 62.400 105.100 62.700 106.800 ;
        RECT 66.500 106.700 66.900 106.800 ;
        RECT 63.000 105.800 63.400 106.600 ;
        RECT 65.700 106.200 66.100 106.300 ;
        RECT 65.700 105.900 68.200 106.200 ;
        RECT 67.800 105.800 68.200 105.900 ;
        RECT 64.600 105.500 67.400 105.600 ;
        RECT 64.600 105.400 67.500 105.500 ;
        RECT 64.600 105.300 69.500 105.400 ;
        RECT 61.400 104.800 62.100 105.100 ;
        RECT 62.400 104.800 62.900 105.100 ;
        RECT 61.800 104.200 62.100 104.800 ;
        RECT 61.800 103.800 62.200 104.200 ;
        RECT 62.500 101.100 62.900 104.800 ;
        RECT 64.600 101.100 65.000 105.300 ;
        RECT 67.100 105.100 69.500 105.300 ;
        RECT 66.200 104.500 68.900 104.800 ;
        RECT 66.200 104.400 66.600 104.500 ;
        RECT 68.500 104.400 68.900 104.500 ;
        RECT 69.200 104.500 69.500 105.100 ;
        RECT 70.200 105.200 70.500 106.800 ;
        RECT 71.000 106.400 71.400 106.500 ;
        RECT 71.000 106.100 72.900 106.400 ;
        RECT 72.500 106.000 72.900 106.100 ;
        RECT 71.700 105.700 72.100 105.800 ;
        RECT 73.400 105.700 73.800 107.400 ;
        RECT 74.200 107.600 74.600 109.900 ;
        RECT 75.800 108.200 76.200 109.900 ;
        RECT 75.800 107.900 76.300 108.200 ;
        RECT 77.400 108.000 77.800 109.900 ;
        RECT 79.000 108.000 79.400 109.900 ;
        RECT 77.400 107.900 79.400 108.000 ;
        RECT 79.800 107.900 80.200 109.900 ;
        RECT 80.600 108.000 81.000 109.900 ;
        RECT 82.200 108.000 82.600 109.900 ;
        RECT 80.600 107.900 82.600 108.000 ;
        RECT 83.000 107.900 83.400 109.900 ;
        RECT 83.800 107.900 84.200 109.900 ;
        RECT 84.600 108.000 85.000 109.900 ;
        RECT 86.200 108.000 86.600 109.900 ;
        RECT 84.600 107.900 86.600 108.000 ;
        RECT 74.200 107.300 75.500 107.600 ;
        RECT 74.300 106.200 74.700 106.600 ;
        RECT 74.200 105.800 74.700 106.200 ;
        RECT 75.200 106.500 75.500 107.300 ;
        RECT 76.000 107.200 76.300 107.900 ;
        RECT 77.500 107.700 79.300 107.900 ;
        RECT 77.800 107.200 78.200 107.400 ;
        RECT 79.800 107.200 80.100 107.900 ;
        RECT 80.700 107.700 82.500 107.900 ;
        RECT 81.000 107.200 81.400 107.400 ;
        RECT 83.000 107.200 83.300 107.900 ;
        RECT 83.900 107.200 84.200 107.900 ;
        RECT 84.700 107.700 86.500 107.900 ;
        RECT 88.600 107.500 89.000 109.900 ;
        RECT 90.800 109.200 91.200 109.900 ;
        RECT 90.200 108.900 91.200 109.200 ;
        RECT 93.000 108.900 93.400 109.900 ;
        RECT 95.100 109.200 95.700 109.900 ;
        RECT 95.000 108.900 95.700 109.200 ;
        RECT 90.200 108.500 90.600 108.900 ;
        RECT 93.000 108.600 93.300 108.900 ;
        RECT 91.000 108.200 91.400 108.600 ;
        RECT 91.900 108.300 93.300 108.600 ;
        RECT 95.000 108.500 95.400 108.900 ;
        RECT 91.900 108.200 92.300 108.300 ;
        RECT 85.800 107.200 86.200 107.400 ;
        RECT 75.800 107.100 76.300 107.200 ;
        RECT 75.800 106.800 76.900 107.100 ;
        RECT 77.400 106.900 78.200 107.200 ;
        RECT 77.400 106.800 77.800 106.900 ;
        RECT 78.900 106.800 80.200 107.200 ;
        RECT 80.600 106.900 81.400 107.200 ;
        RECT 80.600 106.800 81.000 106.900 ;
        RECT 82.100 106.800 83.400 107.200 ;
        RECT 83.800 106.800 85.100 107.200 ;
        RECT 85.800 106.900 86.600 107.200 ;
        RECT 86.200 106.800 86.600 106.900 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 89.000 107.100 89.800 107.200 ;
        RECT 91.100 107.100 91.400 108.200 ;
        RECT 94.200 107.800 94.600 108.200 ;
        RECT 94.200 107.200 94.500 107.800 ;
        RECT 95.900 107.700 96.300 107.800 ;
        RECT 97.400 107.700 97.800 109.900 ;
        RECT 98.200 108.000 98.600 109.900 ;
        RECT 99.800 108.000 100.200 109.900 ;
        RECT 98.200 107.900 100.200 108.000 ;
        RECT 100.600 107.900 101.000 109.900 ;
        RECT 101.700 108.200 102.100 109.900 ;
        RECT 101.700 107.900 102.600 108.200 ;
        RECT 98.300 107.700 100.100 107.900 ;
        RECT 95.900 107.400 97.800 107.700 ;
        RECT 93.900 107.100 94.500 107.200 ;
        RECT 87.800 106.800 94.500 107.100 ;
        RECT 75.200 106.100 75.700 106.500 ;
        RECT 71.700 105.400 73.800 105.700 ;
        RECT 70.200 104.900 71.400 105.200 ;
        RECT 69.900 104.500 70.300 104.600 ;
        RECT 69.200 104.200 70.300 104.500 ;
        RECT 71.100 104.400 71.400 104.900 ;
        RECT 71.100 104.000 71.800 104.400 ;
        RECT 67.900 103.700 68.300 103.800 ;
        RECT 69.300 103.700 69.700 103.800 ;
        RECT 66.200 103.100 66.600 103.500 ;
        RECT 67.900 103.400 69.700 103.700 ;
        RECT 69.000 103.100 69.300 103.400 ;
        RECT 71.000 103.100 71.400 103.500 ;
        RECT 66.200 102.800 67.200 103.100 ;
        RECT 66.800 101.100 67.200 102.800 ;
        RECT 69.000 101.100 69.400 103.100 ;
        RECT 71.100 101.100 71.700 103.100 ;
        RECT 73.400 101.100 73.800 105.400 ;
        RECT 75.200 105.100 75.500 106.100 ;
        RECT 76.000 105.100 76.300 106.800 ;
        RECT 76.600 106.100 76.900 106.800 ;
        RECT 78.200 106.100 78.600 106.600 ;
        RECT 76.600 105.800 78.600 106.100 ;
        RECT 78.900 106.200 79.200 106.800 ;
        RECT 78.900 105.800 79.400 106.200 ;
        RECT 81.400 105.800 81.800 106.600 ;
        RECT 82.100 106.100 82.400 106.800 ;
        RECT 82.100 105.800 84.100 106.100 ;
        RECT 78.900 105.100 79.200 105.800 ;
        RECT 79.800 105.100 80.200 105.200 ;
        RECT 82.100 105.100 82.400 105.800 ;
        RECT 83.800 105.200 84.100 105.800 ;
        RECT 83.000 105.100 83.400 105.200 ;
        RECT 74.200 104.800 75.500 105.100 ;
        RECT 74.200 101.100 74.600 104.800 ;
        RECT 75.800 104.600 76.300 105.100 ;
        RECT 78.700 104.800 79.200 105.100 ;
        RECT 79.500 104.800 80.200 105.100 ;
        RECT 81.900 104.800 82.400 105.100 ;
        RECT 82.700 104.800 83.400 105.100 ;
        RECT 83.800 105.100 84.200 105.200 ;
        RECT 84.800 105.100 85.100 106.800 ;
        RECT 90.500 106.700 90.900 106.800 ;
        RECT 85.400 105.800 85.800 106.600 ;
        RECT 89.700 106.200 90.100 106.300 ;
        RECT 89.700 105.900 92.200 106.200 ;
        RECT 91.800 105.800 92.200 105.900 ;
        RECT 88.600 105.500 91.400 105.600 ;
        RECT 88.600 105.400 91.500 105.500 ;
        RECT 88.600 105.300 93.500 105.400 ;
        RECT 83.800 104.800 84.500 105.100 ;
        RECT 84.800 104.800 85.300 105.100 ;
        RECT 75.800 101.100 76.200 104.600 ;
        RECT 78.700 101.100 79.100 104.800 ;
        RECT 79.500 104.200 79.800 104.800 ;
        RECT 79.400 103.800 80.200 104.200 ;
        RECT 81.900 101.100 82.300 104.800 ;
        RECT 82.700 104.200 83.000 104.800 ;
        RECT 82.600 103.800 83.000 104.200 ;
        RECT 84.200 104.200 84.500 104.800 ;
        RECT 84.200 103.800 84.600 104.200 ;
        RECT 84.900 101.100 85.300 104.800 ;
        RECT 88.600 101.100 89.000 105.300 ;
        RECT 91.100 105.100 93.500 105.300 ;
        RECT 90.200 104.500 92.900 104.800 ;
        RECT 90.200 104.400 90.600 104.500 ;
        RECT 92.500 104.400 92.900 104.500 ;
        RECT 93.200 104.500 93.500 105.100 ;
        RECT 94.200 105.200 94.500 106.800 ;
        RECT 95.000 106.400 95.400 106.500 ;
        RECT 95.000 106.100 96.900 106.400 ;
        RECT 96.500 106.000 96.900 106.100 ;
        RECT 95.700 105.700 96.100 105.800 ;
        RECT 97.400 105.700 97.800 107.400 ;
        RECT 98.600 107.200 99.000 107.400 ;
        RECT 100.600 107.200 100.900 107.900 ;
        RECT 98.200 106.900 99.000 107.200 ;
        RECT 98.200 106.800 98.600 106.900 ;
        RECT 99.700 106.800 101.000 107.200 ;
        RECT 99.000 105.800 99.400 106.600 ;
        RECT 95.700 105.400 97.800 105.700 ;
        RECT 94.200 104.900 95.400 105.200 ;
        RECT 93.900 104.500 94.300 104.600 ;
        RECT 93.200 104.200 94.300 104.500 ;
        RECT 95.100 104.400 95.400 104.900 ;
        RECT 95.100 104.000 95.800 104.400 ;
        RECT 91.900 103.700 92.300 103.800 ;
        RECT 93.300 103.700 93.700 103.800 ;
        RECT 90.200 103.100 90.600 103.500 ;
        RECT 91.900 103.400 93.700 103.700 ;
        RECT 93.000 103.100 93.300 103.400 ;
        RECT 95.000 103.100 95.400 103.500 ;
        RECT 90.200 102.800 91.200 103.100 ;
        RECT 90.800 101.100 91.200 102.800 ;
        RECT 93.000 101.100 93.400 103.100 ;
        RECT 95.100 101.100 95.700 103.100 ;
        RECT 97.400 101.100 97.800 105.400 ;
        RECT 99.700 105.200 100.000 106.800 ;
        RECT 102.200 106.100 102.600 107.900 ;
        RECT 103.000 106.800 103.400 107.600 ;
        RECT 103.800 107.500 104.200 109.900 ;
        RECT 106.000 109.200 106.400 109.900 ;
        RECT 105.400 108.900 106.400 109.200 ;
        RECT 108.200 108.900 108.600 109.900 ;
        RECT 110.300 109.200 110.900 109.900 ;
        RECT 110.200 108.900 110.900 109.200 ;
        RECT 105.400 108.500 105.800 108.900 ;
        RECT 108.200 108.600 108.500 108.900 ;
        RECT 106.200 108.200 106.600 108.600 ;
        RECT 107.100 108.300 108.500 108.600 ;
        RECT 110.200 108.500 110.600 108.900 ;
        RECT 107.100 108.200 107.500 108.300 ;
        RECT 106.300 107.200 106.600 108.200 ;
        RECT 111.100 107.700 111.500 107.800 ;
        RECT 112.600 107.700 113.000 109.900 ;
        RECT 111.100 107.400 113.000 107.700 ;
        RECT 104.200 107.100 105.000 107.200 ;
        RECT 106.200 107.100 106.600 107.200 ;
        RECT 109.100 107.100 109.500 107.200 ;
        RECT 104.200 106.800 109.700 107.100 ;
        RECT 105.700 106.700 106.100 106.800 ;
        RECT 99.000 104.800 100.000 105.200 ;
        RECT 100.600 105.800 102.600 106.100 ;
        RECT 104.900 106.200 105.300 106.300 ;
        RECT 104.900 105.900 107.400 106.200 ;
        RECT 107.000 105.800 107.400 105.900 ;
        RECT 100.600 105.200 100.900 105.800 ;
        RECT 100.600 105.100 101.000 105.200 ;
        RECT 100.300 104.800 101.000 105.100 ;
        RECT 99.500 101.100 99.900 104.800 ;
        RECT 100.300 104.200 100.600 104.800 ;
        RECT 101.400 104.400 101.800 105.200 ;
        RECT 100.200 103.800 100.600 104.200 ;
        RECT 102.200 101.100 102.600 105.800 ;
        RECT 103.800 105.500 106.600 105.600 ;
        RECT 103.800 105.400 106.700 105.500 ;
        RECT 103.800 105.300 108.700 105.400 ;
        RECT 103.800 101.100 104.200 105.300 ;
        RECT 106.300 105.100 108.700 105.300 ;
        RECT 105.400 104.500 108.100 104.800 ;
        RECT 105.400 104.400 105.800 104.500 ;
        RECT 107.700 104.400 108.100 104.500 ;
        RECT 108.400 104.500 108.700 105.100 ;
        RECT 109.400 105.200 109.700 106.800 ;
        RECT 110.200 106.400 110.600 106.500 ;
        RECT 110.200 106.100 112.100 106.400 ;
        RECT 111.700 106.000 112.100 106.100 ;
        RECT 110.900 105.700 111.300 105.800 ;
        RECT 112.600 105.700 113.000 107.400 ;
        RECT 113.400 106.800 113.800 107.600 ;
        RECT 110.900 105.400 113.000 105.700 ;
        RECT 109.400 104.900 110.600 105.200 ;
        RECT 109.100 104.500 109.500 104.600 ;
        RECT 108.400 104.200 109.500 104.500 ;
        RECT 110.300 104.400 110.600 104.900 ;
        RECT 110.300 104.000 111.000 104.400 ;
        RECT 107.100 103.700 107.500 103.800 ;
        RECT 108.500 103.700 108.900 103.800 ;
        RECT 105.400 103.100 105.800 103.500 ;
        RECT 107.100 103.400 108.900 103.700 ;
        RECT 108.200 103.100 108.500 103.400 ;
        RECT 110.200 103.100 110.600 103.500 ;
        RECT 105.400 102.800 106.400 103.100 ;
        RECT 106.000 101.100 106.400 102.800 ;
        RECT 108.200 101.100 108.600 103.100 ;
        RECT 110.300 101.100 110.900 103.100 ;
        RECT 112.600 101.100 113.000 105.400 ;
        RECT 114.200 101.100 114.600 109.900 ;
        RECT 116.600 108.900 117.000 109.900 ;
        RECT 116.600 107.200 116.900 108.900 ;
        RECT 117.400 107.800 117.800 108.600 ;
        RECT 119.000 108.200 119.400 109.900 ;
        RECT 118.900 107.900 119.400 108.200 ;
        RECT 118.900 107.200 119.200 107.900 ;
        RECT 120.600 107.600 121.000 109.900 ;
        RECT 119.700 107.300 121.000 107.600 ;
        RECT 121.400 107.600 121.800 109.900 ;
        RECT 123.000 108.200 123.400 109.900 ;
        RECT 123.000 107.900 123.500 108.200 ;
        RECT 124.600 107.900 125.000 109.900 ;
        RECT 125.400 108.000 125.800 109.900 ;
        RECT 127.000 108.000 127.400 109.900 ;
        RECT 125.400 107.900 127.400 108.000 ;
        RECT 121.400 107.300 122.700 107.600 ;
        RECT 116.600 106.800 117.000 107.200 ;
        RECT 118.900 106.800 119.400 107.200 ;
        RECT 115.800 105.400 116.200 106.200 ;
        RECT 116.600 105.100 116.900 106.800 ;
        RECT 118.900 105.100 119.200 106.800 ;
        RECT 119.700 106.500 120.000 107.300 ;
        RECT 119.500 106.100 120.000 106.500 ;
        RECT 119.700 105.100 120.000 106.100 ;
        RECT 120.500 106.200 120.900 106.600 ;
        RECT 121.500 106.200 121.900 106.600 ;
        RECT 120.500 105.800 121.000 106.200 ;
        RECT 121.400 105.800 121.900 106.200 ;
        RECT 122.400 106.500 122.700 107.300 ;
        RECT 123.200 107.200 123.500 107.900 ;
        RECT 124.700 107.200 125.000 107.900 ;
        RECT 125.500 107.700 127.300 107.900 ;
        RECT 127.800 107.500 128.200 109.900 ;
        RECT 130.000 109.200 130.400 109.900 ;
        RECT 129.400 108.900 130.400 109.200 ;
        RECT 132.200 108.900 132.600 109.900 ;
        RECT 134.300 109.200 134.900 109.900 ;
        RECT 134.200 108.900 134.900 109.200 ;
        RECT 129.400 108.500 129.800 108.900 ;
        RECT 132.200 108.600 132.500 108.900 ;
        RECT 130.200 108.200 130.600 108.600 ;
        RECT 131.100 108.300 132.500 108.600 ;
        RECT 134.200 108.500 134.600 108.900 ;
        RECT 131.100 108.200 131.500 108.300 ;
        RECT 126.600 107.200 127.000 107.400 ;
        RECT 123.000 107.100 123.500 107.200 ;
        RECT 123.800 107.100 124.200 107.200 ;
        RECT 123.000 106.800 124.200 107.100 ;
        RECT 124.600 106.800 125.900 107.200 ;
        RECT 126.600 106.900 127.400 107.200 ;
        RECT 127.000 106.800 127.400 106.900 ;
        RECT 128.200 107.100 129.000 107.200 ;
        RECT 130.300 107.100 130.600 108.200 ;
        RECT 135.100 107.700 135.500 107.800 ;
        RECT 136.600 107.700 137.000 109.900 ;
        RECT 137.400 108.000 137.800 109.900 ;
        RECT 139.000 108.000 139.400 109.900 ;
        RECT 137.400 107.900 139.400 108.000 ;
        RECT 139.800 107.900 140.200 109.900 ;
        RECT 142.500 108.200 142.900 109.900 ;
        RECT 142.500 107.900 143.400 108.200 ;
        RECT 137.500 107.700 139.300 107.900 ;
        RECT 135.100 107.400 137.000 107.700 ;
        RECT 133.100 107.100 133.500 107.200 ;
        RECT 128.200 106.800 133.700 107.100 ;
        RECT 122.400 106.100 122.900 106.500 ;
        RECT 122.400 105.100 122.700 106.100 ;
        RECT 123.200 105.100 123.500 106.800 ;
        RECT 125.600 105.200 125.900 106.800 ;
        RECT 129.700 106.700 130.100 106.800 ;
        RECT 126.200 105.800 126.600 106.600 ;
        RECT 128.900 106.200 129.300 106.300 ;
        RECT 128.900 105.900 131.400 106.200 ;
        RECT 131.000 105.800 131.400 105.900 ;
        RECT 127.800 105.500 130.600 105.600 ;
        RECT 127.800 105.400 130.700 105.500 ;
        RECT 127.800 105.300 132.700 105.400 ;
        RECT 116.100 104.700 117.000 105.100 ;
        RECT 116.100 102.200 116.500 104.700 ;
        RECT 118.900 104.600 119.400 105.100 ;
        RECT 119.700 104.800 121.000 105.100 ;
        RECT 115.800 101.800 116.500 102.200 ;
        RECT 116.100 101.100 116.500 101.800 ;
        RECT 119.000 101.100 119.400 104.600 ;
        RECT 120.600 101.100 121.000 104.800 ;
        RECT 121.400 104.800 122.700 105.100 ;
        RECT 121.400 101.100 121.800 104.800 ;
        RECT 123.000 104.600 123.500 105.100 ;
        RECT 124.600 105.100 125.000 105.200 ;
        RECT 124.600 104.800 125.300 105.100 ;
        RECT 125.600 104.800 126.600 105.200 ;
        RECT 123.000 101.100 123.400 104.600 ;
        RECT 125.000 104.200 125.300 104.800 ;
        RECT 125.000 103.800 125.400 104.200 ;
        RECT 125.700 101.100 126.100 104.800 ;
        RECT 127.800 101.100 128.200 105.300 ;
        RECT 130.300 105.100 132.700 105.300 ;
        RECT 129.400 104.500 132.100 104.800 ;
        RECT 129.400 104.400 129.800 104.500 ;
        RECT 131.700 104.400 132.100 104.500 ;
        RECT 132.400 104.500 132.700 105.100 ;
        RECT 133.400 105.200 133.700 106.800 ;
        RECT 134.200 106.400 134.600 106.500 ;
        RECT 134.200 106.100 136.100 106.400 ;
        RECT 135.700 106.000 136.100 106.100 ;
        RECT 134.900 105.700 135.300 105.800 ;
        RECT 136.600 105.700 137.000 107.400 ;
        RECT 137.800 107.200 138.200 107.400 ;
        RECT 139.800 107.200 140.100 107.900 ;
        RECT 137.400 106.900 138.200 107.200 ;
        RECT 137.400 106.800 137.800 106.900 ;
        RECT 138.900 106.800 140.200 107.200 ;
        RECT 137.400 106.100 137.800 106.200 ;
        RECT 138.200 106.100 138.600 106.600 ;
        RECT 137.400 105.800 138.600 106.100 ;
        RECT 134.900 105.400 137.000 105.700 ;
        RECT 133.400 104.900 134.600 105.200 ;
        RECT 133.100 104.500 133.500 104.600 ;
        RECT 132.400 104.200 133.500 104.500 ;
        RECT 134.300 104.400 134.600 104.900 ;
        RECT 134.300 104.000 135.000 104.400 ;
        RECT 131.100 103.700 131.500 103.800 ;
        RECT 132.500 103.700 132.900 103.800 ;
        RECT 129.400 103.100 129.800 103.500 ;
        RECT 131.100 103.400 132.900 103.700 ;
        RECT 132.200 103.100 132.500 103.400 ;
        RECT 134.200 103.100 134.600 103.500 ;
        RECT 129.400 102.800 130.400 103.100 ;
        RECT 130.000 101.100 130.400 102.800 ;
        RECT 132.200 101.100 132.600 103.100 ;
        RECT 134.300 101.100 134.900 103.100 ;
        RECT 136.600 101.100 137.000 105.400 ;
        RECT 138.900 105.100 139.200 106.800 ;
        RECT 143.000 106.100 143.400 107.900 ;
        RECT 144.600 107.800 145.000 108.600 ;
        RECT 143.800 107.100 144.200 107.600 ;
        RECT 144.600 107.100 144.900 107.800 ;
        RECT 143.800 106.800 144.900 107.100 ;
        RECT 140.600 105.800 143.400 106.100 ;
        RECT 139.800 105.100 140.200 105.200 ;
        RECT 140.600 105.100 140.900 105.800 ;
        RECT 138.700 104.800 139.200 105.100 ;
        RECT 139.500 104.800 140.900 105.100 ;
        RECT 138.700 101.100 139.100 104.800 ;
        RECT 139.500 104.200 139.800 104.800 ;
        RECT 142.200 104.400 142.600 105.200 ;
        RECT 139.400 103.800 139.800 104.200 ;
        RECT 143.000 101.100 143.400 105.800 ;
        RECT 145.400 106.100 145.800 109.900 ;
        RECT 146.200 107.900 146.600 109.900 ;
        RECT 147.000 108.000 147.400 109.900 ;
        RECT 148.600 108.000 149.000 109.900 ;
        RECT 147.000 107.900 149.000 108.000 ;
        RECT 149.400 108.000 149.800 109.900 ;
        RECT 151.000 108.000 151.400 109.900 ;
        RECT 149.400 107.900 151.400 108.000 ;
        RECT 151.800 107.900 152.200 109.900 ;
        RECT 153.900 108.200 154.300 109.900 ;
        RECT 155.800 108.900 156.200 109.900 ;
        RECT 153.400 108.100 154.300 108.200 ;
        RECT 155.000 108.100 155.400 108.200 ;
        RECT 146.300 107.200 146.600 107.900 ;
        RECT 147.100 107.700 148.900 107.900 ;
        RECT 149.500 107.700 151.300 107.900 ;
        RECT 148.200 107.200 148.600 107.400 ;
        RECT 149.800 107.200 150.200 107.400 ;
        RECT 151.800 107.200 152.100 107.900 ;
        RECT 153.400 107.800 155.400 108.100 ;
        RECT 146.200 106.800 147.500 107.200 ;
        RECT 148.200 106.900 149.000 107.200 ;
        RECT 148.600 106.800 149.000 106.900 ;
        RECT 149.400 106.900 150.200 107.200 ;
        RECT 150.900 107.100 152.200 107.200 ;
        RECT 152.600 107.100 153.000 107.600 ;
        RECT 149.400 106.800 149.800 106.900 ;
        RECT 150.900 106.800 153.000 107.100 ;
        RECT 146.200 106.100 146.600 106.200 ;
        RECT 145.400 105.800 146.600 106.100 ;
        RECT 145.400 101.100 145.800 105.800 ;
        RECT 147.200 105.200 147.500 106.800 ;
        RECT 147.800 105.800 148.200 106.600 ;
        RECT 148.600 106.100 149.000 106.200 ;
        RECT 150.200 106.100 150.600 106.600 ;
        RECT 148.600 105.800 150.600 106.100 ;
        RECT 146.200 105.100 146.600 105.200 ;
        RECT 146.200 104.800 146.900 105.100 ;
        RECT 147.200 104.800 148.200 105.200 ;
        RECT 150.900 105.100 151.200 106.800 ;
        RECT 151.800 105.100 152.200 105.200 ;
        RECT 150.700 104.800 151.200 105.100 ;
        RECT 151.500 104.800 152.200 105.100 ;
        RECT 146.600 104.200 146.900 104.800 ;
        RECT 146.600 103.800 147.000 104.200 ;
        RECT 147.300 101.100 147.700 104.800 ;
        RECT 150.700 101.100 151.100 104.800 ;
        RECT 151.500 104.200 151.800 104.800 ;
        RECT 151.400 103.800 151.800 104.200 ;
        RECT 153.400 101.100 153.800 107.800 ;
        RECT 155.800 107.200 156.100 108.900 ;
        RECT 156.600 107.800 157.000 108.600 ;
        RECT 157.400 107.900 157.800 109.900 ;
        RECT 158.200 108.000 158.600 109.900 ;
        RECT 159.800 108.000 160.200 109.900 ;
        RECT 158.200 107.900 160.200 108.000 ;
        RECT 162.200 107.900 162.600 109.900 ;
        RECT 162.900 108.200 163.300 108.600 ;
        RECT 157.500 107.200 157.800 107.900 ;
        RECT 158.300 107.700 160.100 107.900 ;
        RECT 159.400 107.200 159.800 107.400 ;
        RECT 155.800 106.800 156.200 107.200 ;
        RECT 157.400 106.800 158.700 107.200 ;
        RECT 159.400 106.900 160.200 107.200 ;
        RECT 159.800 106.800 160.200 106.900 ;
        RECT 160.600 107.100 161.000 107.200 ;
        RECT 161.400 107.100 161.800 107.200 ;
        RECT 160.600 106.800 161.800 107.100 ;
        RECT 155.000 105.400 155.400 106.200 ;
        RECT 155.800 106.100 156.100 106.800 ;
        RECT 156.600 106.100 157.000 106.200 ;
        RECT 155.800 105.800 157.000 106.100 ;
        RECT 154.200 104.400 154.600 105.200 ;
        RECT 155.800 105.100 156.100 105.800 ;
        RECT 158.400 105.200 158.700 106.800 ;
        RECT 159.000 105.800 159.400 106.600 ;
        RECT 161.400 106.400 161.800 106.800 ;
        RECT 159.800 106.100 160.200 106.200 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 162.200 106.100 162.500 107.900 ;
        RECT 163.000 107.800 163.400 108.200 ;
        RECT 163.800 107.900 164.200 109.900 ;
        RECT 164.600 108.000 165.000 109.900 ;
        RECT 166.200 108.000 166.600 109.900 ;
        RECT 164.600 107.900 166.600 108.000 ;
        RECT 163.900 107.200 164.200 107.900 ;
        RECT 164.700 107.700 166.500 107.900 ;
        RECT 165.800 107.200 166.200 107.400 ;
        RECT 163.800 106.800 165.100 107.200 ;
        RECT 165.800 106.900 166.600 107.200 ;
        RECT 166.200 106.800 166.600 106.900 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 163.800 106.100 164.200 106.200 ;
        RECT 159.800 105.800 161.400 106.100 ;
        RECT 162.200 105.800 164.200 106.100 ;
        RECT 161.000 105.600 161.400 105.800 ;
        RECT 157.400 105.100 157.800 105.200 ;
        RECT 155.300 104.700 156.200 105.100 ;
        RECT 157.400 104.800 158.100 105.100 ;
        RECT 158.400 104.800 159.400 105.200 ;
        RECT 163.000 105.100 163.300 105.800 ;
        RECT 163.800 105.100 164.200 105.200 ;
        RECT 164.800 105.100 165.100 106.800 ;
        RECT 165.400 105.800 165.800 106.600 ;
        RECT 160.600 104.800 162.600 105.100 ;
        RECT 155.300 101.100 155.700 104.700 ;
        RECT 157.800 104.200 158.100 104.800 ;
        RECT 157.800 103.800 158.200 104.200 ;
        RECT 158.500 101.100 158.900 104.800 ;
        RECT 160.600 101.100 161.000 104.800 ;
        RECT 162.200 101.100 162.600 104.800 ;
        RECT 163.000 101.100 163.400 105.100 ;
        RECT 163.800 104.800 164.500 105.100 ;
        RECT 164.800 104.800 165.300 105.100 ;
        RECT 164.200 104.200 164.500 104.800 ;
        RECT 164.200 103.800 164.600 104.200 ;
        RECT 164.900 102.200 165.300 104.800 ;
        RECT 164.900 101.800 165.800 102.200 ;
        RECT 164.900 101.100 165.300 101.800 ;
        RECT 167.000 101.100 167.400 109.900 ;
        RECT 167.800 107.800 168.200 108.600 ;
        RECT 168.600 107.700 169.000 109.900 ;
        RECT 170.700 109.200 171.300 109.900 ;
        RECT 170.700 108.900 171.400 109.200 ;
        RECT 173.000 108.900 173.400 109.900 ;
        RECT 175.200 109.200 175.600 109.900 ;
        RECT 175.200 108.900 176.200 109.200 ;
        RECT 171.000 108.500 171.400 108.900 ;
        RECT 173.100 108.600 173.400 108.900 ;
        RECT 173.100 108.300 174.500 108.600 ;
        RECT 174.100 108.200 174.500 108.300 ;
        RECT 175.000 108.200 175.400 108.600 ;
        RECT 175.800 108.500 176.200 108.900 ;
        RECT 170.100 107.700 170.500 107.800 ;
        RECT 168.600 107.400 170.500 107.700 ;
        RECT 168.600 105.700 169.000 107.400 ;
        RECT 175.000 107.200 175.300 108.200 ;
        RECT 177.400 107.500 177.800 109.900 ;
        RECT 179.500 108.200 179.900 109.900 ;
        RECT 179.000 107.900 179.900 108.200 ;
        RECT 180.600 107.900 181.000 109.900 ;
        RECT 181.400 108.000 181.800 109.900 ;
        RECT 183.000 108.000 183.400 109.900 ;
        RECT 185.100 109.200 185.500 109.900 ;
        RECT 184.600 108.800 185.500 109.200 ;
        RECT 185.100 108.200 185.500 108.800 ;
        RECT 181.400 107.900 183.400 108.000 ;
        RECT 184.600 107.900 185.500 108.200 ;
        RECT 186.200 108.000 186.600 109.900 ;
        RECT 187.800 108.000 188.200 109.900 ;
        RECT 186.200 107.900 188.200 108.000 ;
        RECT 188.600 107.900 189.000 109.900 ;
        RECT 189.700 108.200 190.100 109.900 ;
        RECT 189.700 107.900 190.600 108.200 ;
        RECT 172.100 107.100 172.500 107.200 ;
        RECT 175.000 107.100 175.400 107.200 ;
        RECT 176.600 107.100 177.400 107.200 ;
        RECT 171.900 106.800 177.400 107.100 ;
        RECT 178.200 106.800 178.600 107.600 ;
        RECT 171.000 106.400 171.400 106.500 ;
        RECT 169.500 106.100 171.400 106.400 ;
        RECT 169.500 106.000 169.900 106.100 ;
        RECT 170.300 105.700 170.700 105.800 ;
        RECT 168.600 105.400 170.700 105.700 ;
        RECT 167.800 104.100 168.200 104.200 ;
        RECT 168.600 104.100 169.000 105.400 ;
        RECT 171.900 105.200 172.200 106.800 ;
        RECT 175.500 106.700 175.900 106.800 ;
        RECT 176.300 106.200 176.700 106.300 ;
        RECT 174.200 105.900 176.700 106.200 ;
        RECT 178.200 106.200 178.500 106.800 ;
        RECT 174.200 105.800 174.600 105.900 ;
        RECT 178.200 105.800 178.600 106.200 ;
        RECT 179.000 106.100 179.400 107.900 ;
        RECT 180.700 107.200 181.000 107.900 ;
        RECT 181.500 107.700 183.300 107.900 ;
        RECT 182.600 107.200 183.000 107.400 ;
        RECT 180.600 106.800 181.900 107.200 ;
        RECT 182.600 106.900 183.400 107.200 ;
        RECT 183.000 106.800 183.400 106.900 ;
        RECT 183.800 106.800 184.200 107.600 ;
        RECT 179.000 105.800 180.900 106.100 ;
        RECT 175.000 105.500 177.800 105.600 ;
        RECT 174.900 105.400 177.800 105.500 ;
        RECT 171.000 104.900 172.200 105.200 ;
        RECT 172.900 105.300 177.800 105.400 ;
        RECT 172.900 105.100 175.300 105.300 ;
        RECT 171.000 104.400 171.300 104.900 ;
        RECT 167.800 103.800 169.000 104.100 ;
        RECT 170.600 104.000 171.300 104.400 ;
        RECT 172.100 104.500 172.500 104.600 ;
        RECT 172.900 104.500 173.200 105.100 ;
        RECT 172.100 104.200 173.200 104.500 ;
        RECT 173.500 104.500 176.200 104.800 ;
        RECT 173.500 104.400 173.900 104.500 ;
        RECT 175.800 104.400 176.200 104.500 ;
        RECT 168.600 101.100 169.000 103.800 ;
        RECT 172.700 103.700 173.100 103.800 ;
        RECT 174.100 103.700 174.500 103.800 ;
        RECT 171.000 103.100 171.400 103.500 ;
        RECT 172.700 103.400 174.500 103.700 ;
        RECT 173.100 103.100 173.400 103.400 ;
        RECT 175.800 103.100 176.200 103.500 ;
        RECT 170.700 101.100 171.300 103.100 ;
        RECT 173.000 101.100 173.400 103.100 ;
        RECT 175.200 102.800 176.200 103.100 ;
        RECT 175.200 101.100 175.600 102.800 ;
        RECT 177.400 101.100 177.800 105.300 ;
        RECT 179.000 101.100 179.400 105.800 ;
        RECT 180.600 105.200 180.900 105.800 ;
        RECT 179.800 104.400 180.200 105.200 ;
        RECT 180.600 105.100 181.000 105.200 ;
        RECT 181.600 105.100 181.900 106.800 ;
        RECT 182.200 105.800 182.600 106.600 ;
        RECT 180.600 104.800 181.300 105.100 ;
        RECT 181.600 104.800 182.100 105.100 ;
        RECT 181.000 104.200 181.300 104.800 ;
        RECT 181.000 103.800 181.400 104.200 ;
        RECT 181.700 101.100 182.100 104.800 ;
        RECT 184.600 101.100 185.000 107.900 ;
        RECT 186.300 107.700 188.100 107.900 ;
        RECT 186.600 107.200 187.000 107.400 ;
        RECT 188.600 107.200 188.900 107.900 ;
        RECT 186.200 106.900 187.000 107.200 ;
        RECT 186.200 106.800 186.600 106.900 ;
        RECT 187.700 106.800 189.000 107.200 ;
        RECT 187.000 105.800 187.400 106.600 ;
        RECT 185.400 104.400 185.800 105.200 ;
        RECT 187.700 105.100 188.000 106.800 ;
        RECT 190.200 106.100 190.600 107.900 ;
        RECT 193.400 107.700 193.800 109.900 ;
        RECT 195.500 109.200 196.100 109.900 ;
        RECT 195.500 108.900 196.200 109.200 ;
        RECT 197.800 108.900 198.200 109.900 ;
        RECT 200.000 109.200 200.400 109.900 ;
        RECT 200.000 108.900 201.000 109.200 ;
        RECT 195.800 108.500 196.200 108.900 ;
        RECT 197.900 108.600 198.200 108.900 ;
        RECT 197.900 108.300 199.300 108.600 ;
        RECT 198.900 108.200 199.300 108.300 ;
        RECT 199.800 108.200 200.200 108.600 ;
        RECT 200.600 108.500 201.000 108.900 ;
        RECT 194.900 107.700 195.300 107.800 ;
        RECT 191.000 107.100 191.400 107.600 ;
        RECT 193.400 107.400 195.300 107.700 ;
        RECT 193.400 107.100 193.800 107.400 ;
        RECT 196.900 107.100 197.300 107.200 ;
        RECT 199.800 107.100 200.100 108.200 ;
        RECT 202.200 107.500 202.600 109.900 ;
        RECT 203.800 107.600 204.200 109.900 ;
        RECT 205.400 107.600 205.800 109.900 ;
        RECT 207.000 108.000 207.400 109.900 ;
        RECT 208.600 108.000 209.000 109.900 ;
        RECT 207.000 107.900 209.000 108.000 ;
        RECT 209.400 107.900 209.800 109.900 ;
        RECT 207.100 107.700 208.900 107.900 ;
        RECT 203.800 107.200 205.800 107.600 ;
        RECT 207.400 107.200 207.800 107.400 ;
        RECT 209.400 107.200 209.700 107.900 ;
        RECT 210.200 107.700 210.600 109.900 ;
        RECT 212.300 109.200 212.900 109.900 ;
        RECT 212.300 108.900 213.000 109.200 ;
        RECT 214.600 108.900 215.000 109.900 ;
        RECT 216.800 109.200 217.200 109.900 ;
        RECT 216.800 108.900 217.800 109.200 ;
        RECT 212.600 108.500 213.000 108.900 ;
        RECT 214.700 108.600 215.000 108.900 ;
        RECT 214.700 108.300 216.100 108.600 ;
        RECT 215.700 108.200 216.100 108.300 ;
        RECT 216.600 107.800 217.000 108.600 ;
        RECT 217.400 108.500 217.800 108.900 ;
        RECT 211.700 107.700 212.100 107.800 ;
        RECT 210.200 107.400 212.100 107.700 ;
        RECT 201.400 107.100 202.200 107.200 ;
        RECT 191.000 106.800 193.800 107.100 ;
        RECT 188.600 105.800 190.600 106.100 ;
        RECT 188.600 105.200 188.900 105.800 ;
        RECT 188.600 105.100 189.000 105.200 ;
        RECT 187.500 104.800 188.000 105.100 ;
        RECT 188.300 104.800 189.000 105.100 ;
        RECT 187.500 101.100 187.900 104.800 ;
        RECT 188.300 104.200 188.600 104.800 ;
        RECT 189.400 104.400 189.800 105.200 ;
        RECT 188.200 103.800 188.600 104.200 ;
        RECT 190.200 101.100 190.600 105.800 ;
        RECT 193.400 105.700 193.800 106.800 ;
        RECT 196.700 106.800 202.200 107.100 ;
        RECT 195.800 106.400 196.200 106.500 ;
        RECT 194.300 106.100 196.200 106.400 ;
        RECT 194.300 106.000 194.700 106.100 ;
        RECT 195.100 105.700 195.500 105.800 ;
        RECT 193.400 105.400 195.500 105.700 ;
        RECT 191.800 102.100 192.200 102.200 ;
        RECT 193.400 102.100 193.800 105.400 ;
        RECT 196.700 105.200 197.000 106.800 ;
        RECT 200.300 106.700 200.700 106.800 ;
        RECT 201.100 106.200 201.500 106.300 ;
        RECT 197.400 106.100 197.800 106.200 ;
        RECT 199.000 106.100 201.500 106.200 ;
        RECT 197.400 105.900 201.500 106.100 ;
        RECT 197.400 105.800 199.400 105.900 ;
        RECT 204.600 105.800 205.000 106.200 ;
        RECT 205.400 105.800 205.800 107.200 ;
        RECT 207.000 106.900 207.800 107.200 ;
        RECT 207.000 106.800 207.400 106.900 ;
        RECT 208.500 106.800 209.800 107.200 ;
        RECT 207.800 105.800 208.200 106.600 ;
        RECT 208.500 106.100 208.800 106.800 ;
        RECT 209.400 106.100 209.800 106.200 ;
        RECT 208.500 105.800 209.800 106.100 ;
        RECT 199.800 105.500 202.600 105.600 ;
        RECT 199.700 105.400 202.600 105.500 ;
        RECT 195.800 104.900 197.000 105.200 ;
        RECT 197.700 105.300 202.600 105.400 ;
        RECT 197.700 105.100 200.100 105.300 ;
        RECT 195.800 104.400 196.100 104.900 ;
        RECT 195.400 104.000 196.100 104.400 ;
        RECT 196.900 104.500 197.300 104.600 ;
        RECT 197.700 104.500 198.000 105.100 ;
        RECT 196.900 104.200 198.000 104.500 ;
        RECT 198.300 104.500 201.000 104.800 ;
        RECT 198.300 104.400 198.700 104.500 ;
        RECT 200.600 104.400 201.000 104.500 ;
        RECT 197.500 103.700 197.900 103.800 ;
        RECT 198.900 103.700 199.300 103.800 ;
        RECT 195.800 103.100 196.200 103.500 ;
        RECT 197.500 103.400 199.300 103.700 ;
        RECT 197.900 103.100 198.200 103.400 ;
        RECT 200.600 103.100 201.000 103.500 ;
        RECT 191.800 101.800 193.800 102.100 ;
        RECT 193.400 101.100 193.800 101.800 ;
        RECT 195.500 101.100 196.100 103.100 ;
        RECT 197.800 101.100 198.200 103.100 ;
        RECT 200.000 102.800 201.000 103.100 ;
        RECT 200.000 101.100 200.400 102.800 ;
        RECT 202.200 101.100 202.600 105.300 ;
        RECT 203.800 105.400 205.800 105.800 ;
        RECT 203.800 101.100 204.200 105.400 ;
        RECT 205.400 101.100 205.800 105.400 ;
        RECT 208.500 105.100 208.800 105.800 ;
        RECT 210.200 105.700 210.600 107.400 ;
        RECT 213.700 107.100 214.100 107.200 ;
        RECT 216.600 107.100 216.900 107.800 ;
        RECT 219.000 107.500 219.400 109.900 ;
        RECT 219.800 107.500 220.200 109.900 ;
        RECT 222.000 109.200 222.400 109.900 ;
        RECT 221.400 108.900 222.400 109.200 ;
        RECT 224.200 108.900 224.600 109.900 ;
        RECT 226.300 109.200 226.900 109.900 ;
        RECT 226.200 108.900 226.900 109.200 ;
        RECT 221.400 108.500 221.800 108.900 ;
        RECT 224.200 108.600 224.500 108.900 ;
        RECT 222.200 108.200 222.600 108.600 ;
        RECT 223.100 108.300 224.500 108.600 ;
        RECT 226.200 108.500 226.600 108.900 ;
        RECT 223.100 108.200 223.500 108.300 ;
        RECT 218.200 107.100 219.000 107.200 ;
        RECT 220.200 107.100 221.000 107.200 ;
        RECT 222.300 107.100 222.600 108.200 ;
        RECT 227.100 107.700 227.500 107.800 ;
        RECT 228.600 107.700 229.000 109.900 ;
        RECT 227.100 107.400 229.000 107.700 ;
        RECT 225.100 107.100 225.500 107.200 ;
        RECT 213.500 106.800 225.700 107.100 ;
        RECT 212.600 106.400 213.000 106.500 ;
        RECT 211.100 106.100 213.000 106.400 ;
        RECT 211.100 106.000 211.500 106.100 ;
        RECT 211.900 105.700 212.300 105.800 ;
        RECT 210.200 105.400 212.300 105.700 ;
        RECT 209.400 105.100 209.800 105.200 ;
        RECT 208.300 104.800 208.800 105.100 ;
        RECT 209.100 104.800 209.800 105.100 ;
        RECT 208.300 101.100 208.700 104.800 ;
        RECT 209.100 104.200 209.400 104.800 ;
        RECT 209.000 103.800 209.400 104.200 ;
        RECT 210.200 101.100 210.600 105.400 ;
        RECT 213.500 105.200 213.800 106.800 ;
        RECT 217.100 106.700 217.500 106.800 ;
        RECT 221.700 106.700 222.100 106.800 ;
        RECT 217.900 106.200 218.300 106.300 ;
        RECT 215.000 106.100 215.400 106.200 ;
        RECT 215.800 106.100 218.300 106.200 ;
        RECT 215.000 105.900 218.300 106.100 ;
        RECT 220.900 106.200 221.300 106.300 ;
        RECT 220.900 105.900 223.400 106.200 ;
        RECT 215.000 105.800 216.200 105.900 ;
        RECT 223.000 105.800 223.400 105.900 ;
        RECT 216.600 105.500 219.400 105.600 ;
        RECT 216.500 105.400 219.400 105.500 ;
        RECT 212.600 104.900 213.800 105.200 ;
        RECT 214.500 105.300 219.400 105.400 ;
        RECT 214.500 105.100 216.900 105.300 ;
        RECT 212.600 104.400 212.900 104.900 ;
        RECT 212.200 104.000 212.900 104.400 ;
        RECT 213.700 104.500 214.100 104.600 ;
        RECT 214.500 104.500 214.800 105.100 ;
        RECT 213.700 104.200 214.800 104.500 ;
        RECT 215.100 104.500 217.800 104.800 ;
        RECT 215.100 104.400 215.500 104.500 ;
        RECT 217.400 104.400 217.800 104.500 ;
        RECT 214.300 103.700 214.700 103.800 ;
        RECT 215.700 103.700 216.100 103.800 ;
        RECT 212.600 103.100 213.000 103.500 ;
        RECT 214.300 103.400 216.100 103.700 ;
        RECT 214.700 103.100 215.000 103.400 ;
        RECT 217.400 103.100 217.800 103.500 ;
        RECT 212.300 101.100 212.900 103.100 ;
        RECT 214.600 101.100 215.000 103.100 ;
        RECT 216.800 102.800 217.800 103.100 ;
        RECT 216.800 101.100 217.200 102.800 ;
        RECT 219.000 101.100 219.400 105.300 ;
        RECT 219.800 105.500 222.600 105.600 ;
        RECT 219.800 105.400 222.700 105.500 ;
        RECT 219.800 105.300 224.700 105.400 ;
        RECT 219.800 101.100 220.200 105.300 ;
        RECT 222.300 105.100 224.700 105.300 ;
        RECT 221.400 104.500 224.100 104.800 ;
        RECT 221.400 104.400 221.800 104.500 ;
        RECT 223.700 104.400 224.100 104.500 ;
        RECT 224.400 104.500 224.700 105.100 ;
        RECT 225.400 105.200 225.700 106.800 ;
        RECT 226.200 106.400 226.600 106.500 ;
        RECT 226.200 106.100 228.100 106.400 ;
        RECT 227.700 106.000 228.100 106.100 ;
        RECT 226.900 105.700 227.300 105.800 ;
        RECT 228.600 105.700 229.000 107.400 ;
        RECT 226.900 105.400 229.000 105.700 ;
        RECT 225.400 104.900 226.600 105.200 ;
        RECT 225.100 104.500 225.500 104.600 ;
        RECT 224.400 104.200 225.500 104.500 ;
        RECT 226.300 104.400 226.600 104.900 ;
        RECT 226.300 104.000 227.000 104.400 ;
        RECT 223.100 103.700 223.500 103.800 ;
        RECT 224.500 103.700 224.900 103.800 ;
        RECT 221.400 103.100 221.800 103.500 ;
        RECT 223.100 103.400 224.900 103.700 ;
        RECT 224.200 103.100 224.500 103.400 ;
        RECT 226.200 103.100 226.600 103.500 ;
        RECT 221.400 102.800 222.400 103.100 ;
        RECT 222.000 101.100 222.400 102.800 ;
        RECT 224.200 101.100 224.600 103.100 ;
        RECT 226.300 101.100 226.900 103.100 ;
        RECT 228.600 101.100 229.000 105.400 ;
        RECT 0.600 95.600 1.000 99.900 ;
        RECT 2.700 97.900 3.300 99.900 ;
        RECT 5.000 97.900 5.400 99.900 ;
        RECT 7.200 98.200 7.600 99.900 ;
        RECT 7.200 97.900 8.200 98.200 ;
        RECT 3.000 97.500 3.400 97.900 ;
        RECT 5.100 97.600 5.400 97.900 ;
        RECT 4.700 97.300 6.500 97.600 ;
        RECT 7.800 97.500 8.200 97.900 ;
        RECT 4.700 97.200 5.100 97.300 ;
        RECT 6.100 97.200 6.500 97.300 ;
        RECT 2.600 96.600 3.300 97.000 ;
        RECT 3.000 96.100 3.300 96.600 ;
        RECT 4.100 96.500 5.200 96.800 ;
        RECT 4.100 96.400 4.500 96.500 ;
        RECT 3.000 95.800 4.200 96.100 ;
        RECT 0.600 95.300 2.700 95.600 ;
        RECT 0.600 93.600 1.000 95.300 ;
        RECT 2.300 95.200 2.700 95.300 ;
        RECT 1.500 94.900 1.900 95.000 ;
        RECT 1.500 94.600 3.400 94.900 ;
        RECT 3.000 94.500 3.400 94.600 ;
        RECT 3.900 94.200 4.200 95.800 ;
        RECT 4.900 95.900 5.200 96.500 ;
        RECT 5.500 96.500 5.900 96.600 ;
        RECT 7.800 96.500 8.200 96.600 ;
        RECT 5.500 96.200 8.200 96.500 ;
        RECT 4.900 95.700 7.300 95.900 ;
        RECT 9.400 95.700 9.800 99.900 ;
        RECT 4.900 95.600 9.800 95.700 ;
        RECT 6.900 95.500 9.800 95.600 ;
        RECT 7.000 95.400 9.800 95.500 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 11.000 95.100 11.400 99.900 ;
        RECT 13.000 96.800 13.400 97.200 ;
        RECT 11.800 95.800 12.200 96.600 ;
        RECT 13.000 96.200 13.300 96.800 ;
        RECT 13.700 96.200 14.100 99.900 ;
        RECT 12.600 95.900 13.300 96.200 ;
        RECT 13.600 95.900 14.100 96.200 ;
        RECT 17.100 96.200 17.500 99.900 ;
        RECT 17.800 96.800 18.200 97.200 ;
        RECT 17.900 96.200 18.200 96.800 ;
        RECT 17.100 95.900 17.600 96.200 ;
        RECT 17.900 95.900 18.600 96.200 ;
        RECT 12.600 95.800 13.000 95.900 ;
        RECT 12.600 95.100 12.900 95.800 ;
        RECT 13.600 95.200 13.900 95.900 ;
        RECT 6.200 94.800 8.700 95.100 ;
        RECT 7.000 94.700 7.400 94.800 ;
        RECT 8.300 94.700 8.700 94.800 ;
        RECT 11.000 94.800 12.900 95.100 ;
        RECT 13.400 94.800 13.900 95.200 ;
        RECT 7.500 94.200 7.900 94.300 ;
        RECT 3.900 93.900 9.400 94.200 ;
        RECT 4.100 93.800 5.000 93.900 ;
        RECT 0.600 93.300 2.500 93.600 ;
        RECT 0.600 91.100 1.000 93.300 ;
        RECT 2.100 93.200 2.500 93.300 ;
        RECT 7.000 92.800 7.300 93.900 ;
        RECT 8.600 93.800 9.400 93.900 ;
        RECT 6.100 92.700 6.500 92.800 ;
        RECT 3.000 92.100 3.400 92.500 ;
        RECT 5.100 92.400 6.500 92.700 ;
        RECT 7.000 92.400 7.400 92.800 ;
        RECT 5.100 92.100 5.400 92.400 ;
        RECT 7.800 92.100 8.200 92.500 ;
        RECT 2.700 91.800 3.400 92.100 ;
        RECT 2.700 91.100 3.300 91.800 ;
        RECT 5.000 91.100 5.400 92.100 ;
        RECT 7.200 91.800 8.200 92.100 ;
        RECT 7.200 91.100 7.600 91.800 ;
        RECT 9.400 91.100 9.800 93.500 ;
        RECT 10.200 93.400 10.600 94.200 ;
        RECT 11.000 93.100 11.400 94.800 ;
        RECT 13.600 94.200 13.900 94.800 ;
        RECT 14.200 94.400 14.600 95.200 ;
        RECT 16.600 94.400 17.000 95.200 ;
        RECT 17.300 94.200 17.600 95.900 ;
        RECT 18.200 95.800 18.600 95.900 ;
        RECT 19.000 95.800 19.400 96.600 ;
        RECT 18.200 95.100 18.500 95.800 ;
        RECT 19.800 95.100 20.200 99.900 ;
        RECT 21.400 95.700 21.800 99.900 ;
        RECT 23.600 98.200 24.000 99.900 ;
        RECT 23.000 97.900 24.000 98.200 ;
        RECT 25.800 97.900 26.200 99.900 ;
        RECT 27.900 97.900 28.500 99.900 ;
        RECT 23.000 97.500 23.400 97.900 ;
        RECT 25.800 97.600 26.100 97.900 ;
        RECT 24.700 97.300 26.500 97.600 ;
        RECT 27.800 97.500 28.200 97.900 ;
        RECT 24.700 97.200 25.100 97.300 ;
        RECT 26.100 97.200 26.500 97.300 ;
        RECT 23.000 96.500 23.400 96.600 ;
        RECT 25.300 96.500 25.700 96.600 ;
        RECT 23.000 96.200 25.700 96.500 ;
        RECT 26.000 96.500 27.100 96.800 ;
        RECT 26.000 95.900 26.300 96.500 ;
        RECT 26.700 96.400 27.100 96.500 ;
        RECT 27.900 96.600 28.600 97.000 ;
        RECT 27.900 96.100 28.200 96.600 ;
        RECT 23.900 95.700 26.300 95.900 ;
        RECT 21.400 95.600 26.300 95.700 ;
        RECT 27.000 95.800 28.200 96.100 ;
        RECT 21.400 95.500 24.300 95.600 ;
        RECT 21.400 95.400 24.200 95.500 ;
        RECT 24.600 95.100 25.000 95.200 ;
        RECT 18.200 94.800 20.200 95.100 ;
        RECT 12.600 93.800 13.900 94.200 ;
        RECT 15.000 94.100 15.400 94.200 ;
        RECT 14.600 93.800 15.400 94.100 ;
        RECT 15.800 94.100 16.200 94.200 ;
        RECT 17.300 94.100 18.600 94.200 ;
        RECT 19.000 94.100 19.400 94.200 ;
        RECT 15.800 93.800 16.600 94.100 ;
        RECT 17.300 93.800 19.400 94.100 ;
        RECT 12.700 93.100 13.000 93.800 ;
        RECT 14.600 93.600 15.000 93.800 ;
        RECT 16.200 93.600 16.600 93.800 ;
        RECT 13.500 93.100 15.300 93.300 ;
        RECT 15.900 93.100 17.700 93.300 ;
        RECT 18.200 93.100 18.500 93.800 ;
        RECT 19.800 93.100 20.200 94.800 ;
        RECT 22.500 94.800 25.000 95.100 ;
        RECT 22.500 94.700 22.900 94.800 ;
        RECT 23.800 94.700 24.200 94.800 ;
        RECT 23.300 94.200 23.700 94.300 ;
        RECT 27.000 94.200 27.300 95.800 ;
        RECT 30.200 95.600 30.600 99.900 ;
        RECT 28.500 95.300 30.600 95.600 ;
        RECT 28.500 95.200 28.900 95.300 ;
        RECT 29.300 94.900 29.700 95.000 ;
        RECT 27.800 94.600 29.700 94.900 ;
        RECT 27.800 94.500 28.200 94.600 ;
        RECT 20.600 93.400 21.000 94.200 ;
        RECT 21.800 93.900 27.300 94.200 ;
        RECT 21.800 93.800 22.600 93.900 ;
        RECT 11.000 92.800 11.900 93.100 ;
        RECT 11.500 91.100 11.900 92.800 ;
        RECT 12.600 91.100 13.000 93.100 ;
        RECT 13.400 93.000 15.400 93.100 ;
        RECT 13.400 91.100 13.800 93.000 ;
        RECT 15.000 91.100 15.400 93.000 ;
        RECT 15.800 93.000 17.800 93.100 ;
        RECT 15.800 91.100 16.200 93.000 ;
        RECT 17.400 91.100 17.800 93.000 ;
        RECT 18.200 91.100 18.600 93.100 ;
        RECT 19.300 92.800 20.200 93.100 ;
        RECT 19.300 91.100 19.700 92.800 ;
        RECT 21.400 91.100 21.800 93.500 ;
        RECT 23.900 92.800 24.200 93.900 ;
        RECT 24.600 93.800 25.000 93.900 ;
        RECT 26.700 93.800 27.100 93.900 ;
        RECT 30.200 93.600 30.600 95.300 ;
        RECT 28.700 93.300 30.600 93.600 ;
        RECT 28.700 93.200 29.100 93.300 ;
        RECT 23.000 92.100 23.400 92.500 ;
        RECT 23.800 92.400 24.200 92.800 ;
        RECT 24.700 92.700 25.100 92.800 ;
        RECT 24.700 92.400 26.100 92.700 ;
        RECT 25.800 92.100 26.100 92.400 ;
        RECT 27.800 92.100 28.200 92.500 ;
        RECT 23.000 91.800 24.000 92.100 ;
        RECT 23.600 91.100 24.000 91.800 ;
        RECT 25.800 91.100 26.200 92.100 ;
        RECT 27.800 91.800 28.500 92.100 ;
        RECT 27.900 91.100 28.500 91.800 ;
        RECT 30.200 91.100 30.600 93.300 ;
        RECT 31.000 92.400 31.400 93.200 ;
        RECT 31.800 91.100 32.200 99.900 ;
        RECT 32.600 97.100 33.000 97.200 ;
        RECT 33.400 97.100 33.800 99.900 ;
        RECT 32.600 96.800 33.800 97.100 ;
        RECT 32.600 93.400 33.000 94.200 ;
        RECT 33.400 93.100 33.800 96.800 ;
        RECT 34.200 95.800 34.600 96.600 ;
        RECT 35.800 94.100 36.200 99.900 ;
        RECT 39.500 96.200 39.900 99.900 ;
        RECT 40.200 96.800 40.600 97.200 ;
        RECT 40.300 96.200 40.600 96.800 ;
        RECT 39.500 95.900 40.000 96.200 ;
        RECT 40.300 95.900 41.000 96.200 ;
        RECT 39.000 94.400 39.400 95.200 ;
        RECT 39.700 94.200 40.000 95.900 ;
        RECT 40.600 95.800 41.000 95.900 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 38.200 94.100 38.600 94.200 ;
        RECT 39.700 94.100 41.000 94.200 ;
        RECT 41.400 94.100 41.700 94.800 ;
        RECT 35.800 93.800 39.000 94.100 ;
        RECT 39.700 93.800 41.700 94.100 ;
        RECT 42.200 94.100 42.600 99.900 ;
        RECT 44.300 96.200 45.300 99.900 ;
        RECT 48.300 96.200 48.700 99.900 ;
        RECT 49.000 97.100 49.400 97.200 ;
        RECT 50.200 97.100 50.600 97.200 ;
        RECT 49.000 96.800 50.600 97.100 ;
        RECT 49.100 96.200 49.400 96.800 ;
        RECT 44.300 95.900 45.800 96.200 ;
        RECT 48.300 95.900 48.800 96.200 ;
        RECT 49.100 95.900 49.800 96.200 ;
        RECT 44.600 95.800 45.800 95.900 ;
        RECT 43.800 94.400 44.200 95.200 ;
        RECT 44.600 94.200 44.900 95.800 ;
        RECT 45.400 94.400 45.800 95.200 ;
        RECT 43.000 94.100 43.400 94.200 ;
        RECT 44.600 94.100 45.000 94.200 ;
        RECT 42.200 93.800 43.800 94.100 ;
        RECT 44.600 93.800 45.800 94.100 ;
        RECT 46.200 93.800 46.600 94.600 ;
        RECT 47.800 94.400 48.200 95.200 ;
        RECT 48.500 94.200 48.800 95.900 ;
        RECT 49.400 95.800 49.800 95.900 ;
        RECT 47.000 94.100 47.400 94.200 ;
        RECT 48.500 94.100 49.800 94.200 ;
        RECT 50.200 94.100 50.600 94.200 ;
        RECT 47.000 93.800 47.800 94.100 ;
        RECT 48.500 93.800 50.600 94.100 ;
        RECT 33.400 92.800 34.300 93.100 ;
        RECT 33.900 91.100 34.300 92.800 ;
        RECT 35.000 92.400 35.400 93.200 ;
        RECT 35.800 91.100 36.200 93.800 ;
        RECT 38.600 93.600 39.000 93.800 ;
        RECT 38.300 93.100 40.100 93.300 ;
        RECT 40.600 93.100 40.900 93.800 ;
        RECT 38.200 93.000 40.200 93.100 ;
        RECT 38.200 91.100 38.600 93.000 ;
        RECT 39.800 91.100 40.200 93.000 ;
        RECT 40.600 91.100 41.000 93.100 ;
        RECT 41.400 92.400 41.800 93.200 ;
        RECT 42.200 91.100 42.600 93.800 ;
        RECT 43.400 93.600 43.800 93.800 ;
        RECT 43.100 93.100 44.900 93.300 ;
        RECT 45.500 93.100 45.800 93.800 ;
        RECT 47.400 93.600 47.800 93.800 ;
        RECT 47.100 93.100 48.900 93.300 ;
        RECT 49.400 93.100 49.700 93.800 ;
        RECT 50.200 93.400 50.600 93.800 ;
        RECT 51.000 93.100 51.400 99.900 ;
        RECT 51.800 95.800 52.200 96.600 ;
        RECT 52.600 95.800 53.000 97.200 ;
        RECT 53.400 97.100 53.800 99.900 ;
        RECT 53.400 96.800 54.500 97.100 ;
        RECT 53.400 93.100 53.800 96.800 ;
        RECT 54.200 96.200 54.500 96.800 ;
        RECT 56.300 96.200 56.700 99.900 ;
        RECT 57.000 96.800 57.400 97.200 ;
        RECT 57.100 96.200 57.400 96.800 ;
        RECT 54.200 95.800 54.600 96.200 ;
        RECT 56.300 95.900 56.800 96.200 ;
        RECT 57.100 95.900 57.800 96.200 ;
        RECT 55.800 94.400 56.200 95.200 ;
        RECT 56.500 94.200 56.800 95.900 ;
        RECT 57.400 95.800 57.800 95.900 ;
        RECT 58.200 95.700 58.600 99.900 ;
        RECT 60.400 98.200 60.800 99.900 ;
        RECT 59.800 97.900 60.800 98.200 ;
        RECT 62.600 97.900 63.000 99.900 ;
        RECT 64.700 97.900 65.300 99.900 ;
        RECT 59.800 97.500 60.200 97.900 ;
        RECT 62.600 97.600 62.900 97.900 ;
        RECT 61.500 97.300 63.300 97.600 ;
        RECT 64.600 97.500 65.000 97.900 ;
        RECT 61.500 97.200 61.900 97.300 ;
        RECT 62.900 97.200 63.300 97.300 ;
        RECT 65.100 97.000 65.800 97.200 ;
        RECT 64.700 96.800 65.800 97.000 ;
        RECT 67.000 97.100 67.400 99.900 ;
        RECT 67.800 97.100 68.200 97.200 ;
        RECT 67.000 96.800 68.200 97.100 ;
        RECT 59.800 96.500 60.200 96.600 ;
        RECT 62.100 96.500 62.500 96.600 ;
        RECT 59.800 96.200 62.500 96.500 ;
        RECT 62.800 96.500 63.900 96.800 ;
        RECT 62.800 95.900 63.100 96.500 ;
        RECT 63.500 96.400 63.900 96.500 ;
        RECT 64.700 96.600 65.400 96.800 ;
        RECT 64.700 96.100 65.000 96.600 ;
        RECT 60.700 95.700 63.100 95.900 ;
        RECT 58.200 95.600 63.100 95.700 ;
        RECT 63.800 95.800 65.000 96.100 ;
        RECT 58.200 95.500 61.100 95.600 ;
        RECT 58.200 95.400 61.000 95.500 ;
        RECT 63.800 95.200 64.100 95.800 ;
        RECT 67.000 95.600 67.400 96.800 ;
        RECT 65.300 95.300 67.400 95.600 ;
        RECT 65.300 95.200 65.700 95.300 ;
        RECT 61.400 95.100 61.800 95.200 ;
        RECT 59.300 94.800 61.800 95.100 ;
        RECT 63.800 94.800 64.200 95.200 ;
        RECT 66.100 94.900 66.500 95.000 ;
        RECT 59.300 94.700 59.700 94.800 ;
        RECT 60.100 94.200 60.500 94.300 ;
        RECT 63.800 94.200 64.100 94.800 ;
        RECT 64.600 94.600 66.500 94.900 ;
        RECT 64.600 94.500 65.000 94.600 ;
        RECT 54.200 93.400 54.600 94.200 ;
        RECT 55.000 94.100 55.400 94.200 ;
        RECT 55.000 93.800 55.800 94.100 ;
        RECT 56.500 93.800 57.800 94.200 ;
        RECT 58.600 93.900 64.100 94.200 ;
        RECT 58.600 93.800 59.400 93.900 ;
        RECT 55.400 93.600 55.800 93.800 ;
        RECT 55.100 93.100 56.900 93.300 ;
        RECT 57.400 93.200 57.700 93.800 ;
        RECT 43.000 93.000 45.000 93.100 ;
        RECT 43.000 91.100 43.400 93.000 ;
        RECT 44.600 91.400 45.000 93.000 ;
        RECT 45.400 91.700 45.800 93.100 ;
        RECT 46.200 91.400 46.600 93.100 ;
        RECT 44.600 91.100 46.600 91.400 ;
        RECT 47.000 93.000 49.000 93.100 ;
        RECT 47.000 91.100 47.400 93.000 ;
        RECT 48.600 91.100 49.000 93.000 ;
        RECT 49.400 91.100 49.800 93.100 ;
        RECT 51.000 92.800 51.900 93.100 ;
        RECT 51.500 92.200 51.900 92.800 ;
        RECT 52.900 92.800 53.800 93.100 ;
        RECT 55.000 93.000 57.000 93.100 ;
        RECT 51.500 91.800 52.200 92.200 ;
        RECT 51.500 91.100 51.900 91.800 ;
        RECT 52.900 91.100 53.300 92.800 ;
        RECT 55.000 91.100 55.400 93.000 ;
        RECT 56.600 91.100 57.000 93.000 ;
        RECT 57.400 91.100 57.800 93.200 ;
        RECT 58.200 91.100 58.600 93.500 ;
        RECT 60.700 92.800 61.000 93.900 ;
        RECT 63.500 93.800 63.900 93.900 ;
        RECT 67.000 93.600 67.400 95.300 ;
        RECT 68.600 95.100 69.000 99.900 ;
        RECT 70.600 96.800 71.000 97.200 ;
        RECT 69.400 95.800 69.800 96.600 ;
        RECT 70.600 96.200 70.900 96.800 ;
        RECT 71.300 96.200 71.700 99.900 ;
        RECT 74.200 96.400 74.600 99.900 ;
        RECT 70.200 95.900 70.900 96.200 ;
        RECT 71.200 95.900 71.700 96.200 ;
        RECT 74.100 95.900 74.600 96.400 ;
        RECT 75.800 96.200 76.200 99.900 ;
        RECT 74.900 95.900 76.200 96.200 ;
        RECT 77.900 96.200 78.300 99.900 ;
        RECT 78.600 96.800 79.000 97.200 ;
        RECT 78.700 96.200 79.000 96.800 ;
        RECT 77.900 95.900 78.400 96.200 ;
        RECT 78.700 95.900 79.400 96.200 ;
        RECT 70.200 95.800 70.600 95.900 ;
        RECT 70.200 95.100 70.500 95.800 ;
        RECT 68.600 94.800 70.500 95.100 ;
        RECT 65.400 93.300 67.400 93.600 ;
        RECT 67.800 93.400 68.200 94.200 ;
        RECT 65.400 93.200 65.900 93.300 ;
        RECT 65.400 92.800 65.800 93.200 ;
        RECT 59.800 92.100 60.200 92.500 ;
        RECT 60.600 92.400 61.000 92.800 ;
        RECT 61.500 92.700 61.900 92.800 ;
        RECT 61.500 92.400 62.900 92.700 ;
        RECT 62.600 92.100 62.900 92.400 ;
        RECT 64.600 92.100 65.000 92.500 ;
        RECT 59.800 91.800 60.800 92.100 ;
        RECT 60.400 91.100 60.800 91.800 ;
        RECT 62.600 91.100 63.000 92.100 ;
        RECT 64.600 91.800 65.300 92.100 ;
        RECT 64.700 91.100 65.300 91.800 ;
        RECT 67.000 91.100 67.400 93.300 ;
        RECT 68.600 93.100 69.000 94.800 ;
        RECT 71.200 94.200 71.500 95.900 ;
        RECT 71.800 94.400 72.200 95.200 ;
        RECT 74.100 94.200 74.400 95.900 ;
        RECT 74.900 94.900 75.200 95.900 ;
        RECT 74.700 94.500 75.200 94.900 ;
        RECT 69.400 94.100 69.800 94.200 ;
        RECT 70.200 94.100 71.500 94.200 ;
        RECT 72.600 94.100 73.000 94.200 ;
        RECT 69.400 93.800 71.500 94.100 ;
        RECT 72.200 93.800 73.000 94.100 ;
        RECT 74.100 93.800 74.600 94.200 ;
        RECT 70.300 93.100 70.600 93.800 ;
        RECT 72.200 93.600 72.600 93.800 ;
        RECT 71.100 93.100 72.900 93.300 ;
        RECT 74.100 93.100 74.400 93.800 ;
        RECT 74.900 93.700 75.200 94.500 ;
        RECT 75.700 94.800 76.200 95.200 ;
        RECT 75.700 94.400 76.100 94.800 ;
        RECT 77.400 94.400 77.800 95.200 ;
        RECT 78.100 95.100 78.400 95.900 ;
        RECT 79.000 95.800 79.400 95.900 ;
        RECT 79.800 95.600 80.200 99.900 ;
        RECT 81.900 97.900 82.500 99.900 ;
        RECT 84.200 97.900 84.600 99.900 ;
        RECT 86.400 98.200 86.800 99.900 ;
        RECT 86.400 97.900 87.400 98.200 ;
        RECT 82.200 97.500 82.600 97.900 ;
        RECT 84.300 97.600 84.600 97.900 ;
        RECT 83.900 97.300 85.700 97.600 ;
        RECT 87.000 97.500 87.400 97.900 ;
        RECT 83.900 97.200 84.300 97.300 ;
        RECT 85.300 97.200 85.700 97.300 ;
        RECT 81.800 96.600 82.500 97.000 ;
        RECT 82.200 96.100 82.500 96.600 ;
        RECT 83.300 96.500 84.400 96.800 ;
        RECT 83.300 96.400 83.700 96.500 ;
        RECT 82.200 95.800 83.400 96.100 ;
        RECT 79.800 95.300 81.900 95.600 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 78.100 94.800 79.400 95.100 ;
        RECT 78.100 94.200 78.400 94.800 ;
        RECT 76.600 94.100 77.000 94.200 ;
        RECT 76.600 93.800 77.400 94.100 ;
        RECT 78.100 93.800 79.400 94.200 ;
        RECT 74.900 93.400 76.200 93.700 ;
        RECT 77.000 93.600 77.400 93.800 ;
        RECT 68.600 92.800 69.500 93.100 ;
        RECT 69.100 91.100 69.500 92.800 ;
        RECT 70.200 91.100 70.600 93.100 ;
        RECT 71.000 93.000 73.000 93.100 ;
        RECT 71.000 91.100 71.400 93.000 ;
        RECT 72.600 91.100 73.000 93.000 ;
        RECT 74.100 92.800 74.600 93.100 ;
        RECT 74.200 91.100 74.600 92.800 ;
        RECT 75.800 91.100 76.200 93.400 ;
        RECT 76.700 93.100 78.500 93.300 ;
        RECT 79.000 93.100 79.300 93.800 ;
        RECT 79.800 93.600 80.200 95.300 ;
        RECT 81.500 95.200 81.900 95.300 ;
        RECT 80.700 94.900 81.100 95.000 ;
        RECT 80.700 94.600 82.600 94.900 ;
        RECT 82.200 94.500 82.600 94.600 ;
        RECT 83.100 94.200 83.400 95.800 ;
        RECT 84.100 95.900 84.400 96.500 ;
        RECT 84.700 96.500 85.100 96.600 ;
        RECT 87.000 96.500 87.400 96.600 ;
        RECT 84.700 96.200 87.400 96.500 ;
        RECT 84.100 95.700 86.500 95.900 ;
        RECT 88.600 95.700 89.000 99.900 ;
        RECT 84.100 95.600 89.000 95.700 ;
        RECT 86.100 95.500 89.000 95.600 ;
        RECT 86.200 95.400 89.000 95.500 ;
        RECT 85.400 95.100 85.800 95.200 ;
        RECT 85.400 94.800 87.900 95.100 ;
        RECT 87.500 94.700 87.900 94.800 ;
        RECT 86.700 94.200 87.100 94.300 ;
        RECT 83.100 93.900 88.600 94.200 ;
        RECT 83.300 93.800 83.700 93.900 ;
        RECT 85.400 93.800 85.800 93.900 ;
        RECT 79.800 93.300 81.700 93.600 ;
        RECT 76.600 93.000 78.600 93.100 ;
        RECT 76.600 91.100 77.000 93.000 ;
        RECT 78.200 91.100 78.600 93.000 ;
        RECT 79.000 91.100 79.400 93.100 ;
        RECT 79.800 91.100 80.200 93.300 ;
        RECT 81.300 93.200 81.700 93.300 ;
        RECT 86.200 92.800 86.500 93.900 ;
        RECT 87.800 93.800 88.600 93.900 ;
        RECT 89.400 94.100 89.800 94.200 ;
        RECT 91.000 94.100 91.400 94.200 ;
        RECT 89.400 93.800 91.400 94.100 ;
        RECT 85.300 92.700 85.700 92.800 ;
        RECT 82.200 92.100 82.600 92.500 ;
        RECT 84.300 92.400 85.700 92.700 ;
        RECT 86.200 92.400 86.600 92.800 ;
        RECT 84.300 92.100 84.600 92.400 ;
        RECT 87.000 92.100 87.400 92.500 ;
        RECT 81.900 91.800 82.600 92.100 ;
        RECT 81.900 91.100 82.500 91.800 ;
        RECT 84.200 91.100 84.600 92.100 ;
        RECT 86.400 91.800 87.400 92.100 ;
        RECT 86.400 91.100 86.800 91.800 ;
        RECT 88.600 91.100 89.000 93.500 ;
        RECT 91.000 93.400 91.400 93.800 ;
        RECT 91.800 93.100 92.200 99.900 ;
        RECT 93.400 97.900 93.800 99.900 ;
        RECT 93.500 97.800 93.800 97.900 ;
        RECT 95.000 97.900 95.400 99.900 ;
        RECT 95.000 97.800 95.300 97.900 ;
        RECT 93.500 97.500 95.300 97.800 ;
        RECT 92.600 95.800 93.000 96.600 ;
        RECT 93.500 96.200 93.800 97.500 ;
        RECT 94.200 96.400 94.600 97.200 ;
        RECT 93.400 95.800 93.800 96.200 ;
        RECT 93.500 94.200 93.800 95.800 ;
        RECT 95.800 95.400 96.200 96.200 ;
        RECT 96.600 95.800 97.000 96.600 ;
        RECT 94.600 94.800 95.400 95.200 ;
        RECT 93.500 94.100 94.300 94.200 ;
        RECT 93.500 93.900 94.400 94.100 ;
        RECT 91.800 92.800 92.700 93.100 ;
        RECT 92.300 92.200 92.700 92.800 ;
        RECT 92.300 91.800 93.000 92.200 ;
        RECT 92.300 91.100 92.700 91.800 ;
        RECT 94.000 91.100 94.400 93.900 ;
        RECT 97.400 93.100 97.800 99.900 ;
        RECT 98.200 93.400 98.600 94.200 ;
        RECT 99.000 93.400 99.400 94.200 ;
        RECT 96.900 92.800 97.800 93.100 ;
        RECT 99.800 93.100 100.200 99.900 ;
        RECT 101.800 96.800 102.200 97.200 ;
        RECT 100.600 95.800 101.000 96.600 ;
        RECT 101.800 96.200 102.100 96.800 ;
        RECT 102.500 96.200 102.900 99.900 ;
        RECT 101.400 95.900 102.100 96.200 ;
        RECT 102.400 95.900 102.900 96.200 ;
        RECT 101.400 95.800 101.800 95.900 ;
        RECT 102.400 95.200 102.700 95.900 ;
        RECT 104.600 95.800 105.000 96.600 ;
        RECT 102.200 94.800 102.700 95.200 ;
        RECT 102.400 94.200 102.700 94.800 ;
        RECT 103.000 94.400 103.400 95.200 ;
        RECT 101.400 93.800 102.700 94.200 ;
        RECT 103.800 94.100 104.200 94.200 ;
        RECT 103.400 93.800 104.200 94.100 ;
        RECT 101.500 93.100 101.800 93.800 ;
        RECT 103.400 93.600 103.800 93.800 ;
        RECT 102.300 93.100 104.100 93.300 ;
        RECT 105.400 93.100 105.800 99.900 ;
        RECT 107.000 95.800 107.400 96.600 ;
        RECT 106.200 94.100 106.600 94.200 ;
        RECT 107.000 94.100 107.400 94.200 ;
        RECT 106.200 93.800 107.400 94.100 ;
        RECT 106.200 93.400 106.600 93.800 ;
        RECT 107.800 93.100 108.200 99.900 ;
        RECT 111.300 96.400 111.700 99.900 ;
        RECT 113.400 97.500 113.800 99.500 ;
        RECT 110.900 96.100 111.700 96.400 ;
        RECT 109.400 95.100 109.800 95.200 ;
        RECT 110.200 95.100 110.600 95.600 ;
        RECT 109.400 94.800 110.600 95.100 ;
        RECT 110.900 94.200 111.200 96.100 ;
        RECT 113.500 95.800 113.800 97.500 ;
        RECT 114.200 95.800 114.600 96.600 ;
        RECT 111.900 95.500 113.800 95.800 ;
        RECT 111.900 94.500 112.200 95.500 ;
        RECT 108.600 93.400 109.000 94.200 ;
        RECT 110.200 93.800 111.200 94.200 ;
        RECT 111.500 94.100 112.200 94.500 ;
        RECT 112.600 94.400 113.000 95.200 ;
        RECT 113.400 94.400 113.800 95.200 ;
        RECT 110.900 93.500 111.200 93.800 ;
        RECT 111.700 93.900 112.200 94.100 ;
        RECT 111.700 93.600 113.800 93.900 ;
        RECT 99.800 92.800 100.700 93.100 ;
        RECT 96.900 91.100 97.300 92.800 ;
        RECT 100.300 92.200 100.700 92.800 ;
        RECT 100.300 91.800 101.000 92.200 ;
        RECT 100.300 91.100 100.700 91.800 ;
        RECT 101.400 91.100 101.800 93.100 ;
        RECT 102.200 93.000 104.200 93.100 ;
        RECT 102.200 91.100 102.600 93.000 ;
        RECT 103.800 91.100 104.200 93.000 ;
        RECT 104.900 92.800 105.800 93.100 ;
        RECT 107.300 92.800 108.200 93.100 ;
        RECT 110.900 93.300 111.300 93.500 ;
        RECT 110.900 93.000 111.700 93.300 ;
        RECT 104.900 92.200 105.300 92.800 ;
        RECT 107.300 92.200 107.700 92.800 ;
        RECT 104.600 91.800 105.300 92.200 ;
        RECT 107.000 91.800 107.700 92.200 ;
        RECT 104.900 91.100 105.300 91.800 ;
        RECT 107.300 91.100 107.700 91.800 ;
        RECT 111.300 91.500 111.700 93.000 ;
        RECT 113.500 92.500 113.800 93.600 ;
        RECT 115.000 93.100 115.400 99.900 ;
        RECT 117.400 96.400 117.800 99.900 ;
        RECT 117.300 95.900 117.800 96.400 ;
        RECT 119.000 96.200 119.400 99.900 ;
        RECT 120.600 96.400 121.000 99.900 ;
        RECT 118.100 95.900 119.400 96.200 ;
        RECT 120.500 95.900 121.000 96.400 ;
        RECT 122.200 96.200 122.600 99.900 ;
        RECT 121.300 95.900 122.600 96.200 ;
        RECT 117.300 94.200 117.600 95.900 ;
        RECT 118.100 94.900 118.400 95.900 ;
        RECT 117.900 94.500 118.400 94.900 ;
        RECT 115.800 93.400 116.200 94.200 ;
        RECT 117.300 93.800 117.800 94.200 ;
        RECT 113.400 91.500 113.800 92.500 ;
        RECT 114.500 92.800 115.400 93.100 ;
        RECT 117.300 93.100 117.600 93.800 ;
        RECT 118.100 93.700 118.400 94.500 ;
        RECT 118.900 95.100 119.400 95.200 ;
        RECT 119.800 95.100 120.200 95.200 ;
        RECT 118.900 94.800 120.200 95.100 ;
        RECT 118.900 94.400 119.300 94.800 ;
        RECT 120.500 94.200 120.800 95.900 ;
        RECT 121.300 94.900 121.600 95.900 ;
        RECT 123.000 95.800 123.400 96.600 ;
        RECT 121.100 94.500 121.600 94.900 ;
        RECT 120.500 93.800 121.000 94.200 ;
        RECT 118.100 93.400 119.400 93.700 ;
        RECT 117.300 92.800 117.800 93.100 ;
        RECT 114.500 92.200 114.900 92.800 ;
        RECT 114.500 91.800 115.400 92.200 ;
        RECT 114.500 91.100 114.900 91.800 ;
        RECT 117.400 91.100 117.800 92.800 ;
        RECT 119.000 91.100 119.400 93.400 ;
        RECT 120.500 93.100 120.800 93.800 ;
        RECT 121.300 93.700 121.600 94.500 ;
        RECT 122.100 94.800 122.600 95.200 ;
        RECT 122.100 94.400 122.500 94.800 ;
        RECT 121.300 93.400 122.600 93.700 ;
        RECT 120.500 92.800 121.000 93.100 ;
        RECT 120.600 91.100 121.000 92.800 ;
        RECT 122.200 91.100 122.600 93.400 ;
        RECT 123.800 93.100 124.200 99.900 ;
        RECT 125.400 99.600 127.400 99.900 ;
        RECT 125.400 95.900 125.800 99.600 ;
        RECT 126.200 95.900 126.600 99.300 ;
        RECT 127.000 96.200 127.400 99.600 ;
        RECT 128.600 96.200 129.000 99.900 ;
        RECT 127.000 95.900 129.000 96.200 ;
        RECT 126.300 95.600 126.600 95.900 ;
        RECT 124.600 95.100 125.000 95.200 ;
        RECT 125.400 95.100 125.800 95.600 ;
        RECT 126.300 95.300 127.300 95.600 ;
        RECT 124.600 94.800 125.800 95.100 ;
        RECT 127.000 95.200 127.300 95.300 ;
        RECT 128.200 95.200 128.600 95.400 ;
        RECT 127.000 94.800 127.400 95.200 ;
        RECT 128.200 94.900 129.000 95.200 ;
        RECT 128.600 94.800 129.000 94.900 ;
        RECT 126.300 94.400 126.700 94.800 ;
        RECT 126.300 94.200 126.600 94.400 ;
        RECT 124.600 94.100 125.000 94.200 ;
        RECT 125.400 94.100 125.800 94.200 ;
        RECT 124.600 93.800 125.800 94.100 ;
        RECT 126.200 93.800 126.600 94.200 ;
        RECT 124.600 93.400 125.000 93.800 ;
        RECT 127.000 93.100 127.300 94.800 ;
        RECT 127.800 93.800 128.200 94.600 ;
        RECT 123.300 92.800 124.200 93.100 ;
        RECT 123.300 92.200 123.700 92.800 ;
        RECT 123.300 91.800 124.200 92.200 ;
        RECT 123.300 91.100 123.700 91.800 ;
        RECT 126.700 91.100 127.500 93.100 ;
        RECT 129.400 91.100 129.800 99.900 ;
        RECT 131.000 95.800 131.400 96.600 ;
        RECT 131.800 96.100 132.200 99.900 ;
        RECT 133.800 96.800 134.200 97.200 ;
        RECT 133.800 96.200 134.100 96.800 ;
        RECT 134.500 96.200 134.900 99.900 ;
        RECT 133.400 96.100 134.100 96.200 ;
        RECT 131.800 95.900 134.100 96.100 ;
        RECT 134.400 95.900 134.900 96.200 ;
        RECT 131.800 95.800 133.800 95.900 ;
        RECT 130.200 92.400 130.600 93.200 ;
        RECT 131.800 93.100 132.200 95.800 ;
        RECT 132.600 95.100 133.000 95.200 ;
        RECT 134.400 95.100 134.700 95.900 ;
        RECT 138.200 95.700 138.600 99.900 ;
        RECT 140.400 98.200 140.800 99.900 ;
        RECT 139.800 97.900 140.800 98.200 ;
        RECT 142.600 97.900 143.000 99.900 ;
        RECT 144.700 97.900 145.300 99.900 ;
        RECT 139.800 97.500 140.200 97.900 ;
        RECT 142.600 97.600 142.900 97.900 ;
        RECT 141.500 97.300 143.300 97.600 ;
        RECT 144.600 97.500 145.000 97.900 ;
        RECT 141.500 97.200 141.900 97.300 ;
        RECT 142.900 97.200 143.300 97.300 ;
        RECT 139.800 96.500 140.200 96.600 ;
        RECT 142.100 96.500 142.500 96.600 ;
        RECT 139.800 96.200 142.500 96.500 ;
        RECT 142.800 96.500 143.900 96.800 ;
        RECT 142.800 95.900 143.100 96.500 ;
        RECT 143.500 96.400 143.900 96.500 ;
        RECT 144.700 96.600 145.400 97.000 ;
        RECT 144.700 96.100 145.000 96.600 ;
        RECT 140.700 95.700 143.100 95.900 ;
        RECT 138.200 95.600 143.100 95.700 ;
        RECT 143.800 95.800 145.000 96.100 ;
        RECT 138.200 95.500 141.100 95.600 ;
        RECT 138.200 95.400 141.000 95.500 ;
        RECT 143.800 95.200 144.100 95.800 ;
        RECT 147.000 95.600 147.400 99.900 ;
        RECT 148.200 96.800 148.600 97.200 ;
        RECT 148.200 96.200 148.500 96.800 ;
        RECT 148.900 96.200 149.300 99.900 ;
        RECT 152.100 99.200 152.500 99.900 ;
        RECT 152.100 98.800 153.000 99.200 ;
        RECT 151.400 96.800 151.800 97.200 ;
        RECT 151.400 96.200 151.700 96.800 ;
        RECT 152.100 96.200 152.500 98.800 ;
        RECT 155.000 96.400 155.400 99.900 ;
        RECT 147.800 95.900 148.500 96.200 ;
        RECT 148.800 95.900 149.300 96.200 ;
        RECT 151.000 95.900 151.700 96.200 ;
        RECT 152.000 95.900 152.500 96.200 ;
        RECT 154.900 95.900 155.400 96.400 ;
        RECT 156.600 96.200 157.000 99.900 ;
        RECT 155.700 95.900 157.000 96.200 ;
        RECT 157.400 96.200 157.800 99.900 ;
        RECT 159.000 96.400 159.400 99.900 ;
        RECT 157.400 95.900 158.700 96.200 ;
        RECT 159.000 95.900 159.500 96.400 ;
        RECT 147.800 95.800 148.200 95.900 ;
        RECT 145.300 95.300 147.400 95.600 ;
        RECT 145.300 95.200 145.700 95.300 ;
        RECT 132.600 94.800 134.700 95.100 ;
        RECT 134.400 94.200 134.700 94.800 ;
        RECT 135.000 95.100 135.400 95.200 ;
        RECT 135.800 95.100 136.200 95.200 ;
        RECT 141.400 95.100 141.800 95.200 ;
        RECT 142.200 95.100 142.600 95.200 ;
        RECT 135.000 94.800 136.200 95.100 ;
        RECT 139.300 94.800 142.600 95.100 ;
        RECT 143.800 94.800 144.200 95.200 ;
        RECT 146.100 94.900 146.500 95.000 ;
        RECT 135.000 94.400 135.400 94.800 ;
        RECT 139.300 94.700 139.700 94.800 ;
        RECT 140.100 94.200 140.500 94.300 ;
        RECT 143.800 94.200 144.100 94.800 ;
        RECT 144.600 94.600 146.500 94.900 ;
        RECT 144.600 94.500 145.000 94.600 ;
        RECT 132.600 93.400 133.000 94.200 ;
        RECT 133.400 93.800 134.700 94.200 ;
        RECT 135.800 94.100 136.200 94.200 ;
        RECT 135.400 93.800 136.200 94.100 ;
        RECT 138.600 93.900 144.100 94.200 ;
        RECT 138.600 93.800 139.400 93.900 ;
        RECT 133.500 93.100 133.800 93.800 ;
        RECT 135.400 93.600 135.800 93.800 ;
        RECT 134.300 93.100 136.100 93.300 ;
        RECT 131.300 92.800 132.200 93.100 ;
        RECT 131.300 91.100 131.700 92.800 ;
        RECT 133.400 91.100 133.800 93.100 ;
        RECT 134.200 93.000 136.200 93.100 ;
        RECT 134.200 91.100 134.600 93.000 ;
        RECT 135.800 91.100 136.200 93.000 ;
        RECT 138.200 91.100 138.600 93.500 ;
        RECT 140.700 92.800 141.000 93.900 ;
        RECT 143.500 93.800 143.900 93.900 ;
        RECT 147.000 93.600 147.400 95.300 ;
        RECT 147.800 95.100 148.200 95.200 ;
        RECT 148.800 95.100 149.100 95.900 ;
        RECT 151.000 95.800 151.400 95.900 ;
        RECT 147.800 94.800 149.100 95.100 ;
        RECT 148.800 94.200 149.100 94.800 ;
        RECT 149.400 94.400 149.800 95.200 ;
        RECT 152.000 94.200 152.300 95.900 ;
        RECT 152.600 94.400 153.000 95.200 ;
        RECT 154.900 94.200 155.200 95.900 ;
        RECT 155.700 94.900 156.000 95.900 ;
        RECT 155.500 94.500 156.000 94.900 ;
        RECT 147.800 93.800 149.100 94.200 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 149.800 93.800 150.600 94.100 ;
        RECT 151.000 93.800 152.300 94.200 ;
        RECT 153.400 94.100 153.800 94.200 ;
        RECT 154.200 94.100 154.600 94.200 ;
        RECT 153.000 93.800 154.600 94.100 ;
        RECT 154.900 93.800 155.400 94.200 ;
        RECT 145.500 93.300 147.400 93.600 ;
        RECT 145.500 93.200 145.900 93.300 ;
        RECT 139.800 92.100 140.200 92.500 ;
        RECT 140.600 92.400 141.000 92.800 ;
        RECT 141.500 92.700 141.900 92.800 ;
        RECT 141.500 92.400 142.900 92.700 ;
        RECT 142.600 92.100 142.900 92.400 ;
        RECT 144.600 92.100 145.000 92.500 ;
        RECT 139.800 91.800 140.800 92.100 ;
        RECT 140.400 91.100 140.800 91.800 ;
        RECT 142.600 91.100 143.000 92.100 ;
        RECT 144.600 91.800 145.300 92.100 ;
        RECT 144.700 91.100 145.300 91.800 ;
        RECT 147.000 91.100 147.400 93.300 ;
        RECT 147.900 93.100 148.200 93.800 ;
        RECT 149.800 93.600 150.200 93.800 ;
        RECT 148.700 93.100 150.500 93.300 ;
        RECT 151.100 93.100 151.400 93.800 ;
        RECT 153.000 93.600 153.400 93.800 ;
        RECT 151.900 93.100 153.700 93.300 ;
        RECT 154.900 93.100 155.200 93.800 ;
        RECT 155.700 93.700 156.000 94.500 ;
        RECT 156.500 95.100 157.000 95.200 ;
        RECT 157.400 95.100 157.900 95.200 ;
        RECT 156.500 94.800 157.900 95.100 ;
        RECT 156.500 94.400 156.900 94.800 ;
        RECT 157.500 94.400 157.900 94.800 ;
        RECT 158.400 94.900 158.700 95.900 ;
        RECT 158.400 94.500 158.900 94.900 ;
        RECT 158.400 93.700 158.700 94.500 ;
        RECT 159.200 94.200 159.500 95.900 ;
        RECT 160.600 95.700 161.000 99.900 ;
        RECT 162.800 98.200 163.200 99.900 ;
        RECT 162.200 97.900 163.200 98.200 ;
        RECT 165.000 97.900 165.400 99.900 ;
        RECT 167.100 97.900 167.700 99.900 ;
        RECT 162.200 97.500 162.600 97.900 ;
        RECT 165.000 97.600 165.300 97.900 ;
        RECT 163.900 97.300 165.700 97.600 ;
        RECT 167.000 97.500 167.400 97.900 ;
        RECT 163.900 97.200 164.300 97.300 ;
        RECT 165.300 97.200 165.700 97.300 ;
        RECT 162.200 96.500 162.600 96.600 ;
        RECT 164.500 96.500 164.900 96.600 ;
        RECT 162.200 96.200 164.900 96.500 ;
        RECT 165.200 96.500 166.300 96.800 ;
        RECT 165.200 95.900 165.500 96.500 ;
        RECT 165.900 96.400 166.300 96.500 ;
        RECT 167.100 96.600 167.800 97.000 ;
        RECT 167.100 96.100 167.400 96.600 ;
        RECT 163.100 95.700 165.500 95.900 ;
        RECT 160.600 95.600 165.500 95.700 ;
        RECT 166.200 95.800 167.400 96.100 ;
        RECT 160.600 95.500 163.500 95.600 ;
        RECT 160.600 95.400 163.400 95.500 ;
        RECT 166.200 95.200 166.500 95.800 ;
        RECT 169.400 95.600 169.800 99.900 ;
        RECT 167.700 95.300 169.800 95.600 ;
        RECT 170.200 95.700 170.600 99.900 ;
        RECT 172.400 98.200 172.800 99.900 ;
        RECT 171.800 97.900 172.800 98.200 ;
        RECT 174.600 97.900 175.000 99.900 ;
        RECT 176.700 97.900 177.300 99.900 ;
        RECT 171.800 97.500 172.200 97.900 ;
        RECT 174.600 97.600 174.900 97.900 ;
        RECT 173.500 97.300 175.300 97.600 ;
        RECT 176.600 97.500 177.000 97.900 ;
        RECT 173.500 97.200 173.900 97.300 ;
        RECT 174.900 97.200 175.300 97.300 ;
        RECT 171.800 96.500 172.200 96.600 ;
        RECT 174.100 96.500 174.500 96.600 ;
        RECT 171.800 96.200 174.500 96.500 ;
        RECT 174.800 96.500 175.900 96.800 ;
        RECT 174.800 95.900 175.100 96.500 ;
        RECT 175.500 96.400 175.900 96.500 ;
        RECT 176.700 96.600 177.400 97.000 ;
        RECT 176.700 96.100 177.000 96.600 ;
        RECT 172.700 95.700 175.100 95.900 ;
        RECT 170.200 95.600 175.100 95.700 ;
        RECT 175.800 95.800 177.000 96.100 ;
        RECT 170.200 95.500 173.100 95.600 ;
        RECT 170.200 95.400 173.000 95.500 ;
        RECT 167.700 95.200 168.100 95.300 ;
        RECT 163.800 95.100 164.200 95.200 ;
        RECT 161.700 94.800 164.200 95.100 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 168.500 94.900 168.900 95.000 ;
        RECT 161.700 94.700 162.100 94.800 ;
        RECT 163.000 94.700 163.400 94.800 ;
        RECT 162.500 94.200 162.900 94.300 ;
        RECT 166.200 94.200 166.500 94.800 ;
        RECT 167.000 94.600 168.900 94.900 ;
        RECT 167.000 94.500 167.400 94.600 ;
        RECT 159.000 93.800 159.500 94.200 ;
        RECT 161.000 93.900 166.500 94.200 ;
        RECT 161.000 93.800 161.800 93.900 ;
        RECT 155.700 93.400 157.000 93.700 ;
        RECT 147.800 91.100 148.200 93.100 ;
        RECT 148.600 93.000 150.600 93.100 ;
        RECT 148.600 91.100 149.000 93.000 ;
        RECT 150.200 91.100 150.600 93.000 ;
        RECT 151.000 91.100 151.400 93.100 ;
        RECT 151.800 93.000 153.800 93.100 ;
        RECT 151.800 91.100 152.200 93.000 ;
        RECT 153.400 91.100 153.800 93.000 ;
        RECT 154.900 92.800 155.400 93.100 ;
        RECT 155.000 91.100 155.400 92.800 ;
        RECT 156.600 91.100 157.000 93.400 ;
        RECT 157.400 93.400 158.700 93.700 ;
        RECT 157.400 91.100 157.800 93.400 ;
        RECT 159.200 93.100 159.500 93.800 ;
        RECT 159.000 92.800 159.500 93.100 ;
        RECT 159.000 91.100 159.400 92.800 ;
        RECT 160.600 91.100 161.000 93.500 ;
        RECT 163.100 92.800 163.400 93.900 ;
        RECT 165.900 93.800 166.300 93.900 ;
        RECT 169.400 93.600 169.800 95.300 ;
        RECT 175.800 95.200 176.100 95.800 ;
        RECT 179.000 95.600 179.400 99.900 ;
        RECT 181.100 97.200 181.500 99.900 ;
        RECT 180.600 96.800 181.500 97.200 ;
        RECT 181.800 96.800 182.200 97.200 ;
        RECT 181.100 96.200 181.500 96.800 ;
        RECT 181.900 96.200 182.200 96.800 ;
        RECT 181.100 95.900 181.600 96.200 ;
        RECT 181.900 95.900 182.600 96.200 ;
        RECT 177.300 95.300 179.400 95.600 ;
        RECT 177.300 95.200 177.700 95.300 ;
        RECT 173.400 95.100 173.800 95.200 ;
        RECT 174.200 95.100 174.600 95.200 ;
        RECT 171.300 94.800 174.600 95.100 ;
        RECT 175.800 94.800 176.200 95.200 ;
        RECT 178.100 94.900 178.500 95.000 ;
        RECT 171.300 94.700 171.700 94.800 ;
        RECT 172.100 94.200 172.500 94.300 ;
        RECT 175.800 94.200 176.100 94.800 ;
        RECT 176.600 94.600 178.500 94.900 ;
        RECT 176.600 94.500 177.000 94.600 ;
        RECT 170.600 93.900 176.100 94.200 ;
        RECT 170.600 93.800 171.400 93.900 ;
        RECT 167.900 93.300 169.800 93.600 ;
        RECT 167.900 93.200 168.300 93.300 ;
        RECT 162.200 92.100 162.600 92.500 ;
        RECT 163.000 92.400 163.400 92.800 ;
        RECT 163.900 92.700 164.300 92.800 ;
        RECT 163.900 92.400 165.300 92.700 ;
        RECT 165.000 92.100 165.300 92.400 ;
        RECT 167.000 92.100 167.400 92.500 ;
        RECT 162.200 91.800 163.200 92.100 ;
        RECT 162.800 91.100 163.200 91.800 ;
        RECT 165.000 91.100 165.400 92.100 ;
        RECT 167.000 91.800 167.700 92.100 ;
        RECT 167.100 91.100 167.700 91.800 ;
        RECT 169.400 91.100 169.800 93.300 ;
        RECT 170.200 91.100 170.600 93.500 ;
        RECT 172.700 92.800 173.000 93.900 ;
        RECT 175.500 93.800 175.900 93.900 ;
        RECT 179.000 93.600 179.400 95.300 ;
        RECT 179.800 95.100 180.200 95.200 ;
        RECT 180.600 95.100 181.000 95.200 ;
        RECT 179.800 94.800 181.000 95.100 ;
        RECT 180.600 94.400 181.000 94.800 ;
        RECT 181.300 94.200 181.600 95.900 ;
        RECT 182.200 95.800 182.600 95.900 ;
        RECT 183.000 95.800 183.400 96.600 ;
        RECT 182.200 95.100 182.500 95.800 ;
        RECT 183.800 95.100 184.200 99.900 ;
        RECT 186.200 96.400 186.600 99.900 ;
        RECT 182.200 94.800 184.200 95.100 ;
        RECT 179.800 94.100 180.200 94.200 ;
        RECT 179.800 93.800 180.600 94.100 ;
        RECT 181.300 93.800 182.600 94.200 ;
        RECT 180.200 93.600 180.600 93.800 ;
        RECT 177.500 93.300 179.400 93.600 ;
        RECT 177.500 93.200 177.900 93.300 ;
        RECT 171.800 92.100 172.200 92.500 ;
        RECT 172.600 92.400 173.000 92.800 ;
        RECT 173.500 92.700 173.900 92.800 ;
        RECT 173.500 92.400 174.900 92.700 ;
        RECT 174.600 92.100 174.900 92.400 ;
        RECT 176.600 92.100 177.000 92.500 ;
        RECT 171.800 91.800 172.800 92.100 ;
        RECT 172.400 91.100 172.800 91.800 ;
        RECT 174.600 91.100 175.000 92.100 ;
        RECT 176.600 91.800 177.300 92.100 ;
        RECT 176.700 91.100 177.300 91.800 ;
        RECT 179.000 91.100 179.400 93.300 ;
        RECT 179.900 93.100 181.700 93.300 ;
        RECT 182.200 93.100 182.500 93.800 ;
        RECT 183.800 93.100 184.200 94.800 ;
        RECT 186.100 95.900 186.600 96.400 ;
        RECT 187.800 96.200 188.200 99.900 ;
        RECT 186.900 95.900 188.200 96.200 ;
        RECT 186.100 94.200 186.400 95.900 ;
        RECT 186.900 94.900 187.200 95.900 ;
        RECT 186.700 94.500 187.200 94.900 ;
        RECT 184.600 93.400 185.000 94.200 ;
        RECT 186.100 93.800 186.600 94.200 ;
        RECT 179.800 93.000 181.800 93.100 ;
        RECT 179.800 91.100 180.200 93.000 ;
        RECT 181.400 91.100 181.800 93.000 ;
        RECT 182.200 91.100 182.600 93.100 ;
        RECT 183.300 92.800 184.200 93.100 ;
        RECT 186.100 93.100 186.400 93.800 ;
        RECT 186.900 93.700 187.200 94.500 ;
        RECT 187.700 94.800 188.200 95.200 ;
        RECT 187.700 94.400 188.100 94.800 ;
        RECT 186.900 93.400 188.200 93.700 ;
        RECT 188.600 93.400 189.000 94.200 ;
        RECT 186.100 92.800 186.600 93.100 ;
        RECT 183.300 91.100 183.700 92.800 ;
        RECT 186.200 91.100 186.600 92.800 ;
        RECT 187.800 91.100 188.200 93.400 ;
        RECT 189.400 93.100 189.800 99.900 ;
        RECT 191.800 97.100 192.200 97.200 ;
        RECT 190.200 96.800 192.200 97.100 ;
        RECT 190.200 95.800 190.600 96.800 ;
        RECT 192.600 96.200 193.000 99.900 ;
        RECT 194.200 96.200 194.600 99.900 ;
        RECT 192.600 95.900 194.600 96.200 ;
        RECT 195.000 95.900 195.400 99.900 ;
        RECT 196.200 96.800 196.600 97.200 ;
        RECT 196.200 96.200 196.500 96.800 ;
        RECT 196.900 96.200 197.300 99.900 ;
        RECT 195.800 95.900 196.500 96.200 ;
        RECT 196.800 95.900 197.300 96.200 ;
        RECT 199.000 96.200 199.400 99.900 ;
        RECT 200.600 96.200 201.000 99.900 ;
        RECT 199.000 95.900 201.000 96.200 ;
        RECT 201.400 95.900 201.800 99.900 ;
        RECT 202.600 96.800 203.000 97.200 ;
        RECT 202.600 96.200 202.900 96.800 ;
        RECT 203.300 96.200 203.700 99.900 ;
        RECT 202.200 95.900 202.900 96.200 ;
        RECT 203.200 95.900 203.700 96.200 ;
        RECT 193.000 95.200 193.400 95.400 ;
        RECT 195.000 95.200 195.300 95.900 ;
        RECT 195.800 95.800 196.200 95.900 ;
        RECT 191.800 95.100 192.200 95.200 ;
        RECT 192.600 95.100 193.400 95.200 ;
        RECT 191.800 94.900 193.400 95.100 ;
        RECT 194.200 95.100 195.400 95.200 ;
        RECT 195.800 95.100 196.200 95.200 ;
        RECT 194.200 94.900 196.200 95.100 ;
        RECT 191.800 94.800 193.000 94.900 ;
        RECT 191.800 94.100 192.200 94.200 ;
        RECT 193.400 94.100 193.800 94.600 ;
        RECT 191.800 93.800 193.800 94.100 ;
        RECT 194.200 93.100 194.500 94.900 ;
        RECT 195.000 94.800 196.200 94.900 ;
        RECT 196.800 94.200 197.100 95.900 ;
        RECT 199.400 95.200 199.800 95.400 ;
        RECT 201.400 95.200 201.700 95.900 ;
        RECT 202.200 95.800 202.600 95.900 ;
        RECT 197.400 95.100 197.800 95.200 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 197.400 94.800 198.600 95.100 ;
        RECT 199.000 94.900 199.800 95.200 ;
        RECT 200.600 95.100 201.800 95.200 ;
        RECT 202.200 95.100 202.600 95.200 ;
        RECT 200.600 94.900 202.600 95.100 ;
        RECT 199.000 94.800 199.400 94.900 ;
        RECT 197.400 94.400 197.800 94.800 ;
        RECT 195.800 93.800 197.100 94.200 ;
        RECT 198.200 94.100 198.600 94.200 ;
        RECT 199.000 94.100 199.300 94.800 ;
        RECT 197.800 93.800 199.300 94.100 ;
        RECT 199.800 93.800 200.200 94.600 ;
        RECT 195.000 93.100 195.400 93.200 ;
        RECT 195.900 93.100 196.200 93.800 ;
        RECT 197.800 93.600 198.200 93.800 ;
        RECT 196.700 93.100 198.500 93.300 ;
        RECT 200.600 93.100 200.900 94.900 ;
        RECT 201.400 94.800 202.600 94.900 ;
        RECT 203.200 94.200 203.500 95.900 ;
        RECT 205.400 95.700 205.800 99.900 ;
        RECT 207.600 98.200 208.000 99.900 ;
        RECT 207.000 97.900 208.000 98.200 ;
        RECT 209.800 97.900 210.200 99.900 ;
        RECT 211.900 97.900 212.500 99.900 ;
        RECT 207.000 97.500 207.400 97.900 ;
        RECT 209.800 97.600 210.100 97.900 ;
        RECT 208.700 97.300 210.500 97.600 ;
        RECT 211.800 97.500 212.200 97.900 ;
        RECT 208.700 97.200 209.100 97.300 ;
        RECT 210.100 97.200 210.500 97.300 ;
        RECT 207.000 96.500 207.400 96.600 ;
        RECT 209.300 96.500 209.700 96.600 ;
        RECT 207.000 96.200 209.700 96.500 ;
        RECT 210.000 96.500 211.100 96.800 ;
        RECT 210.000 95.900 210.300 96.500 ;
        RECT 210.700 96.400 211.100 96.500 ;
        RECT 211.900 96.600 212.600 97.000 ;
        RECT 211.900 96.100 212.200 96.600 ;
        RECT 207.900 95.700 210.300 95.900 ;
        RECT 205.400 95.600 210.300 95.700 ;
        RECT 211.000 95.800 212.200 96.100 ;
        RECT 205.400 95.500 208.300 95.600 ;
        RECT 205.400 95.400 208.200 95.500 ;
        RECT 211.000 95.200 211.300 95.800 ;
        RECT 214.200 95.600 214.600 99.900 ;
        RECT 212.500 95.300 214.600 95.600 ;
        RECT 215.000 95.700 215.400 99.900 ;
        RECT 217.200 98.200 217.600 99.900 ;
        RECT 216.600 97.900 217.600 98.200 ;
        RECT 219.400 97.900 219.800 99.900 ;
        RECT 221.500 97.900 222.100 99.900 ;
        RECT 216.600 97.500 217.000 97.900 ;
        RECT 219.400 97.600 219.700 97.900 ;
        RECT 218.300 97.300 220.100 97.600 ;
        RECT 221.400 97.500 221.800 97.900 ;
        RECT 218.300 97.200 218.700 97.300 ;
        RECT 219.700 97.200 220.100 97.300 ;
        RECT 221.900 97.000 222.600 97.200 ;
        RECT 221.500 96.800 222.600 97.000 ;
        RECT 216.600 96.500 217.000 96.600 ;
        RECT 218.900 96.500 219.300 96.600 ;
        RECT 216.600 96.200 219.300 96.500 ;
        RECT 219.600 96.500 220.700 96.800 ;
        RECT 219.600 95.900 219.900 96.500 ;
        RECT 220.300 96.400 220.700 96.500 ;
        RECT 221.500 96.600 222.200 96.800 ;
        RECT 221.500 96.100 221.800 96.600 ;
        RECT 217.500 95.700 219.900 95.900 ;
        RECT 215.000 95.600 219.900 95.700 ;
        RECT 220.600 95.800 221.800 96.100 ;
        RECT 215.000 95.500 217.900 95.600 ;
        RECT 215.000 95.400 217.800 95.500 ;
        RECT 212.500 95.200 212.900 95.300 ;
        RECT 203.800 94.400 204.200 95.200 ;
        RECT 208.600 95.100 209.000 95.200 ;
        RECT 206.500 94.800 209.000 95.100 ;
        RECT 211.000 94.800 211.400 95.200 ;
        RECT 213.300 94.900 213.700 95.000 ;
        RECT 206.500 94.700 206.900 94.800 ;
        RECT 207.800 94.700 208.200 94.800 ;
        RECT 207.300 94.200 207.700 94.300 ;
        RECT 211.000 94.200 211.300 94.800 ;
        RECT 211.800 94.600 213.700 94.900 ;
        RECT 211.800 94.500 212.200 94.600 ;
        RECT 202.200 93.800 203.500 94.200 ;
        RECT 204.600 94.100 205.000 94.200 ;
        RECT 204.200 93.800 205.000 94.100 ;
        RECT 205.800 93.900 211.300 94.200 ;
        RECT 205.800 93.800 206.600 93.900 ;
        RECT 201.400 93.100 201.800 93.200 ;
        RECT 202.300 93.100 202.600 93.800 ;
        RECT 204.200 93.600 204.600 93.800 ;
        RECT 203.100 93.100 204.900 93.300 ;
        RECT 189.400 92.800 190.300 93.100 ;
        RECT 189.900 92.200 190.300 92.800 ;
        RECT 189.400 91.800 190.300 92.200 ;
        RECT 189.900 91.100 190.300 91.800 ;
        RECT 194.200 91.100 194.600 93.100 ;
        RECT 195.000 92.800 196.200 93.100 ;
        RECT 194.900 92.400 195.300 92.800 ;
        RECT 195.800 91.100 196.200 92.800 ;
        RECT 196.600 93.000 198.600 93.100 ;
        RECT 196.600 91.100 197.000 93.000 ;
        RECT 198.200 91.100 198.600 93.000 ;
        RECT 200.600 91.100 201.000 93.100 ;
        RECT 201.400 92.800 202.600 93.100 ;
        RECT 201.300 92.400 201.700 92.800 ;
        RECT 202.200 91.100 202.600 92.800 ;
        RECT 203.000 93.000 205.000 93.100 ;
        RECT 203.000 91.100 203.400 93.000 ;
        RECT 204.600 91.100 205.000 93.000 ;
        RECT 205.400 91.100 205.800 93.500 ;
        RECT 207.900 92.800 208.200 93.900 ;
        RECT 210.700 93.800 211.100 93.900 ;
        RECT 214.200 93.600 214.600 95.300 ;
        RECT 220.600 95.200 220.900 95.800 ;
        RECT 223.800 95.600 224.200 99.900 ;
        RECT 224.600 96.200 225.000 99.900 ;
        RECT 227.000 96.200 227.400 99.900 ;
        RECT 224.600 95.900 225.700 96.200 ;
        RECT 227.000 95.900 228.100 96.200 ;
        RECT 222.100 95.300 224.200 95.600 ;
        RECT 222.100 95.200 222.500 95.300 ;
        RECT 218.200 95.100 218.600 95.200 ;
        RECT 216.100 94.800 218.600 95.100 ;
        RECT 220.600 94.800 221.000 95.200 ;
        RECT 223.800 95.100 224.200 95.300 ;
        RECT 225.400 95.600 225.700 95.900 ;
        RECT 227.800 95.600 228.100 95.900 ;
        RECT 225.400 95.200 226.000 95.600 ;
        RECT 227.800 95.200 228.400 95.600 ;
        RECT 224.600 95.100 225.000 95.200 ;
        RECT 222.900 94.900 223.300 95.000 ;
        RECT 216.100 94.700 216.500 94.800 ;
        RECT 217.400 94.700 217.800 94.800 ;
        RECT 216.900 94.200 217.300 94.300 ;
        RECT 220.600 94.200 220.900 94.800 ;
        RECT 221.400 94.600 223.300 94.900 ;
        RECT 223.800 94.800 225.000 95.100 ;
        RECT 221.400 94.500 221.800 94.600 ;
        RECT 215.400 93.900 220.900 94.200 ;
        RECT 215.400 93.800 216.200 93.900 ;
        RECT 212.700 93.300 214.600 93.600 ;
        RECT 212.700 93.200 213.100 93.300 ;
        RECT 207.000 92.100 207.400 92.500 ;
        RECT 207.800 92.400 208.200 92.800 ;
        RECT 208.700 92.700 209.100 92.800 ;
        RECT 208.700 92.400 210.100 92.700 ;
        RECT 209.800 92.100 210.100 92.400 ;
        RECT 211.800 92.100 212.200 92.500 ;
        RECT 207.000 91.800 208.000 92.100 ;
        RECT 207.600 91.100 208.000 91.800 ;
        RECT 209.800 91.100 210.200 92.100 ;
        RECT 211.800 91.800 212.500 92.100 ;
        RECT 211.900 91.100 212.500 91.800 ;
        RECT 214.200 91.100 214.600 93.300 ;
        RECT 215.000 91.100 215.400 93.500 ;
        RECT 217.500 92.800 217.800 93.900 ;
        RECT 220.300 93.800 220.700 93.900 ;
        RECT 223.800 93.600 224.200 94.800 ;
        RECT 224.600 94.400 225.000 94.800 ;
        RECT 225.400 93.700 225.700 95.200 ;
        RECT 227.000 94.400 227.400 95.200 ;
        RECT 227.800 93.700 228.100 95.200 ;
        RECT 222.300 93.300 224.200 93.600 ;
        RECT 222.300 93.200 222.700 93.300 ;
        RECT 216.600 92.100 217.000 92.500 ;
        RECT 217.400 92.400 217.800 92.800 ;
        RECT 218.300 92.700 218.700 92.800 ;
        RECT 218.300 92.400 219.700 92.700 ;
        RECT 219.400 92.100 219.700 92.400 ;
        RECT 221.400 92.100 221.800 92.500 ;
        RECT 216.600 91.800 217.600 92.100 ;
        RECT 217.200 91.100 217.600 91.800 ;
        RECT 219.400 91.100 219.800 92.100 ;
        RECT 221.400 91.800 222.100 92.100 ;
        RECT 221.500 91.100 222.100 91.800 ;
        RECT 223.800 91.100 224.200 93.300 ;
        RECT 224.600 93.400 225.700 93.700 ;
        RECT 227.000 93.400 228.100 93.700 ;
        RECT 224.600 91.100 225.000 93.400 ;
        RECT 227.000 91.100 227.400 93.400 ;
        RECT 0.600 87.500 1.000 89.900 ;
        RECT 2.800 89.200 3.200 89.900 ;
        RECT 2.200 88.900 3.200 89.200 ;
        RECT 5.000 88.900 5.400 89.900 ;
        RECT 7.100 89.200 7.700 89.900 ;
        RECT 7.000 88.900 7.700 89.200 ;
        RECT 2.200 88.500 2.600 88.900 ;
        RECT 5.000 88.600 5.300 88.900 ;
        RECT 3.000 88.200 3.400 88.600 ;
        RECT 3.900 88.300 5.300 88.600 ;
        RECT 7.000 88.500 7.400 88.900 ;
        RECT 3.900 88.200 4.300 88.300 ;
        RECT 1.000 87.100 1.800 87.200 ;
        RECT 3.100 87.100 3.400 88.200 ;
        RECT 7.900 87.700 8.300 87.800 ;
        RECT 9.400 87.700 9.800 89.900 ;
        RECT 10.200 87.900 10.600 89.900 ;
        RECT 11.000 88.000 11.400 89.900 ;
        RECT 12.600 88.000 13.000 89.900 ;
        RECT 11.000 87.900 13.000 88.000 ;
        RECT 13.400 87.900 13.800 89.900 ;
        RECT 14.200 88.000 14.600 89.900 ;
        RECT 15.800 88.000 16.200 89.900 ;
        RECT 14.200 87.900 16.200 88.000 ;
        RECT 16.600 88.000 17.000 89.900 ;
        RECT 18.200 88.000 18.600 89.900 ;
        RECT 16.600 87.900 18.600 88.000 ;
        RECT 19.000 87.900 19.400 89.900 ;
        RECT 19.800 87.900 20.200 89.900 ;
        RECT 20.600 88.000 21.000 89.900 ;
        RECT 22.200 88.000 22.600 89.900 ;
        RECT 20.600 87.900 22.600 88.000 ;
        RECT 23.000 88.000 23.400 89.900 ;
        RECT 24.600 88.000 25.000 89.900 ;
        RECT 23.000 87.900 25.000 88.000 ;
        RECT 25.400 87.900 25.800 89.900 ;
        RECT 26.200 88.000 26.600 89.900 ;
        RECT 27.800 88.000 28.200 89.900 ;
        RECT 26.200 87.900 28.200 88.000 ;
        RECT 28.600 87.900 29.000 89.900 ;
        RECT 7.900 87.400 9.800 87.700 ;
        RECT 4.600 87.100 5.000 87.200 ;
        RECT 5.900 87.100 6.300 87.200 ;
        RECT 1.000 86.800 6.500 87.100 ;
        RECT 2.500 86.700 2.900 86.800 ;
        RECT 1.700 86.200 2.100 86.300 ;
        RECT 6.200 86.200 6.500 86.800 ;
        RECT 7.000 86.400 7.400 86.500 ;
        RECT 1.700 86.100 4.200 86.200 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 1.700 85.900 5.000 86.100 ;
        RECT 3.800 85.800 5.000 85.900 ;
        RECT 6.200 85.800 6.600 86.200 ;
        RECT 7.000 86.100 8.900 86.400 ;
        RECT 8.500 86.000 8.900 86.100 ;
        RECT 0.600 85.500 3.400 85.600 ;
        RECT 0.600 85.400 3.500 85.500 ;
        RECT 0.600 85.300 5.500 85.400 ;
        RECT 0.600 81.100 1.000 85.300 ;
        RECT 3.100 85.100 5.500 85.300 ;
        RECT 2.200 84.500 4.900 84.800 ;
        RECT 2.200 84.400 2.600 84.500 ;
        RECT 4.500 84.400 4.900 84.500 ;
        RECT 5.200 84.500 5.500 85.100 ;
        RECT 6.200 85.200 6.500 85.800 ;
        RECT 7.700 85.700 8.100 85.800 ;
        RECT 9.400 85.700 9.800 87.400 ;
        RECT 10.300 87.200 10.600 87.900 ;
        RECT 11.100 87.700 12.900 87.900 ;
        RECT 12.200 87.200 12.600 87.400 ;
        RECT 13.500 87.200 13.800 87.900 ;
        RECT 14.300 87.700 16.100 87.900 ;
        RECT 16.700 87.700 18.500 87.900 ;
        RECT 15.400 87.200 15.800 87.400 ;
        RECT 17.000 87.200 17.400 87.400 ;
        RECT 19.000 87.200 19.300 87.900 ;
        RECT 19.900 87.200 20.200 87.900 ;
        RECT 20.700 87.700 22.500 87.900 ;
        RECT 23.100 87.700 24.900 87.900 ;
        RECT 21.800 87.200 22.200 87.400 ;
        RECT 23.400 87.200 23.800 87.400 ;
        RECT 25.400 87.200 25.700 87.900 ;
        RECT 26.300 87.700 28.100 87.900 ;
        RECT 26.600 87.200 27.000 87.400 ;
        RECT 28.600 87.200 28.900 87.900 ;
        RECT 29.400 87.500 29.800 89.900 ;
        RECT 31.600 89.200 32.000 89.900 ;
        RECT 31.000 88.900 32.000 89.200 ;
        RECT 33.800 88.900 34.200 89.900 ;
        RECT 35.900 89.200 36.500 89.900 ;
        RECT 35.800 88.900 36.500 89.200 ;
        RECT 31.000 88.500 31.400 88.900 ;
        RECT 33.800 88.600 34.100 88.900 ;
        RECT 31.800 88.200 32.200 88.600 ;
        RECT 32.700 88.300 34.100 88.600 ;
        RECT 35.800 88.500 36.200 88.900 ;
        RECT 32.700 88.200 33.100 88.300 ;
        RECT 10.200 86.800 11.500 87.200 ;
        RECT 12.200 86.900 13.000 87.200 ;
        RECT 12.600 86.800 13.000 86.900 ;
        RECT 13.400 86.800 14.700 87.200 ;
        RECT 15.400 87.100 16.200 87.200 ;
        RECT 16.600 87.100 17.400 87.200 ;
        RECT 15.400 86.900 17.400 87.100 ;
        RECT 15.800 86.800 17.000 86.900 ;
        RECT 18.100 86.800 19.400 87.200 ;
        RECT 19.800 86.800 21.100 87.200 ;
        RECT 21.800 87.100 22.600 87.200 ;
        RECT 23.000 87.100 23.800 87.200 ;
        RECT 21.800 86.900 23.800 87.100 ;
        RECT 22.200 86.800 23.400 86.900 ;
        RECT 24.500 86.800 25.800 87.200 ;
        RECT 26.200 86.900 27.000 87.200 ;
        RECT 26.200 86.800 26.600 86.900 ;
        RECT 27.700 86.800 29.000 87.200 ;
        RECT 29.800 87.100 30.600 87.200 ;
        RECT 31.900 87.100 32.200 88.200 ;
        RECT 36.700 87.700 37.100 87.800 ;
        RECT 38.200 87.700 38.600 89.900 ;
        RECT 41.900 88.200 42.300 89.900 ;
        RECT 36.700 87.400 38.600 87.700 ;
        RECT 41.400 87.800 42.500 88.200 ;
        RECT 34.700 87.100 35.100 87.200 ;
        RECT 29.800 86.800 35.300 87.100 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 11.200 86.100 11.500 86.800 ;
        RECT 10.200 85.800 11.500 86.100 ;
        RECT 11.800 86.100 12.200 86.600 ;
        RECT 14.400 86.200 14.700 86.800 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 11.800 85.800 13.000 86.100 ;
        RECT 14.200 85.800 14.700 86.200 ;
        RECT 15.000 86.100 15.400 86.600 ;
        RECT 17.400 86.100 17.800 86.600 ;
        RECT 15.000 85.800 17.800 86.100 ;
        RECT 18.100 86.100 18.400 86.800 ;
        RECT 18.100 85.800 20.100 86.100 ;
        RECT 7.700 85.400 9.800 85.700 ;
        RECT 6.200 84.900 7.400 85.200 ;
        RECT 5.900 84.500 6.300 84.600 ;
        RECT 5.200 84.200 6.300 84.500 ;
        RECT 7.100 84.400 7.400 84.900 ;
        RECT 7.100 84.000 7.800 84.400 ;
        RECT 3.900 83.700 4.300 83.800 ;
        RECT 5.300 83.700 5.700 83.800 ;
        RECT 2.200 83.100 2.600 83.500 ;
        RECT 3.900 83.400 5.700 83.700 ;
        RECT 5.000 83.100 5.300 83.400 ;
        RECT 7.000 83.100 7.400 83.500 ;
        RECT 2.200 82.800 3.200 83.100 ;
        RECT 2.800 81.100 3.200 82.800 ;
        RECT 5.000 81.100 5.400 83.100 ;
        RECT 7.100 81.100 7.700 83.100 ;
        RECT 9.400 81.100 9.800 85.400 ;
        RECT 10.200 85.100 10.600 85.200 ;
        RECT 11.200 85.100 11.500 85.800 ;
        RECT 13.400 85.100 13.800 85.200 ;
        RECT 14.400 85.100 14.700 85.800 ;
        RECT 18.100 85.100 18.400 85.800 ;
        RECT 19.800 85.200 20.100 85.800 ;
        RECT 19.000 85.100 19.400 85.200 ;
        RECT 10.200 84.800 10.900 85.100 ;
        RECT 11.200 84.800 11.700 85.100 ;
        RECT 13.400 84.800 14.100 85.100 ;
        RECT 14.400 84.800 14.900 85.100 ;
        RECT 10.600 84.200 10.900 84.800 ;
        RECT 10.600 83.800 11.000 84.200 ;
        RECT 11.300 81.100 11.700 84.800 ;
        RECT 13.800 84.200 14.100 84.800 ;
        RECT 13.800 83.800 14.200 84.200 ;
        RECT 14.500 81.100 14.900 84.800 ;
        RECT 17.900 84.800 18.400 85.100 ;
        RECT 18.700 84.800 19.400 85.100 ;
        RECT 19.800 85.100 20.200 85.200 ;
        RECT 20.800 85.100 21.100 86.800 ;
        RECT 21.400 85.800 21.800 86.600 ;
        RECT 23.800 85.800 24.200 86.600 ;
        RECT 24.500 86.100 24.800 86.800 ;
        RECT 25.400 86.100 25.800 86.200 ;
        RECT 24.500 85.800 25.800 86.100 ;
        RECT 27.000 85.800 27.400 86.600 ;
        RECT 24.500 85.100 24.800 85.800 ;
        RECT 27.700 85.200 28.000 86.800 ;
        RECT 31.300 86.700 31.700 86.800 ;
        RECT 30.500 86.200 30.900 86.300 ;
        RECT 31.800 86.200 32.200 86.300 ;
        RECT 30.500 85.900 33.000 86.200 ;
        RECT 32.600 85.800 33.000 85.900 ;
        RECT 29.400 85.500 32.200 85.600 ;
        RECT 29.400 85.400 32.300 85.500 ;
        RECT 29.400 85.300 34.300 85.400 ;
        RECT 25.400 85.100 25.800 85.200 ;
        RECT 19.800 84.800 20.500 85.100 ;
        RECT 20.800 84.800 21.300 85.100 ;
        RECT 17.900 81.100 18.300 84.800 ;
        RECT 18.700 84.200 19.000 84.800 ;
        RECT 20.200 84.200 20.500 84.800 ;
        RECT 18.600 83.800 19.400 84.200 ;
        RECT 20.200 83.800 20.600 84.200 ;
        RECT 20.900 82.200 21.300 84.800 ;
        RECT 24.300 84.800 24.800 85.100 ;
        RECT 25.100 84.800 25.800 85.100 ;
        RECT 27.000 84.800 28.000 85.200 ;
        RECT 28.600 85.100 29.000 85.200 ;
        RECT 28.300 84.800 29.000 85.100 ;
        RECT 20.900 81.800 21.800 82.200 ;
        RECT 20.900 81.100 21.300 81.800 ;
        RECT 24.300 81.100 24.700 84.800 ;
        RECT 25.100 84.200 25.400 84.800 ;
        RECT 25.000 83.800 25.400 84.200 ;
        RECT 27.500 81.100 27.900 84.800 ;
        RECT 28.300 84.200 28.600 84.800 ;
        RECT 28.200 83.800 28.600 84.200 ;
        RECT 29.400 81.100 29.800 85.300 ;
        RECT 31.900 85.100 34.300 85.300 ;
        RECT 31.000 84.500 33.700 84.800 ;
        RECT 31.000 84.400 31.400 84.500 ;
        RECT 33.300 84.400 33.700 84.500 ;
        RECT 34.000 84.500 34.300 85.100 ;
        RECT 35.000 85.200 35.300 86.800 ;
        RECT 35.800 86.400 36.200 86.500 ;
        RECT 35.800 86.100 37.700 86.400 ;
        RECT 37.300 86.000 37.700 86.100 ;
        RECT 36.500 85.700 36.900 85.800 ;
        RECT 38.200 85.700 38.600 87.400 ;
        RECT 40.600 86.800 41.000 87.600 ;
        RECT 36.500 85.400 38.600 85.700 ;
        RECT 35.000 84.900 36.200 85.200 ;
        RECT 34.700 84.500 35.100 84.600 ;
        RECT 34.000 84.200 35.100 84.500 ;
        RECT 35.900 84.400 36.200 84.900 ;
        RECT 35.900 84.000 36.600 84.400 ;
        RECT 32.700 83.700 33.100 83.800 ;
        RECT 34.100 83.700 34.500 83.800 ;
        RECT 31.000 83.100 31.400 83.500 ;
        RECT 32.700 83.400 34.500 83.700 ;
        RECT 33.800 83.100 34.100 83.400 ;
        RECT 35.800 83.100 36.200 83.500 ;
        RECT 31.000 82.800 32.000 83.100 ;
        RECT 31.600 81.100 32.000 82.800 ;
        RECT 33.800 81.100 34.200 83.100 ;
        RECT 35.900 81.100 36.500 83.100 ;
        RECT 38.200 81.100 38.600 85.400 ;
        RECT 41.400 81.100 41.800 87.800 ;
        RECT 42.200 87.200 42.500 87.800 ;
        RECT 43.000 87.500 43.400 89.900 ;
        RECT 45.200 89.200 45.600 89.900 ;
        RECT 44.600 88.900 45.600 89.200 ;
        RECT 47.400 88.900 47.800 89.900 ;
        RECT 49.500 89.200 50.100 89.900 ;
        RECT 49.400 88.900 50.100 89.200 ;
        RECT 44.600 88.500 45.000 88.900 ;
        RECT 47.400 88.600 47.700 88.900 ;
        RECT 45.400 88.200 45.800 88.600 ;
        RECT 46.300 88.300 47.700 88.600 ;
        RECT 49.400 88.500 49.800 88.900 ;
        RECT 46.300 88.200 46.700 88.300 ;
        RECT 42.200 86.800 42.600 87.200 ;
        RECT 43.400 87.100 44.200 87.200 ;
        RECT 45.500 87.100 45.800 88.200 ;
        RECT 50.300 87.700 50.700 87.800 ;
        RECT 51.800 87.700 52.200 89.900 ;
        RECT 52.600 88.000 53.000 89.900 ;
        RECT 54.200 88.000 54.600 89.900 ;
        RECT 52.600 87.900 54.600 88.000 ;
        RECT 55.000 87.900 55.400 89.900 ;
        RECT 56.100 88.200 56.500 89.900 ;
        RECT 56.100 87.900 57.000 88.200 ;
        RECT 52.700 87.700 54.500 87.900 ;
        RECT 50.300 87.400 52.200 87.700 ;
        RECT 48.300 87.100 49.000 87.200 ;
        RECT 43.400 86.800 49.000 87.100 ;
        RECT 44.900 86.700 45.300 86.800 ;
        RECT 44.100 86.200 44.500 86.300 ;
        RECT 44.100 85.900 46.600 86.200 ;
        RECT 46.200 85.800 46.600 85.900 ;
        RECT 43.000 85.500 45.800 85.600 ;
        RECT 43.000 85.400 45.900 85.500 ;
        RECT 43.000 85.300 47.900 85.400 ;
        RECT 42.200 84.400 42.600 85.200 ;
        RECT 43.000 81.100 43.400 85.300 ;
        RECT 45.500 85.100 47.900 85.300 ;
        RECT 44.600 84.500 47.300 84.800 ;
        RECT 44.600 84.400 45.000 84.500 ;
        RECT 46.900 84.400 47.300 84.500 ;
        RECT 47.600 84.500 47.900 85.100 ;
        RECT 48.600 85.200 48.900 86.800 ;
        RECT 49.400 86.400 49.800 86.500 ;
        RECT 49.400 86.100 51.300 86.400 ;
        RECT 50.900 86.000 51.300 86.100 ;
        RECT 50.100 85.700 50.500 85.800 ;
        RECT 51.800 85.700 52.200 87.400 ;
        RECT 53.000 87.200 53.400 87.400 ;
        RECT 55.000 87.200 55.300 87.900 ;
        RECT 52.600 86.900 53.400 87.200 ;
        RECT 52.600 86.800 53.000 86.900 ;
        RECT 54.100 86.800 55.400 87.200 ;
        RECT 53.400 85.800 53.800 86.600 ;
        RECT 54.100 86.200 54.400 86.800 ;
        RECT 54.100 85.800 54.600 86.200 ;
        RECT 56.600 86.100 57.000 87.900 ;
        RECT 58.200 87.800 58.600 88.600 ;
        RECT 57.400 87.100 57.800 87.600 ;
        RECT 58.200 87.100 58.500 87.800 ;
        RECT 57.400 86.800 58.500 87.100 ;
        RECT 55.000 85.800 57.000 86.100 ;
        RECT 50.100 85.400 52.200 85.700 ;
        RECT 48.600 84.900 49.800 85.200 ;
        RECT 48.300 84.500 48.700 84.600 ;
        RECT 47.600 84.200 48.700 84.500 ;
        RECT 49.500 84.400 49.800 84.900 ;
        RECT 49.500 84.000 50.200 84.400 ;
        RECT 46.300 83.700 46.700 83.800 ;
        RECT 47.700 83.700 48.100 83.800 ;
        RECT 44.600 83.100 45.000 83.500 ;
        RECT 46.300 83.400 48.100 83.700 ;
        RECT 47.400 83.100 47.700 83.400 ;
        RECT 49.400 83.100 49.800 83.500 ;
        RECT 44.600 82.800 45.600 83.100 ;
        RECT 45.200 81.100 45.600 82.800 ;
        RECT 47.400 81.100 47.800 83.100 ;
        RECT 49.500 81.100 50.100 83.100 ;
        RECT 51.800 81.100 52.200 85.400 ;
        RECT 54.100 85.100 54.400 85.800 ;
        RECT 55.000 85.200 55.300 85.800 ;
        RECT 55.000 85.100 55.400 85.200 ;
        RECT 53.900 84.800 54.400 85.100 ;
        RECT 54.700 84.800 55.400 85.100 ;
        RECT 53.900 81.100 54.300 84.800 ;
        RECT 54.700 84.200 55.000 84.800 ;
        RECT 55.800 84.400 56.200 85.200 ;
        RECT 54.600 83.800 55.000 84.200 ;
        RECT 56.600 81.100 57.000 85.800 ;
        RECT 59.000 81.100 59.400 89.900 ;
        RECT 59.800 88.000 60.200 89.900 ;
        RECT 61.400 89.600 63.400 89.900 ;
        RECT 61.400 88.000 61.800 89.600 ;
        RECT 59.800 87.900 61.800 88.000 ;
        RECT 62.200 87.900 62.600 89.300 ;
        RECT 63.000 87.900 63.400 89.600 ;
        RECT 59.900 87.700 61.700 87.900 ;
        RECT 60.200 87.200 60.600 87.400 ;
        RECT 62.300 87.200 62.600 87.900 ;
        RECT 59.800 86.900 60.600 87.200 ;
        RECT 61.400 86.900 62.600 87.200 ;
        RECT 59.800 86.800 60.200 86.900 ;
        RECT 61.400 86.800 61.800 86.900 ;
        RECT 60.600 85.800 61.000 86.600 ;
        RECT 61.400 85.100 61.700 86.800 ;
        RECT 62.200 85.800 62.600 86.600 ;
        RECT 63.000 86.400 63.400 87.200 ;
        RECT 63.800 86.100 64.200 89.900 ;
        RECT 64.600 87.800 65.000 88.600 ;
        RECT 65.400 88.000 65.800 89.900 ;
        RECT 67.000 88.000 67.400 89.900 ;
        RECT 65.400 87.900 67.400 88.000 ;
        RECT 67.800 87.900 68.200 89.900 ;
        RECT 65.500 87.700 67.300 87.900 ;
        RECT 65.800 87.200 66.200 87.400 ;
        RECT 67.800 87.200 68.100 87.900 ;
        RECT 69.400 87.600 69.800 89.900 ;
        RECT 71.000 87.600 71.400 89.900 ;
        RECT 72.600 87.600 73.000 89.900 ;
        RECT 74.200 87.600 74.600 89.900 ;
        RECT 68.600 87.200 69.800 87.600 ;
        RECT 70.300 87.200 71.400 87.600 ;
        RECT 71.900 87.200 73.000 87.600 ;
        RECT 73.700 87.200 74.600 87.600 ;
        RECT 65.400 86.900 66.200 87.200 ;
        RECT 65.400 86.800 65.800 86.900 ;
        RECT 66.900 86.800 68.200 87.200 ;
        RECT 64.600 86.100 65.000 86.200 ;
        RECT 63.800 85.800 65.000 86.100 ;
        RECT 66.200 85.800 66.600 86.600 ;
        RECT 61.100 82.200 62.100 85.100 ;
        RECT 61.100 81.800 62.600 82.200 ;
        RECT 61.100 81.100 62.100 81.800 ;
        RECT 63.800 81.100 64.200 85.800 ;
        RECT 66.900 85.100 67.200 86.800 ;
        RECT 67.800 86.200 68.100 86.800 ;
        RECT 67.800 85.800 68.200 86.200 ;
        RECT 68.600 85.800 69.000 87.200 ;
        RECT 70.300 86.900 70.700 87.200 ;
        RECT 71.900 86.900 72.300 87.200 ;
        RECT 73.700 86.900 74.100 87.200 ;
        RECT 77.600 87.100 78.000 89.900 ;
        RECT 79.000 87.700 79.400 89.900 ;
        RECT 81.100 89.200 81.700 89.900 ;
        RECT 81.100 88.900 81.800 89.200 ;
        RECT 83.400 88.900 83.800 89.900 ;
        RECT 85.600 89.200 86.000 89.900 ;
        RECT 85.600 88.900 86.600 89.200 ;
        RECT 81.400 88.500 81.800 88.900 ;
        RECT 83.500 88.600 83.800 88.900 ;
        RECT 83.500 88.300 84.900 88.600 ;
        RECT 84.500 88.200 84.900 88.300 ;
        RECT 85.400 87.800 85.800 88.600 ;
        RECT 86.200 88.500 86.600 88.900 ;
        RECT 80.500 87.700 80.900 87.800 ;
        RECT 79.000 87.400 80.900 87.700 ;
        RECT 77.600 86.900 78.500 87.100 ;
        RECT 69.400 86.500 70.700 86.900 ;
        RECT 71.100 86.500 72.300 86.900 ;
        RECT 72.800 86.500 74.100 86.900 ;
        RECT 77.700 86.800 78.500 86.900 ;
        RECT 70.300 85.800 70.700 86.500 ;
        RECT 71.900 85.800 72.300 86.500 ;
        RECT 73.700 85.800 74.100 86.500 ;
        RECT 76.600 85.800 77.400 86.200 ;
        RECT 68.600 85.400 69.800 85.800 ;
        RECT 70.300 85.400 71.400 85.800 ;
        RECT 71.900 85.400 73.000 85.800 ;
        RECT 73.700 85.400 74.600 85.800 ;
        RECT 67.800 85.100 68.200 85.200 ;
        RECT 66.700 84.800 67.200 85.100 ;
        RECT 67.500 84.800 68.200 85.100 ;
        RECT 66.700 81.100 67.100 84.800 ;
        RECT 67.500 84.200 67.800 84.800 ;
        RECT 67.400 83.800 67.800 84.200 ;
        RECT 69.400 81.100 69.800 85.400 ;
        RECT 71.000 81.100 71.400 85.400 ;
        RECT 72.600 81.100 73.000 85.400 ;
        RECT 74.200 81.100 74.600 85.400 ;
        RECT 75.800 84.800 76.200 85.600 ;
        RECT 78.200 85.200 78.500 86.800 ;
        RECT 79.000 85.700 79.400 87.400 ;
        RECT 82.500 87.100 82.900 87.200 ;
        RECT 85.400 87.100 85.700 87.800 ;
        RECT 87.800 87.500 88.200 89.900 ;
        RECT 90.200 88.000 90.600 89.900 ;
        RECT 91.800 88.000 92.200 89.900 ;
        RECT 90.200 87.900 92.200 88.000 ;
        RECT 92.600 87.900 93.000 89.900 ;
        RECT 94.700 88.200 95.100 89.900 ;
        RECT 94.200 87.900 95.100 88.200 ;
        RECT 95.800 88.000 96.200 89.900 ;
        RECT 97.400 88.000 97.800 89.900 ;
        RECT 95.800 87.900 97.800 88.000 ;
        RECT 98.200 87.900 98.600 89.900 ;
        RECT 90.300 87.700 92.100 87.900 ;
        RECT 90.600 87.200 91.000 87.400 ;
        RECT 92.600 87.200 92.900 87.900 ;
        RECT 87.000 87.100 87.800 87.200 ;
        RECT 82.300 86.800 87.800 87.100 ;
        RECT 90.200 86.900 91.000 87.200 ;
        RECT 90.200 86.800 90.600 86.900 ;
        RECT 91.700 86.800 93.000 87.200 ;
        RECT 93.400 86.800 93.800 87.600 ;
        RECT 81.400 86.400 81.800 86.500 ;
        RECT 79.900 86.100 81.800 86.400 ;
        RECT 82.300 86.200 82.600 86.800 ;
        RECT 85.900 86.700 86.300 86.800 ;
        RECT 85.400 86.200 85.800 86.300 ;
        RECT 86.700 86.200 87.100 86.300 ;
        RECT 79.900 86.000 80.300 86.100 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 84.600 85.900 87.100 86.200 ;
        RECT 84.600 85.800 85.000 85.900 ;
        RECT 91.000 85.800 91.400 86.600 ;
        RECT 80.700 85.700 81.100 85.800 ;
        RECT 79.000 85.400 81.100 85.700 ;
        RECT 78.200 84.800 78.600 85.200 ;
        RECT 77.400 83.800 77.800 84.600 ;
        RECT 78.200 83.500 78.500 84.800 ;
        RECT 76.700 83.200 78.500 83.500 ;
        RECT 76.700 83.100 77.000 83.200 ;
        RECT 76.600 81.100 77.000 83.100 ;
        RECT 78.200 83.100 78.500 83.200 ;
        RECT 78.200 81.100 78.600 83.100 ;
        RECT 79.000 81.100 79.400 85.400 ;
        RECT 82.300 85.200 82.600 85.800 ;
        RECT 85.400 85.500 88.200 85.600 ;
        RECT 85.300 85.400 88.200 85.500 ;
        RECT 81.400 84.900 82.600 85.200 ;
        RECT 83.300 85.300 88.200 85.400 ;
        RECT 83.300 85.100 85.700 85.300 ;
        RECT 81.400 84.400 81.700 84.900 ;
        RECT 81.000 84.000 81.700 84.400 ;
        RECT 82.500 84.500 82.900 84.600 ;
        RECT 83.300 84.500 83.600 85.100 ;
        RECT 82.500 84.200 83.600 84.500 ;
        RECT 83.900 84.500 86.600 84.800 ;
        RECT 83.900 84.400 84.300 84.500 ;
        RECT 86.200 84.400 86.600 84.500 ;
        RECT 83.100 83.700 83.500 83.800 ;
        RECT 84.500 83.700 84.900 83.800 ;
        RECT 81.400 83.100 81.800 83.500 ;
        RECT 83.100 83.400 84.900 83.700 ;
        RECT 83.500 83.100 83.800 83.400 ;
        RECT 86.200 83.100 86.600 83.500 ;
        RECT 81.100 81.100 81.700 83.100 ;
        RECT 83.400 81.100 83.800 83.100 ;
        RECT 85.600 82.800 86.600 83.100 ;
        RECT 85.600 81.100 86.000 82.800 ;
        RECT 87.800 81.100 88.200 85.300 ;
        RECT 91.700 85.200 92.000 86.800 ;
        RECT 91.000 84.800 92.000 85.200 ;
        RECT 92.600 85.100 93.000 85.200 ;
        RECT 92.300 84.800 93.000 85.100 ;
        RECT 91.500 81.100 91.900 84.800 ;
        RECT 92.300 84.200 92.600 84.800 ;
        RECT 92.200 83.800 92.600 84.200 ;
        RECT 93.400 84.100 93.800 84.200 ;
        RECT 94.200 84.100 94.600 87.900 ;
        RECT 95.900 87.700 97.700 87.900 ;
        RECT 96.200 87.200 96.600 87.400 ;
        RECT 98.200 87.200 98.500 87.900 ;
        RECT 99.000 87.500 99.400 89.900 ;
        RECT 101.200 89.200 101.600 89.900 ;
        RECT 100.600 88.900 101.600 89.200 ;
        RECT 103.400 88.900 103.800 89.900 ;
        RECT 105.500 89.200 106.100 89.900 ;
        RECT 105.400 88.900 106.100 89.200 ;
        RECT 100.600 88.500 101.000 88.900 ;
        RECT 103.400 88.600 103.700 88.900 ;
        RECT 101.400 88.200 101.800 88.600 ;
        RECT 102.300 88.300 103.700 88.600 ;
        RECT 105.400 88.500 105.800 88.900 ;
        RECT 102.300 88.200 102.700 88.300 ;
        RECT 95.800 86.900 96.600 87.200 ;
        RECT 95.800 86.800 96.200 86.900 ;
        RECT 97.300 86.800 98.600 87.200 ;
        RECT 99.400 87.100 100.200 87.200 ;
        RECT 101.500 87.100 101.800 88.200 ;
        RECT 106.300 87.700 106.700 87.800 ;
        RECT 107.800 87.700 108.200 89.900 ;
        RECT 108.600 88.000 109.000 89.900 ;
        RECT 110.200 88.000 110.600 89.900 ;
        RECT 108.600 87.900 110.600 88.000 ;
        RECT 111.000 87.900 111.400 89.900 ;
        RECT 113.400 87.900 113.800 89.900 ;
        RECT 114.100 88.200 114.500 88.600 ;
        RECT 108.700 87.700 110.500 87.900 ;
        RECT 106.300 87.400 108.200 87.700 ;
        RECT 104.300 87.100 104.700 87.200 ;
        RECT 99.400 86.800 104.900 87.100 ;
        RECT 96.600 85.800 97.000 86.600 ;
        RECT 95.000 84.400 95.400 85.200 ;
        RECT 97.300 85.100 97.600 86.800 ;
        RECT 98.200 86.200 98.500 86.800 ;
        RECT 100.900 86.700 101.300 86.800 ;
        RECT 100.100 86.200 100.500 86.300 ;
        RECT 101.400 86.200 101.800 86.300 ;
        RECT 104.600 86.200 104.900 86.800 ;
        RECT 105.400 86.400 105.800 86.500 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 100.100 85.900 102.600 86.200 ;
        RECT 102.200 85.800 102.600 85.900 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 105.400 86.100 107.300 86.400 ;
        RECT 106.900 86.000 107.300 86.100 ;
        RECT 99.000 85.500 101.800 85.600 ;
        RECT 99.000 85.400 101.900 85.500 ;
        RECT 99.000 85.300 103.900 85.400 ;
        RECT 98.200 85.100 98.600 85.200 ;
        RECT 97.100 84.800 97.600 85.100 ;
        RECT 97.900 84.800 98.600 85.100 ;
        RECT 93.400 83.800 94.600 84.100 ;
        RECT 94.200 81.100 94.600 83.800 ;
        RECT 97.100 81.100 97.500 84.800 ;
        RECT 97.900 84.200 98.200 84.800 ;
        RECT 97.800 83.800 98.200 84.200 ;
        RECT 99.000 81.100 99.400 85.300 ;
        RECT 101.500 85.100 103.900 85.300 ;
        RECT 100.600 84.500 103.300 84.800 ;
        RECT 100.600 84.400 101.000 84.500 ;
        RECT 102.900 84.400 103.300 84.500 ;
        RECT 103.600 84.500 103.900 85.100 ;
        RECT 104.600 85.200 104.900 85.800 ;
        RECT 106.100 85.700 106.500 85.800 ;
        RECT 107.800 85.700 108.200 87.400 ;
        RECT 109.000 87.200 109.400 87.400 ;
        RECT 111.000 87.200 111.300 87.900 ;
        RECT 108.600 86.900 109.400 87.200 ;
        RECT 108.600 86.800 109.000 86.900 ;
        RECT 110.100 86.800 111.400 87.200 ;
        RECT 109.400 85.800 109.800 86.600 ;
        RECT 110.100 86.100 110.400 86.800 ;
        RECT 112.600 86.400 113.000 87.200 ;
        RECT 111.800 86.100 112.200 86.200 ;
        RECT 113.400 86.100 113.700 87.900 ;
        RECT 114.200 87.800 114.600 88.200 ;
        RECT 115.000 88.000 115.400 89.900 ;
        RECT 116.600 88.000 117.000 89.900 ;
        RECT 115.000 87.900 117.000 88.000 ;
        RECT 117.400 87.900 117.800 89.900 ;
        RECT 118.200 88.000 118.600 89.900 ;
        RECT 119.800 88.000 120.200 89.900 ;
        RECT 118.200 87.900 120.200 88.000 ;
        RECT 120.600 87.900 121.000 89.900 ;
        RECT 115.100 87.700 116.900 87.900 ;
        RECT 115.400 87.200 115.800 87.400 ;
        RECT 117.400 87.200 117.700 87.900 ;
        RECT 118.300 87.700 120.100 87.900 ;
        RECT 118.600 87.200 119.000 87.400 ;
        RECT 120.600 87.200 120.900 87.900 ;
        RECT 121.400 87.500 121.800 89.900 ;
        RECT 123.600 89.200 124.000 89.900 ;
        RECT 123.000 88.900 124.000 89.200 ;
        RECT 125.800 88.900 126.200 89.900 ;
        RECT 127.900 89.200 128.500 89.900 ;
        RECT 127.800 88.900 128.500 89.200 ;
        RECT 123.000 88.500 123.400 88.900 ;
        RECT 125.800 88.600 126.100 88.900 ;
        RECT 123.800 88.200 124.200 88.600 ;
        RECT 124.700 88.300 126.100 88.600 ;
        RECT 127.800 88.500 128.200 88.900 ;
        RECT 124.700 88.200 125.100 88.300 ;
        RECT 114.200 87.100 114.600 87.200 ;
        RECT 115.000 87.100 115.800 87.200 ;
        RECT 114.200 86.900 115.800 87.100 ;
        RECT 114.200 86.800 115.400 86.900 ;
        RECT 116.500 86.800 117.800 87.200 ;
        RECT 118.200 86.900 119.000 87.200 ;
        RECT 118.200 86.800 118.600 86.900 ;
        RECT 119.700 86.800 121.000 87.200 ;
        RECT 121.800 87.100 122.600 87.200 ;
        RECT 123.900 87.100 124.200 88.200 ;
        RECT 128.700 87.700 129.100 87.800 ;
        RECT 130.200 87.700 130.600 89.900 ;
        RECT 128.700 87.400 130.600 87.700 ;
        RECT 126.700 87.100 127.100 87.200 ;
        RECT 121.800 86.800 127.300 87.100 ;
        RECT 114.200 86.100 114.600 86.200 ;
        RECT 115.800 86.100 116.200 86.600 ;
        RECT 110.100 85.800 112.600 86.100 ;
        RECT 113.400 85.800 116.200 86.100 ;
        RECT 116.500 86.200 116.800 86.800 ;
        RECT 116.500 85.800 117.000 86.200 ;
        RECT 119.000 85.800 119.400 86.600 ;
        RECT 106.100 85.400 108.200 85.700 ;
        RECT 104.600 84.900 105.800 85.200 ;
        RECT 104.300 84.500 104.700 84.600 ;
        RECT 103.600 84.200 104.700 84.500 ;
        RECT 105.500 84.400 105.800 84.900 ;
        RECT 105.500 84.000 106.200 84.400 ;
        RECT 102.300 83.700 102.700 83.800 ;
        RECT 103.700 83.700 104.100 83.800 ;
        RECT 100.600 83.100 101.000 83.500 ;
        RECT 102.300 83.400 104.100 83.700 ;
        RECT 103.400 83.100 103.700 83.400 ;
        RECT 105.400 83.100 105.800 83.500 ;
        RECT 100.600 82.800 101.600 83.100 ;
        RECT 101.200 81.100 101.600 82.800 ;
        RECT 103.400 81.100 103.800 83.100 ;
        RECT 105.500 81.100 106.100 83.100 ;
        RECT 107.800 81.100 108.200 85.400 ;
        RECT 110.100 85.100 110.400 85.800 ;
        RECT 112.200 85.600 112.600 85.800 ;
        RECT 111.000 85.100 111.400 85.200 ;
        RECT 114.200 85.100 114.500 85.800 ;
        RECT 116.500 85.100 116.800 85.800 ;
        RECT 117.400 85.100 117.800 85.200 ;
        RECT 119.700 85.100 120.000 86.800 ;
        RECT 123.300 86.700 123.700 86.800 ;
        RECT 122.500 86.200 122.900 86.300 ;
        RECT 122.500 85.900 125.000 86.200 ;
        RECT 124.600 85.800 125.000 85.900 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 127.000 86.100 127.300 86.800 ;
        RECT 127.800 86.400 128.200 86.500 ;
        RECT 127.800 86.100 129.700 86.400 ;
        RECT 126.200 85.800 127.300 86.100 ;
        RECT 129.300 86.000 129.700 86.100 ;
        RECT 121.400 85.500 124.200 85.600 ;
        RECT 121.400 85.400 124.300 85.500 ;
        RECT 121.400 85.300 126.300 85.400 ;
        RECT 120.600 85.100 121.000 85.200 ;
        RECT 109.900 84.800 110.400 85.100 ;
        RECT 110.700 84.800 111.400 85.100 ;
        RECT 111.800 84.800 113.800 85.100 ;
        RECT 109.900 81.100 110.300 84.800 ;
        RECT 110.700 84.200 111.000 84.800 ;
        RECT 110.600 83.800 111.000 84.200 ;
        RECT 111.800 81.100 112.200 84.800 ;
        RECT 113.400 81.100 113.800 84.800 ;
        RECT 114.200 81.100 114.600 85.100 ;
        RECT 116.300 84.800 116.800 85.100 ;
        RECT 117.100 84.800 117.800 85.100 ;
        RECT 119.500 84.800 120.000 85.100 ;
        RECT 120.300 84.800 121.000 85.100 ;
        RECT 116.300 81.100 116.700 84.800 ;
        RECT 117.100 84.200 117.400 84.800 ;
        RECT 117.000 83.800 117.400 84.200 ;
        RECT 119.500 81.100 119.900 84.800 ;
        RECT 120.300 84.200 120.600 84.800 ;
        RECT 120.200 83.800 120.600 84.200 ;
        RECT 121.400 81.100 121.800 85.300 ;
        RECT 123.900 85.100 126.300 85.300 ;
        RECT 123.000 84.500 125.700 84.800 ;
        RECT 123.000 84.400 123.400 84.500 ;
        RECT 125.300 84.400 125.700 84.500 ;
        RECT 126.000 84.500 126.300 85.100 ;
        RECT 127.000 85.200 127.300 85.800 ;
        RECT 128.500 85.700 128.900 85.800 ;
        RECT 130.200 85.700 130.600 87.400 ;
        RECT 128.500 85.400 130.600 85.700 ;
        RECT 127.000 84.900 128.200 85.200 ;
        RECT 126.700 84.500 127.100 84.600 ;
        RECT 126.000 84.200 127.100 84.500 ;
        RECT 127.900 84.400 128.200 84.900 ;
        RECT 127.900 84.000 128.600 84.400 ;
        RECT 124.700 83.700 125.100 83.800 ;
        RECT 126.100 83.700 126.500 83.800 ;
        RECT 123.000 83.100 123.400 83.500 ;
        RECT 124.700 83.400 126.500 83.700 ;
        RECT 125.800 83.100 126.100 83.400 ;
        RECT 127.800 83.100 128.200 83.500 ;
        RECT 123.000 82.800 124.000 83.100 ;
        RECT 123.600 81.100 124.000 82.800 ;
        RECT 125.800 81.100 126.200 83.100 ;
        RECT 127.900 81.100 128.500 83.100 ;
        RECT 130.200 81.100 130.600 85.400 ;
        RECT 131.000 87.700 131.400 89.900 ;
        RECT 133.100 89.200 133.700 89.900 ;
        RECT 133.100 88.900 133.800 89.200 ;
        RECT 135.400 88.900 135.800 89.900 ;
        RECT 137.600 89.200 138.000 89.900 ;
        RECT 137.600 88.900 138.600 89.200 ;
        RECT 133.400 88.500 133.800 88.900 ;
        RECT 135.500 88.600 135.800 88.900 ;
        RECT 135.500 88.300 136.900 88.600 ;
        RECT 136.500 88.200 136.900 88.300 ;
        RECT 137.400 88.200 137.800 88.600 ;
        RECT 138.200 88.500 138.600 88.900 ;
        RECT 132.500 87.700 132.900 87.800 ;
        RECT 131.000 87.400 132.900 87.700 ;
        RECT 131.000 85.700 131.400 87.400 ;
        RECT 134.500 87.100 134.900 87.200 ;
        RECT 137.400 87.100 137.700 88.200 ;
        RECT 139.800 87.500 140.200 89.900 ;
        RECT 143.500 88.200 143.900 89.900 ;
        RECT 143.000 87.900 143.900 88.200 ;
        RECT 144.600 87.900 145.000 89.900 ;
        RECT 145.400 88.000 145.800 89.900 ;
        RECT 147.000 88.000 147.400 89.900 ;
        RECT 145.400 87.900 147.400 88.000 ;
        RECT 148.100 89.200 148.500 89.900 ;
        RECT 148.100 88.800 149.000 89.200 ;
        RECT 148.100 88.200 148.500 88.800 ;
        RECT 150.500 88.200 150.900 89.900 ;
        RECT 148.100 87.900 149.000 88.200 ;
        RECT 150.500 87.900 151.400 88.200 ;
        RECT 139.000 87.100 139.800 87.200 ;
        RECT 134.300 86.800 139.800 87.100 ;
        RECT 140.600 87.100 141.000 87.200 ;
        RECT 142.200 87.100 142.600 87.600 ;
        RECT 140.600 86.800 142.600 87.100 ;
        RECT 133.400 86.400 133.800 86.500 ;
        RECT 131.900 86.100 133.800 86.400 ;
        RECT 134.300 86.200 134.600 86.800 ;
        RECT 137.900 86.700 138.300 86.800 ;
        RECT 137.400 86.200 137.800 86.300 ;
        RECT 138.700 86.200 139.100 86.300 ;
        RECT 131.900 86.000 132.300 86.100 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 136.600 85.900 139.100 86.200 ;
        RECT 143.000 86.100 143.400 87.900 ;
        RECT 144.700 87.200 145.000 87.900 ;
        RECT 145.500 87.700 147.300 87.900 ;
        RECT 146.600 87.200 147.000 87.400 ;
        RECT 143.800 87.100 144.200 87.200 ;
        RECT 144.600 87.100 145.900 87.200 ;
        RECT 143.800 86.800 145.900 87.100 ;
        RECT 146.600 86.900 147.400 87.200 ;
        RECT 147.000 86.800 147.400 86.900 ;
        RECT 136.600 85.800 137.000 85.900 ;
        RECT 143.000 85.800 144.900 86.100 ;
        RECT 132.700 85.700 133.100 85.800 ;
        RECT 131.000 85.400 133.100 85.700 ;
        RECT 131.000 81.100 131.400 85.400 ;
        RECT 134.300 85.200 134.600 85.800 ;
        RECT 137.400 85.500 140.200 85.600 ;
        RECT 137.300 85.400 140.200 85.500 ;
        RECT 133.400 84.900 134.600 85.200 ;
        RECT 135.300 85.300 140.200 85.400 ;
        RECT 135.300 85.100 137.700 85.300 ;
        RECT 133.400 84.400 133.700 84.900 ;
        RECT 133.000 84.000 133.700 84.400 ;
        RECT 134.500 84.500 134.900 84.600 ;
        RECT 135.300 84.500 135.600 85.100 ;
        RECT 134.500 84.200 135.600 84.500 ;
        RECT 135.900 84.500 138.600 84.800 ;
        RECT 135.900 84.400 136.300 84.500 ;
        RECT 138.200 84.400 138.600 84.500 ;
        RECT 135.100 83.700 135.500 83.800 ;
        RECT 136.500 83.700 136.900 83.800 ;
        RECT 133.400 83.100 133.800 83.500 ;
        RECT 135.100 83.400 136.900 83.700 ;
        RECT 135.500 83.100 135.800 83.400 ;
        RECT 138.200 83.100 138.600 83.500 ;
        RECT 133.100 81.100 133.700 83.100 ;
        RECT 135.400 81.100 135.800 83.100 ;
        RECT 137.600 82.800 138.600 83.100 ;
        RECT 137.600 81.100 138.000 82.800 ;
        RECT 139.800 81.100 140.200 85.300 ;
        RECT 143.000 81.100 143.400 85.800 ;
        RECT 144.600 85.200 144.900 85.800 ;
        RECT 143.800 84.400 144.200 85.200 ;
        RECT 144.600 85.100 145.000 85.200 ;
        RECT 145.600 85.100 145.900 86.800 ;
        RECT 146.200 85.800 146.600 86.600 ;
        RECT 144.600 84.800 145.300 85.100 ;
        RECT 145.600 84.800 146.100 85.100 ;
        RECT 145.000 84.200 145.300 84.800 ;
        RECT 145.000 83.800 145.400 84.200 ;
        RECT 145.700 81.100 146.100 84.800 ;
        RECT 147.800 84.400 148.200 85.200 ;
        RECT 148.600 81.100 149.000 87.900 ;
        RECT 149.400 86.800 149.800 87.600 ;
        RECT 149.400 85.100 149.800 85.200 ;
        RECT 150.200 85.100 150.600 85.200 ;
        RECT 149.400 84.800 150.600 85.100 ;
        RECT 150.200 84.400 150.600 84.800 ;
        RECT 151.000 81.100 151.400 87.900 ;
        RECT 154.200 87.900 154.600 89.900 ;
        RECT 157.400 87.900 157.800 89.900 ;
        RECT 160.600 87.900 161.000 89.900 ;
        RECT 161.300 88.200 161.700 88.600 ;
        RECT 151.800 86.800 152.200 87.600 ;
        RECT 153.400 86.400 153.800 87.200 ;
        RECT 152.600 86.100 153.000 86.200 ;
        RECT 154.200 86.100 154.500 87.900 ;
        RECT 156.600 86.400 157.000 87.200 ;
        RECT 155.000 86.100 155.400 86.200 ;
        RECT 152.600 85.800 153.400 86.100 ;
        RECT 154.200 85.800 155.400 86.100 ;
        RECT 155.800 86.100 156.200 86.200 ;
        RECT 157.400 86.100 157.700 87.900 ;
        RECT 159.800 86.400 160.200 87.200 ;
        RECT 158.200 86.100 158.600 86.200 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 160.600 86.100 160.900 87.900 ;
        RECT 161.400 87.800 161.800 88.200 ;
        RECT 163.800 87.900 164.200 89.900 ;
        RECT 164.500 88.200 164.900 88.600 ;
        RECT 163.000 86.400 163.400 87.200 ;
        RECT 161.400 86.100 161.800 86.200 ;
        RECT 155.800 85.800 156.600 86.100 ;
        RECT 157.400 85.800 159.800 86.100 ;
        RECT 160.600 85.800 161.800 86.100 ;
        RECT 162.200 86.100 162.600 86.200 ;
        RECT 163.800 86.100 164.100 87.900 ;
        RECT 164.600 87.800 165.000 88.200 ;
        RECT 165.400 87.900 165.800 89.900 ;
        RECT 166.200 88.000 166.600 89.900 ;
        RECT 167.800 88.000 168.200 89.900 ;
        RECT 166.200 87.900 168.200 88.000 ;
        RECT 165.500 87.200 165.800 87.900 ;
        RECT 166.300 87.700 168.100 87.900 ;
        RECT 168.600 87.800 169.000 89.900 ;
        RECT 169.400 88.000 169.800 89.900 ;
        RECT 171.000 88.000 171.400 89.900 ;
        RECT 169.400 87.900 171.400 88.000 ;
        RECT 167.400 87.200 167.800 87.400 ;
        RECT 168.700 87.200 169.000 87.800 ;
        RECT 169.500 87.700 171.300 87.900 ;
        RECT 171.800 87.600 172.200 89.900 ;
        RECT 174.200 87.900 174.600 89.900 ;
        RECT 175.000 88.000 175.400 89.900 ;
        RECT 176.600 88.000 177.000 89.900 ;
        RECT 177.500 88.200 177.900 88.600 ;
        RECT 175.000 87.900 177.000 88.000 ;
        RECT 170.600 87.200 171.000 87.400 ;
        RECT 171.800 87.300 172.900 87.600 ;
        RECT 165.400 86.800 166.700 87.200 ;
        RECT 167.400 86.900 168.200 87.200 ;
        RECT 167.800 86.800 168.200 86.900 ;
        RECT 168.600 86.800 169.900 87.200 ;
        RECT 170.600 86.900 171.400 87.200 ;
        RECT 171.000 86.800 171.400 86.900 ;
        RECT 164.600 86.100 165.000 86.200 ;
        RECT 162.200 85.800 163.000 86.100 ;
        RECT 163.800 85.800 165.000 86.100 ;
        RECT 153.000 85.600 153.400 85.800 ;
        RECT 155.000 85.200 155.300 85.800 ;
        RECT 156.200 85.600 156.600 85.800 ;
        RECT 152.600 84.800 154.600 85.100 ;
        RECT 152.600 81.100 153.000 84.800 ;
        RECT 154.200 81.100 154.600 84.800 ;
        RECT 155.000 81.100 155.400 85.200 ;
        RECT 158.200 85.100 158.500 85.800 ;
        RECT 159.400 85.600 159.800 85.800 ;
        RECT 161.400 85.100 161.700 85.800 ;
        RECT 162.600 85.600 163.000 85.800 ;
        RECT 164.600 85.100 164.900 85.800 ;
        RECT 165.400 85.100 165.800 85.200 ;
        RECT 166.400 85.100 166.700 86.800 ;
        RECT 167.000 85.800 167.400 86.600 ;
        RECT 168.600 85.800 169.000 86.200 ;
        RECT 168.600 85.200 168.900 85.800 ;
        RECT 168.600 85.100 169.000 85.200 ;
        RECT 169.600 85.100 169.900 86.800 ;
        RECT 170.200 85.800 170.600 86.600 ;
        RECT 171.800 85.800 172.200 86.600 ;
        RECT 172.600 85.800 172.900 87.300 ;
        RECT 174.300 87.200 174.600 87.900 ;
        RECT 175.100 87.700 176.900 87.900 ;
        RECT 177.400 87.800 177.800 88.200 ;
        RECT 178.200 87.900 178.600 89.900 ;
        RECT 180.600 88.000 181.000 89.900 ;
        RECT 182.200 88.000 182.600 89.900 ;
        RECT 180.600 87.900 182.600 88.000 ;
        RECT 183.000 87.900 183.400 89.900 ;
        RECT 184.100 88.200 184.500 89.900 ;
        RECT 176.200 87.200 176.600 87.400 ;
        RECT 174.200 86.800 175.500 87.200 ;
        RECT 176.200 86.900 177.000 87.200 ;
        RECT 176.600 86.800 177.000 86.900 ;
        RECT 172.600 85.400 173.200 85.800 ;
        RECT 172.600 85.100 172.900 85.400 ;
        RECT 175.200 85.200 175.500 86.800 ;
        RECT 175.800 86.100 176.200 86.600 ;
        RECT 178.300 86.200 178.600 87.900 ;
        RECT 180.700 87.700 182.500 87.900 ;
        RECT 181.000 87.200 181.400 87.400 ;
        RECT 183.000 87.200 183.300 87.900 ;
        RECT 183.800 87.800 185.000 88.200 ;
        RECT 188.100 88.000 188.500 89.500 ;
        RECT 190.200 88.500 190.600 89.500 ;
        RECT 183.800 87.200 184.100 87.800 ;
        RECT 179.000 86.400 179.400 87.200 ;
        RECT 180.600 86.900 181.400 87.200 ;
        RECT 180.600 86.800 181.000 86.900 ;
        RECT 182.100 86.800 183.400 87.200 ;
        RECT 183.800 86.800 184.200 87.200 ;
        RECT 176.600 86.100 177.000 86.200 ;
        RECT 175.800 85.800 177.000 86.100 ;
        RECT 177.400 86.100 177.800 86.200 ;
        RECT 178.200 86.100 178.600 86.200 ;
        RECT 179.800 86.100 180.200 86.200 ;
        RECT 177.400 85.800 178.600 86.100 ;
        RECT 179.400 85.800 180.200 86.100 ;
        RECT 181.400 85.800 181.800 86.600 ;
        RECT 155.800 84.800 157.800 85.100 ;
        RECT 155.800 81.100 156.200 84.800 ;
        RECT 157.400 81.100 157.800 84.800 ;
        RECT 158.200 81.100 158.600 85.100 ;
        RECT 159.000 84.800 161.000 85.100 ;
        RECT 159.000 81.100 159.400 84.800 ;
        RECT 160.600 81.100 161.000 84.800 ;
        RECT 161.400 81.100 161.800 85.100 ;
        RECT 162.200 84.800 164.200 85.100 ;
        RECT 162.200 81.100 162.600 84.800 ;
        RECT 163.800 81.100 164.200 84.800 ;
        RECT 164.600 81.100 165.000 85.100 ;
        RECT 165.400 84.800 166.100 85.100 ;
        RECT 166.400 84.800 166.900 85.100 ;
        RECT 168.600 84.800 169.300 85.100 ;
        RECT 169.600 84.800 170.100 85.100 ;
        RECT 165.800 84.200 166.100 84.800 ;
        RECT 165.800 83.800 166.200 84.200 ;
        RECT 166.500 81.100 166.900 84.800 ;
        RECT 169.000 84.200 169.300 84.800 ;
        RECT 169.000 83.800 169.400 84.200 ;
        RECT 169.700 81.100 170.100 84.800 ;
        RECT 171.800 84.800 172.900 85.100 ;
        RECT 174.200 85.100 174.600 85.200 ;
        RECT 174.200 84.800 174.900 85.100 ;
        RECT 175.200 84.800 176.200 85.200 ;
        RECT 177.500 85.100 177.800 85.800 ;
        RECT 179.400 85.600 179.800 85.800 ;
        RECT 182.100 85.100 182.400 86.800 ;
        RECT 183.000 85.100 183.400 85.200 ;
        RECT 171.800 81.100 172.200 84.800 ;
        RECT 174.600 84.200 174.900 84.800 ;
        RECT 174.600 83.800 175.000 84.200 ;
        RECT 175.300 81.100 175.700 84.800 ;
        RECT 177.400 81.100 177.800 85.100 ;
        RECT 178.200 84.800 180.200 85.100 ;
        RECT 178.200 81.100 178.600 84.800 ;
        RECT 179.800 81.100 180.200 84.800 ;
        RECT 181.900 84.800 182.400 85.100 ;
        RECT 182.700 84.800 183.400 85.100 ;
        RECT 181.900 81.100 182.300 84.800 ;
        RECT 182.700 84.200 183.000 84.800 ;
        RECT 183.800 84.400 184.200 85.200 ;
        RECT 182.600 83.800 183.000 84.200 ;
        RECT 184.600 81.100 185.000 87.800 ;
        RECT 187.700 87.700 188.500 88.000 ;
        RECT 185.400 86.800 185.800 87.600 ;
        RECT 187.700 87.500 188.100 87.700 ;
        RECT 187.700 87.200 188.000 87.500 ;
        RECT 190.300 87.400 190.600 88.500 ;
        RECT 192.600 88.000 193.000 89.900 ;
        RECT 194.200 88.000 194.600 89.900 ;
        RECT 192.600 87.900 194.600 88.000 ;
        RECT 195.000 87.900 195.400 89.900 ;
        RECT 196.100 88.200 196.500 89.900 ;
        RECT 196.100 87.900 197.000 88.200 ;
        RECT 192.700 87.700 194.500 87.900 ;
        RECT 187.000 86.800 188.000 87.200 ;
        RECT 188.500 87.100 190.600 87.400 ;
        RECT 193.000 87.200 193.400 87.400 ;
        RECT 195.000 87.200 195.300 87.900 ;
        RECT 188.500 86.900 189.000 87.100 ;
        RECT 187.000 85.400 187.400 86.200 ;
        RECT 187.700 84.900 188.000 86.800 ;
        RECT 188.300 86.500 189.000 86.900 ;
        RECT 192.600 86.900 193.400 87.200 ;
        RECT 194.100 87.100 195.400 87.200 ;
        RECT 195.800 87.100 196.200 87.200 ;
        RECT 192.600 86.800 193.000 86.900 ;
        RECT 194.100 86.800 196.200 87.100 ;
        RECT 188.700 85.500 189.000 86.500 ;
        RECT 189.400 85.800 189.800 86.600 ;
        RECT 190.200 86.100 190.600 86.600 ;
        RECT 192.600 86.100 193.000 86.200 ;
        RECT 190.200 85.800 193.000 86.100 ;
        RECT 193.400 85.800 193.800 86.600 ;
        RECT 188.700 85.200 190.600 85.500 ;
        RECT 187.700 84.600 188.500 84.900 ;
        RECT 188.100 82.200 188.500 84.600 ;
        RECT 190.300 83.500 190.600 85.200 ;
        RECT 194.100 85.100 194.400 86.800 ;
        RECT 196.600 86.100 197.000 87.900 ;
        RECT 198.200 87.700 198.600 89.900 ;
        RECT 200.300 89.200 200.900 89.900 ;
        RECT 200.300 88.900 201.000 89.200 ;
        RECT 202.600 88.900 203.000 89.900 ;
        RECT 204.800 89.200 205.200 89.900 ;
        RECT 204.800 88.900 205.800 89.200 ;
        RECT 200.600 88.500 201.000 88.900 ;
        RECT 202.700 88.600 203.000 88.900 ;
        RECT 202.700 88.300 204.100 88.600 ;
        RECT 203.700 88.200 204.100 88.300 ;
        RECT 204.600 88.200 205.000 88.600 ;
        RECT 205.400 88.500 205.800 88.900 ;
        RECT 199.700 87.700 200.100 87.800 ;
        RECT 197.400 87.100 197.800 87.600 ;
        RECT 198.200 87.400 200.100 87.700 ;
        RECT 198.200 87.100 198.600 87.400 ;
        RECT 197.400 86.800 198.600 87.100 ;
        RECT 201.400 87.100 202.100 87.200 ;
        RECT 204.600 87.100 204.900 88.200 ;
        RECT 207.000 87.500 207.400 89.900 ;
        RECT 207.800 88.500 208.200 89.500 ;
        RECT 207.800 87.400 208.100 88.500 ;
        RECT 209.900 88.000 210.300 89.500 ;
        RECT 209.900 87.700 210.700 88.000 ;
        RECT 210.300 87.500 210.700 87.700 ;
        RECT 206.200 87.100 207.000 87.200 ;
        RECT 207.800 87.100 209.900 87.400 ;
        RECT 201.400 86.800 207.000 87.100 ;
        RECT 209.400 86.900 209.900 87.100 ;
        RECT 210.400 87.200 210.700 87.500 ;
        RECT 212.600 87.700 213.000 89.900 ;
        RECT 214.700 89.200 215.300 89.900 ;
        RECT 214.700 88.900 215.400 89.200 ;
        RECT 217.000 88.900 217.400 89.900 ;
        RECT 219.200 89.200 219.600 89.900 ;
        RECT 219.200 88.900 220.200 89.200 ;
        RECT 215.000 88.500 215.400 88.900 ;
        RECT 217.100 88.600 217.400 88.900 ;
        RECT 217.100 88.300 218.500 88.600 ;
        RECT 218.100 88.200 218.500 88.300 ;
        RECT 219.000 88.200 219.400 88.600 ;
        RECT 219.800 88.500 220.200 88.900 ;
        RECT 214.100 87.700 214.500 87.800 ;
        RECT 212.600 87.400 214.600 87.700 ;
        RECT 195.000 85.800 197.000 86.100 ;
        RECT 195.000 85.200 195.300 85.800 ;
        RECT 195.000 85.100 195.400 85.200 ;
        RECT 188.100 81.800 189.000 82.200 ;
        RECT 188.100 81.100 188.500 81.800 ;
        RECT 190.200 81.500 190.600 83.500 ;
        RECT 193.900 84.800 194.400 85.100 ;
        RECT 194.700 84.800 195.400 85.100 ;
        RECT 193.900 81.100 194.300 84.800 ;
        RECT 194.700 84.200 195.000 84.800 ;
        RECT 195.800 84.400 196.200 85.200 ;
        RECT 194.600 83.800 195.000 84.200 ;
        RECT 196.600 81.100 197.000 85.800 ;
        RECT 198.200 85.700 198.600 86.800 ;
        RECT 200.600 86.400 201.000 86.500 ;
        RECT 199.100 86.100 201.000 86.400 ;
        RECT 199.100 86.000 199.500 86.100 ;
        RECT 199.900 85.700 200.300 85.800 ;
        RECT 198.200 85.400 200.300 85.700 ;
        RECT 198.200 81.100 198.600 85.400 ;
        RECT 201.500 85.200 201.800 86.800 ;
        RECT 205.100 86.700 205.500 86.800 ;
        RECT 205.900 86.200 206.300 86.300 ;
        RECT 203.800 85.900 206.300 86.200 ;
        RECT 203.800 85.800 204.200 85.900 ;
        RECT 207.800 85.800 208.200 86.600 ;
        RECT 208.600 85.800 209.000 86.600 ;
        RECT 209.400 86.500 210.100 86.900 ;
        RECT 210.400 86.800 211.400 87.200 ;
        RECT 204.600 85.500 207.400 85.600 ;
        RECT 209.400 85.500 209.700 86.500 ;
        RECT 204.500 85.400 207.400 85.500 ;
        RECT 200.600 84.900 201.800 85.200 ;
        RECT 202.500 85.300 207.400 85.400 ;
        RECT 202.500 85.100 204.900 85.300 ;
        RECT 200.600 84.400 200.900 84.900 ;
        RECT 200.200 84.000 200.900 84.400 ;
        RECT 201.700 84.500 202.100 84.600 ;
        RECT 202.500 84.500 202.800 85.100 ;
        RECT 201.700 84.200 202.800 84.500 ;
        RECT 203.100 84.500 205.800 84.800 ;
        RECT 203.100 84.400 203.500 84.500 ;
        RECT 205.400 84.400 205.800 84.500 ;
        RECT 202.300 83.700 202.700 83.800 ;
        RECT 203.700 83.700 204.100 83.800 ;
        RECT 200.600 83.100 201.000 83.500 ;
        RECT 202.300 83.400 204.100 83.700 ;
        RECT 202.700 83.100 203.000 83.400 ;
        RECT 205.400 83.100 205.800 83.500 ;
        RECT 200.300 81.100 200.900 83.100 ;
        RECT 202.600 81.100 203.000 83.100 ;
        RECT 204.800 82.800 205.800 83.100 ;
        RECT 204.800 81.100 205.200 82.800 ;
        RECT 207.000 81.100 207.400 85.300 ;
        RECT 207.800 85.200 209.700 85.500 ;
        RECT 207.800 83.500 208.100 85.200 ;
        RECT 210.400 84.900 210.700 86.800 ;
        RECT 211.000 86.100 211.400 86.200 ;
        RECT 212.600 86.100 213.000 87.400 ;
        RECT 214.200 86.800 214.600 87.400 ;
        RECT 216.100 87.100 216.500 87.200 ;
        RECT 219.000 87.100 219.300 88.200 ;
        RECT 221.400 87.500 221.800 89.900 ;
        RECT 223.500 88.200 223.900 89.900 ;
        RECT 223.000 87.900 223.900 88.200 ;
        RECT 224.600 87.900 225.000 89.900 ;
        RECT 225.400 88.000 225.800 89.900 ;
        RECT 227.000 88.000 227.400 89.900 ;
        RECT 229.100 89.200 229.500 89.900 ;
        RECT 228.600 88.800 229.500 89.200 ;
        RECT 229.100 88.200 229.500 88.800 ;
        RECT 225.400 87.900 227.400 88.000 ;
        RECT 228.600 87.900 229.500 88.200 ;
        RECT 220.600 87.100 221.400 87.200 ;
        RECT 215.900 86.800 221.400 87.100 ;
        RECT 222.200 86.800 222.600 87.600 ;
        RECT 215.000 86.400 215.400 86.500 ;
        RECT 211.000 85.800 213.000 86.100 ;
        RECT 213.500 86.100 215.400 86.400 ;
        RECT 213.500 86.000 213.900 86.100 ;
        RECT 211.000 85.400 211.400 85.800 ;
        RECT 212.600 85.700 213.000 85.800 ;
        RECT 214.300 85.700 214.700 85.800 ;
        RECT 212.600 85.400 214.700 85.700 ;
        RECT 209.900 84.600 210.700 84.900 ;
        RECT 207.800 81.500 208.200 83.500 ;
        RECT 209.900 82.200 210.300 84.600 ;
        RECT 209.400 81.800 210.300 82.200 ;
        RECT 209.900 81.100 210.300 81.800 ;
        RECT 212.600 81.100 213.000 85.400 ;
        RECT 215.900 85.200 216.200 86.800 ;
        RECT 219.500 86.700 219.900 86.800 ;
        RECT 219.000 86.200 219.400 86.300 ;
        RECT 220.300 86.200 220.700 86.300 ;
        RECT 218.200 85.900 220.700 86.200 ;
        RECT 223.000 86.100 223.400 87.900 ;
        RECT 224.700 87.200 225.000 87.900 ;
        RECT 225.500 87.700 227.300 87.900 ;
        RECT 226.600 87.200 227.000 87.400 ;
        RECT 224.600 86.800 225.900 87.200 ;
        RECT 226.600 86.900 227.400 87.200 ;
        RECT 227.000 86.800 227.400 86.900 ;
        RECT 227.800 86.800 228.200 87.600 ;
        RECT 218.200 85.800 218.600 85.900 ;
        RECT 223.000 85.800 224.900 86.100 ;
        RECT 219.000 85.500 221.800 85.600 ;
        RECT 218.900 85.400 221.800 85.500 ;
        RECT 215.000 84.900 216.200 85.200 ;
        RECT 216.900 85.300 221.800 85.400 ;
        RECT 216.900 85.100 219.300 85.300 ;
        RECT 215.000 84.400 215.300 84.900 ;
        RECT 214.600 84.200 215.300 84.400 ;
        RECT 216.100 84.500 216.500 84.600 ;
        RECT 216.900 84.500 217.200 85.100 ;
        RECT 216.100 84.200 217.200 84.500 ;
        RECT 217.500 84.500 220.200 84.800 ;
        RECT 217.500 84.400 217.900 84.500 ;
        RECT 219.800 84.400 220.200 84.500 ;
        RECT 214.200 84.000 215.300 84.200 ;
        RECT 214.200 83.800 214.900 84.000 ;
        RECT 216.700 83.700 217.100 83.800 ;
        RECT 218.100 83.700 218.500 83.800 ;
        RECT 215.000 83.100 215.400 83.500 ;
        RECT 216.700 83.400 218.500 83.700 ;
        RECT 217.100 83.100 217.400 83.400 ;
        RECT 219.800 83.100 220.200 83.500 ;
        RECT 214.700 81.100 215.300 83.100 ;
        RECT 217.000 81.100 217.400 83.100 ;
        RECT 219.200 82.800 220.200 83.100 ;
        RECT 219.200 81.100 219.600 82.800 ;
        RECT 221.400 81.100 221.800 85.300 ;
        RECT 223.000 81.100 223.400 85.800 ;
        RECT 224.600 85.200 224.900 85.800 ;
        RECT 223.800 84.400 224.200 85.200 ;
        RECT 224.600 85.100 225.000 85.200 ;
        RECT 225.600 85.100 225.900 86.800 ;
        RECT 226.200 85.800 226.600 86.600 ;
        RECT 224.600 84.800 225.300 85.100 ;
        RECT 225.600 84.800 226.100 85.100 ;
        RECT 225.000 84.200 225.300 84.800 ;
        RECT 225.000 83.800 225.400 84.200 ;
        RECT 225.700 81.100 226.100 84.800 ;
        RECT 228.600 81.100 229.000 87.900 ;
        RECT 229.400 84.400 229.800 85.200 ;
        RECT 0.600 75.700 1.000 79.900 ;
        RECT 2.800 78.200 3.200 79.900 ;
        RECT 2.200 77.900 3.200 78.200 ;
        RECT 5.000 77.900 5.400 79.900 ;
        RECT 7.100 77.900 7.700 79.900 ;
        RECT 2.200 77.500 2.600 77.900 ;
        RECT 5.000 77.600 5.300 77.900 ;
        RECT 3.900 77.300 5.700 77.600 ;
        RECT 7.000 77.500 7.400 77.900 ;
        RECT 3.900 77.200 4.300 77.300 ;
        RECT 5.300 77.200 5.700 77.300 ;
        RECT 2.200 76.500 2.600 76.600 ;
        RECT 4.500 76.500 4.900 76.600 ;
        RECT 2.200 76.200 4.900 76.500 ;
        RECT 5.200 76.500 6.300 76.800 ;
        RECT 5.200 75.900 5.500 76.500 ;
        RECT 5.900 76.400 6.300 76.500 ;
        RECT 7.100 76.600 7.800 77.000 ;
        RECT 7.100 76.100 7.400 76.600 ;
        RECT 3.100 75.700 5.500 75.900 ;
        RECT 0.600 75.600 5.500 75.700 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 0.600 75.500 3.500 75.600 ;
        RECT 0.600 75.400 3.400 75.500 ;
        RECT 6.200 75.200 6.500 75.800 ;
        RECT 9.400 75.600 9.800 79.900 ;
        RECT 11.500 77.200 11.900 79.900 ;
        RECT 11.000 76.800 11.900 77.200 ;
        RECT 12.200 76.800 12.600 77.200 ;
        RECT 11.500 76.200 11.900 76.800 ;
        RECT 12.300 76.200 12.600 76.800 ;
        RECT 11.500 75.900 12.000 76.200 ;
        RECT 12.300 75.900 13.000 76.200 ;
        RECT 7.700 75.300 9.800 75.600 ;
        RECT 7.700 75.200 8.100 75.300 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 1.700 74.800 5.000 75.100 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 8.500 74.900 8.900 75.000 ;
        RECT 1.700 74.700 2.100 74.800 ;
        RECT 2.500 74.200 2.900 74.300 ;
        RECT 6.200 74.200 6.500 74.800 ;
        RECT 7.000 74.600 8.900 74.900 ;
        RECT 7.000 74.500 7.400 74.600 ;
        RECT 1.000 73.900 6.500 74.200 ;
        RECT 1.000 73.800 1.800 73.900 ;
        RECT 0.600 71.100 1.000 73.500 ;
        RECT 3.100 72.800 3.400 73.900 ;
        RECT 5.400 73.800 6.300 73.900 ;
        RECT 9.400 73.600 9.800 75.300 ;
        RECT 11.000 74.400 11.400 75.200 ;
        RECT 11.700 74.200 12.000 75.900 ;
        RECT 12.600 75.800 13.000 75.900 ;
        RECT 13.400 75.800 13.800 76.600 ;
        RECT 12.600 75.100 12.900 75.800 ;
        RECT 14.200 75.100 14.600 79.900 ;
        RECT 17.100 76.200 17.500 79.900 ;
        RECT 17.800 76.800 18.200 77.200 ;
        RECT 17.900 76.200 18.200 76.800 ;
        RECT 17.100 75.900 17.600 76.200 ;
        RECT 17.900 75.900 18.600 76.200 ;
        RECT 12.600 74.800 14.600 75.100 ;
        RECT 10.200 74.100 10.600 74.200 ;
        RECT 10.200 73.800 11.000 74.100 ;
        RECT 11.700 73.800 13.000 74.200 ;
        RECT 10.600 73.600 11.000 73.800 ;
        RECT 7.900 73.300 9.800 73.600 ;
        RECT 7.900 73.200 8.300 73.300 ;
        RECT 2.200 72.100 2.600 72.500 ;
        RECT 3.000 72.400 3.400 72.800 ;
        RECT 3.900 72.700 4.300 72.800 ;
        RECT 3.900 72.400 5.300 72.700 ;
        RECT 5.000 72.100 5.300 72.400 ;
        RECT 7.000 72.100 7.400 72.500 ;
        RECT 2.200 71.800 3.200 72.100 ;
        RECT 2.800 71.100 3.200 71.800 ;
        RECT 5.000 71.100 5.400 72.100 ;
        RECT 7.000 71.800 7.700 72.100 ;
        RECT 7.100 71.100 7.700 71.800 ;
        RECT 9.400 71.100 9.800 73.300 ;
        RECT 10.300 73.100 12.100 73.300 ;
        RECT 12.600 73.100 12.900 73.800 ;
        RECT 14.200 73.100 14.600 74.800 ;
        RECT 16.600 74.400 17.000 75.200 ;
        RECT 17.300 74.200 17.600 75.900 ;
        RECT 18.200 75.800 18.600 75.900 ;
        RECT 19.000 75.800 19.400 76.600 ;
        RECT 18.200 75.100 18.500 75.800 ;
        RECT 19.800 75.100 20.200 79.900 ;
        RECT 21.400 75.700 21.800 79.900 ;
        RECT 23.600 78.200 24.000 79.900 ;
        RECT 23.000 77.900 24.000 78.200 ;
        RECT 25.800 77.900 26.200 79.900 ;
        RECT 27.900 77.900 28.500 79.900 ;
        RECT 23.000 77.500 23.400 77.900 ;
        RECT 25.800 77.600 26.100 77.900 ;
        RECT 24.700 77.300 26.500 77.600 ;
        RECT 27.800 77.500 28.200 77.900 ;
        RECT 24.700 77.200 25.100 77.300 ;
        RECT 26.100 77.200 26.500 77.300 ;
        RECT 23.000 76.500 23.400 76.600 ;
        RECT 25.300 76.500 25.700 76.600 ;
        RECT 23.000 76.200 25.700 76.500 ;
        RECT 26.000 76.500 27.100 76.800 ;
        RECT 26.000 75.900 26.300 76.500 ;
        RECT 26.700 76.400 27.100 76.500 ;
        RECT 27.900 76.600 28.600 77.000 ;
        RECT 27.900 76.100 28.200 76.600 ;
        RECT 23.900 75.700 26.300 75.900 ;
        RECT 21.400 75.600 26.300 75.700 ;
        RECT 27.000 75.800 28.200 76.100 ;
        RECT 21.400 75.500 24.300 75.600 ;
        RECT 21.400 75.400 24.200 75.500 ;
        RECT 27.000 75.200 27.300 75.800 ;
        RECT 30.200 75.600 30.600 79.900 ;
        RECT 32.300 75.900 33.300 79.900 ;
        RECT 28.500 75.300 30.600 75.600 ;
        RECT 28.500 75.200 28.900 75.300 ;
        RECT 24.600 75.100 25.000 75.200 ;
        RECT 18.200 74.800 20.200 75.100 ;
        RECT 15.000 73.400 15.400 74.200 ;
        RECT 15.800 74.100 16.200 74.200 ;
        RECT 15.800 73.800 16.600 74.100 ;
        RECT 17.300 73.800 18.600 74.200 ;
        RECT 16.200 73.600 16.600 73.800 ;
        RECT 15.900 73.100 17.700 73.300 ;
        RECT 18.200 73.100 18.500 73.800 ;
        RECT 19.800 73.100 20.200 74.800 ;
        RECT 22.500 74.800 25.000 75.100 ;
        RECT 27.000 74.800 27.400 75.200 ;
        RECT 29.300 74.900 29.700 75.000 ;
        RECT 22.500 74.700 22.900 74.800 ;
        RECT 23.800 74.700 24.200 74.800 ;
        RECT 23.300 74.200 23.700 74.300 ;
        RECT 27.000 74.200 27.300 74.800 ;
        RECT 27.800 74.600 29.700 74.900 ;
        RECT 27.800 74.500 28.200 74.600 ;
        RECT 20.600 73.400 21.000 74.200 ;
        RECT 21.800 73.900 27.300 74.200 ;
        RECT 21.800 73.800 22.600 73.900 ;
        RECT 10.200 73.000 12.200 73.100 ;
        RECT 10.200 71.100 10.600 73.000 ;
        RECT 11.800 71.100 12.200 73.000 ;
        RECT 12.600 71.100 13.000 73.100 ;
        RECT 13.700 72.800 14.600 73.100 ;
        RECT 15.800 73.000 17.800 73.100 ;
        RECT 13.700 71.100 14.100 72.800 ;
        RECT 15.800 71.100 16.200 73.000 ;
        RECT 17.400 71.100 17.800 73.000 ;
        RECT 18.200 71.100 18.600 73.100 ;
        RECT 19.300 72.800 20.200 73.100 ;
        RECT 19.300 71.100 19.700 72.800 ;
        RECT 21.400 71.100 21.800 73.500 ;
        RECT 23.900 72.800 24.200 73.900 ;
        RECT 26.700 73.800 27.100 73.900 ;
        RECT 30.200 73.600 30.600 75.300 ;
        RECT 31.000 73.800 31.400 74.600 ;
        RECT 31.800 74.400 32.200 75.200 ;
        RECT 32.700 74.200 33.000 75.900 ;
        RECT 33.400 74.400 33.800 75.200 ;
        RECT 32.600 74.100 33.000 74.200 ;
        RECT 34.200 74.100 34.600 74.200 ;
        RECT 35.000 74.100 35.400 79.900 ;
        RECT 31.800 73.800 33.000 74.100 ;
        RECT 33.800 73.800 35.400 74.100 ;
        RECT 28.700 73.300 30.600 73.600 ;
        RECT 28.700 73.200 29.100 73.300 ;
        RECT 23.000 72.100 23.400 72.500 ;
        RECT 23.800 72.400 24.200 72.800 ;
        RECT 24.700 72.700 25.100 72.800 ;
        RECT 24.700 72.400 26.100 72.700 ;
        RECT 25.800 72.100 26.100 72.400 ;
        RECT 27.800 72.100 28.200 72.500 ;
        RECT 23.000 71.800 24.000 72.100 ;
        RECT 23.600 71.100 24.000 71.800 ;
        RECT 25.800 71.100 26.200 72.100 ;
        RECT 27.800 71.800 28.500 72.100 ;
        RECT 27.900 71.100 28.500 71.800 ;
        RECT 30.200 71.100 30.600 73.300 ;
        RECT 31.800 73.100 32.100 73.800 ;
        RECT 33.800 73.600 34.200 73.800 ;
        RECT 32.700 73.100 34.500 73.300 ;
        RECT 31.000 71.400 31.400 73.100 ;
        RECT 31.800 71.700 32.200 73.100 ;
        RECT 32.600 73.000 34.600 73.100 ;
        RECT 32.600 71.400 33.000 73.000 ;
        RECT 31.000 71.100 33.000 71.400 ;
        RECT 34.200 71.100 34.600 73.000 ;
        RECT 35.000 71.100 35.400 73.800 ;
        RECT 35.800 72.400 36.200 73.200 ;
        RECT 36.600 72.400 37.000 73.200 ;
        RECT 37.400 72.100 37.800 79.900 ;
        RECT 41.100 75.900 42.100 79.900 ;
        RECT 45.100 79.200 45.500 79.900 ;
        RECT 44.600 78.800 45.500 79.200 ;
        RECT 45.100 76.200 45.500 78.800 ;
        RECT 45.800 76.800 46.200 77.200 ;
        RECT 45.900 76.200 46.200 76.800 ;
        RECT 48.300 76.200 48.700 79.900 ;
        RECT 49.000 76.800 49.400 77.200 ;
        RECT 49.100 76.200 49.400 76.800 ;
        RECT 50.200 76.200 50.600 79.900 ;
        RECT 51.800 76.400 52.200 79.900 ;
        RECT 53.800 76.800 54.200 77.200 ;
        RECT 45.100 75.900 45.600 76.200 ;
        RECT 45.900 75.900 46.600 76.200 ;
        RECT 48.300 75.900 48.800 76.200 ;
        RECT 49.100 75.900 49.800 76.200 ;
        RECT 50.200 75.900 51.500 76.200 ;
        RECT 51.800 75.900 52.300 76.400 ;
        RECT 53.800 76.200 54.100 76.800 ;
        RECT 54.500 76.200 54.900 79.900 ;
        RECT 39.000 74.100 39.400 74.200 ;
        RECT 39.800 74.100 40.200 74.600 ;
        RECT 40.600 74.400 41.000 75.200 ;
        RECT 41.500 74.200 41.800 75.900 ;
        RECT 42.200 74.400 42.600 75.200 ;
        RECT 44.600 74.400 45.000 75.200 ;
        RECT 45.300 74.200 45.600 75.900 ;
        RECT 46.200 75.800 46.600 75.900 ;
        RECT 47.800 74.400 48.200 75.200 ;
        RECT 48.500 74.200 48.800 75.900 ;
        RECT 49.400 75.800 49.800 75.900 ;
        RECT 50.200 74.800 50.700 75.200 ;
        RECT 50.300 74.400 50.700 74.800 ;
        RECT 51.200 74.900 51.500 75.900 ;
        RECT 51.200 74.500 51.700 74.900 ;
        RECT 41.400 74.100 41.800 74.200 ;
        RECT 43.000 74.100 43.400 74.200 ;
        RECT 39.000 73.800 40.200 74.100 ;
        RECT 40.600 73.800 41.800 74.100 ;
        RECT 42.600 73.800 43.400 74.100 ;
        RECT 43.800 74.100 44.200 74.200 ;
        RECT 43.800 73.800 44.600 74.100 ;
        RECT 45.300 73.800 46.600 74.200 ;
        RECT 47.000 74.100 47.400 74.200 ;
        RECT 47.000 73.800 47.800 74.100 ;
        RECT 48.500 73.800 49.800 74.200 ;
        RECT 40.600 73.100 40.900 73.800 ;
        RECT 42.600 73.600 43.000 73.800 ;
        RECT 44.200 73.600 44.600 73.800 ;
        RECT 41.500 73.100 43.300 73.300 ;
        RECT 43.900 73.100 45.700 73.300 ;
        RECT 46.200 73.100 46.500 73.800 ;
        RECT 47.400 73.600 47.800 73.800 ;
        RECT 47.100 73.100 48.900 73.300 ;
        RECT 49.400 73.100 49.700 73.800 ;
        RECT 51.200 73.700 51.500 74.500 ;
        RECT 52.000 74.200 52.300 75.900 ;
        RECT 53.400 75.900 54.100 76.200 ;
        RECT 54.400 75.900 54.900 76.200 ;
        RECT 53.400 75.800 53.800 75.900 ;
        RECT 54.400 74.200 54.700 75.900 ;
        RECT 56.600 75.800 57.000 76.600 ;
        RECT 57.400 76.100 57.800 79.900 ;
        RECT 60.300 76.200 60.700 79.900 ;
        RECT 61.000 76.800 61.400 77.200 ;
        RECT 61.100 76.200 61.400 76.800 ;
        RECT 62.600 76.800 63.000 77.200 ;
        RECT 62.600 76.200 62.900 76.800 ;
        RECT 63.300 76.200 63.700 79.900 ;
        RECT 58.200 76.100 58.600 76.200 ;
        RECT 57.400 75.800 58.600 76.100 ;
        RECT 60.300 75.900 60.800 76.200 ;
        RECT 61.100 75.900 61.800 76.200 ;
        RECT 55.000 75.100 55.400 75.200 ;
        RECT 55.800 75.100 56.200 75.200 ;
        RECT 56.600 75.100 56.900 75.800 ;
        RECT 55.000 74.800 56.900 75.100 ;
        RECT 55.000 74.400 55.400 74.800 ;
        RECT 51.800 74.100 52.300 74.200 ;
        RECT 52.600 74.100 53.000 74.200 ;
        RECT 51.800 73.800 53.000 74.100 ;
        RECT 53.400 73.800 54.700 74.200 ;
        RECT 55.800 74.100 56.200 74.200 ;
        RECT 55.400 73.800 56.200 74.100 ;
        RECT 50.200 73.400 51.500 73.700 ;
        RECT 38.200 72.100 38.600 72.200 ;
        RECT 37.400 71.800 38.600 72.100 ;
        RECT 37.400 71.100 37.800 71.800 ;
        RECT 39.800 71.400 40.200 73.100 ;
        RECT 40.600 71.700 41.000 73.100 ;
        RECT 41.400 73.000 43.400 73.100 ;
        RECT 41.400 71.400 41.800 73.000 ;
        RECT 39.800 71.100 41.800 71.400 ;
        RECT 43.000 71.100 43.400 73.000 ;
        RECT 43.800 73.000 45.800 73.100 ;
        RECT 43.800 71.100 44.200 73.000 ;
        RECT 45.400 71.100 45.800 73.000 ;
        RECT 46.200 71.100 46.600 73.100 ;
        RECT 47.000 73.000 49.000 73.100 ;
        RECT 47.000 71.100 47.400 73.000 ;
        RECT 48.600 71.100 49.000 73.000 ;
        RECT 49.400 71.100 49.800 73.100 ;
        RECT 50.200 71.100 50.600 73.400 ;
        RECT 52.000 73.100 52.300 73.800 ;
        RECT 53.500 73.100 53.800 73.800 ;
        RECT 55.400 73.600 55.800 73.800 ;
        RECT 54.300 73.100 56.100 73.300 ;
        RECT 57.400 73.100 57.800 75.800 ;
        RECT 59.800 74.400 60.200 75.200 ;
        RECT 60.500 74.200 60.800 75.900 ;
        RECT 61.400 75.800 61.800 75.900 ;
        RECT 62.200 75.900 62.900 76.200 ;
        RECT 63.200 75.900 63.700 76.200 ;
        RECT 66.700 76.200 67.100 79.900 ;
        RECT 67.400 76.800 67.800 77.200 ;
        RECT 67.500 76.200 67.800 76.800 ;
        RECT 66.700 75.900 67.200 76.200 ;
        RECT 67.500 75.900 68.200 76.200 ;
        RECT 62.200 75.800 62.600 75.900 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 61.400 74.200 61.700 74.800 ;
        RECT 63.200 74.200 63.500 75.900 ;
        RECT 63.800 74.400 64.200 75.200 ;
        RECT 66.200 74.400 66.600 75.200 ;
        RECT 66.900 74.200 67.200 75.900 ;
        RECT 67.800 75.800 68.200 75.900 ;
        RECT 68.600 75.800 69.000 76.600 ;
        RECT 67.800 75.100 68.100 75.800 ;
        RECT 69.400 75.100 69.800 79.900 ;
        RECT 67.800 74.800 69.800 75.100 ;
        RECT 58.200 73.400 58.600 74.200 ;
        RECT 59.000 74.100 59.400 74.200 ;
        RECT 59.000 73.800 59.800 74.100 ;
        RECT 60.500 73.800 61.800 74.200 ;
        RECT 62.200 73.800 63.500 74.200 ;
        RECT 64.600 74.100 65.000 74.200 ;
        RECT 64.200 73.800 65.000 74.100 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 65.400 73.800 66.200 74.100 ;
        RECT 66.900 73.800 68.200 74.200 ;
        RECT 59.400 73.600 59.800 73.800 ;
        RECT 59.100 73.100 60.900 73.300 ;
        RECT 61.400 73.100 61.700 73.800 ;
        RECT 62.300 73.100 62.600 73.800 ;
        RECT 64.200 73.600 64.600 73.800 ;
        RECT 65.800 73.600 66.200 73.800 ;
        RECT 63.100 73.100 64.900 73.300 ;
        RECT 65.500 73.100 67.300 73.300 ;
        RECT 67.800 73.100 68.100 73.800 ;
        RECT 69.400 73.100 69.800 74.800 ;
        RECT 71.000 75.600 71.400 79.900 ;
        RECT 73.100 77.900 73.700 79.900 ;
        RECT 75.400 77.900 75.800 79.900 ;
        RECT 77.600 78.200 78.000 79.900 ;
        RECT 77.600 77.900 78.600 78.200 ;
        RECT 73.400 77.500 73.800 77.900 ;
        RECT 75.500 77.600 75.800 77.900 ;
        RECT 75.100 77.300 76.900 77.600 ;
        RECT 78.200 77.500 78.600 77.900 ;
        RECT 75.100 77.200 75.500 77.300 ;
        RECT 76.500 77.200 76.900 77.300 ;
        RECT 73.000 76.600 73.700 77.000 ;
        RECT 73.400 76.100 73.700 76.600 ;
        RECT 74.500 76.500 75.600 76.800 ;
        RECT 74.500 76.400 74.900 76.500 ;
        RECT 73.400 75.800 74.600 76.100 ;
        RECT 71.000 75.300 73.100 75.600 ;
        RECT 70.200 74.100 70.600 74.200 ;
        RECT 71.000 74.100 71.400 75.300 ;
        RECT 72.700 75.200 73.100 75.300 ;
        RECT 74.300 75.200 74.600 75.800 ;
        RECT 75.300 75.900 75.600 76.500 ;
        RECT 75.900 76.500 76.300 76.600 ;
        RECT 78.200 76.500 78.600 76.600 ;
        RECT 75.900 76.200 78.600 76.500 ;
        RECT 75.300 75.700 77.700 75.900 ;
        RECT 79.800 75.700 80.200 79.900 ;
        RECT 81.900 76.300 82.300 79.900 ;
        RECT 81.400 75.900 82.300 76.300 ;
        RECT 84.300 76.200 84.700 79.900 ;
        RECT 85.000 76.800 85.400 77.200 ;
        RECT 85.100 76.200 85.400 76.800 ;
        RECT 84.300 75.900 84.800 76.200 ;
        RECT 85.100 75.900 85.800 76.200 ;
        RECT 75.300 75.600 80.200 75.700 ;
        RECT 77.300 75.500 80.200 75.600 ;
        RECT 77.400 75.400 80.200 75.500 ;
        RECT 71.900 74.900 72.300 75.000 ;
        RECT 71.900 74.600 73.800 74.900 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 80.600 75.100 81.000 75.200 ;
        RECT 81.500 75.100 81.800 75.900 ;
        RECT 75.000 74.800 79.100 75.100 ;
        RECT 80.600 74.800 81.800 75.100 ;
        RECT 82.200 75.100 82.600 75.600 ;
        RECT 83.000 75.100 83.400 75.200 ;
        RECT 82.200 74.800 83.400 75.100 ;
        RECT 73.400 74.500 73.800 74.600 ;
        RECT 70.200 73.800 71.400 74.100 ;
        RECT 74.300 74.200 74.600 74.800 ;
        RECT 78.700 74.700 79.100 74.800 ;
        RECT 77.900 74.200 78.300 74.300 ;
        RECT 81.500 74.200 81.800 74.800 ;
        RECT 83.800 74.400 84.200 75.200 ;
        RECT 84.500 74.200 84.800 75.900 ;
        RECT 85.400 75.800 85.800 75.900 ;
        RECT 86.200 75.800 86.600 76.600 ;
        RECT 85.400 75.100 85.700 75.800 ;
        RECT 87.000 75.100 87.400 79.900 ;
        RECT 85.400 74.800 87.400 75.100 ;
        RECT 74.300 73.900 79.800 74.200 ;
        RECT 74.500 73.800 74.900 73.900 ;
        RECT 70.200 73.400 70.600 73.800 ;
        RECT 71.000 73.600 71.400 73.800 ;
        RECT 51.800 72.800 52.300 73.100 ;
        RECT 51.800 71.100 52.200 72.800 ;
        RECT 53.400 71.100 53.800 73.100 ;
        RECT 54.200 73.000 56.200 73.100 ;
        RECT 54.200 71.100 54.600 73.000 ;
        RECT 55.800 71.100 56.200 73.000 ;
        RECT 56.900 72.800 57.800 73.100 ;
        RECT 59.000 73.000 61.000 73.100 ;
        RECT 56.900 71.100 57.300 72.800 ;
        RECT 59.000 71.100 59.400 73.000 ;
        RECT 60.600 71.100 61.000 73.000 ;
        RECT 61.400 71.100 61.800 73.100 ;
        RECT 62.200 71.100 62.600 73.100 ;
        RECT 63.000 73.000 65.000 73.100 ;
        RECT 63.000 71.100 63.400 73.000 ;
        RECT 64.600 71.100 65.000 73.000 ;
        RECT 65.400 73.000 67.400 73.100 ;
        RECT 65.400 71.100 65.800 73.000 ;
        RECT 67.000 71.100 67.400 73.000 ;
        RECT 67.800 71.100 68.200 73.100 ;
        RECT 68.900 72.800 69.800 73.100 ;
        RECT 71.000 73.300 72.900 73.600 ;
        RECT 68.900 71.100 69.300 72.800 ;
        RECT 71.000 71.100 71.400 73.300 ;
        RECT 72.500 73.200 72.900 73.300 ;
        RECT 77.400 72.800 77.700 73.900 ;
        RECT 79.000 73.800 79.800 73.900 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 83.000 74.100 83.400 74.200 ;
        RECT 84.500 74.100 85.800 74.200 ;
        RECT 86.200 74.100 86.600 74.200 ;
        RECT 83.000 73.800 83.800 74.100 ;
        RECT 84.500 73.800 86.600 74.100 ;
        RECT 76.500 72.700 76.900 72.800 ;
        RECT 73.400 72.100 73.800 72.500 ;
        RECT 75.500 72.400 76.900 72.700 ;
        RECT 77.400 72.400 77.800 72.800 ;
        RECT 75.500 72.100 75.800 72.400 ;
        RECT 78.200 72.100 78.600 72.500 ;
        RECT 73.100 71.800 73.800 72.100 ;
        RECT 73.100 71.100 73.700 71.800 ;
        RECT 75.400 71.100 75.800 72.100 ;
        RECT 77.600 71.800 78.600 72.100 ;
        RECT 77.600 71.100 78.000 71.800 ;
        RECT 79.800 71.100 80.200 73.500 ;
        RECT 80.600 72.400 81.000 73.200 ;
        RECT 81.500 72.100 81.800 73.800 ;
        RECT 83.400 73.600 83.800 73.800 ;
        RECT 83.100 73.100 84.900 73.300 ;
        RECT 85.400 73.100 85.700 73.800 ;
        RECT 87.000 73.100 87.400 74.800 ;
        RECT 90.200 75.600 90.600 79.900 ;
        RECT 92.300 77.900 92.900 79.900 ;
        RECT 94.600 77.900 95.000 79.900 ;
        RECT 96.800 78.200 97.200 79.900 ;
        RECT 96.800 77.900 97.800 78.200 ;
        RECT 92.600 77.500 93.000 77.900 ;
        RECT 94.700 77.600 95.000 77.900 ;
        RECT 94.300 77.300 96.100 77.600 ;
        RECT 97.400 77.500 97.800 77.900 ;
        RECT 94.300 77.200 94.700 77.300 ;
        RECT 95.700 77.200 96.100 77.300 ;
        RECT 92.200 76.600 92.900 77.000 ;
        RECT 92.600 76.100 92.900 76.600 ;
        RECT 93.700 76.500 94.800 76.800 ;
        RECT 93.700 76.400 94.100 76.500 ;
        RECT 92.600 75.800 93.800 76.100 ;
        RECT 90.200 75.300 92.300 75.600 ;
        RECT 87.800 74.100 88.200 74.200 ;
        RECT 89.400 74.100 89.800 74.200 ;
        RECT 87.800 73.800 89.800 74.100 ;
        RECT 87.800 73.400 88.200 73.800 ;
        RECT 90.200 73.600 90.600 75.300 ;
        RECT 91.900 75.200 92.300 75.300 ;
        RECT 93.500 75.200 93.800 75.800 ;
        RECT 94.500 75.900 94.800 76.500 ;
        RECT 95.100 76.500 95.500 76.600 ;
        RECT 97.400 76.500 97.800 76.600 ;
        RECT 95.100 76.200 97.800 76.500 ;
        RECT 94.500 75.700 96.900 75.900 ;
        RECT 99.000 75.700 99.400 79.900 ;
        RECT 94.500 75.600 99.400 75.700 ;
        RECT 96.500 75.500 99.400 75.600 ;
        RECT 99.800 77.500 100.200 79.500 ;
        RECT 99.800 75.800 100.100 77.500 ;
        RECT 101.900 76.400 102.300 79.900 ;
        RECT 105.400 77.900 105.800 79.900 ;
        RECT 105.500 77.800 105.800 77.900 ;
        RECT 107.000 77.900 107.400 79.900 ;
        RECT 107.000 77.800 107.300 77.900 ;
        RECT 105.500 77.500 107.300 77.800 ;
        RECT 106.200 76.400 106.600 77.200 ;
        RECT 101.900 76.100 102.700 76.400 ;
        RECT 107.000 76.200 107.300 77.500 ;
        RECT 99.800 75.500 101.700 75.800 ;
        RECT 96.600 75.400 99.400 75.500 ;
        RECT 91.100 74.900 91.500 75.000 ;
        RECT 91.100 74.600 93.000 74.900 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 95.800 75.100 96.200 75.200 ;
        RECT 95.800 74.800 98.300 75.100 ;
        RECT 92.600 74.500 93.000 74.600 ;
        RECT 93.500 74.200 93.800 74.800 ;
        RECT 97.900 74.700 98.300 74.800 ;
        RECT 99.800 74.400 100.200 75.200 ;
        RECT 100.600 74.400 101.000 75.200 ;
        RECT 101.400 74.500 101.700 75.500 ;
        RECT 97.100 74.200 97.500 74.300 ;
        RECT 93.500 73.900 99.000 74.200 ;
        RECT 101.400 74.100 102.100 74.500 ;
        RECT 102.400 74.200 102.700 76.100 ;
        RECT 103.000 74.800 103.400 75.600 ;
        RECT 104.600 75.400 105.000 76.200 ;
        RECT 107.000 75.800 107.400 76.200 ;
        RECT 107.800 75.800 108.200 76.600 ;
        RECT 105.400 74.800 106.200 75.200 ;
        RECT 107.000 74.200 107.300 75.800 ;
        RECT 102.400 74.100 103.400 74.200 ;
        RECT 103.800 74.100 104.200 74.200 ;
        RECT 106.500 74.100 107.300 74.200 ;
        RECT 101.400 73.900 101.900 74.100 ;
        RECT 93.700 73.800 94.100 73.900 ;
        RECT 81.400 71.100 81.800 72.100 ;
        RECT 83.000 73.000 85.000 73.100 ;
        RECT 83.000 71.100 83.400 73.000 ;
        RECT 84.600 71.100 85.000 73.000 ;
        RECT 85.400 71.100 85.800 73.100 ;
        RECT 86.500 72.800 87.400 73.100 ;
        RECT 90.200 73.300 92.200 73.600 ;
        RECT 86.500 71.100 86.900 72.800 ;
        RECT 89.400 72.100 89.800 72.200 ;
        RECT 90.200 72.100 90.600 73.300 ;
        RECT 91.700 73.200 92.200 73.300 ;
        RECT 91.800 72.800 92.200 73.200 ;
        RECT 96.600 72.800 96.900 73.900 ;
        RECT 98.200 73.800 99.000 73.900 ;
        RECT 99.800 73.600 101.900 73.900 ;
        RECT 102.400 73.800 104.200 74.100 ;
        RECT 106.400 73.900 107.300 74.100 ;
        RECT 107.800 74.100 108.200 74.200 ;
        RECT 108.600 74.100 109.000 79.900 ;
        RECT 111.500 79.200 111.900 79.900 ;
        RECT 111.000 78.800 111.900 79.200 ;
        RECT 111.500 76.200 111.900 78.800 ;
        RECT 114.200 77.900 114.600 79.900 ;
        RECT 114.300 77.800 114.600 77.900 ;
        RECT 115.800 77.900 116.200 79.900 ;
        RECT 115.800 77.800 116.100 77.900 ;
        RECT 114.300 77.500 116.100 77.800 ;
        RECT 112.200 76.800 112.600 77.200 ;
        RECT 112.300 76.200 112.600 76.800 ;
        RECT 115.000 76.400 115.400 77.200 ;
        RECT 115.800 76.200 116.100 77.500 ;
        RECT 117.400 76.400 117.800 79.900 ;
        RECT 111.500 75.900 112.000 76.200 ;
        RECT 112.300 75.900 113.000 76.200 ;
        RECT 111.000 74.400 111.400 75.200 ;
        RECT 111.700 74.200 112.000 75.900 ;
        RECT 112.600 75.800 113.000 75.900 ;
        RECT 113.400 75.400 113.800 76.200 ;
        RECT 115.800 75.800 116.200 76.200 ;
        RECT 117.300 75.900 117.800 76.400 ;
        RECT 119.000 76.200 119.400 79.900 ;
        RECT 118.100 75.900 119.400 76.200 ;
        RECT 114.200 74.800 115.000 75.200 ;
        RECT 115.800 74.200 116.100 75.800 ;
        RECT 95.700 72.700 96.100 72.800 ;
        RECT 92.600 72.100 93.000 72.500 ;
        RECT 94.700 72.400 96.100 72.700 ;
        RECT 96.600 72.400 97.000 72.800 ;
        RECT 94.700 72.100 95.000 72.400 ;
        RECT 97.400 72.100 97.800 72.500 ;
        RECT 89.400 71.800 90.600 72.100 ;
        RECT 90.200 71.100 90.600 71.800 ;
        RECT 92.300 71.800 93.000 72.100 ;
        RECT 92.300 71.100 92.900 71.800 ;
        RECT 94.600 71.100 95.000 72.100 ;
        RECT 96.800 71.800 97.800 72.100 ;
        RECT 96.800 71.100 97.200 71.800 ;
        RECT 99.000 71.100 99.400 73.500 ;
        RECT 99.800 72.500 100.100 73.600 ;
        RECT 102.400 73.500 102.700 73.800 ;
        RECT 102.300 73.300 102.700 73.500 ;
        RECT 101.900 73.000 102.700 73.300 ;
        RECT 99.800 71.500 100.200 72.500 ;
        RECT 101.900 71.500 102.300 73.000 ;
        RECT 106.400 72.200 106.800 73.900 ;
        RECT 107.800 73.800 109.000 74.100 ;
        RECT 108.600 73.100 109.000 73.800 ;
        RECT 109.400 73.400 109.800 74.200 ;
        RECT 110.200 74.100 110.600 74.200 ;
        RECT 110.200 73.800 111.000 74.100 ;
        RECT 111.700 73.800 113.000 74.200 ;
        RECT 115.300 74.100 116.100 74.200 ;
        RECT 115.200 73.900 116.100 74.100 ;
        RECT 117.300 74.200 117.600 75.900 ;
        RECT 118.100 74.900 118.400 75.900 ;
        RECT 119.800 75.800 120.200 76.200 ;
        RECT 117.900 74.500 118.400 74.900 ;
        RECT 110.600 73.600 111.000 73.800 ;
        RECT 110.300 73.100 112.100 73.300 ;
        RECT 112.600 73.100 112.900 73.800 ;
        RECT 106.200 71.800 106.800 72.200 ;
        RECT 106.400 71.100 106.800 71.800 ;
        RECT 108.100 72.800 109.000 73.100 ;
        RECT 110.200 73.000 112.200 73.100 ;
        RECT 108.100 71.100 108.500 72.800 ;
        RECT 110.200 71.100 110.600 73.000 ;
        RECT 111.800 71.100 112.200 73.000 ;
        RECT 112.600 71.100 113.000 73.100 ;
        RECT 115.200 71.100 115.600 73.900 ;
        RECT 117.300 73.800 117.800 74.200 ;
        RECT 117.300 73.100 117.600 73.800 ;
        RECT 118.100 73.700 118.400 74.500 ;
        RECT 118.900 75.100 119.400 75.200 ;
        RECT 119.800 75.100 120.100 75.800 ;
        RECT 118.900 74.800 120.100 75.100 ;
        RECT 118.900 74.400 119.300 74.800 ;
        RECT 118.100 73.400 119.400 73.700 ;
        RECT 119.800 73.400 120.200 74.200 ;
        RECT 117.300 72.800 117.800 73.100 ;
        RECT 117.400 71.100 117.800 72.800 ;
        RECT 119.000 71.100 119.400 73.400 ;
        RECT 120.600 73.100 121.000 79.900 ;
        RECT 121.400 75.800 121.800 76.600 ;
        RECT 123.000 76.400 123.400 79.900 ;
        RECT 122.900 75.900 123.400 76.400 ;
        RECT 124.600 76.200 125.000 79.900 ;
        RECT 123.700 75.900 125.000 76.200 ;
        RECT 122.900 74.200 123.200 75.900 ;
        RECT 123.700 74.900 124.000 75.900 ;
        RECT 125.400 75.700 125.800 79.900 ;
        RECT 127.600 78.200 128.000 79.900 ;
        RECT 127.000 77.900 128.000 78.200 ;
        RECT 129.800 77.900 130.200 79.900 ;
        RECT 131.900 77.900 132.500 79.900 ;
        RECT 127.000 77.500 127.400 77.900 ;
        RECT 129.800 77.600 130.100 77.900 ;
        RECT 128.700 77.300 130.500 77.600 ;
        RECT 131.800 77.500 132.200 77.900 ;
        RECT 128.700 77.200 129.100 77.300 ;
        RECT 130.100 77.200 130.500 77.300 ;
        RECT 127.000 76.500 127.400 76.600 ;
        RECT 129.300 76.500 129.700 76.600 ;
        RECT 127.000 76.200 129.700 76.500 ;
        RECT 130.000 76.500 131.100 76.800 ;
        RECT 130.000 75.900 130.300 76.500 ;
        RECT 130.700 76.400 131.100 76.500 ;
        RECT 131.900 76.600 132.600 77.000 ;
        RECT 131.900 76.100 132.200 76.600 ;
        RECT 127.900 75.700 130.300 75.900 ;
        RECT 125.400 75.600 130.300 75.700 ;
        RECT 131.000 75.800 132.200 76.100 ;
        RECT 125.400 75.500 128.300 75.600 ;
        RECT 125.400 75.400 128.200 75.500 ;
        RECT 131.000 75.200 131.300 75.800 ;
        RECT 134.200 75.600 134.600 79.900 ;
        RECT 136.300 76.200 136.700 79.900 ;
        RECT 137.000 76.800 137.400 77.200 ;
        RECT 137.100 76.200 137.400 76.800 ;
        RECT 136.300 75.900 136.800 76.200 ;
        RECT 137.100 75.900 137.800 76.200 ;
        RECT 132.500 75.300 134.600 75.600 ;
        RECT 132.500 75.200 132.900 75.300 ;
        RECT 123.500 74.500 124.000 74.900 ;
        RECT 122.200 74.100 122.600 74.200 ;
        RECT 122.900 74.100 123.400 74.200 ;
        RECT 122.200 73.800 123.400 74.100 ;
        RECT 122.900 73.100 123.200 73.800 ;
        RECT 123.700 73.700 124.000 74.500 ;
        RECT 124.500 74.800 125.000 75.200 ;
        RECT 128.600 75.100 129.000 75.200 ;
        RECT 130.200 75.100 130.600 75.200 ;
        RECT 126.500 74.800 130.600 75.100 ;
        RECT 131.000 74.800 131.400 75.200 ;
        RECT 133.300 74.900 133.700 75.000 ;
        RECT 124.500 74.400 124.900 74.800 ;
        RECT 126.500 74.700 126.900 74.800 ;
        RECT 127.300 74.200 127.700 74.300 ;
        RECT 131.000 74.200 131.300 74.800 ;
        RECT 131.800 74.600 133.700 74.900 ;
        RECT 131.800 74.500 132.200 74.600 ;
        RECT 125.800 73.900 131.300 74.200 ;
        RECT 125.800 73.800 126.600 73.900 ;
        RECT 123.700 73.400 125.000 73.700 ;
        RECT 120.600 72.800 121.500 73.100 ;
        RECT 122.900 72.800 123.400 73.100 ;
        RECT 121.100 72.200 121.500 72.800 ;
        RECT 121.100 71.800 121.800 72.200 ;
        RECT 121.100 71.100 121.500 71.800 ;
        RECT 123.000 71.100 123.400 72.800 ;
        RECT 124.600 71.100 125.000 73.400 ;
        RECT 125.400 71.100 125.800 73.500 ;
        RECT 127.900 72.800 128.200 73.900 ;
        RECT 130.700 73.800 131.100 73.900 ;
        RECT 134.200 73.600 134.600 75.300 ;
        RECT 136.500 75.200 136.800 75.900 ;
        RECT 137.400 75.800 137.800 75.900 ;
        RECT 138.200 75.800 138.600 76.600 ;
        RECT 135.000 75.100 135.400 75.200 ;
        RECT 135.800 75.100 136.200 75.200 ;
        RECT 135.000 74.800 136.200 75.100 ;
        RECT 135.800 74.400 136.200 74.800 ;
        RECT 136.500 74.800 137.000 75.200 ;
        RECT 137.400 75.100 137.700 75.800 ;
        RECT 139.000 75.100 139.400 79.900 ;
        RECT 143.500 76.200 143.900 79.900 ;
        RECT 144.200 76.800 144.600 77.200 ;
        RECT 144.300 76.200 144.600 76.800 ;
        RECT 143.500 75.900 144.000 76.200 ;
        RECT 144.300 75.900 145.000 76.200 ;
        RECT 143.700 75.200 144.000 75.900 ;
        RECT 144.600 75.800 145.000 75.900 ;
        RECT 145.400 75.800 145.800 76.600 ;
        RECT 137.400 74.800 139.400 75.100 ;
        RECT 136.500 74.200 136.800 74.800 ;
        RECT 135.000 74.100 135.400 74.200 ;
        RECT 135.000 73.800 135.800 74.100 ;
        RECT 136.500 73.800 137.800 74.200 ;
        RECT 135.400 73.600 135.800 73.800 ;
        RECT 132.700 73.300 134.600 73.600 ;
        RECT 132.700 73.200 133.100 73.300 ;
        RECT 127.000 72.100 127.400 72.500 ;
        RECT 127.800 72.400 128.200 72.800 ;
        RECT 128.700 72.700 129.100 72.800 ;
        RECT 128.700 72.400 130.100 72.700 ;
        RECT 129.800 72.100 130.100 72.400 ;
        RECT 131.800 72.100 132.200 72.500 ;
        RECT 127.000 71.800 128.000 72.100 ;
        RECT 127.600 71.100 128.000 71.800 ;
        RECT 129.800 71.100 130.200 72.100 ;
        RECT 131.800 71.800 132.500 72.100 ;
        RECT 131.900 71.100 132.500 71.800 ;
        RECT 134.200 71.100 134.600 73.300 ;
        RECT 135.100 73.100 136.900 73.300 ;
        RECT 137.400 73.100 137.700 73.800 ;
        RECT 139.000 73.100 139.400 74.800 ;
        RECT 143.000 74.400 143.400 75.200 ;
        RECT 143.700 74.800 144.200 75.200 ;
        RECT 144.600 75.100 144.900 75.800 ;
        RECT 146.200 75.100 146.600 79.900 ;
        RECT 147.800 75.700 148.200 79.900 ;
        RECT 150.000 78.200 150.400 79.900 ;
        RECT 149.400 77.900 150.400 78.200 ;
        RECT 152.200 77.900 152.600 79.900 ;
        RECT 154.300 77.900 154.900 79.900 ;
        RECT 149.400 77.500 149.800 77.900 ;
        RECT 152.200 77.600 152.500 77.900 ;
        RECT 151.100 77.300 152.900 77.600 ;
        RECT 154.200 77.500 154.600 77.900 ;
        RECT 151.100 77.200 151.500 77.300 ;
        RECT 152.500 77.200 152.900 77.300 ;
        RECT 149.400 76.500 149.800 76.600 ;
        RECT 151.700 76.500 152.100 76.600 ;
        RECT 149.400 76.200 152.100 76.500 ;
        RECT 152.400 76.500 153.500 76.800 ;
        RECT 152.400 75.900 152.700 76.500 ;
        RECT 153.100 76.400 153.500 76.500 ;
        RECT 154.300 76.600 155.000 77.000 ;
        RECT 154.300 76.100 154.600 76.600 ;
        RECT 150.300 75.700 152.700 75.900 ;
        RECT 147.800 75.600 152.700 75.700 ;
        RECT 153.400 75.800 154.600 76.100 ;
        RECT 147.800 75.500 150.700 75.600 ;
        RECT 147.800 75.400 150.600 75.500 ;
        RECT 151.000 75.100 151.400 75.200 ;
        RECT 144.600 74.800 146.600 75.100 ;
        RECT 143.700 74.200 144.000 74.800 ;
        RECT 139.800 73.400 140.200 74.200 ;
        RECT 142.200 74.100 142.600 74.200 ;
        RECT 142.200 73.800 143.000 74.100 ;
        RECT 143.700 73.800 145.000 74.200 ;
        RECT 142.600 73.600 143.000 73.800 ;
        RECT 142.300 73.100 144.100 73.300 ;
        RECT 144.600 73.100 144.900 73.800 ;
        RECT 146.200 73.100 146.600 74.800 ;
        RECT 148.900 74.800 151.400 75.100 ;
        RECT 148.900 74.700 149.300 74.800 ;
        RECT 150.200 74.700 150.600 74.800 ;
        RECT 149.700 74.200 150.100 74.300 ;
        RECT 153.400 74.200 153.700 75.800 ;
        RECT 156.600 75.600 157.000 79.900 ;
        RECT 154.900 75.300 157.000 75.600 ;
        RECT 154.900 75.200 155.300 75.300 ;
        RECT 155.700 74.900 156.100 75.000 ;
        RECT 154.200 74.600 156.100 74.900 ;
        RECT 154.200 74.500 154.600 74.600 ;
        RECT 147.000 73.400 147.400 74.200 ;
        RECT 148.200 73.900 153.700 74.200 ;
        RECT 148.200 73.800 149.000 73.900 ;
        RECT 135.000 73.000 137.000 73.100 ;
        RECT 135.000 71.100 135.400 73.000 ;
        RECT 136.600 71.100 137.000 73.000 ;
        RECT 137.400 71.100 137.800 73.100 ;
        RECT 138.500 72.800 139.400 73.100 ;
        RECT 142.200 73.000 144.200 73.100 ;
        RECT 138.500 71.100 138.900 72.800 ;
        RECT 142.200 71.100 142.600 73.000 ;
        RECT 143.800 71.100 144.200 73.000 ;
        RECT 144.600 71.100 145.000 73.100 ;
        RECT 145.700 72.800 146.600 73.100 ;
        RECT 145.700 71.100 146.100 72.800 ;
        RECT 147.800 71.100 148.200 73.500 ;
        RECT 150.300 72.800 150.600 73.900 ;
        RECT 153.100 73.800 153.500 73.900 ;
        RECT 156.600 73.600 157.000 75.300 ;
        RECT 155.100 73.300 157.000 73.600 ;
        RECT 155.100 73.200 155.500 73.300 ;
        RECT 149.400 72.100 149.800 72.500 ;
        RECT 150.200 72.400 150.600 72.800 ;
        RECT 151.100 72.700 151.500 72.800 ;
        RECT 151.100 72.400 152.500 72.700 ;
        RECT 152.200 72.100 152.500 72.400 ;
        RECT 154.200 72.100 154.600 72.500 ;
        RECT 149.400 71.800 150.400 72.100 ;
        RECT 150.000 71.100 150.400 71.800 ;
        RECT 152.200 71.100 152.600 72.100 ;
        RECT 154.200 71.800 154.900 72.100 ;
        RECT 154.300 71.100 154.900 71.800 ;
        RECT 156.600 71.100 157.000 73.300 ;
        RECT 158.200 75.600 158.600 79.900 ;
        RECT 159.800 75.600 160.200 79.900 ;
        RECT 158.200 75.200 160.200 75.600 ;
        RECT 161.400 75.700 161.800 79.900 ;
        RECT 163.600 78.200 164.000 79.900 ;
        RECT 163.000 77.900 164.000 78.200 ;
        RECT 165.800 77.900 166.200 79.900 ;
        RECT 167.900 77.900 168.500 79.900 ;
        RECT 163.000 77.500 163.400 77.900 ;
        RECT 165.800 77.600 166.100 77.900 ;
        RECT 164.700 77.300 166.500 77.600 ;
        RECT 167.800 77.500 168.200 77.900 ;
        RECT 164.700 77.200 165.100 77.300 ;
        RECT 166.100 77.200 166.500 77.300 ;
        RECT 163.000 76.500 163.400 76.600 ;
        RECT 165.300 76.500 165.700 76.600 ;
        RECT 163.000 76.200 165.700 76.500 ;
        RECT 166.000 76.500 167.100 76.800 ;
        RECT 166.000 75.900 166.300 76.500 ;
        RECT 166.700 76.400 167.100 76.500 ;
        RECT 167.900 76.600 168.600 77.000 ;
        RECT 167.900 76.100 168.200 76.600 ;
        RECT 163.900 75.700 166.300 75.900 ;
        RECT 161.400 75.600 166.300 75.700 ;
        RECT 167.000 75.800 168.200 76.100 ;
        RECT 161.400 75.500 164.300 75.600 ;
        RECT 161.400 75.400 164.200 75.500 ;
        RECT 158.200 73.800 158.600 75.200 ;
        RECT 164.600 75.100 165.000 75.200 ;
        RECT 162.500 74.800 165.000 75.100 ;
        RECT 162.500 74.700 162.900 74.800 ;
        RECT 163.300 74.200 163.700 74.300 ;
        RECT 167.000 74.200 167.300 75.800 ;
        RECT 170.200 75.600 170.600 79.900 ;
        RECT 171.000 76.200 171.400 79.900 ;
        RECT 173.800 76.800 174.200 77.200 ;
        RECT 173.800 76.200 174.100 76.800 ;
        RECT 174.500 76.200 174.900 79.900 ;
        RECT 171.000 75.900 172.100 76.200 ;
        RECT 168.500 75.300 170.600 75.600 ;
        RECT 168.500 75.200 168.900 75.300 ;
        RECT 170.200 75.100 170.600 75.300 ;
        RECT 171.800 75.600 172.100 75.900 ;
        RECT 173.400 75.900 174.100 76.200 ;
        RECT 174.400 75.900 174.900 76.200 ;
        RECT 176.600 76.200 177.000 79.900 ;
        RECT 178.200 76.400 178.600 79.900 ;
        RECT 179.800 77.900 180.200 79.900 ;
        RECT 179.900 77.800 180.200 77.900 ;
        RECT 181.400 77.900 181.800 79.900 ;
        RECT 181.400 77.800 181.700 77.900 ;
        RECT 179.900 77.500 181.700 77.800 ;
        RECT 176.600 75.900 177.900 76.200 ;
        RECT 178.200 75.900 178.700 76.400 ;
        RECT 179.900 76.200 180.200 77.500 ;
        RECT 180.600 76.400 181.000 77.200 ;
        RECT 173.400 75.800 173.800 75.900 ;
        RECT 171.800 75.200 172.400 75.600 ;
        RECT 174.400 75.200 174.700 75.900 ;
        RECT 171.000 75.100 171.400 75.200 ;
        RECT 169.300 74.900 169.700 75.000 ;
        RECT 167.800 74.600 169.700 74.900 ;
        RECT 170.200 74.800 171.400 75.100 ;
        RECT 167.800 74.500 168.200 74.600 ;
        RECT 158.200 73.400 160.200 73.800 ;
        RECT 160.600 73.400 161.000 74.200 ;
        RECT 161.800 73.900 167.300 74.200 ;
        RECT 161.800 73.800 162.600 73.900 ;
        RECT 158.200 71.100 158.600 73.400 ;
        RECT 159.800 71.100 160.200 73.400 ;
        RECT 161.400 71.100 161.800 73.500 ;
        RECT 163.900 72.800 164.200 73.900 ;
        RECT 165.400 73.800 165.800 73.900 ;
        RECT 166.700 73.800 167.100 73.900 ;
        RECT 170.200 73.600 170.600 74.800 ;
        RECT 171.000 74.400 171.400 74.800 ;
        RECT 171.800 73.700 172.100 75.200 ;
        RECT 174.200 74.800 174.700 75.200 ;
        RECT 174.400 74.200 174.700 74.800 ;
        RECT 175.000 74.400 175.400 75.200 ;
        RECT 176.600 74.800 177.100 75.200 ;
        RECT 176.700 74.400 177.100 74.800 ;
        RECT 177.600 74.900 177.900 75.900 ;
        RECT 177.600 74.500 178.100 74.900 ;
        RECT 173.400 73.800 174.700 74.200 ;
        RECT 175.800 74.100 176.200 74.200 ;
        RECT 175.400 73.800 176.200 74.100 ;
        RECT 168.700 73.300 170.600 73.600 ;
        RECT 168.700 73.200 169.100 73.300 ;
        RECT 163.000 72.100 163.400 72.500 ;
        RECT 163.800 72.400 164.200 72.800 ;
        RECT 164.700 72.700 165.100 72.800 ;
        RECT 164.700 72.400 166.100 72.700 ;
        RECT 165.800 72.100 166.100 72.400 ;
        RECT 167.800 72.100 168.200 72.500 ;
        RECT 163.000 71.800 164.000 72.100 ;
        RECT 163.600 71.100 164.000 71.800 ;
        RECT 165.800 71.100 166.200 72.100 ;
        RECT 167.800 71.800 168.500 72.100 ;
        RECT 167.900 71.100 168.500 71.800 ;
        RECT 170.200 71.100 170.600 73.300 ;
        RECT 171.000 73.400 172.100 73.700 ;
        RECT 171.000 71.100 171.400 73.400 ;
        RECT 173.500 73.100 173.800 73.800 ;
        RECT 175.400 73.600 175.800 73.800 ;
        RECT 177.600 73.700 177.900 74.500 ;
        RECT 178.400 74.200 178.700 75.900 ;
        RECT 179.800 75.800 180.200 76.200 ;
        RECT 178.200 73.800 178.700 74.200 ;
        RECT 179.900 74.200 180.200 75.800 ;
        RECT 182.200 75.400 182.600 76.200 ;
        RECT 183.800 76.100 184.200 79.900 ;
        RECT 185.400 77.500 185.800 79.500 ;
        RECT 187.500 79.200 187.900 79.900 ;
        RECT 187.000 78.800 187.900 79.200 ;
        RECT 183.000 75.800 184.200 76.100 ;
        RECT 184.600 75.800 185.000 76.600 ;
        RECT 185.400 75.800 185.700 77.500 ;
        RECT 187.500 76.400 187.900 78.800 ;
        RECT 192.900 79.200 193.300 79.900 ;
        RECT 192.900 78.800 193.800 79.200 ;
        RECT 192.200 76.800 192.600 77.200 ;
        RECT 187.500 76.100 188.300 76.400 ;
        RECT 192.200 76.200 192.500 76.800 ;
        RECT 192.900 76.200 193.300 78.800 ;
        RECT 183.000 75.200 183.300 75.800 ;
        RECT 181.000 74.800 181.800 75.200 ;
        RECT 183.000 74.800 183.400 75.200 ;
        RECT 179.900 74.100 180.700 74.200 ;
        RECT 179.900 73.900 180.800 74.100 ;
        RECT 176.600 73.400 177.900 73.700 ;
        RECT 174.300 73.100 176.100 73.300 ;
        RECT 173.400 71.100 173.800 73.100 ;
        RECT 174.200 73.000 176.200 73.100 ;
        RECT 174.200 71.100 174.600 73.000 ;
        RECT 175.800 71.100 176.200 73.000 ;
        RECT 176.600 71.100 177.000 73.400 ;
        RECT 178.400 73.100 178.700 73.800 ;
        RECT 178.200 72.800 178.700 73.100 ;
        RECT 178.200 71.100 178.600 72.800 ;
        RECT 180.400 71.100 180.800 73.900 ;
        RECT 183.000 73.400 183.400 74.200 ;
        RECT 183.800 73.100 184.200 75.800 ;
        RECT 185.400 75.500 187.300 75.800 ;
        RECT 185.400 74.400 185.800 75.200 ;
        RECT 186.200 74.400 186.600 75.200 ;
        RECT 187.000 74.500 187.300 75.500 ;
        RECT 187.000 74.100 187.700 74.500 ;
        RECT 188.000 74.200 188.300 76.100 ;
        RECT 191.800 75.900 192.500 76.200 ;
        RECT 192.800 75.900 193.300 76.200 ;
        RECT 191.800 75.800 192.200 75.900 ;
        RECT 188.600 74.800 189.000 75.600 ;
        RECT 192.800 74.200 193.100 75.900 ;
        RECT 193.400 74.400 193.800 75.200 ;
        RECT 187.000 73.900 187.500 74.100 ;
        RECT 185.400 73.600 187.500 73.900 ;
        RECT 188.000 73.800 189.000 74.200 ;
        RECT 191.800 73.800 193.100 74.200 ;
        RECT 194.200 74.100 194.600 74.200 ;
        RECT 195.000 74.100 195.400 79.900 ;
        RECT 198.500 76.400 198.900 79.900 ;
        RECT 200.600 77.500 201.000 79.500 ;
        RECT 198.100 76.100 198.900 76.400 ;
        RECT 196.600 75.100 197.000 75.200 ;
        RECT 197.400 75.100 197.800 75.600 ;
        RECT 196.600 74.800 197.800 75.100 ;
        RECT 198.100 74.200 198.400 76.100 ;
        RECT 200.700 75.800 201.000 77.500 ;
        RECT 203.300 76.400 203.700 79.900 ;
        RECT 205.400 77.500 205.800 79.500 ;
        RECT 199.100 75.500 201.000 75.800 ;
        RECT 202.900 76.100 203.700 76.400 ;
        RECT 199.100 74.500 199.400 75.500 ;
        RECT 193.800 73.800 195.400 74.100 ;
        RECT 197.400 73.800 198.400 74.200 ;
        RECT 198.700 74.100 199.400 74.500 ;
        RECT 199.800 74.400 200.200 75.200 ;
        RECT 200.600 74.400 201.000 75.200 ;
        RECT 202.200 74.800 202.600 75.600 ;
        RECT 202.900 74.200 203.200 76.100 ;
        RECT 205.500 75.800 205.800 77.500 ;
        RECT 203.900 75.500 205.800 75.800 ;
        RECT 206.200 75.600 206.600 79.900 ;
        RECT 208.300 77.900 208.900 79.900 ;
        RECT 210.600 77.900 211.000 79.900 ;
        RECT 212.800 78.200 213.200 79.900 ;
        RECT 212.800 77.900 213.800 78.200 ;
        RECT 208.600 77.500 209.000 77.900 ;
        RECT 210.700 77.600 211.000 77.900 ;
        RECT 210.300 77.300 212.100 77.600 ;
        RECT 213.400 77.500 213.800 77.900 ;
        RECT 210.300 77.200 210.700 77.300 ;
        RECT 211.700 77.200 212.100 77.300 ;
        RECT 208.200 76.600 208.900 77.000 ;
        RECT 208.600 76.100 208.900 76.600 ;
        RECT 209.700 76.500 210.800 76.800 ;
        RECT 209.700 76.400 210.100 76.500 ;
        RECT 208.600 75.800 209.800 76.100 ;
        RECT 203.900 74.500 204.200 75.500 ;
        RECT 206.200 75.300 208.300 75.600 ;
        RECT 183.800 72.800 184.700 73.100 ;
        RECT 184.300 71.100 184.700 72.800 ;
        RECT 185.400 72.500 185.700 73.600 ;
        RECT 188.000 73.500 188.300 73.800 ;
        RECT 187.900 73.300 188.300 73.500 ;
        RECT 187.500 73.000 188.300 73.300 ;
        RECT 191.900 73.100 192.200 73.800 ;
        RECT 193.800 73.600 194.200 73.800 ;
        RECT 192.700 73.100 194.500 73.300 ;
        RECT 185.400 71.500 185.800 72.500 ;
        RECT 187.500 71.500 187.900 73.000 ;
        RECT 191.800 71.100 192.200 73.100 ;
        RECT 192.600 73.000 194.600 73.100 ;
        RECT 192.600 71.100 193.000 73.000 ;
        RECT 194.200 71.100 194.600 73.000 ;
        RECT 195.000 71.100 195.400 73.800 ;
        RECT 198.100 73.500 198.400 73.800 ;
        RECT 198.900 73.900 199.400 74.100 ;
        RECT 201.400 74.100 201.800 74.200 ;
        RECT 202.200 74.100 203.200 74.200 ;
        RECT 203.500 74.100 204.200 74.500 ;
        RECT 204.600 74.400 205.000 75.200 ;
        RECT 205.400 74.400 205.800 75.200 ;
        RECT 198.900 73.600 201.000 73.900 ;
        RECT 201.400 73.800 203.200 74.100 ;
        RECT 198.100 73.300 198.500 73.500 ;
        RECT 195.800 72.400 196.200 73.200 ;
        RECT 198.100 73.000 198.900 73.300 ;
        RECT 198.500 71.500 198.900 73.000 ;
        RECT 200.700 72.500 201.000 73.600 ;
        RECT 202.900 73.500 203.200 73.800 ;
        RECT 203.700 73.900 204.200 74.100 ;
        RECT 203.700 73.600 205.800 73.900 ;
        RECT 202.900 73.300 203.300 73.500 ;
        RECT 202.900 73.000 203.700 73.300 ;
        RECT 200.600 71.500 201.000 72.500 ;
        RECT 203.300 71.500 203.700 73.000 ;
        RECT 205.500 72.500 205.800 73.600 ;
        RECT 205.400 71.500 205.800 72.500 ;
        RECT 206.200 73.600 206.600 75.300 ;
        RECT 207.900 75.200 208.300 75.300 ;
        RECT 207.100 74.900 207.500 75.000 ;
        RECT 207.100 74.600 209.000 74.900 ;
        RECT 208.600 74.500 209.000 74.600 ;
        RECT 209.500 74.200 209.800 75.800 ;
        RECT 210.500 75.900 210.800 76.500 ;
        RECT 211.100 76.500 211.500 76.600 ;
        RECT 213.400 76.500 213.800 76.600 ;
        RECT 211.100 76.200 213.800 76.500 ;
        RECT 210.500 75.700 212.900 75.900 ;
        RECT 215.000 75.700 215.400 79.900 ;
        RECT 210.500 75.600 215.400 75.700 ;
        RECT 212.500 75.500 215.400 75.600 ;
        RECT 212.600 75.400 215.400 75.500 ;
        RECT 211.800 75.100 212.200 75.200 ;
        RECT 216.600 75.100 217.000 79.900 ;
        RECT 218.600 76.800 219.000 77.200 ;
        RECT 217.400 75.800 217.800 76.600 ;
        RECT 218.600 76.200 218.900 76.800 ;
        RECT 219.300 76.200 219.700 79.900 ;
        RECT 218.200 75.900 218.900 76.200 ;
        RECT 219.200 75.900 219.700 76.200 ;
        RECT 218.200 75.800 218.600 75.900 ;
        RECT 218.200 75.100 218.500 75.800 ;
        RECT 211.800 74.800 214.300 75.100 ;
        RECT 212.600 74.700 213.000 74.800 ;
        RECT 213.900 74.700 214.300 74.800 ;
        RECT 216.600 74.800 218.500 75.100 ;
        RECT 213.100 74.200 213.500 74.300 ;
        RECT 209.500 73.900 215.000 74.200 ;
        RECT 209.700 73.800 210.100 73.900 ;
        RECT 206.200 73.300 208.100 73.600 ;
        RECT 206.200 71.100 206.600 73.300 ;
        RECT 207.700 73.200 208.100 73.300 ;
        RECT 212.600 72.800 212.900 73.900 ;
        RECT 214.200 73.800 215.000 73.900 ;
        RECT 211.700 72.700 212.100 72.800 ;
        RECT 208.600 72.100 209.000 72.500 ;
        RECT 210.700 72.400 212.100 72.700 ;
        RECT 212.600 72.400 213.000 72.800 ;
        RECT 210.700 72.100 211.000 72.400 ;
        RECT 213.400 72.100 213.800 72.500 ;
        RECT 208.300 71.800 209.000 72.100 ;
        RECT 208.300 71.100 208.900 71.800 ;
        RECT 210.600 71.100 211.000 72.100 ;
        RECT 212.800 71.800 213.800 72.100 ;
        RECT 212.800 71.100 213.200 71.800 ;
        RECT 215.000 71.100 215.400 73.500 ;
        RECT 215.800 73.400 216.200 74.200 ;
        RECT 216.600 73.100 217.000 74.800 ;
        RECT 219.200 74.200 219.500 75.900 ;
        RECT 222.200 75.600 222.600 79.900 ;
        RECT 223.800 75.600 224.200 79.900 ;
        RECT 225.400 75.600 225.800 79.900 ;
        RECT 227.000 75.600 227.400 79.900 ;
        RECT 228.600 76.200 229.000 79.900 ;
        RECT 228.600 75.900 229.700 76.200 ;
        RECT 229.400 75.600 229.700 75.900 ;
        RECT 222.200 75.200 223.100 75.600 ;
        RECT 223.800 75.200 224.900 75.600 ;
        RECT 225.400 75.200 226.500 75.600 ;
        RECT 227.000 75.200 228.200 75.600 ;
        RECT 229.400 75.200 230.000 75.600 ;
        RECT 219.800 74.400 220.200 75.200 ;
        RECT 222.700 74.500 223.100 75.200 ;
        RECT 224.500 74.500 224.900 75.200 ;
        RECT 226.100 74.500 226.500 75.200 ;
        RECT 217.400 74.100 217.800 74.200 ;
        RECT 218.200 74.100 219.500 74.200 ;
        RECT 220.600 74.100 221.000 74.200 ;
        RECT 217.400 73.800 219.500 74.100 ;
        RECT 220.200 73.800 221.000 74.100 ;
        RECT 222.700 74.100 224.000 74.500 ;
        RECT 224.500 74.100 225.700 74.500 ;
        RECT 226.100 74.100 227.400 74.500 ;
        RECT 222.700 73.800 223.100 74.100 ;
        RECT 224.500 73.800 224.900 74.100 ;
        RECT 226.100 73.800 226.500 74.100 ;
        RECT 227.800 73.800 228.200 75.200 ;
        RECT 228.600 74.400 229.000 75.200 ;
        RECT 218.300 73.100 218.600 73.800 ;
        RECT 220.200 73.600 220.600 73.800 ;
        RECT 222.200 73.400 223.100 73.800 ;
        RECT 223.800 73.400 224.900 73.800 ;
        RECT 225.400 73.400 226.500 73.800 ;
        RECT 227.000 73.400 228.200 73.800 ;
        RECT 229.400 73.700 229.700 75.200 ;
        RECT 228.600 73.400 229.700 73.700 ;
        RECT 219.100 73.100 220.900 73.300 ;
        RECT 216.600 72.800 217.500 73.100 ;
        RECT 217.100 71.100 217.500 72.800 ;
        RECT 218.200 71.100 218.600 73.100 ;
        RECT 219.000 73.000 221.000 73.100 ;
        RECT 219.000 71.100 219.400 73.000 ;
        RECT 220.600 71.100 221.000 73.000 ;
        RECT 222.200 71.100 222.600 73.400 ;
        RECT 223.800 71.100 224.200 73.400 ;
        RECT 225.400 71.100 225.800 73.400 ;
        RECT 227.000 71.100 227.400 73.400 ;
        RECT 228.600 71.100 229.000 73.400 ;
        RECT 1.400 67.600 1.800 69.900 ;
        RECT 3.000 67.600 3.400 69.900 ;
        RECT 1.400 67.200 3.400 67.600 ;
        RECT 4.600 67.500 5.000 69.900 ;
        RECT 6.800 69.200 7.200 69.900 ;
        RECT 6.200 68.900 7.200 69.200 ;
        RECT 9.000 68.900 9.400 69.900 ;
        RECT 11.100 69.200 11.700 69.900 ;
        RECT 11.000 68.900 11.700 69.200 ;
        RECT 6.200 68.500 6.600 68.900 ;
        RECT 9.000 68.600 9.300 68.900 ;
        RECT 7.000 68.200 7.400 68.600 ;
        RECT 7.900 68.300 9.300 68.600 ;
        RECT 11.000 68.500 11.400 68.900 ;
        RECT 7.900 68.200 8.300 68.300 ;
        RECT 3.000 65.800 3.400 67.200 ;
        RECT 5.000 67.100 5.800 67.200 ;
        RECT 7.100 67.100 7.400 68.200 ;
        RECT 11.900 67.700 12.300 67.800 ;
        RECT 13.400 67.700 13.800 69.900 ;
        RECT 14.200 67.900 14.600 69.900 ;
        RECT 15.000 68.000 15.400 69.900 ;
        RECT 16.600 68.000 17.000 69.900 ;
        RECT 15.000 67.900 17.000 68.000 ;
        RECT 11.900 67.400 13.800 67.700 ;
        RECT 7.800 67.100 8.200 67.200 ;
        RECT 9.900 67.100 10.300 67.200 ;
        RECT 5.000 66.800 10.500 67.100 ;
        RECT 6.500 66.700 6.900 66.800 ;
        RECT 5.700 66.200 6.100 66.300 ;
        RECT 5.700 66.100 8.200 66.200 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 5.700 65.900 9.000 66.100 ;
        RECT 7.800 65.800 9.000 65.900 ;
        RECT 1.400 65.400 3.400 65.800 ;
        RECT 1.400 61.100 1.800 65.400 ;
        RECT 3.000 61.100 3.400 65.400 ;
        RECT 4.600 65.500 7.400 65.600 ;
        RECT 4.600 65.400 7.500 65.500 ;
        RECT 4.600 65.300 9.500 65.400 ;
        RECT 4.600 61.100 5.000 65.300 ;
        RECT 7.100 65.100 9.500 65.300 ;
        RECT 6.200 64.500 8.900 64.800 ;
        RECT 6.200 64.400 6.600 64.500 ;
        RECT 8.500 64.400 8.900 64.500 ;
        RECT 9.200 64.500 9.500 65.100 ;
        RECT 10.200 65.200 10.500 66.800 ;
        RECT 11.000 66.400 11.400 66.500 ;
        RECT 11.000 66.100 12.900 66.400 ;
        RECT 12.500 66.000 12.900 66.100 ;
        RECT 11.700 65.700 12.100 65.800 ;
        RECT 13.400 65.700 13.800 67.400 ;
        RECT 14.300 67.200 14.600 67.900 ;
        RECT 15.100 67.700 16.900 67.900 ;
        RECT 17.400 67.800 17.800 68.600 ;
        RECT 16.200 67.200 16.600 67.400 ;
        RECT 17.400 67.200 17.700 67.800 ;
        RECT 14.200 66.800 15.500 67.200 ;
        RECT 16.200 66.900 17.000 67.200 ;
        RECT 16.600 66.800 17.000 66.900 ;
        RECT 17.400 66.800 17.800 67.200 ;
        RECT 18.200 67.100 18.600 69.900 ;
        RECT 19.000 68.000 19.400 69.900 ;
        RECT 20.600 68.000 21.000 69.900 ;
        RECT 19.000 67.900 21.000 68.000 ;
        RECT 21.400 67.900 21.800 69.900 ;
        RECT 19.100 67.700 20.900 67.900 ;
        RECT 19.400 67.200 19.800 67.400 ;
        RECT 21.400 67.200 21.700 67.900 ;
        RECT 22.200 67.500 22.600 69.900 ;
        RECT 24.400 69.200 24.800 69.900 ;
        RECT 23.800 68.900 24.800 69.200 ;
        RECT 26.600 68.900 27.000 69.900 ;
        RECT 28.700 69.200 29.300 69.900 ;
        RECT 28.600 68.900 29.300 69.200 ;
        RECT 23.800 68.500 24.200 68.900 ;
        RECT 26.600 68.600 26.900 68.900 ;
        RECT 24.600 68.200 25.000 68.600 ;
        RECT 25.500 68.300 26.900 68.600 ;
        RECT 28.600 68.500 29.000 68.900 ;
        RECT 25.500 68.200 25.900 68.300 ;
        RECT 19.000 67.100 19.800 67.200 ;
        RECT 18.200 66.900 19.800 67.100 ;
        RECT 18.200 66.800 19.400 66.900 ;
        RECT 20.500 66.800 21.800 67.200 ;
        RECT 22.600 67.100 23.400 67.200 ;
        RECT 24.700 67.100 25.000 68.200 ;
        RECT 29.500 67.700 29.900 67.800 ;
        RECT 31.000 67.700 31.400 69.900 ;
        RECT 31.800 68.000 32.200 69.900 ;
        RECT 33.400 68.000 33.800 69.900 ;
        RECT 31.800 67.900 33.800 68.000 ;
        RECT 34.200 67.900 34.600 69.900 ;
        RECT 35.800 68.200 36.200 69.900 ;
        RECT 31.900 67.700 33.700 67.900 ;
        RECT 29.500 67.400 31.400 67.700 ;
        RECT 27.500 67.100 27.900 67.200 ;
        RECT 22.600 66.800 28.100 67.100 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 15.200 66.100 15.500 66.800 ;
        RECT 14.200 65.800 15.500 66.100 ;
        RECT 15.800 65.800 16.200 66.600 ;
        RECT 11.700 65.400 13.800 65.700 ;
        RECT 10.200 64.900 11.400 65.200 ;
        RECT 9.900 64.500 10.300 64.600 ;
        RECT 9.200 64.200 10.300 64.500 ;
        RECT 11.100 64.400 11.400 64.900 ;
        RECT 11.100 64.000 11.800 64.400 ;
        RECT 7.900 63.700 8.300 63.800 ;
        RECT 9.300 63.700 9.700 63.800 ;
        RECT 6.200 63.100 6.600 63.500 ;
        RECT 7.900 63.400 9.700 63.700 ;
        RECT 9.000 63.100 9.300 63.400 ;
        RECT 11.000 63.100 11.400 63.500 ;
        RECT 6.200 62.800 7.200 63.100 ;
        RECT 6.800 61.100 7.200 62.800 ;
        RECT 9.000 61.100 9.400 63.100 ;
        RECT 11.100 61.100 11.700 63.100 ;
        RECT 13.400 61.100 13.800 65.400 ;
        RECT 14.200 65.100 14.600 65.200 ;
        RECT 15.200 65.100 15.500 65.800 ;
        RECT 14.200 64.800 14.900 65.100 ;
        RECT 15.200 64.800 15.700 65.100 ;
        RECT 14.600 64.200 14.900 64.800 ;
        RECT 14.600 63.800 15.000 64.200 ;
        RECT 15.300 61.100 15.700 64.800 ;
        RECT 18.200 61.100 18.600 66.800 ;
        RECT 19.800 65.800 20.200 66.600 ;
        RECT 20.500 65.100 20.800 66.800 ;
        RECT 21.400 66.200 21.700 66.800 ;
        RECT 24.100 66.700 24.500 66.800 ;
        RECT 23.300 66.200 23.700 66.300 ;
        RECT 21.400 65.800 21.800 66.200 ;
        RECT 23.300 65.900 25.800 66.200 ;
        RECT 25.400 65.800 25.800 65.900 ;
        RECT 27.000 66.100 27.400 66.200 ;
        RECT 27.800 66.100 28.100 66.800 ;
        RECT 28.600 66.400 29.000 66.500 ;
        RECT 28.600 66.100 30.500 66.400 ;
        RECT 27.000 65.800 28.100 66.100 ;
        RECT 30.100 66.000 30.500 66.100 ;
        RECT 22.200 65.500 25.000 65.600 ;
        RECT 22.200 65.400 25.100 65.500 ;
        RECT 22.200 65.300 27.100 65.400 ;
        RECT 21.400 65.100 21.800 65.200 ;
        RECT 20.300 64.800 20.800 65.100 ;
        RECT 21.100 64.800 21.800 65.100 ;
        RECT 20.300 61.100 20.700 64.800 ;
        RECT 21.100 64.200 21.400 64.800 ;
        RECT 21.000 63.800 21.400 64.200 ;
        RECT 22.200 61.100 22.600 65.300 ;
        RECT 24.700 65.100 27.100 65.300 ;
        RECT 23.800 64.500 26.500 64.800 ;
        RECT 23.800 64.400 24.200 64.500 ;
        RECT 26.100 64.400 26.500 64.500 ;
        RECT 26.800 64.500 27.100 65.100 ;
        RECT 27.800 65.200 28.100 65.800 ;
        RECT 29.300 65.700 29.700 65.800 ;
        RECT 31.000 65.700 31.400 67.400 ;
        RECT 32.200 67.200 32.600 67.400 ;
        RECT 34.200 67.200 34.500 67.900 ;
        RECT 35.700 67.800 36.200 68.200 ;
        RECT 35.700 67.200 36.000 67.800 ;
        RECT 37.400 67.600 37.800 69.900 ;
        RECT 39.800 67.900 40.200 69.900 ;
        RECT 40.600 68.000 41.000 69.900 ;
        RECT 42.200 68.000 42.600 69.900 ;
        RECT 40.600 67.900 42.600 68.000 ;
        RECT 36.500 67.300 37.800 67.600 ;
        RECT 31.800 66.900 32.600 67.200 ;
        RECT 33.300 67.100 34.600 67.200 ;
        RECT 31.800 66.800 32.200 66.900 ;
        RECT 33.300 66.800 35.300 67.100 ;
        RECT 32.600 65.800 33.000 66.600 ;
        RECT 29.300 65.400 31.400 65.700 ;
        RECT 27.800 64.900 29.000 65.200 ;
        RECT 27.500 64.500 27.900 64.600 ;
        RECT 26.800 64.200 27.900 64.500 ;
        RECT 28.700 64.400 29.000 64.900 ;
        RECT 28.700 64.000 29.400 64.400 ;
        RECT 25.500 63.700 25.900 63.800 ;
        RECT 26.900 63.700 27.300 63.800 ;
        RECT 23.800 63.100 24.200 63.500 ;
        RECT 25.500 63.400 27.300 63.700 ;
        RECT 26.600 63.100 26.900 63.400 ;
        RECT 28.600 63.100 29.000 63.500 ;
        RECT 23.800 62.800 24.800 63.100 ;
        RECT 24.400 61.100 24.800 62.800 ;
        RECT 26.600 61.100 27.000 63.100 ;
        RECT 28.700 61.100 29.300 63.100 ;
        RECT 31.000 61.100 31.400 65.400 ;
        RECT 33.300 65.100 33.600 66.800 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 35.700 66.800 36.200 67.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 34.200 65.100 34.600 65.200 ;
        RECT 33.100 64.800 33.600 65.100 ;
        RECT 33.900 64.800 34.600 65.100 ;
        RECT 35.700 65.100 36.000 66.800 ;
        RECT 36.500 66.500 36.800 67.300 ;
        RECT 39.900 67.200 40.200 67.900 ;
        RECT 40.700 67.700 42.500 67.900 ;
        RECT 43.000 67.600 43.400 69.900 ;
        RECT 44.600 68.200 45.000 69.900 ;
        RECT 47.500 68.200 47.900 69.900 ;
        RECT 49.900 69.200 50.300 69.900 ;
        RECT 49.900 68.800 50.600 69.200 ;
        RECT 49.900 68.200 50.300 68.800 ;
        RECT 44.600 67.900 45.100 68.200 ;
        RECT 41.800 67.200 42.200 67.400 ;
        RECT 43.000 67.300 44.300 67.600 ;
        RECT 39.800 66.800 41.100 67.200 ;
        RECT 41.800 66.900 42.600 67.200 ;
        RECT 42.200 66.800 42.600 66.900 ;
        RECT 36.300 66.100 36.800 66.500 ;
        RECT 36.500 65.100 36.800 66.100 ;
        RECT 37.300 66.200 37.700 66.600 ;
        RECT 37.300 65.800 37.800 66.200 ;
        RECT 39.800 65.100 40.200 65.200 ;
        RECT 40.800 65.100 41.100 66.800 ;
        RECT 41.400 65.800 41.800 66.600 ;
        RECT 43.100 66.200 43.500 66.600 ;
        RECT 43.000 65.800 43.500 66.200 ;
        RECT 44.000 66.500 44.300 67.300 ;
        RECT 44.800 67.200 45.100 67.900 ;
        RECT 47.000 67.900 47.900 68.200 ;
        RECT 49.400 67.900 50.300 68.200 ;
        RECT 44.600 66.800 45.100 67.200 ;
        RECT 46.200 66.800 46.600 67.600 ;
        RECT 44.000 66.100 44.500 66.500 ;
        RECT 44.000 65.100 44.300 66.100 ;
        RECT 44.800 65.100 45.100 66.800 ;
        RECT 33.100 61.100 33.500 64.800 ;
        RECT 33.900 64.200 34.200 64.800 ;
        RECT 35.700 64.600 36.200 65.100 ;
        RECT 36.500 64.800 37.800 65.100 ;
        RECT 39.800 64.800 40.500 65.100 ;
        RECT 40.800 64.800 41.300 65.100 ;
        RECT 33.800 63.800 34.200 64.200 ;
        RECT 35.800 61.100 36.200 64.600 ;
        RECT 37.400 61.100 37.800 64.800 ;
        RECT 40.200 64.200 40.500 64.800 ;
        RECT 40.200 63.800 40.600 64.200 ;
        RECT 40.900 61.100 41.300 64.800 ;
        RECT 43.000 64.800 44.300 65.100 ;
        RECT 43.000 61.100 43.400 64.800 ;
        RECT 44.600 64.600 45.100 65.100 ;
        RECT 44.600 61.100 45.000 64.600 ;
        RECT 47.000 61.100 47.400 67.900 ;
        RECT 48.600 66.800 49.000 67.600 ;
        RECT 47.800 65.100 48.200 65.200 ;
        RECT 48.600 65.100 49.000 65.200 ;
        RECT 47.800 64.800 49.000 65.100 ;
        RECT 47.800 64.400 48.200 64.800 ;
        RECT 49.400 61.100 49.800 67.900 ;
        RECT 51.000 67.500 51.400 69.900 ;
        RECT 53.200 69.200 53.600 69.900 ;
        RECT 52.600 68.900 53.600 69.200 ;
        RECT 55.400 68.900 55.800 69.900 ;
        RECT 57.500 69.200 58.100 69.900 ;
        RECT 57.400 68.900 58.100 69.200 ;
        RECT 52.600 68.500 53.000 68.900 ;
        RECT 55.400 68.600 55.700 68.900 ;
        RECT 53.400 68.200 53.800 68.600 ;
        RECT 54.300 68.300 55.700 68.600 ;
        RECT 57.400 68.500 57.800 68.900 ;
        RECT 54.300 68.200 54.700 68.300 ;
        RECT 51.400 67.100 52.200 67.200 ;
        RECT 53.500 67.100 53.800 68.200 ;
        RECT 58.300 67.700 58.700 67.800 ;
        RECT 59.800 67.700 60.200 69.900 ;
        RECT 60.900 68.200 61.300 69.900 ;
        RECT 64.300 68.200 64.700 69.900 ;
        RECT 66.700 69.200 67.100 69.900 ;
        RECT 66.700 68.800 67.400 69.200 ;
        RECT 66.700 68.200 67.100 68.800 ;
        RECT 60.900 67.900 61.800 68.200 ;
        RECT 58.300 67.400 60.200 67.700 ;
        RECT 56.300 67.100 56.700 67.200 ;
        RECT 51.400 66.800 56.900 67.100 ;
        RECT 52.900 66.700 53.300 66.800 ;
        RECT 52.100 66.200 52.500 66.300 ;
        RECT 53.400 66.200 53.800 66.300 ;
        RECT 56.600 66.200 56.900 66.800 ;
        RECT 57.400 66.400 57.800 66.500 ;
        RECT 52.100 65.900 54.600 66.200 ;
        RECT 54.200 65.800 54.600 65.900 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 57.400 66.100 59.300 66.400 ;
        RECT 58.900 66.000 59.300 66.100 ;
        RECT 51.000 65.500 53.800 65.600 ;
        RECT 51.000 65.400 53.900 65.500 ;
        RECT 51.000 65.300 55.900 65.400 ;
        RECT 50.200 63.800 50.600 65.200 ;
        RECT 51.000 61.100 51.400 65.300 ;
        RECT 53.500 65.100 55.900 65.300 ;
        RECT 52.600 64.500 55.300 64.800 ;
        RECT 52.600 64.400 53.000 64.500 ;
        RECT 54.900 64.400 55.300 64.500 ;
        RECT 55.600 64.500 55.900 65.100 ;
        RECT 56.600 65.200 56.900 65.800 ;
        RECT 58.100 65.700 58.500 65.800 ;
        RECT 59.800 65.700 60.200 67.400 ;
        RECT 58.100 65.400 60.200 65.700 ;
        RECT 56.600 64.900 57.800 65.200 ;
        RECT 56.300 64.500 56.700 64.600 ;
        RECT 55.600 64.200 56.700 64.500 ;
        RECT 57.500 64.400 57.800 64.900 ;
        RECT 57.500 64.000 58.200 64.400 ;
        RECT 54.300 63.700 54.700 63.800 ;
        RECT 55.700 63.700 56.100 63.800 ;
        RECT 52.600 63.100 53.000 63.500 ;
        RECT 54.300 63.400 56.100 63.700 ;
        RECT 55.400 63.100 55.700 63.400 ;
        RECT 57.400 63.100 57.800 63.500 ;
        RECT 52.600 62.800 53.600 63.100 ;
        RECT 53.200 61.100 53.600 62.800 ;
        RECT 55.400 61.100 55.800 63.100 ;
        RECT 57.500 61.100 58.100 63.100 ;
        RECT 59.800 61.100 60.200 65.400 ;
        RECT 60.600 64.400 61.000 65.200 ;
        RECT 61.400 61.100 61.800 67.900 ;
        RECT 63.800 67.900 64.700 68.200 ;
        RECT 66.200 67.900 67.100 68.200 ;
        RECT 67.800 68.500 68.200 69.500 ;
        RECT 62.200 66.800 62.600 67.600 ;
        RECT 63.000 66.800 63.400 67.600 ;
        RECT 63.800 67.100 64.200 67.900 ;
        RECT 63.800 66.800 64.900 67.100 ;
        RECT 65.400 66.800 65.800 67.600 ;
        RECT 63.800 61.100 64.200 66.800 ;
        RECT 64.600 66.200 64.900 66.800 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 64.600 64.400 65.000 65.200 ;
        RECT 66.200 61.100 66.600 67.900 ;
        RECT 67.800 67.400 68.100 68.500 ;
        RECT 69.900 68.000 70.300 69.500 ;
        RECT 72.600 68.000 73.000 69.900 ;
        RECT 74.200 68.000 74.600 69.900 ;
        RECT 69.900 67.700 70.700 68.000 ;
        RECT 72.600 67.900 74.600 68.000 ;
        RECT 75.000 67.900 75.400 69.900 ;
        RECT 76.100 68.200 76.500 69.900 ;
        RECT 76.100 67.900 77.000 68.200 ;
        RECT 72.700 67.700 74.500 67.900 ;
        RECT 70.300 67.500 70.700 67.700 ;
        RECT 67.800 67.100 69.900 67.400 ;
        RECT 69.400 66.900 69.900 67.100 ;
        RECT 70.400 67.200 70.700 67.500 ;
        RECT 73.000 67.200 73.400 67.400 ;
        RECT 75.000 67.200 75.300 67.900 ;
        RECT 67.800 65.800 68.200 66.600 ;
        RECT 68.600 65.800 69.000 66.600 ;
        RECT 69.400 66.500 70.100 66.900 ;
        RECT 70.400 66.800 71.400 67.200 ;
        RECT 72.600 66.900 73.400 67.200 ;
        RECT 72.600 66.800 73.000 66.900 ;
        RECT 74.100 66.800 75.400 67.200 ;
        RECT 69.400 65.500 69.700 66.500 ;
        RECT 67.800 65.200 69.700 65.500 ;
        RECT 67.000 63.800 67.400 65.200 ;
        RECT 67.800 63.500 68.100 65.200 ;
        RECT 70.400 64.900 70.700 66.800 ;
        RECT 71.000 65.400 71.400 66.200 ;
        RECT 73.400 65.800 73.800 66.600 ;
        RECT 74.100 65.100 74.400 66.800 ;
        RECT 76.600 66.100 77.000 67.900 ;
        RECT 77.400 66.800 77.800 67.600 ;
        RECT 78.200 67.500 78.600 69.900 ;
        RECT 80.400 69.200 80.800 69.900 ;
        RECT 79.800 68.900 80.800 69.200 ;
        RECT 82.600 68.900 83.000 69.900 ;
        RECT 84.700 69.200 85.300 69.900 ;
        RECT 84.600 68.900 85.300 69.200 ;
        RECT 87.000 69.100 87.400 69.900 ;
        RECT 87.800 69.100 88.200 69.200 ;
        RECT 79.800 68.500 80.200 68.900 ;
        RECT 82.600 68.600 82.900 68.900 ;
        RECT 80.600 68.200 81.000 68.600 ;
        RECT 81.500 68.300 82.900 68.600 ;
        RECT 84.600 68.500 85.000 68.900 ;
        RECT 87.000 68.800 88.200 69.100 ;
        RECT 81.500 68.200 81.900 68.300 ;
        RECT 78.600 67.100 79.400 67.200 ;
        RECT 80.700 67.100 81.000 68.200 ;
        RECT 85.500 67.700 85.900 67.800 ;
        RECT 87.000 67.700 87.400 68.800 ;
        RECT 91.300 68.000 91.700 69.500 ;
        RECT 93.400 68.500 93.800 69.500 ;
        RECT 85.500 67.400 87.400 67.700 ;
        RECT 82.200 67.100 82.600 67.200 ;
        RECT 83.500 67.100 83.900 67.200 ;
        RECT 78.600 66.800 84.100 67.100 ;
        RECT 80.100 66.700 80.500 66.800 ;
        RECT 75.000 65.800 77.000 66.100 ;
        RECT 79.300 66.200 79.700 66.300 ;
        RECT 80.600 66.200 81.000 66.300 ;
        RECT 79.300 65.900 81.800 66.200 ;
        RECT 81.400 65.800 81.800 65.900 ;
        RECT 75.000 65.200 75.300 65.800 ;
        RECT 75.000 65.100 75.400 65.200 ;
        RECT 69.900 64.600 70.700 64.900 ;
        RECT 73.900 64.800 74.400 65.100 ;
        RECT 74.700 64.800 75.400 65.100 ;
        RECT 67.800 61.500 68.200 63.500 ;
        RECT 69.900 62.200 70.300 64.600 ;
        RECT 69.900 61.800 70.600 62.200 ;
        RECT 69.900 61.100 70.300 61.800 ;
        RECT 73.900 61.100 74.300 64.800 ;
        RECT 74.700 64.200 75.000 64.800 ;
        RECT 75.800 64.400 76.200 65.200 ;
        RECT 74.600 63.800 75.000 64.200 ;
        RECT 76.600 61.100 77.000 65.800 ;
        RECT 78.200 65.500 81.000 65.600 ;
        RECT 78.200 65.400 81.100 65.500 ;
        RECT 78.200 65.300 83.100 65.400 ;
        RECT 78.200 61.100 78.600 65.300 ;
        RECT 80.700 65.100 83.100 65.300 ;
        RECT 79.800 64.500 82.500 64.800 ;
        RECT 79.800 64.400 80.200 64.500 ;
        RECT 82.100 64.400 82.500 64.500 ;
        RECT 82.800 64.500 83.100 65.100 ;
        RECT 83.800 65.200 84.100 66.800 ;
        RECT 84.600 66.400 85.000 66.500 ;
        RECT 84.600 66.100 86.500 66.400 ;
        RECT 86.100 66.000 86.500 66.100 ;
        RECT 85.300 65.700 85.700 65.800 ;
        RECT 87.000 65.700 87.400 67.400 ;
        RECT 90.900 67.700 91.700 68.000 ;
        RECT 90.900 67.500 91.300 67.700 ;
        RECT 90.900 67.200 91.200 67.500 ;
        RECT 93.500 67.400 93.800 68.500 ;
        RECT 94.500 69.200 94.900 69.900 ;
        RECT 94.500 68.800 95.400 69.200 ;
        RECT 94.500 68.200 94.900 68.800 ;
        RECT 94.500 67.900 95.400 68.200 ;
        RECT 96.600 67.900 97.000 69.900 ;
        RECT 97.400 68.000 97.800 69.900 ;
        RECT 99.000 68.000 99.400 69.900 ;
        RECT 97.400 67.900 99.400 68.000 ;
        RECT 101.400 67.900 101.800 69.900 ;
        RECT 102.100 68.200 102.500 68.600 ;
        RECT 90.200 66.800 91.200 67.200 ;
        RECT 91.700 67.100 93.800 67.400 ;
        RECT 91.700 66.900 92.200 67.100 ;
        RECT 87.800 66.100 88.200 66.200 ;
        RECT 90.200 66.100 90.600 66.200 ;
        RECT 87.800 65.800 90.600 66.100 ;
        RECT 85.300 65.400 87.400 65.700 ;
        RECT 90.200 65.400 90.600 65.800 ;
        RECT 83.800 64.900 85.000 65.200 ;
        RECT 83.500 64.500 83.900 64.600 ;
        RECT 82.800 64.200 83.900 64.500 ;
        RECT 84.700 64.400 85.000 64.900 ;
        RECT 84.700 64.000 85.400 64.400 ;
        RECT 81.500 63.700 81.900 63.800 ;
        RECT 82.900 63.700 83.300 63.800 ;
        RECT 79.800 63.100 80.200 63.500 ;
        RECT 81.500 63.400 83.300 63.700 ;
        RECT 82.600 63.100 82.900 63.400 ;
        RECT 84.600 63.100 85.000 63.500 ;
        RECT 79.800 62.800 80.800 63.100 ;
        RECT 80.400 61.100 80.800 62.800 ;
        RECT 82.600 61.100 83.000 63.100 ;
        RECT 84.700 61.100 85.300 63.100 ;
        RECT 87.000 61.100 87.400 65.400 ;
        RECT 90.900 64.900 91.200 66.800 ;
        RECT 91.500 66.500 92.200 66.900 ;
        RECT 91.900 65.500 92.200 66.500 ;
        RECT 92.600 65.800 93.000 66.600 ;
        RECT 93.400 65.800 93.800 66.600 ;
        RECT 91.900 65.200 93.800 65.500 ;
        RECT 90.900 64.600 91.700 64.900 ;
        RECT 91.300 62.200 91.700 64.600 ;
        RECT 93.500 63.500 93.800 65.200 ;
        RECT 94.200 64.400 94.600 65.200 ;
        RECT 91.300 61.800 92.200 62.200 ;
        RECT 91.300 61.100 91.700 61.800 ;
        RECT 93.400 61.500 93.800 63.500 ;
        RECT 95.000 61.100 95.400 67.900 ;
        RECT 95.800 66.800 96.200 67.600 ;
        RECT 96.700 67.200 97.000 67.900 ;
        RECT 97.500 67.700 99.300 67.900 ;
        RECT 98.600 67.200 99.000 67.400 ;
        RECT 96.600 66.800 97.900 67.200 ;
        RECT 98.600 66.900 99.400 67.200 ;
        RECT 99.000 66.800 99.400 66.900 ;
        RECT 97.600 65.200 97.900 66.800 ;
        RECT 98.200 65.800 98.600 66.600 ;
        RECT 100.600 66.400 101.000 67.200 ;
        RECT 99.000 66.100 99.400 66.200 ;
        RECT 99.800 66.100 100.200 66.200 ;
        RECT 101.400 66.100 101.700 67.900 ;
        RECT 102.200 67.800 102.600 68.200 ;
        RECT 103.000 67.900 103.400 69.900 ;
        RECT 103.800 68.000 104.200 69.900 ;
        RECT 105.400 68.000 105.800 69.900 ;
        RECT 103.800 67.900 105.800 68.000 ;
        RECT 106.200 68.000 106.600 69.900 ;
        RECT 107.800 68.000 108.200 69.900 ;
        RECT 106.200 67.900 108.200 68.000 ;
        RECT 108.600 67.900 109.000 69.900 ;
        RECT 109.700 69.200 110.100 69.900 ;
        RECT 113.100 69.200 113.500 69.900 ;
        RECT 109.400 68.800 110.100 69.200 ;
        RECT 112.600 68.800 113.500 69.200 ;
        RECT 109.700 68.200 110.100 68.800 ;
        RECT 113.100 68.200 113.500 68.800 ;
        RECT 115.500 68.200 115.900 69.900 ;
        RECT 109.700 67.900 110.600 68.200 ;
        RECT 103.100 67.200 103.400 67.900 ;
        RECT 103.900 67.700 105.700 67.900 ;
        RECT 106.300 67.700 108.100 67.900 ;
        RECT 105.000 67.200 105.400 67.400 ;
        RECT 106.600 67.200 107.000 67.400 ;
        RECT 108.600 67.200 108.900 67.900 ;
        RECT 102.200 67.100 102.600 67.200 ;
        RECT 103.000 67.100 104.300 67.200 ;
        RECT 102.200 66.800 104.300 67.100 ;
        RECT 105.000 66.900 105.800 67.200 ;
        RECT 105.400 66.800 105.800 66.900 ;
        RECT 106.200 66.900 107.000 67.200 ;
        RECT 106.200 66.800 106.600 66.900 ;
        RECT 107.700 66.800 109.000 67.200 ;
        RECT 102.200 66.100 102.600 66.200 ;
        RECT 103.000 66.100 103.400 66.200 ;
        RECT 99.000 65.800 100.600 66.100 ;
        RECT 101.400 65.800 103.400 66.100 ;
        RECT 100.200 65.600 100.600 65.800 ;
        RECT 95.800 65.100 96.200 65.200 ;
        RECT 96.600 65.100 97.000 65.200 ;
        RECT 95.800 64.800 97.300 65.100 ;
        RECT 97.600 64.800 98.600 65.200 ;
        RECT 102.200 65.100 102.500 65.800 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 104.000 65.100 104.300 66.800 ;
        RECT 104.600 65.800 105.000 66.600 ;
        RECT 107.000 65.800 107.400 66.600 ;
        RECT 107.700 65.100 108.000 66.800 ;
        RECT 108.600 65.100 109.000 65.200 ;
        RECT 99.800 64.800 101.800 65.100 ;
        RECT 97.000 64.200 97.300 64.800 ;
        RECT 97.000 63.800 97.400 64.200 ;
        RECT 97.700 61.100 98.100 64.800 ;
        RECT 99.800 61.100 100.200 64.800 ;
        RECT 101.400 61.100 101.800 64.800 ;
        RECT 102.200 61.100 102.600 65.100 ;
        RECT 103.000 64.800 103.700 65.100 ;
        RECT 104.000 64.800 104.500 65.100 ;
        RECT 103.400 64.200 103.700 64.800 ;
        RECT 103.400 63.800 103.800 64.200 ;
        RECT 104.100 61.100 104.500 64.800 ;
        RECT 107.500 64.800 108.000 65.100 ;
        RECT 108.300 64.800 109.000 65.100 ;
        RECT 107.500 61.100 107.900 64.800 ;
        RECT 108.300 64.200 108.600 64.800 ;
        RECT 109.400 64.400 109.800 65.200 ;
        RECT 108.200 63.800 108.600 64.200 ;
        RECT 110.200 61.100 110.600 67.900 ;
        RECT 112.600 67.900 113.500 68.200 ;
        RECT 115.000 67.900 115.900 68.200 ;
        RECT 116.600 67.900 117.000 69.900 ;
        RECT 117.400 68.000 117.800 69.900 ;
        RECT 119.000 68.000 119.400 69.900 ;
        RECT 117.400 67.900 119.400 68.000 ;
        RECT 119.800 68.000 120.200 69.900 ;
        RECT 121.400 68.000 121.800 69.900 ;
        RECT 119.800 67.900 121.800 68.000 ;
        RECT 122.200 67.900 122.600 69.900 ;
        RECT 124.600 67.900 125.000 69.900 ;
        RECT 125.300 68.200 125.700 68.600 ;
        RECT 111.000 66.800 111.400 67.600 ;
        RECT 111.800 66.800 112.200 67.600 ;
        RECT 112.600 61.100 113.000 67.900 ;
        RECT 114.200 66.800 114.600 67.600 ;
        RECT 115.000 66.100 115.400 67.900 ;
        RECT 116.700 67.200 117.000 67.900 ;
        RECT 117.500 67.700 119.300 67.900 ;
        RECT 119.900 67.700 121.700 67.900 ;
        RECT 118.600 67.200 119.000 67.400 ;
        RECT 120.200 67.200 120.600 67.400 ;
        RECT 122.200 67.200 122.500 67.900 ;
        RECT 116.600 66.800 117.900 67.200 ;
        RECT 118.600 66.900 119.400 67.200 ;
        RECT 119.000 66.800 119.400 66.900 ;
        RECT 119.800 66.900 120.600 67.200 ;
        RECT 119.800 66.800 120.200 66.900 ;
        RECT 121.300 66.800 122.600 67.200 ;
        RECT 115.000 65.800 116.900 66.100 ;
        RECT 113.400 65.100 113.800 65.200 ;
        RECT 114.200 65.100 114.600 65.200 ;
        RECT 113.400 64.800 114.600 65.100 ;
        RECT 113.400 64.400 113.800 64.800 ;
        RECT 115.000 61.100 115.400 65.800 ;
        RECT 116.600 65.200 116.900 65.800 ;
        RECT 115.800 64.400 116.200 65.200 ;
        RECT 116.600 65.100 117.000 65.200 ;
        RECT 117.600 65.100 117.900 66.800 ;
        RECT 118.200 65.800 118.600 66.600 ;
        RECT 120.600 65.800 121.000 66.600 ;
        RECT 121.300 66.100 121.600 66.800 ;
        RECT 123.800 66.400 124.200 67.200 ;
        RECT 123.000 66.100 123.400 66.200 ;
        RECT 124.600 66.100 124.900 67.900 ;
        RECT 125.400 67.800 125.800 68.200 ;
        RECT 126.200 68.000 126.600 69.900 ;
        RECT 127.800 68.000 128.200 69.900 ;
        RECT 126.200 67.900 128.200 68.000 ;
        RECT 128.600 67.900 129.000 69.900 ;
        RECT 126.300 67.700 128.100 67.900 ;
        RECT 126.600 67.200 127.000 67.400 ;
        RECT 128.600 67.200 128.900 67.900 ;
        RECT 129.400 67.700 129.800 69.900 ;
        RECT 131.500 69.200 132.100 69.900 ;
        RECT 131.500 68.900 132.200 69.200 ;
        RECT 133.800 68.900 134.200 69.900 ;
        RECT 136.000 69.200 136.400 69.900 ;
        RECT 136.000 68.900 137.000 69.200 ;
        RECT 131.800 68.500 132.200 68.900 ;
        RECT 133.900 68.600 134.200 68.900 ;
        RECT 133.900 68.300 135.300 68.600 ;
        RECT 134.900 68.200 135.300 68.300 ;
        RECT 135.800 68.200 136.200 68.600 ;
        RECT 136.600 68.500 137.000 68.900 ;
        RECT 130.900 67.700 131.300 67.800 ;
        RECT 129.400 67.400 131.300 67.700 ;
        RECT 126.200 66.900 127.000 67.200 ;
        RECT 126.200 66.800 126.600 66.900 ;
        RECT 127.700 66.800 129.000 67.200 ;
        RECT 125.400 66.100 125.800 66.200 ;
        RECT 127.000 66.100 127.400 66.600 ;
        RECT 121.300 65.800 123.800 66.100 ;
        RECT 124.600 65.800 127.400 66.100 ;
        RECT 121.300 65.100 121.600 65.800 ;
        RECT 123.400 65.600 123.800 65.800 ;
        RECT 122.200 65.100 122.600 65.200 ;
        RECT 125.400 65.100 125.700 65.800 ;
        RECT 127.700 65.100 128.000 66.800 ;
        RECT 128.600 66.200 128.900 66.800 ;
        RECT 128.600 65.800 129.000 66.200 ;
        RECT 129.400 65.700 129.800 67.400 ;
        RECT 132.900 67.100 133.300 67.200 ;
        RECT 135.800 67.100 136.100 68.200 ;
        RECT 138.200 67.500 138.600 69.900 ;
        RECT 142.200 67.900 142.600 69.900 ;
        RECT 142.900 68.200 143.300 68.600 ;
        RECT 137.400 67.100 138.200 67.200 ;
        RECT 132.700 66.800 138.200 67.100 ;
        RECT 139.000 67.100 139.400 67.200 ;
        RECT 141.400 67.100 141.800 67.200 ;
        RECT 139.000 66.800 141.800 67.100 ;
        RECT 131.800 66.400 132.200 66.500 ;
        RECT 130.300 66.100 132.200 66.400 ;
        RECT 132.700 66.200 133.000 66.800 ;
        RECT 136.300 66.700 136.700 66.800 ;
        RECT 141.400 66.400 141.800 66.800 ;
        RECT 137.100 66.200 137.500 66.300 ;
        RECT 130.300 66.000 130.700 66.100 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 135.000 66.100 137.500 66.200 ;
        RECT 134.200 65.900 137.500 66.100 ;
        RECT 140.600 66.100 141.000 66.200 ;
        RECT 142.200 66.100 142.500 67.900 ;
        RECT 143.000 67.800 143.400 68.200 ;
        RECT 145.600 67.100 146.000 69.900 ;
        RECT 147.000 68.000 147.400 69.900 ;
        RECT 148.600 68.000 149.000 69.900 ;
        RECT 147.000 67.900 149.000 68.000 ;
        RECT 149.400 67.900 149.800 69.900 ;
        RECT 150.200 68.500 150.600 69.500 ;
        RECT 147.100 67.700 148.900 67.900 ;
        RECT 147.400 67.200 147.800 67.400 ;
        RECT 149.400 67.200 149.700 67.900 ;
        RECT 150.200 67.400 150.500 68.500 ;
        RECT 152.300 68.000 152.700 69.500 ;
        RECT 152.300 67.700 153.100 68.000 ;
        RECT 152.700 67.500 153.100 67.700 ;
        RECT 145.600 66.900 146.500 67.100 ;
        RECT 145.700 66.800 146.500 66.900 ;
        RECT 147.000 66.900 147.800 67.200 ;
        RECT 147.000 66.800 147.400 66.900 ;
        RECT 148.500 66.800 149.800 67.200 ;
        RECT 150.200 67.100 152.300 67.400 ;
        RECT 151.800 66.900 152.300 67.100 ;
        RECT 152.800 67.200 153.100 67.500 ;
        RECT 156.600 67.900 157.000 69.900 ;
        RECT 159.800 67.900 160.200 69.900 ;
        RECT 160.500 68.200 160.900 68.600 ;
        RECT 143.000 66.100 143.400 66.200 ;
        RECT 134.200 65.800 135.400 65.900 ;
        RECT 140.600 65.800 141.400 66.100 ;
        RECT 142.200 65.800 143.400 66.100 ;
        RECT 144.600 65.800 145.400 66.200 ;
        RECT 131.100 65.700 131.500 65.800 ;
        RECT 129.400 65.400 131.500 65.700 ;
        RECT 128.600 65.100 129.000 65.200 ;
        RECT 116.600 64.800 117.300 65.100 ;
        RECT 117.600 64.800 118.100 65.100 ;
        RECT 117.000 64.200 117.300 64.800 ;
        RECT 117.000 63.800 117.400 64.200 ;
        RECT 117.700 61.100 118.100 64.800 ;
        RECT 121.100 64.800 121.600 65.100 ;
        RECT 121.900 64.800 122.600 65.100 ;
        RECT 123.000 64.800 125.000 65.100 ;
        RECT 121.100 61.100 121.500 64.800 ;
        RECT 121.900 64.200 122.200 64.800 ;
        RECT 121.800 63.800 122.200 64.200 ;
        RECT 123.000 61.100 123.400 64.800 ;
        RECT 124.600 61.100 125.000 64.800 ;
        RECT 125.400 61.100 125.800 65.100 ;
        RECT 127.500 64.800 128.000 65.100 ;
        RECT 128.300 64.800 129.000 65.100 ;
        RECT 127.500 61.100 127.900 64.800 ;
        RECT 128.300 64.200 128.600 64.800 ;
        RECT 128.200 63.800 128.600 64.200 ;
        RECT 129.400 61.100 129.800 65.400 ;
        RECT 132.700 65.200 133.000 65.800 ;
        RECT 141.000 65.600 141.400 65.800 ;
        RECT 135.800 65.500 138.600 65.600 ;
        RECT 135.700 65.400 138.600 65.500 ;
        RECT 131.800 64.900 133.000 65.200 ;
        RECT 133.700 65.300 138.600 65.400 ;
        RECT 133.700 65.100 136.100 65.300 ;
        RECT 131.800 64.400 132.100 64.900 ;
        RECT 131.400 64.200 132.100 64.400 ;
        RECT 132.900 64.500 133.300 64.600 ;
        RECT 133.700 64.500 134.000 65.100 ;
        RECT 132.900 64.200 134.000 64.500 ;
        RECT 134.300 64.500 137.000 64.800 ;
        RECT 134.300 64.400 134.700 64.500 ;
        RECT 136.600 64.400 137.000 64.500 ;
        RECT 131.000 64.000 132.100 64.200 ;
        RECT 131.000 63.800 131.700 64.000 ;
        RECT 133.500 63.700 133.900 63.800 ;
        RECT 134.900 63.700 135.300 63.800 ;
        RECT 131.800 63.100 132.200 63.500 ;
        RECT 133.500 63.400 135.300 63.700 ;
        RECT 133.900 63.100 134.200 63.400 ;
        RECT 136.600 63.100 137.000 63.500 ;
        RECT 131.500 61.100 132.100 63.100 ;
        RECT 133.800 61.100 134.200 63.100 ;
        RECT 136.000 62.800 137.000 63.100 ;
        RECT 136.000 61.100 136.400 62.800 ;
        RECT 138.200 61.100 138.600 65.300 ;
        RECT 143.000 65.100 143.300 65.800 ;
        RECT 140.600 64.800 142.600 65.100 ;
        RECT 140.600 61.100 141.000 64.800 ;
        RECT 142.200 61.100 142.600 64.800 ;
        RECT 143.000 64.100 143.400 65.100 ;
        RECT 143.800 64.800 144.200 65.600 ;
        RECT 146.200 65.200 146.500 66.800 ;
        RECT 147.800 65.800 148.200 66.600 ;
        RECT 146.200 64.800 146.600 65.200 ;
        RECT 148.500 65.100 148.800 66.800 ;
        RECT 150.200 65.800 150.600 66.600 ;
        RECT 151.000 65.800 151.400 66.600 ;
        RECT 151.800 66.500 152.500 66.900 ;
        RECT 152.800 66.800 153.800 67.200 ;
        RECT 151.800 65.500 152.100 66.500 ;
        RECT 150.200 65.200 152.100 65.500 ;
        RECT 149.400 65.100 149.800 65.200 ;
        RECT 148.300 64.800 148.800 65.100 ;
        RECT 149.100 64.800 149.800 65.100 ;
        RECT 145.400 64.100 145.800 64.600 ;
        RECT 143.000 63.800 145.800 64.100 ;
        RECT 143.000 61.100 143.400 63.800 ;
        RECT 146.200 63.500 146.500 64.800 ;
        RECT 144.700 63.200 146.500 63.500 ;
        RECT 144.700 63.100 145.000 63.200 ;
        RECT 144.600 61.100 145.000 63.100 ;
        RECT 146.200 63.100 146.500 63.200 ;
        RECT 146.200 61.100 146.600 63.100 ;
        RECT 148.300 61.100 148.700 64.800 ;
        RECT 149.100 64.200 149.400 64.800 ;
        RECT 149.000 63.800 149.400 64.200 ;
        RECT 150.200 63.500 150.500 65.200 ;
        RECT 152.800 64.900 153.100 66.800 ;
        RECT 155.800 66.400 156.200 67.200 ;
        RECT 153.400 65.400 153.800 66.200 ;
        RECT 155.000 66.100 155.400 66.200 ;
        RECT 156.600 66.100 156.900 67.900 ;
        RECT 159.000 66.400 159.400 67.200 ;
        RECT 157.400 66.100 157.800 66.200 ;
        RECT 158.200 66.100 158.600 66.200 ;
        RECT 159.800 66.100 160.100 67.900 ;
        RECT 160.600 67.800 161.000 68.200 ;
        RECT 163.000 67.900 163.400 69.900 ;
        RECT 164.600 67.900 165.000 69.900 ;
        RECT 165.400 68.000 165.800 69.900 ;
        RECT 167.000 68.000 167.400 69.900 ;
        RECT 165.400 67.900 167.400 68.000 ;
        RECT 169.400 67.900 169.800 69.900 ;
        RECT 170.100 68.200 170.500 68.600 ;
        RECT 170.200 68.100 170.600 68.200 ;
        RECT 171.000 68.100 171.400 69.900 ;
        RECT 162.200 66.400 162.600 67.200 ;
        RECT 160.600 66.100 161.000 66.200 ;
        RECT 155.000 65.800 155.800 66.100 ;
        RECT 156.600 65.800 159.000 66.100 ;
        RECT 159.800 65.800 161.000 66.100 ;
        RECT 161.400 66.100 161.800 66.200 ;
        RECT 163.000 66.100 163.300 67.900 ;
        RECT 164.700 67.200 165.000 67.900 ;
        RECT 165.500 67.700 167.300 67.900 ;
        RECT 166.600 67.200 167.000 67.400 ;
        RECT 164.600 66.800 165.900 67.200 ;
        RECT 166.600 66.900 167.400 67.200 ;
        RECT 167.000 66.800 167.400 66.900 ;
        RECT 163.800 66.100 164.200 66.200 ;
        RECT 161.400 65.800 162.200 66.100 ;
        RECT 163.000 65.800 164.200 66.100 ;
        RECT 155.400 65.600 155.800 65.800 ;
        RECT 157.400 65.100 157.700 65.800 ;
        RECT 158.600 65.600 159.000 65.800 ;
        RECT 160.600 65.100 160.900 65.800 ;
        RECT 161.800 65.600 162.200 65.800 ;
        RECT 163.800 65.100 164.100 65.800 ;
        RECT 164.600 65.100 165.000 65.200 ;
        RECT 165.600 65.100 165.900 66.800 ;
        RECT 166.200 65.800 166.600 66.600 ;
        RECT 168.600 66.400 169.000 67.200 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 169.400 66.100 169.700 67.900 ;
        RECT 170.200 67.800 171.400 68.100 ;
        RECT 171.800 68.000 172.200 69.900 ;
        RECT 173.400 68.000 173.800 69.900 ;
        RECT 171.800 67.900 173.800 68.000 ;
        RECT 171.100 67.200 171.400 67.800 ;
        RECT 171.900 67.700 173.700 67.900 ;
        RECT 174.200 67.500 174.600 69.900 ;
        RECT 176.400 69.200 176.800 69.900 ;
        RECT 175.800 68.900 176.800 69.200 ;
        RECT 178.600 68.900 179.000 69.900 ;
        RECT 180.700 69.200 181.300 69.900 ;
        RECT 180.600 68.900 181.300 69.200 ;
        RECT 175.800 68.500 176.200 68.900 ;
        RECT 178.600 68.600 178.900 68.900 ;
        RECT 176.600 68.200 177.000 68.600 ;
        RECT 177.500 68.300 178.900 68.600 ;
        RECT 180.600 68.500 181.000 68.900 ;
        RECT 177.500 68.200 177.900 68.300 ;
        RECT 173.000 67.200 173.400 67.400 ;
        RECT 171.000 66.800 172.300 67.200 ;
        RECT 173.000 66.900 173.800 67.200 ;
        RECT 173.400 66.800 173.800 66.900 ;
        RECT 174.600 67.100 175.400 67.200 ;
        RECT 176.700 67.100 177.000 68.200 ;
        RECT 181.500 67.700 181.900 67.800 ;
        RECT 183.000 67.700 183.400 69.900 ;
        RECT 184.100 69.200 184.500 69.900 ;
        RECT 187.500 69.200 187.900 69.900 ;
        RECT 183.800 68.800 184.500 69.200 ;
        RECT 187.000 68.800 187.900 69.200 ;
        RECT 184.100 68.200 184.500 68.800 ;
        RECT 187.500 68.200 187.900 68.800 ;
        RECT 184.100 67.900 185.000 68.200 ;
        RECT 181.500 67.400 183.400 67.700 ;
        RECT 177.400 67.100 177.800 67.200 ;
        RECT 179.500 67.100 179.900 67.200 ;
        RECT 174.600 66.800 180.100 67.100 ;
        RECT 170.200 66.100 170.600 66.200 ;
        RECT 167.800 65.800 168.600 66.100 ;
        RECT 169.400 65.800 170.600 66.100 ;
        RECT 168.200 65.600 168.600 65.800 ;
        RECT 170.200 65.100 170.500 65.800 ;
        RECT 171.000 65.100 171.400 65.200 ;
        RECT 172.000 65.100 172.300 66.800 ;
        RECT 176.100 66.700 176.500 66.800 ;
        RECT 172.600 65.800 173.000 66.600 ;
        RECT 175.300 66.200 175.700 66.300 ;
        RECT 176.600 66.200 177.000 66.300 ;
        RECT 175.300 65.900 177.800 66.200 ;
        RECT 177.400 65.800 177.800 65.900 ;
        RECT 174.200 65.500 177.000 65.600 ;
        RECT 174.200 65.400 177.100 65.500 ;
        RECT 174.200 65.300 179.100 65.400 ;
        RECT 152.300 64.600 153.100 64.900 ;
        RECT 155.000 64.800 157.000 65.100 ;
        RECT 150.200 61.500 150.600 63.500 ;
        RECT 152.300 62.200 152.700 64.600 ;
        RECT 151.800 61.800 152.700 62.200 ;
        RECT 152.300 61.100 152.700 61.800 ;
        RECT 155.000 61.100 155.400 64.800 ;
        RECT 156.600 61.100 157.000 64.800 ;
        RECT 157.400 61.100 157.800 65.100 ;
        RECT 158.200 64.800 160.200 65.100 ;
        RECT 158.200 61.100 158.600 64.800 ;
        RECT 159.800 61.100 160.200 64.800 ;
        RECT 160.600 61.100 161.000 65.100 ;
        RECT 161.400 64.800 163.400 65.100 ;
        RECT 161.400 61.100 161.800 64.800 ;
        RECT 163.000 61.100 163.400 64.800 ;
        RECT 163.800 61.100 164.200 65.100 ;
        RECT 164.600 64.800 165.300 65.100 ;
        RECT 165.600 64.800 166.100 65.100 ;
        RECT 165.000 64.200 165.300 64.800 ;
        RECT 165.000 63.800 165.400 64.200 ;
        RECT 165.700 61.100 166.100 64.800 ;
        RECT 167.800 64.800 169.800 65.100 ;
        RECT 167.800 61.100 168.200 64.800 ;
        RECT 169.400 61.100 169.800 64.800 ;
        RECT 170.200 61.100 170.600 65.100 ;
        RECT 171.000 64.800 171.700 65.100 ;
        RECT 172.000 64.800 172.500 65.100 ;
        RECT 171.400 64.200 171.700 64.800 ;
        RECT 171.400 63.800 171.800 64.200 ;
        RECT 172.100 61.100 172.500 64.800 ;
        RECT 174.200 61.100 174.600 65.300 ;
        RECT 176.700 65.100 179.100 65.300 ;
        RECT 175.800 64.500 178.500 64.800 ;
        RECT 175.800 64.400 176.200 64.500 ;
        RECT 178.100 64.400 178.500 64.500 ;
        RECT 178.800 64.500 179.100 65.100 ;
        RECT 179.800 65.200 180.100 66.800 ;
        RECT 180.600 66.400 181.000 66.500 ;
        RECT 180.600 66.100 182.500 66.400 ;
        RECT 182.100 66.000 182.500 66.100 ;
        RECT 181.300 65.700 181.700 65.800 ;
        RECT 183.000 65.700 183.400 67.400 ;
        RECT 181.300 65.400 183.400 65.700 ;
        RECT 179.800 64.900 181.000 65.200 ;
        RECT 179.500 64.500 179.900 64.600 ;
        RECT 178.800 64.200 179.900 64.500 ;
        RECT 180.700 64.400 181.000 64.900 ;
        RECT 180.700 64.000 181.400 64.400 ;
        RECT 177.500 63.700 177.900 63.800 ;
        RECT 178.900 63.700 179.300 63.800 ;
        RECT 175.800 63.100 176.200 63.500 ;
        RECT 177.500 63.400 179.300 63.700 ;
        RECT 178.600 63.100 178.900 63.400 ;
        RECT 180.600 63.100 181.000 63.500 ;
        RECT 175.800 62.800 176.800 63.100 ;
        RECT 176.400 61.100 176.800 62.800 ;
        RECT 178.600 61.100 179.000 63.100 ;
        RECT 180.700 61.100 181.300 63.100 ;
        RECT 183.000 61.100 183.400 65.400 ;
        RECT 183.800 64.400 184.200 65.200 ;
        RECT 184.600 61.100 185.000 67.900 ;
        RECT 187.000 67.900 187.900 68.200 ;
        RECT 185.400 66.800 185.800 67.600 ;
        RECT 186.200 66.800 186.600 67.600 ;
        RECT 187.000 61.100 187.400 67.900 ;
        RECT 188.600 67.600 189.000 69.900 ;
        RECT 190.200 68.200 190.600 69.900 ;
        RECT 190.200 67.900 190.700 68.200 ;
        RECT 188.600 67.300 189.900 67.600 ;
        RECT 188.700 66.200 189.100 66.600 ;
        RECT 188.600 65.800 189.100 66.200 ;
        RECT 189.600 66.500 189.900 67.300 ;
        RECT 190.400 67.200 190.700 67.900 ;
        RECT 190.200 66.800 190.700 67.200 ;
        RECT 189.600 66.100 190.100 66.500 ;
        RECT 187.800 64.400 188.200 65.200 ;
        RECT 189.600 65.100 189.900 66.100 ;
        RECT 190.400 65.100 190.700 66.800 ;
        RECT 188.600 64.800 189.900 65.100 ;
        RECT 188.600 61.100 189.000 64.800 ;
        RECT 190.200 64.600 190.700 65.100 ;
        RECT 193.400 67.700 193.800 69.900 ;
        RECT 195.500 69.200 196.100 69.900 ;
        RECT 195.500 68.900 196.200 69.200 ;
        RECT 197.800 68.900 198.200 69.900 ;
        RECT 200.000 69.200 200.400 69.900 ;
        RECT 200.000 68.900 201.000 69.200 ;
        RECT 195.800 68.500 196.200 68.900 ;
        RECT 197.900 68.600 198.200 68.900 ;
        RECT 197.900 68.300 199.300 68.600 ;
        RECT 198.900 68.200 199.300 68.300 ;
        RECT 199.800 68.200 200.200 68.600 ;
        RECT 200.600 68.500 201.000 68.900 ;
        RECT 194.900 67.700 195.300 67.800 ;
        RECT 193.400 67.400 195.300 67.700 ;
        RECT 193.400 65.700 193.800 67.400 ;
        RECT 196.900 67.100 197.300 67.200 ;
        RECT 199.800 67.100 200.100 68.200 ;
        RECT 202.200 67.500 202.600 69.900 ;
        RECT 203.000 68.000 203.400 69.900 ;
        RECT 204.600 68.000 205.000 69.900 ;
        RECT 203.000 67.900 205.000 68.000 ;
        RECT 205.400 67.900 205.800 69.900 ;
        RECT 207.500 68.200 207.900 69.900 ;
        RECT 207.000 67.900 207.900 68.200 ;
        RECT 208.600 67.900 209.000 69.900 ;
        RECT 209.400 68.000 209.800 69.900 ;
        RECT 211.000 68.000 211.400 69.900 ;
        RECT 209.400 67.900 211.400 68.000 ;
        RECT 203.100 67.700 204.900 67.900 ;
        RECT 203.400 67.200 203.800 67.400 ;
        RECT 205.400 67.200 205.700 67.900 ;
        RECT 201.400 67.100 202.200 67.200 ;
        RECT 196.700 66.800 202.200 67.100 ;
        RECT 203.000 66.900 203.800 67.200 ;
        RECT 203.000 66.800 203.400 66.900 ;
        RECT 204.500 66.800 205.800 67.200 ;
        RECT 206.200 66.800 206.600 67.600 ;
        RECT 195.800 66.400 196.200 66.500 ;
        RECT 194.300 66.100 196.200 66.400 ;
        RECT 194.300 66.000 194.700 66.100 ;
        RECT 195.100 65.700 195.500 65.800 ;
        RECT 193.400 65.400 195.500 65.700 ;
        RECT 190.200 61.100 190.600 64.600 ;
        RECT 193.400 61.100 193.800 65.400 ;
        RECT 196.700 65.200 197.000 66.800 ;
        RECT 200.300 66.700 200.700 66.800 ;
        RECT 199.800 66.200 200.200 66.300 ;
        RECT 201.100 66.200 201.500 66.300 ;
        RECT 199.000 65.900 201.500 66.200 ;
        RECT 199.000 65.800 199.400 65.900 ;
        RECT 203.800 65.800 204.200 66.600 ;
        RECT 204.500 66.200 204.800 66.800 ;
        RECT 204.500 65.800 205.000 66.200 ;
        RECT 199.800 65.500 202.600 65.600 ;
        RECT 199.700 65.400 202.600 65.500 ;
        RECT 195.800 64.900 197.000 65.200 ;
        RECT 197.700 65.300 202.600 65.400 ;
        RECT 197.700 65.100 200.100 65.300 ;
        RECT 195.800 64.400 196.100 64.900 ;
        RECT 195.400 64.000 196.100 64.400 ;
        RECT 196.900 64.500 197.300 64.600 ;
        RECT 197.700 64.500 198.000 65.100 ;
        RECT 196.900 64.200 198.000 64.500 ;
        RECT 198.300 64.500 201.000 64.800 ;
        RECT 198.300 64.400 198.700 64.500 ;
        RECT 200.600 64.400 201.000 64.500 ;
        RECT 197.500 63.700 197.900 63.800 ;
        RECT 198.900 63.700 199.300 63.800 ;
        RECT 195.800 63.100 196.200 63.500 ;
        RECT 197.500 63.400 199.300 63.700 ;
        RECT 197.900 63.100 198.200 63.400 ;
        RECT 200.600 63.100 201.000 63.500 ;
        RECT 195.500 61.100 196.100 63.100 ;
        RECT 197.800 61.100 198.200 63.100 ;
        RECT 200.000 62.800 201.000 63.100 ;
        RECT 200.000 61.100 200.400 62.800 ;
        RECT 202.200 61.100 202.600 65.300 ;
        RECT 204.500 65.100 204.800 65.800 ;
        RECT 205.400 65.100 205.800 65.200 ;
        RECT 207.000 65.100 207.400 67.900 ;
        RECT 208.700 67.200 209.000 67.900 ;
        RECT 209.500 67.700 211.300 67.900 ;
        RECT 211.800 67.700 212.200 69.900 ;
        RECT 213.900 69.200 214.500 69.900 ;
        RECT 213.900 68.900 214.600 69.200 ;
        RECT 216.200 68.900 216.600 69.900 ;
        RECT 218.400 69.200 218.800 69.900 ;
        RECT 218.400 68.900 219.400 69.200 ;
        RECT 214.200 68.500 214.600 68.900 ;
        RECT 216.300 68.600 216.600 68.900 ;
        RECT 216.300 68.300 217.700 68.600 ;
        RECT 217.300 68.200 217.700 68.300 ;
        RECT 218.200 68.200 218.600 68.600 ;
        RECT 219.000 68.500 219.400 68.900 ;
        RECT 213.300 67.700 213.700 67.800 ;
        RECT 211.800 67.400 213.700 67.700 ;
        RECT 210.600 67.200 211.000 67.400 ;
        RECT 208.600 66.800 209.900 67.200 ;
        RECT 210.600 66.900 211.400 67.200 ;
        RECT 211.000 66.800 211.400 66.900 ;
        RECT 208.600 66.100 209.000 66.200 ;
        RECT 209.600 66.100 209.900 66.800 ;
        RECT 208.600 65.800 209.900 66.100 ;
        RECT 210.200 65.800 210.600 66.600 ;
        RECT 204.300 64.800 204.800 65.100 ;
        RECT 205.100 64.800 207.400 65.100 ;
        RECT 204.300 61.100 204.700 64.800 ;
        RECT 205.100 64.200 205.400 64.800 ;
        RECT 205.000 63.800 205.400 64.200 ;
        RECT 207.000 61.100 207.400 64.800 ;
        RECT 207.800 64.400 208.200 65.200 ;
        RECT 208.600 65.100 209.000 65.200 ;
        RECT 209.600 65.100 209.900 65.800 ;
        RECT 211.800 65.700 212.200 67.400 ;
        RECT 215.300 67.100 215.700 67.200 ;
        RECT 218.200 67.100 218.500 68.200 ;
        RECT 220.600 67.500 221.000 69.900 ;
        RECT 221.400 67.500 221.800 69.900 ;
        RECT 223.600 69.200 224.000 69.900 ;
        RECT 223.000 68.900 224.000 69.200 ;
        RECT 225.800 68.900 226.200 69.900 ;
        RECT 227.900 69.200 228.500 69.900 ;
        RECT 227.800 68.900 228.500 69.200 ;
        RECT 223.000 68.500 223.400 68.900 ;
        RECT 225.800 68.600 226.100 68.900 ;
        RECT 223.800 68.200 224.200 68.600 ;
        RECT 224.700 68.300 226.100 68.600 ;
        RECT 227.800 68.500 228.200 68.900 ;
        RECT 224.700 68.200 225.100 68.300 ;
        RECT 219.800 67.100 220.600 67.200 ;
        RECT 221.800 67.100 222.600 67.200 ;
        RECT 223.900 67.100 224.200 68.200 ;
        RECT 227.000 68.100 227.400 68.200 ;
        RECT 227.000 67.800 229.000 68.100 ;
        RECT 228.600 67.700 229.100 67.800 ;
        RECT 230.200 67.700 230.600 69.900 ;
        RECT 228.600 67.400 230.600 67.700 ;
        RECT 225.400 67.100 225.800 67.200 ;
        RECT 226.700 67.100 227.100 67.200 ;
        RECT 215.100 66.800 227.300 67.100 ;
        RECT 214.200 66.400 214.600 66.500 ;
        RECT 212.700 66.100 214.600 66.400 ;
        RECT 212.700 66.000 213.100 66.100 ;
        RECT 213.500 65.700 213.900 65.800 ;
        RECT 211.800 65.400 213.900 65.700 ;
        RECT 208.600 64.800 209.300 65.100 ;
        RECT 209.600 64.800 210.100 65.100 ;
        RECT 209.000 64.200 209.300 64.800 ;
        RECT 209.000 63.800 209.400 64.200 ;
        RECT 209.700 61.100 210.100 64.800 ;
        RECT 211.800 61.100 212.200 65.400 ;
        RECT 215.100 65.200 215.400 66.800 ;
        RECT 218.700 66.700 219.100 66.800 ;
        RECT 223.300 66.700 223.700 66.800 ;
        RECT 219.500 66.200 219.900 66.300 ;
        RECT 217.400 65.900 219.900 66.200 ;
        RECT 222.500 66.200 222.900 66.300 ;
        RECT 222.500 65.900 225.000 66.200 ;
        RECT 217.400 65.800 217.800 65.900 ;
        RECT 224.600 65.800 225.000 65.900 ;
        RECT 218.200 65.500 221.000 65.600 ;
        RECT 218.100 65.400 221.000 65.500 ;
        RECT 214.200 64.900 215.400 65.200 ;
        RECT 216.100 65.300 221.000 65.400 ;
        RECT 216.100 65.100 218.500 65.300 ;
        RECT 214.200 64.400 214.500 64.900 ;
        RECT 213.800 64.200 214.500 64.400 ;
        RECT 215.300 64.500 215.700 64.600 ;
        RECT 216.100 64.500 216.400 65.100 ;
        RECT 215.300 64.200 216.400 64.500 ;
        RECT 216.700 64.500 219.400 64.800 ;
        RECT 216.700 64.400 217.100 64.500 ;
        RECT 219.000 64.400 219.400 64.500 ;
        RECT 213.400 64.000 214.500 64.200 ;
        RECT 213.400 63.800 214.100 64.000 ;
        RECT 215.900 63.700 216.300 63.800 ;
        RECT 217.300 63.700 217.700 63.800 ;
        RECT 214.200 63.100 214.600 63.500 ;
        RECT 215.900 63.400 217.700 63.700 ;
        RECT 216.300 63.100 216.600 63.400 ;
        RECT 219.000 63.100 219.400 63.500 ;
        RECT 213.900 61.100 214.500 63.100 ;
        RECT 216.200 61.100 216.600 63.100 ;
        RECT 218.400 62.800 219.400 63.100 ;
        RECT 218.400 61.100 218.800 62.800 ;
        RECT 220.600 61.100 221.000 65.300 ;
        RECT 221.400 65.500 224.200 65.600 ;
        RECT 221.400 65.400 224.300 65.500 ;
        RECT 221.400 65.300 226.300 65.400 ;
        RECT 221.400 61.100 221.800 65.300 ;
        RECT 223.900 65.100 226.300 65.300 ;
        RECT 223.000 64.500 225.700 64.800 ;
        RECT 223.000 64.400 223.400 64.500 ;
        RECT 225.300 64.400 225.700 64.500 ;
        RECT 226.000 64.500 226.300 65.100 ;
        RECT 227.000 65.200 227.300 66.800 ;
        RECT 227.800 66.400 228.200 66.500 ;
        RECT 227.800 66.100 229.700 66.400 ;
        RECT 229.300 66.000 229.700 66.100 ;
        RECT 228.500 65.700 228.900 65.800 ;
        RECT 230.200 65.700 230.600 67.400 ;
        RECT 228.500 65.400 230.600 65.700 ;
        RECT 227.000 64.900 228.200 65.200 ;
        RECT 226.700 64.500 227.100 64.600 ;
        RECT 226.000 64.200 227.100 64.500 ;
        RECT 227.900 64.400 228.200 64.900 ;
        RECT 227.900 64.000 228.600 64.400 ;
        RECT 224.700 63.700 225.100 63.800 ;
        RECT 226.100 63.700 226.500 63.800 ;
        RECT 223.000 63.100 223.400 63.500 ;
        RECT 224.700 63.400 226.500 63.700 ;
        RECT 225.800 63.100 226.100 63.400 ;
        RECT 227.800 63.100 228.200 63.500 ;
        RECT 223.000 62.800 224.000 63.100 ;
        RECT 223.600 61.100 224.000 62.800 ;
        RECT 225.800 61.100 226.200 63.100 ;
        RECT 227.900 61.100 228.500 63.100 ;
        RECT 230.200 61.100 230.600 65.400 ;
        RECT 0.600 56.200 1.000 59.900 ;
        RECT 2.200 56.400 2.600 59.900 ;
        RECT 0.600 55.900 1.900 56.200 ;
        RECT 2.200 55.900 2.700 56.400 ;
        RECT 0.600 54.800 1.100 55.200 ;
        RECT 0.700 54.400 1.100 54.800 ;
        RECT 1.600 54.900 1.900 55.900 ;
        RECT 1.600 54.500 2.100 54.900 ;
        RECT 1.600 53.700 1.900 54.500 ;
        RECT 2.400 54.200 2.700 55.900 ;
        RECT 3.800 55.700 4.200 59.900 ;
        RECT 6.000 58.200 6.400 59.900 ;
        RECT 5.400 57.900 6.400 58.200 ;
        RECT 8.200 57.900 8.600 59.900 ;
        RECT 10.300 57.900 10.900 59.900 ;
        RECT 5.400 57.500 5.800 57.900 ;
        RECT 8.200 57.600 8.500 57.900 ;
        RECT 7.100 57.300 8.900 57.600 ;
        RECT 10.200 57.500 10.600 57.900 ;
        RECT 7.100 57.200 7.500 57.300 ;
        RECT 8.500 57.200 8.900 57.300 ;
        RECT 5.400 56.500 5.800 56.600 ;
        RECT 7.700 56.500 8.100 56.600 ;
        RECT 5.400 56.200 8.100 56.500 ;
        RECT 8.400 56.500 9.500 56.800 ;
        RECT 8.400 55.900 8.700 56.500 ;
        RECT 9.100 56.400 9.500 56.500 ;
        RECT 10.300 56.600 11.000 57.000 ;
        RECT 10.300 56.100 10.600 56.600 ;
        RECT 6.300 55.700 8.700 55.900 ;
        RECT 3.800 55.600 8.700 55.700 ;
        RECT 9.400 55.800 10.600 56.100 ;
        RECT 3.800 55.500 6.700 55.600 ;
        RECT 3.800 55.400 6.600 55.500 ;
        RECT 2.200 54.100 2.700 54.200 ;
        RECT 3.000 54.800 3.400 55.200 ;
        RECT 7.000 55.100 7.400 55.200 ;
        RECT 4.900 54.800 7.400 55.100 ;
        RECT 3.000 54.100 3.300 54.800 ;
        RECT 4.900 54.700 5.300 54.800 ;
        RECT 5.700 54.200 6.100 54.300 ;
        RECT 9.400 54.200 9.700 55.800 ;
        RECT 12.600 55.600 13.000 59.900 ;
        RECT 10.900 55.300 13.000 55.600 ;
        RECT 10.900 55.200 11.300 55.300 ;
        RECT 11.700 54.900 12.100 55.000 ;
        RECT 10.200 54.600 12.100 54.900 ;
        RECT 10.200 54.500 10.600 54.600 ;
        RECT 2.200 53.800 3.300 54.100 ;
        RECT 4.200 53.900 9.700 54.200 ;
        RECT 4.200 53.800 5.000 53.900 ;
        RECT 0.600 53.400 1.900 53.700 ;
        RECT 0.600 51.100 1.000 53.400 ;
        RECT 2.400 53.100 2.700 53.800 ;
        RECT 2.200 52.800 2.700 53.100 ;
        RECT 2.200 51.100 2.600 52.800 ;
        RECT 3.800 51.100 4.200 53.500 ;
        RECT 6.300 52.800 6.600 53.900 ;
        RECT 7.800 53.800 8.200 53.900 ;
        RECT 9.100 53.800 9.500 53.900 ;
        RECT 12.600 53.600 13.000 55.300 ;
        RECT 11.100 53.300 13.000 53.600 ;
        RECT 13.400 53.400 13.800 54.200 ;
        RECT 11.100 53.200 11.500 53.300 ;
        RECT 5.400 52.100 5.800 52.500 ;
        RECT 6.200 52.400 6.600 52.800 ;
        RECT 7.100 52.700 7.500 52.800 ;
        RECT 7.100 52.400 8.500 52.700 ;
        RECT 8.200 52.100 8.500 52.400 ;
        RECT 10.200 52.100 10.600 52.500 ;
        RECT 5.400 51.800 6.400 52.100 ;
        RECT 6.000 51.100 6.400 51.800 ;
        RECT 8.200 51.100 8.600 52.100 ;
        RECT 10.200 51.800 10.900 52.100 ;
        RECT 10.300 51.100 10.900 51.800 ;
        RECT 12.600 51.100 13.000 53.300 ;
        RECT 14.200 53.100 14.600 59.900 ;
        RECT 17.100 57.200 17.500 59.900 ;
        RECT 16.600 56.800 17.500 57.200 ;
        RECT 17.800 56.800 18.200 57.200 ;
        RECT 15.000 55.800 15.400 56.600 ;
        RECT 17.100 56.200 17.500 56.800 ;
        RECT 17.900 56.200 18.200 56.800 ;
        RECT 17.100 55.900 17.600 56.200 ;
        RECT 17.900 55.900 18.600 56.200 ;
        RECT 16.600 54.400 17.000 55.200 ;
        RECT 17.300 54.200 17.600 55.900 ;
        RECT 18.200 55.800 18.600 55.900 ;
        RECT 19.000 55.800 19.400 56.600 ;
        RECT 18.200 55.100 18.500 55.800 ;
        RECT 19.800 55.100 20.200 59.900 ;
        RECT 22.200 55.600 22.600 59.900 ;
        RECT 23.800 55.600 24.200 59.900 ;
        RECT 25.400 55.600 25.800 59.900 ;
        RECT 27.000 55.600 27.400 59.900 ;
        RECT 22.200 55.200 23.100 55.600 ;
        RECT 23.800 55.200 24.900 55.600 ;
        RECT 25.400 55.200 26.500 55.600 ;
        RECT 27.000 55.200 28.200 55.600 ;
        RECT 18.200 54.800 20.200 55.100 ;
        RECT 15.800 54.100 16.200 54.200 ;
        RECT 15.800 53.800 16.600 54.100 ;
        RECT 17.300 53.800 18.600 54.200 ;
        RECT 16.200 53.600 16.600 53.800 ;
        RECT 15.900 53.100 17.700 53.300 ;
        RECT 18.200 53.100 18.500 53.800 ;
        RECT 19.800 53.100 20.200 54.800 ;
        RECT 20.600 54.800 21.000 55.200 ;
        RECT 20.600 54.200 20.900 54.800 ;
        RECT 22.700 54.500 23.100 55.200 ;
        RECT 24.500 54.500 24.900 55.200 ;
        RECT 26.100 54.500 26.500 55.200 ;
        RECT 20.600 53.400 21.000 54.200 ;
        RECT 22.700 54.100 24.000 54.500 ;
        RECT 24.500 54.100 25.700 54.500 ;
        RECT 26.100 54.100 27.400 54.500 ;
        RECT 22.700 53.800 23.100 54.100 ;
        RECT 24.500 53.800 24.900 54.100 ;
        RECT 26.100 53.800 26.500 54.100 ;
        RECT 27.800 53.800 28.200 55.200 ;
        RECT 22.200 53.400 23.100 53.800 ;
        RECT 23.800 53.400 24.900 53.800 ;
        RECT 25.400 53.400 26.500 53.800 ;
        RECT 27.000 53.400 28.200 53.800 ;
        RECT 28.600 53.400 29.000 54.200 ;
        RECT 14.200 52.800 15.100 53.100 ;
        RECT 14.700 51.100 15.100 52.800 ;
        RECT 15.800 53.000 17.800 53.100 ;
        RECT 15.800 51.100 16.200 53.000 ;
        RECT 17.400 51.100 17.800 53.000 ;
        RECT 18.200 51.100 18.600 53.100 ;
        RECT 19.300 52.800 20.200 53.100 ;
        RECT 19.300 51.100 19.700 52.800 ;
        RECT 22.200 51.100 22.600 53.400 ;
        RECT 23.800 51.100 24.200 53.400 ;
        RECT 25.400 51.100 25.800 53.400 ;
        RECT 27.000 51.100 27.400 53.400 ;
        RECT 29.400 53.100 29.800 59.900 ;
        RECT 32.300 59.200 32.700 59.900 ;
        RECT 31.800 58.800 32.700 59.200 ;
        RECT 30.200 55.800 30.600 56.600 ;
        RECT 32.300 56.200 32.700 58.800 ;
        RECT 33.000 56.800 33.400 57.200 ;
        RECT 33.100 56.200 33.400 56.800 ;
        RECT 32.300 55.900 32.800 56.200 ;
        RECT 33.100 56.100 33.800 56.200 ;
        RECT 34.200 56.100 34.600 56.200 ;
        RECT 33.100 55.900 34.600 56.100 ;
        RECT 31.800 54.400 32.200 55.200 ;
        RECT 32.500 54.200 32.800 55.900 ;
        RECT 33.400 55.800 34.600 55.900 ;
        RECT 35.800 55.700 36.200 59.900 ;
        RECT 38.000 58.200 38.400 59.900 ;
        RECT 37.400 57.900 38.400 58.200 ;
        RECT 40.200 57.900 40.600 59.900 ;
        RECT 42.300 57.900 42.900 59.900 ;
        RECT 37.400 57.500 37.800 57.900 ;
        RECT 40.200 57.600 40.500 57.900 ;
        RECT 39.100 57.300 40.900 57.600 ;
        RECT 42.200 57.500 42.600 57.900 ;
        RECT 39.100 57.200 39.500 57.300 ;
        RECT 40.500 57.200 40.900 57.300 ;
        RECT 37.400 56.500 37.800 56.600 ;
        RECT 39.700 56.500 40.100 56.600 ;
        RECT 37.400 56.200 40.100 56.500 ;
        RECT 40.400 56.500 41.500 56.800 ;
        RECT 40.400 55.900 40.700 56.500 ;
        RECT 41.100 56.400 41.500 56.500 ;
        RECT 42.300 56.600 43.000 57.000 ;
        RECT 42.300 56.100 42.600 56.600 ;
        RECT 38.300 55.700 40.700 55.900 ;
        RECT 35.800 55.600 40.700 55.700 ;
        RECT 41.400 55.800 42.600 56.100 ;
        RECT 35.800 55.500 38.700 55.600 ;
        RECT 35.800 55.400 38.600 55.500 ;
        RECT 39.000 55.100 39.400 55.200 ;
        RECT 39.800 55.100 40.200 55.200 ;
        RECT 36.900 54.800 40.200 55.100 ;
        RECT 36.900 54.700 37.300 54.800 ;
        RECT 37.700 54.200 38.100 54.300 ;
        RECT 41.400 54.200 41.700 55.800 ;
        RECT 44.600 55.600 45.000 59.900 ;
        RECT 46.700 56.200 47.100 59.900 ;
        RECT 47.400 56.800 47.800 57.200 ;
        RECT 47.500 56.200 47.800 56.800 ;
        RECT 46.700 55.900 47.200 56.200 ;
        RECT 47.500 55.900 48.200 56.200 ;
        RECT 42.900 55.300 45.000 55.600 ;
        RECT 42.900 55.200 43.300 55.300 ;
        RECT 43.700 54.900 44.100 55.000 ;
        RECT 42.200 54.600 44.100 54.900 ;
        RECT 42.200 54.500 42.600 54.600 ;
        RECT 31.000 54.100 31.400 54.200 ;
        RECT 31.000 53.800 31.800 54.100 ;
        RECT 32.500 53.800 33.800 54.200 ;
        RECT 36.200 53.900 41.700 54.200 ;
        RECT 36.200 53.800 37.000 53.900 ;
        RECT 31.400 53.600 31.800 53.800 ;
        RECT 31.100 53.100 32.900 53.300 ;
        RECT 33.400 53.100 33.700 53.800 ;
        RECT 29.400 52.800 30.300 53.100 ;
        RECT 29.900 51.100 30.300 52.800 ;
        RECT 31.000 53.000 33.000 53.100 ;
        RECT 31.000 51.100 31.400 53.000 ;
        RECT 32.600 51.100 33.000 53.000 ;
        RECT 33.400 51.100 33.800 53.100 ;
        RECT 35.800 51.100 36.200 53.500 ;
        RECT 38.300 52.800 38.600 53.900 ;
        RECT 41.100 53.800 41.500 53.900 ;
        RECT 44.600 53.600 45.000 55.300 ;
        RECT 46.900 55.200 47.200 55.900 ;
        RECT 47.800 55.800 48.200 55.900 ;
        RECT 48.600 55.800 49.000 56.600 ;
        RECT 45.400 55.100 45.800 55.200 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 45.400 54.800 46.600 55.100 ;
        RECT 46.200 54.400 46.600 54.800 ;
        RECT 46.900 54.800 47.400 55.200 ;
        RECT 47.800 55.100 48.100 55.800 ;
        RECT 49.400 55.100 49.800 59.900 ;
        RECT 47.800 54.800 49.800 55.100 ;
        RECT 46.900 54.200 47.200 54.800 ;
        RECT 45.400 54.100 45.800 54.200 ;
        RECT 45.400 53.800 46.200 54.100 ;
        RECT 46.900 53.800 48.200 54.200 ;
        RECT 45.800 53.600 46.200 53.800 ;
        RECT 43.100 53.300 45.000 53.600 ;
        RECT 43.100 53.200 43.500 53.300 ;
        RECT 37.400 52.100 37.800 52.500 ;
        RECT 38.200 52.400 38.600 52.800 ;
        RECT 39.100 52.700 39.500 52.800 ;
        RECT 39.100 52.400 40.500 52.700 ;
        RECT 40.200 52.100 40.500 52.400 ;
        RECT 42.200 52.100 42.600 52.500 ;
        RECT 37.400 51.800 38.400 52.100 ;
        RECT 38.000 51.100 38.400 51.800 ;
        RECT 40.200 51.100 40.600 52.100 ;
        RECT 42.200 51.800 42.900 52.100 ;
        RECT 42.300 51.100 42.900 51.800 ;
        RECT 44.600 51.100 45.000 53.300 ;
        RECT 45.500 53.100 47.300 53.300 ;
        RECT 47.800 53.100 48.100 53.800 ;
        RECT 49.400 53.100 49.800 54.800 ;
        RECT 51.800 55.100 52.200 59.900 ;
        RECT 53.900 59.200 54.300 59.900 ;
        RECT 53.400 58.800 54.300 59.200 ;
        RECT 53.900 56.200 54.300 58.800 ;
        RECT 57.100 57.200 57.500 59.900 ;
        RECT 54.600 56.800 55.000 57.200 ;
        RECT 56.600 56.800 57.500 57.200 ;
        RECT 57.800 56.800 58.200 57.200 ;
        RECT 54.700 56.200 55.000 56.800 ;
        RECT 57.100 56.200 57.500 56.800 ;
        RECT 57.900 56.200 58.200 56.800 ;
        RECT 60.300 56.200 60.700 59.900 ;
        RECT 61.000 56.800 61.400 57.200 ;
        RECT 61.100 56.200 61.400 56.800 ;
        RECT 53.900 55.900 54.400 56.200 ;
        RECT 54.700 55.900 55.400 56.200 ;
        RECT 57.100 55.900 57.600 56.200 ;
        RECT 57.900 55.900 58.600 56.200 ;
        RECT 60.300 55.900 60.800 56.200 ;
        RECT 61.100 55.900 61.800 56.200 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 51.800 54.800 53.000 55.100 ;
        RECT 50.200 53.400 50.600 54.200 ;
        RECT 45.400 53.000 47.400 53.100 ;
        RECT 45.400 51.100 45.800 53.000 ;
        RECT 47.000 51.100 47.400 53.000 ;
        RECT 47.800 51.100 48.200 53.100 ;
        RECT 48.900 52.800 49.800 53.100 ;
        RECT 48.900 51.100 49.300 52.800 ;
        RECT 51.000 52.400 51.400 53.200 ;
        RECT 51.800 51.100 52.200 54.800 ;
        RECT 53.400 54.400 53.800 55.200 ;
        RECT 54.100 54.200 54.400 55.900 ;
        RECT 55.000 55.800 55.400 55.900 ;
        RECT 56.600 54.400 57.000 55.200 ;
        RECT 57.300 54.200 57.600 55.900 ;
        RECT 58.200 55.800 58.600 55.900 ;
        RECT 59.800 54.400 60.200 55.200 ;
        RECT 60.500 54.200 60.800 55.900 ;
        RECT 61.400 55.800 61.800 55.900 ;
        RECT 62.200 55.700 62.600 59.900 ;
        RECT 64.400 58.200 64.800 59.900 ;
        RECT 63.800 57.900 64.800 58.200 ;
        RECT 66.600 57.900 67.000 59.900 ;
        RECT 68.700 57.900 69.300 59.900 ;
        RECT 63.800 57.500 64.200 57.900 ;
        RECT 66.600 57.600 66.900 57.900 ;
        RECT 65.500 57.300 67.300 57.600 ;
        RECT 68.600 57.500 69.000 57.900 ;
        RECT 65.500 57.200 65.900 57.300 ;
        RECT 66.900 57.200 67.300 57.300 ;
        RECT 63.800 56.500 64.200 56.600 ;
        RECT 66.100 56.500 66.500 56.600 ;
        RECT 63.800 56.200 66.500 56.500 ;
        RECT 66.800 56.500 67.900 56.800 ;
        RECT 66.800 55.900 67.100 56.500 ;
        RECT 67.500 56.400 67.900 56.500 ;
        RECT 68.700 56.600 69.400 57.000 ;
        RECT 68.700 56.100 69.000 56.600 ;
        RECT 64.700 55.700 67.100 55.900 ;
        RECT 62.200 55.600 67.100 55.700 ;
        RECT 67.800 55.800 69.000 56.100 ;
        RECT 62.200 55.500 65.100 55.600 ;
        RECT 62.200 55.400 65.000 55.500 ;
        RECT 65.400 55.100 65.800 55.200 ;
        RECT 63.300 54.800 65.800 55.100 ;
        RECT 63.300 54.700 63.700 54.800 ;
        RECT 64.600 54.700 65.000 54.800 ;
        RECT 64.100 54.200 64.500 54.300 ;
        RECT 67.800 54.200 68.100 55.800 ;
        RECT 71.000 55.600 71.400 59.900 ;
        RECT 71.800 56.200 72.200 59.900 ;
        RECT 73.400 56.400 73.800 59.900 ;
        RECT 71.800 55.900 73.100 56.200 ;
        RECT 73.400 55.900 73.900 56.400 ;
        RECT 69.300 55.300 71.400 55.600 ;
        RECT 69.300 55.200 69.700 55.300 ;
        RECT 70.100 54.900 70.500 55.000 ;
        RECT 68.600 54.600 70.500 54.900 ;
        RECT 68.600 54.500 69.000 54.600 ;
        RECT 52.600 54.100 53.000 54.200 ;
        RECT 52.600 53.800 53.400 54.100 ;
        RECT 54.100 53.800 55.400 54.200 ;
        RECT 55.800 54.100 56.200 54.200 ;
        RECT 55.800 53.800 56.600 54.100 ;
        RECT 57.300 53.800 58.600 54.200 ;
        RECT 59.000 54.100 59.400 54.200 ;
        RECT 59.000 53.800 59.800 54.100 ;
        RECT 60.500 53.800 61.800 54.200 ;
        RECT 62.600 53.900 68.100 54.200 ;
        RECT 62.600 53.800 63.400 53.900 ;
        RECT 53.000 53.600 53.400 53.800 ;
        RECT 52.700 53.100 54.500 53.300 ;
        RECT 55.000 53.100 55.300 53.800 ;
        RECT 56.200 53.600 56.600 53.800 ;
        RECT 55.900 53.100 57.700 53.300 ;
        RECT 58.200 53.100 58.500 53.800 ;
        RECT 59.400 53.600 59.800 53.800 ;
        RECT 59.100 53.100 60.900 53.300 ;
        RECT 61.400 53.100 61.700 53.800 ;
        RECT 52.600 53.000 54.600 53.100 ;
        RECT 52.600 51.100 53.000 53.000 ;
        RECT 54.200 51.100 54.600 53.000 ;
        RECT 55.000 51.100 55.400 53.100 ;
        RECT 55.800 53.000 57.800 53.100 ;
        RECT 55.800 51.100 56.200 53.000 ;
        RECT 57.400 51.100 57.800 53.000 ;
        RECT 58.200 51.100 58.600 53.100 ;
        RECT 59.000 53.000 61.000 53.100 ;
        RECT 59.000 51.100 59.400 53.000 ;
        RECT 60.600 51.100 61.000 53.000 ;
        RECT 61.400 51.100 61.800 53.100 ;
        RECT 62.200 51.100 62.600 53.500 ;
        RECT 64.700 52.800 65.000 53.900 ;
        RECT 66.200 53.800 66.600 53.900 ;
        RECT 67.500 53.800 67.900 53.900 ;
        RECT 71.000 53.600 71.400 55.300 ;
        RECT 71.800 54.800 72.300 55.200 ;
        RECT 71.900 54.400 72.300 54.800 ;
        RECT 72.800 54.900 73.100 55.900 ;
        RECT 72.800 54.500 73.300 54.900 ;
        RECT 72.800 53.700 73.100 54.500 ;
        RECT 73.600 54.200 73.900 55.900 ;
        RECT 73.400 53.800 73.900 54.200 ;
        RECT 74.200 54.100 74.600 54.200 ;
        RECT 75.000 54.100 75.400 54.200 ;
        RECT 74.200 53.800 75.400 54.100 ;
        RECT 69.500 53.300 71.400 53.600 ;
        RECT 69.500 53.200 69.900 53.300 ;
        RECT 63.800 52.100 64.200 52.500 ;
        RECT 64.600 52.400 65.000 52.800 ;
        RECT 65.500 52.700 65.900 52.800 ;
        RECT 65.500 52.400 66.900 52.700 ;
        RECT 66.600 52.100 66.900 52.400 ;
        RECT 68.600 52.100 69.000 52.500 ;
        RECT 63.800 51.800 64.800 52.100 ;
        RECT 64.400 51.100 64.800 51.800 ;
        RECT 66.600 51.100 67.000 52.100 ;
        RECT 68.600 51.800 69.300 52.100 ;
        RECT 68.700 51.100 69.300 51.800 ;
        RECT 71.000 51.100 71.400 53.300 ;
        RECT 71.800 53.400 73.100 53.700 ;
        RECT 71.800 51.100 72.200 53.400 ;
        RECT 73.600 53.100 73.900 53.800 ;
        RECT 75.000 53.400 75.400 53.800 ;
        RECT 73.400 52.800 73.900 53.100 ;
        RECT 75.800 53.100 76.200 59.900 ;
        RECT 77.400 57.500 77.800 59.500 ;
        RECT 76.600 55.800 77.000 56.600 ;
        RECT 77.400 55.800 77.700 57.500 ;
        RECT 79.500 56.400 79.900 59.900 ;
        RECT 84.100 59.200 84.500 59.900 ;
        RECT 84.100 58.800 85.000 59.200 ;
        RECT 84.100 56.400 84.500 58.800 ;
        RECT 86.200 57.500 86.600 59.500 ;
        RECT 79.500 56.100 80.300 56.400 ;
        RECT 77.400 55.500 79.300 55.800 ;
        RECT 77.400 54.400 77.800 55.200 ;
        RECT 78.200 54.400 78.600 55.200 ;
        RECT 79.000 54.500 79.300 55.500 ;
        RECT 79.000 54.100 79.700 54.500 ;
        RECT 80.000 54.200 80.300 56.100 ;
        RECT 83.700 56.100 84.500 56.400 ;
        RECT 80.600 54.800 81.000 55.600 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 83.000 54.800 83.400 55.600 ;
        RECT 80.000 54.100 81.000 54.200 ;
        RECT 81.400 54.100 81.700 54.800 ;
        RECT 83.700 54.200 84.000 56.100 ;
        RECT 86.300 55.800 86.600 57.500 ;
        RECT 84.700 55.500 86.600 55.800 ;
        RECT 88.600 57.500 89.000 59.500 ;
        RECT 90.700 59.200 91.100 59.900 ;
        RECT 90.700 58.800 91.400 59.200 ;
        RECT 88.600 55.800 88.900 57.500 ;
        RECT 90.700 56.400 91.100 58.800 ;
        RECT 90.700 56.100 91.500 56.400 ;
        RECT 88.600 55.500 90.500 55.800 ;
        RECT 84.700 54.500 85.000 55.500 ;
        RECT 79.000 53.900 79.500 54.100 ;
        RECT 77.400 53.600 79.500 53.900 ;
        RECT 80.000 53.800 81.700 54.100 ;
        RECT 83.000 53.800 84.000 54.200 ;
        RECT 84.300 54.100 85.000 54.500 ;
        RECT 85.400 54.400 85.800 55.200 ;
        RECT 86.200 55.100 86.600 55.200 ;
        RECT 88.600 55.100 89.000 55.200 ;
        RECT 86.200 54.800 89.000 55.100 ;
        RECT 86.200 54.400 86.600 54.800 ;
        RECT 88.600 54.400 89.000 54.800 ;
        RECT 89.400 54.400 89.800 55.200 ;
        RECT 90.200 54.500 90.500 55.500 ;
        RECT 75.800 52.800 76.700 53.100 ;
        RECT 73.400 51.100 73.800 52.800 ;
        RECT 76.300 52.200 76.700 52.800 ;
        RECT 75.800 51.800 76.700 52.200 ;
        RECT 76.300 51.100 76.700 51.800 ;
        RECT 77.400 52.500 77.700 53.600 ;
        RECT 80.000 53.500 80.300 53.800 ;
        RECT 79.900 53.300 80.300 53.500 ;
        RECT 79.500 53.000 80.300 53.300 ;
        RECT 83.700 53.500 84.000 53.800 ;
        RECT 84.500 53.900 85.000 54.100 ;
        RECT 90.200 54.100 90.900 54.500 ;
        RECT 91.200 54.200 91.500 56.100 ;
        RECT 93.400 55.700 93.800 59.900 ;
        RECT 95.600 58.200 96.000 59.900 ;
        RECT 95.000 57.900 96.000 58.200 ;
        RECT 97.800 57.900 98.200 59.900 ;
        RECT 99.900 57.900 100.500 59.900 ;
        RECT 95.000 57.500 95.400 57.900 ;
        RECT 97.800 57.600 98.100 57.900 ;
        RECT 96.700 57.300 98.500 57.600 ;
        RECT 99.800 57.500 100.200 57.900 ;
        RECT 96.700 57.200 97.100 57.300 ;
        RECT 98.100 57.200 98.500 57.300 ;
        RECT 95.000 56.500 95.400 56.600 ;
        RECT 97.300 56.500 97.700 56.600 ;
        RECT 95.000 56.200 97.700 56.500 ;
        RECT 98.000 56.500 99.100 56.800 ;
        RECT 98.000 55.900 98.300 56.500 ;
        RECT 98.700 56.400 99.100 56.500 ;
        RECT 99.900 56.600 100.600 57.000 ;
        RECT 99.900 56.100 100.200 56.600 ;
        RECT 95.900 55.700 98.300 55.900 ;
        RECT 93.400 55.600 98.300 55.700 ;
        RECT 99.000 55.800 100.200 56.100 ;
        RECT 91.800 54.800 92.200 55.600 ;
        RECT 93.400 55.500 96.300 55.600 ;
        RECT 93.400 55.400 96.200 55.500 ;
        RECT 96.600 55.100 97.000 55.200 ;
        RECT 94.500 54.800 97.000 55.100 ;
        RECT 94.500 54.700 94.900 54.800 ;
        RECT 95.300 54.200 95.700 54.300 ;
        RECT 99.000 54.200 99.300 55.800 ;
        RECT 102.200 55.600 102.600 59.900 ;
        RECT 103.000 55.800 103.400 56.600 ;
        RECT 100.500 55.300 102.600 55.600 ;
        RECT 100.500 55.200 100.900 55.300 ;
        RECT 101.300 54.900 101.700 55.000 ;
        RECT 99.800 54.600 101.700 54.900 ;
        RECT 99.800 54.500 100.200 54.600 ;
        RECT 90.200 53.900 90.700 54.100 ;
        RECT 84.500 53.600 86.600 53.900 ;
        RECT 83.700 53.300 84.100 53.500 ;
        RECT 83.700 53.000 84.500 53.300 ;
        RECT 77.400 51.500 77.800 52.500 ;
        RECT 79.500 51.500 79.900 53.000 ;
        RECT 84.100 51.500 84.500 53.000 ;
        RECT 86.300 52.500 86.600 53.600 ;
        RECT 86.200 51.500 86.600 52.500 ;
        RECT 88.600 53.600 90.700 53.900 ;
        RECT 91.200 53.800 92.200 54.200 ;
        RECT 93.800 53.900 99.300 54.200 ;
        RECT 93.800 53.800 94.600 53.900 ;
        RECT 88.600 52.500 88.900 53.600 ;
        RECT 91.200 53.500 91.500 53.800 ;
        RECT 91.100 53.300 91.500 53.500 ;
        RECT 90.700 53.000 91.500 53.300 ;
        RECT 88.600 51.500 89.000 52.500 ;
        RECT 90.700 51.500 91.100 53.000 ;
        RECT 93.400 51.100 93.800 53.500 ;
        RECT 95.900 52.800 96.200 53.900 ;
        RECT 98.700 53.800 99.100 53.900 ;
        RECT 102.200 53.600 102.600 55.300 ;
        RECT 100.700 53.300 102.600 53.600 ;
        RECT 100.700 53.200 101.100 53.300 ;
        RECT 95.000 52.100 95.400 52.500 ;
        RECT 95.800 52.400 96.200 52.800 ;
        RECT 96.700 52.700 97.100 52.800 ;
        RECT 96.700 52.400 98.100 52.700 ;
        RECT 97.800 52.100 98.100 52.400 ;
        RECT 99.800 52.100 100.200 52.500 ;
        RECT 95.000 51.800 96.000 52.100 ;
        RECT 95.600 51.100 96.000 51.800 ;
        RECT 97.800 51.100 98.200 52.100 ;
        RECT 99.800 51.800 100.500 52.100 ;
        RECT 99.900 51.100 100.500 51.800 ;
        RECT 102.200 51.100 102.600 53.300 ;
        RECT 103.800 53.100 104.200 59.900 ;
        RECT 106.200 57.100 106.600 59.900 ;
        RECT 107.000 57.100 107.400 57.200 ;
        RECT 106.200 56.800 107.400 57.100 ;
        RECT 104.600 56.100 105.000 56.200 ;
        RECT 105.400 56.100 105.800 56.600 ;
        RECT 104.600 55.800 105.800 56.100 ;
        RECT 104.600 53.400 105.000 54.200 ;
        RECT 106.200 53.100 106.600 56.800 ;
        RECT 107.000 53.400 107.400 54.200 ;
        RECT 103.300 52.800 104.200 53.100 ;
        RECT 105.700 52.800 106.600 53.100 ;
        RECT 103.300 51.100 103.700 52.800 ;
        RECT 105.700 51.100 106.100 52.800 ;
        RECT 107.800 52.400 108.200 53.200 ;
        RECT 108.600 51.100 109.000 59.900 ;
        RECT 110.500 59.200 110.900 59.900 ;
        RECT 110.500 58.800 111.400 59.200 ;
        RECT 109.800 56.800 110.200 57.200 ;
        RECT 109.800 56.200 110.100 56.800 ;
        RECT 110.500 56.200 110.900 58.800 ;
        RECT 109.400 55.900 110.100 56.200 ;
        RECT 110.400 55.900 110.900 56.200 ;
        RECT 112.600 56.200 113.000 59.900 ;
        RECT 114.200 56.400 114.600 59.900 ;
        RECT 115.800 57.500 116.200 59.500 ;
        RECT 112.600 55.900 113.900 56.200 ;
        RECT 114.200 55.900 114.700 56.400 ;
        RECT 109.400 55.800 109.800 55.900 ;
        RECT 110.400 54.200 110.700 55.900 ;
        RECT 111.000 54.400 111.400 55.200 ;
        RECT 112.600 54.800 113.100 55.200 ;
        RECT 112.700 54.400 113.100 54.800 ;
        RECT 113.600 54.900 113.900 55.900 ;
        RECT 113.600 54.500 114.100 54.900 ;
        RECT 109.400 53.800 110.700 54.200 ;
        RECT 111.800 54.100 112.200 54.200 ;
        RECT 111.400 53.800 112.200 54.100 ;
        RECT 109.500 53.100 109.800 53.800 ;
        RECT 111.400 53.600 111.800 53.800 ;
        RECT 113.600 53.700 113.900 54.500 ;
        RECT 114.400 54.200 114.700 55.900 ;
        RECT 115.800 55.800 116.100 57.500 ;
        RECT 117.900 57.200 118.300 59.900 ;
        RECT 120.600 57.900 121.000 59.900 ;
        RECT 120.700 57.800 121.000 57.900 ;
        RECT 122.200 57.900 122.600 59.900 ;
        RECT 122.200 57.800 122.500 57.900 ;
        RECT 120.700 57.500 122.500 57.800 ;
        RECT 117.900 56.800 118.600 57.200 ;
        RECT 117.900 56.400 118.300 56.800 ;
        RECT 117.900 56.100 118.700 56.400 ;
        RECT 120.700 56.200 121.000 57.500 ;
        RECT 121.400 56.400 121.800 57.200 ;
        RECT 115.800 55.500 117.700 55.800 ;
        RECT 115.800 55.100 116.200 55.200 ;
        RECT 114.200 54.100 114.700 54.200 ;
        RECT 115.000 54.800 116.200 55.100 ;
        RECT 115.000 54.100 115.300 54.800 ;
        RECT 115.800 54.400 116.200 54.800 ;
        RECT 116.600 54.400 117.000 55.200 ;
        RECT 117.400 54.500 117.700 55.500 ;
        RECT 114.200 53.800 115.300 54.100 ;
        RECT 117.400 54.100 118.100 54.500 ;
        RECT 118.400 54.200 118.700 56.100 ;
        RECT 120.600 55.800 121.000 56.200 ;
        RECT 119.000 55.100 119.400 55.600 ;
        RECT 119.800 55.100 120.200 55.200 ;
        RECT 119.000 54.800 120.200 55.100 ;
        RECT 120.700 54.200 121.000 55.800 ;
        RECT 123.000 55.400 123.400 56.200 ;
        RECT 123.800 55.800 124.200 56.600 ;
        RECT 124.600 56.100 125.000 59.900 ;
        RECT 126.200 56.200 126.600 59.900 ;
        RECT 127.800 56.400 128.200 59.900 ;
        RECT 130.200 57.900 130.600 59.900 ;
        RECT 130.300 57.800 130.600 57.900 ;
        RECT 131.800 57.900 132.200 59.900 ;
        RECT 131.800 57.800 132.100 57.900 ;
        RECT 130.300 57.500 132.100 57.800 ;
        RECT 131.000 56.400 131.400 57.200 ;
        RECT 125.400 56.100 125.800 56.200 ;
        RECT 124.600 55.800 125.800 56.100 ;
        RECT 126.200 55.900 127.500 56.200 ;
        RECT 127.800 55.900 128.300 56.400 ;
        RECT 131.800 56.200 132.100 57.500 ;
        RECT 133.400 57.100 133.800 59.900 ;
        RECT 132.600 56.800 133.800 57.100 ;
        RECT 132.600 56.200 132.900 56.800 ;
        RECT 121.800 54.800 122.600 55.200 ;
        RECT 117.400 53.900 117.900 54.100 ;
        RECT 112.600 53.400 113.900 53.700 ;
        RECT 110.300 53.100 112.100 53.300 ;
        RECT 109.400 51.100 109.800 53.100 ;
        RECT 110.200 53.000 112.200 53.100 ;
        RECT 110.200 51.100 110.600 53.000 ;
        RECT 111.800 51.100 112.200 53.000 ;
        RECT 112.600 51.100 113.000 53.400 ;
        RECT 114.400 53.100 114.700 53.800 ;
        RECT 114.200 52.800 114.700 53.100 ;
        RECT 115.800 53.600 117.900 53.900 ;
        RECT 118.400 53.800 119.400 54.200 ;
        RECT 120.700 54.100 121.500 54.200 ;
        RECT 120.700 53.900 121.600 54.100 ;
        RECT 114.200 51.100 114.600 52.800 ;
        RECT 115.800 52.500 116.100 53.600 ;
        RECT 118.400 53.500 118.700 53.800 ;
        RECT 118.300 53.300 118.700 53.500 ;
        RECT 117.900 53.000 118.700 53.300 ;
        RECT 115.800 51.500 116.200 52.500 ;
        RECT 117.900 51.500 118.300 53.000 ;
        RECT 121.200 51.100 121.600 53.900 ;
        RECT 124.600 53.100 125.000 55.800 ;
        RECT 126.200 54.800 126.700 55.200 ;
        RECT 126.300 54.400 126.700 54.800 ;
        RECT 127.200 54.900 127.500 55.900 ;
        RECT 127.200 54.500 127.700 54.900 ;
        RECT 125.400 53.400 125.800 54.200 ;
        RECT 127.200 53.700 127.500 54.500 ;
        RECT 128.000 54.200 128.300 55.900 ;
        RECT 129.400 55.400 129.800 56.200 ;
        RECT 131.800 55.800 132.200 56.200 ;
        RECT 132.600 55.800 133.000 56.200 ;
        RECT 130.200 54.800 131.000 55.200 ;
        RECT 131.800 54.200 132.100 55.800 ;
        RECT 127.800 53.800 128.300 54.200 ;
        RECT 131.300 54.100 132.100 54.200 ;
        RECT 126.200 53.400 127.500 53.700 ;
        RECT 124.100 52.800 125.000 53.100 ;
        RECT 124.100 51.100 124.500 52.800 ;
        RECT 126.200 51.100 126.600 53.400 ;
        RECT 128.000 53.100 128.300 53.800 ;
        RECT 127.800 52.800 128.300 53.100 ;
        RECT 131.200 53.900 132.100 54.100 ;
        RECT 127.800 51.100 128.200 52.800 ;
        RECT 131.200 51.100 131.600 53.900 ;
        RECT 132.600 53.400 133.000 54.200 ;
        RECT 133.400 53.100 133.800 56.800 ;
        RECT 135.000 57.500 135.400 59.500 ;
        RECT 134.200 55.800 134.600 56.600 ;
        RECT 135.000 55.800 135.300 57.500 ;
        RECT 137.100 56.400 137.500 59.900 ;
        RECT 137.100 56.100 137.900 56.400 ;
        RECT 135.000 55.500 136.900 55.800 ;
        RECT 135.000 54.400 135.400 55.200 ;
        RECT 135.800 54.400 136.200 55.200 ;
        RECT 136.600 54.500 136.900 55.500 ;
        RECT 136.600 54.100 137.300 54.500 ;
        RECT 137.600 54.200 137.900 56.100 ;
        RECT 138.200 54.800 138.600 55.600 ;
        RECT 136.600 53.900 137.100 54.100 ;
        RECT 135.000 53.600 137.100 53.900 ;
        RECT 137.600 53.800 138.600 54.200 ;
        RECT 133.400 52.800 134.300 53.100 ;
        RECT 133.900 51.100 134.300 52.800 ;
        RECT 135.000 52.500 135.300 53.600 ;
        RECT 137.600 53.500 137.900 53.800 ;
        RECT 137.500 53.300 137.900 53.500 ;
        RECT 137.100 53.200 137.900 53.300 ;
        RECT 136.600 53.000 137.900 53.200 ;
        RECT 136.600 52.800 137.500 53.000 ;
        RECT 135.000 51.500 135.400 52.500 ;
        RECT 137.100 51.500 137.500 52.800 ;
        RECT 141.400 51.100 141.800 59.900 ;
        RECT 143.300 59.200 143.700 59.900 ;
        RECT 143.000 58.800 143.700 59.200 ;
        RECT 143.300 56.200 143.700 58.800 ;
        RECT 143.000 55.900 143.700 56.200 ;
        RECT 143.000 55.200 143.300 55.900 ;
        RECT 145.400 55.600 145.800 59.900 ;
        RECT 147.300 59.200 147.700 59.900 ;
        RECT 147.300 58.800 148.200 59.200 ;
        RECT 146.600 56.800 147.000 57.200 ;
        RECT 146.600 56.200 146.900 56.800 ;
        RECT 147.300 56.200 147.700 58.800 ;
        RECT 146.200 55.900 146.900 56.200 ;
        RECT 147.200 55.900 147.700 56.200 ;
        RECT 146.200 55.800 146.600 55.900 ;
        RECT 143.800 55.400 145.800 55.600 ;
        RECT 143.700 55.300 145.800 55.400 ;
        RECT 143.000 54.800 143.400 55.200 ;
        RECT 143.700 55.000 144.100 55.300 ;
        RECT 142.200 52.400 142.600 53.200 ;
        RECT 143.000 53.100 143.300 54.800 ;
        RECT 143.700 53.500 144.000 55.000 ;
        RECT 144.400 54.200 144.800 54.600 ;
        RECT 147.200 54.200 147.500 55.900 ;
        RECT 149.400 55.800 149.800 56.600 ;
        RECT 147.800 54.400 148.200 55.200 ;
        RECT 144.500 53.800 145.000 54.200 ;
        RECT 146.200 53.800 147.500 54.200 ;
        RECT 148.600 54.100 149.000 54.200 ;
        RECT 148.200 53.800 149.000 54.100 ;
        RECT 143.700 53.200 144.900 53.500 ;
        RECT 143.000 51.100 143.400 53.100 ;
        RECT 144.600 52.100 144.900 53.200 ;
        RECT 145.400 52.400 145.800 53.200 ;
        RECT 146.300 53.100 146.600 53.800 ;
        RECT 148.200 53.600 148.600 53.800 ;
        RECT 147.100 53.100 148.900 53.300 ;
        RECT 150.200 53.100 150.600 59.900 ;
        RECT 151.800 55.700 152.200 59.900 ;
        RECT 154.000 58.200 154.400 59.900 ;
        RECT 153.400 57.900 154.400 58.200 ;
        RECT 156.200 57.900 156.600 59.900 ;
        RECT 158.300 57.900 158.900 59.900 ;
        RECT 153.400 57.500 153.800 57.900 ;
        RECT 156.200 57.600 156.500 57.900 ;
        RECT 155.100 57.300 156.900 57.600 ;
        RECT 158.200 57.500 158.600 57.900 ;
        RECT 155.100 57.200 155.500 57.300 ;
        RECT 156.500 57.200 156.900 57.300 ;
        RECT 153.400 56.500 153.800 56.600 ;
        RECT 155.700 56.500 156.100 56.600 ;
        RECT 153.400 56.200 156.100 56.500 ;
        RECT 156.400 56.500 157.500 56.800 ;
        RECT 156.400 55.900 156.700 56.500 ;
        RECT 157.100 56.400 157.500 56.500 ;
        RECT 158.300 56.600 159.000 57.000 ;
        RECT 158.300 56.100 158.600 56.600 ;
        RECT 154.300 55.700 156.700 55.900 ;
        RECT 151.800 55.600 156.700 55.700 ;
        RECT 157.400 55.800 158.600 56.100 ;
        RECT 151.800 55.500 154.700 55.600 ;
        RECT 151.800 55.400 154.600 55.500 ;
        RECT 155.000 55.100 155.400 55.200 ;
        RECT 152.900 54.800 155.400 55.100 ;
        RECT 152.900 54.700 153.300 54.800 ;
        RECT 153.700 54.200 154.100 54.300 ;
        RECT 157.400 54.200 157.700 55.800 ;
        RECT 160.600 55.600 161.000 59.900 ;
        RECT 158.900 55.300 161.000 55.600 ;
        RECT 158.900 55.200 159.300 55.300 ;
        RECT 159.700 54.900 160.100 55.000 ;
        RECT 158.200 54.600 160.100 54.900 ;
        RECT 158.200 54.500 158.600 54.600 ;
        RECT 151.000 53.400 151.400 54.200 ;
        RECT 152.200 53.900 157.700 54.200 ;
        RECT 152.200 53.800 153.000 53.900 ;
        RECT 144.600 51.100 145.000 52.100 ;
        RECT 146.200 51.100 146.600 53.100 ;
        RECT 147.000 53.000 149.000 53.100 ;
        RECT 147.000 51.100 147.400 53.000 ;
        RECT 148.600 51.100 149.000 53.000 ;
        RECT 149.700 52.800 150.600 53.100 ;
        RECT 149.700 52.200 150.100 52.800 ;
        RECT 149.700 51.800 150.600 52.200 ;
        RECT 149.700 51.100 150.100 51.800 ;
        RECT 151.800 51.100 152.200 53.500 ;
        RECT 154.300 53.200 154.600 53.900 ;
        RECT 157.100 53.800 157.700 53.900 ;
        RECT 153.400 52.100 153.800 52.500 ;
        RECT 154.200 52.400 154.600 53.200 ;
        RECT 157.400 53.200 157.700 53.800 ;
        RECT 160.600 53.600 161.000 55.300 ;
        RECT 162.200 55.100 162.600 59.900 ;
        RECT 164.900 57.200 165.300 59.900 ;
        RECT 167.000 57.500 167.400 59.500 ;
        RECT 164.200 56.800 164.600 57.200 ;
        RECT 164.900 56.800 165.800 57.200 ;
        RECT 163.000 55.800 163.400 56.600 ;
        RECT 164.200 56.200 164.500 56.800 ;
        RECT 164.900 56.200 165.300 56.800 ;
        RECT 163.800 55.900 164.500 56.200 ;
        RECT 164.800 55.900 165.300 56.200 ;
        RECT 163.800 55.800 164.200 55.900 ;
        RECT 163.800 55.100 164.100 55.800 ;
        RECT 162.200 54.800 164.100 55.100 ;
        RECT 159.100 53.300 161.000 53.600 ;
        RECT 161.400 53.400 161.800 54.200 ;
        RECT 159.100 53.200 159.500 53.300 ;
        RECT 157.400 52.800 157.800 53.200 ;
        RECT 155.100 52.700 155.500 52.800 ;
        RECT 155.100 52.400 156.500 52.700 ;
        RECT 156.200 52.100 156.500 52.400 ;
        RECT 158.200 52.100 158.600 52.500 ;
        RECT 153.400 51.800 154.400 52.100 ;
        RECT 154.000 51.100 154.400 51.800 ;
        RECT 156.200 51.100 156.600 52.100 ;
        RECT 158.200 51.800 158.900 52.100 ;
        RECT 158.300 51.100 158.900 51.800 ;
        RECT 160.600 51.100 161.000 53.300 ;
        RECT 162.200 53.100 162.600 54.800 ;
        RECT 164.800 54.200 165.100 55.900 ;
        RECT 167.000 55.800 167.300 57.500 ;
        RECT 169.100 56.400 169.500 59.900 ;
        RECT 169.100 56.100 169.900 56.400 ;
        RECT 167.000 55.500 168.900 55.800 ;
        RECT 165.400 54.400 165.800 55.200 ;
        RECT 167.000 54.400 167.400 55.200 ;
        RECT 167.800 54.400 168.200 55.200 ;
        RECT 168.600 54.500 168.900 55.500 ;
        RECT 163.800 53.800 165.100 54.200 ;
        RECT 166.200 54.100 166.600 54.200 ;
        RECT 165.800 53.800 166.600 54.100 ;
        RECT 168.600 54.100 169.300 54.500 ;
        RECT 169.600 54.200 169.900 56.100 ;
        RECT 171.800 55.700 172.200 59.900 ;
        RECT 174.000 58.200 174.400 59.900 ;
        RECT 173.400 57.900 174.400 58.200 ;
        RECT 176.200 57.900 176.600 59.900 ;
        RECT 178.300 57.900 178.900 59.900 ;
        RECT 173.400 57.500 173.800 57.900 ;
        RECT 176.200 57.600 176.500 57.900 ;
        RECT 175.100 57.300 176.900 57.600 ;
        RECT 178.200 57.500 178.600 57.900 ;
        RECT 175.100 57.200 175.500 57.300 ;
        RECT 176.500 57.200 176.900 57.300 ;
        RECT 173.400 56.500 173.800 56.600 ;
        RECT 175.700 56.500 176.100 56.600 ;
        RECT 173.400 56.200 176.100 56.500 ;
        RECT 176.400 56.500 177.500 56.800 ;
        RECT 176.400 55.900 176.700 56.500 ;
        RECT 177.100 56.400 177.500 56.500 ;
        RECT 178.300 56.600 179.000 57.000 ;
        RECT 178.300 56.100 178.600 56.600 ;
        RECT 174.300 55.700 176.700 55.900 ;
        RECT 171.800 55.600 176.700 55.700 ;
        RECT 177.400 55.800 178.600 56.100 ;
        RECT 170.200 54.800 170.600 55.600 ;
        RECT 171.800 55.500 174.700 55.600 ;
        RECT 171.800 55.400 174.600 55.500 ;
        RECT 177.400 55.200 177.700 55.800 ;
        RECT 180.600 55.600 181.000 59.900 ;
        RECT 182.200 56.400 182.600 59.900 ;
        RECT 178.900 55.300 181.000 55.600 ;
        RECT 178.900 55.200 179.300 55.300 ;
        RECT 175.000 55.100 175.400 55.200 ;
        RECT 172.900 54.800 175.400 55.100 ;
        RECT 177.400 54.800 177.800 55.200 ;
        RECT 179.700 54.900 180.100 55.000 ;
        RECT 172.900 54.700 173.300 54.800 ;
        RECT 174.200 54.700 174.600 54.800 ;
        RECT 173.700 54.200 174.100 54.300 ;
        RECT 177.400 54.200 177.700 54.800 ;
        RECT 178.200 54.600 180.100 54.900 ;
        RECT 178.200 54.500 178.600 54.600 ;
        RECT 168.600 53.900 169.100 54.100 ;
        RECT 163.900 53.100 164.200 53.800 ;
        RECT 165.800 53.600 166.200 53.800 ;
        RECT 167.000 53.600 169.100 53.900 ;
        RECT 169.600 53.800 170.600 54.200 ;
        RECT 172.200 53.900 177.700 54.200 ;
        RECT 172.200 53.800 173.000 53.900 ;
        RECT 164.700 53.100 166.500 53.300 ;
        RECT 162.200 52.800 163.100 53.100 ;
        RECT 162.700 51.100 163.100 52.800 ;
        RECT 163.800 51.100 164.200 53.100 ;
        RECT 164.600 53.000 166.600 53.100 ;
        RECT 164.600 51.100 165.000 53.000 ;
        RECT 166.200 51.100 166.600 53.000 ;
        RECT 167.000 52.500 167.300 53.600 ;
        RECT 169.600 53.500 169.900 53.800 ;
        RECT 169.500 53.300 169.900 53.500 ;
        RECT 169.100 53.000 169.900 53.300 ;
        RECT 167.000 51.500 167.400 52.500 ;
        RECT 169.100 52.200 169.500 53.000 ;
        RECT 168.600 51.800 169.500 52.200 ;
        RECT 169.100 51.500 169.500 51.800 ;
        RECT 171.800 51.100 172.200 53.500 ;
        RECT 174.300 52.800 174.600 53.900 ;
        RECT 177.100 53.800 177.500 53.900 ;
        RECT 180.600 53.600 181.000 55.300 ;
        RECT 179.100 53.300 181.000 53.600 ;
        RECT 179.100 53.200 179.500 53.300 ;
        RECT 173.400 52.100 173.800 52.500 ;
        RECT 174.200 52.400 174.600 52.800 ;
        RECT 175.100 52.700 175.500 52.800 ;
        RECT 175.100 52.400 176.500 52.700 ;
        RECT 176.200 52.100 176.500 52.400 ;
        RECT 178.200 52.100 178.600 52.500 ;
        RECT 173.400 51.800 174.400 52.100 ;
        RECT 174.000 51.100 174.400 51.800 ;
        RECT 176.200 51.100 176.600 52.100 ;
        RECT 178.200 51.800 178.900 52.100 ;
        RECT 178.300 51.100 178.900 51.800 ;
        RECT 180.600 51.100 181.000 53.300 ;
        RECT 182.100 55.900 182.600 56.400 ;
        RECT 183.800 56.200 184.200 59.900 ;
        RECT 182.900 55.900 184.200 56.200 ;
        RECT 184.600 57.500 185.000 59.500 ;
        RECT 186.700 59.200 187.100 59.900 ;
        RECT 186.200 58.800 187.100 59.200 ;
        RECT 182.100 54.200 182.400 55.900 ;
        RECT 182.900 54.900 183.200 55.900 ;
        RECT 184.600 55.800 184.900 57.500 ;
        RECT 186.700 56.400 187.100 58.800 ;
        RECT 186.700 56.100 187.500 56.400 ;
        RECT 184.600 55.500 186.500 55.800 ;
        RECT 182.700 54.500 183.200 54.900 ;
        RECT 182.100 53.800 182.600 54.200 ;
        RECT 182.100 53.100 182.400 53.800 ;
        RECT 182.900 53.700 183.200 54.500 ;
        RECT 183.700 54.800 184.200 55.200 ;
        RECT 183.700 54.400 184.100 54.800 ;
        RECT 184.600 54.400 185.000 55.200 ;
        RECT 185.400 54.400 185.800 55.200 ;
        RECT 186.200 54.500 186.500 55.500 ;
        RECT 186.200 54.100 186.900 54.500 ;
        RECT 187.200 54.200 187.500 56.100 ;
        RECT 187.800 55.100 188.200 55.600 ;
        RECT 189.400 55.100 189.800 55.200 ;
        RECT 187.800 54.800 189.800 55.100 ;
        RECT 190.200 55.100 190.600 59.900 ;
        RECT 193.800 56.800 194.200 57.200 ;
        RECT 191.000 55.800 191.400 56.600 ;
        RECT 193.800 56.200 194.100 56.800 ;
        RECT 194.500 56.200 194.900 59.900 ;
        RECT 193.400 55.900 194.100 56.200 ;
        RECT 194.400 55.900 194.900 56.200 ;
        RECT 196.600 56.200 197.000 59.900 ;
        RECT 198.200 56.400 198.600 59.900 ;
        RECT 196.600 55.900 197.900 56.200 ;
        RECT 198.200 55.900 198.700 56.400 ;
        RECT 193.400 55.800 193.800 55.900 ;
        RECT 193.400 55.100 193.700 55.800 ;
        RECT 190.200 54.800 193.700 55.100 ;
        RECT 186.200 53.900 186.700 54.100 ;
        RECT 182.900 53.400 184.200 53.700 ;
        RECT 182.100 52.800 182.600 53.100 ;
        RECT 182.200 51.100 182.600 52.800 ;
        RECT 183.800 51.100 184.200 53.400 ;
        RECT 184.600 53.600 186.700 53.900 ;
        RECT 187.200 53.800 188.200 54.200 ;
        RECT 184.600 52.500 184.900 53.600 ;
        RECT 187.200 53.500 187.500 53.800 ;
        RECT 187.100 53.300 187.500 53.500 ;
        RECT 189.400 53.400 189.800 54.200 ;
        RECT 186.700 53.000 187.500 53.300 ;
        RECT 190.200 53.100 190.600 54.800 ;
        RECT 194.400 54.200 194.700 55.900 ;
        RECT 195.000 54.400 195.400 55.200 ;
        RECT 196.600 54.800 197.100 55.200 ;
        RECT 196.700 54.400 197.100 54.800 ;
        RECT 197.600 54.900 197.900 55.900 ;
        RECT 197.600 54.500 198.100 54.900 ;
        RECT 193.400 53.800 194.700 54.200 ;
        RECT 195.800 54.100 196.200 54.200 ;
        RECT 195.400 53.800 196.200 54.100 ;
        RECT 193.500 53.100 193.800 53.800 ;
        RECT 195.400 53.600 195.800 53.800 ;
        RECT 197.600 53.700 197.900 54.500 ;
        RECT 198.400 54.200 198.700 55.900 ;
        RECT 198.200 53.800 198.700 54.200 ;
        RECT 196.600 53.400 197.900 53.700 ;
        RECT 194.300 53.100 196.100 53.300 ;
        RECT 184.600 51.500 185.000 52.500 ;
        RECT 186.700 51.500 187.100 53.000 ;
        RECT 190.200 52.800 191.100 53.100 ;
        RECT 190.700 51.100 191.100 52.800 ;
        RECT 193.400 51.100 193.800 53.100 ;
        RECT 194.200 53.000 196.200 53.100 ;
        RECT 194.200 51.100 194.600 53.000 ;
        RECT 195.800 51.100 196.200 53.000 ;
        RECT 196.600 51.100 197.000 53.400 ;
        RECT 198.400 53.100 198.700 53.800 ;
        RECT 198.200 52.800 198.700 53.100 ;
        RECT 198.200 51.100 198.600 52.800 ;
        RECT 199.800 51.100 200.200 59.900 ;
        RECT 201.400 57.500 201.800 59.500 ;
        RECT 201.400 55.800 201.700 57.500 ;
        RECT 203.500 56.400 203.900 59.900 ;
        RECT 206.200 57.500 206.600 59.500 ;
        RECT 203.500 56.100 204.300 56.400 ;
        RECT 201.400 55.500 203.300 55.800 ;
        RECT 201.400 54.400 201.800 55.200 ;
        RECT 202.200 54.400 202.600 55.200 ;
        RECT 203.000 54.500 203.300 55.500 ;
        RECT 203.000 54.100 203.700 54.500 ;
        RECT 204.000 54.200 204.300 56.100 ;
        RECT 206.200 55.800 206.500 57.500 ;
        RECT 208.300 56.400 208.700 59.900 ;
        RECT 211.800 56.400 212.200 59.900 ;
        RECT 208.300 56.100 209.100 56.400 ;
        RECT 204.600 54.800 205.000 55.600 ;
        RECT 206.200 55.500 208.100 55.800 ;
        RECT 206.200 54.400 206.600 55.200 ;
        RECT 207.000 54.400 207.400 55.200 ;
        RECT 207.800 54.500 208.100 55.500 ;
        RECT 208.800 55.200 209.100 56.100 ;
        RECT 211.700 55.900 212.200 56.400 ;
        RECT 213.400 56.200 213.800 59.900 ;
        RECT 212.500 55.900 213.800 56.200 ;
        RECT 215.500 56.200 215.900 59.900 ;
        RECT 216.200 56.800 216.600 57.200 ;
        RECT 216.300 56.200 216.600 56.800 ;
        RECT 215.500 55.900 216.000 56.200 ;
        RECT 216.300 55.900 217.000 56.200 ;
        RECT 208.600 54.800 209.100 55.200 ;
        RECT 209.400 55.100 209.800 55.600 ;
        RECT 211.000 55.100 211.400 55.200 ;
        RECT 209.400 54.800 211.400 55.100 ;
        RECT 203.000 53.900 203.500 54.100 ;
        RECT 201.400 53.600 203.500 53.900 ;
        RECT 204.000 53.800 205.000 54.200 ;
        RECT 207.800 54.100 208.500 54.500 ;
        RECT 208.800 54.200 209.100 54.800 ;
        RECT 211.700 54.200 212.000 55.900 ;
        RECT 212.500 54.900 212.800 55.900 ;
        RECT 212.300 54.500 212.800 54.900 ;
        RECT 207.800 53.900 208.300 54.100 ;
        RECT 200.600 52.400 201.000 53.200 ;
        RECT 201.400 52.500 201.700 53.600 ;
        RECT 204.000 53.500 204.300 53.800 ;
        RECT 203.900 53.300 204.300 53.500 ;
        RECT 203.500 53.200 204.300 53.300 ;
        RECT 203.000 53.000 204.300 53.200 ;
        RECT 206.200 53.600 208.300 53.900 ;
        RECT 208.800 53.800 209.800 54.200 ;
        RECT 211.700 53.800 212.200 54.200 ;
        RECT 203.000 52.800 203.900 53.000 ;
        RECT 201.400 51.500 201.800 52.500 ;
        RECT 203.500 51.500 203.900 52.800 ;
        RECT 206.200 52.500 206.500 53.600 ;
        RECT 208.800 53.500 209.100 53.800 ;
        RECT 208.700 53.300 209.100 53.500 ;
        RECT 208.300 53.000 209.100 53.300 ;
        RECT 211.700 53.100 212.000 53.800 ;
        RECT 212.500 53.700 212.800 54.500 ;
        RECT 213.300 54.800 213.800 55.200 ;
        RECT 213.300 54.400 213.700 54.800 ;
        RECT 215.000 54.400 215.400 55.200 ;
        RECT 215.700 55.100 216.000 55.900 ;
        RECT 216.600 55.800 217.000 55.900 ;
        RECT 217.400 55.600 217.800 59.900 ;
        RECT 219.500 57.900 220.100 59.900 ;
        RECT 221.800 57.900 222.200 59.900 ;
        RECT 224.000 58.200 224.400 59.900 ;
        RECT 224.000 57.900 225.000 58.200 ;
        RECT 219.800 57.500 220.200 57.900 ;
        RECT 221.900 57.600 222.200 57.900 ;
        RECT 221.500 57.300 223.300 57.600 ;
        RECT 224.600 57.500 225.000 57.900 ;
        RECT 221.500 57.200 221.900 57.300 ;
        RECT 222.900 57.200 223.300 57.300 ;
        RECT 219.400 56.600 220.100 57.000 ;
        RECT 219.800 56.100 220.100 56.600 ;
        RECT 220.900 56.500 222.000 56.800 ;
        RECT 220.900 56.400 221.300 56.500 ;
        RECT 219.800 55.800 221.000 56.100 ;
        RECT 217.400 55.300 219.500 55.600 ;
        RECT 216.600 55.100 217.000 55.200 ;
        RECT 215.700 54.800 217.000 55.100 ;
        RECT 215.700 54.200 216.000 54.800 ;
        RECT 214.200 54.100 214.600 54.200 ;
        RECT 214.200 53.800 215.000 54.100 ;
        RECT 215.700 53.800 217.000 54.200 ;
        RECT 212.500 53.400 213.800 53.700 ;
        RECT 214.600 53.600 215.000 53.800 ;
        RECT 206.200 51.500 206.600 52.500 ;
        RECT 208.300 51.500 208.700 53.000 ;
        RECT 211.700 52.800 212.200 53.100 ;
        RECT 211.800 51.100 212.200 52.800 ;
        RECT 213.400 51.100 213.800 53.400 ;
        RECT 214.300 53.100 216.100 53.300 ;
        RECT 216.600 53.100 216.900 53.800 ;
        RECT 217.400 53.600 217.800 55.300 ;
        RECT 219.100 55.200 219.500 55.300 ;
        RECT 218.300 54.900 218.700 55.000 ;
        RECT 218.300 54.600 220.200 54.900 ;
        RECT 219.800 54.500 220.200 54.600 ;
        RECT 220.700 54.200 221.000 55.800 ;
        RECT 221.700 55.900 222.000 56.500 ;
        RECT 222.300 56.500 222.700 56.600 ;
        RECT 224.600 56.500 225.000 56.600 ;
        RECT 222.300 56.200 225.000 56.500 ;
        RECT 221.700 55.700 224.100 55.900 ;
        RECT 226.200 55.700 226.600 59.900 ;
        RECT 227.000 56.200 227.400 59.900 ;
        RECT 228.600 56.400 229.000 59.900 ;
        RECT 227.000 55.900 228.300 56.200 ;
        RECT 228.600 55.900 229.100 56.400 ;
        RECT 221.700 55.600 226.600 55.700 ;
        RECT 223.700 55.500 226.600 55.600 ;
        RECT 223.800 55.400 226.600 55.500 ;
        RECT 222.200 55.100 222.600 55.200 ;
        RECT 223.000 55.100 223.400 55.200 ;
        RECT 222.200 54.800 225.500 55.100 ;
        RECT 227.000 54.800 227.500 55.200 ;
        RECT 225.100 54.700 225.500 54.800 ;
        RECT 227.100 54.400 227.500 54.800 ;
        RECT 228.000 54.900 228.300 55.900 ;
        RECT 228.000 54.500 228.500 54.900 ;
        RECT 224.300 54.200 224.700 54.300 ;
        RECT 220.700 53.900 226.200 54.200 ;
        RECT 220.900 53.800 221.300 53.900 ;
        RECT 217.400 53.300 219.300 53.600 ;
        RECT 214.200 53.000 216.200 53.100 ;
        RECT 214.200 51.100 214.600 53.000 ;
        RECT 215.800 51.100 216.200 53.000 ;
        RECT 216.600 51.100 217.000 53.100 ;
        RECT 217.400 51.100 217.800 53.300 ;
        RECT 218.900 53.200 219.300 53.300 ;
        RECT 223.800 52.800 224.100 53.900 ;
        RECT 225.400 53.800 226.200 53.900 ;
        RECT 228.000 53.700 228.300 54.500 ;
        RECT 228.800 54.200 229.100 55.900 ;
        RECT 228.600 54.100 229.100 54.200 ;
        RECT 229.400 54.100 229.800 54.200 ;
        RECT 228.600 53.800 229.800 54.100 ;
        RECT 222.900 52.700 223.300 52.800 ;
        RECT 219.800 52.100 220.200 52.500 ;
        RECT 221.900 52.400 223.300 52.700 ;
        RECT 223.800 52.400 224.200 52.800 ;
        RECT 221.900 52.100 222.200 52.400 ;
        RECT 224.600 52.100 225.000 52.500 ;
        RECT 219.500 51.800 220.200 52.100 ;
        RECT 219.500 51.100 220.100 51.800 ;
        RECT 221.800 51.100 222.200 52.100 ;
        RECT 224.000 51.800 225.000 52.100 ;
        RECT 224.000 51.100 224.400 51.800 ;
        RECT 226.200 51.100 226.600 53.500 ;
        RECT 227.000 53.400 228.300 53.700 ;
        RECT 227.000 51.100 227.400 53.400 ;
        RECT 228.800 53.100 229.100 53.800 ;
        RECT 228.600 52.800 229.100 53.100 ;
        RECT 228.600 51.100 229.000 52.800 ;
        RECT 0.600 47.500 1.000 49.900 ;
        RECT 2.800 49.200 3.200 49.900 ;
        RECT 2.200 48.900 3.200 49.200 ;
        RECT 5.000 48.900 5.400 49.900 ;
        RECT 7.100 49.200 7.700 49.900 ;
        RECT 7.000 48.900 7.700 49.200 ;
        RECT 2.200 48.500 2.600 48.900 ;
        RECT 5.000 48.600 5.300 48.900 ;
        RECT 3.000 48.200 3.400 48.600 ;
        RECT 3.900 48.300 5.300 48.600 ;
        RECT 7.000 48.500 7.400 48.900 ;
        RECT 3.900 48.200 4.300 48.300 ;
        RECT 1.000 47.100 1.800 47.200 ;
        RECT 3.100 47.100 3.400 48.200 ;
        RECT 7.900 47.700 8.300 47.800 ;
        RECT 9.400 47.700 9.800 49.900 ;
        RECT 11.500 48.200 11.900 49.900 ;
        RECT 7.900 47.400 9.800 47.700 ;
        RECT 11.000 47.900 11.900 48.200 ;
        RECT 5.900 47.100 6.300 47.200 ;
        RECT 9.400 47.100 9.800 47.400 ;
        RECT 10.200 47.100 10.600 47.600 ;
        RECT 1.000 46.800 6.500 47.100 ;
        RECT 2.500 46.700 2.900 46.800 ;
        RECT 1.700 46.200 2.100 46.300 ;
        RECT 6.200 46.200 6.500 46.800 ;
        RECT 9.400 46.800 10.600 47.100 ;
        RECT 7.000 46.400 7.400 46.500 ;
        RECT 1.700 45.900 4.200 46.200 ;
        RECT 3.800 45.800 4.200 45.900 ;
        RECT 6.200 45.800 6.600 46.200 ;
        RECT 7.000 46.100 8.900 46.400 ;
        RECT 8.500 46.000 8.900 46.100 ;
        RECT 0.600 45.500 3.400 45.600 ;
        RECT 0.600 45.400 3.500 45.500 ;
        RECT 0.600 45.300 5.500 45.400 ;
        RECT 0.600 41.100 1.000 45.300 ;
        RECT 3.100 45.100 5.500 45.300 ;
        RECT 2.200 44.500 4.900 44.800 ;
        RECT 2.200 44.400 2.600 44.500 ;
        RECT 4.500 44.400 4.900 44.500 ;
        RECT 5.200 44.500 5.500 45.100 ;
        RECT 6.200 45.200 6.500 45.800 ;
        RECT 7.700 45.700 8.100 45.800 ;
        RECT 9.400 45.700 9.800 46.800 ;
        RECT 10.200 46.200 10.500 46.800 ;
        RECT 10.200 45.800 10.600 46.200 ;
        RECT 11.000 46.100 11.400 47.900 ;
        RECT 12.600 47.800 13.000 49.900 ;
        RECT 13.400 48.000 13.800 49.900 ;
        RECT 15.000 48.000 15.400 49.900 ;
        RECT 17.100 49.200 17.500 49.900 ;
        RECT 17.100 48.800 17.800 49.200 ;
        RECT 17.100 48.200 17.500 48.800 ;
        RECT 13.400 47.900 15.400 48.000 ;
        RECT 16.600 47.900 17.500 48.200 ;
        RECT 12.700 47.200 13.000 47.800 ;
        RECT 13.500 47.700 15.300 47.900 ;
        RECT 14.600 47.200 15.000 47.400 ;
        RECT 12.600 46.800 13.900 47.200 ;
        RECT 14.600 46.900 15.400 47.200 ;
        RECT 15.000 46.800 15.400 46.900 ;
        RECT 15.800 46.800 16.200 47.600 ;
        RECT 11.000 45.800 12.900 46.100 ;
        RECT 7.700 45.400 9.800 45.700 ;
        RECT 6.200 44.900 7.400 45.200 ;
        RECT 5.900 44.500 6.300 44.600 ;
        RECT 5.200 44.200 6.300 44.500 ;
        RECT 7.100 44.400 7.400 44.900 ;
        RECT 7.100 44.000 7.800 44.400 ;
        RECT 3.900 43.700 4.300 43.800 ;
        RECT 5.300 43.700 5.700 43.800 ;
        RECT 2.200 43.100 2.600 43.500 ;
        RECT 3.900 43.400 5.700 43.700 ;
        RECT 5.000 43.100 5.300 43.400 ;
        RECT 7.000 43.100 7.400 43.500 ;
        RECT 2.200 42.800 3.200 43.100 ;
        RECT 2.800 41.100 3.200 42.800 ;
        RECT 5.000 41.100 5.400 43.100 ;
        RECT 7.100 41.100 7.700 43.100 ;
        RECT 9.400 41.100 9.800 45.400 ;
        RECT 11.000 41.100 11.400 45.800 ;
        RECT 12.600 45.200 12.900 45.800 ;
        RECT 11.800 44.400 12.200 45.200 ;
        RECT 12.600 45.100 13.000 45.200 ;
        RECT 13.600 45.100 13.900 46.800 ;
        RECT 14.200 45.800 14.600 46.600 ;
        RECT 12.600 44.800 13.300 45.100 ;
        RECT 13.600 44.800 14.100 45.100 ;
        RECT 13.000 44.200 13.300 44.800 ;
        RECT 13.000 43.800 13.400 44.200 ;
        RECT 13.700 41.100 14.100 44.800 ;
        RECT 16.600 41.100 17.000 47.900 ;
        RECT 18.200 47.500 18.600 49.900 ;
        RECT 20.400 49.200 20.800 49.900 ;
        RECT 19.800 48.900 20.800 49.200 ;
        RECT 22.600 48.900 23.000 49.900 ;
        RECT 24.700 49.200 25.300 49.900 ;
        RECT 24.600 48.900 25.300 49.200 ;
        RECT 19.800 48.500 20.200 48.900 ;
        RECT 22.600 48.600 22.900 48.900 ;
        RECT 20.600 48.200 21.000 48.600 ;
        RECT 21.500 48.300 22.900 48.600 ;
        RECT 24.600 48.500 25.000 48.900 ;
        RECT 21.500 48.200 21.900 48.300 ;
        RECT 18.600 47.100 19.400 47.200 ;
        RECT 20.700 47.100 21.000 48.200 ;
        RECT 25.500 47.700 25.900 47.800 ;
        RECT 27.000 47.700 27.400 49.900 ;
        RECT 29.100 48.200 29.500 49.900 ;
        RECT 25.500 47.400 27.400 47.700 ;
        RECT 28.600 47.900 29.500 48.200 ;
        RECT 21.400 47.100 21.800 47.200 ;
        RECT 23.500 47.100 23.900 47.200 ;
        RECT 27.000 47.100 27.400 47.400 ;
        RECT 27.800 47.100 28.200 47.600 ;
        RECT 18.600 46.800 24.100 47.100 ;
        RECT 20.100 46.700 20.500 46.800 ;
        RECT 19.300 46.200 19.700 46.300 ;
        RECT 19.300 46.100 21.800 46.200 ;
        RECT 22.200 46.100 22.600 46.200 ;
        RECT 19.300 45.900 22.600 46.100 ;
        RECT 21.400 45.800 22.600 45.900 ;
        RECT 18.200 45.500 21.000 45.600 ;
        RECT 18.200 45.400 21.100 45.500 ;
        RECT 18.200 45.300 23.100 45.400 ;
        RECT 17.400 44.400 17.800 45.200 ;
        RECT 18.200 41.100 18.600 45.300 ;
        RECT 20.700 45.100 23.100 45.300 ;
        RECT 19.800 44.500 22.500 44.800 ;
        RECT 19.800 44.400 20.200 44.500 ;
        RECT 22.100 44.400 22.500 44.500 ;
        RECT 22.800 44.500 23.100 45.100 ;
        RECT 23.800 45.200 24.100 46.800 ;
        RECT 27.000 46.800 28.200 47.100 ;
        RECT 24.600 46.400 25.000 46.500 ;
        RECT 24.600 46.100 26.500 46.400 ;
        RECT 26.100 46.000 26.500 46.100 ;
        RECT 25.300 45.700 25.700 45.800 ;
        RECT 27.000 45.700 27.400 46.800 ;
        RECT 25.300 45.400 27.400 45.700 ;
        RECT 23.800 44.900 25.000 45.200 ;
        RECT 23.500 44.500 23.900 44.600 ;
        RECT 22.800 44.200 23.900 44.500 ;
        RECT 24.700 44.400 25.000 44.900 ;
        RECT 24.700 44.000 25.400 44.400 ;
        RECT 21.500 43.700 21.900 43.800 ;
        RECT 22.900 43.700 23.300 43.800 ;
        RECT 19.800 43.100 20.200 43.500 ;
        RECT 21.500 43.400 23.300 43.700 ;
        RECT 22.600 43.100 22.900 43.400 ;
        RECT 24.600 43.100 25.000 43.500 ;
        RECT 19.800 42.800 20.800 43.100 ;
        RECT 20.400 41.100 20.800 42.800 ;
        RECT 22.600 41.100 23.000 43.100 ;
        RECT 24.700 41.100 25.300 43.100 ;
        RECT 27.000 41.100 27.400 45.400 ;
        RECT 28.600 46.100 29.000 47.900 ;
        RECT 30.200 47.800 30.600 49.900 ;
        RECT 31.000 48.000 31.400 49.900 ;
        RECT 32.600 48.000 33.000 49.900 ;
        RECT 34.700 49.200 35.100 49.900 ;
        RECT 34.200 48.800 35.100 49.200 ;
        RECT 34.700 48.200 35.100 48.800 ;
        RECT 31.000 47.900 33.000 48.000 ;
        RECT 34.200 47.900 35.100 48.200 ;
        RECT 30.300 47.200 30.600 47.800 ;
        RECT 31.100 47.700 32.900 47.900 ;
        RECT 32.200 47.200 32.600 47.400 ;
        RECT 30.200 46.800 31.500 47.200 ;
        RECT 32.200 46.900 33.000 47.200 ;
        RECT 32.600 46.800 33.000 46.900 ;
        RECT 33.400 46.800 33.800 47.600 ;
        RECT 28.600 45.800 30.500 46.100 ;
        RECT 28.600 41.100 29.000 45.800 ;
        RECT 30.200 45.200 30.500 45.800 ;
        RECT 29.400 44.400 29.800 45.200 ;
        RECT 30.200 45.100 30.600 45.200 ;
        RECT 31.200 45.100 31.500 46.800 ;
        RECT 31.800 46.100 32.200 46.600 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 31.800 45.800 33.000 46.100 ;
        RECT 30.200 44.800 30.900 45.100 ;
        RECT 31.200 44.800 31.700 45.100 ;
        RECT 30.600 44.200 30.900 44.800 ;
        RECT 30.600 43.800 31.000 44.200 ;
        RECT 31.300 41.100 31.700 44.800 ;
        RECT 34.200 41.100 34.600 47.900 ;
        RECT 37.400 47.500 37.800 49.900 ;
        RECT 39.600 49.200 40.000 49.900 ;
        RECT 39.000 48.900 40.000 49.200 ;
        RECT 41.800 48.900 42.200 49.900 ;
        RECT 43.900 49.200 44.500 49.900 ;
        RECT 43.800 48.900 44.500 49.200 ;
        RECT 39.000 48.500 39.400 48.900 ;
        RECT 41.800 48.600 42.100 48.900 ;
        RECT 39.800 48.200 40.200 48.600 ;
        RECT 40.700 48.300 42.100 48.600 ;
        RECT 43.800 48.500 44.200 48.900 ;
        RECT 40.700 48.200 41.100 48.300 ;
        RECT 39.900 47.200 40.200 48.200 ;
        RECT 44.700 47.700 45.100 47.800 ;
        RECT 46.200 47.700 46.600 49.900 ;
        RECT 47.000 48.000 47.400 49.900 ;
        RECT 48.600 48.000 49.000 49.900 ;
        RECT 47.000 47.900 49.000 48.000 ;
        RECT 49.400 47.900 49.800 49.900 ;
        RECT 50.500 48.200 50.900 49.900 ;
        RECT 50.500 47.900 51.400 48.200 ;
        RECT 47.100 47.700 48.900 47.900 ;
        RECT 44.700 47.400 46.600 47.700 ;
        RECT 37.800 47.100 38.600 47.200 ;
        RECT 39.800 47.100 40.200 47.200 ;
        RECT 42.700 47.100 43.100 47.200 ;
        RECT 37.800 46.800 43.300 47.100 ;
        RECT 39.300 46.700 39.700 46.800 ;
        RECT 38.500 46.200 38.900 46.300 ;
        RECT 38.500 45.900 41.000 46.200 ;
        RECT 40.600 45.800 41.000 45.900 ;
        RECT 37.400 45.500 40.200 45.600 ;
        RECT 37.400 45.400 40.300 45.500 ;
        RECT 37.400 45.300 42.300 45.400 ;
        RECT 35.000 44.400 35.400 45.200 ;
        RECT 37.400 41.100 37.800 45.300 ;
        RECT 39.900 45.100 42.300 45.300 ;
        RECT 39.000 44.500 41.700 44.800 ;
        RECT 39.000 44.400 39.400 44.500 ;
        RECT 41.300 44.400 41.700 44.500 ;
        RECT 42.000 44.500 42.300 45.100 ;
        RECT 43.000 45.200 43.300 46.800 ;
        RECT 43.800 46.400 44.200 46.500 ;
        RECT 43.800 46.100 45.700 46.400 ;
        RECT 45.300 46.000 45.700 46.100 ;
        RECT 44.500 45.700 44.900 45.800 ;
        RECT 46.200 45.700 46.600 47.400 ;
        RECT 47.400 47.200 47.800 47.400 ;
        RECT 49.400 47.200 49.700 47.900 ;
        RECT 47.000 46.900 47.800 47.200 ;
        RECT 47.000 46.800 47.400 46.900 ;
        RECT 48.500 46.800 49.800 47.200 ;
        RECT 47.800 45.800 48.200 46.600 ;
        RECT 48.500 46.200 48.800 46.800 ;
        RECT 48.500 45.800 49.000 46.200 ;
        RECT 51.000 46.100 51.400 47.900 ;
        RECT 52.600 47.700 53.000 49.900 ;
        RECT 54.700 49.200 55.300 49.900 ;
        RECT 54.700 48.900 55.400 49.200 ;
        RECT 57.000 48.900 57.400 49.900 ;
        RECT 59.200 49.200 59.600 49.900 ;
        RECT 59.200 48.900 60.200 49.200 ;
        RECT 55.000 48.500 55.400 48.900 ;
        RECT 57.100 48.600 57.400 48.900 ;
        RECT 57.100 48.300 58.500 48.600 ;
        RECT 58.100 48.200 58.500 48.300 ;
        RECT 59.000 48.200 59.400 48.600 ;
        RECT 59.800 48.500 60.200 48.900 ;
        RECT 54.100 47.700 54.500 47.800 ;
        RECT 51.800 46.800 52.200 47.600 ;
        RECT 52.600 47.400 54.500 47.700 ;
        RECT 49.400 45.800 51.400 46.100 ;
        RECT 44.500 45.400 46.600 45.700 ;
        RECT 43.000 44.900 44.200 45.200 ;
        RECT 42.700 44.500 43.100 44.600 ;
        RECT 42.000 44.200 43.100 44.500 ;
        RECT 43.900 44.400 44.200 44.900 ;
        RECT 43.900 44.200 44.600 44.400 ;
        RECT 43.900 44.000 45.000 44.200 ;
        RECT 44.300 43.800 45.000 44.000 ;
        RECT 40.700 43.700 41.100 43.800 ;
        RECT 42.100 43.700 42.500 43.800 ;
        RECT 39.000 43.100 39.400 43.500 ;
        RECT 40.700 43.400 42.500 43.700 ;
        RECT 41.800 43.100 42.100 43.400 ;
        RECT 43.800 43.100 44.200 43.500 ;
        RECT 39.000 42.800 40.000 43.100 ;
        RECT 39.600 41.100 40.000 42.800 ;
        RECT 41.800 41.100 42.200 43.100 ;
        RECT 43.900 41.100 44.500 43.100 ;
        RECT 46.200 41.100 46.600 45.400 ;
        RECT 48.500 45.100 48.800 45.800 ;
        RECT 49.400 45.200 49.700 45.800 ;
        RECT 49.400 45.100 49.800 45.200 ;
        RECT 48.300 44.800 48.800 45.100 ;
        RECT 49.100 44.800 49.800 45.100 ;
        RECT 48.300 41.100 48.700 44.800 ;
        RECT 49.100 44.200 49.400 44.800 ;
        RECT 50.200 44.400 50.600 45.200 ;
        RECT 49.000 43.800 49.400 44.200 ;
        RECT 51.000 41.100 51.400 45.800 ;
        RECT 52.600 45.700 53.000 47.400 ;
        RECT 56.100 47.100 56.500 47.200 ;
        RECT 59.000 47.100 59.300 48.200 ;
        RECT 61.400 47.500 61.800 49.900 ;
        RECT 62.200 47.900 62.600 49.900 ;
        RECT 63.000 48.000 63.400 49.900 ;
        RECT 64.600 48.000 65.000 49.900 ;
        RECT 63.000 47.900 65.000 48.000 ;
        RECT 62.300 47.200 62.600 47.900 ;
        RECT 63.100 47.700 64.900 47.900 ;
        RECT 65.400 47.500 65.800 49.900 ;
        RECT 67.600 49.200 68.000 49.900 ;
        RECT 67.000 48.900 68.000 49.200 ;
        RECT 69.800 48.900 70.200 49.900 ;
        RECT 71.900 49.200 72.500 49.900 ;
        RECT 71.800 48.900 72.500 49.200 ;
        RECT 67.000 48.500 67.400 48.900 ;
        RECT 69.800 48.600 70.100 48.900 ;
        RECT 67.800 48.200 68.200 48.600 ;
        RECT 68.700 48.300 70.100 48.600 ;
        RECT 71.800 48.500 72.200 48.900 ;
        RECT 68.700 48.200 69.100 48.300 ;
        RECT 64.200 47.200 64.600 47.400 ;
        RECT 60.600 47.100 61.400 47.200 ;
        RECT 55.900 46.800 61.400 47.100 ;
        RECT 62.200 46.800 63.500 47.200 ;
        RECT 64.200 46.900 65.000 47.200 ;
        RECT 64.600 46.800 65.000 46.900 ;
        RECT 65.800 47.100 66.600 47.200 ;
        RECT 67.900 47.100 68.200 48.200 ;
        RECT 72.700 47.700 73.100 47.800 ;
        RECT 74.200 47.700 74.600 49.900 ;
        RECT 75.000 47.900 75.400 49.900 ;
        RECT 75.800 48.000 76.200 49.900 ;
        RECT 77.400 48.000 77.800 49.900 ;
        RECT 75.800 47.900 77.800 48.000 ;
        RECT 78.200 48.000 78.600 49.900 ;
        RECT 79.800 48.000 80.200 49.900 ;
        RECT 78.200 47.900 80.200 48.000 ;
        RECT 80.600 47.900 81.000 49.900 ;
        RECT 81.700 48.200 82.100 49.900 ;
        RECT 81.700 47.900 82.600 48.200 ;
        RECT 72.700 47.400 74.600 47.700 ;
        RECT 70.700 47.100 71.100 47.200 ;
        RECT 65.800 46.800 71.300 47.100 ;
        RECT 55.000 46.400 55.400 46.500 ;
        RECT 53.500 46.100 55.400 46.400 ;
        RECT 55.900 46.200 56.200 46.800 ;
        RECT 59.500 46.700 59.900 46.800 ;
        RECT 59.000 46.200 59.400 46.300 ;
        RECT 60.300 46.200 60.700 46.300 ;
        RECT 63.200 46.200 63.500 46.800 ;
        RECT 67.300 46.700 67.700 46.800 ;
        RECT 53.500 46.000 53.900 46.100 ;
        RECT 55.800 45.800 56.200 46.200 ;
        RECT 58.200 45.900 60.700 46.200 ;
        RECT 58.200 45.800 58.600 45.900 ;
        RECT 63.000 45.800 63.500 46.200 ;
        RECT 63.800 45.800 64.200 46.600 ;
        RECT 66.500 46.200 66.900 46.300 ;
        RECT 71.000 46.200 71.300 46.800 ;
        RECT 71.800 46.400 72.200 46.500 ;
        RECT 66.500 46.100 69.000 46.200 ;
        RECT 69.400 46.100 69.800 46.200 ;
        RECT 66.500 45.900 69.800 46.100 ;
        RECT 68.600 45.800 69.800 45.900 ;
        RECT 71.000 45.800 71.400 46.200 ;
        RECT 71.800 46.100 73.700 46.400 ;
        RECT 73.300 46.000 73.700 46.100 ;
        RECT 54.300 45.700 54.700 45.800 ;
        RECT 52.600 45.400 54.700 45.700 ;
        RECT 52.600 41.100 53.000 45.400 ;
        RECT 55.900 45.200 56.200 45.800 ;
        RECT 59.000 45.500 61.800 45.600 ;
        RECT 58.900 45.400 61.800 45.500 ;
        RECT 55.000 44.900 56.200 45.200 ;
        RECT 56.900 45.300 61.800 45.400 ;
        RECT 56.900 45.100 59.300 45.300 ;
        RECT 55.000 44.400 55.300 44.900 ;
        RECT 54.600 44.000 55.300 44.400 ;
        RECT 56.100 44.500 56.500 44.600 ;
        RECT 56.900 44.500 57.200 45.100 ;
        RECT 56.100 44.200 57.200 44.500 ;
        RECT 57.500 44.500 60.200 44.800 ;
        RECT 57.500 44.400 57.900 44.500 ;
        RECT 59.800 44.400 60.200 44.500 ;
        RECT 56.700 43.700 57.100 43.800 ;
        RECT 58.100 43.700 58.500 43.800 ;
        RECT 55.000 43.100 55.400 43.500 ;
        RECT 56.700 43.400 58.500 43.700 ;
        RECT 57.100 43.100 57.400 43.400 ;
        RECT 59.800 43.100 60.200 43.500 ;
        RECT 54.700 41.100 55.300 43.100 ;
        RECT 57.000 41.100 57.400 43.100 ;
        RECT 59.200 42.800 60.200 43.100 ;
        RECT 59.200 41.100 59.600 42.800 ;
        RECT 61.400 41.100 61.800 45.300 ;
        RECT 62.200 45.100 62.600 45.200 ;
        RECT 63.200 45.100 63.500 45.800 ;
        RECT 65.400 45.500 68.200 45.600 ;
        RECT 65.400 45.400 68.300 45.500 ;
        RECT 65.400 45.300 70.300 45.400 ;
        RECT 62.200 44.800 62.900 45.100 ;
        RECT 63.200 44.800 63.700 45.100 ;
        RECT 62.600 44.200 62.900 44.800 ;
        RECT 62.600 43.800 63.000 44.200 ;
        RECT 63.300 41.100 63.700 44.800 ;
        RECT 65.400 41.100 65.800 45.300 ;
        RECT 67.900 45.100 70.300 45.300 ;
        RECT 67.000 44.500 69.700 44.800 ;
        RECT 67.000 44.400 67.400 44.500 ;
        RECT 69.300 44.400 69.700 44.500 ;
        RECT 70.000 44.500 70.300 45.100 ;
        RECT 71.000 45.200 71.300 45.800 ;
        RECT 72.500 45.700 72.900 45.800 ;
        RECT 74.200 45.700 74.600 47.400 ;
        RECT 75.100 47.200 75.400 47.900 ;
        RECT 75.900 47.700 77.700 47.900 ;
        RECT 78.300 47.700 80.100 47.900 ;
        RECT 77.000 47.200 77.400 47.400 ;
        RECT 78.600 47.200 79.000 47.400 ;
        RECT 80.600 47.200 80.900 47.900 ;
        RECT 75.000 46.800 76.300 47.200 ;
        RECT 77.000 47.100 77.800 47.200 ;
        RECT 78.200 47.100 79.000 47.200 ;
        RECT 77.000 46.900 79.000 47.100 ;
        RECT 77.400 46.800 78.600 46.900 ;
        RECT 79.700 46.800 81.000 47.200 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 76.000 46.100 76.300 46.800 ;
        RECT 75.000 45.800 76.300 46.100 ;
        RECT 76.600 45.800 77.000 46.600 ;
        RECT 79.000 45.800 79.400 46.600 ;
        RECT 72.500 45.400 74.600 45.700 ;
        RECT 71.000 44.900 72.200 45.200 ;
        RECT 70.700 44.500 71.100 44.600 ;
        RECT 70.000 44.200 71.100 44.500 ;
        RECT 71.900 44.400 72.200 44.900 ;
        RECT 71.900 44.000 72.600 44.400 ;
        RECT 68.700 43.700 69.100 43.800 ;
        RECT 70.100 43.700 70.500 43.800 ;
        RECT 67.000 43.100 67.400 43.500 ;
        RECT 68.700 43.400 70.500 43.700 ;
        RECT 69.800 43.100 70.100 43.400 ;
        RECT 71.800 43.100 72.200 43.500 ;
        RECT 67.000 42.800 68.000 43.100 ;
        RECT 67.600 41.100 68.000 42.800 ;
        RECT 69.800 41.100 70.200 43.100 ;
        RECT 71.900 41.100 72.500 43.100 ;
        RECT 74.200 41.100 74.600 45.400 ;
        RECT 75.000 45.100 75.400 45.200 ;
        RECT 76.000 45.100 76.300 45.800 ;
        RECT 79.700 45.100 80.000 46.800 ;
        RECT 82.200 46.100 82.600 47.900 ;
        RECT 83.800 47.700 84.200 49.900 ;
        RECT 85.900 49.200 86.500 49.900 ;
        RECT 85.900 48.900 86.600 49.200 ;
        RECT 88.200 48.900 88.600 49.900 ;
        RECT 90.400 49.200 90.800 49.900 ;
        RECT 90.400 48.900 91.400 49.200 ;
        RECT 86.200 48.500 86.600 48.900 ;
        RECT 88.300 48.600 88.600 48.900 ;
        RECT 88.300 48.300 89.700 48.600 ;
        RECT 89.300 48.200 89.700 48.300 ;
        RECT 90.200 48.200 90.600 48.600 ;
        RECT 91.000 48.500 91.400 48.900 ;
        RECT 85.300 47.700 85.700 47.800 ;
        RECT 83.000 47.100 83.400 47.600 ;
        RECT 83.800 47.400 85.700 47.700 ;
        RECT 83.800 47.100 84.200 47.400 ;
        RECT 90.200 47.200 90.500 48.200 ;
        RECT 92.600 47.500 93.000 49.900 ;
        RECT 95.000 48.000 95.400 49.900 ;
        RECT 96.600 48.000 97.000 49.900 ;
        RECT 95.000 47.900 97.000 48.000 ;
        RECT 97.400 47.900 97.800 49.900 ;
        RECT 98.500 48.200 98.900 49.900 ;
        RECT 98.500 47.900 99.400 48.200 ;
        RECT 95.100 47.700 96.900 47.900 ;
        RECT 95.400 47.200 95.800 47.400 ;
        RECT 97.400 47.200 97.700 47.900 ;
        RECT 87.300 47.100 87.700 47.200 ;
        RECT 90.200 47.100 90.600 47.200 ;
        RECT 91.800 47.100 92.600 47.200 ;
        RECT 94.200 47.100 94.600 47.200 ;
        RECT 83.000 46.800 84.200 47.100 ;
        RECT 80.600 45.800 82.600 46.100 ;
        RECT 80.600 45.200 80.900 45.800 ;
        RECT 80.600 45.100 81.000 45.200 ;
        RECT 75.000 44.800 75.700 45.100 ;
        RECT 76.000 44.800 76.500 45.100 ;
        RECT 75.400 44.200 75.700 44.800 ;
        RECT 75.400 43.800 75.800 44.200 ;
        RECT 76.100 41.100 76.500 44.800 ;
        RECT 79.500 44.800 80.000 45.100 ;
        RECT 80.300 44.800 81.000 45.100 ;
        RECT 79.500 41.100 79.900 44.800 ;
        RECT 80.300 44.200 80.600 44.800 ;
        RECT 81.400 44.400 81.800 45.200 ;
        RECT 80.200 43.800 80.600 44.200 ;
        RECT 82.200 41.100 82.600 45.800 ;
        RECT 83.800 45.700 84.200 46.800 ;
        RECT 87.100 46.800 94.600 47.100 ;
        RECT 95.000 46.900 95.800 47.200 ;
        RECT 96.500 47.100 97.800 47.200 ;
        RECT 98.200 47.100 98.600 47.200 ;
        RECT 95.000 46.800 95.400 46.900 ;
        RECT 96.500 46.800 98.600 47.100 ;
        RECT 86.200 46.400 86.600 46.500 ;
        RECT 84.700 46.100 86.600 46.400 ;
        RECT 84.700 46.000 85.100 46.100 ;
        RECT 85.500 45.700 85.900 45.800 ;
        RECT 83.800 45.400 85.900 45.700 ;
        RECT 83.800 41.100 84.200 45.400 ;
        RECT 87.100 45.200 87.400 46.800 ;
        RECT 90.700 46.700 91.100 46.800 ;
        RECT 91.500 46.200 91.900 46.300 ;
        RECT 87.800 46.100 88.200 46.200 ;
        RECT 89.400 46.100 91.900 46.200 ;
        RECT 87.800 45.900 91.900 46.100 ;
        RECT 87.800 45.800 89.800 45.900 ;
        RECT 95.800 45.800 96.200 46.600 ;
        RECT 90.200 45.500 93.000 45.600 ;
        RECT 90.100 45.400 93.000 45.500 ;
        RECT 86.200 44.900 87.400 45.200 ;
        RECT 88.100 45.300 93.000 45.400 ;
        RECT 88.100 45.100 90.500 45.300 ;
        RECT 86.200 44.400 86.500 44.900 ;
        RECT 85.800 44.000 86.500 44.400 ;
        RECT 87.300 44.500 87.700 44.600 ;
        RECT 88.100 44.500 88.400 45.100 ;
        RECT 87.300 44.200 88.400 44.500 ;
        RECT 88.700 44.500 91.400 44.800 ;
        RECT 88.700 44.400 89.100 44.500 ;
        RECT 91.000 44.400 91.400 44.500 ;
        RECT 87.900 43.700 88.300 43.800 ;
        RECT 89.300 43.700 89.700 43.800 ;
        RECT 86.200 43.100 86.600 43.500 ;
        RECT 87.900 43.400 89.700 43.700 ;
        RECT 88.300 43.100 88.600 43.400 ;
        RECT 91.000 43.100 91.400 43.500 ;
        RECT 85.900 41.100 86.500 43.100 ;
        RECT 88.200 41.100 88.600 43.100 ;
        RECT 90.400 42.800 91.400 43.100 ;
        RECT 90.400 41.100 90.800 42.800 ;
        RECT 92.600 41.100 93.000 45.300 ;
        RECT 96.500 45.100 96.800 46.800 ;
        RECT 99.000 46.100 99.400 47.900 ;
        RECT 99.800 46.800 100.200 47.600 ;
        RECT 100.600 47.500 101.000 49.900 ;
        RECT 102.800 49.200 103.200 49.900 ;
        RECT 102.200 48.900 103.200 49.200 ;
        RECT 105.000 48.900 105.400 49.900 ;
        RECT 107.100 49.200 107.700 49.900 ;
        RECT 107.000 48.900 107.700 49.200 ;
        RECT 102.200 48.500 102.600 48.900 ;
        RECT 105.000 48.600 105.300 48.900 ;
        RECT 103.000 48.200 103.400 48.600 ;
        RECT 103.900 48.300 105.300 48.600 ;
        RECT 107.000 48.500 107.400 48.900 ;
        RECT 103.900 48.200 104.300 48.300 ;
        RECT 101.000 47.100 101.800 47.200 ;
        RECT 103.100 47.100 103.400 48.200 ;
        RECT 107.900 47.700 108.300 47.800 ;
        RECT 109.400 47.700 109.800 49.900 ;
        RECT 110.200 47.800 110.600 48.600 ;
        RECT 107.900 47.400 109.800 47.700 ;
        RECT 105.900 47.100 106.300 47.200 ;
        RECT 101.000 46.800 106.500 47.100 ;
        RECT 102.500 46.700 102.900 46.800 ;
        RECT 97.400 45.800 99.400 46.100 ;
        RECT 101.700 46.200 102.100 46.300 ;
        RECT 103.000 46.200 103.400 46.300 ;
        RECT 101.700 45.900 104.200 46.200 ;
        RECT 103.800 45.800 104.200 45.900 ;
        RECT 97.400 45.200 97.700 45.800 ;
        RECT 97.400 45.100 97.800 45.200 ;
        RECT 96.300 44.800 96.800 45.100 ;
        RECT 97.100 44.800 97.800 45.100 ;
        RECT 96.300 41.100 96.700 44.800 ;
        RECT 97.100 44.200 97.400 44.800 ;
        RECT 98.200 44.400 98.600 45.200 ;
        RECT 97.000 43.800 97.400 44.200 ;
        RECT 99.000 41.100 99.400 45.800 ;
        RECT 100.600 45.500 103.400 45.600 ;
        RECT 100.600 45.400 103.500 45.500 ;
        RECT 100.600 45.300 105.500 45.400 ;
        RECT 100.600 41.100 101.000 45.300 ;
        RECT 103.100 45.100 105.500 45.300 ;
        RECT 102.200 44.500 104.900 44.800 ;
        RECT 102.200 44.400 102.600 44.500 ;
        RECT 104.500 44.400 104.900 44.500 ;
        RECT 105.200 44.500 105.500 45.100 ;
        RECT 106.200 45.200 106.500 46.800 ;
        RECT 107.000 46.400 107.400 46.500 ;
        RECT 107.000 46.100 108.900 46.400 ;
        RECT 108.500 46.000 108.900 46.100 ;
        RECT 107.700 45.700 108.100 45.800 ;
        RECT 109.400 45.700 109.800 47.400 ;
        RECT 107.700 45.400 109.800 45.700 ;
        RECT 106.200 44.900 107.400 45.200 ;
        RECT 105.900 44.500 106.300 44.600 ;
        RECT 105.200 44.200 106.300 44.500 ;
        RECT 107.100 44.400 107.400 44.900 ;
        RECT 107.100 44.000 107.800 44.400 ;
        RECT 103.900 43.700 104.300 43.800 ;
        RECT 105.300 43.700 105.700 43.800 ;
        RECT 102.200 43.100 102.600 43.500 ;
        RECT 103.900 43.400 105.700 43.700 ;
        RECT 105.000 43.100 105.300 43.400 ;
        RECT 107.000 43.100 107.400 43.500 ;
        RECT 102.200 42.800 103.200 43.100 ;
        RECT 102.800 41.100 103.200 42.800 ;
        RECT 105.000 41.100 105.400 43.100 ;
        RECT 107.100 41.100 107.700 43.100 ;
        RECT 109.400 41.100 109.800 45.400 ;
        RECT 111.000 41.100 111.400 49.900 ;
        RECT 113.700 48.000 114.100 49.500 ;
        RECT 115.800 48.500 116.200 49.500 ;
        RECT 113.300 47.700 114.100 48.000 ;
        RECT 113.300 47.500 113.700 47.700 ;
        RECT 113.300 47.200 113.600 47.500 ;
        RECT 115.900 47.400 116.200 48.500 ;
        RECT 112.600 46.800 113.600 47.200 ;
        RECT 114.100 47.100 116.200 47.400 ;
        RECT 116.600 48.500 117.000 49.500 ;
        RECT 116.600 47.400 116.900 48.500 ;
        RECT 118.700 48.000 119.100 49.500 ;
        RECT 121.700 49.200 122.100 49.900 ;
        RECT 124.100 49.200 124.500 49.900 ;
        RECT 121.700 48.800 122.600 49.200 ;
        RECT 123.800 48.800 124.500 49.200 ;
        RECT 121.700 48.200 122.100 48.800 ;
        RECT 124.100 48.200 124.500 48.800 ;
        RECT 118.700 47.700 119.500 48.000 ;
        RECT 121.700 47.900 122.600 48.200 ;
        RECT 124.100 47.900 125.000 48.200 ;
        RECT 119.100 47.500 119.500 47.700 ;
        RECT 116.600 47.100 118.700 47.400 ;
        RECT 114.100 46.900 114.600 47.100 ;
        RECT 112.600 45.400 113.000 46.200 ;
        RECT 113.300 44.900 113.600 46.800 ;
        RECT 113.900 46.500 114.600 46.900 ;
        RECT 118.200 46.900 118.700 47.100 ;
        RECT 119.200 47.200 119.500 47.500 ;
        RECT 114.300 45.500 114.600 46.500 ;
        RECT 115.000 45.800 115.400 46.600 ;
        RECT 115.800 45.800 116.200 46.600 ;
        RECT 116.600 45.800 117.000 46.600 ;
        RECT 117.400 45.800 117.800 46.600 ;
        RECT 118.200 46.500 118.900 46.900 ;
        RECT 119.200 46.800 120.200 47.200 ;
        RECT 118.200 45.500 118.500 46.500 ;
        RECT 114.300 45.200 116.200 45.500 ;
        RECT 113.300 44.600 114.100 44.900 ;
        RECT 113.700 43.200 114.100 44.600 ;
        RECT 115.900 43.500 116.200 45.200 ;
        RECT 113.700 42.800 114.600 43.200 ;
        RECT 113.700 41.100 114.100 42.800 ;
        RECT 115.800 41.500 116.200 43.500 ;
        RECT 116.600 45.200 118.500 45.500 ;
        RECT 116.600 43.500 116.900 45.200 ;
        RECT 119.200 44.900 119.500 46.800 ;
        RECT 119.800 46.100 120.200 46.200 ;
        RECT 120.600 46.100 121.000 46.200 ;
        RECT 119.800 45.800 121.000 46.100 ;
        RECT 119.800 45.400 120.200 45.800 ;
        RECT 118.700 44.600 119.500 44.900 ;
        RECT 116.600 41.500 117.000 43.500 ;
        RECT 118.700 41.100 119.100 44.600 ;
        RECT 121.400 44.400 121.800 45.200 ;
        RECT 122.200 41.100 122.600 47.900 ;
        RECT 123.000 46.800 123.400 47.600 ;
        RECT 123.000 45.100 123.400 45.200 ;
        RECT 123.800 45.100 124.200 45.200 ;
        RECT 123.000 44.800 124.200 45.100 ;
        RECT 123.800 44.400 124.200 44.800 ;
        RECT 124.600 41.100 125.000 47.900 ;
        RECT 126.200 47.700 126.600 49.900 ;
        RECT 128.300 49.200 128.900 49.900 ;
        RECT 128.300 48.900 129.000 49.200 ;
        RECT 130.600 48.900 131.000 49.900 ;
        RECT 132.800 49.200 133.200 49.900 ;
        RECT 132.800 48.900 133.800 49.200 ;
        RECT 128.600 48.500 129.000 48.900 ;
        RECT 130.700 48.600 131.000 48.900 ;
        RECT 130.700 48.300 132.100 48.600 ;
        RECT 131.700 48.200 132.100 48.300 ;
        RECT 132.600 48.200 133.000 48.600 ;
        RECT 133.400 48.500 133.800 48.900 ;
        RECT 127.700 47.700 128.100 47.800 ;
        RECT 125.400 46.800 125.800 47.600 ;
        RECT 126.200 47.400 128.100 47.700 ;
        RECT 126.200 45.700 126.600 47.400 ;
        RECT 129.700 47.100 130.100 47.200 ;
        RECT 132.600 47.100 132.900 48.200 ;
        RECT 135.000 47.500 135.400 49.900 ;
        RECT 137.100 48.200 137.500 49.900 ;
        RECT 136.600 47.900 137.500 48.200 ;
        RECT 138.200 47.900 138.600 49.900 ;
        RECT 139.000 48.000 139.400 49.900 ;
        RECT 140.600 48.000 141.000 49.900 ;
        RECT 139.000 47.900 141.000 48.000 ;
        RECT 134.200 47.100 135.000 47.200 ;
        RECT 129.500 46.800 135.000 47.100 ;
        RECT 135.800 46.800 136.200 47.600 ;
        RECT 128.600 46.400 129.000 46.500 ;
        RECT 127.100 46.100 129.000 46.400 ;
        RECT 127.100 46.000 127.500 46.100 ;
        RECT 127.900 45.700 128.300 45.800 ;
        RECT 126.200 45.400 128.300 45.700 ;
        RECT 126.200 41.100 126.600 45.400 ;
        RECT 129.500 45.200 129.800 46.800 ;
        RECT 133.100 46.700 133.500 46.800 ;
        RECT 133.900 46.200 134.300 46.300 ;
        RECT 131.800 45.900 134.300 46.200 ;
        RECT 136.600 46.100 137.000 47.900 ;
        RECT 138.300 47.200 138.600 47.900 ;
        RECT 139.100 47.700 140.900 47.900 ;
        RECT 140.200 47.200 140.600 47.400 ;
        RECT 138.200 46.800 139.500 47.200 ;
        RECT 140.200 46.900 141.000 47.200 ;
        RECT 140.600 46.800 141.000 46.900 ;
        RECT 143.000 46.800 143.400 47.600 ;
        RECT 131.800 45.800 132.200 45.900 ;
        RECT 136.600 45.800 138.500 46.100 ;
        RECT 132.600 45.500 135.400 45.600 ;
        RECT 132.500 45.400 135.400 45.500 ;
        RECT 128.600 44.900 129.800 45.200 ;
        RECT 130.500 45.300 135.400 45.400 ;
        RECT 130.500 45.100 132.900 45.300 ;
        RECT 128.600 44.400 128.900 44.900 ;
        RECT 128.200 44.000 128.900 44.400 ;
        RECT 129.700 44.500 130.100 44.600 ;
        RECT 130.500 44.500 130.800 45.100 ;
        RECT 129.700 44.200 130.800 44.500 ;
        RECT 131.100 44.500 133.800 44.800 ;
        RECT 131.100 44.400 131.500 44.500 ;
        RECT 133.400 44.400 133.800 44.500 ;
        RECT 130.300 43.700 130.700 43.800 ;
        RECT 131.700 43.700 132.100 43.800 ;
        RECT 128.600 43.100 129.000 43.500 ;
        RECT 130.300 43.400 132.100 43.700 ;
        RECT 130.700 43.100 131.000 43.400 ;
        RECT 133.400 43.100 133.800 43.500 ;
        RECT 128.300 41.100 128.900 43.100 ;
        RECT 130.600 41.100 131.000 43.100 ;
        RECT 132.800 42.800 133.800 43.100 ;
        RECT 132.800 41.100 133.200 42.800 ;
        RECT 135.000 41.100 135.400 45.300 ;
        RECT 136.600 41.100 137.000 45.800 ;
        RECT 138.200 45.200 138.500 45.800 ;
        RECT 137.400 44.400 137.800 45.200 ;
        RECT 138.200 45.100 138.600 45.200 ;
        RECT 139.200 45.100 139.500 46.800 ;
        RECT 139.800 45.800 140.200 46.600 ;
        RECT 138.200 44.800 138.900 45.100 ;
        RECT 139.200 44.800 139.700 45.100 ;
        RECT 138.600 44.200 138.900 44.800 ;
        RECT 138.600 43.800 139.000 44.200 ;
        RECT 139.300 41.100 139.700 44.800 ;
        RECT 143.800 41.100 144.200 49.900 ;
        RECT 145.700 49.200 146.100 49.900 ;
        RECT 145.700 48.800 146.600 49.200 ;
        RECT 145.700 48.200 146.100 48.800 ;
        RECT 145.700 47.900 146.600 48.200 ;
        RECT 147.800 48.000 148.200 49.900 ;
        RECT 149.400 48.000 149.800 49.900 ;
        RECT 147.800 47.900 149.800 48.000 ;
        RECT 150.200 47.900 150.600 49.900 ;
        RECT 145.400 44.400 145.800 45.200 ;
        RECT 146.200 41.100 146.600 47.900 ;
        RECT 147.900 47.700 149.700 47.900 ;
        RECT 147.000 46.800 147.400 47.600 ;
        RECT 148.200 47.200 148.600 47.400 ;
        RECT 150.200 47.200 150.500 47.900 ;
        RECT 151.000 47.500 151.400 49.900 ;
        RECT 153.200 49.200 153.600 49.900 ;
        RECT 152.600 48.900 153.600 49.200 ;
        RECT 155.400 48.900 155.800 49.900 ;
        RECT 157.500 49.200 158.100 49.900 ;
        RECT 157.400 48.900 158.100 49.200 ;
        RECT 152.600 48.500 153.000 48.900 ;
        RECT 155.400 48.600 155.700 48.900 ;
        RECT 153.400 48.200 153.800 48.600 ;
        RECT 154.300 48.300 155.700 48.600 ;
        RECT 157.400 48.500 157.800 48.900 ;
        RECT 154.300 48.200 154.700 48.300 ;
        RECT 147.800 46.900 148.600 47.200 ;
        RECT 147.800 46.800 148.200 46.900 ;
        RECT 149.300 46.800 150.600 47.200 ;
        RECT 151.400 47.100 152.200 47.200 ;
        RECT 153.500 47.100 153.800 48.200 ;
        RECT 158.300 47.700 158.700 47.800 ;
        RECT 159.800 47.700 160.200 49.900 ;
        RECT 158.300 47.400 160.200 47.700 ;
        RECT 154.200 47.100 154.600 47.200 ;
        RECT 156.300 47.100 156.700 47.200 ;
        RECT 151.400 46.800 156.900 47.100 ;
        RECT 148.600 45.800 149.000 46.600 ;
        RECT 149.300 46.200 149.600 46.800 ;
        RECT 152.900 46.700 153.300 46.800 ;
        RECT 152.100 46.200 152.500 46.300 ;
        RECT 153.400 46.200 153.800 46.300 ;
        RECT 149.300 45.800 149.800 46.200 ;
        RECT 152.100 45.900 154.600 46.200 ;
        RECT 154.200 45.800 154.600 45.900 ;
        RECT 149.300 45.100 149.600 45.800 ;
        RECT 151.000 45.500 153.800 45.600 ;
        RECT 151.000 45.400 153.900 45.500 ;
        RECT 151.000 45.300 155.900 45.400 ;
        RECT 150.200 45.100 150.600 45.200 ;
        RECT 149.100 44.800 149.600 45.100 ;
        RECT 149.900 44.800 150.600 45.100 ;
        RECT 149.100 41.100 149.500 44.800 ;
        RECT 149.900 44.200 150.200 44.800 ;
        RECT 149.800 43.800 150.200 44.200 ;
        RECT 151.000 41.100 151.400 45.300 ;
        RECT 153.500 45.100 155.900 45.300 ;
        RECT 152.600 44.500 155.300 44.800 ;
        RECT 152.600 44.400 153.000 44.500 ;
        RECT 154.900 44.400 155.300 44.500 ;
        RECT 155.600 44.500 155.900 45.100 ;
        RECT 156.600 45.200 156.900 46.800 ;
        RECT 157.400 46.400 157.800 46.500 ;
        RECT 157.400 46.100 159.300 46.400 ;
        RECT 158.900 46.000 159.300 46.100 ;
        RECT 158.100 45.700 158.500 45.800 ;
        RECT 159.800 45.700 160.200 47.400 ;
        RECT 160.600 47.600 161.000 49.900 ;
        RECT 163.000 48.000 163.400 49.900 ;
        RECT 164.600 48.000 165.000 49.900 ;
        RECT 163.000 47.900 165.000 48.000 ;
        RECT 165.400 47.900 165.800 49.900 ;
        RECT 166.500 48.200 166.900 49.900 ;
        RECT 166.500 47.900 167.400 48.200 ;
        RECT 163.100 47.700 164.900 47.900 ;
        RECT 160.600 47.300 161.700 47.600 ;
        RECT 160.600 45.800 161.000 46.600 ;
        RECT 161.400 45.800 161.700 47.300 ;
        RECT 163.400 47.200 163.800 47.400 ;
        RECT 165.400 47.200 165.700 47.900 ;
        RECT 163.000 46.900 163.800 47.200 ;
        RECT 164.500 47.100 165.800 47.200 ;
        RECT 166.200 47.100 166.600 47.200 ;
        RECT 163.000 46.800 163.400 46.900 ;
        RECT 164.500 46.800 166.600 47.100 ;
        RECT 163.800 45.800 164.200 46.600 ;
        RECT 158.100 45.400 160.200 45.700 ;
        RECT 156.600 44.900 157.800 45.200 ;
        RECT 156.300 44.500 156.700 44.600 ;
        RECT 155.600 44.200 156.700 44.500 ;
        RECT 157.500 44.400 157.800 44.900 ;
        RECT 157.500 44.000 158.200 44.400 ;
        RECT 154.300 43.700 154.700 43.800 ;
        RECT 155.700 43.700 156.100 43.800 ;
        RECT 152.600 43.100 153.000 43.500 ;
        RECT 154.300 43.400 156.100 43.700 ;
        RECT 155.400 43.100 155.700 43.400 ;
        RECT 157.400 43.100 157.800 43.500 ;
        RECT 152.600 42.800 153.600 43.100 ;
        RECT 153.200 41.100 153.600 42.800 ;
        RECT 155.400 41.100 155.800 43.100 ;
        RECT 157.500 41.100 158.100 43.100 ;
        RECT 159.800 41.100 160.200 45.400 ;
        RECT 161.400 45.400 162.000 45.800 ;
        RECT 161.400 45.100 161.700 45.400 ;
        RECT 164.500 45.100 164.800 46.800 ;
        RECT 167.000 46.100 167.400 47.900 ;
        RECT 168.600 47.700 169.000 49.900 ;
        RECT 170.700 49.200 171.300 49.900 ;
        RECT 170.700 48.900 171.400 49.200 ;
        RECT 173.000 48.900 173.400 49.900 ;
        RECT 175.200 49.200 175.600 49.900 ;
        RECT 175.200 48.900 176.200 49.200 ;
        RECT 171.000 48.500 171.400 48.900 ;
        RECT 173.100 48.600 173.400 48.900 ;
        RECT 173.100 48.300 174.500 48.600 ;
        RECT 174.100 48.200 174.500 48.300 ;
        RECT 175.000 48.200 175.400 48.600 ;
        RECT 175.800 48.500 176.200 48.900 ;
        RECT 170.200 47.800 170.600 48.200 ;
        RECT 170.100 47.700 170.600 47.800 ;
        RECT 167.800 47.100 168.200 47.600 ;
        RECT 168.600 47.400 170.600 47.700 ;
        RECT 168.600 47.100 169.000 47.400 ;
        RECT 172.100 47.100 172.500 47.200 ;
        RECT 175.000 47.100 175.300 48.200 ;
        RECT 177.400 47.500 177.800 49.900 ;
        RECT 179.000 48.200 179.400 49.900 ;
        RECT 178.900 47.900 179.400 48.200 ;
        RECT 178.900 47.200 179.200 47.900 ;
        RECT 180.600 47.600 181.000 49.900 ;
        RECT 179.700 47.300 181.000 47.600 ;
        RECT 181.400 48.500 181.800 49.500 ;
        RECT 183.500 49.200 183.900 49.500 ;
        RECT 183.000 48.800 183.900 49.200 ;
        RECT 181.400 47.400 181.700 48.500 ;
        RECT 183.500 48.000 183.900 48.800 ;
        RECT 183.500 47.700 184.300 48.000 ;
        RECT 183.900 47.500 184.300 47.700 ;
        RECT 176.600 47.100 177.400 47.200 ;
        RECT 167.800 46.800 169.000 47.100 ;
        RECT 165.400 45.800 167.400 46.100 ;
        RECT 165.400 45.200 165.700 45.800 ;
        RECT 165.400 45.100 165.800 45.200 ;
        RECT 160.600 44.800 161.700 45.100 ;
        RECT 164.300 44.800 164.800 45.100 ;
        RECT 165.100 44.800 165.800 45.100 ;
        RECT 160.600 41.100 161.000 44.800 ;
        RECT 164.300 41.100 164.700 44.800 ;
        RECT 165.100 44.200 165.400 44.800 ;
        RECT 166.200 44.400 166.600 45.200 ;
        RECT 165.000 43.800 165.400 44.200 ;
        RECT 167.000 41.100 167.400 45.800 ;
        RECT 168.600 45.700 169.000 46.800 ;
        RECT 171.900 46.800 177.400 47.100 ;
        RECT 178.900 46.800 179.400 47.200 ;
        RECT 171.000 46.400 171.400 46.500 ;
        RECT 169.500 46.100 171.400 46.400 ;
        RECT 171.900 46.100 172.200 46.800 ;
        RECT 175.500 46.700 175.900 46.800 ;
        RECT 176.300 46.200 176.700 46.300 ;
        RECT 172.600 46.100 173.000 46.200 ;
        RECT 169.500 46.000 169.900 46.100 ;
        RECT 171.800 45.800 173.000 46.100 ;
        RECT 174.200 45.900 176.700 46.200 ;
        RECT 174.200 45.800 174.600 45.900 ;
        RECT 170.300 45.700 170.700 45.800 ;
        RECT 168.600 45.400 170.700 45.700 ;
        RECT 168.600 41.100 169.000 45.400 ;
        RECT 171.900 45.200 172.200 45.800 ;
        RECT 175.000 45.500 177.800 45.600 ;
        RECT 174.900 45.400 177.800 45.500 ;
        RECT 171.000 44.900 172.200 45.200 ;
        RECT 172.900 45.300 177.800 45.400 ;
        RECT 172.900 45.100 175.300 45.300 ;
        RECT 171.000 44.400 171.300 44.900 ;
        RECT 170.600 44.000 171.300 44.400 ;
        RECT 172.100 44.500 172.500 44.600 ;
        RECT 172.900 44.500 173.200 45.100 ;
        RECT 172.100 44.200 173.200 44.500 ;
        RECT 173.500 44.500 176.200 44.800 ;
        RECT 173.500 44.400 173.900 44.500 ;
        RECT 175.800 44.400 176.200 44.500 ;
        RECT 172.700 43.700 173.100 43.800 ;
        RECT 174.100 43.700 174.500 43.800 ;
        RECT 171.000 43.100 171.400 43.500 ;
        RECT 172.700 43.400 174.500 43.700 ;
        RECT 173.100 43.100 173.400 43.400 ;
        RECT 175.800 43.100 176.200 43.500 ;
        RECT 170.700 41.100 171.300 43.100 ;
        RECT 173.000 41.100 173.400 43.100 ;
        RECT 175.200 42.800 176.200 43.100 ;
        RECT 175.200 41.100 175.600 42.800 ;
        RECT 177.400 41.100 177.800 45.300 ;
        RECT 178.900 45.100 179.200 46.800 ;
        RECT 179.700 46.500 180.000 47.300 ;
        RECT 181.400 47.100 183.500 47.400 ;
        RECT 183.000 46.900 183.500 47.100 ;
        RECT 184.000 47.200 184.300 47.500 ;
        RECT 186.200 47.700 186.600 49.900 ;
        RECT 188.300 49.200 188.900 49.900 ;
        RECT 188.300 48.900 189.000 49.200 ;
        RECT 190.600 48.900 191.000 49.900 ;
        RECT 192.800 49.200 193.200 49.900 ;
        RECT 192.800 48.900 193.800 49.200 ;
        RECT 188.600 48.500 189.000 48.900 ;
        RECT 190.700 48.600 191.000 48.900 ;
        RECT 190.700 48.300 192.100 48.600 ;
        RECT 191.700 48.200 192.100 48.300 ;
        RECT 192.600 48.200 193.000 48.600 ;
        RECT 193.400 48.500 193.800 48.900 ;
        RECT 187.700 47.700 188.100 47.800 ;
        RECT 186.200 47.400 188.100 47.700 ;
        RECT 179.500 46.100 180.000 46.500 ;
        RECT 179.700 45.100 180.000 46.100 ;
        RECT 180.500 46.200 180.900 46.600 ;
        RECT 180.500 45.800 181.000 46.200 ;
        RECT 181.400 45.800 181.800 46.600 ;
        RECT 182.200 45.800 182.600 46.600 ;
        RECT 183.000 46.500 183.700 46.900 ;
        RECT 184.000 46.800 185.000 47.200 ;
        RECT 183.000 45.500 183.300 46.500 ;
        RECT 181.400 45.200 183.300 45.500 ;
        RECT 178.900 44.600 179.400 45.100 ;
        RECT 179.700 44.800 181.000 45.100 ;
        RECT 179.000 41.100 179.400 44.600 ;
        RECT 180.600 41.100 181.000 44.800 ;
        RECT 181.400 43.500 181.700 45.200 ;
        RECT 184.000 44.900 184.300 46.800 ;
        RECT 184.600 45.400 185.000 46.200 ;
        RECT 186.200 45.700 186.600 47.400 ;
        RECT 189.700 47.100 190.100 47.200 ;
        RECT 191.800 47.100 192.200 47.200 ;
        RECT 192.600 47.100 192.900 48.200 ;
        RECT 195.000 47.500 195.400 49.900 ;
        RECT 197.400 47.600 197.800 49.900 ;
        RECT 199.000 48.200 199.400 49.900 ;
        RECT 201.400 48.200 201.800 49.900 ;
        RECT 199.000 47.900 199.500 48.200 ;
        RECT 197.400 47.300 198.700 47.600 ;
        RECT 194.200 47.100 195.000 47.200 ;
        RECT 189.500 46.800 195.000 47.100 ;
        RECT 188.600 46.400 189.000 46.500 ;
        RECT 187.100 46.100 189.000 46.400 ;
        RECT 187.100 46.000 187.500 46.100 ;
        RECT 187.900 45.700 188.300 45.800 ;
        RECT 186.200 45.400 188.300 45.700 ;
        RECT 183.500 44.600 184.300 44.900 ;
        RECT 181.400 41.500 181.800 43.500 ;
        RECT 183.500 41.100 183.900 44.600 ;
        RECT 186.200 41.100 186.600 45.400 ;
        RECT 189.500 45.200 189.800 46.800 ;
        RECT 193.100 46.700 193.500 46.800 ;
        RECT 192.600 46.200 193.000 46.300 ;
        RECT 193.900 46.200 194.300 46.300 ;
        RECT 197.500 46.200 197.900 46.600 ;
        RECT 191.800 45.900 194.300 46.200 ;
        RECT 196.600 46.100 197.000 46.200 ;
        RECT 197.400 46.100 197.900 46.200 ;
        RECT 191.800 45.800 192.200 45.900 ;
        RECT 196.600 45.800 197.900 46.100 ;
        RECT 198.400 46.500 198.700 47.300 ;
        RECT 199.200 47.200 199.500 47.900 ;
        RECT 199.000 46.800 199.500 47.200 ;
        RECT 198.400 46.100 198.900 46.500 ;
        RECT 192.600 45.500 195.400 45.600 ;
        RECT 192.500 45.400 195.400 45.500 ;
        RECT 188.600 44.900 189.800 45.200 ;
        RECT 190.500 45.300 195.400 45.400 ;
        RECT 190.500 45.100 192.900 45.300 ;
        RECT 188.600 44.400 188.900 44.900 ;
        RECT 188.200 44.000 188.900 44.400 ;
        RECT 189.700 44.500 190.100 44.600 ;
        RECT 190.500 44.500 190.800 45.100 ;
        RECT 189.700 44.200 190.800 44.500 ;
        RECT 191.100 44.500 193.800 44.800 ;
        RECT 191.100 44.400 191.500 44.500 ;
        RECT 193.400 44.400 193.800 44.500 ;
        RECT 190.300 43.700 190.700 43.800 ;
        RECT 191.700 43.700 192.100 43.800 ;
        RECT 188.600 43.100 189.000 43.500 ;
        RECT 190.300 43.400 192.100 43.700 ;
        RECT 190.700 43.100 191.000 43.400 ;
        RECT 193.400 43.100 193.800 43.500 ;
        RECT 188.300 41.100 188.900 43.100 ;
        RECT 190.600 41.100 191.000 43.100 ;
        RECT 192.800 42.800 193.800 43.100 ;
        RECT 192.800 41.100 193.200 42.800 ;
        RECT 195.000 41.100 195.400 45.300 ;
        RECT 198.400 45.100 198.700 46.100 ;
        RECT 199.200 45.100 199.500 46.800 ;
        RECT 197.400 44.800 198.700 45.100 ;
        RECT 197.400 41.100 197.800 44.800 ;
        RECT 199.000 44.600 199.500 45.100 ;
        RECT 201.300 47.900 201.800 48.200 ;
        RECT 201.300 47.200 201.600 47.900 ;
        RECT 203.000 47.600 203.400 49.900 ;
        RECT 205.700 48.000 206.100 49.500 ;
        RECT 207.800 48.500 208.200 49.500 ;
        RECT 202.100 47.300 203.400 47.600 ;
        RECT 205.300 47.700 206.100 48.000 ;
        RECT 205.300 47.500 205.700 47.700 ;
        RECT 201.300 46.800 201.800 47.200 ;
        RECT 201.300 45.100 201.600 46.800 ;
        RECT 202.100 46.500 202.400 47.300 ;
        RECT 205.300 47.200 205.600 47.500 ;
        RECT 207.900 47.400 208.200 48.500 ;
        RECT 209.900 48.200 210.300 49.900 ;
        RECT 209.400 47.900 210.300 48.200 ;
        RECT 211.000 47.900 211.400 49.900 ;
        RECT 211.800 48.000 212.200 49.900 ;
        RECT 213.400 48.000 213.800 49.900 ;
        RECT 215.500 49.200 215.900 49.900 ;
        RECT 215.500 48.800 216.200 49.200 ;
        RECT 215.500 48.200 215.900 48.800 ;
        RECT 211.800 47.900 213.800 48.000 ;
        RECT 215.000 47.900 215.900 48.200 ;
        RECT 216.600 48.000 217.000 49.900 ;
        RECT 218.200 48.000 218.600 49.900 ;
        RECT 216.600 47.900 218.600 48.000 ;
        RECT 219.000 47.900 219.400 49.900 ;
        RECT 204.600 46.800 205.600 47.200 ;
        RECT 206.100 47.100 208.200 47.400 ;
        RECT 206.100 46.900 206.600 47.100 ;
        RECT 201.900 46.100 202.400 46.500 ;
        RECT 202.100 45.100 202.400 46.100 ;
        RECT 202.900 46.200 203.300 46.600 ;
        RECT 202.900 45.800 203.400 46.200 ;
        RECT 204.600 45.400 205.000 46.200 ;
        RECT 201.300 44.600 201.800 45.100 ;
        RECT 202.100 44.800 203.400 45.100 ;
        RECT 199.000 41.100 199.400 44.600 ;
        RECT 201.400 41.100 201.800 44.600 ;
        RECT 203.000 41.100 203.400 44.800 ;
        RECT 205.300 44.900 205.600 46.800 ;
        RECT 205.900 46.500 206.600 46.900 ;
        RECT 208.600 46.800 209.000 47.600 ;
        RECT 206.300 45.500 206.600 46.500 ;
        RECT 207.000 45.800 207.400 46.600 ;
        RECT 207.800 45.800 208.200 46.600 ;
        RECT 209.400 46.100 209.800 47.900 ;
        RECT 211.100 47.200 211.400 47.900 ;
        RECT 211.900 47.700 213.700 47.900 ;
        RECT 213.000 47.200 213.400 47.400 ;
        RECT 211.000 46.800 212.300 47.200 ;
        RECT 213.000 46.900 213.800 47.200 ;
        RECT 213.400 46.800 213.800 46.900 ;
        RECT 214.200 46.800 214.600 47.600 ;
        RECT 212.000 46.200 212.300 46.800 ;
        RECT 209.400 45.800 211.300 46.100 ;
        RECT 211.800 45.800 212.300 46.200 ;
        RECT 212.600 45.800 213.000 46.600 ;
        RECT 206.300 45.200 208.200 45.500 ;
        RECT 205.300 44.600 206.100 44.900 ;
        RECT 205.700 41.100 206.100 44.600 ;
        RECT 207.900 43.500 208.200 45.200 ;
        RECT 207.800 41.500 208.200 43.500 ;
        RECT 209.400 41.100 209.800 45.800 ;
        RECT 211.000 45.200 211.300 45.800 ;
        RECT 210.200 44.400 210.600 45.200 ;
        RECT 211.000 45.100 211.400 45.200 ;
        RECT 212.000 45.100 212.300 45.800 ;
        RECT 211.000 44.800 211.700 45.100 ;
        RECT 212.000 44.800 212.500 45.100 ;
        RECT 211.400 44.200 211.700 44.800 ;
        RECT 211.400 43.800 211.800 44.200 ;
        RECT 212.100 41.100 212.500 44.800 ;
        RECT 215.000 41.100 215.400 47.900 ;
        RECT 216.700 47.700 218.500 47.900 ;
        RECT 217.000 47.200 217.400 47.400 ;
        RECT 219.000 47.200 219.300 47.900 ;
        RECT 219.800 47.700 220.200 49.900 ;
        RECT 221.900 49.200 222.500 49.900 ;
        RECT 221.900 48.900 222.600 49.200 ;
        RECT 224.200 48.900 224.600 49.900 ;
        RECT 226.400 49.200 226.800 49.900 ;
        RECT 226.400 48.900 227.400 49.200 ;
        RECT 222.200 48.500 222.600 48.900 ;
        RECT 224.300 48.600 224.600 48.900 ;
        RECT 224.300 48.300 225.700 48.600 ;
        RECT 225.300 48.200 225.700 48.300 ;
        RECT 226.200 48.200 226.600 48.600 ;
        RECT 227.000 48.500 227.400 48.900 ;
        RECT 221.300 47.700 221.700 47.800 ;
        RECT 219.800 47.400 221.700 47.700 ;
        RECT 216.600 46.900 217.400 47.200 ;
        RECT 216.600 46.800 217.000 46.900 ;
        RECT 218.100 46.800 219.400 47.200 ;
        RECT 217.400 45.800 217.800 46.600 ;
        RECT 218.100 46.100 218.400 46.800 ;
        RECT 219.000 46.100 219.400 46.200 ;
        RECT 218.100 45.800 219.400 46.100 ;
        RECT 215.800 44.400 216.200 45.200 ;
        RECT 218.100 45.100 218.400 45.800 ;
        RECT 219.800 45.700 220.200 47.400 ;
        RECT 220.600 46.800 221.000 47.400 ;
        RECT 223.300 47.100 223.700 47.200 ;
        RECT 225.400 47.100 225.800 47.200 ;
        RECT 226.200 47.100 226.500 48.200 ;
        RECT 228.600 47.500 229.000 49.900 ;
        RECT 227.800 47.100 228.600 47.200 ;
        RECT 223.100 46.800 228.600 47.100 ;
        RECT 222.200 46.400 222.600 46.500 ;
        RECT 220.700 46.100 222.600 46.400 ;
        RECT 220.700 46.000 221.100 46.100 ;
        RECT 221.500 45.700 221.900 45.800 ;
        RECT 219.800 45.400 221.900 45.700 ;
        RECT 219.000 45.100 219.400 45.200 ;
        RECT 217.900 44.800 218.400 45.100 ;
        RECT 218.700 44.800 219.400 45.100 ;
        RECT 217.900 41.100 218.300 44.800 ;
        RECT 218.700 44.200 219.000 44.800 ;
        RECT 218.600 43.800 219.000 44.200 ;
        RECT 219.800 41.100 220.200 45.400 ;
        RECT 223.100 45.200 223.400 46.800 ;
        RECT 226.700 46.700 227.100 46.800 ;
        RECT 227.500 46.200 227.900 46.300 ;
        RECT 224.600 46.100 225.000 46.200 ;
        RECT 225.400 46.100 227.900 46.200 ;
        RECT 224.600 45.900 227.900 46.100 ;
        RECT 224.600 45.800 225.800 45.900 ;
        RECT 226.200 45.500 229.000 45.600 ;
        RECT 226.100 45.400 229.000 45.500 ;
        RECT 222.200 44.900 223.400 45.200 ;
        RECT 224.100 45.300 229.000 45.400 ;
        RECT 224.100 45.100 226.500 45.300 ;
        RECT 222.200 44.400 222.500 44.900 ;
        RECT 221.800 44.000 222.500 44.400 ;
        RECT 223.300 44.500 223.700 44.600 ;
        RECT 224.100 44.500 224.400 45.100 ;
        RECT 223.300 44.200 224.400 44.500 ;
        RECT 224.700 44.500 227.400 44.800 ;
        RECT 224.700 44.400 225.100 44.500 ;
        RECT 227.000 44.400 227.400 44.500 ;
        RECT 223.900 43.700 224.300 43.800 ;
        RECT 225.300 43.700 225.700 43.800 ;
        RECT 222.200 43.100 222.600 43.500 ;
        RECT 223.900 43.400 225.700 43.700 ;
        RECT 224.300 43.100 224.600 43.400 ;
        RECT 227.000 43.100 227.400 43.500 ;
        RECT 221.900 41.100 222.500 43.100 ;
        RECT 224.200 41.100 224.600 43.100 ;
        RECT 226.400 42.800 227.400 43.100 ;
        RECT 226.400 41.100 226.800 42.800 ;
        RECT 228.600 41.100 229.000 45.300 ;
        RECT 0.600 35.800 1.000 36.600 ;
        RECT 1.400 33.100 1.800 39.900 ;
        RECT 2.200 34.100 2.600 34.200 ;
        RECT 2.200 33.800 3.300 34.100 ;
        RECT 2.200 33.400 2.600 33.800 ;
        RECT 0.900 32.800 1.800 33.100 ;
        RECT 3.000 33.200 3.300 33.800 ;
        RECT 0.900 32.200 1.300 32.800 ;
        RECT 3.000 32.400 3.400 33.200 ;
        RECT 0.600 31.800 1.300 32.200 ;
        RECT 0.900 31.100 1.300 31.800 ;
        RECT 3.800 31.100 4.200 39.900 ;
        RECT 5.900 36.200 6.300 39.900 ;
        RECT 6.600 36.800 7.000 37.200 ;
        RECT 6.700 36.200 7.000 36.800 ;
        RECT 5.900 35.900 6.400 36.200 ;
        RECT 6.700 35.900 7.400 36.200 ;
        RECT 5.400 34.400 5.800 35.200 ;
        RECT 6.100 34.200 6.400 35.900 ;
        RECT 7.000 35.800 7.400 35.900 ;
        RECT 7.800 35.800 8.200 36.600 ;
        RECT 7.000 35.100 7.300 35.800 ;
        RECT 8.600 35.100 9.000 39.900 ;
        RECT 7.000 34.800 9.000 35.100 ;
        RECT 4.600 34.100 5.000 34.200 ;
        RECT 4.600 33.800 5.400 34.100 ;
        RECT 6.100 33.800 7.400 34.200 ;
        RECT 5.000 33.600 5.400 33.800 ;
        RECT 4.700 33.100 6.500 33.300 ;
        RECT 7.000 33.100 7.300 33.800 ;
        RECT 8.600 33.100 9.000 34.800 ;
        RECT 9.400 34.100 9.800 34.200 ;
        RECT 11.000 34.100 11.400 39.900 ;
        RECT 13.100 39.200 14.100 39.900 ;
        RECT 13.100 38.800 14.600 39.200 ;
        RECT 13.100 35.900 14.100 38.800 ;
        RECT 11.800 34.100 12.200 34.600 ;
        RECT 12.600 34.400 13.000 35.200 ;
        RECT 13.500 34.200 13.800 35.900 ;
        RECT 15.800 35.700 16.200 39.900 ;
        RECT 18.000 38.200 18.400 39.900 ;
        RECT 17.400 37.900 18.400 38.200 ;
        RECT 20.200 37.900 20.600 39.900 ;
        RECT 22.300 37.900 22.900 39.900 ;
        RECT 17.400 37.500 17.800 37.900 ;
        RECT 20.200 37.600 20.500 37.900 ;
        RECT 19.100 37.300 20.900 37.600 ;
        RECT 22.200 37.500 22.600 37.900 ;
        RECT 19.100 37.200 19.500 37.300 ;
        RECT 20.500 37.200 20.900 37.300 ;
        RECT 17.400 36.500 17.800 36.600 ;
        RECT 19.700 36.500 20.100 36.600 ;
        RECT 17.400 36.200 20.100 36.500 ;
        RECT 20.400 36.500 21.500 36.800 ;
        RECT 20.400 35.900 20.700 36.500 ;
        RECT 21.100 36.400 21.500 36.500 ;
        RECT 22.300 36.600 23.000 37.000 ;
        RECT 22.300 36.100 22.600 36.600 ;
        RECT 18.300 35.700 20.700 35.900 ;
        RECT 15.800 35.600 20.700 35.700 ;
        RECT 21.400 35.800 22.600 36.100 ;
        RECT 15.800 35.500 18.700 35.600 ;
        RECT 15.800 35.400 18.600 35.500 ;
        RECT 21.400 35.200 21.700 35.800 ;
        RECT 24.600 35.600 25.000 39.900 ;
        RECT 22.900 35.300 25.000 35.600 ;
        RECT 22.900 35.200 23.300 35.300 ;
        RECT 14.200 34.400 14.600 35.200 ;
        RECT 19.000 35.100 19.400 35.200 ;
        RECT 16.900 34.800 19.400 35.100 ;
        RECT 21.400 34.800 21.800 35.200 ;
        RECT 23.700 34.900 24.100 35.000 ;
        RECT 16.900 34.700 17.300 34.800 ;
        RECT 17.700 34.200 18.100 34.300 ;
        RECT 21.400 34.200 21.700 34.800 ;
        RECT 22.200 34.600 24.100 34.900 ;
        RECT 22.200 34.500 22.600 34.600 ;
        RECT 13.400 34.100 13.800 34.200 ;
        RECT 15.000 34.100 15.400 34.200 ;
        RECT 9.400 33.800 10.500 34.100 ;
        RECT 9.400 33.400 9.800 33.800 ;
        RECT 4.600 33.000 6.600 33.100 ;
        RECT 4.600 31.100 5.000 33.000 ;
        RECT 6.200 31.100 6.600 33.000 ;
        RECT 7.000 31.100 7.400 33.100 ;
        RECT 8.100 32.800 9.000 33.100 ;
        RECT 10.200 33.200 10.500 33.800 ;
        RECT 11.000 33.800 12.200 34.100 ;
        RECT 12.600 33.800 13.800 34.100 ;
        RECT 14.600 33.800 15.400 34.100 ;
        RECT 16.200 33.900 21.700 34.200 ;
        RECT 16.200 33.800 17.000 33.900 ;
        RECT 8.100 31.100 8.500 32.800 ;
        RECT 10.200 32.400 10.600 33.200 ;
        RECT 11.000 31.100 11.400 33.800 ;
        RECT 12.600 33.100 12.900 33.800 ;
        RECT 14.600 33.600 15.000 33.800 ;
        RECT 13.500 33.100 15.300 33.300 ;
        RECT 11.800 31.400 12.200 33.100 ;
        RECT 12.600 31.700 13.000 33.100 ;
        RECT 13.400 33.000 15.400 33.100 ;
        RECT 13.400 31.400 13.800 33.000 ;
        RECT 11.800 31.100 13.800 31.400 ;
        RECT 15.000 31.100 15.400 33.000 ;
        RECT 15.800 31.100 16.200 33.500 ;
        RECT 18.300 32.800 18.600 33.900 ;
        RECT 21.100 33.800 21.500 33.900 ;
        RECT 24.600 33.600 25.000 35.300 ;
        RECT 23.100 33.300 25.000 33.600 ;
        RECT 23.100 33.200 23.500 33.300 ;
        RECT 24.600 33.100 25.000 33.300 ;
        RECT 25.400 33.100 25.800 33.200 ;
        RECT 24.600 32.800 25.800 33.100 ;
        RECT 17.400 32.100 17.800 32.500 ;
        RECT 18.200 32.400 18.600 32.800 ;
        RECT 19.100 32.700 19.500 32.800 ;
        RECT 19.100 32.400 20.500 32.700 ;
        RECT 20.200 32.100 20.500 32.400 ;
        RECT 22.200 32.100 22.600 32.500 ;
        RECT 17.400 31.800 18.400 32.100 ;
        RECT 18.000 31.100 18.400 31.800 ;
        RECT 20.200 31.100 20.600 32.100 ;
        RECT 22.200 31.800 22.900 32.100 ;
        RECT 22.300 31.100 22.900 31.800 ;
        RECT 24.600 31.100 25.000 32.800 ;
        RECT 25.400 32.400 25.800 32.800 ;
        RECT 26.200 31.100 26.600 39.900 ;
        RECT 28.300 39.200 29.300 39.900 ;
        RECT 28.300 38.800 29.800 39.200 ;
        RECT 28.300 35.900 29.300 38.800 ;
        RECT 27.000 33.800 27.400 34.600 ;
        RECT 27.800 34.400 28.200 35.200 ;
        RECT 28.700 34.200 29.000 35.900 ;
        RECT 29.400 35.100 29.800 35.200 ;
        RECT 31.000 35.100 31.400 39.900 ;
        RECT 32.600 35.700 33.000 39.900 ;
        RECT 34.800 38.200 35.200 39.900 ;
        RECT 34.200 37.900 35.200 38.200 ;
        RECT 37.000 37.900 37.400 39.900 ;
        RECT 39.100 37.900 39.700 39.900 ;
        RECT 34.200 37.500 34.600 37.900 ;
        RECT 37.000 37.600 37.300 37.900 ;
        RECT 35.900 37.300 37.700 37.600 ;
        RECT 39.000 37.500 39.400 37.900 ;
        RECT 35.900 37.200 36.300 37.300 ;
        RECT 37.300 37.200 37.700 37.300 ;
        RECT 39.500 37.000 40.200 37.200 ;
        RECT 39.100 36.800 40.200 37.000 ;
        RECT 34.200 36.500 34.600 36.600 ;
        RECT 36.500 36.500 36.900 36.600 ;
        RECT 34.200 36.200 36.900 36.500 ;
        RECT 37.200 36.500 38.300 36.800 ;
        RECT 37.200 35.900 37.500 36.500 ;
        RECT 37.900 36.400 38.300 36.500 ;
        RECT 39.100 36.600 39.800 36.800 ;
        RECT 39.100 36.100 39.400 36.600 ;
        RECT 35.100 35.700 37.500 35.900 ;
        RECT 32.600 35.600 37.500 35.700 ;
        RECT 38.200 35.800 39.400 36.100 ;
        RECT 32.600 35.500 35.500 35.600 ;
        RECT 32.600 35.400 35.400 35.500 ;
        RECT 35.800 35.100 36.200 35.200 ;
        RECT 37.400 35.100 37.800 35.200 ;
        RECT 29.400 34.800 31.400 35.100 ;
        RECT 29.400 34.400 29.800 34.800 ;
        RECT 28.600 34.100 29.000 34.200 ;
        RECT 30.200 34.100 30.600 34.200 ;
        RECT 27.800 33.800 29.000 34.100 ;
        RECT 29.800 33.800 30.600 34.100 ;
        RECT 27.800 33.100 28.100 33.800 ;
        RECT 29.800 33.600 30.200 33.800 ;
        RECT 28.700 33.100 30.500 33.300 ;
        RECT 27.000 31.400 27.400 33.100 ;
        RECT 27.800 31.700 28.200 33.100 ;
        RECT 28.600 33.000 30.600 33.100 ;
        RECT 28.600 31.400 29.000 33.000 ;
        RECT 27.000 31.100 29.000 31.400 ;
        RECT 30.200 31.100 30.600 33.000 ;
        RECT 31.000 31.100 31.400 34.800 ;
        RECT 33.700 34.800 37.800 35.100 ;
        RECT 33.700 34.700 34.100 34.800 ;
        RECT 34.500 34.200 34.900 34.300 ;
        RECT 38.200 34.200 38.500 35.800 ;
        RECT 41.400 35.600 41.800 39.900 ;
        RECT 43.000 39.100 43.400 39.200 ;
        RECT 43.800 39.100 44.200 39.900 ;
        RECT 43.000 38.800 44.200 39.100 ;
        RECT 39.700 35.300 41.800 35.600 ;
        RECT 39.700 35.200 40.100 35.300 ;
        RECT 40.500 34.900 40.900 35.000 ;
        RECT 39.000 34.600 40.900 34.900 ;
        RECT 39.000 34.500 39.400 34.600 ;
        RECT 33.000 33.900 38.500 34.200 ;
        RECT 33.000 33.800 33.800 33.900 ;
        RECT 31.800 32.400 32.200 33.200 ;
        RECT 32.600 31.100 33.000 33.500 ;
        RECT 35.100 32.800 35.400 33.900 ;
        RECT 37.900 33.800 38.300 33.900 ;
        RECT 41.400 33.600 41.800 35.300 ;
        RECT 39.900 33.300 41.800 33.600 ;
        RECT 39.900 33.200 40.300 33.300 ;
        RECT 34.200 32.100 34.600 32.500 ;
        RECT 35.000 32.400 35.400 32.800 ;
        RECT 35.900 32.700 36.300 32.800 ;
        RECT 35.900 32.400 37.300 32.700 ;
        RECT 37.000 32.100 37.300 32.400 ;
        RECT 39.000 32.100 39.400 32.500 ;
        RECT 34.200 31.800 35.200 32.100 ;
        RECT 34.800 31.100 35.200 31.800 ;
        RECT 37.000 31.100 37.400 32.100 ;
        RECT 39.000 31.800 39.700 32.100 ;
        RECT 39.100 31.100 39.700 31.800 ;
        RECT 41.400 31.100 41.800 33.300 ;
        RECT 43.800 31.100 44.200 38.800 ;
        RECT 46.200 35.100 46.600 39.900 ;
        RECT 48.200 36.800 48.600 37.200 ;
        RECT 47.000 35.800 47.400 36.600 ;
        RECT 48.200 36.200 48.500 36.800 ;
        RECT 48.900 36.200 49.300 39.900 ;
        RECT 47.800 35.900 48.500 36.200 ;
        RECT 48.800 35.900 49.300 36.200 ;
        RECT 51.000 36.200 51.400 39.900 ;
        RECT 52.600 36.400 53.000 39.900 ;
        RECT 56.100 39.200 56.500 39.900 ;
        RECT 56.100 38.800 57.000 39.200 ;
        RECT 56.100 36.400 56.500 38.800 ;
        RECT 58.200 37.500 58.600 39.500 ;
        RECT 51.000 35.900 52.300 36.200 ;
        RECT 52.600 35.900 53.100 36.400 ;
        RECT 47.800 35.800 48.200 35.900 ;
        RECT 47.800 35.100 48.100 35.800 ;
        RECT 46.200 34.800 48.100 35.100 ;
        RECT 44.600 34.100 45.000 34.200 ;
        RECT 45.400 34.100 45.800 34.200 ;
        RECT 44.600 33.800 45.800 34.100 ;
        RECT 44.600 33.200 44.900 33.800 ;
        RECT 45.400 33.400 45.800 33.800 ;
        RECT 44.600 32.400 45.000 33.200 ;
        RECT 46.200 33.100 46.600 34.800 ;
        RECT 48.800 34.200 49.100 35.900 ;
        RECT 49.400 34.400 49.800 35.200 ;
        RECT 51.000 34.800 51.500 35.200 ;
        RECT 51.100 34.400 51.500 34.800 ;
        RECT 52.000 34.900 52.300 35.900 ;
        RECT 52.000 34.500 52.500 34.900 ;
        RECT 47.800 33.800 49.100 34.200 ;
        RECT 50.200 34.100 50.600 34.200 ;
        RECT 49.800 33.800 50.600 34.100 ;
        RECT 47.900 33.100 48.200 33.800 ;
        RECT 49.800 33.600 50.200 33.800 ;
        RECT 52.000 33.700 52.300 34.500 ;
        RECT 52.800 34.200 53.100 35.900 ;
        RECT 55.700 36.100 56.500 36.400 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 55.000 35.100 55.400 35.600 ;
        RECT 54.200 34.800 55.400 35.100 ;
        RECT 55.700 34.200 56.000 36.100 ;
        RECT 58.300 35.800 58.600 37.500 ;
        RECT 56.700 35.500 58.600 35.800 ;
        RECT 56.700 34.500 57.000 35.500 ;
        RECT 52.600 33.800 53.100 34.200 ;
        RECT 55.000 33.800 56.000 34.200 ;
        RECT 56.300 34.100 57.000 34.500 ;
        RECT 57.400 34.400 57.800 35.200 ;
        RECT 58.200 34.400 58.600 35.200 ;
        RECT 51.000 33.400 52.300 33.700 ;
        RECT 48.700 33.100 50.500 33.300 ;
        RECT 46.200 32.800 47.100 33.100 ;
        RECT 46.700 31.100 47.100 32.800 ;
        RECT 47.800 31.100 48.200 33.100 ;
        RECT 48.600 33.000 50.600 33.100 ;
        RECT 48.600 31.100 49.000 33.000 ;
        RECT 50.200 31.100 50.600 33.000 ;
        RECT 51.000 31.100 51.400 33.400 ;
        RECT 52.800 33.100 53.100 33.800 ;
        RECT 52.600 32.800 53.100 33.100 ;
        RECT 55.700 33.500 56.000 33.800 ;
        RECT 56.500 33.900 57.000 34.100 ;
        RECT 56.500 33.600 58.600 33.900 ;
        RECT 55.700 33.300 56.100 33.500 ;
        RECT 55.700 33.000 56.500 33.300 ;
        RECT 52.600 31.100 53.000 32.800 ;
        RECT 56.100 31.500 56.500 33.000 ;
        RECT 58.300 32.500 58.600 33.600 ;
        RECT 59.000 33.400 59.400 34.200 ;
        RECT 59.800 33.100 60.200 39.900 ;
        RECT 60.600 35.800 61.000 36.600 ;
        RECT 62.700 36.200 63.100 39.900 ;
        RECT 63.400 36.800 63.800 37.200 ;
        RECT 63.500 36.200 63.800 36.800 ;
        RECT 62.700 35.900 63.200 36.200 ;
        RECT 63.500 35.900 64.200 36.200 ;
        RECT 62.200 34.400 62.600 35.200 ;
        RECT 62.900 34.200 63.200 35.900 ;
        RECT 63.800 35.800 64.200 35.900 ;
        RECT 64.600 35.800 65.000 36.600 ;
        RECT 63.800 35.100 64.100 35.800 ;
        RECT 65.400 35.100 65.800 39.900 ;
        RECT 68.900 39.200 69.300 39.900 ;
        RECT 68.900 38.800 69.800 39.200 ;
        RECT 68.900 36.400 69.300 38.800 ;
        RECT 71.000 37.500 71.400 39.500 ;
        RECT 73.100 39.200 73.500 39.900 ;
        RECT 72.600 38.800 73.500 39.200 ;
        RECT 68.500 36.100 69.300 36.400 ;
        RECT 67.800 35.100 68.200 35.600 ;
        RECT 63.800 34.800 65.800 35.100 ;
        RECT 61.400 34.100 61.800 34.200 ;
        RECT 61.400 33.800 62.200 34.100 ;
        RECT 62.900 33.800 64.200 34.200 ;
        RECT 61.800 33.600 62.200 33.800 ;
        RECT 61.500 33.100 63.300 33.300 ;
        RECT 63.800 33.100 64.100 33.800 ;
        RECT 65.400 33.100 65.800 34.800 ;
        RECT 67.000 34.800 68.200 35.100 ;
        RECT 66.200 34.100 66.600 34.200 ;
        RECT 67.000 34.100 67.300 34.800 ;
        RECT 68.500 34.200 68.800 36.100 ;
        RECT 71.100 35.800 71.400 37.500 ;
        RECT 73.100 36.200 73.500 38.800 ;
        RECT 73.800 36.800 74.200 37.200 ;
        RECT 73.900 36.200 74.200 36.800 ;
        RECT 73.100 35.900 73.600 36.200 ;
        RECT 73.900 36.100 74.600 36.200 ;
        RECT 75.800 36.100 76.200 39.900 ;
        RECT 73.900 35.900 76.200 36.100 ;
        RECT 69.500 35.500 71.400 35.800 ;
        RECT 69.500 34.500 69.800 35.500 ;
        RECT 66.200 33.800 67.300 34.100 ;
        RECT 67.800 33.800 68.800 34.200 ;
        RECT 69.100 34.100 69.800 34.500 ;
        RECT 70.200 34.400 70.600 35.200 ;
        RECT 71.000 34.400 71.400 35.200 ;
        RECT 72.600 34.400 73.000 35.200 ;
        RECT 73.300 34.200 73.600 35.900 ;
        RECT 74.200 35.800 76.200 35.900 ;
        RECT 76.600 35.800 77.000 37.200 ;
        RECT 78.700 36.200 79.100 39.900 ;
        RECT 79.400 36.800 79.800 37.200 ;
        RECT 79.500 36.200 79.800 36.800 ;
        RECT 78.700 35.900 79.200 36.200 ;
        RECT 79.500 35.900 80.200 36.200 ;
        RECT 66.200 33.400 66.600 33.800 ;
        RECT 68.500 33.500 68.800 33.800 ;
        RECT 69.300 33.900 69.800 34.100 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 69.300 33.600 71.400 33.900 ;
        RECT 71.800 33.800 72.600 34.100 ;
        RECT 73.300 33.800 74.600 34.200 ;
        RECT 72.200 33.600 72.600 33.800 ;
        RECT 59.800 32.800 60.700 33.100 ;
        RECT 58.200 31.500 58.600 32.500 ;
        RECT 60.300 31.100 60.700 32.800 ;
        RECT 61.400 33.000 63.400 33.100 ;
        RECT 61.400 31.100 61.800 33.000 ;
        RECT 63.000 31.100 63.400 33.000 ;
        RECT 63.800 31.100 64.200 33.100 ;
        RECT 64.900 32.800 65.800 33.100 ;
        RECT 68.500 33.300 68.900 33.500 ;
        RECT 68.500 33.000 69.300 33.300 ;
        RECT 64.900 31.100 65.300 32.800 ;
        RECT 68.900 31.500 69.300 33.000 ;
        RECT 71.100 32.500 71.400 33.600 ;
        RECT 71.900 33.100 73.700 33.300 ;
        RECT 74.200 33.100 74.500 33.800 ;
        RECT 75.000 33.400 75.400 34.200 ;
        RECT 75.800 33.100 76.200 35.800 ;
        RECT 78.200 34.400 78.600 35.200 ;
        RECT 78.900 34.200 79.200 35.900 ;
        RECT 79.800 35.800 80.200 35.900 ;
        RECT 80.600 35.800 81.000 36.600 ;
        RECT 79.800 35.100 80.100 35.800 ;
        RECT 81.400 35.100 81.800 39.900 ;
        RECT 84.900 39.200 85.300 39.900 ;
        RECT 84.900 38.800 85.800 39.200 ;
        RECT 84.900 36.400 85.300 38.800 ;
        RECT 87.000 37.500 87.400 39.500 ;
        RECT 84.500 36.100 85.300 36.400 ;
        RECT 79.800 34.800 81.800 35.100 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 83.800 35.100 84.200 35.600 ;
        RECT 83.000 34.800 84.200 35.100 ;
        RECT 77.400 34.100 77.800 34.200 ;
        RECT 77.400 33.800 78.200 34.100 ;
        RECT 78.900 33.800 80.200 34.200 ;
        RECT 77.800 33.600 78.200 33.800 ;
        RECT 77.500 33.100 79.300 33.300 ;
        RECT 79.800 33.100 80.100 33.800 ;
        RECT 81.400 33.100 81.800 34.800 ;
        RECT 84.500 34.200 84.800 36.100 ;
        RECT 87.100 35.800 87.400 37.500 ;
        RECT 85.500 35.500 87.400 35.800 ;
        RECT 89.400 35.600 89.800 39.900 ;
        RECT 91.500 37.900 92.100 39.900 ;
        RECT 93.800 37.900 94.200 39.900 ;
        RECT 96.000 38.200 96.400 39.900 ;
        RECT 96.000 37.900 97.000 38.200 ;
        RECT 91.800 37.500 92.200 37.900 ;
        RECT 93.900 37.600 94.200 37.900 ;
        RECT 93.500 37.300 95.300 37.600 ;
        RECT 96.600 37.500 97.000 37.900 ;
        RECT 93.500 37.200 93.900 37.300 ;
        RECT 94.900 37.200 95.300 37.300 ;
        RECT 91.400 36.600 92.100 37.000 ;
        RECT 91.800 36.100 92.100 36.600 ;
        RECT 92.900 36.500 94.000 36.800 ;
        RECT 92.900 36.400 93.300 36.500 ;
        RECT 91.800 35.800 93.000 36.100 ;
        RECT 85.500 34.500 85.800 35.500 ;
        RECT 89.400 35.300 91.500 35.600 ;
        RECT 82.200 33.400 82.600 34.200 ;
        RECT 83.800 33.800 84.800 34.200 ;
        RECT 85.100 34.100 85.800 34.500 ;
        RECT 86.200 34.400 86.600 35.200 ;
        RECT 87.000 34.400 87.400 35.200 ;
        RECT 84.500 33.500 84.800 33.800 ;
        RECT 85.300 33.900 85.800 34.100 ;
        RECT 85.300 33.600 87.400 33.900 ;
        RECT 71.000 31.500 71.400 32.500 ;
        RECT 71.800 33.000 73.800 33.100 ;
        RECT 71.800 31.100 72.200 33.000 ;
        RECT 73.400 31.100 73.800 33.000 ;
        RECT 74.200 31.100 74.600 33.100 ;
        RECT 75.800 32.800 76.700 33.100 ;
        RECT 76.300 31.100 76.700 32.800 ;
        RECT 77.400 33.000 79.400 33.100 ;
        RECT 77.400 31.100 77.800 33.000 ;
        RECT 79.000 31.100 79.400 33.000 ;
        RECT 79.800 31.100 80.200 33.100 ;
        RECT 80.900 32.800 81.800 33.100 ;
        RECT 84.500 33.300 84.900 33.500 ;
        RECT 84.500 33.000 85.300 33.300 ;
        RECT 80.900 31.100 81.300 32.800 ;
        RECT 84.900 31.500 85.300 33.000 ;
        RECT 87.100 32.500 87.400 33.600 ;
        RECT 87.000 31.500 87.400 32.500 ;
        RECT 89.400 33.600 89.800 35.300 ;
        RECT 91.100 35.200 91.500 35.300 ;
        RECT 90.300 34.900 90.700 35.000 ;
        RECT 90.300 34.600 92.200 34.900 ;
        RECT 91.800 34.500 92.200 34.600 ;
        RECT 92.700 34.200 93.000 35.800 ;
        RECT 93.700 35.900 94.000 36.500 ;
        RECT 94.300 36.500 94.700 36.600 ;
        RECT 96.600 36.500 97.000 36.600 ;
        RECT 94.300 36.200 97.000 36.500 ;
        RECT 93.700 35.700 96.100 35.900 ;
        RECT 98.200 35.700 98.600 39.900 ;
        RECT 93.700 35.600 98.600 35.700 ;
        RECT 95.700 35.500 98.600 35.600 ;
        RECT 95.800 35.400 98.600 35.500 ;
        RECT 95.000 35.100 95.400 35.200 ;
        RECT 99.800 35.100 100.200 39.900 ;
        RECT 102.500 37.200 102.900 39.900 ;
        RECT 101.800 36.800 102.200 37.200 ;
        RECT 102.500 36.800 103.400 37.200 ;
        RECT 100.600 35.800 101.000 36.600 ;
        RECT 101.800 36.200 102.100 36.800 ;
        RECT 102.500 36.200 102.900 36.800 ;
        RECT 101.400 35.900 102.100 36.200 ;
        RECT 102.400 35.900 102.900 36.200 ;
        RECT 101.400 35.800 101.800 35.900 ;
        RECT 101.400 35.100 101.700 35.800 ;
        RECT 95.000 34.800 97.500 35.100 ;
        RECT 95.800 34.700 96.200 34.800 ;
        RECT 97.100 34.700 97.500 34.800 ;
        RECT 99.800 34.800 101.700 35.100 ;
        RECT 96.300 34.200 96.700 34.300 ;
        RECT 92.700 33.900 98.200 34.200 ;
        RECT 92.900 33.800 93.300 33.900 ;
        RECT 89.400 33.300 91.300 33.600 ;
        RECT 89.400 31.100 89.800 33.300 ;
        RECT 90.900 33.200 91.300 33.300 ;
        RECT 95.800 32.800 96.100 33.900 ;
        RECT 97.400 33.800 98.200 33.900 ;
        RECT 94.900 32.700 95.300 32.800 ;
        RECT 91.800 32.100 92.200 32.500 ;
        RECT 93.900 32.400 95.300 32.700 ;
        RECT 95.800 32.400 96.200 32.800 ;
        RECT 93.900 32.100 94.200 32.400 ;
        RECT 96.600 32.100 97.000 32.500 ;
        RECT 91.500 31.800 92.200 32.100 ;
        RECT 91.500 31.100 92.100 31.800 ;
        RECT 93.800 31.100 94.200 32.100 ;
        RECT 96.000 31.800 97.000 32.100 ;
        RECT 96.000 31.100 96.400 31.800 ;
        RECT 98.200 31.100 98.600 33.500 ;
        RECT 99.000 33.400 99.400 34.200 ;
        RECT 99.800 33.100 100.200 34.800 ;
        RECT 102.400 34.200 102.700 35.900 ;
        RECT 104.600 35.800 105.000 36.600 ;
        RECT 103.000 35.100 103.400 35.200 ;
        RECT 103.800 35.100 104.200 35.200 ;
        RECT 103.000 34.800 104.200 35.100 ;
        RECT 103.000 34.400 103.400 34.800 ;
        RECT 101.400 33.800 102.700 34.200 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 103.400 33.800 104.200 34.100 ;
        RECT 101.500 33.100 101.800 33.800 ;
        RECT 103.400 33.600 103.800 33.800 ;
        RECT 102.300 33.100 104.100 33.300 ;
        RECT 105.400 33.100 105.800 39.900 ;
        RECT 107.000 37.500 107.400 39.500 ;
        RECT 109.100 39.200 109.500 39.900 ;
        RECT 109.100 38.800 109.800 39.200 ;
        RECT 107.000 35.800 107.300 37.500 ;
        RECT 109.100 36.400 109.500 38.800 ;
        RECT 109.100 36.100 109.900 36.400 ;
        RECT 107.000 35.500 108.900 35.800 ;
        RECT 107.000 34.400 107.400 35.200 ;
        RECT 107.800 34.400 108.200 35.200 ;
        RECT 108.600 34.500 108.900 35.500 ;
        RECT 106.200 33.400 106.600 34.200 ;
        RECT 108.600 34.100 109.300 34.500 ;
        RECT 109.600 34.200 109.900 36.100 ;
        RECT 110.200 34.800 110.600 35.600 ;
        RECT 112.600 35.100 113.000 39.900 ;
        RECT 114.600 36.800 115.000 37.200 ;
        RECT 113.400 35.800 113.800 36.600 ;
        RECT 114.600 36.200 114.900 36.800 ;
        RECT 115.300 36.200 115.700 39.900 ;
        RECT 118.700 39.200 119.100 39.900 ;
        RECT 118.200 38.800 119.100 39.200 ;
        RECT 114.200 35.900 114.900 36.200 ;
        RECT 115.200 35.900 115.700 36.200 ;
        RECT 118.700 36.200 119.100 38.800 ;
        RECT 122.500 39.200 122.900 39.900 ;
        RECT 122.500 38.800 123.400 39.200 ;
        RECT 119.400 36.800 119.800 37.200 ;
        RECT 119.500 36.200 119.800 36.800 ;
        RECT 122.500 36.400 122.900 38.800 ;
        RECT 124.600 37.500 125.000 39.500 ;
        RECT 118.700 35.900 119.200 36.200 ;
        RECT 119.500 35.900 120.200 36.200 ;
        RECT 114.200 35.800 114.600 35.900 ;
        RECT 114.200 35.100 114.500 35.800 ;
        RECT 112.600 34.800 114.500 35.100 ;
        RECT 108.600 33.900 109.100 34.100 ;
        RECT 107.000 33.600 109.100 33.900 ;
        RECT 109.600 33.800 110.600 34.200 ;
        RECT 111.000 34.100 111.400 34.200 ;
        RECT 111.800 34.100 112.200 34.200 ;
        RECT 111.000 33.800 112.200 34.100 ;
        RECT 99.800 32.800 100.700 33.100 ;
        RECT 100.300 31.100 100.700 32.800 ;
        RECT 101.400 31.100 101.800 33.100 ;
        RECT 102.200 33.000 104.200 33.100 ;
        RECT 102.200 31.100 102.600 33.000 ;
        RECT 103.800 31.100 104.200 33.000 ;
        RECT 104.900 32.800 105.800 33.100 ;
        RECT 104.900 32.200 105.300 32.800 ;
        RECT 107.000 32.500 107.300 33.600 ;
        RECT 109.600 33.500 109.900 33.800 ;
        RECT 109.500 33.300 109.900 33.500 ;
        RECT 111.800 33.400 112.200 33.800 ;
        RECT 109.100 33.000 109.900 33.300 ;
        RECT 112.600 33.100 113.000 34.800 ;
        RECT 115.200 34.200 115.500 35.900 ;
        RECT 115.800 34.400 116.200 35.200 ;
        RECT 118.200 34.400 118.600 35.200 ;
        RECT 118.900 34.200 119.200 35.900 ;
        RECT 119.800 35.800 120.200 35.900 ;
        RECT 122.100 36.100 122.900 36.400 ;
        RECT 119.800 35.100 120.200 35.200 ;
        RECT 121.400 35.100 121.800 35.600 ;
        RECT 119.800 34.800 121.800 35.100 ;
        RECT 122.100 34.200 122.400 36.100 ;
        RECT 124.700 35.800 125.000 37.500 ;
        RECT 123.100 35.500 125.000 35.800 ;
        RECT 125.400 37.500 125.800 39.500 ;
        RECT 125.400 35.800 125.700 37.500 ;
        RECT 127.500 36.400 127.900 39.900 ;
        RECT 130.200 37.500 130.600 39.500 ;
        RECT 132.300 39.200 132.700 39.900 ;
        RECT 132.300 38.800 133.000 39.200 ;
        RECT 127.500 36.100 128.300 36.400 ;
        RECT 125.400 35.500 127.300 35.800 ;
        RECT 123.100 34.500 123.400 35.500 ;
        RECT 114.200 33.800 115.500 34.200 ;
        RECT 116.600 34.100 117.000 34.200 ;
        RECT 116.200 33.800 117.000 34.100 ;
        RECT 117.400 34.100 117.800 34.200 ;
        RECT 117.400 33.800 118.200 34.100 ;
        RECT 118.900 33.800 120.200 34.200 ;
        RECT 121.400 33.800 122.400 34.200 ;
        RECT 122.700 34.100 123.400 34.500 ;
        RECT 123.800 34.400 124.200 35.200 ;
        RECT 124.600 34.400 125.000 35.200 ;
        RECT 125.400 34.400 125.800 35.200 ;
        RECT 126.200 34.400 126.600 35.200 ;
        RECT 127.000 34.500 127.300 35.500 ;
        RECT 114.300 33.100 114.600 33.800 ;
        RECT 116.200 33.600 116.600 33.800 ;
        RECT 117.800 33.600 118.200 33.800 ;
        RECT 115.100 33.100 116.900 33.300 ;
        RECT 117.500 33.100 119.300 33.300 ;
        RECT 119.800 33.100 120.100 33.800 ;
        RECT 122.100 33.500 122.400 33.800 ;
        RECT 122.900 33.900 123.400 34.100 ;
        RECT 127.000 34.100 127.700 34.500 ;
        RECT 128.000 34.200 128.300 36.100 ;
        RECT 130.200 35.800 130.500 37.500 ;
        RECT 132.300 36.400 132.700 38.800 ;
        RECT 132.300 36.100 133.100 36.400 ;
        RECT 128.600 35.100 129.000 35.600 ;
        RECT 130.200 35.500 132.100 35.800 ;
        RECT 129.400 35.100 129.800 35.200 ;
        RECT 128.600 34.800 129.800 35.100 ;
        RECT 130.200 34.400 130.600 35.200 ;
        RECT 131.000 34.400 131.400 35.200 ;
        RECT 131.800 34.500 132.100 35.500 ;
        RECT 127.000 33.900 127.500 34.100 ;
        RECT 122.900 33.600 125.000 33.900 ;
        RECT 122.100 33.300 122.500 33.500 ;
        RECT 104.900 31.800 105.800 32.200 ;
        RECT 104.900 31.100 105.300 31.800 ;
        RECT 107.000 31.500 107.400 32.500 ;
        RECT 109.100 31.500 109.500 33.000 ;
        RECT 112.600 32.800 113.500 33.100 ;
        RECT 113.100 31.100 113.500 32.800 ;
        RECT 114.200 31.100 114.600 33.100 ;
        RECT 115.000 33.000 117.000 33.100 ;
        RECT 115.000 31.100 115.400 33.000 ;
        RECT 116.600 31.100 117.000 33.000 ;
        RECT 117.400 33.000 119.400 33.100 ;
        RECT 117.400 31.100 117.800 33.000 ;
        RECT 119.000 31.100 119.400 33.000 ;
        RECT 119.800 31.100 120.200 33.100 ;
        RECT 122.100 33.000 122.900 33.300 ;
        RECT 122.500 31.500 122.900 33.000 ;
        RECT 124.700 32.500 125.000 33.600 ;
        RECT 124.600 31.500 125.000 32.500 ;
        RECT 125.400 33.600 127.500 33.900 ;
        RECT 128.000 33.800 129.000 34.200 ;
        RECT 131.800 34.100 132.500 34.500 ;
        RECT 132.800 34.200 133.100 36.100 ;
        RECT 133.400 34.800 133.800 35.600 ;
        RECT 135.800 35.100 136.200 39.900 ;
        RECT 137.800 36.800 138.200 37.200 ;
        RECT 136.600 35.800 137.000 36.600 ;
        RECT 137.800 36.200 138.100 36.800 ;
        RECT 138.500 36.200 138.900 39.900 ;
        RECT 137.400 35.900 138.100 36.200 ;
        RECT 137.400 35.800 137.800 35.900 ;
        RECT 138.400 35.800 139.400 36.200 ;
        RECT 137.400 35.100 137.700 35.800 ;
        RECT 135.800 34.800 137.700 35.100 ;
        RECT 131.800 33.900 132.300 34.100 ;
        RECT 125.400 32.500 125.700 33.600 ;
        RECT 128.000 33.500 128.300 33.800 ;
        RECT 127.900 33.300 128.300 33.500 ;
        RECT 127.500 33.000 128.300 33.300 ;
        RECT 130.200 33.600 132.300 33.900 ;
        RECT 132.800 33.800 133.800 34.200 ;
        RECT 125.400 31.500 125.800 32.500 ;
        RECT 127.500 31.500 127.900 33.000 ;
        RECT 130.200 32.500 130.500 33.600 ;
        RECT 132.800 33.500 133.100 33.800 ;
        RECT 132.700 33.300 133.100 33.500 ;
        RECT 135.000 33.400 135.400 34.200 ;
        RECT 132.300 33.000 133.100 33.300 ;
        RECT 135.800 33.100 136.200 34.800 ;
        RECT 138.400 34.200 138.700 35.800 ;
        RECT 142.200 35.600 142.600 39.900 ;
        RECT 144.300 37.900 144.900 39.900 ;
        RECT 146.600 37.900 147.000 39.900 ;
        RECT 148.800 38.200 149.200 39.900 ;
        RECT 148.800 37.900 149.800 38.200 ;
        RECT 144.600 37.500 145.000 37.900 ;
        RECT 146.700 37.600 147.000 37.900 ;
        RECT 146.300 37.300 148.100 37.600 ;
        RECT 149.400 37.500 149.800 37.900 ;
        RECT 146.300 37.200 146.700 37.300 ;
        RECT 147.700 37.200 148.100 37.300 ;
        RECT 144.200 36.600 144.900 37.000 ;
        RECT 144.600 36.100 144.900 36.600 ;
        RECT 145.700 36.500 146.800 36.800 ;
        RECT 145.700 36.400 146.100 36.500 ;
        RECT 144.600 35.800 145.800 36.100 ;
        RECT 142.200 35.300 144.300 35.600 ;
        RECT 139.000 34.400 139.400 35.200 ;
        RECT 137.400 33.800 138.700 34.200 ;
        RECT 139.800 34.100 140.200 34.200 ;
        RECT 139.400 33.800 140.200 34.100 ;
        RECT 137.500 33.100 137.800 33.800 ;
        RECT 139.400 33.600 139.800 33.800 ;
        RECT 142.200 33.600 142.600 35.300 ;
        RECT 143.900 35.200 144.300 35.300 ;
        RECT 145.500 35.200 145.800 35.800 ;
        RECT 146.500 35.900 146.800 36.500 ;
        RECT 147.100 36.500 147.500 36.600 ;
        RECT 149.400 36.500 149.800 36.600 ;
        RECT 147.100 36.200 149.800 36.500 ;
        RECT 146.500 35.700 148.900 35.900 ;
        RECT 151.000 35.700 151.400 39.900 ;
        RECT 153.100 35.900 154.100 39.900 ;
        RECT 157.700 39.200 158.100 39.900 ;
        RECT 157.400 38.800 158.100 39.200 ;
        RECT 157.700 36.400 158.100 38.800 ;
        RECT 159.800 37.500 160.200 39.500 ;
        RECT 157.300 36.100 158.100 36.400 ;
        RECT 146.500 35.600 151.400 35.700 ;
        RECT 148.500 35.500 151.400 35.600 ;
        RECT 148.600 35.400 151.400 35.500 ;
        RECT 143.100 34.900 143.500 35.000 ;
        RECT 143.100 34.600 145.000 34.900 ;
        RECT 145.400 34.800 145.800 35.200 ;
        RECT 147.800 35.100 148.200 35.200 ;
        RECT 147.800 34.800 150.300 35.100 ;
        RECT 144.600 34.500 145.000 34.600 ;
        RECT 145.500 34.200 145.800 34.800 ;
        RECT 149.900 34.700 150.300 34.800 ;
        RECT 152.600 34.400 153.000 35.200 ;
        RECT 149.100 34.200 149.500 34.300 ;
        RECT 153.400 34.200 153.700 35.900 ;
        RECT 154.200 34.400 154.600 35.200 ;
        RECT 155.800 35.100 156.200 35.200 ;
        RECT 156.600 35.100 157.000 35.600 ;
        RECT 155.800 34.800 157.000 35.100 ;
        RECT 145.500 33.900 151.000 34.200 ;
        RECT 145.700 33.800 146.100 33.900 ;
        RECT 142.200 33.300 144.100 33.600 ;
        RECT 138.300 33.100 140.100 33.300 ;
        RECT 130.200 31.500 130.600 32.500 ;
        RECT 132.300 31.500 132.700 33.000 ;
        RECT 135.800 32.800 136.700 33.100 ;
        RECT 136.300 31.100 136.700 32.800 ;
        RECT 137.400 31.100 137.800 33.100 ;
        RECT 138.200 33.000 140.200 33.100 ;
        RECT 138.200 31.100 138.600 33.000 ;
        RECT 139.800 31.100 140.200 33.000 ;
        RECT 142.200 31.100 142.600 33.300 ;
        RECT 143.700 33.200 144.100 33.300 ;
        RECT 148.600 32.800 148.900 33.900 ;
        RECT 150.200 33.800 151.000 33.900 ;
        RECT 151.800 34.100 152.200 34.200 ;
        RECT 153.400 34.100 153.800 34.200 ;
        RECT 151.800 33.800 152.600 34.100 ;
        RECT 153.400 33.800 154.600 34.100 ;
        RECT 155.000 33.800 155.400 34.600 ;
        RECT 157.300 34.200 157.600 36.100 ;
        RECT 159.900 35.800 160.200 37.500 ;
        RECT 158.300 35.500 160.200 35.800 ;
        RECT 158.300 34.500 158.600 35.500 ;
        RECT 156.600 33.800 157.600 34.200 ;
        RECT 157.900 34.100 158.600 34.500 ;
        RECT 159.000 34.400 159.400 35.200 ;
        RECT 159.800 35.100 160.200 35.200 ;
        RECT 160.600 35.100 161.000 35.200 ;
        RECT 159.800 34.800 161.000 35.100 ;
        RECT 159.800 34.400 160.200 34.800 ;
        RECT 152.200 33.600 152.600 33.800 ;
        RECT 147.700 32.700 148.100 32.800 ;
        RECT 144.600 32.100 145.000 32.500 ;
        RECT 146.700 32.400 148.100 32.700 ;
        RECT 148.600 32.400 149.000 32.800 ;
        RECT 146.700 32.100 147.000 32.400 ;
        RECT 149.400 32.100 149.800 32.500 ;
        RECT 144.300 31.800 145.000 32.100 ;
        RECT 144.300 31.100 144.900 31.800 ;
        RECT 146.600 31.100 147.000 32.100 ;
        RECT 148.800 31.800 149.800 32.100 ;
        RECT 148.800 31.100 149.200 31.800 ;
        RECT 151.000 31.100 151.400 33.500 ;
        RECT 151.900 33.100 153.700 33.300 ;
        RECT 154.300 33.100 154.600 33.800 ;
        RECT 157.300 33.500 157.600 33.800 ;
        RECT 158.100 33.900 158.600 34.100 ;
        RECT 158.100 33.600 160.200 33.900 ;
        RECT 157.300 33.300 157.700 33.500 ;
        RECT 151.800 33.000 153.800 33.100 ;
        RECT 151.800 31.100 152.200 33.000 ;
        RECT 153.400 31.400 153.800 33.000 ;
        RECT 154.200 31.700 154.600 33.100 ;
        RECT 155.000 31.400 155.400 33.100 ;
        RECT 157.300 33.000 158.100 33.300 ;
        RECT 157.700 31.500 158.100 33.000 ;
        RECT 159.900 32.500 160.200 33.600 ;
        RECT 160.600 33.400 161.000 34.200 ;
        RECT 161.400 33.100 161.800 39.900 ;
        RECT 163.000 37.100 163.400 37.200 ;
        RECT 163.800 37.100 164.200 39.900 ;
        RECT 163.000 36.800 164.200 37.100 ;
        RECT 162.200 35.800 162.600 36.600 ;
        RECT 163.000 33.400 163.400 34.200 ;
        RECT 163.800 33.100 164.200 36.800 ;
        RECT 164.600 35.800 165.000 36.600 ;
        RECT 166.700 36.200 167.100 39.900 ;
        RECT 167.400 36.800 167.800 37.200 ;
        RECT 167.500 36.200 167.800 36.800 ;
        RECT 166.700 35.900 167.200 36.200 ;
        RECT 167.500 35.900 168.200 36.200 ;
        RECT 164.600 35.100 164.900 35.800 ;
        RECT 166.200 35.100 166.600 35.200 ;
        RECT 164.600 34.800 166.600 35.100 ;
        RECT 166.200 34.400 166.600 34.800 ;
        RECT 166.900 34.200 167.200 35.900 ;
        RECT 167.800 35.800 168.200 35.900 ;
        RECT 165.400 34.100 165.800 34.200 ;
        RECT 165.400 33.800 166.200 34.100 ;
        RECT 166.900 33.800 168.200 34.200 ;
        RECT 165.800 33.600 166.200 33.800 ;
        RECT 165.500 33.100 167.300 33.300 ;
        RECT 167.800 33.200 168.100 33.800 ;
        RECT 161.400 32.800 162.300 33.100 ;
        RECT 163.800 32.800 164.700 33.100 ;
        RECT 159.800 31.500 160.200 32.500 ;
        RECT 161.900 32.200 162.300 32.800 ;
        RECT 161.400 31.800 162.300 32.200 ;
        RECT 153.400 31.100 155.400 31.400 ;
        RECT 161.900 31.100 162.300 31.800 ;
        RECT 164.300 31.100 164.700 32.800 ;
        RECT 165.400 33.000 167.400 33.100 ;
        RECT 165.400 31.100 165.800 33.000 ;
        RECT 167.000 31.100 167.400 33.000 ;
        RECT 167.800 31.100 168.200 33.200 ;
        RECT 168.600 31.100 169.000 39.900 ;
        RECT 171.000 36.400 171.400 39.900 ;
        RECT 170.900 35.900 171.400 36.400 ;
        RECT 172.600 36.200 173.000 39.900 ;
        RECT 171.700 35.900 173.000 36.200 ;
        RECT 170.900 34.200 171.200 35.900 ;
        RECT 171.700 34.900 172.000 35.900 ;
        RECT 171.500 34.500 172.000 34.900 ;
        RECT 170.900 33.800 171.400 34.200 ;
        RECT 169.400 32.400 169.800 33.200 ;
        RECT 170.900 33.100 171.200 33.800 ;
        RECT 171.700 33.700 172.000 34.500 ;
        RECT 172.500 35.100 173.000 35.200 ;
        RECT 173.400 35.100 173.800 35.200 ;
        RECT 172.500 34.800 173.800 35.100 ;
        RECT 174.200 35.100 174.600 39.900 ;
        RECT 176.200 36.800 176.600 37.200 ;
        RECT 175.000 35.800 175.400 36.600 ;
        RECT 176.200 36.200 176.500 36.800 ;
        RECT 176.900 36.200 177.300 39.900 ;
        RECT 175.800 35.900 176.500 36.200 ;
        RECT 176.800 35.900 177.300 36.200 ;
        RECT 179.000 37.500 179.400 39.500 ;
        RECT 175.800 35.800 176.200 35.900 ;
        RECT 175.800 35.100 176.100 35.800 ;
        RECT 174.200 34.800 176.100 35.100 ;
        RECT 172.500 34.400 172.900 34.800 ;
        RECT 171.700 33.400 173.000 33.700 ;
        RECT 173.400 33.400 173.800 34.200 ;
        RECT 170.900 32.800 171.400 33.100 ;
        RECT 171.000 31.100 171.400 32.800 ;
        RECT 172.600 31.100 173.000 33.400 ;
        RECT 174.200 33.100 174.600 34.800 ;
        RECT 176.800 34.200 177.100 35.900 ;
        RECT 179.000 35.800 179.300 37.500 ;
        RECT 181.100 36.400 181.500 39.900 ;
        RECT 181.100 36.100 181.900 36.400 ;
        RECT 179.000 35.500 180.900 35.800 ;
        RECT 177.400 34.400 177.800 35.200 ;
        RECT 179.000 34.400 179.400 35.200 ;
        RECT 179.800 34.400 180.200 35.200 ;
        RECT 180.600 34.500 180.900 35.500 ;
        RECT 175.800 33.800 177.100 34.200 ;
        RECT 178.200 34.100 178.600 34.200 ;
        RECT 177.800 33.800 178.600 34.100 ;
        RECT 180.600 34.100 181.300 34.500 ;
        RECT 181.600 34.200 181.900 36.100 ;
        RECT 182.200 35.100 182.600 35.600 ;
        RECT 183.000 35.100 183.400 35.200 ;
        RECT 182.200 34.800 183.400 35.100 ;
        RECT 180.600 33.900 181.100 34.100 ;
        RECT 175.900 33.100 176.200 33.800 ;
        RECT 177.800 33.600 178.200 33.800 ;
        RECT 179.000 33.600 181.100 33.900 ;
        RECT 181.600 33.800 182.600 34.200 ;
        RECT 176.700 33.100 178.500 33.300 ;
        RECT 174.200 32.800 175.100 33.100 ;
        RECT 174.700 31.100 175.100 32.800 ;
        RECT 175.800 31.100 176.200 33.100 ;
        RECT 176.600 33.000 178.600 33.100 ;
        RECT 176.600 31.100 177.000 33.000 ;
        RECT 178.200 31.100 178.600 33.000 ;
        RECT 179.000 32.500 179.300 33.600 ;
        RECT 181.600 33.500 181.900 33.800 ;
        RECT 181.500 33.300 181.900 33.500 ;
        RECT 181.100 33.000 181.900 33.300 ;
        RECT 179.000 31.500 179.400 32.500 ;
        RECT 181.100 31.500 181.500 33.000 ;
        RECT 183.800 31.100 184.200 39.900 ;
        RECT 185.400 35.600 185.800 39.900 ;
        RECT 187.500 37.900 188.100 39.900 ;
        RECT 189.800 37.900 190.200 39.900 ;
        RECT 192.000 38.200 192.400 39.900 ;
        RECT 192.000 37.900 193.000 38.200 ;
        RECT 187.800 37.500 188.200 37.900 ;
        RECT 189.900 37.600 190.200 37.900 ;
        RECT 189.500 37.300 191.300 37.600 ;
        RECT 192.600 37.500 193.000 37.900 ;
        RECT 189.500 37.200 189.900 37.300 ;
        RECT 190.900 37.200 191.300 37.300 ;
        RECT 187.400 36.600 188.100 37.000 ;
        RECT 187.800 36.100 188.100 36.600 ;
        RECT 188.900 36.500 190.000 36.800 ;
        RECT 188.900 36.400 189.300 36.500 ;
        RECT 187.800 35.800 189.000 36.100 ;
        RECT 185.400 35.300 187.500 35.600 ;
        RECT 185.400 33.600 185.800 35.300 ;
        RECT 187.100 35.200 187.500 35.300 ;
        RECT 186.300 34.900 186.700 35.000 ;
        RECT 186.300 34.600 188.200 34.900 ;
        RECT 187.800 34.500 188.200 34.600 ;
        RECT 188.700 34.200 189.000 35.800 ;
        RECT 189.700 35.900 190.000 36.500 ;
        RECT 190.300 36.500 190.700 36.600 ;
        RECT 192.600 36.500 193.000 36.600 ;
        RECT 190.300 36.200 193.000 36.500 ;
        RECT 189.700 35.700 192.100 35.900 ;
        RECT 194.200 35.700 194.600 39.900 ;
        RECT 197.900 36.200 198.300 39.900 ;
        RECT 198.600 36.800 199.000 37.200 ;
        RECT 198.700 36.200 199.000 36.800 ;
        RECT 201.100 36.200 201.500 39.900 ;
        RECT 201.800 36.800 202.200 37.200 ;
        RECT 201.900 36.200 202.200 36.800 ;
        RECT 197.900 35.900 198.400 36.200 ;
        RECT 198.700 35.900 199.400 36.200 ;
        RECT 201.100 35.900 201.600 36.200 ;
        RECT 201.900 35.900 202.600 36.200 ;
        RECT 189.700 35.600 194.600 35.700 ;
        RECT 191.700 35.500 194.600 35.600 ;
        RECT 191.800 35.400 194.600 35.500 ;
        RECT 198.100 35.200 198.400 35.900 ;
        RECT 199.000 35.800 199.400 35.900 ;
        RECT 191.000 35.100 191.400 35.200 ;
        RECT 191.000 34.800 193.500 35.100 ;
        RECT 193.100 34.700 193.500 34.800 ;
        RECT 197.400 34.400 197.800 35.200 ;
        RECT 198.100 34.800 198.600 35.200 ;
        RECT 192.300 34.200 192.700 34.300 ;
        RECT 198.100 34.200 198.400 34.800 ;
        RECT 200.600 34.400 201.000 35.200 ;
        RECT 201.300 34.200 201.600 35.900 ;
        RECT 202.200 35.800 202.600 35.900 ;
        RECT 203.000 35.800 203.400 36.600 ;
        RECT 202.200 35.100 202.500 35.800 ;
        RECT 203.800 35.100 204.200 39.900 ;
        RECT 202.200 34.800 204.200 35.100 ;
        RECT 188.700 33.900 194.200 34.200 ;
        RECT 188.900 33.800 189.300 33.900 ;
        RECT 191.800 33.800 192.200 33.900 ;
        RECT 193.400 33.800 194.200 33.900 ;
        RECT 196.600 34.100 197.000 34.200 ;
        RECT 196.600 33.800 197.400 34.100 ;
        RECT 198.100 33.800 199.400 34.200 ;
        RECT 199.800 34.100 200.200 34.200 ;
        RECT 199.800 33.800 200.600 34.100 ;
        RECT 201.300 33.800 202.600 34.200 ;
        RECT 185.400 33.300 187.300 33.600 ;
        RECT 184.600 32.400 185.000 33.200 ;
        RECT 185.400 31.100 185.800 33.300 ;
        RECT 186.900 33.200 187.300 33.300 ;
        RECT 191.800 32.800 192.100 33.800 ;
        RECT 197.000 33.600 197.400 33.800 ;
        RECT 190.900 32.700 191.300 32.800 ;
        RECT 187.800 32.100 188.200 32.500 ;
        RECT 189.900 32.400 191.300 32.700 ;
        RECT 191.800 32.400 192.200 32.800 ;
        RECT 189.900 32.100 190.200 32.400 ;
        RECT 192.600 32.100 193.000 32.500 ;
        RECT 187.500 31.800 188.200 32.100 ;
        RECT 187.500 31.100 188.100 31.800 ;
        RECT 189.800 31.100 190.200 32.100 ;
        RECT 192.000 31.800 193.000 32.100 ;
        RECT 192.000 31.100 192.400 31.800 ;
        RECT 194.200 31.100 194.600 33.500 ;
        RECT 196.700 33.100 198.500 33.300 ;
        RECT 199.000 33.100 199.300 33.800 ;
        RECT 200.200 33.600 200.600 33.800 ;
        RECT 199.900 33.100 201.700 33.300 ;
        RECT 202.200 33.100 202.500 33.800 ;
        RECT 203.800 33.100 204.200 34.800 ;
        RECT 205.400 35.600 205.800 39.900 ;
        RECT 207.500 37.900 208.100 39.900 ;
        RECT 209.800 37.900 210.200 39.900 ;
        RECT 212.000 38.200 212.400 39.900 ;
        RECT 212.000 37.900 213.000 38.200 ;
        RECT 207.800 37.500 208.200 37.900 ;
        RECT 209.900 37.600 210.200 37.900 ;
        RECT 209.500 37.300 211.300 37.600 ;
        RECT 212.600 37.500 213.000 37.900 ;
        RECT 209.500 37.200 209.900 37.300 ;
        RECT 210.900 37.200 211.300 37.300 ;
        RECT 207.400 36.600 208.100 37.000 ;
        RECT 207.800 36.100 208.100 36.600 ;
        RECT 208.900 36.500 210.000 36.800 ;
        RECT 208.900 36.400 209.300 36.500 ;
        RECT 207.800 35.800 209.000 36.100 ;
        RECT 205.400 35.300 207.500 35.600 ;
        RECT 204.600 33.400 205.000 34.200 ;
        RECT 205.400 33.600 205.800 35.300 ;
        RECT 207.100 35.200 207.500 35.300 ;
        RECT 206.300 34.900 206.700 35.000 ;
        RECT 206.300 34.600 208.200 34.900 ;
        RECT 207.800 34.500 208.200 34.600 ;
        RECT 208.700 34.200 209.000 35.800 ;
        RECT 209.700 35.900 210.000 36.500 ;
        RECT 210.300 36.500 210.700 36.600 ;
        RECT 212.600 36.500 213.000 36.600 ;
        RECT 210.300 36.200 213.000 36.500 ;
        RECT 209.700 35.700 212.100 35.900 ;
        RECT 214.200 35.700 214.600 39.900 ;
        RECT 216.300 36.200 216.700 39.900 ;
        RECT 217.000 36.800 217.400 37.200 ;
        RECT 217.100 36.200 217.400 36.800 ;
        RECT 216.300 35.900 216.800 36.200 ;
        RECT 217.100 35.900 217.800 36.200 ;
        RECT 209.700 35.600 214.600 35.700 ;
        RECT 211.700 35.500 214.600 35.600 ;
        RECT 211.800 35.400 214.600 35.500 ;
        RECT 211.000 35.100 211.400 35.200 ;
        RECT 211.000 34.800 213.500 35.100 ;
        RECT 211.800 34.700 212.200 34.800 ;
        RECT 213.100 34.700 213.500 34.800 ;
        RECT 215.800 34.400 216.200 35.200 ;
        RECT 212.300 34.200 212.700 34.300 ;
        RECT 216.500 34.200 216.800 35.900 ;
        RECT 217.400 35.800 217.800 35.900 ;
        RECT 218.200 35.800 218.600 36.600 ;
        RECT 217.400 35.100 217.700 35.800 ;
        RECT 219.000 35.100 219.400 39.900 ;
        RECT 219.800 37.100 220.200 37.200 ;
        RECT 220.600 37.100 221.000 39.900 ;
        RECT 222.700 37.900 223.300 39.900 ;
        RECT 225.000 37.900 225.400 39.900 ;
        RECT 227.200 38.200 227.600 39.900 ;
        RECT 227.200 37.900 228.200 38.200 ;
        RECT 223.000 37.500 223.400 37.900 ;
        RECT 225.100 37.600 225.400 37.900 ;
        RECT 224.700 37.300 226.500 37.600 ;
        RECT 227.800 37.500 228.200 37.900 ;
        RECT 224.700 37.200 225.100 37.300 ;
        RECT 226.100 37.200 226.500 37.300 ;
        RECT 219.800 36.800 221.000 37.100 ;
        RECT 217.400 34.800 219.400 35.100 ;
        RECT 208.700 33.900 214.200 34.200 ;
        RECT 208.900 33.800 209.300 33.900 ;
        RECT 196.600 33.000 198.600 33.100 ;
        RECT 196.600 31.100 197.000 33.000 ;
        RECT 198.200 31.100 198.600 33.000 ;
        RECT 199.000 31.100 199.400 33.100 ;
        RECT 199.800 33.000 201.800 33.100 ;
        RECT 199.800 31.100 200.200 33.000 ;
        RECT 201.400 31.100 201.800 33.000 ;
        RECT 202.200 31.100 202.600 33.100 ;
        RECT 203.300 32.800 204.200 33.100 ;
        RECT 205.400 33.300 207.300 33.600 ;
        RECT 203.300 31.100 203.700 32.800 ;
        RECT 205.400 31.100 205.800 33.300 ;
        RECT 206.900 33.200 207.300 33.300 ;
        RECT 211.800 32.800 212.100 33.900 ;
        RECT 213.400 33.800 214.200 33.900 ;
        RECT 215.000 34.100 215.400 34.200 ;
        RECT 216.500 34.100 217.800 34.200 ;
        RECT 218.200 34.100 218.600 34.200 ;
        RECT 215.000 33.800 215.800 34.100 ;
        RECT 216.500 33.800 218.600 34.100 ;
        RECT 215.400 33.600 215.800 33.800 ;
        RECT 210.900 32.700 211.300 32.800 ;
        RECT 207.800 32.100 208.200 32.500 ;
        RECT 209.900 32.400 211.300 32.700 ;
        RECT 211.800 32.400 212.200 32.800 ;
        RECT 209.900 32.100 210.200 32.400 ;
        RECT 212.600 32.100 213.000 32.500 ;
        RECT 207.500 31.800 208.200 32.100 ;
        RECT 207.500 31.100 208.100 31.800 ;
        RECT 209.800 31.100 210.200 32.100 ;
        RECT 212.000 31.800 213.000 32.100 ;
        RECT 212.000 31.100 212.400 31.800 ;
        RECT 214.200 31.100 214.600 33.500 ;
        RECT 215.100 33.100 216.900 33.300 ;
        RECT 217.400 33.100 217.700 33.800 ;
        RECT 219.000 33.100 219.400 34.800 ;
        RECT 220.600 35.600 221.000 36.800 ;
        RECT 222.600 36.600 223.300 37.000 ;
        RECT 223.000 36.100 223.300 36.600 ;
        RECT 224.100 36.500 225.200 36.800 ;
        RECT 224.100 36.400 224.500 36.500 ;
        RECT 223.000 35.800 224.200 36.100 ;
        RECT 220.600 35.300 222.700 35.600 ;
        RECT 219.800 33.400 220.200 34.200 ;
        RECT 220.600 33.600 221.000 35.300 ;
        RECT 222.300 35.200 222.700 35.300 ;
        RECT 223.900 35.100 224.200 35.800 ;
        RECT 224.900 35.900 225.200 36.500 ;
        RECT 225.500 36.500 225.900 36.600 ;
        RECT 227.800 36.500 228.200 36.600 ;
        RECT 225.500 36.200 228.200 36.500 ;
        RECT 224.900 35.700 227.300 35.900 ;
        RECT 229.400 35.700 229.800 39.900 ;
        RECT 224.900 35.600 229.800 35.700 ;
        RECT 226.900 35.500 229.800 35.600 ;
        RECT 227.000 35.400 229.800 35.500 ;
        RECT 224.600 35.100 225.000 35.200 ;
        RECT 221.500 34.900 221.900 35.000 ;
        RECT 221.500 34.600 223.400 34.900 ;
        RECT 223.800 34.800 225.000 35.100 ;
        RECT 226.200 35.100 226.600 35.200 ;
        RECT 226.200 34.800 228.700 35.100 ;
        RECT 223.000 34.500 223.400 34.600 ;
        RECT 223.900 34.200 224.200 34.800 ;
        RECT 228.300 34.700 228.700 34.800 ;
        RECT 227.500 34.200 227.900 34.300 ;
        RECT 223.900 33.900 229.400 34.200 ;
        RECT 224.100 33.800 224.500 33.900 ;
        RECT 215.000 33.000 217.000 33.100 ;
        RECT 215.000 31.100 215.400 33.000 ;
        RECT 216.600 31.100 217.000 33.000 ;
        RECT 217.400 31.100 217.800 33.100 ;
        RECT 218.500 32.800 219.400 33.100 ;
        RECT 220.600 33.300 222.500 33.600 ;
        RECT 218.500 31.100 218.900 32.800 ;
        RECT 220.600 31.100 221.000 33.300 ;
        RECT 222.100 33.200 222.500 33.300 ;
        RECT 227.000 32.800 227.300 33.900 ;
        RECT 228.600 33.800 229.400 33.900 ;
        RECT 226.100 32.700 226.500 32.800 ;
        RECT 223.000 32.100 223.400 32.500 ;
        RECT 225.100 32.400 226.500 32.700 ;
        RECT 227.000 32.400 227.400 32.800 ;
        RECT 225.100 32.100 225.400 32.400 ;
        RECT 227.800 32.100 228.200 32.500 ;
        RECT 222.700 31.800 223.400 32.100 ;
        RECT 222.700 31.100 223.300 31.800 ;
        RECT 225.000 31.100 225.400 32.100 ;
        RECT 227.200 31.800 228.200 32.100 ;
        RECT 227.200 31.100 227.600 31.800 ;
        RECT 229.400 31.100 229.800 33.500 ;
        RECT 0.600 27.900 1.000 29.900 ;
        RECT 1.400 28.000 1.800 29.900 ;
        RECT 3.000 28.000 3.400 29.900 ;
        RECT 1.400 27.900 3.400 28.000 ;
        RECT 0.700 27.200 1.000 27.900 ;
        RECT 1.500 27.700 3.300 27.900 ;
        RECT 3.800 27.700 4.200 29.900 ;
        RECT 5.900 29.200 6.500 29.900 ;
        RECT 5.900 28.900 6.600 29.200 ;
        RECT 8.200 28.900 8.600 29.900 ;
        RECT 10.400 29.200 10.800 29.900 ;
        RECT 10.400 28.900 11.400 29.200 ;
        RECT 6.200 28.500 6.600 28.900 ;
        RECT 8.300 28.600 8.600 28.900 ;
        RECT 8.300 28.300 9.700 28.600 ;
        RECT 9.300 28.200 9.700 28.300 ;
        RECT 10.200 28.200 10.600 28.600 ;
        RECT 11.000 28.500 11.400 28.900 ;
        RECT 5.300 27.700 5.700 27.800 ;
        RECT 3.800 27.400 5.700 27.700 ;
        RECT 2.600 27.200 3.000 27.400 ;
        RECT 0.600 26.800 1.900 27.200 ;
        RECT 2.600 26.900 3.400 27.200 ;
        RECT 3.000 26.800 3.400 26.900 ;
        RECT 1.600 25.200 1.900 26.800 ;
        RECT 2.200 25.800 2.600 26.600 ;
        RECT 3.800 25.700 4.200 27.400 ;
        RECT 7.300 27.100 7.700 27.200 ;
        RECT 10.200 27.100 10.500 28.200 ;
        RECT 12.600 27.500 13.000 29.900 ;
        RECT 13.400 27.700 13.800 29.900 ;
        RECT 15.500 29.200 16.100 29.900 ;
        RECT 15.500 28.900 16.200 29.200 ;
        RECT 17.800 28.900 18.200 29.900 ;
        RECT 20.000 29.200 20.400 29.900 ;
        RECT 20.000 28.900 21.000 29.200 ;
        RECT 15.800 28.500 16.200 28.900 ;
        RECT 17.900 28.600 18.200 28.900 ;
        RECT 17.900 28.300 19.300 28.600 ;
        RECT 18.900 28.200 19.300 28.300 ;
        RECT 19.800 28.200 20.200 28.600 ;
        RECT 20.600 28.500 21.000 28.900 ;
        RECT 14.900 27.700 15.300 27.800 ;
        RECT 13.400 27.400 15.300 27.700 ;
        RECT 11.800 27.100 12.600 27.200 ;
        RECT 7.100 26.800 12.600 27.100 ;
        RECT 6.200 26.400 6.600 26.500 ;
        RECT 4.700 26.100 6.600 26.400 ;
        RECT 4.700 26.000 5.100 26.100 ;
        RECT 5.500 25.700 5.900 25.800 ;
        RECT 3.800 25.400 5.900 25.700 ;
        RECT 0.600 25.100 1.000 25.200 ;
        RECT 0.600 24.800 1.300 25.100 ;
        RECT 1.600 24.800 2.600 25.200 ;
        RECT 1.000 24.200 1.300 24.800 ;
        RECT 1.000 23.800 1.400 24.200 ;
        RECT 1.700 21.100 2.100 24.800 ;
        RECT 3.800 21.100 4.200 25.400 ;
        RECT 7.100 25.200 7.400 26.800 ;
        RECT 10.700 26.700 11.100 26.800 ;
        RECT 11.500 26.200 11.900 26.300 ;
        RECT 9.400 25.900 11.900 26.200 ;
        RECT 9.400 25.800 9.800 25.900 ;
        RECT 13.400 25.700 13.800 27.400 ;
        RECT 16.900 27.100 17.300 27.200 ;
        RECT 19.000 27.100 19.400 27.200 ;
        RECT 19.800 27.100 20.100 28.200 ;
        RECT 22.200 27.500 22.600 29.900 ;
        RECT 23.000 27.800 23.400 28.600 ;
        RECT 21.400 27.100 22.200 27.200 ;
        RECT 16.700 26.800 22.200 27.100 ;
        RECT 15.800 26.400 16.200 26.500 ;
        RECT 14.300 26.100 16.200 26.400 ;
        RECT 14.300 26.000 14.700 26.100 ;
        RECT 15.100 25.700 15.500 25.800 ;
        RECT 10.200 25.500 13.000 25.600 ;
        RECT 10.100 25.400 13.000 25.500 ;
        RECT 6.200 24.900 7.400 25.200 ;
        RECT 8.100 25.300 13.000 25.400 ;
        RECT 8.100 25.100 10.500 25.300 ;
        RECT 6.200 24.400 6.500 24.900 ;
        RECT 5.800 24.200 6.500 24.400 ;
        RECT 7.300 24.500 7.700 24.600 ;
        RECT 8.100 24.500 8.400 25.100 ;
        RECT 7.300 24.200 8.400 24.500 ;
        RECT 8.700 24.500 11.400 24.800 ;
        RECT 8.700 24.400 9.100 24.500 ;
        RECT 11.000 24.400 11.400 24.500 ;
        RECT 5.400 24.000 6.500 24.200 ;
        RECT 5.400 23.800 6.100 24.000 ;
        RECT 7.900 23.700 8.300 23.800 ;
        RECT 9.300 23.700 9.700 23.800 ;
        RECT 6.200 23.100 6.600 23.500 ;
        RECT 7.900 23.400 9.700 23.700 ;
        RECT 8.300 23.100 8.600 23.400 ;
        RECT 11.000 23.100 11.400 23.500 ;
        RECT 5.900 21.100 6.500 23.100 ;
        RECT 8.200 21.100 8.600 23.100 ;
        RECT 10.400 22.800 11.400 23.100 ;
        RECT 10.400 21.100 10.800 22.800 ;
        RECT 12.600 21.100 13.000 25.300 ;
        RECT 13.400 25.400 15.500 25.700 ;
        RECT 13.400 21.100 13.800 25.400 ;
        RECT 16.700 25.200 17.000 26.800 ;
        RECT 20.300 26.700 20.700 26.800 ;
        RECT 21.100 26.200 21.500 26.300 ;
        RECT 17.400 26.100 17.800 26.200 ;
        RECT 19.000 26.100 21.500 26.200 ;
        RECT 17.400 25.900 21.500 26.100 ;
        RECT 17.400 25.800 19.400 25.900 ;
        RECT 19.800 25.500 22.600 25.600 ;
        RECT 19.700 25.400 22.600 25.500 ;
        RECT 15.800 24.900 17.000 25.200 ;
        RECT 17.700 25.300 22.600 25.400 ;
        RECT 17.700 25.100 20.100 25.300 ;
        RECT 15.800 24.400 16.100 24.900 ;
        RECT 15.400 24.000 16.100 24.400 ;
        RECT 16.900 24.500 17.300 24.600 ;
        RECT 17.700 24.500 18.000 25.100 ;
        RECT 16.900 24.200 18.000 24.500 ;
        RECT 18.300 24.500 21.000 24.800 ;
        RECT 18.300 24.400 18.700 24.500 ;
        RECT 20.600 24.400 21.000 24.500 ;
        RECT 17.500 23.700 17.900 23.800 ;
        RECT 18.900 23.700 19.300 23.800 ;
        RECT 15.800 23.100 16.200 23.500 ;
        RECT 17.500 23.400 19.300 23.700 ;
        RECT 17.900 23.100 18.200 23.400 ;
        RECT 20.600 23.100 21.000 23.500 ;
        RECT 15.500 21.100 16.100 23.100 ;
        RECT 17.800 21.100 18.200 23.100 ;
        RECT 20.000 22.800 21.000 23.100 ;
        RECT 20.000 21.100 20.400 22.800 ;
        RECT 22.200 21.100 22.600 25.300 ;
        RECT 23.800 21.100 24.200 29.900 ;
        RECT 25.900 28.200 26.300 29.900 ;
        RECT 25.400 27.900 26.300 28.200 ;
        RECT 27.000 27.900 27.400 29.900 ;
        RECT 27.800 28.000 28.200 29.900 ;
        RECT 29.400 28.000 29.800 29.900 ;
        RECT 27.800 27.900 29.800 28.000 ;
        RECT 24.600 26.800 25.000 27.600 ;
        RECT 25.400 26.100 25.800 27.900 ;
        RECT 27.100 27.200 27.400 27.900 ;
        RECT 27.900 27.700 29.700 27.900 ;
        RECT 31.000 27.600 31.400 29.900 ;
        RECT 32.600 27.600 33.000 29.900 ;
        RECT 34.200 27.600 34.600 29.900 ;
        RECT 35.800 27.600 36.200 29.900 ;
        RECT 29.000 27.200 29.400 27.400 ;
        RECT 30.200 27.200 31.400 27.600 ;
        RECT 31.900 27.200 33.000 27.600 ;
        RECT 33.500 27.200 34.600 27.600 ;
        RECT 35.300 27.200 36.200 27.600 ;
        RECT 39.000 27.700 39.400 29.900 ;
        RECT 41.100 29.200 41.700 29.900 ;
        RECT 41.100 28.900 41.800 29.200 ;
        RECT 43.400 28.900 43.800 29.900 ;
        RECT 45.600 29.200 46.000 29.900 ;
        RECT 45.600 28.900 46.600 29.200 ;
        RECT 41.400 28.500 41.800 28.900 ;
        RECT 43.500 28.600 43.800 28.900 ;
        RECT 43.500 28.300 44.900 28.600 ;
        RECT 44.500 28.200 44.900 28.300 ;
        RECT 45.400 28.200 45.800 28.600 ;
        RECT 46.200 28.500 46.600 28.900 ;
        RECT 40.500 27.700 40.900 27.800 ;
        RECT 39.000 27.400 40.900 27.700 ;
        RECT 27.000 26.800 28.300 27.200 ;
        RECT 29.000 26.900 29.800 27.200 ;
        RECT 29.400 26.800 29.800 26.900 ;
        RECT 25.400 25.800 27.300 26.100 ;
        RECT 25.400 21.100 25.800 25.800 ;
        RECT 27.000 25.200 27.300 25.800 ;
        RECT 26.200 24.400 26.600 25.200 ;
        RECT 27.000 25.100 27.400 25.200 ;
        RECT 28.000 25.100 28.300 26.800 ;
        RECT 28.600 25.800 29.000 26.600 ;
        RECT 30.200 25.800 30.600 27.200 ;
        RECT 31.900 26.900 32.300 27.200 ;
        RECT 33.500 26.900 33.900 27.200 ;
        RECT 35.300 26.900 35.700 27.200 ;
        RECT 31.000 26.500 32.300 26.900 ;
        RECT 32.700 26.500 33.900 26.900 ;
        RECT 34.400 26.500 35.700 26.900 ;
        RECT 31.900 25.800 32.300 26.500 ;
        RECT 33.500 25.800 33.900 26.500 ;
        RECT 35.300 25.800 35.700 26.500 ;
        RECT 30.200 25.400 31.400 25.800 ;
        RECT 31.900 25.400 33.000 25.800 ;
        RECT 33.500 25.400 34.600 25.800 ;
        RECT 35.300 25.400 36.200 25.800 ;
        RECT 27.000 24.800 27.700 25.100 ;
        RECT 28.000 24.800 28.500 25.100 ;
        RECT 27.400 24.200 27.700 24.800 ;
        RECT 27.400 23.800 27.800 24.200 ;
        RECT 28.100 21.100 28.500 24.800 ;
        RECT 31.000 21.100 31.400 25.400 ;
        RECT 32.600 21.100 33.000 25.400 ;
        RECT 34.200 21.100 34.600 25.400 ;
        RECT 35.800 21.100 36.200 25.400 ;
        RECT 39.000 25.700 39.400 27.400 ;
        RECT 42.500 27.100 42.900 27.200 ;
        RECT 45.400 27.100 45.700 28.200 ;
        RECT 47.800 27.500 48.200 29.900 ;
        RECT 48.600 28.000 49.000 29.900 ;
        RECT 50.200 28.000 50.600 29.900 ;
        RECT 48.600 27.900 50.600 28.000 ;
        RECT 51.000 27.900 51.400 29.900 ;
        RECT 53.100 28.200 53.500 29.900 ;
        RECT 55.500 28.200 55.900 29.900 ;
        RECT 52.600 27.900 53.500 28.200 ;
        RECT 55.000 27.900 55.900 28.200 ;
        RECT 56.600 27.900 57.000 29.900 ;
        RECT 57.400 28.000 57.800 29.900 ;
        RECT 59.000 28.000 59.400 29.900 ;
        RECT 57.400 27.900 59.400 28.000 ;
        RECT 48.700 27.700 50.500 27.900 ;
        RECT 49.000 27.200 49.400 27.400 ;
        RECT 51.000 27.200 51.300 27.900 ;
        RECT 47.000 27.100 47.800 27.200 ;
        RECT 42.300 26.800 47.800 27.100 ;
        RECT 48.600 26.900 49.400 27.200 ;
        RECT 48.600 26.800 49.000 26.900 ;
        RECT 50.100 26.800 51.400 27.200 ;
        RECT 51.800 26.800 52.200 27.600 ;
        RECT 41.400 26.400 41.800 26.500 ;
        RECT 39.900 26.100 41.800 26.400 ;
        RECT 42.300 26.200 42.600 26.800 ;
        RECT 45.900 26.700 46.300 26.800 ;
        RECT 45.400 26.200 45.800 26.300 ;
        RECT 46.700 26.200 47.100 26.300 ;
        RECT 39.900 26.000 40.300 26.100 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 44.600 25.900 47.100 26.200 ;
        RECT 44.600 25.800 45.000 25.900 ;
        RECT 49.400 25.800 49.800 26.600 ;
        RECT 40.700 25.700 41.100 25.800 ;
        RECT 39.000 25.400 41.100 25.700 ;
        RECT 39.000 21.100 39.400 25.400 ;
        RECT 42.300 25.200 42.600 25.800 ;
        RECT 45.400 25.500 48.200 25.600 ;
        RECT 45.300 25.400 48.200 25.500 ;
        RECT 41.400 24.900 42.600 25.200 ;
        RECT 43.300 25.300 48.200 25.400 ;
        RECT 43.300 25.100 45.700 25.300 ;
        RECT 41.400 24.400 41.700 24.900 ;
        RECT 41.000 24.000 41.700 24.400 ;
        RECT 42.500 24.500 42.900 24.600 ;
        RECT 43.300 24.500 43.600 25.100 ;
        RECT 42.500 24.200 43.600 24.500 ;
        RECT 43.900 24.500 46.600 24.800 ;
        RECT 43.900 24.400 44.300 24.500 ;
        RECT 46.200 24.400 46.600 24.500 ;
        RECT 43.100 23.700 43.500 23.800 ;
        RECT 44.500 23.700 44.900 23.800 ;
        RECT 41.400 23.100 41.800 23.500 ;
        RECT 43.100 23.400 44.900 23.700 ;
        RECT 43.500 23.100 43.800 23.400 ;
        RECT 46.200 23.100 46.600 23.500 ;
        RECT 41.100 21.100 41.700 23.100 ;
        RECT 43.400 21.100 43.800 23.100 ;
        RECT 45.600 22.800 46.600 23.100 ;
        RECT 45.600 21.100 46.000 22.800 ;
        RECT 47.800 21.100 48.200 25.300 ;
        RECT 50.100 25.100 50.400 26.800 ;
        RECT 51.000 25.100 51.400 25.200 ;
        RECT 52.600 25.100 53.000 27.900 ;
        RECT 54.200 26.800 54.600 27.600 ;
        RECT 55.000 26.100 55.400 27.900 ;
        RECT 56.700 27.200 57.000 27.900 ;
        RECT 57.500 27.700 59.300 27.900 ;
        RECT 59.800 27.500 60.200 29.900 ;
        RECT 62.000 29.200 62.400 29.900 ;
        RECT 61.400 28.900 62.400 29.200 ;
        RECT 64.200 28.900 64.600 29.900 ;
        RECT 66.300 29.200 66.900 29.900 ;
        RECT 66.200 28.900 66.900 29.200 ;
        RECT 61.400 28.500 61.800 28.900 ;
        RECT 64.200 28.600 64.500 28.900 ;
        RECT 62.200 28.200 62.600 28.600 ;
        RECT 63.100 28.300 64.500 28.600 ;
        RECT 66.200 28.500 66.600 28.900 ;
        RECT 63.100 28.200 63.500 28.300 ;
        RECT 58.600 27.200 59.000 27.400 ;
        RECT 56.600 26.800 57.900 27.200 ;
        RECT 58.600 26.900 59.400 27.200 ;
        RECT 59.000 26.800 59.400 26.900 ;
        RECT 60.200 27.100 61.000 27.200 ;
        RECT 62.300 27.100 62.600 28.200 ;
        RECT 67.100 27.700 67.500 27.800 ;
        RECT 68.600 27.700 69.000 29.900 ;
        RECT 67.100 27.400 69.000 27.700 ;
        RECT 65.100 27.100 65.500 27.200 ;
        RECT 60.200 26.800 65.700 27.100 ;
        RECT 57.600 26.200 57.900 26.800 ;
        RECT 61.700 26.700 62.100 26.800 ;
        RECT 55.000 25.800 56.900 26.100 ;
        RECT 57.400 25.800 57.900 26.200 ;
        RECT 58.200 25.800 58.600 26.600 ;
        RECT 60.900 26.200 61.300 26.300 ;
        RECT 60.900 26.100 63.400 26.200 ;
        RECT 63.800 26.100 64.200 26.200 ;
        RECT 60.900 25.900 64.200 26.100 ;
        RECT 63.000 25.800 64.200 25.900 ;
        RECT 49.900 24.800 50.400 25.100 ;
        RECT 50.700 24.800 53.000 25.100 ;
        RECT 49.900 21.100 50.300 24.800 ;
        RECT 50.700 24.200 51.000 24.800 ;
        RECT 50.600 23.800 51.000 24.200 ;
        RECT 52.600 21.100 53.000 24.800 ;
        RECT 53.400 24.400 53.800 25.200 ;
        RECT 55.000 21.100 55.400 25.800 ;
        RECT 56.600 25.200 56.900 25.800 ;
        RECT 55.800 24.400 56.200 25.200 ;
        RECT 56.600 25.100 57.000 25.200 ;
        RECT 57.600 25.100 57.900 25.800 ;
        RECT 59.800 25.500 62.600 25.600 ;
        RECT 59.800 25.400 62.700 25.500 ;
        RECT 59.800 25.300 64.700 25.400 ;
        RECT 56.600 24.800 57.300 25.100 ;
        RECT 57.600 24.800 58.100 25.100 ;
        RECT 57.000 24.200 57.300 24.800 ;
        RECT 57.000 23.800 57.400 24.200 ;
        RECT 57.700 21.100 58.100 24.800 ;
        RECT 59.800 21.100 60.200 25.300 ;
        RECT 62.300 25.100 64.700 25.300 ;
        RECT 61.400 24.500 64.100 24.800 ;
        RECT 61.400 24.400 61.800 24.500 ;
        RECT 63.700 24.400 64.100 24.500 ;
        RECT 64.400 24.500 64.700 25.100 ;
        RECT 65.400 25.200 65.700 26.800 ;
        RECT 66.200 26.400 66.600 26.500 ;
        RECT 66.200 26.100 68.100 26.400 ;
        RECT 67.700 26.000 68.100 26.100 ;
        RECT 66.900 25.700 67.300 25.800 ;
        RECT 68.600 25.700 69.000 27.400 ;
        RECT 66.900 25.400 69.000 25.700 ;
        RECT 65.400 24.900 66.600 25.200 ;
        RECT 65.100 24.500 65.500 24.600 ;
        RECT 64.400 24.200 65.500 24.500 ;
        RECT 66.300 24.400 66.600 24.900 ;
        RECT 66.300 24.000 67.000 24.400 ;
        RECT 63.100 23.700 63.500 23.800 ;
        RECT 64.500 23.700 64.900 23.800 ;
        RECT 61.400 23.100 61.800 23.500 ;
        RECT 63.100 23.400 64.900 23.700 ;
        RECT 64.200 23.100 64.500 23.400 ;
        RECT 66.200 23.100 66.600 23.500 ;
        RECT 61.400 22.800 62.400 23.100 ;
        RECT 62.000 21.100 62.400 22.800 ;
        RECT 64.200 21.100 64.600 23.100 ;
        RECT 66.300 21.100 66.900 23.100 ;
        RECT 68.600 21.100 69.000 25.400 ;
        RECT 69.400 27.700 69.800 29.900 ;
        RECT 71.500 29.200 72.100 29.900 ;
        RECT 71.500 28.900 72.200 29.200 ;
        RECT 73.800 28.900 74.200 29.900 ;
        RECT 76.000 29.200 76.400 29.900 ;
        RECT 76.000 28.900 77.000 29.200 ;
        RECT 71.800 28.500 72.200 28.900 ;
        RECT 73.900 28.600 74.200 28.900 ;
        RECT 73.900 28.300 75.300 28.600 ;
        RECT 74.900 28.200 75.300 28.300 ;
        RECT 75.800 28.200 76.200 28.600 ;
        RECT 76.600 28.500 77.000 28.900 ;
        RECT 70.900 27.700 71.300 27.800 ;
        RECT 69.400 27.400 71.300 27.700 ;
        RECT 69.400 25.700 69.800 27.400 ;
        RECT 72.900 27.100 73.300 27.200 ;
        RECT 75.800 27.100 76.100 28.200 ;
        RECT 78.200 27.500 78.600 29.900 ;
        RECT 80.300 28.200 80.700 29.900 ;
        RECT 79.800 27.900 80.700 28.200 ;
        RECT 81.400 27.900 81.800 29.900 ;
        RECT 82.200 28.000 82.600 29.900 ;
        RECT 83.800 28.000 84.200 29.900 ;
        RECT 82.200 27.900 84.200 28.000 ;
        RECT 77.400 27.100 78.200 27.200 ;
        RECT 72.700 26.800 78.200 27.100 ;
        RECT 79.000 26.800 79.400 27.600 ;
        RECT 71.800 26.400 72.200 26.500 ;
        RECT 70.300 26.100 72.200 26.400 ;
        RECT 72.700 26.200 73.000 26.800 ;
        RECT 76.300 26.700 76.700 26.800 ;
        RECT 75.800 26.200 76.200 26.300 ;
        RECT 77.100 26.200 77.500 26.300 ;
        RECT 70.300 26.000 70.700 26.100 ;
        RECT 72.600 25.800 73.000 26.200 ;
        RECT 75.000 25.900 77.500 26.200 ;
        RECT 79.800 26.100 80.200 27.900 ;
        RECT 81.500 27.200 81.800 27.900 ;
        RECT 82.300 27.700 84.100 27.900 ;
        RECT 86.200 27.700 86.600 29.900 ;
        RECT 88.300 29.200 88.900 29.900 ;
        RECT 88.300 28.900 89.000 29.200 ;
        RECT 90.600 28.900 91.000 29.900 ;
        RECT 92.800 29.200 93.200 29.900 ;
        RECT 92.800 28.900 93.800 29.200 ;
        RECT 88.600 28.500 89.000 28.900 ;
        RECT 90.700 28.600 91.000 28.900 ;
        RECT 90.700 28.300 92.100 28.600 ;
        RECT 91.700 28.200 92.100 28.300 ;
        RECT 92.600 28.200 93.000 28.600 ;
        RECT 93.400 28.500 93.800 28.900 ;
        RECT 87.700 27.700 88.100 27.800 ;
        RECT 86.200 27.400 88.100 27.700 ;
        RECT 83.400 27.200 83.800 27.400 ;
        RECT 80.600 27.100 81.000 27.200 ;
        RECT 81.400 27.100 82.700 27.200 ;
        RECT 80.600 26.800 82.700 27.100 ;
        RECT 83.400 26.900 84.200 27.200 ;
        RECT 83.800 26.800 84.200 26.900 ;
        RECT 75.000 25.800 75.400 25.900 ;
        RECT 79.800 25.800 81.700 26.100 ;
        RECT 71.100 25.700 71.500 25.800 ;
        RECT 69.400 25.400 71.500 25.700 ;
        RECT 69.400 21.100 69.800 25.400 ;
        RECT 72.700 25.200 73.000 25.800 ;
        RECT 75.800 25.500 78.600 25.600 ;
        RECT 75.700 25.400 78.600 25.500 ;
        RECT 71.800 24.900 73.000 25.200 ;
        RECT 73.700 25.300 78.600 25.400 ;
        RECT 73.700 25.100 76.100 25.300 ;
        RECT 71.800 24.400 72.100 24.900 ;
        RECT 71.400 24.000 72.100 24.400 ;
        RECT 72.900 24.500 73.300 24.600 ;
        RECT 73.700 24.500 74.000 25.100 ;
        RECT 72.900 24.200 74.000 24.500 ;
        RECT 74.300 24.500 77.000 24.800 ;
        RECT 74.300 24.400 74.700 24.500 ;
        RECT 76.600 24.400 77.000 24.500 ;
        RECT 73.500 23.700 73.900 23.800 ;
        RECT 74.900 23.700 75.300 23.800 ;
        RECT 71.800 23.100 72.200 23.500 ;
        RECT 73.500 23.400 75.300 23.700 ;
        RECT 73.900 23.100 74.200 23.400 ;
        RECT 76.600 23.100 77.000 23.500 ;
        RECT 71.500 21.100 72.100 23.100 ;
        RECT 73.800 21.100 74.200 23.100 ;
        RECT 76.000 22.800 77.000 23.100 ;
        RECT 76.000 21.100 76.400 22.800 ;
        RECT 78.200 21.100 78.600 25.300 ;
        RECT 79.800 21.100 80.200 25.800 ;
        RECT 81.400 25.200 81.700 25.800 ;
        RECT 80.600 24.400 81.000 25.200 ;
        RECT 81.400 25.100 81.800 25.200 ;
        RECT 82.400 25.100 82.700 26.800 ;
        RECT 83.000 26.100 83.400 26.600 ;
        RECT 84.600 26.100 85.000 26.200 ;
        RECT 83.000 25.800 85.000 26.100 ;
        RECT 86.200 25.700 86.600 27.400 ;
        RECT 89.700 27.100 90.100 27.200 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 92.600 27.100 92.900 28.200 ;
        RECT 95.000 27.500 95.400 29.900 ;
        RECT 97.100 29.200 97.500 29.900 ;
        RECT 99.500 29.200 99.900 29.900 ;
        RECT 100.900 29.200 101.300 29.900 ;
        RECT 97.100 28.800 97.800 29.200 ;
        RECT 99.500 28.800 100.200 29.200 ;
        RECT 100.600 28.800 101.300 29.200 ;
        RECT 97.100 28.200 97.500 28.800 ;
        RECT 99.500 28.200 99.900 28.800 ;
        RECT 96.600 27.900 97.500 28.200 ;
        RECT 99.000 27.900 99.900 28.200 ;
        RECT 100.900 28.200 101.300 28.800 ;
        RECT 100.900 27.900 101.800 28.200 ;
        RECT 103.000 28.000 103.400 29.900 ;
        RECT 104.600 28.000 105.000 29.900 ;
        RECT 103.000 27.900 105.000 28.000 ;
        RECT 105.400 27.900 105.800 29.900 ;
        RECT 94.200 27.100 95.000 27.200 ;
        RECT 89.500 26.800 95.000 27.100 ;
        RECT 95.800 26.800 96.200 27.600 ;
        RECT 88.600 26.400 89.000 26.500 ;
        RECT 87.100 26.100 89.000 26.400 ;
        RECT 89.500 26.200 89.800 26.800 ;
        RECT 93.100 26.700 93.500 26.800 ;
        RECT 93.900 26.200 94.300 26.300 ;
        RECT 87.100 26.000 87.500 26.100 ;
        RECT 89.400 25.800 89.800 26.200 ;
        RECT 91.000 26.100 91.400 26.200 ;
        RECT 91.800 26.100 94.300 26.200 ;
        RECT 91.000 25.900 94.300 26.100 ;
        RECT 91.000 25.800 92.200 25.900 ;
        RECT 87.900 25.700 88.300 25.800 ;
        RECT 86.200 25.400 88.300 25.700 ;
        RECT 81.400 24.800 82.100 25.100 ;
        RECT 82.400 24.800 82.900 25.100 ;
        RECT 81.800 24.200 82.100 24.800 ;
        RECT 81.800 23.800 82.200 24.200 ;
        RECT 82.500 21.100 82.900 24.800 ;
        RECT 86.200 21.100 86.600 25.400 ;
        RECT 89.500 25.200 89.800 25.800 ;
        RECT 92.600 25.500 95.400 25.600 ;
        RECT 92.500 25.400 95.400 25.500 ;
        RECT 88.600 24.900 89.800 25.200 ;
        RECT 90.500 25.300 95.400 25.400 ;
        RECT 90.500 25.100 92.900 25.300 ;
        RECT 88.600 24.400 88.900 24.900 ;
        RECT 88.200 24.000 88.900 24.400 ;
        RECT 89.700 24.500 90.100 24.600 ;
        RECT 90.500 24.500 90.800 25.100 ;
        RECT 89.700 24.200 90.800 24.500 ;
        RECT 91.100 24.500 93.800 24.800 ;
        RECT 91.100 24.400 91.500 24.500 ;
        RECT 93.400 24.400 93.800 24.500 ;
        RECT 90.300 23.700 90.700 23.800 ;
        RECT 91.700 23.700 92.100 23.800 ;
        RECT 88.600 23.100 89.000 23.500 ;
        RECT 90.300 23.400 92.100 23.700 ;
        RECT 90.700 23.100 91.000 23.400 ;
        RECT 93.400 23.100 93.800 23.500 ;
        RECT 88.300 21.100 88.900 23.100 ;
        RECT 90.600 21.100 91.000 23.100 ;
        RECT 92.800 22.800 93.800 23.100 ;
        RECT 92.800 21.100 93.200 22.800 ;
        RECT 95.000 21.100 95.400 25.300 ;
        RECT 96.600 21.100 97.000 27.900 ;
        RECT 97.400 27.100 97.800 27.200 ;
        RECT 98.200 27.100 98.600 27.600 ;
        RECT 97.400 26.800 98.600 27.100 ;
        RECT 97.400 24.400 97.800 25.200 ;
        RECT 99.000 21.100 99.400 27.900 ;
        RECT 99.800 25.100 100.200 25.200 ;
        RECT 100.600 25.100 101.000 25.200 ;
        RECT 99.800 24.800 101.000 25.100 ;
        RECT 99.800 24.400 100.200 24.800 ;
        RECT 100.600 24.400 101.000 24.800 ;
        RECT 101.400 21.100 101.800 27.900 ;
        RECT 103.100 27.700 104.900 27.900 ;
        RECT 102.200 26.800 102.600 27.600 ;
        RECT 103.400 27.200 103.800 27.400 ;
        RECT 105.400 27.200 105.700 27.900 ;
        RECT 106.200 27.500 106.600 29.900 ;
        RECT 108.400 29.200 108.800 29.900 ;
        RECT 107.800 28.900 108.800 29.200 ;
        RECT 110.600 28.900 111.000 29.900 ;
        RECT 112.700 29.200 113.300 29.900 ;
        RECT 112.600 28.900 113.300 29.200 ;
        RECT 107.800 28.500 108.200 28.900 ;
        RECT 110.600 28.600 110.900 28.900 ;
        RECT 108.600 28.200 109.000 28.600 ;
        RECT 109.500 28.300 110.900 28.600 ;
        RECT 112.600 28.500 113.000 28.900 ;
        RECT 109.500 28.200 109.900 28.300 ;
        RECT 103.000 26.900 103.800 27.200 ;
        RECT 103.000 26.800 103.400 26.900 ;
        RECT 104.500 26.800 105.800 27.200 ;
        RECT 106.600 27.100 107.400 27.200 ;
        RECT 108.700 27.100 109.000 28.200 ;
        RECT 113.500 27.700 113.900 27.800 ;
        RECT 115.000 27.700 115.400 29.900 ;
        RECT 113.500 27.400 115.400 27.700 ;
        RECT 111.500 27.100 111.900 27.200 ;
        RECT 106.600 26.800 112.100 27.100 ;
        RECT 103.800 25.800 104.200 26.600 ;
        RECT 104.500 26.200 104.800 26.800 ;
        RECT 108.100 26.700 108.500 26.800 ;
        RECT 107.300 26.200 107.700 26.300 ;
        RECT 108.600 26.200 109.000 26.300 ;
        RECT 111.800 26.200 112.100 26.800 ;
        RECT 112.600 26.400 113.000 26.500 ;
        RECT 104.500 25.800 105.000 26.200 ;
        RECT 107.300 25.900 109.800 26.200 ;
        RECT 109.400 25.800 109.800 25.900 ;
        RECT 111.800 25.800 112.200 26.200 ;
        RECT 112.600 26.100 114.500 26.400 ;
        RECT 114.100 26.000 114.500 26.100 ;
        RECT 104.500 25.100 104.800 25.800 ;
        RECT 106.200 25.500 109.000 25.600 ;
        RECT 106.200 25.400 109.100 25.500 ;
        RECT 106.200 25.300 111.100 25.400 ;
        RECT 105.400 25.100 105.800 25.200 ;
        RECT 104.300 24.800 104.800 25.100 ;
        RECT 105.100 24.800 105.800 25.100 ;
        RECT 104.300 21.100 104.700 24.800 ;
        RECT 105.100 24.200 105.400 24.800 ;
        RECT 105.000 23.800 105.400 24.200 ;
        RECT 106.200 21.100 106.600 25.300 ;
        RECT 108.700 25.100 111.100 25.300 ;
        RECT 107.800 24.500 110.500 24.800 ;
        RECT 107.800 24.400 108.200 24.500 ;
        RECT 110.100 24.400 110.500 24.500 ;
        RECT 110.800 24.500 111.100 25.100 ;
        RECT 111.800 25.200 112.100 25.800 ;
        RECT 113.300 25.700 113.700 25.800 ;
        RECT 115.000 25.700 115.400 27.400 ;
        RECT 113.300 25.400 115.400 25.700 ;
        RECT 111.800 24.900 113.000 25.200 ;
        RECT 111.500 24.500 111.900 24.600 ;
        RECT 110.800 24.200 111.900 24.500 ;
        RECT 112.700 24.400 113.000 24.900 ;
        RECT 112.700 24.000 113.400 24.400 ;
        RECT 109.500 23.700 109.900 23.800 ;
        RECT 110.900 23.700 111.300 23.800 ;
        RECT 107.800 23.100 108.200 23.500 ;
        RECT 109.500 23.400 111.300 23.700 ;
        RECT 110.600 23.100 110.900 23.400 ;
        RECT 112.600 23.100 113.000 23.500 ;
        RECT 107.800 22.800 108.800 23.100 ;
        RECT 108.400 21.100 108.800 22.800 ;
        RECT 110.600 21.100 111.000 23.100 ;
        RECT 112.700 21.100 113.300 23.100 ;
        RECT 115.000 21.100 115.400 25.400 ;
        RECT 115.800 27.700 116.200 29.900 ;
        RECT 117.900 29.200 118.500 29.900 ;
        RECT 117.900 28.900 118.600 29.200 ;
        RECT 120.200 28.900 120.600 29.900 ;
        RECT 122.400 29.200 122.800 29.900 ;
        RECT 122.400 28.900 123.400 29.200 ;
        RECT 118.200 28.500 118.600 28.900 ;
        RECT 120.300 28.600 120.600 28.900 ;
        RECT 120.300 28.300 121.700 28.600 ;
        RECT 121.300 28.200 121.700 28.300 ;
        RECT 122.200 28.200 122.600 28.600 ;
        RECT 123.000 28.500 123.400 28.900 ;
        RECT 117.300 27.700 117.700 27.800 ;
        RECT 115.800 27.400 117.700 27.700 ;
        RECT 115.800 25.700 116.200 27.400 ;
        RECT 122.200 27.200 122.500 28.200 ;
        RECT 124.600 27.500 125.000 29.900 ;
        RECT 125.700 29.200 126.100 29.900 ;
        RECT 125.400 28.800 126.100 29.200 ;
        RECT 125.700 28.200 126.100 28.800 ;
        RECT 125.700 27.900 126.600 28.200 ;
        RECT 119.300 27.100 119.700 27.200 ;
        RECT 122.200 27.100 122.600 27.200 ;
        RECT 123.800 27.100 124.600 27.200 ;
        RECT 119.100 26.800 124.600 27.100 ;
        RECT 118.200 26.400 118.600 26.500 ;
        RECT 116.700 26.100 118.600 26.400 ;
        RECT 116.700 26.000 117.100 26.100 ;
        RECT 117.500 25.700 117.900 25.800 ;
        RECT 115.800 25.400 117.900 25.700 ;
        RECT 115.800 21.100 116.200 25.400 ;
        RECT 119.100 25.200 119.400 26.800 ;
        RECT 122.700 26.700 123.100 26.800 ;
        RECT 123.500 26.200 123.900 26.300 ;
        RECT 121.400 25.900 123.900 26.200 ;
        RECT 121.400 25.800 121.800 25.900 ;
        RECT 122.200 25.500 125.000 25.600 ;
        RECT 122.100 25.400 125.000 25.500 ;
        RECT 118.200 24.900 119.400 25.200 ;
        RECT 120.100 25.300 125.000 25.400 ;
        RECT 120.100 25.100 122.500 25.300 ;
        RECT 118.200 24.400 118.500 24.900 ;
        RECT 117.800 24.000 118.500 24.400 ;
        RECT 119.300 24.500 119.700 24.600 ;
        RECT 120.100 24.500 120.400 25.100 ;
        RECT 119.300 24.200 120.400 24.500 ;
        RECT 120.700 24.500 123.400 24.800 ;
        RECT 120.700 24.400 121.100 24.500 ;
        RECT 123.000 24.400 123.400 24.500 ;
        RECT 119.900 23.700 120.300 23.800 ;
        RECT 121.300 23.700 121.700 23.800 ;
        RECT 118.200 23.100 118.600 23.500 ;
        RECT 119.900 23.400 121.700 23.700 ;
        RECT 120.300 23.100 120.600 23.400 ;
        RECT 123.000 23.100 123.400 23.500 ;
        RECT 117.900 21.100 118.500 23.100 ;
        RECT 120.200 21.100 120.600 23.100 ;
        RECT 122.400 22.800 123.400 23.100 ;
        RECT 122.400 21.100 122.800 22.800 ;
        RECT 124.600 21.100 125.000 25.300 ;
        RECT 125.400 24.400 125.800 25.200 ;
        RECT 126.200 21.100 126.600 27.900 ;
        RECT 128.600 27.600 129.000 29.900 ;
        RECT 130.200 27.600 130.600 29.900 ;
        RECT 131.800 27.600 132.200 29.900 ;
        RECT 133.400 27.600 133.800 29.900 ;
        RECT 135.800 27.600 136.200 29.900 ;
        RECT 137.400 27.600 137.800 29.900 ;
        RECT 139.000 27.600 139.400 29.900 ;
        RECT 140.600 27.600 141.000 29.900 ;
        RECT 145.100 28.200 145.500 29.900 ;
        RECT 144.600 27.900 145.500 28.200 ;
        RECT 146.200 27.900 146.600 29.900 ;
        RECT 147.000 28.000 147.400 29.900 ;
        RECT 148.600 28.000 149.000 29.900 ;
        RECT 147.000 27.900 149.000 28.000 ;
        RECT 127.000 26.800 127.400 27.600 ;
        RECT 128.600 27.200 129.500 27.600 ;
        RECT 130.200 27.200 131.300 27.600 ;
        RECT 131.800 27.200 132.900 27.600 ;
        RECT 133.400 27.200 134.600 27.600 ;
        RECT 135.800 27.200 136.700 27.600 ;
        RECT 137.400 27.200 138.500 27.600 ;
        RECT 139.000 27.200 140.100 27.600 ;
        RECT 140.600 27.200 141.800 27.600 ;
        RECT 129.100 26.900 129.500 27.200 ;
        RECT 130.900 26.900 131.300 27.200 ;
        RECT 132.500 26.900 132.900 27.200 ;
        RECT 129.100 26.500 130.400 26.900 ;
        RECT 130.900 26.500 132.100 26.900 ;
        RECT 132.500 26.500 133.800 26.900 ;
        RECT 129.100 25.800 129.500 26.500 ;
        RECT 130.900 25.800 131.300 26.500 ;
        RECT 132.500 25.800 132.900 26.500 ;
        RECT 134.200 25.800 134.600 27.200 ;
        RECT 136.300 26.900 136.700 27.200 ;
        RECT 138.100 26.900 138.500 27.200 ;
        RECT 139.700 26.900 140.100 27.200 ;
        RECT 136.300 26.500 137.600 26.900 ;
        RECT 138.100 26.500 139.300 26.900 ;
        RECT 139.700 26.500 141.000 26.900 ;
        RECT 136.300 25.800 136.700 26.500 ;
        RECT 138.100 25.800 138.500 26.500 ;
        RECT 139.700 25.800 140.100 26.500 ;
        RECT 141.400 25.800 141.800 27.200 ;
        RECT 143.800 26.800 144.200 27.600 ;
        RECT 128.600 25.400 129.500 25.800 ;
        RECT 130.200 25.400 131.300 25.800 ;
        RECT 131.800 25.400 132.900 25.800 ;
        RECT 133.400 25.400 134.600 25.800 ;
        RECT 135.800 25.400 136.700 25.800 ;
        RECT 137.400 25.400 138.500 25.800 ;
        RECT 139.000 25.400 140.100 25.800 ;
        RECT 140.600 25.400 141.800 25.800 ;
        RECT 144.600 26.100 145.000 27.900 ;
        RECT 146.300 27.200 146.600 27.900 ;
        RECT 147.100 27.700 148.900 27.900 ;
        RECT 149.400 27.700 149.800 29.900 ;
        RECT 151.500 29.200 152.100 29.900 ;
        RECT 151.500 28.900 152.200 29.200 ;
        RECT 153.800 28.900 154.200 29.900 ;
        RECT 156.000 29.200 156.400 29.900 ;
        RECT 156.000 28.900 157.000 29.200 ;
        RECT 151.800 28.500 152.200 28.900 ;
        RECT 153.900 28.600 154.200 28.900 ;
        RECT 153.900 28.300 155.300 28.600 ;
        RECT 154.900 28.200 155.300 28.300 ;
        RECT 155.800 28.200 156.200 28.600 ;
        RECT 156.600 28.500 157.000 28.900 ;
        RECT 150.900 27.700 151.300 27.800 ;
        RECT 149.400 27.400 151.300 27.700 ;
        RECT 148.200 27.200 148.600 27.400 ;
        RECT 146.200 26.800 147.500 27.200 ;
        RECT 148.200 26.900 149.000 27.200 ;
        RECT 148.600 26.800 149.000 26.900 ;
        RECT 144.600 25.800 146.500 26.100 ;
        RECT 128.600 21.100 129.000 25.400 ;
        RECT 130.200 21.100 130.600 25.400 ;
        RECT 131.800 21.100 132.200 25.400 ;
        RECT 133.400 21.100 133.800 25.400 ;
        RECT 135.800 21.100 136.200 25.400 ;
        RECT 137.400 21.100 137.800 25.400 ;
        RECT 139.000 21.100 139.400 25.400 ;
        RECT 140.600 21.100 141.000 25.400 ;
        RECT 144.600 21.100 145.000 25.800 ;
        RECT 146.200 25.200 146.500 25.800 ;
        RECT 147.200 25.200 147.500 26.800 ;
        RECT 147.800 25.800 148.200 26.600 ;
        RECT 149.400 25.700 149.800 27.400 ;
        RECT 152.900 27.100 153.300 27.200 ;
        RECT 155.800 27.100 156.100 28.200 ;
        RECT 158.200 27.500 158.600 29.900 ;
        RECT 159.000 28.000 159.400 29.900 ;
        RECT 160.600 28.000 161.000 29.900 ;
        RECT 159.000 27.900 161.000 28.000 ;
        RECT 161.400 27.900 161.800 29.900 ;
        RECT 162.200 28.000 162.600 29.900 ;
        RECT 163.800 28.000 164.200 29.900 ;
        RECT 162.200 27.900 164.200 28.000 ;
        RECT 164.600 27.900 165.000 29.900 ;
        RECT 165.700 28.200 166.100 29.900 ;
        RECT 165.700 27.900 166.600 28.200 ;
        RECT 159.100 27.700 160.900 27.900 ;
        RECT 159.400 27.200 159.800 27.400 ;
        RECT 161.400 27.200 161.700 27.900 ;
        RECT 162.300 27.700 164.100 27.900 ;
        RECT 162.600 27.200 163.000 27.400 ;
        RECT 164.600 27.200 164.900 27.900 ;
        RECT 157.400 27.100 158.200 27.200 ;
        RECT 152.700 26.800 158.200 27.100 ;
        RECT 159.000 26.900 159.800 27.200 ;
        RECT 159.000 26.800 159.400 26.900 ;
        RECT 160.500 26.800 161.800 27.200 ;
        RECT 162.200 26.900 163.000 27.200 ;
        RECT 162.200 26.800 162.600 26.900 ;
        RECT 163.700 26.800 165.000 27.200 ;
        RECT 151.800 26.400 152.200 26.500 ;
        RECT 150.300 26.100 152.200 26.400 ;
        RECT 152.700 26.100 153.000 26.800 ;
        RECT 156.300 26.700 156.700 26.800 ;
        RECT 157.100 26.200 157.500 26.300 ;
        RECT 153.400 26.100 153.800 26.200 ;
        RECT 150.300 26.000 150.700 26.100 ;
        RECT 152.600 25.800 153.800 26.100 ;
        RECT 155.000 25.900 157.500 26.200 ;
        RECT 155.000 25.800 155.400 25.900 ;
        RECT 159.800 25.800 160.200 26.600 ;
        RECT 151.100 25.700 151.500 25.800 ;
        RECT 149.400 25.400 151.500 25.700 ;
        RECT 145.400 24.400 145.800 25.200 ;
        RECT 146.200 25.100 146.600 25.200 ;
        RECT 146.200 24.800 146.900 25.100 ;
        RECT 147.200 24.800 148.200 25.200 ;
        RECT 146.600 24.200 146.900 24.800 ;
        RECT 146.600 23.800 147.000 24.200 ;
        RECT 147.300 21.100 147.700 24.800 ;
        RECT 149.400 21.100 149.800 25.400 ;
        RECT 152.700 25.200 153.000 25.800 ;
        RECT 155.800 25.500 158.600 25.600 ;
        RECT 155.700 25.400 158.600 25.500 ;
        RECT 151.800 24.900 153.000 25.200 ;
        RECT 153.700 25.300 158.600 25.400 ;
        RECT 153.700 25.100 156.100 25.300 ;
        RECT 151.800 24.400 152.100 24.900 ;
        RECT 151.400 24.000 152.100 24.400 ;
        RECT 152.900 24.500 153.300 24.600 ;
        RECT 153.700 24.500 154.000 25.100 ;
        RECT 152.900 24.200 154.000 24.500 ;
        RECT 154.300 24.500 157.000 24.800 ;
        RECT 154.300 24.400 154.700 24.500 ;
        RECT 156.600 24.400 157.000 24.500 ;
        RECT 153.500 23.700 153.900 23.800 ;
        RECT 154.900 23.700 155.300 23.800 ;
        RECT 151.800 23.100 152.200 23.500 ;
        RECT 153.500 23.400 155.300 23.700 ;
        RECT 153.900 23.100 154.200 23.400 ;
        RECT 156.600 23.100 157.000 23.500 ;
        RECT 151.500 21.100 152.100 23.100 ;
        RECT 153.800 21.100 154.200 23.100 ;
        RECT 156.000 22.800 157.000 23.100 ;
        RECT 156.000 21.100 156.400 22.800 ;
        RECT 158.200 21.100 158.600 25.300 ;
        RECT 160.500 25.100 160.800 26.800 ;
        RECT 163.000 25.800 163.400 26.600 ;
        RECT 161.400 25.100 161.800 25.200 ;
        RECT 163.700 25.100 164.000 26.800 ;
        RECT 166.200 26.100 166.600 27.900 ;
        RECT 167.800 27.700 168.200 29.900 ;
        RECT 169.900 29.200 170.500 29.900 ;
        RECT 169.900 28.900 170.600 29.200 ;
        RECT 172.200 28.900 172.600 29.900 ;
        RECT 174.400 29.200 174.800 29.900 ;
        RECT 174.400 28.900 175.400 29.200 ;
        RECT 170.200 28.500 170.600 28.900 ;
        RECT 172.300 28.600 172.600 28.900 ;
        RECT 172.300 28.300 173.700 28.600 ;
        RECT 173.300 28.200 173.700 28.300 ;
        RECT 174.200 28.200 174.600 28.600 ;
        RECT 175.000 28.500 175.400 28.900 ;
        RECT 169.300 27.700 169.700 27.800 ;
        RECT 167.000 26.800 167.400 27.600 ;
        RECT 167.800 27.400 169.700 27.700 ;
        RECT 164.600 25.800 166.600 26.100 ;
        RECT 164.600 25.200 164.900 25.800 ;
        RECT 164.600 25.100 165.000 25.200 ;
        RECT 160.300 24.800 160.800 25.100 ;
        RECT 161.100 24.800 161.800 25.100 ;
        RECT 163.500 24.800 164.000 25.100 ;
        RECT 164.300 24.800 165.000 25.100 ;
        RECT 160.300 21.100 160.700 24.800 ;
        RECT 161.100 24.200 161.400 24.800 ;
        RECT 161.000 23.800 161.400 24.200 ;
        RECT 163.500 21.100 163.900 24.800 ;
        RECT 164.300 24.200 164.600 24.800 ;
        RECT 165.400 24.400 165.800 25.200 ;
        RECT 164.200 23.800 164.600 24.200 ;
        RECT 166.200 21.100 166.600 25.800 ;
        RECT 167.800 25.700 168.200 27.400 ;
        RECT 171.300 27.100 171.700 27.200 ;
        RECT 174.200 27.100 174.500 28.200 ;
        RECT 176.600 27.500 177.000 29.900 ;
        RECT 177.400 27.700 177.800 29.900 ;
        RECT 179.500 29.200 180.100 29.900 ;
        RECT 179.500 28.900 180.200 29.200 ;
        RECT 181.800 28.900 182.200 29.900 ;
        RECT 184.000 29.200 184.400 29.900 ;
        RECT 184.000 28.900 185.000 29.200 ;
        RECT 179.800 28.500 180.200 28.900 ;
        RECT 181.900 28.600 182.200 28.900 ;
        RECT 181.900 28.300 183.300 28.600 ;
        RECT 182.900 28.200 183.300 28.300 ;
        RECT 183.800 28.200 184.200 28.600 ;
        RECT 184.600 28.500 185.000 28.900 ;
        RECT 178.900 27.700 179.300 27.800 ;
        RECT 177.400 27.400 179.300 27.700 ;
        RECT 175.800 27.100 176.600 27.200 ;
        RECT 171.100 26.800 176.600 27.100 ;
        RECT 170.200 26.400 170.600 26.500 ;
        RECT 168.700 26.100 170.600 26.400 ;
        RECT 171.100 26.200 171.400 26.800 ;
        RECT 174.700 26.700 175.100 26.800 ;
        RECT 175.500 26.200 175.900 26.300 ;
        RECT 168.700 26.000 169.100 26.100 ;
        RECT 171.000 25.800 171.400 26.200 ;
        RECT 172.600 26.100 173.000 26.200 ;
        RECT 173.400 26.100 175.900 26.200 ;
        RECT 172.600 25.900 175.900 26.100 ;
        RECT 172.600 25.800 173.800 25.900 ;
        RECT 169.500 25.700 169.900 25.800 ;
        RECT 167.800 25.400 169.900 25.700 ;
        RECT 167.800 21.100 168.200 25.400 ;
        RECT 171.100 25.200 171.400 25.800 ;
        RECT 177.400 25.700 177.800 27.400 ;
        RECT 180.900 27.100 181.300 27.200 ;
        RECT 183.800 27.100 184.100 28.200 ;
        RECT 186.200 27.500 186.600 29.900 ;
        RECT 188.600 27.500 189.000 29.900 ;
        RECT 190.800 29.200 191.200 29.900 ;
        RECT 190.200 28.900 191.200 29.200 ;
        RECT 193.000 28.900 193.400 29.900 ;
        RECT 195.100 29.200 195.700 29.900 ;
        RECT 195.000 28.900 195.700 29.200 ;
        RECT 190.200 28.500 190.600 28.900 ;
        RECT 193.000 28.600 193.300 28.900 ;
        RECT 191.000 28.200 191.400 28.600 ;
        RECT 191.900 28.300 193.300 28.600 ;
        RECT 195.000 28.500 195.400 28.900 ;
        RECT 191.900 28.200 192.300 28.300 ;
        RECT 185.400 27.100 186.200 27.200 ;
        RECT 189.000 27.100 189.800 27.200 ;
        RECT 191.100 27.100 191.400 28.200 ;
        RECT 195.900 27.700 196.300 27.800 ;
        RECT 197.400 27.700 197.800 29.900 ;
        RECT 198.500 29.200 198.900 29.900 ;
        RECT 198.500 28.800 199.400 29.200 ;
        RECT 198.500 28.200 198.900 28.800 ;
        RECT 198.500 27.900 199.400 28.200 ;
        RECT 195.900 27.400 197.800 27.700 ;
        RECT 193.900 27.100 194.300 27.200 ;
        RECT 180.700 26.800 194.500 27.100 ;
        RECT 179.800 26.400 180.200 26.500 ;
        RECT 178.300 26.100 180.200 26.400 ;
        RECT 180.700 26.200 181.000 26.800 ;
        RECT 184.300 26.700 184.700 26.800 ;
        RECT 190.500 26.700 190.900 26.800 ;
        RECT 185.100 26.200 185.500 26.300 ;
        RECT 178.300 26.000 178.700 26.100 ;
        RECT 180.600 25.800 181.000 26.200 ;
        RECT 181.400 26.100 181.800 26.200 ;
        RECT 183.000 26.100 185.500 26.200 ;
        RECT 181.400 25.900 185.500 26.100 ;
        RECT 189.700 26.200 190.100 26.300 ;
        RECT 191.000 26.200 191.400 26.300 ;
        RECT 189.700 25.900 192.200 26.200 ;
        RECT 181.400 25.800 183.400 25.900 ;
        RECT 191.800 25.800 192.200 25.900 ;
        RECT 179.100 25.700 179.500 25.800 ;
        RECT 174.200 25.500 177.000 25.600 ;
        RECT 174.100 25.400 177.000 25.500 ;
        RECT 170.200 24.900 171.400 25.200 ;
        RECT 172.100 25.300 177.000 25.400 ;
        RECT 172.100 25.100 174.500 25.300 ;
        RECT 170.200 24.400 170.500 24.900 ;
        RECT 169.800 24.000 170.500 24.400 ;
        RECT 171.300 24.500 171.700 24.600 ;
        RECT 172.100 24.500 172.400 25.100 ;
        RECT 171.300 24.200 172.400 24.500 ;
        RECT 172.700 24.500 175.400 24.800 ;
        RECT 172.700 24.400 173.100 24.500 ;
        RECT 175.000 24.400 175.400 24.500 ;
        RECT 171.900 23.700 172.300 23.800 ;
        RECT 173.300 23.700 173.700 23.800 ;
        RECT 170.200 23.100 170.600 23.500 ;
        RECT 171.900 23.400 173.700 23.700 ;
        RECT 172.300 23.100 172.600 23.400 ;
        RECT 175.000 23.100 175.400 23.500 ;
        RECT 169.900 21.100 170.500 23.100 ;
        RECT 172.200 21.100 172.600 23.100 ;
        RECT 174.400 22.800 175.400 23.100 ;
        RECT 174.400 21.100 174.800 22.800 ;
        RECT 176.600 21.100 177.000 25.300 ;
        RECT 177.400 25.400 179.500 25.700 ;
        RECT 177.400 21.100 177.800 25.400 ;
        RECT 180.700 25.200 181.000 25.800 ;
        RECT 183.800 25.500 186.600 25.600 ;
        RECT 183.700 25.400 186.600 25.500 ;
        RECT 179.800 24.900 181.000 25.200 ;
        RECT 181.700 25.300 186.600 25.400 ;
        RECT 181.700 25.100 184.100 25.300 ;
        RECT 179.800 24.400 180.100 24.900 ;
        RECT 179.400 24.000 180.100 24.400 ;
        RECT 180.900 24.500 181.300 24.600 ;
        RECT 181.700 24.500 182.000 25.100 ;
        RECT 180.900 24.200 182.000 24.500 ;
        RECT 182.300 24.500 185.000 24.800 ;
        RECT 182.300 24.400 182.700 24.500 ;
        RECT 184.600 24.400 185.000 24.500 ;
        RECT 181.500 23.700 181.900 23.800 ;
        RECT 182.900 23.700 183.300 23.800 ;
        RECT 179.800 23.100 180.200 23.500 ;
        RECT 181.500 23.400 183.300 23.700 ;
        RECT 181.900 23.100 182.200 23.400 ;
        RECT 184.600 23.100 185.000 23.500 ;
        RECT 179.500 21.100 180.100 23.100 ;
        RECT 181.800 21.100 182.200 23.100 ;
        RECT 184.000 22.800 185.000 23.100 ;
        RECT 184.000 21.100 184.400 22.800 ;
        RECT 186.200 21.100 186.600 25.300 ;
        RECT 188.600 25.500 191.400 25.600 ;
        RECT 188.600 25.400 191.500 25.500 ;
        RECT 188.600 25.300 193.500 25.400 ;
        RECT 188.600 21.100 189.000 25.300 ;
        RECT 191.100 25.100 193.500 25.300 ;
        RECT 190.200 24.500 192.900 24.800 ;
        RECT 190.200 24.400 190.600 24.500 ;
        RECT 192.500 24.400 192.900 24.500 ;
        RECT 193.200 24.500 193.500 25.100 ;
        RECT 194.200 25.200 194.500 26.800 ;
        RECT 195.000 26.400 195.400 26.500 ;
        RECT 195.000 26.100 196.900 26.400 ;
        RECT 196.500 26.000 196.900 26.100 ;
        RECT 195.700 25.700 196.100 25.800 ;
        RECT 197.400 25.700 197.800 27.400 ;
        RECT 195.700 25.400 197.800 25.700 ;
        RECT 194.200 24.900 195.400 25.200 ;
        RECT 193.900 24.500 194.300 24.600 ;
        RECT 193.200 24.200 194.300 24.500 ;
        RECT 195.100 24.400 195.400 24.900 ;
        RECT 195.100 24.000 195.800 24.400 ;
        RECT 191.900 23.700 192.300 23.800 ;
        RECT 193.300 23.700 193.700 23.800 ;
        RECT 190.200 23.100 190.600 23.500 ;
        RECT 191.900 23.400 193.700 23.700 ;
        RECT 193.000 23.100 193.300 23.400 ;
        RECT 195.000 23.100 195.400 23.500 ;
        RECT 190.200 22.800 191.200 23.100 ;
        RECT 190.800 21.100 191.200 22.800 ;
        RECT 193.000 21.100 193.400 23.100 ;
        RECT 195.100 21.100 195.700 23.100 ;
        RECT 197.400 21.100 197.800 25.400 ;
        RECT 198.200 24.400 198.600 25.200 ;
        RECT 199.000 21.100 199.400 27.900 ;
        RECT 200.600 27.600 201.000 29.900 ;
        RECT 202.200 28.200 202.600 29.900 ;
        RECT 202.200 27.900 202.700 28.200 ;
        RECT 203.800 28.000 204.200 29.900 ;
        RECT 205.400 28.000 205.800 29.900 ;
        RECT 203.800 27.900 205.800 28.000 ;
        RECT 206.200 27.900 206.600 29.900 ;
        RECT 207.300 28.200 207.700 29.900 ;
        RECT 207.300 27.900 208.200 28.200 ;
        RECT 199.800 26.800 200.200 27.600 ;
        RECT 200.600 27.300 201.900 27.600 ;
        RECT 200.700 26.200 201.100 26.600 ;
        RECT 200.600 25.800 201.100 26.200 ;
        RECT 201.600 26.500 201.900 27.300 ;
        RECT 202.400 27.200 202.700 27.900 ;
        RECT 203.900 27.700 205.700 27.900 ;
        RECT 204.200 27.200 204.600 27.400 ;
        RECT 206.200 27.200 206.500 27.900 ;
        RECT 202.200 26.800 202.700 27.200 ;
        RECT 203.800 26.900 204.600 27.200 ;
        RECT 205.300 27.100 206.600 27.200 ;
        RECT 207.000 27.100 207.400 27.200 ;
        RECT 203.800 26.800 204.200 26.900 ;
        RECT 205.300 26.800 207.400 27.100 ;
        RECT 201.600 26.100 202.100 26.500 ;
        RECT 201.600 25.100 201.900 26.100 ;
        RECT 202.400 25.100 202.700 26.800 ;
        RECT 204.600 25.800 205.000 26.600 ;
        RECT 205.300 25.100 205.600 26.800 ;
        RECT 207.800 26.100 208.200 27.900 ;
        RECT 209.400 27.700 209.800 29.900 ;
        RECT 211.500 29.200 212.100 29.900 ;
        RECT 211.500 28.900 212.200 29.200 ;
        RECT 213.800 28.900 214.200 29.900 ;
        RECT 216.000 29.200 216.400 29.900 ;
        RECT 216.000 28.900 217.000 29.200 ;
        RECT 211.800 28.500 212.200 28.900 ;
        RECT 213.900 28.600 214.200 28.900 ;
        RECT 213.900 28.300 215.300 28.600 ;
        RECT 214.900 28.200 215.300 28.300 ;
        RECT 215.800 28.200 216.200 28.600 ;
        RECT 216.600 28.500 217.000 28.900 ;
        RECT 210.900 27.700 211.300 27.800 ;
        RECT 208.600 27.100 209.000 27.600 ;
        RECT 209.400 27.400 211.300 27.700 ;
        RECT 209.400 27.100 209.800 27.400 ;
        RECT 215.800 27.200 216.100 28.200 ;
        RECT 218.200 27.500 218.600 29.900 ;
        RECT 219.300 29.200 219.700 29.900 ;
        RECT 219.000 28.800 219.700 29.200 ;
        RECT 219.300 28.200 219.700 28.800 ;
        RECT 219.300 27.900 220.200 28.200 ;
        RECT 212.900 27.100 213.800 27.200 ;
        RECT 215.800 27.100 216.200 27.200 ;
        RECT 217.400 27.100 218.200 27.200 ;
        RECT 208.600 26.800 209.800 27.100 ;
        RECT 206.200 25.800 208.200 26.100 ;
        RECT 206.200 25.200 206.500 25.800 ;
        RECT 206.200 25.100 206.600 25.200 ;
        RECT 200.600 24.800 201.900 25.100 ;
        RECT 200.600 21.100 201.000 24.800 ;
        RECT 202.200 24.600 202.700 25.100 ;
        RECT 205.100 24.800 205.600 25.100 ;
        RECT 205.900 24.800 206.600 25.100 ;
        RECT 202.200 21.100 202.600 24.600 ;
        RECT 205.100 21.100 205.500 24.800 ;
        RECT 205.900 24.200 206.200 24.800 ;
        RECT 207.000 24.400 207.400 25.200 ;
        RECT 205.800 23.800 206.200 24.200 ;
        RECT 207.800 21.100 208.200 25.800 ;
        RECT 209.400 25.700 209.800 26.800 ;
        RECT 212.700 26.800 218.200 27.100 ;
        RECT 211.800 26.400 212.200 26.500 ;
        RECT 210.300 26.100 212.200 26.400 ;
        RECT 210.300 26.000 210.700 26.100 ;
        RECT 211.100 25.700 211.500 25.800 ;
        RECT 209.400 25.400 211.500 25.700 ;
        RECT 209.400 21.100 209.800 25.400 ;
        RECT 212.700 25.200 213.000 26.800 ;
        RECT 216.300 26.700 216.700 26.800 ;
        RECT 217.100 26.200 217.500 26.300 ;
        RECT 215.000 25.900 217.500 26.200 ;
        RECT 215.000 25.800 215.400 25.900 ;
        RECT 215.800 25.500 218.600 25.600 ;
        RECT 215.700 25.400 218.600 25.500 ;
        RECT 211.800 24.900 213.000 25.200 ;
        RECT 213.700 25.300 218.600 25.400 ;
        RECT 213.700 25.100 216.100 25.300 ;
        RECT 211.800 24.400 212.100 24.900 ;
        RECT 211.400 24.000 212.100 24.400 ;
        RECT 212.900 24.500 213.300 24.600 ;
        RECT 213.700 24.500 214.000 25.100 ;
        RECT 212.900 24.200 214.000 24.500 ;
        RECT 214.300 24.500 217.000 24.800 ;
        RECT 214.300 24.400 214.700 24.500 ;
        RECT 216.600 24.400 217.000 24.500 ;
        RECT 213.500 23.700 213.900 23.800 ;
        RECT 214.900 23.700 215.300 23.800 ;
        RECT 211.800 23.100 212.200 23.500 ;
        RECT 213.500 23.400 215.300 23.700 ;
        RECT 213.900 23.100 214.200 23.400 ;
        RECT 216.600 23.100 217.000 23.500 ;
        RECT 211.500 21.100 212.100 23.100 ;
        RECT 213.800 21.100 214.200 23.100 ;
        RECT 216.000 22.800 217.000 23.100 ;
        RECT 216.000 21.100 216.400 22.800 ;
        RECT 218.200 21.100 218.600 25.300 ;
        RECT 219.000 24.400 219.400 25.200 ;
        RECT 219.800 21.100 220.200 27.900 ;
        RECT 221.400 27.700 221.800 29.900 ;
        RECT 223.500 29.200 224.100 29.900 ;
        RECT 223.500 28.900 224.200 29.200 ;
        RECT 225.800 28.900 226.200 29.900 ;
        RECT 228.000 29.200 228.400 29.900 ;
        RECT 228.000 28.900 229.000 29.200 ;
        RECT 223.800 28.500 224.200 28.900 ;
        RECT 225.900 28.600 226.200 28.900 ;
        RECT 225.900 28.300 227.300 28.600 ;
        RECT 226.900 28.200 227.300 28.300 ;
        RECT 227.800 28.200 228.200 28.600 ;
        RECT 228.600 28.500 229.000 28.900 ;
        RECT 222.900 27.700 223.300 27.800 ;
        RECT 220.600 26.800 221.000 27.600 ;
        RECT 221.400 27.400 223.300 27.700 ;
        RECT 221.400 25.700 221.800 27.400 ;
        RECT 224.900 27.100 225.300 27.200 ;
        RECT 227.800 27.100 228.100 28.200 ;
        RECT 230.200 27.500 230.600 29.900 ;
        RECT 229.400 27.100 230.200 27.200 ;
        RECT 224.700 26.800 230.200 27.100 ;
        RECT 223.800 26.400 224.200 26.500 ;
        RECT 222.300 26.100 224.200 26.400 ;
        RECT 224.700 26.200 225.000 26.800 ;
        RECT 228.300 26.700 228.700 26.800 ;
        RECT 229.100 26.200 229.500 26.300 ;
        RECT 222.300 26.000 222.700 26.100 ;
        RECT 224.600 25.800 225.000 26.200 ;
        RECT 227.000 25.900 229.500 26.200 ;
        RECT 227.000 25.800 227.400 25.900 ;
        RECT 223.100 25.700 223.500 25.800 ;
        RECT 221.400 25.400 223.500 25.700 ;
        RECT 221.400 21.100 221.800 25.400 ;
        RECT 224.700 25.200 225.000 25.800 ;
        RECT 227.800 25.500 230.600 25.600 ;
        RECT 227.700 25.400 230.600 25.500 ;
        RECT 223.800 24.900 225.000 25.200 ;
        RECT 225.700 25.300 230.600 25.400 ;
        RECT 225.700 25.100 228.100 25.300 ;
        RECT 223.800 24.400 224.100 24.900 ;
        RECT 223.400 24.000 224.100 24.400 ;
        RECT 224.900 24.500 225.300 24.600 ;
        RECT 225.700 24.500 226.000 25.100 ;
        RECT 224.900 24.200 226.000 24.500 ;
        RECT 226.300 24.500 229.000 24.800 ;
        RECT 226.300 24.400 226.700 24.500 ;
        RECT 228.600 24.400 229.000 24.500 ;
        RECT 225.500 23.700 225.900 23.800 ;
        RECT 226.900 23.700 227.300 23.800 ;
        RECT 223.800 23.100 224.200 23.500 ;
        RECT 225.500 23.400 227.300 23.700 ;
        RECT 225.900 23.100 226.200 23.400 ;
        RECT 228.600 23.100 229.000 23.500 ;
        RECT 223.500 21.100 224.100 23.100 ;
        RECT 225.800 21.100 226.200 23.100 ;
        RECT 228.000 22.800 229.000 23.100 ;
        RECT 228.000 21.100 228.400 22.800 ;
        RECT 230.200 21.100 230.600 25.300 ;
        RECT 0.600 15.700 1.000 19.900 ;
        RECT 2.800 18.200 3.200 19.900 ;
        RECT 2.200 17.900 3.200 18.200 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.100 17.900 7.700 19.900 ;
        RECT 2.200 17.500 2.600 17.900 ;
        RECT 5.000 17.600 5.300 17.900 ;
        RECT 3.900 17.300 5.700 17.600 ;
        RECT 7.000 17.500 7.400 17.900 ;
        RECT 3.900 17.200 4.300 17.300 ;
        RECT 5.300 17.200 5.700 17.300 ;
        RECT 2.200 16.500 2.600 16.600 ;
        RECT 4.500 16.500 4.900 16.600 ;
        RECT 2.200 16.200 4.900 16.500 ;
        RECT 5.200 16.500 6.300 16.800 ;
        RECT 5.200 15.900 5.500 16.500 ;
        RECT 5.900 16.400 6.300 16.500 ;
        RECT 7.100 16.600 7.800 17.000 ;
        RECT 7.100 16.100 7.400 16.600 ;
        RECT 3.100 15.700 5.500 15.900 ;
        RECT 0.600 15.600 5.500 15.700 ;
        RECT 6.200 15.800 7.400 16.100 ;
        RECT 0.600 15.500 3.500 15.600 ;
        RECT 0.600 15.400 3.400 15.500 ;
        RECT 3.800 15.100 4.200 15.200 ;
        RECT 1.700 14.800 4.200 15.100 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 6.200 15.100 6.500 15.800 ;
        RECT 9.400 15.600 9.800 19.900 ;
        RECT 11.500 16.200 11.900 19.900 ;
        RECT 12.200 16.800 12.600 17.200 ;
        RECT 12.300 16.200 12.600 16.800 ;
        RECT 11.500 15.900 12.000 16.200 ;
        RECT 12.300 15.900 13.000 16.200 ;
        RECT 7.700 15.300 9.800 15.600 ;
        RECT 7.700 15.200 8.100 15.300 ;
        RECT 5.400 14.800 6.500 15.100 ;
        RECT 8.500 14.900 8.900 15.000 ;
        RECT 1.700 14.700 2.100 14.800 ;
        RECT 3.000 14.700 3.400 14.800 ;
        RECT 2.500 14.200 2.900 14.300 ;
        RECT 6.200 14.200 6.500 14.800 ;
        RECT 7.000 14.600 8.900 14.900 ;
        RECT 7.000 14.500 7.400 14.600 ;
        RECT 1.000 13.900 6.500 14.200 ;
        RECT 1.000 13.800 1.800 13.900 ;
        RECT 0.600 11.100 1.000 13.500 ;
        RECT 3.100 12.800 3.400 13.900 ;
        RECT 5.900 13.800 6.300 13.900 ;
        RECT 9.400 13.600 9.800 15.300 ;
        RECT 11.000 14.400 11.400 15.200 ;
        RECT 11.700 14.200 12.000 15.900 ;
        RECT 12.600 15.800 13.000 15.900 ;
        RECT 13.400 15.700 13.800 19.900 ;
        RECT 15.600 18.200 16.000 19.900 ;
        RECT 15.000 17.900 16.000 18.200 ;
        RECT 17.800 17.900 18.200 19.900 ;
        RECT 19.900 17.900 20.500 19.900 ;
        RECT 15.000 17.500 15.400 17.900 ;
        RECT 17.800 17.600 18.100 17.900 ;
        RECT 16.700 17.300 18.500 17.600 ;
        RECT 19.800 17.500 20.200 17.900 ;
        RECT 16.700 17.200 17.100 17.300 ;
        RECT 18.100 17.200 18.500 17.300 ;
        RECT 15.000 16.500 15.400 16.600 ;
        RECT 17.300 16.500 17.700 16.600 ;
        RECT 15.000 16.200 17.700 16.500 ;
        RECT 18.000 16.500 19.100 16.800 ;
        RECT 18.000 15.900 18.300 16.500 ;
        RECT 18.700 16.400 19.100 16.500 ;
        RECT 19.900 16.600 20.600 17.000 ;
        RECT 19.900 16.100 20.200 16.600 ;
        RECT 15.900 15.700 18.300 15.900 ;
        RECT 13.400 15.600 18.300 15.700 ;
        RECT 19.000 15.800 20.200 16.100 ;
        RECT 13.400 15.500 16.300 15.600 ;
        RECT 13.400 15.400 16.200 15.500 ;
        RECT 19.000 15.200 19.300 15.800 ;
        RECT 22.200 15.600 22.600 19.900 ;
        RECT 20.500 15.300 22.600 15.600 ;
        RECT 20.500 15.200 20.900 15.300 ;
        RECT 16.600 15.100 17.000 15.200 ;
        RECT 14.500 14.800 17.000 15.100 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 21.300 14.900 21.700 15.000 ;
        RECT 14.500 14.700 14.900 14.800 ;
        RECT 15.800 14.700 16.200 14.800 ;
        RECT 15.300 14.200 15.700 14.300 ;
        RECT 19.000 14.200 19.300 14.800 ;
        RECT 19.800 14.600 21.700 14.900 ;
        RECT 19.800 14.500 20.200 14.600 ;
        RECT 10.200 14.100 10.600 14.200 ;
        RECT 10.200 13.800 11.000 14.100 ;
        RECT 11.700 13.800 13.000 14.200 ;
        RECT 13.800 13.900 19.300 14.200 ;
        RECT 13.800 13.800 14.600 13.900 ;
        RECT 10.600 13.600 11.000 13.800 ;
        RECT 7.800 13.300 9.800 13.600 ;
        RECT 7.800 13.200 8.300 13.300 ;
        RECT 6.200 13.100 6.600 13.200 ;
        RECT 7.800 13.100 8.200 13.200 ;
        RECT 6.200 12.800 8.200 13.100 ;
        RECT 2.200 12.100 2.600 12.500 ;
        RECT 3.000 12.400 3.400 12.800 ;
        RECT 3.900 12.700 4.300 12.800 ;
        RECT 3.900 12.400 5.300 12.700 ;
        RECT 5.000 12.100 5.300 12.400 ;
        RECT 7.000 12.100 7.400 12.500 ;
        RECT 2.200 11.800 3.200 12.100 ;
        RECT 2.800 11.100 3.200 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.000 11.800 7.700 12.100 ;
        RECT 7.100 11.100 7.700 11.800 ;
        RECT 9.400 11.100 9.800 13.300 ;
        RECT 10.300 13.100 12.100 13.300 ;
        RECT 12.600 13.100 12.900 13.800 ;
        RECT 10.200 13.000 12.200 13.100 ;
        RECT 10.200 11.100 10.600 13.000 ;
        RECT 11.800 11.100 12.200 13.000 ;
        RECT 12.600 11.100 13.000 13.100 ;
        RECT 13.400 11.100 13.800 13.500 ;
        RECT 15.900 12.800 16.200 13.900 ;
        RECT 18.700 13.800 19.100 13.900 ;
        RECT 22.200 13.600 22.600 15.300 ;
        RECT 20.600 13.300 22.600 13.600 ;
        RECT 20.600 13.200 21.100 13.300 ;
        RECT 19.000 13.100 19.400 13.200 ;
        RECT 20.600 13.100 21.000 13.200 ;
        RECT 19.000 12.800 21.000 13.100 ;
        RECT 22.200 13.100 22.600 13.300 ;
        RECT 23.000 13.100 23.400 13.200 ;
        RECT 22.200 12.800 23.400 13.100 ;
        RECT 15.000 12.100 15.400 12.500 ;
        RECT 15.800 12.400 16.200 12.800 ;
        RECT 16.700 12.700 17.100 12.800 ;
        RECT 16.700 12.400 18.100 12.700 ;
        RECT 17.800 12.100 18.100 12.400 ;
        RECT 19.800 12.100 20.200 12.500 ;
        RECT 15.000 11.800 16.000 12.100 ;
        RECT 15.600 11.100 16.000 11.800 ;
        RECT 17.800 11.100 18.200 12.100 ;
        RECT 19.800 11.800 20.500 12.100 ;
        RECT 19.900 11.100 20.500 11.800 ;
        RECT 22.200 11.100 22.600 12.800 ;
        RECT 23.000 12.400 23.400 12.800 ;
        RECT 23.800 11.100 24.200 19.900 ;
        RECT 24.600 15.700 25.000 19.900 ;
        RECT 26.800 18.200 27.200 19.900 ;
        RECT 26.200 17.900 27.200 18.200 ;
        RECT 29.000 17.900 29.400 19.900 ;
        RECT 31.100 17.900 31.700 19.900 ;
        RECT 26.200 17.500 26.600 17.900 ;
        RECT 29.000 17.600 29.300 17.900 ;
        RECT 27.900 17.300 29.700 17.600 ;
        RECT 31.000 17.500 31.400 17.900 ;
        RECT 27.900 17.200 28.300 17.300 ;
        RECT 29.300 17.200 29.700 17.300 ;
        RECT 26.200 16.500 26.600 16.600 ;
        RECT 28.500 16.500 28.900 16.600 ;
        RECT 26.200 16.200 28.900 16.500 ;
        RECT 29.200 16.500 30.300 16.800 ;
        RECT 29.200 15.900 29.500 16.500 ;
        RECT 29.900 16.400 30.300 16.500 ;
        RECT 31.100 16.600 31.800 17.000 ;
        RECT 31.100 16.100 31.400 16.600 ;
        RECT 27.100 15.700 29.500 15.900 ;
        RECT 24.600 15.600 29.500 15.700 ;
        RECT 30.200 15.800 31.400 16.100 ;
        RECT 24.600 15.500 27.500 15.600 ;
        RECT 24.600 15.400 27.400 15.500 ;
        RECT 30.200 15.200 30.500 15.800 ;
        RECT 33.400 15.600 33.800 19.900 ;
        RECT 34.600 16.800 35.000 17.200 ;
        RECT 34.600 16.200 34.900 16.800 ;
        RECT 35.300 16.200 35.700 19.900 ;
        RECT 40.900 19.200 41.300 19.900 ;
        RECT 40.600 18.800 41.300 19.200 ;
        RECT 40.900 16.400 41.300 18.800 ;
        RECT 43.000 17.500 43.400 19.500 ;
        RECT 34.200 15.900 34.900 16.200 ;
        RECT 35.200 15.900 35.700 16.200 ;
        RECT 40.500 16.100 41.300 16.400 ;
        RECT 34.200 15.800 34.600 15.900 ;
        RECT 31.700 15.300 33.800 15.600 ;
        RECT 31.700 15.200 32.100 15.300 ;
        RECT 27.800 15.100 28.200 15.200 ;
        RECT 28.600 15.100 29.000 15.200 ;
        RECT 25.700 14.800 29.000 15.100 ;
        RECT 30.200 14.800 30.600 15.200 ;
        RECT 32.500 14.900 32.900 15.000 ;
        RECT 25.700 14.700 26.100 14.800 ;
        RECT 26.500 14.200 26.900 14.300 ;
        RECT 30.200 14.200 30.500 14.800 ;
        RECT 31.000 14.600 32.900 14.900 ;
        RECT 31.000 14.500 31.400 14.600 ;
        RECT 25.000 13.900 30.500 14.200 ;
        RECT 25.000 13.800 25.800 13.900 ;
        RECT 24.600 11.100 25.000 13.500 ;
        RECT 27.100 12.800 27.400 13.900 ;
        RECT 29.900 13.800 30.300 13.900 ;
        RECT 33.400 13.600 33.800 15.300 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 35.200 15.100 35.500 15.900 ;
        RECT 34.200 14.800 35.500 15.100 ;
        RECT 35.200 14.200 35.500 14.800 ;
        RECT 35.800 15.100 36.200 15.200 ;
        RECT 37.400 15.100 37.800 15.200 ;
        RECT 35.800 14.800 37.800 15.100 ;
        RECT 39.000 15.100 39.400 15.200 ;
        RECT 39.800 15.100 40.200 15.600 ;
        RECT 39.000 14.800 40.200 15.100 ;
        RECT 35.800 14.400 36.200 14.800 ;
        RECT 40.500 14.200 40.800 16.100 ;
        RECT 43.100 15.800 43.400 17.500 ;
        RECT 43.800 16.200 44.200 19.900 ;
        RECT 45.400 16.400 45.800 19.900 ;
        RECT 43.800 15.900 45.100 16.200 ;
        RECT 45.400 15.900 45.900 16.400 ;
        RECT 41.500 15.500 43.400 15.800 ;
        RECT 41.500 14.500 41.800 15.500 ;
        RECT 34.200 13.800 35.500 14.200 ;
        RECT 36.600 14.100 37.000 14.200 ;
        RECT 36.200 13.800 37.000 14.100 ;
        RECT 39.800 13.800 40.800 14.200 ;
        RECT 41.100 14.100 41.800 14.500 ;
        RECT 42.200 14.400 42.600 15.200 ;
        RECT 43.000 14.400 43.400 15.200 ;
        RECT 43.800 14.800 44.300 15.200 ;
        RECT 43.900 14.400 44.300 14.800 ;
        RECT 44.800 14.900 45.100 15.900 ;
        RECT 44.800 14.500 45.300 14.900 ;
        RECT 31.900 13.300 33.800 13.600 ;
        RECT 31.900 13.200 32.300 13.300 ;
        RECT 26.200 12.100 26.600 12.500 ;
        RECT 27.000 12.400 27.400 12.800 ;
        RECT 27.900 12.700 28.300 12.800 ;
        RECT 27.900 12.400 29.300 12.700 ;
        RECT 29.000 12.100 29.300 12.400 ;
        RECT 31.000 12.100 31.400 12.500 ;
        RECT 26.200 11.800 27.200 12.100 ;
        RECT 26.800 11.100 27.200 11.800 ;
        RECT 29.000 11.100 29.400 12.100 ;
        RECT 31.000 11.800 31.700 12.100 ;
        RECT 31.100 11.100 31.700 11.800 ;
        RECT 33.400 11.100 33.800 13.300 ;
        RECT 34.300 13.100 34.600 13.800 ;
        RECT 36.200 13.600 36.600 13.800 ;
        RECT 40.500 13.500 40.800 13.800 ;
        RECT 41.300 13.900 41.800 14.100 ;
        RECT 41.300 13.600 43.400 13.900 ;
        RECT 44.800 13.700 45.100 14.500 ;
        RECT 45.600 14.200 45.900 15.900 ;
        RECT 47.000 15.700 47.400 19.900 ;
        RECT 49.200 18.200 49.600 19.900 ;
        RECT 48.600 17.900 49.600 18.200 ;
        RECT 51.400 17.900 51.800 19.900 ;
        RECT 53.500 17.900 54.100 19.900 ;
        RECT 48.600 17.500 49.000 17.900 ;
        RECT 51.400 17.600 51.700 17.900 ;
        RECT 50.300 17.300 52.100 17.600 ;
        RECT 53.400 17.500 53.800 17.900 ;
        RECT 50.300 17.200 50.700 17.300 ;
        RECT 51.700 17.200 52.100 17.300 ;
        RECT 48.600 16.500 49.000 16.600 ;
        RECT 50.900 16.500 51.300 16.600 ;
        RECT 48.600 16.200 51.300 16.500 ;
        RECT 51.600 16.500 52.700 16.800 ;
        RECT 51.600 15.900 51.900 16.500 ;
        RECT 52.300 16.400 52.700 16.500 ;
        RECT 53.500 16.600 54.200 17.000 ;
        RECT 53.500 16.100 53.800 16.600 ;
        RECT 49.500 15.700 51.900 15.900 ;
        RECT 47.000 15.600 51.900 15.700 ;
        RECT 52.600 15.800 53.800 16.100 ;
        RECT 47.000 15.500 49.900 15.600 ;
        RECT 47.000 15.400 49.800 15.500 ;
        RECT 45.400 14.100 45.900 14.200 ;
        RECT 46.200 14.800 46.600 15.200 ;
        RECT 50.200 15.100 50.600 15.200 ;
        RECT 51.800 15.100 52.200 15.200 ;
        RECT 48.100 14.800 52.200 15.100 ;
        RECT 46.200 14.100 46.500 14.800 ;
        RECT 48.100 14.700 48.500 14.800 ;
        RECT 48.900 14.200 49.300 14.300 ;
        RECT 52.600 14.200 52.900 15.800 ;
        RECT 55.800 15.600 56.200 19.900 ;
        RECT 57.900 16.200 58.300 19.900 ;
        RECT 58.600 16.800 59.000 17.200 ;
        RECT 58.700 16.200 59.000 16.800 ;
        RECT 57.900 15.900 58.400 16.200 ;
        RECT 58.700 15.900 59.400 16.200 ;
        RECT 54.100 15.300 56.200 15.600 ;
        RECT 54.100 15.200 54.500 15.300 ;
        RECT 54.900 14.900 55.300 15.000 ;
        RECT 53.400 14.600 55.300 14.900 ;
        RECT 53.400 14.500 53.800 14.600 ;
        RECT 45.400 13.800 46.500 14.100 ;
        RECT 47.400 13.900 52.900 14.200 ;
        RECT 47.400 13.800 48.200 13.900 ;
        RECT 40.500 13.300 40.900 13.500 ;
        RECT 35.100 13.100 36.900 13.300 ;
        RECT 34.200 11.100 34.600 13.100 ;
        RECT 35.000 13.000 37.000 13.100 ;
        RECT 40.500 13.000 41.300 13.300 ;
        RECT 35.000 11.100 35.400 13.000 ;
        RECT 36.600 11.100 37.000 13.000 ;
        RECT 40.900 11.500 41.300 13.000 ;
        RECT 43.100 12.500 43.400 13.600 ;
        RECT 43.000 11.500 43.400 12.500 ;
        RECT 43.800 13.400 45.100 13.700 ;
        RECT 43.800 11.100 44.200 13.400 ;
        RECT 45.600 13.100 45.900 13.800 ;
        RECT 45.400 12.800 45.900 13.100 ;
        RECT 45.400 11.100 45.800 12.800 ;
        RECT 47.000 11.100 47.400 13.500 ;
        RECT 49.500 12.800 49.800 13.900 ;
        RECT 52.300 13.800 52.700 13.900 ;
        RECT 55.800 13.600 56.200 15.300 ;
        RECT 57.400 14.400 57.800 15.200 ;
        RECT 58.100 14.200 58.400 15.900 ;
        RECT 59.000 15.800 59.400 15.900 ;
        RECT 59.800 15.800 60.200 16.600 ;
        RECT 59.000 15.100 59.300 15.800 ;
        RECT 60.600 15.100 61.000 19.900 ;
        RECT 59.000 14.800 61.000 15.100 ;
        RECT 56.600 14.100 57.000 14.200 ;
        RECT 56.600 13.800 57.400 14.100 ;
        RECT 58.100 13.800 59.400 14.200 ;
        RECT 57.000 13.600 57.400 13.800 ;
        RECT 54.300 13.300 56.200 13.600 ;
        RECT 54.300 13.200 54.700 13.300 ;
        RECT 48.600 12.100 49.000 12.500 ;
        RECT 49.400 12.400 49.800 12.800 ;
        RECT 50.300 12.700 50.700 12.800 ;
        RECT 50.300 12.400 51.700 12.700 ;
        RECT 51.400 12.100 51.700 12.400 ;
        RECT 53.400 12.100 53.800 12.500 ;
        RECT 48.600 11.800 49.600 12.100 ;
        RECT 49.200 11.100 49.600 11.800 ;
        RECT 51.400 11.100 51.800 12.100 ;
        RECT 53.400 11.800 54.100 12.100 ;
        RECT 53.500 11.100 54.100 11.800 ;
        RECT 55.800 11.100 56.200 13.300 ;
        RECT 56.700 13.100 58.500 13.300 ;
        RECT 59.000 13.100 59.300 13.800 ;
        RECT 60.600 13.100 61.000 14.800 ;
        RECT 61.400 14.100 61.800 14.200 ;
        RECT 61.400 13.800 62.500 14.100 ;
        RECT 61.400 13.400 61.800 13.800 ;
        RECT 56.600 13.000 58.600 13.100 ;
        RECT 56.600 11.100 57.000 13.000 ;
        RECT 58.200 11.100 58.600 13.000 ;
        RECT 59.000 11.100 59.400 13.100 ;
        RECT 60.100 12.800 61.000 13.100 ;
        RECT 62.200 13.200 62.500 13.800 ;
        RECT 60.100 11.100 60.500 12.800 ;
        RECT 62.200 12.400 62.600 13.200 ;
        RECT 63.000 11.100 63.400 19.900 ;
        RECT 65.100 16.200 65.500 19.900 ;
        RECT 65.800 16.800 66.200 17.200 ;
        RECT 65.900 16.200 66.200 16.800 ;
        RECT 65.100 15.900 65.600 16.200 ;
        RECT 65.900 15.900 66.600 16.200 ;
        RECT 64.600 14.400 65.000 15.200 ;
        RECT 65.300 14.200 65.600 15.900 ;
        RECT 66.200 15.800 66.600 15.900 ;
        RECT 67.000 15.800 67.400 16.600 ;
        RECT 66.200 15.100 66.500 15.800 ;
        RECT 67.800 15.100 68.200 19.900 ;
        RECT 69.400 15.700 69.800 19.900 ;
        RECT 71.600 18.200 72.000 19.900 ;
        RECT 71.000 17.900 72.000 18.200 ;
        RECT 73.800 17.900 74.200 19.900 ;
        RECT 75.900 17.900 76.500 19.900 ;
        RECT 71.000 17.500 71.400 17.900 ;
        RECT 73.800 17.600 74.100 17.900 ;
        RECT 72.700 17.300 74.500 17.600 ;
        RECT 75.800 17.500 76.200 17.900 ;
        RECT 72.700 17.200 73.100 17.300 ;
        RECT 74.100 17.200 74.500 17.300 ;
        RECT 71.000 16.500 71.400 16.600 ;
        RECT 73.300 16.500 73.700 16.600 ;
        RECT 71.000 16.200 73.700 16.500 ;
        RECT 74.000 16.500 75.100 16.800 ;
        RECT 74.000 15.900 74.300 16.500 ;
        RECT 74.700 16.400 75.100 16.500 ;
        RECT 75.900 16.600 76.600 17.000 ;
        RECT 75.900 16.100 76.200 16.600 ;
        RECT 71.900 15.700 74.300 15.900 ;
        RECT 69.400 15.600 74.300 15.700 ;
        RECT 75.000 15.800 76.200 16.100 ;
        RECT 69.400 15.500 72.300 15.600 ;
        RECT 69.400 15.400 72.200 15.500 ;
        RECT 72.600 15.100 73.000 15.200 ;
        RECT 66.200 14.800 68.200 15.100 ;
        RECT 63.800 14.100 64.200 14.200 ;
        RECT 65.300 14.100 66.600 14.200 ;
        RECT 67.000 14.100 67.400 14.200 ;
        RECT 63.800 13.800 64.600 14.100 ;
        RECT 65.300 13.800 67.400 14.100 ;
        RECT 64.200 13.600 64.600 13.800 ;
        RECT 63.900 13.100 65.700 13.300 ;
        RECT 66.200 13.100 66.500 13.800 ;
        RECT 67.800 13.100 68.200 14.800 ;
        RECT 70.500 14.800 73.000 15.100 ;
        RECT 70.500 14.700 70.900 14.800 ;
        RECT 71.800 14.700 72.200 14.800 ;
        RECT 71.300 14.200 71.700 14.300 ;
        RECT 75.000 14.200 75.300 15.800 ;
        RECT 78.200 15.600 78.600 19.900 ;
        RECT 76.500 15.300 78.600 15.600 ;
        RECT 76.500 15.200 76.900 15.300 ;
        RECT 77.300 14.900 77.700 15.000 ;
        RECT 75.800 14.600 77.700 14.900 ;
        RECT 75.800 14.500 76.200 14.600 ;
        RECT 68.600 13.400 69.000 14.200 ;
        RECT 69.800 13.900 75.300 14.200 ;
        RECT 69.800 13.800 70.600 13.900 ;
        RECT 63.800 13.000 65.800 13.100 ;
        RECT 63.800 11.100 64.200 13.000 ;
        RECT 65.400 11.100 65.800 13.000 ;
        RECT 66.200 11.100 66.600 13.100 ;
        RECT 67.300 12.800 68.200 13.100 ;
        RECT 67.300 11.100 67.700 12.800 ;
        RECT 69.400 11.100 69.800 13.500 ;
        RECT 71.900 13.200 72.200 13.900 ;
        RECT 72.600 13.800 73.000 13.900 ;
        RECT 74.700 13.800 75.100 13.900 ;
        RECT 76.600 13.600 77.000 14.200 ;
        RECT 78.200 13.600 78.600 15.300 ;
        RECT 76.600 13.300 78.600 13.600 ;
        RECT 79.000 13.400 79.400 14.200 ;
        RECT 76.700 13.200 77.100 13.300 ;
        RECT 71.000 12.100 71.400 12.500 ;
        RECT 71.800 12.400 72.200 13.200 ;
        RECT 72.700 12.700 73.100 12.800 ;
        RECT 72.700 12.400 74.100 12.700 ;
        RECT 73.800 12.100 74.100 12.400 ;
        RECT 75.800 12.100 76.200 12.500 ;
        RECT 71.000 11.800 72.000 12.100 ;
        RECT 71.600 11.100 72.000 11.800 ;
        RECT 73.800 11.100 74.200 12.100 ;
        RECT 75.800 11.800 76.500 12.100 ;
        RECT 75.900 11.100 76.500 11.800 ;
        RECT 78.200 11.100 78.600 13.300 ;
        RECT 79.800 11.100 80.200 19.900 ;
        RECT 80.600 13.400 81.000 14.200 ;
        RECT 81.400 11.100 81.800 19.900 ;
        RECT 83.500 16.200 83.900 19.900 ;
        RECT 84.200 16.800 84.600 17.200 ;
        RECT 84.300 16.200 84.600 16.800 ;
        RECT 83.500 15.900 84.000 16.200 ;
        RECT 84.300 15.900 85.000 16.200 ;
        RECT 83.000 14.400 83.400 15.200 ;
        RECT 83.700 14.200 84.000 15.900 ;
        RECT 84.600 15.800 85.000 15.900 ;
        RECT 85.400 15.800 85.800 16.600 ;
        RECT 84.600 15.100 84.900 15.800 ;
        RECT 86.200 15.100 86.600 19.900 ;
        RECT 89.400 15.700 89.800 19.900 ;
        RECT 91.600 18.200 92.000 19.900 ;
        RECT 91.000 17.900 92.000 18.200 ;
        RECT 93.800 17.900 94.200 19.900 ;
        RECT 95.900 17.900 96.500 19.900 ;
        RECT 91.000 17.500 91.400 17.900 ;
        RECT 93.800 17.600 94.100 17.900 ;
        RECT 92.700 17.300 94.500 17.600 ;
        RECT 95.800 17.500 96.200 17.900 ;
        RECT 92.700 17.200 93.100 17.300 ;
        RECT 94.100 17.200 94.500 17.300 ;
        RECT 91.000 16.500 91.400 16.600 ;
        RECT 93.300 16.500 93.700 16.600 ;
        RECT 91.000 16.200 93.700 16.500 ;
        RECT 94.000 16.500 95.100 16.800 ;
        RECT 94.000 15.900 94.300 16.500 ;
        RECT 94.700 16.400 95.100 16.500 ;
        RECT 95.900 16.600 96.600 17.000 ;
        RECT 95.900 16.100 96.200 16.600 ;
        RECT 91.900 15.700 94.300 15.900 ;
        RECT 89.400 15.600 94.300 15.700 ;
        RECT 95.000 15.800 96.200 16.100 ;
        RECT 89.400 15.500 92.300 15.600 ;
        RECT 89.400 15.400 92.200 15.500 ;
        RECT 92.600 15.100 93.000 15.200 ;
        RECT 84.600 14.800 86.600 15.100 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 83.700 14.100 85.000 14.200 ;
        RECT 85.400 14.100 85.800 14.200 ;
        RECT 82.200 13.800 83.000 14.100 ;
        RECT 83.700 13.800 85.800 14.100 ;
        RECT 82.600 13.600 83.000 13.800 ;
        RECT 82.300 13.100 84.100 13.300 ;
        RECT 84.600 13.100 84.900 13.800 ;
        RECT 86.200 13.100 86.600 14.800 ;
        RECT 90.500 14.800 93.000 15.100 ;
        RECT 90.500 14.700 90.900 14.800 ;
        RECT 91.300 14.200 91.700 14.300 ;
        RECT 95.000 14.200 95.300 15.800 ;
        RECT 98.200 15.600 98.600 19.900 ;
        RECT 96.500 15.300 98.600 15.600 ;
        RECT 96.500 15.200 96.900 15.300 ;
        RECT 97.300 14.900 97.700 15.000 ;
        RECT 95.800 14.600 97.700 14.900 ;
        RECT 95.800 14.500 96.200 14.600 ;
        RECT 87.000 14.100 87.400 14.200 ;
        RECT 88.600 14.100 89.000 14.200 ;
        RECT 87.000 13.800 89.000 14.100 ;
        RECT 89.800 13.900 95.300 14.200 ;
        RECT 89.800 13.800 90.600 13.900 ;
        RECT 91.800 13.800 92.200 13.900 ;
        RECT 94.700 13.800 95.100 13.900 ;
        RECT 87.000 13.400 87.400 13.800 ;
        RECT 82.200 13.000 84.200 13.100 ;
        RECT 82.200 11.100 82.600 13.000 ;
        RECT 83.800 11.100 84.200 13.000 ;
        RECT 84.600 11.100 85.000 13.100 ;
        RECT 85.700 12.800 86.600 13.100 ;
        RECT 85.700 11.100 86.100 12.800 ;
        RECT 89.400 11.100 89.800 13.500 ;
        RECT 91.900 12.800 92.200 13.800 ;
        RECT 98.200 13.600 98.600 15.300 ;
        RECT 96.700 13.300 98.600 13.600 ;
        RECT 96.700 13.200 97.100 13.300 ;
        RECT 91.000 12.100 91.400 12.500 ;
        RECT 91.800 12.400 92.200 12.800 ;
        RECT 92.700 12.700 93.100 12.800 ;
        RECT 92.700 12.400 94.100 12.700 ;
        RECT 93.800 12.100 94.100 12.400 ;
        RECT 95.800 12.100 96.200 12.500 ;
        RECT 91.000 11.800 92.000 12.100 ;
        RECT 91.600 11.100 92.000 11.800 ;
        RECT 93.800 11.100 94.200 12.100 ;
        RECT 95.800 11.800 96.500 12.100 ;
        RECT 95.900 11.100 96.500 11.800 ;
        RECT 98.200 11.100 98.600 13.300 ;
        RECT 99.000 12.400 99.400 13.200 ;
        RECT 99.800 11.100 100.200 19.900 ;
        RECT 100.600 15.700 101.000 19.900 ;
        RECT 102.800 18.200 103.200 19.900 ;
        RECT 102.200 17.900 103.200 18.200 ;
        RECT 105.000 17.900 105.400 19.900 ;
        RECT 107.100 17.900 107.700 19.900 ;
        RECT 102.200 17.500 102.600 17.900 ;
        RECT 105.000 17.600 105.300 17.900 ;
        RECT 103.900 17.300 105.700 17.600 ;
        RECT 107.000 17.500 107.400 17.900 ;
        RECT 103.900 17.200 104.300 17.300 ;
        RECT 105.300 17.200 105.700 17.300 ;
        RECT 102.200 16.500 102.600 16.600 ;
        RECT 104.500 16.500 104.900 16.600 ;
        RECT 102.200 16.200 104.900 16.500 ;
        RECT 105.200 16.500 106.300 16.800 ;
        RECT 105.200 15.900 105.500 16.500 ;
        RECT 105.900 16.400 106.300 16.500 ;
        RECT 107.100 16.600 107.800 17.000 ;
        RECT 107.100 16.100 107.400 16.600 ;
        RECT 103.100 15.700 105.500 15.900 ;
        RECT 100.600 15.600 105.500 15.700 ;
        RECT 106.200 15.800 107.400 16.100 ;
        RECT 100.600 15.500 103.500 15.600 ;
        RECT 100.600 15.400 103.400 15.500 ;
        RECT 106.200 15.200 106.500 15.800 ;
        RECT 109.400 15.600 109.800 19.900 ;
        RECT 111.500 16.200 111.900 19.900 ;
        RECT 112.200 16.800 112.600 17.200 ;
        RECT 112.300 16.200 112.600 16.800 ;
        RECT 111.000 15.800 112.000 16.200 ;
        RECT 112.300 15.900 113.000 16.200 ;
        RECT 107.700 15.300 109.800 15.600 ;
        RECT 107.700 15.200 108.100 15.300 ;
        RECT 103.800 15.100 104.200 15.200 ;
        RECT 101.700 14.800 104.200 15.100 ;
        RECT 106.200 14.800 106.600 15.200 ;
        RECT 108.500 14.900 108.900 15.000 ;
        RECT 101.700 14.700 102.100 14.800 ;
        RECT 102.500 14.200 102.900 14.300 ;
        RECT 106.200 14.200 106.500 14.800 ;
        RECT 107.000 14.600 108.900 14.900 ;
        RECT 107.000 14.500 107.400 14.600 ;
        RECT 101.000 13.900 106.500 14.200 ;
        RECT 101.000 13.800 101.800 13.900 ;
        RECT 100.600 11.100 101.000 13.500 ;
        RECT 103.100 12.800 103.400 13.900 ;
        RECT 105.900 13.800 106.300 13.900 ;
        RECT 109.400 13.600 109.800 15.300 ;
        RECT 110.200 15.100 110.600 15.200 ;
        RECT 111.000 15.100 111.400 15.200 ;
        RECT 110.200 14.800 111.400 15.100 ;
        RECT 111.000 14.400 111.400 14.800 ;
        RECT 111.700 14.200 112.000 15.800 ;
        RECT 112.600 15.800 113.000 15.900 ;
        RECT 113.400 15.800 113.800 16.600 ;
        RECT 112.600 15.100 112.900 15.800 ;
        RECT 114.200 15.100 114.600 19.900 ;
        RECT 115.800 17.500 116.200 19.500 ;
        RECT 117.900 19.200 118.300 19.900 ;
        RECT 117.900 18.800 118.600 19.200 ;
        RECT 115.800 15.800 116.100 17.500 ;
        RECT 117.900 16.400 118.300 18.800 ;
        RECT 117.900 16.100 118.700 16.400 ;
        RECT 115.800 15.500 117.700 15.800 ;
        RECT 112.600 14.800 114.600 15.100 ;
        RECT 110.200 14.100 110.600 14.200 ;
        RECT 110.200 13.800 111.000 14.100 ;
        RECT 111.700 13.800 113.000 14.200 ;
        RECT 110.600 13.600 111.000 13.800 ;
        RECT 107.900 13.300 109.800 13.600 ;
        RECT 107.900 13.200 108.300 13.300 ;
        RECT 102.200 12.100 102.600 12.500 ;
        RECT 103.000 12.400 103.400 12.800 ;
        RECT 103.900 12.700 104.300 12.800 ;
        RECT 103.900 12.400 105.300 12.700 ;
        RECT 105.000 12.100 105.300 12.400 ;
        RECT 107.000 12.100 107.400 12.500 ;
        RECT 102.200 11.800 103.200 12.100 ;
        RECT 102.800 11.100 103.200 11.800 ;
        RECT 105.000 11.100 105.400 12.100 ;
        RECT 107.000 11.800 107.700 12.100 ;
        RECT 107.100 11.100 107.700 11.800 ;
        RECT 109.400 11.100 109.800 13.300 ;
        RECT 110.300 13.100 112.100 13.300 ;
        RECT 112.600 13.100 112.900 13.800 ;
        RECT 114.200 13.100 114.600 14.800 ;
        RECT 115.800 14.400 116.200 15.200 ;
        RECT 116.600 14.400 117.000 15.200 ;
        RECT 117.400 14.500 117.700 15.500 ;
        RECT 115.000 13.400 115.400 14.200 ;
        RECT 117.400 14.100 118.100 14.500 ;
        RECT 118.400 14.200 118.700 16.100 ;
        RECT 121.900 16.200 122.300 19.900 ;
        RECT 122.600 16.800 123.000 17.200 ;
        RECT 122.700 16.200 123.000 16.800 ;
        RECT 121.900 15.900 122.400 16.200 ;
        RECT 122.700 15.900 123.400 16.200 ;
        RECT 119.000 14.800 119.400 15.600 ;
        RECT 121.400 14.400 121.800 15.200 ;
        RECT 122.100 14.200 122.400 15.900 ;
        RECT 123.000 15.800 123.400 15.900 ;
        RECT 123.800 15.800 124.200 16.600 ;
        RECT 123.000 15.100 123.300 15.800 ;
        RECT 124.600 15.100 125.000 19.900 ;
        RECT 126.200 16.200 126.600 19.900 ;
        RECT 127.800 16.400 128.200 19.900 ;
        RECT 126.200 15.900 127.500 16.200 ;
        RECT 127.800 15.900 128.300 16.400 ;
        RECT 123.000 14.800 125.000 15.100 ;
        RECT 126.200 14.800 126.700 15.200 ;
        RECT 117.400 13.900 117.900 14.100 ;
        RECT 115.800 13.600 117.900 13.900 ;
        RECT 118.400 13.800 119.400 14.200 ;
        RECT 120.600 14.100 121.000 14.200 ;
        RECT 120.600 13.800 121.400 14.100 ;
        RECT 122.100 13.800 123.400 14.200 ;
        RECT 110.200 13.000 112.200 13.100 ;
        RECT 110.200 11.100 110.600 13.000 ;
        RECT 111.800 11.100 112.200 13.000 ;
        RECT 112.600 11.100 113.000 13.100 ;
        RECT 113.700 12.800 114.600 13.100 ;
        RECT 113.700 11.100 114.100 12.800 ;
        RECT 115.800 12.500 116.100 13.600 ;
        RECT 118.400 13.500 118.700 13.800 ;
        RECT 121.000 13.600 121.400 13.800 ;
        RECT 118.300 13.300 118.700 13.500 ;
        RECT 117.900 13.000 118.700 13.300 ;
        RECT 120.700 13.100 122.500 13.300 ;
        RECT 123.000 13.100 123.300 13.800 ;
        RECT 124.600 13.100 125.000 14.800 ;
        RECT 126.300 14.400 126.700 14.800 ;
        RECT 127.200 14.900 127.500 15.900 ;
        RECT 127.200 14.500 127.700 14.900 ;
        RECT 125.400 13.400 125.800 14.200 ;
        RECT 127.200 13.700 127.500 14.500 ;
        RECT 128.000 14.200 128.300 15.900 ;
        RECT 127.800 13.800 128.300 14.200 ;
        RECT 126.200 13.400 127.500 13.700 ;
        RECT 120.600 13.000 122.600 13.100 ;
        RECT 115.800 11.500 116.200 12.500 ;
        RECT 117.900 11.500 118.300 13.000 ;
        RECT 120.600 11.100 121.000 13.000 ;
        RECT 122.200 11.100 122.600 13.000 ;
        RECT 123.000 11.100 123.400 13.100 ;
        RECT 124.100 12.800 125.000 13.100 ;
        RECT 124.100 11.100 124.500 12.800 ;
        RECT 126.200 11.100 126.600 13.400 ;
        RECT 128.000 13.100 128.300 13.800 ;
        RECT 129.400 13.400 129.800 14.200 ;
        RECT 127.800 12.800 128.300 13.100 ;
        RECT 130.200 13.100 130.600 19.900 ;
        RECT 133.700 19.200 134.100 19.900 ;
        RECT 133.700 18.800 134.600 19.200 ;
        RECT 131.000 15.800 131.400 16.600 ;
        RECT 133.700 16.400 134.100 18.800 ;
        RECT 135.800 17.500 136.200 19.500 ;
        RECT 133.300 16.100 134.100 16.400 ;
        RECT 132.600 14.800 133.000 15.600 ;
        RECT 133.300 14.200 133.600 16.100 ;
        RECT 135.900 15.800 136.200 17.500 ;
        RECT 134.300 15.500 136.200 15.800 ;
        RECT 134.300 14.500 134.600 15.500 ;
        RECT 132.600 13.800 133.600 14.200 ;
        RECT 133.900 14.100 134.600 14.500 ;
        RECT 135.000 14.400 135.400 15.200 ;
        RECT 135.800 14.400 136.200 15.200 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 137.400 15.100 137.800 19.900 ;
        RECT 141.000 16.800 141.400 17.200 ;
        RECT 138.200 15.800 138.600 16.600 ;
        RECT 141.000 16.200 141.300 16.800 ;
        RECT 141.700 16.200 142.100 19.900 ;
        RECT 145.700 19.200 146.100 19.900 ;
        RECT 145.700 18.800 146.600 19.200 ;
        RECT 145.700 16.400 146.100 18.800 ;
        RECT 147.800 17.500 148.200 19.500 ;
        RECT 140.600 15.900 141.300 16.200 ;
        RECT 141.600 15.900 142.100 16.200 ;
        RECT 145.300 16.100 146.100 16.400 ;
        RECT 140.600 15.800 141.000 15.900 ;
        RECT 140.600 15.100 140.900 15.800 ;
        RECT 137.400 14.800 140.900 15.100 ;
        RECT 133.300 13.500 133.600 13.800 ;
        RECT 134.100 13.900 134.600 14.100 ;
        RECT 136.600 14.200 136.900 14.800 ;
        RECT 134.100 13.600 136.200 13.900 ;
        RECT 133.300 13.300 133.700 13.500 ;
        RECT 130.200 12.800 131.100 13.100 ;
        RECT 133.300 13.000 134.100 13.300 ;
        RECT 127.800 11.100 128.200 12.800 ;
        RECT 130.700 12.200 131.100 12.800 ;
        RECT 130.200 11.800 131.100 12.200 ;
        RECT 130.700 11.100 131.100 11.800 ;
        RECT 133.700 11.500 134.100 13.000 ;
        RECT 135.900 12.500 136.200 13.600 ;
        RECT 136.600 13.400 137.000 14.200 ;
        RECT 137.400 13.100 137.800 14.800 ;
        RECT 141.600 14.200 141.900 15.900 ;
        RECT 142.200 14.400 142.600 15.200 ;
        RECT 143.800 15.100 144.200 15.200 ;
        RECT 144.600 15.100 145.000 15.600 ;
        RECT 143.800 14.800 145.000 15.100 ;
        RECT 145.300 14.200 145.600 16.100 ;
        RECT 147.900 15.800 148.200 17.500 ;
        RECT 146.300 15.500 148.200 15.800 ;
        RECT 148.600 15.700 149.000 19.900 ;
        RECT 150.800 18.200 151.200 19.900 ;
        RECT 150.200 17.900 151.200 18.200 ;
        RECT 153.000 17.900 153.400 19.900 ;
        RECT 155.100 17.900 155.700 19.900 ;
        RECT 150.200 17.500 150.600 17.900 ;
        RECT 153.000 17.600 153.300 17.900 ;
        RECT 151.900 17.300 153.700 17.600 ;
        RECT 155.000 17.500 155.400 17.900 ;
        RECT 151.900 17.200 152.300 17.300 ;
        RECT 153.300 17.200 153.700 17.300 ;
        RECT 150.200 16.500 150.600 16.600 ;
        RECT 152.500 16.500 152.900 16.600 ;
        RECT 150.200 16.200 152.900 16.500 ;
        RECT 153.200 16.500 154.300 16.800 ;
        RECT 153.200 15.900 153.500 16.500 ;
        RECT 153.900 16.400 154.300 16.500 ;
        RECT 155.100 16.600 155.800 17.000 ;
        RECT 155.100 16.100 155.400 16.600 ;
        RECT 151.100 15.700 153.500 15.900 ;
        RECT 148.600 15.600 153.500 15.700 ;
        RECT 154.200 15.800 155.400 16.100 ;
        RECT 148.600 15.500 151.500 15.600 ;
        RECT 146.300 14.500 146.600 15.500 ;
        RECT 148.600 15.400 151.400 15.500 ;
        RECT 140.600 13.800 141.900 14.200 ;
        RECT 143.000 14.100 143.400 14.200 ;
        RECT 142.600 13.800 143.400 14.100 ;
        RECT 144.600 13.800 145.600 14.200 ;
        RECT 145.900 14.100 146.600 14.500 ;
        RECT 147.000 14.400 147.400 15.200 ;
        RECT 147.800 14.400 148.200 15.200 ;
        RECT 151.800 15.100 152.200 15.200 ;
        RECT 152.600 15.100 153.000 15.200 ;
        RECT 149.700 14.800 153.000 15.100 ;
        RECT 149.700 14.700 150.100 14.800 ;
        RECT 150.500 14.200 150.900 14.300 ;
        RECT 154.200 14.200 154.500 15.800 ;
        RECT 157.400 15.600 157.800 19.900 ;
        RECT 155.700 15.300 157.800 15.600 ;
        RECT 158.200 15.700 158.600 19.900 ;
        RECT 160.400 18.200 160.800 19.900 ;
        RECT 159.800 17.900 160.800 18.200 ;
        RECT 162.600 17.900 163.000 19.900 ;
        RECT 164.700 17.900 165.300 19.900 ;
        RECT 159.800 17.500 160.200 17.900 ;
        RECT 162.600 17.600 162.900 17.900 ;
        RECT 161.500 17.300 163.300 17.600 ;
        RECT 164.600 17.500 165.000 17.900 ;
        RECT 161.500 17.200 161.900 17.300 ;
        RECT 162.900 17.200 163.300 17.300 ;
        RECT 167.000 17.100 167.400 19.900 ;
        RECT 167.800 17.100 168.200 17.200 ;
        RECT 159.800 16.500 160.200 16.600 ;
        RECT 162.100 16.500 162.500 16.600 ;
        RECT 159.800 16.200 162.500 16.500 ;
        RECT 162.800 16.500 163.900 16.800 ;
        RECT 162.800 15.900 163.100 16.500 ;
        RECT 163.500 16.400 163.900 16.500 ;
        RECT 164.700 16.600 165.400 17.000 ;
        RECT 167.000 16.800 168.200 17.100 ;
        RECT 164.700 16.100 165.000 16.600 ;
        RECT 160.700 15.700 163.100 15.900 ;
        RECT 158.200 15.600 163.100 15.700 ;
        RECT 163.800 15.800 165.000 16.100 ;
        RECT 158.200 15.500 161.100 15.600 ;
        RECT 158.200 15.400 161.000 15.500 ;
        RECT 155.700 15.200 156.100 15.300 ;
        RECT 156.500 14.900 156.900 15.000 ;
        RECT 155.000 14.600 156.900 14.900 ;
        RECT 155.000 14.500 155.400 14.600 ;
        RECT 140.700 13.100 141.000 13.800 ;
        RECT 142.600 13.600 143.000 13.800 ;
        RECT 145.300 13.500 145.600 13.800 ;
        RECT 146.100 13.900 146.600 14.100 ;
        RECT 149.000 13.900 154.500 14.200 ;
        RECT 146.100 13.600 148.200 13.900 ;
        RECT 149.000 13.800 149.800 13.900 ;
        RECT 145.300 13.300 145.700 13.500 ;
        RECT 141.500 13.100 143.300 13.300 ;
        RECT 137.400 12.800 138.300 13.100 ;
        RECT 135.800 11.500 136.200 12.500 ;
        RECT 137.900 11.100 138.300 12.800 ;
        RECT 140.600 11.100 141.000 13.100 ;
        RECT 141.400 13.000 143.400 13.100 ;
        RECT 145.300 13.000 146.100 13.300 ;
        RECT 141.400 11.100 141.800 13.000 ;
        RECT 143.000 11.100 143.400 13.000 ;
        RECT 145.700 11.500 146.100 13.000 ;
        RECT 147.900 12.500 148.200 13.600 ;
        RECT 147.800 11.500 148.200 12.500 ;
        RECT 148.600 11.100 149.000 13.500 ;
        RECT 151.100 12.800 151.400 13.900 ;
        RECT 153.900 13.800 154.300 13.900 ;
        RECT 157.400 13.600 157.800 15.300 ;
        RECT 161.400 15.100 161.800 15.200 ;
        RECT 159.300 14.800 161.800 15.100 ;
        RECT 159.300 14.700 159.700 14.800 ;
        RECT 160.100 14.200 160.500 14.300 ;
        RECT 163.800 14.200 164.100 15.800 ;
        RECT 167.000 15.600 167.400 16.800 ;
        RECT 165.300 15.300 167.400 15.600 ;
        RECT 165.300 15.200 165.700 15.300 ;
        RECT 166.100 14.900 166.500 15.000 ;
        RECT 164.600 14.600 166.500 14.900 ;
        RECT 164.600 14.500 165.000 14.600 ;
        RECT 158.600 13.900 164.100 14.200 ;
        RECT 158.600 13.800 159.400 13.900 ;
        RECT 160.600 13.800 161.000 13.900 ;
        RECT 163.500 13.800 163.900 13.900 ;
        RECT 155.900 13.300 157.800 13.600 ;
        RECT 155.900 13.200 156.300 13.300 ;
        RECT 150.200 12.100 150.600 12.500 ;
        RECT 151.000 12.400 151.400 12.800 ;
        RECT 151.900 12.700 152.300 12.800 ;
        RECT 151.900 12.400 153.300 12.700 ;
        RECT 153.000 12.100 153.300 12.400 ;
        RECT 155.000 12.100 155.400 12.500 ;
        RECT 150.200 11.800 151.200 12.100 ;
        RECT 150.800 11.100 151.200 11.800 ;
        RECT 153.000 11.100 153.400 12.100 ;
        RECT 155.000 11.800 155.700 12.100 ;
        RECT 155.100 11.100 155.700 11.800 ;
        RECT 157.400 11.100 157.800 13.300 ;
        RECT 158.200 11.100 158.600 13.500 ;
        RECT 160.700 12.800 161.000 13.800 ;
        RECT 167.000 13.600 167.400 15.300 ;
        RECT 168.600 15.100 169.000 19.900 ;
        RECT 170.600 16.800 171.000 17.200 ;
        RECT 169.400 15.800 169.800 16.600 ;
        RECT 170.600 16.200 170.900 16.800 ;
        RECT 171.300 16.200 171.700 19.900 ;
        RECT 170.200 15.900 170.900 16.200 ;
        RECT 171.200 15.900 171.700 16.200 ;
        RECT 170.200 15.800 170.600 15.900 ;
        RECT 170.200 15.100 170.500 15.800 ;
        RECT 168.600 14.800 170.500 15.100 ;
        RECT 165.500 13.300 167.400 13.600 ;
        RECT 167.800 13.400 168.200 14.200 ;
        RECT 165.500 13.200 165.900 13.300 ;
        RECT 159.800 12.100 160.200 12.500 ;
        RECT 160.600 12.400 161.000 12.800 ;
        RECT 161.500 12.700 161.900 12.800 ;
        RECT 161.500 12.400 162.900 12.700 ;
        RECT 162.600 12.100 162.900 12.400 ;
        RECT 164.600 12.100 165.000 12.500 ;
        RECT 159.800 11.800 160.800 12.100 ;
        RECT 160.400 11.100 160.800 11.800 ;
        RECT 162.600 11.100 163.000 12.100 ;
        RECT 164.600 11.800 165.300 12.100 ;
        RECT 164.700 11.100 165.300 11.800 ;
        RECT 167.000 11.100 167.400 13.300 ;
        RECT 168.600 13.100 169.000 14.800 ;
        RECT 171.200 14.200 171.500 15.900 ;
        RECT 173.400 15.700 173.800 19.900 ;
        RECT 175.600 18.200 176.000 19.900 ;
        RECT 175.000 17.900 176.000 18.200 ;
        RECT 177.800 17.900 178.200 19.900 ;
        RECT 179.900 17.900 180.500 19.900 ;
        RECT 175.000 17.500 175.400 17.900 ;
        RECT 177.800 17.600 178.100 17.900 ;
        RECT 176.700 17.300 178.500 17.600 ;
        RECT 179.800 17.500 180.200 17.900 ;
        RECT 176.700 17.200 177.100 17.300 ;
        RECT 178.100 17.200 178.500 17.300 ;
        RECT 180.300 17.000 181.000 17.200 ;
        RECT 179.900 16.800 181.000 17.000 ;
        RECT 175.000 16.500 175.400 16.600 ;
        RECT 177.300 16.500 177.700 16.600 ;
        RECT 175.000 16.200 177.700 16.500 ;
        RECT 178.000 16.500 179.100 16.800 ;
        RECT 178.000 15.900 178.300 16.500 ;
        RECT 178.700 16.400 179.100 16.500 ;
        RECT 179.900 16.600 180.600 16.800 ;
        RECT 179.900 16.100 180.200 16.600 ;
        RECT 175.900 15.700 178.300 15.900 ;
        RECT 173.400 15.600 178.300 15.700 ;
        RECT 179.000 15.800 180.200 16.100 ;
        RECT 173.400 15.500 176.300 15.600 ;
        RECT 173.400 15.400 176.200 15.500 ;
        RECT 171.800 15.100 172.200 15.200 ;
        RECT 172.600 15.100 173.000 15.200 ;
        RECT 176.600 15.100 177.000 15.200 ;
        RECT 171.800 14.800 173.000 15.100 ;
        RECT 174.500 14.800 177.000 15.100 ;
        RECT 171.800 14.400 172.200 14.800 ;
        RECT 174.500 14.700 174.900 14.800 ;
        RECT 175.300 14.200 175.700 14.300 ;
        RECT 179.000 14.200 179.300 15.800 ;
        RECT 182.200 15.600 182.600 19.900 ;
        RECT 180.500 15.300 182.600 15.600 ;
        RECT 180.500 15.200 180.900 15.300 ;
        RECT 181.300 14.900 181.700 15.000 ;
        RECT 179.800 14.600 181.700 14.900 ;
        RECT 179.800 14.500 180.200 14.600 ;
        RECT 169.400 14.100 169.800 14.200 ;
        RECT 170.200 14.100 171.500 14.200 ;
        RECT 172.600 14.100 173.000 14.200 ;
        RECT 169.400 13.800 171.500 14.100 ;
        RECT 172.200 13.800 173.000 14.100 ;
        RECT 173.800 13.900 179.300 14.200 ;
        RECT 173.800 13.800 174.600 13.900 ;
        RECT 170.300 13.100 170.600 13.800 ;
        RECT 172.200 13.600 172.600 13.800 ;
        RECT 171.100 13.100 172.900 13.300 ;
        RECT 168.600 12.800 169.500 13.100 ;
        RECT 169.100 11.100 169.500 12.800 ;
        RECT 170.200 11.100 170.600 13.100 ;
        RECT 171.000 13.000 173.000 13.100 ;
        RECT 171.000 11.100 171.400 13.000 ;
        RECT 172.600 11.100 173.000 13.000 ;
        RECT 173.400 11.100 173.800 13.500 ;
        RECT 175.900 12.800 176.200 13.900 ;
        RECT 178.700 13.800 179.100 13.900 ;
        RECT 182.200 13.600 182.600 15.300 ;
        RECT 180.700 13.300 182.600 13.600 ;
        RECT 180.700 13.200 181.100 13.300 ;
        RECT 175.000 12.100 175.400 12.500 ;
        RECT 175.800 12.400 176.200 12.800 ;
        RECT 176.700 12.700 177.100 12.800 ;
        RECT 176.700 12.400 178.100 12.700 ;
        RECT 177.800 12.100 178.100 12.400 ;
        RECT 179.800 12.100 180.200 12.500 ;
        RECT 175.000 11.800 176.000 12.100 ;
        RECT 175.600 11.100 176.000 11.800 ;
        RECT 177.800 11.100 178.200 12.100 ;
        RECT 179.800 11.800 180.500 12.100 ;
        RECT 179.900 11.100 180.500 11.800 ;
        RECT 182.200 11.100 182.600 13.300 ;
        RECT 183.800 11.100 184.200 19.900 ;
        RECT 186.700 19.200 187.100 19.900 ;
        RECT 186.700 18.800 187.400 19.200 ;
        RECT 186.700 16.300 187.100 18.800 ;
        RECT 186.200 15.900 187.100 16.300 ;
        RECT 186.300 14.200 186.600 15.900 ;
        RECT 187.000 14.800 187.400 15.600 ;
        RECT 184.600 14.100 185.000 14.200 ;
        RECT 184.600 13.800 185.700 14.100 ;
        RECT 186.200 13.800 186.600 14.200 ;
        RECT 184.600 13.400 185.000 13.800 ;
        RECT 185.400 13.200 185.700 13.800 ;
        RECT 185.400 12.400 185.800 13.200 ;
        RECT 186.300 12.100 186.600 13.800 ;
        RECT 186.200 11.100 186.600 12.100 ;
        RECT 188.600 11.100 189.000 19.900 ;
        RECT 191.800 15.600 192.200 19.900 ;
        RECT 193.900 17.900 194.500 19.900 ;
        RECT 196.200 17.900 196.600 19.900 ;
        RECT 198.400 18.200 198.800 19.900 ;
        RECT 198.400 17.900 199.400 18.200 ;
        RECT 194.200 17.500 194.600 17.900 ;
        RECT 196.300 17.600 196.600 17.900 ;
        RECT 195.900 17.300 197.700 17.600 ;
        RECT 199.000 17.500 199.400 17.900 ;
        RECT 195.900 17.200 196.300 17.300 ;
        RECT 197.300 17.200 197.700 17.300 ;
        RECT 193.400 17.000 194.100 17.200 ;
        RECT 193.400 16.800 194.500 17.000 ;
        RECT 193.800 16.600 194.500 16.800 ;
        RECT 194.200 16.100 194.500 16.600 ;
        RECT 195.300 16.500 196.400 16.800 ;
        RECT 195.300 16.400 195.700 16.500 ;
        RECT 194.200 15.800 195.400 16.100 ;
        RECT 191.800 15.300 193.900 15.600 ;
        RECT 189.400 14.100 189.800 14.200 ;
        RECT 191.800 14.100 192.200 15.300 ;
        RECT 193.500 15.200 193.900 15.300 ;
        RECT 192.700 14.900 193.100 15.000 ;
        RECT 192.700 14.600 194.600 14.900 ;
        RECT 194.200 14.500 194.600 14.600 ;
        RECT 189.400 13.800 192.200 14.100 ;
        RECT 195.100 14.200 195.400 15.800 ;
        RECT 196.100 15.900 196.400 16.500 ;
        RECT 196.700 16.500 197.100 16.600 ;
        RECT 199.000 16.500 199.400 16.600 ;
        RECT 196.700 16.200 199.400 16.500 ;
        RECT 196.100 15.700 198.500 15.900 ;
        RECT 200.600 15.700 201.000 19.900 ;
        RECT 196.100 15.600 201.000 15.700 ;
        RECT 198.100 15.500 201.000 15.600 ;
        RECT 201.400 17.500 201.800 19.500 ;
        RECT 203.500 19.200 203.900 19.900 ;
        RECT 203.500 18.800 204.200 19.200 ;
        RECT 201.400 15.800 201.700 17.500 ;
        RECT 203.500 16.400 203.900 18.800 ;
        RECT 203.500 16.100 204.300 16.400 ;
        RECT 201.400 15.500 203.300 15.800 ;
        RECT 198.200 15.400 201.000 15.500 ;
        RECT 195.800 15.100 196.200 15.200 ;
        RECT 197.400 15.100 197.800 15.200 ;
        RECT 195.800 14.800 199.900 15.100 ;
        RECT 199.500 14.700 199.900 14.800 ;
        RECT 201.400 14.400 201.800 15.200 ;
        RECT 202.200 14.400 202.600 15.200 ;
        RECT 203.000 14.500 203.300 15.500 ;
        RECT 198.700 14.200 199.100 14.300 ;
        RECT 195.100 13.900 200.600 14.200 ;
        RECT 203.000 14.100 203.700 14.500 ;
        RECT 204.000 14.200 204.300 16.100 ;
        RECT 204.600 15.100 205.000 15.600 ;
        RECT 207.000 15.100 207.400 19.900 ;
        RECT 209.000 16.800 209.400 17.200 ;
        RECT 207.800 15.800 208.200 16.600 ;
        RECT 209.000 16.200 209.300 16.800 ;
        RECT 209.700 16.200 210.100 19.900 ;
        RECT 208.600 15.900 209.300 16.200 ;
        RECT 209.600 15.900 210.100 16.200 ;
        RECT 213.100 16.200 213.500 19.900 ;
        RECT 213.800 16.800 214.200 17.200 ;
        RECT 213.900 16.200 214.200 16.800 ;
        RECT 213.100 15.900 213.600 16.200 ;
        RECT 213.900 15.900 214.600 16.200 ;
        RECT 208.600 15.800 209.000 15.900 ;
        RECT 208.600 15.100 208.900 15.800 ;
        RECT 204.600 14.800 206.500 15.100 ;
        RECT 206.200 14.200 206.500 14.800 ;
        RECT 207.000 14.800 208.900 15.100 ;
        RECT 203.000 13.900 203.500 14.100 ;
        RECT 195.300 13.800 195.700 13.900 ;
        RECT 189.400 13.400 189.800 13.800 ;
        RECT 191.800 13.600 192.200 13.800 ;
        RECT 191.800 13.300 193.700 13.600 ;
        RECT 191.800 11.100 192.200 13.300 ;
        RECT 193.300 13.200 193.700 13.300 ;
        RECT 198.200 13.200 198.500 13.900 ;
        RECT 199.800 13.800 200.600 13.900 ;
        RECT 201.400 13.600 203.500 13.900 ;
        RECT 204.000 13.800 205.000 14.200 ;
        RECT 197.300 12.700 197.700 12.800 ;
        RECT 194.200 12.100 194.600 12.500 ;
        RECT 196.300 12.400 197.700 12.700 ;
        RECT 198.200 12.400 198.600 13.200 ;
        RECT 196.300 12.100 196.600 12.400 ;
        RECT 199.000 12.100 199.400 12.500 ;
        RECT 193.900 11.800 194.600 12.100 ;
        RECT 193.900 11.100 194.500 11.800 ;
        RECT 196.200 11.100 196.600 12.100 ;
        RECT 198.400 11.800 199.400 12.100 ;
        RECT 198.400 11.100 198.800 11.800 ;
        RECT 200.600 11.100 201.000 13.500 ;
        RECT 201.400 12.500 201.700 13.600 ;
        RECT 204.000 13.500 204.300 13.800 ;
        RECT 203.900 13.300 204.300 13.500 ;
        RECT 206.200 13.400 206.600 14.200 ;
        RECT 203.500 13.000 204.300 13.300 ;
        RECT 207.000 13.100 207.400 14.800 ;
        RECT 209.600 14.200 209.900 15.900 ;
        RECT 210.200 14.400 210.600 15.200 ;
        RECT 212.600 14.400 213.000 15.200 ;
        RECT 213.300 14.200 213.600 15.900 ;
        RECT 214.200 15.800 214.600 15.900 ;
        RECT 215.000 15.800 215.400 16.600 ;
        RECT 214.200 15.100 214.500 15.800 ;
        RECT 215.800 15.100 216.200 19.900 ;
        RECT 218.200 15.600 218.600 19.900 ;
        RECT 219.800 15.600 220.200 19.900 ;
        RECT 221.400 15.600 221.800 19.900 ;
        RECT 223.000 15.600 223.400 19.900 ;
        RECT 218.200 15.200 219.100 15.600 ;
        RECT 219.800 15.200 220.900 15.600 ;
        RECT 221.400 15.200 222.500 15.600 ;
        RECT 223.000 15.200 224.200 15.600 ;
        RECT 214.200 14.800 216.200 15.100 ;
        RECT 208.600 13.800 209.900 14.200 ;
        RECT 211.000 14.100 211.400 14.200 ;
        RECT 211.800 14.100 212.200 14.200 ;
        RECT 210.600 13.800 212.600 14.100 ;
        RECT 213.300 13.800 214.600 14.200 ;
        RECT 208.700 13.100 209.000 13.800 ;
        RECT 210.600 13.600 211.000 13.800 ;
        RECT 212.200 13.600 212.600 13.800 ;
        RECT 209.500 13.100 211.300 13.300 ;
        RECT 211.900 13.100 213.700 13.300 ;
        RECT 214.200 13.100 214.500 13.800 ;
        RECT 215.800 13.100 216.200 14.800 ;
        RECT 218.700 14.500 219.100 15.200 ;
        RECT 220.500 14.500 220.900 15.200 ;
        RECT 222.100 14.500 222.500 15.200 ;
        RECT 216.600 13.400 217.000 14.200 ;
        RECT 218.700 14.100 220.000 14.500 ;
        RECT 220.500 14.100 221.700 14.500 ;
        RECT 222.100 14.100 223.400 14.500 ;
        RECT 218.700 13.800 219.100 14.100 ;
        RECT 220.500 13.800 220.900 14.100 ;
        RECT 222.100 13.800 222.500 14.100 ;
        RECT 223.800 13.800 224.200 15.200 ;
        RECT 225.400 15.100 225.800 19.900 ;
        RECT 228.100 19.200 228.500 19.900 ;
        RECT 228.100 18.800 229.000 19.200 ;
        RECT 227.400 16.800 227.800 17.200 ;
        RECT 226.200 15.800 226.600 16.600 ;
        RECT 227.400 16.200 227.700 16.800 ;
        RECT 228.100 16.200 228.500 18.800 ;
        RECT 227.000 15.900 227.700 16.200 ;
        RECT 228.000 15.900 228.500 16.200 ;
        RECT 227.000 15.800 227.400 15.900 ;
        RECT 227.000 15.100 227.300 15.800 ;
        RECT 225.400 14.800 227.300 15.100 ;
        RECT 218.200 13.400 219.100 13.800 ;
        RECT 219.800 13.400 220.900 13.800 ;
        RECT 221.400 13.400 222.500 13.800 ;
        RECT 223.000 13.400 224.200 13.800 ;
        RECT 224.600 13.400 225.000 14.200 ;
        RECT 201.400 11.500 201.800 12.500 ;
        RECT 203.500 11.500 203.900 13.000 ;
        RECT 207.000 12.800 207.900 13.100 ;
        RECT 207.500 11.100 207.900 12.800 ;
        RECT 208.600 11.100 209.000 13.100 ;
        RECT 209.400 13.000 211.400 13.100 ;
        RECT 209.400 11.100 209.800 13.000 ;
        RECT 211.000 11.100 211.400 13.000 ;
        RECT 211.800 13.000 213.800 13.100 ;
        RECT 211.800 11.100 212.200 13.000 ;
        RECT 213.400 11.100 213.800 13.000 ;
        RECT 214.200 11.100 214.600 13.100 ;
        RECT 215.300 12.800 216.200 13.100 ;
        RECT 215.300 11.100 215.700 12.800 ;
        RECT 218.200 11.100 218.600 13.400 ;
        RECT 219.800 11.100 220.200 13.400 ;
        RECT 221.400 11.100 221.800 13.400 ;
        RECT 223.000 11.100 223.400 13.400 ;
        RECT 225.400 13.100 225.800 14.800 ;
        RECT 228.000 14.200 228.300 15.900 ;
        RECT 228.600 14.400 229.000 15.200 ;
        RECT 227.000 13.800 228.300 14.200 ;
        RECT 229.400 14.100 229.800 14.200 ;
        RECT 229.000 13.800 229.800 14.100 ;
        RECT 227.100 13.100 227.400 13.800 ;
        RECT 229.000 13.600 229.400 13.800 ;
        RECT 227.900 13.100 229.700 13.300 ;
        RECT 225.400 12.800 226.300 13.100 ;
        RECT 225.900 11.100 226.300 12.800 ;
        RECT 227.000 11.100 227.400 13.100 ;
        RECT 227.800 13.000 229.800 13.100 ;
        RECT 227.800 11.100 228.200 13.000 ;
        RECT 229.400 11.100 229.800 13.000 ;
        RECT 0.600 7.900 1.000 9.900 ;
        RECT 1.400 8.000 1.800 9.900 ;
        RECT 3.000 8.000 3.400 9.900 ;
        RECT 1.400 7.900 3.400 8.000 ;
        RECT 4.100 8.200 4.500 9.900 ;
        RECT 7.000 8.200 7.400 9.900 ;
        RECT 4.100 7.900 5.000 8.200 ;
        RECT 0.700 7.200 1.000 7.900 ;
        RECT 1.500 7.700 3.300 7.900 ;
        RECT 2.600 7.200 3.000 7.400 ;
        RECT 0.600 6.800 1.900 7.200 ;
        RECT 2.600 7.100 3.400 7.200 ;
        RECT 3.800 7.100 4.200 7.200 ;
        RECT 2.600 6.900 4.200 7.100 ;
        RECT 3.000 6.800 4.200 6.900 ;
        RECT 0.600 5.100 1.000 5.200 ;
        RECT 1.600 5.100 1.900 6.800 ;
        RECT 2.200 6.100 2.600 6.600 ;
        RECT 4.600 6.100 5.000 7.900 ;
        RECT 6.900 7.900 7.400 8.200 ;
        RECT 5.400 6.800 5.800 7.600 ;
        RECT 6.900 7.200 7.200 7.900 ;
        RECT 8.600 7.600 9.000 9.900 ;
        RECT 7.700 7.300 9.000 7.600 ;
        RECT 10.200 7.600 10.600 9.900 ;
        RECT 11.800 7.600 12.200 9.900 ;
        RECT 13.700 9.200 14.100 9.900 ;
        RECT 13.700 8.800 14.600 9.200 ;
        RECT 13.700 8.200 14.100 8.800 ;
        RECT 13.700 7.900 14.600 8.200 ;
        RECT 6.900 7.100 7.400 7.200 ;
        RECT 6.200 6.800 7.400 7.100 ;
        RECT 6.200 6.200 6.500 6.800 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 2.200 5.800 4.100 6.100 ;
        RECT 3.800 5.200 4.100 5.800 ;
        RECT 4.600 5.800 5.800 6.100 ;
        RECT 6.200 5.800 6.600 6.200 ;
        RECT 0.600 4.800 1.300 5.100 ;
        RECT 1.600 4.800 2.100 5.100 ;
        RECT 1.000 4.200 1.300 4.800 ;
        RECT 1.000 3.800 1.400 4.200 ;
        RECT 1.700 1.100 2.100 4.800 ;
        RECT 3.800 4.400 4.200 5.200 ;
        RECT 4.600 1.100 5.000 5.800 ;
        RECT 6.900 5.100 7.200 6.800 ;
        RECT 7.700 6.500 8.000 7.300 ;
        RECT 10.200 7.200 12.200 7.600 ;
        RECT 7.500 6.100 8.000 6.500 ;
        RECT 7.700 5.100 8.000 6.100 ;
        RECT 8.500 6.200 8.900 6.600 ;
        RECT 8.500 6.100 9.000 6.200 ;
        RECT 8.500 5.800 10.600 6.100 ;
        RECT 11.800 5.800 12.200 7.200 ;
        RECT 10.200 5.400 12.200 5.800 ;
        RECT 6.900 4.600 7.400 5.100 ;
        RECT 7.700 4.800 9.000 5.100 ;
        RECT 7.000 1.100 7.400 4.600 ;
        RECT 8.600 1.100 9.000 4.800 ;
        RECT 10.200 1.100 10.600 5.400 ;
        RECT 11.800 1.100 12.200 5.400 ;
        RECT 13.400 4.400 13.800 5.200 ;
        RECT 14.200 1.100 14.600 7.900 ;
        RECT 16.600 7.600 17.000 9.900 ;
        RECT 18.200 7.600 18.600 9.900 ;
        RECT 15.000 6.800 15.400 7.600 ;
        RECT 16.600 7.200 18.600 7.600 ;
        RECT 19.800 7.600 20.200 9.900 ;
        RECT 21.400 8.200 21.800 9.900 ;
        RECT 21.400 7.900 21.900 8.200 ;
        RECT 19.800 7.300 21.100 7.600 ;
        RECT 18.200 5.800 18.600 7.200 ;
        RECT 19.900 6.200 20.300 6.600 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 19.800 6.100 20.300 6.200 ;
        RECT 19.000 5.800 20.300 6.100 ;
        RECT 20.800 6.500 21.100 7.300 ;
        RECT 21.600 7.200 21.900 7.900 ;
        RECT 23.800 7.600 24.200 9.900 ;
        RECT 25.400 7.600 25.800 9.900 ;
        RECT 27.000 7.600 27.400 9.900 ;
        RECT 28.600 7.600 29.000 9.900 ;
        RECT 23.800 7.200 24.700 7.600 ;
        RECT 25.400 7.200 26.500 7.600 ;
        RECT 27.000 7.200 28.100 7.600 ;
        RECT 28.600 7.200 29.800 7.600 ;
        RECT 30.200 7.500 30.600 9.900 ;
        RECT 32.400 9.200 32.800 9.900 ;
        RECT 31.800 8.900 32.800 9.200 ;
        RECT 34.600 8.900 35.000 9.900 ;
        RECT 36.700 9.200 37.300 9.900 ;
        RECT 36.600 8.900 37.300 9.200 ;
        RECT 31.800 8.500 32.200 8.900 ;
        RECT 34.600 8.600 34.900 8.900 ;
        RECT 32.600 8.200 33.000 8.600 ;
        RECT 33.500 8.300 34.900 8.600 ;
        RECT 36.600 8.500 37.000 8.900 ;
        RECT 33.500 8.200 33.900 8.300 ;
        RECT 21.400 6.800 21.900 7.200 ;
        RECT 20.800 6.100 21.300 6.500 ;
        RECT 16.600 5.400 18.600 5.800 ;
        RECT 16.600 1.100 17.000 5.400 ;
        RECT 18.200 1.100 18.600 5.400 ;
        RECT 20.800 5.100 21.100 6.100 ;
        RECT 21.600 5.100 21.900 6.800 ;
        RECT 24.300 6.900 24.700 7.200 ;
        RECT 26.100 6.900 26.500 7.200 ;
        RECT 27.700 6.900 28.100 7.200 ;
        RECT 24.300 6.500 25.600 6.900 ;
        RECT 26.100 6.500 27.300 6.900 ;
        RECT 27.700 6.500 29.000 6.900 ;
        RECT 24.300 5.800 24.700 6.500 ;
        RECT 26.100 5.800 26.500 6.500 ;
        RECT 27.700 5.800 28.100 6.500 ;
        RECT 29.400 5.800 29.800 7.200 ;
        RECT 30.600 7.100 31.400 7.200 ;
        RECT 32.700 7.100 33.000 8.200 ;
        RECT 37.500 7.700 37.900 7.800 ;
        RECT 39.000 7.700 39.400 9.900 ;
        RECT 39.800 9.100 40.200 9.200 ;
        RECT 41.700 9.100 42.100 9.900 ;
        RECT 39.800 8.800 42.100 9.100 ;
        RECT 41.700 8.200 42.100 8.800 ;
        RECT 45.100 8.200 45.500 9.900 ;
        RECT 41.700 7.900 42.600 8.200 ;
        RECT 37.500 7.400 39.400 7.700 ;
        RECT 35.500 7.100 36.200 7.200 ;
        RECT 30.600 6.800 36.200 7.100 ;
        RECT 32.100 6.700 32.500 6.800 ;
        RECT 31.300 6.200 31.700 6.300 ;
        RECT 31.300 6.100 33.800 6.200 ;
        RECT 35.000 6.100 35.400 6.200 ;
        RECT 31.300 5.900 35.400 6.100 ;
        RECT 33.400 5.800 35.400 5.900 ;
        RECT 19.800 4.800 21.100 5.100 ;
        RECT 19.800 1.100 20.200 4.800 ;
        RECT 21.400 4.600 21.900 5.100 ;
        RECT 23.800 5.400 24.700 5.800 ;
        RECT 25.400 5.400 26.500 5.800 ;
        RECT 27.000 5.400 28.100 5.800 ;
        RECT 28.600 5.400 29.800 5.800 ;
        RECT 30.200 5.500 33.000 5.600 ;
        RECT 30.200 5.400 33.100 5.500 ;
        RECT 21.400 1.100 21.800 4.600 ;
        RECT 23.800 1.100 24.200 5.400 ;
        RECT 25.400 1.100 25.800 5.400 ;
        RECT 27.000 1.100 27.400 5.400 ;
        RECT 28.600 1.100 29.000 5.400 ;
        RECT 30.200 5.300 35.100 5.400 ;
        RECT 30.200 1.100 30.600 5.300 ;
        RECT 32.700 5.100 35.100 5.300 ;
        RECT 31.800 4.500 34.500 4.800 ;
        RECT 31.800 4.400 32.200 4.500 ;
        RECT 34.100 4.400 34.500 4.500 ;
        RECT 34.800 4.500 35.100 5.100 ;
        RECT 35.800 5.200 36.100 6.800 ;
        RECT 36.600 6.400 37.000 6.500 ;
        RECT 36.600 6.100 38.500 6.400 ;
        RECT 38.100 6.000 38.500 6.100 ;
        RECT 37.300 5.700 37.700 5.800 ;
        RECT 39.000 5.700 39.400 7.400 ;
        RECT 37.300 5.400 39.400 5.700 ;
        RECT 35.800 4.900 37.000 5.200 ;
        RECT 35.500 4.500 35.900 4.600 ;
        RECT 34.800 4.200 35.900 4.500 ;
        RECT 36.700 4.400 37.000 4.900 ;
        RECT 36.700 4.000 37.400 4.400 ;
        RECT 33.500 3.700 33.900 3.800 ;
        RECT 34.900 3.700 35.300 3.800 ;
        RECT 31.800 3.100 32.200 3.500 ;
        RECT 33.500 3.400 35.300 3.700 ;
        RECT 34.600 3.100 34.900 3.400 ;
        RECT 36.600 3.100 37.000 3.500 ;
        RECT 31.800 2.800 32.800 3.100 ;
        RECT 32.400 1.100 32.800 2.800 ;
        RECT 34.600 1.100 35.000 3.100 ;
        RECT 36.700 1.100 37.300 3.100 ;
        RECT 39.000 1.100 39.400 5.400 ;
        RECT 41.400 4.400 41.800 5.200 ;
        RECT 42.200 1.100 42.600 7.900 ;
        RECT 44.600 7.900 45.500 8.200 ;
        RECT 46.200 7.900 46.600 9.900 ;
        RECT 47.000 8.000 47.400 9.900 ;
        RECT 48.600 8.000 49.000 9.900 ;
        RECT 47.000 7.900 49.000 8.000 ;
        RECT 43.000 6.800 43.400 7.600 ;
        RECT 43.800 6.800 44.200 7.600 ;
        RECT 44.600 6.100 45.000 7.900 ;
        RECT 46.300 7.200 46.600 7.900 ;
        RECT 47.100 7.700 48.900 7.900 ;
        RECT 49.400 7.700 49.800 9.900 ;
        RECT 51.500 9.200 52.100 9.900 ;
        RECT 51.500 8.900 52.200 9.200 ;
        RECT 53.800 8.900 54.200 9.900 ;
        RECT 56.000 9.200 56.400 9.900 ;
        RECT 56.000 8.900 57.000 9.200 ;
        RECT 51.800 8.500 52.200 8.900 ;
        RECT 53.900 8.600 54.200 8.900 ;
        RECT 53.900 8.300 55.300 8.600 ;
        RECT 54.900 8.200 55.300 8.300 ;
        RECT 55.800 8.200 56.200 8.600 ;
        RECT 56.600 8.500 57.000 8.900 ;
        RECT 50.900 7.700 51.300 7.800 ;
        RECT 49.400 7.400 51.300 7.700 ;
        RECT 48.200 7.200 48.600 7.400 ;
        RECT 46.200 6.800 47.500 7.200 ;
        RECT 48.200 6.900 49.000 7.200 ;
        RECT 48.600 6.800 49.000 6.900 ;
        RECT 44.600 5.800 46.500 6.100 ;
        RECT 44.600 1.100 45.000 5.800 ;
        RECT 46.200 5.200 46.500 5.800 ;
        RECT 45.400 4.400 45.800 5.200 ;
        RECT 46.200 5.100 46.600 5.200 ;
        RECT 47.200 5.100 47.500 6.800 ;
        RECT 47.800 5.800 48.200 6.600 ;
        RECT 49.400 5.700 49.800 7.400 ;
        RECT 52.900 7.100 53.300 7.200 ;
        RECT 55.800 7.100 56.100 8.200 ;
        RECT 58.200 7.500 58.600 9.900 ;
        RECT 59.000 7.500 59.400 9.900 ;
        RECT 61.200 9.200 61.600 9.900 ;
        RECT 60.600 8.900 61.600 9.200 ;
        RECT 63.400 8.900 63.800 9.900 ;
        RECT 65.500 9.200 66.100 9.900 ;
        RECT 65.400 8.900 66.100 9.200 ;
        RECT 60.600 8.500 61.000 8.900 ;
        RECT 63.400 8.600 63.700 8.900 ;
        RECT 61.400 8.200 61.800 8.600 ;
        RECT 62.300 8.300 63.700 8.600 ;
        RECT 65.400 8.500 65.800 8.900 ;
        RECT 62.300 8.200 62.700 8.300 ;
        RECT 57.400 7.100 58.200 7.200 ;
        RECT 59.400 7.100 60.200 7.200 ;
        RECT 61.500 7.100 61.800 8.200 ;
        RECT 64.600 7.800 65.000 8.200 ;
        RECT 64.600 7.200 64.900 7.800 ;
        RECT 66.300 7.700 66.700 7.800 ;
        RECT 67.800 7.700 68.200 9.900 ;
        RECT 66.300 7.400 68.200 7.700 ;
        RECT 68.600 7.500 69.000 9.900 ;
        RECT 70.800 9.200 71.200 9.900 ;
        RECT 70.200 8.900 71.200 9.200 ;
        RECT 73.000 8.900 73.400 9.900 ;
        RECT 75.100 9.200 75.700 9.900 ;
        RECT 75.000 8.900 75.700 9.200 ;
        RECT 70.200 8.500 70.600 8.900 ;
        RECT 73.000 8.600 73.300 8.900 ;
        RECT 71.000 8.200 71.400 8.600 ;
        RECT 71.900 8.300 73.300 8.600 ;
        RECT 75.000 8.500 75.400 8.900 ;
        RECT 71.900 8.200 72.300 8.300 ;
        RECT 64.300 7.100 64.900 7.200 ;
        RECT 52.700 6.800 64.900 7.100 ;
        RECT 51.800 6.400 52.200 6.500 ;
        RECT 50.300 6.100 52.200 6.400 ;
        RECT 52.700 6.200 53.000 6.800 ;
        RECT 56.300 6.700 56.700 6.800 ;
        RECT 60.900 6.700 61.300 6.800 ;
        RECT 55.800 6.200 56.200 6.300 ;
        RECT 57.100 6.200 57.500 6.300 ;
        RECT 50.300 6.000 50.700 6.100 ;
        RECT 52.600 5.800 53.000 6.200 ;
        RECT 55.000 5.900 57.500 6.200 ;
        RECT 60.100 6.200 60.500 6.300 ;
        RECT 60.100 5.900 62.600 6.200 ;
        RECT 55.000 5.800 55.400 5.900 ;
        RECT 62.200 5.800 62.600 5.900 ;
        RECT 51.100 5.700 51.500 5.800 ;
        RECT 49.400 5.400 51.500 5.700 ;
        RECT 46.200 4.800 46.900 5.100 ;
        RECT 47.200 4.800 47.700 5.100 ;
        RECT 46.600 4.200 46.900 4.800 ;
        RECT 46.600 3.800 47.000 4.200 ;
        RECT 47.300 1.100 47.700 4.800 ;
        RECT 49.400 1.100 49.800 5.400 ;
        RECT 52.700 5.200 53.000 5.800 ;
        RECT 55.800 5.500 58.600 5.600 ;
        RECT 55.700 5.400 58.600 5.500 ;
        RECT 51.800 4.900 53.000 5.200 ;
        RECT 53.700 5.300 58.600 5.400 ;
        RECT 53.700 5.100 56.100 5.300 ;
        RECT 51.800 4.400 52.100 4.900 ;
        RECT 51.400 4.000 52.100 4.400 ;
        RECT 52.900 4.500 53.300 4.600 ;
        RECT 53.700 4.500 54.000 5.100 ;
        RECT 52.900 4.200 54.000 4.500 ;
        RECT 54.300 4.500 57.000 4.800 ;
        RECT 54.300 4.400 54.700 4.500 ;
        RECT 56.600 4.400 57.000 4.500 ;
        RECT 53.500 3.700 53.900 3.800 ;
        RECT 54.900 3.700 55.300 3.800 ;
        RECT 51.800 3.100 52.200 3.500 ;
        RECT 53.500 3.400 55.300 3.700 ;
        RECT 53.900 3.100 54.200 3.400 ;
        RECT 56.600 3.100 57.000 3.500 ;
        RECT 51.500 1.100 52.100 3.100 ;
        RECT 53.800 1.100 54.200 3.100 ;
        RECT 56.000 2.800 57.000 3.100 ;
        RECT 56.000 1.100 56.400 2.800 ;
        RECT 58.200 1.100 58.600 5.300 ;
        RECT 59.000 5.500 61.800 5.600 ;
        RECT 59.000 5.400 61.900 5.500 ;
        RECT 59.000 5.300 63.900 5.400 ;
        RECT 59.000 1.100 59.400 5.300 ;
        RECT 61.500 5.100 63.900 5.300 ;
        RECT 60.600 4.500 63.300 4.800 ;
        RECT 60.600 4.400 61.000 4.500 ;
        RECT 62.900 4.400 63.300 4.500 ;
        RECT 63.600 4.500 63.900 5.100 ;
        RECT 64.600 5.200 64.900 6.800 ;
        RECT 65.400 6.400 65.800 6.500 ;
        RECT 65.400 6.100 67.300 6.400 ;
        RECT 66.900 6.000 67.300 6.100 ;
        RECT 66.100 5.700 66.500 5.800 ;
        RECT 67.800 5.700 68.200 7.400 ;
        RECT 69.000 7.100 69.800 7.200 ;
        RECT 71.100 7.100 71.400 8.200 ;
        RECT 75.900 7.700 76.300 7.800 ;
        RECT 77.400 7.700 77.800 9.900 ;
        RECT 78.300 8.200 78.700 8.600 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 79.000 7.900 79.400 9.900 ;
        RECT 75.900 7.400 77.800 7.700 ;
        RECT 71.800 7.100 72.200 7.200 ;
        RECT 73.900 7.100 74.300 7.200 ;
        RECT 69.000 6.800 74.500 7.100 ;
        RECT 70.500 6.700 70.900 6.800 ;
        RECT 69.700 6.200 70.100 6.300 ;
        RECT 69.700 6.100 72.200 6.200 ;
        RECT 72.600 6.100 73.000 6.200 ;
        RECT 69.700 5.900 73.000 6.100 ;
        RECT 71.800 5.800 73.000 5.900 ;
        RECT 66.100 5.400 68.200 5.700 ;
        RECT 64.600 4.900 65.800 5.200 ;
        RECT 64.300 4.500 64.700 4.600 ;
        RECT 63.600 4.200 64.700 4.500 ;
        RECT 65.500 4.400 65.800 4.900 ;
        RECT 65.500 4.000 66.200 4.400 ;
        RECT 62.300 3.700 62.700 3.800 ;
        RECT 63.700 3.700 64.100 3.800 ;
        RECT 60.600 3.100 61.000 3.500 ;
        RECT 62.300 3.400 64.100 3.700 ;
        RECT 63.400 3.100 63.700 3.400 ;
        RECT 65.400 3.100 65.800 3.500 ;
        RECT 60.600 2.800 61.600 3.100 ;
        RECT 61.200 1.100 61.600 2.800 ;
        RECT 63.400 1.100 63.800 3.100 ;
        RECT 65.500 1.100 66.100 3.100 ;
        RECT 67.800 1.100 68.200 5.400 ;
        RECT 68.600 5.500 71.400 5.600 ;
        RECT 68.600 5.400 71.500 5.500 ;
        RECT 68.600 5.300 73.500 5.400 ;
        RECT 68.600 1.100 69.000 5.300 ;
        RECT 71.100 5.100 73.500 5.300 ;
        RECT 70.200 4.500 72.900 4.800 ;
        RECT 70.200 4.400 70.600 4.500 ;
        RECT 72.500 4.400 72.900 4.500 ;
        RECT 73.200 4.500 73.500 5.100 ;
        RECT 74.200 5.200 74.500 6.800 ;
        RECT 75.000 6.400 75.400 6.500 ;
        RECT 75.000 6.100 76.900 6.400 ;
        RECT 76.500 6.000 76.900 6.100 ;
        RECT 75.700 5.700 76.100 5.800 ;
        RECT 77.400 5.700 77.800 7.400 ;
        RECT 78.200 6.100 78.600 6.200 ;
        RECT 79.100 6.100 79.400 7.900 ;
        RECT 83.000 7.900 83.400 9.900 ;
        RECT 85.400 8.900 85.800 9.900 ;
        RECT 87.800 8.900 88.200 9.900 ;
        RECT 83.700 8.200 84.100 8.600 ;
        RECT 83.800 8.100 84.200 8.200 ;
        RECT 85.400 8.100 85.700 8.900 ;
        RECT 79.800 6.400 80.200 7.200 ;
        RECT 82.200 6.400 82.600 7.200 ;
        RECT 78.200 5.800 79.400 6.100 ;
        RECT 83.000 6.200 83.300 7.900 ;
        RECT 83.800 7.800 85.700 8.100 ;
        RECT 85.400 7.200 85.700 7.800 ;
        RECT 87.900 7.200 88.200 8.900 ;
        RECT 91.000 8.000 91.400 9.900 ;
        RECT 92.600 8.000 93.000 9.900 ;
        RECT 91.000 7.900 93.000 8.000 ;
        RECT 93.400 7.900 93.800 9.900 ;
        RECT 94.500 8.200 94.900 9.900 ;
        RECT 94.500 7.900 95.400 8.200 ;
        RECT 91.100 7.700 92.900 7.900 ;
        RECT 91.400 7.200 91.800 7.400 ;
        RECT 93.400 7.200 93.700 7.900 ;
        RECT 85.400 6.800 85.800 7.200 ;
        RECT 87.800 7.100 88.200 7.200 ;
        RECT 87.000 6.800 88.200 7.100 ;
        RECT 90.200 7.100 90.600 7.200 ;
        RECT 91.000 7.100 91.800 7.200 ;
        RECT 90.200 6.900 91.800 7.100 ;
        RECT 90.200 6.800 91.400 6.900 ;
        RECT 92.500 6.800 93.800 7.200 ;
        RECT 83.000 6.100 83.400 6.200 ;
        RECT 83.800 6.100 84.200 6.200 ;
        RECT 83.000 5.800 84.200 6.100 ;
        RECT 75.700 5.400 77.800 5.700 ;
        RECT 74.200 4.900 75.400 5.200 ;
        RECT 73.900 4.500 74.300 4.600 ;
        RECT 73.200 4.200 74.300 4.500 ;
        RECT 75.100 4.400 75.400 4.900 ;
        RECT 75.100 4.000 75.800 4.400 ;
        RECT 71.900 3.700 72.300 3.800 ;
        RECT 73.300 3.700 73.700 3.800 ;
        RECT 70.200 3.100 70.600 3.500 ;
        RECT 71.900 3.400 73.700 3.700 ;
        RECT 73.000 3.100 73.300 3.400 ;
        RECT 75.000 3.100 75.400 3.500 ;
        RECT 70.200 2.800 71.200 3.100 ;
        RECT 70.800 1.100 71.200 2.800 ;
        RECT 73.000 1.100 73.400 3.100 ;
        RECT 75.100 1.100 75.700 3.100 ;
        RECT 77.400 1.100 77.800 5.400 ;
        RECT 78.300 5.200 78.600 5.800 ;
        RECT 78.200 1.100 78.600 5.200 ;
        RECT 83.800 5.100 84.100 5.800 ;
        RECT 85.400 5.100 85.700 6.800 ;
        RECT 87.000 6.200 87.300 6.800 ;
        RECT 87.000 5.800 87.400 6.200 ;
        RECT 87.900 5.100 88.200 6.800 ;
        RECT 91.800 5.800 92.200 6.600 ;
        RECT 92.500 5.100 92.800 6.800 ;
        RECT 95.000 6.100 95.400 7.900 ;
        RECT 95.800 6.800 96.200 7.600 ;
        RECT 96.600 7.500 97.000 9.900 ;
        RECT 98.800 9.200 99.200 9.900 ;
        RECT 98.200 8.900 99.200 9.200 ;
        RECT 101.000 8.900 101.400 9.900 ;
        RECT 103.100 9.200 103.700 9.900 ;
        RECT 103.000 8.900 103.700 9.200 ;
        RECT 98.200 8.500 98.600 8.900 ;
        RECT 101.000 8.600 101.300 8.900 ;
        RECT 99.000 8.200 99.400 8.600 ;
        RECT 99.900 8.300 101.300 8.600 ;
        RECT 103.000 8.500 103.400 8.900 ;
        RECT 99.900 8.200 100.300 8.300 ;
        RECT 97.000 7.100 97.800 7.200 ;
        RECT 99.100 7.100 99.400 8.200 ;
        RECT 103.900 7.700 104.300 7.800 ;
        RECT 105.400 7.700 105.800 9.900 ;
        RECT 103.900 7.400 105.800 7.700 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 101.900 7.100 102.300 7.200 ;
        RECT 97.000 6.800 102.500 7.100 ;
        RECT 98.500 6.700 98.900 6.800 ;
        RECT 93.400 5.800 95.400 6.100 ;
        RECT 97.700 6.200 98.100 6.300 ;
        RECT 99.000 6.200 99.400 6.300 ;
        RECT 97.700 5.900 100.200 6.200 ;
        RECT 99.800 5.800 100.200 5.900 ;
        RECT 93.400 5.200 93.700 5.800 ;
        RECT 93.400 5.100 93.800 5.200 ;
        RECT 79.000 4.800 81.000 5.100 ;
        RECT 79.000 1.100 79.400 4.800 ;
        RECT 80.600 1.100 81.000 4.800 ;
        RECT 81.400 4.800 83.400 5.100 ;
        RECT 81.400 1.100 81.800 4.800 ;
        RECT 83.000 1.100 83.400 4.800 ;
        RECT 83.800 1.100 84.200 5.100 ;
        RECT 84.900 4.700 85.800 5.100 ;
        RECT 87.800 4.700 88.700 5.100 ;
        RECT 84.900 1.100 85.300 4.700 ;
        RECT 88.300 1.100 88.700 4.700 ;
        RECT 92.300 4.800 92.800 5.100 ;
        RECT 93.100 4.800 93.800 5.100 ;
        RECT 92.300 1.100 92.700 4.800 ;
        RECT 93.100 4.200 93.400 4.800 ;
        RECT 94.200 4.400 94.600 5.200 ;
        RECT 93.000 3.800 93.400 4.200 ;
        RECT 95.000 1.100 95.400 5.800 ;
        RECT 96.600 5.500 99.400 5.600 ;
        RECT 96.600 5.400 99.500 5.500 ;
        RECT 96.600 5.300 101.500 5.400 ;
        RECT 96.600 1.100 97.000 5.300 ;
        RECT 99.100 5.100 101.500 5.300 ;
        RECT 98.200 4.500 100.900 4.800 ;
        RECT 98.200 4.400 98.600 4.500 ;
        RECT 100.500 4.400 100.900 4.500 ;
        RECT 101.200 4.500 101.500 5.100 ;
        RECT 102.200 5.200 102.500 6.800 ;
        RECT 103.000 6.400 103.400 6.500 ;
        RECT 103.000 6.100 104.900 6.400 ;
        RECT 104.500 6.000 104.900 6.100 ;
        RECT 103.700 5.700 104.100 5.800 ;
        RECT 105.400 5.700 105.800 7.400 ;
        RECT 103.700 5.400 105.800 5.700 ;
        RECT 102.200 4.900 103.400 5.200 ;
        RECT 101.900 4.500 102.300 4.600 ;
        RECT 101.200 4.200 102.300 4.500 ;
        RECT 103.100 4.400 103.400 4.900 ;
        RECT 103.100 4.000 103.800 4.400 ;
        RECT 99.900 3.700 100.300 3.800 ;
        RECT 101.300 3.700 101.700 3.800 ;
        RECT 98.200 3.100 98.600 3.500 ;
        RECT 99.900 3.400 101.700 3.700 ;
        RECT 101.000 3.100 101.300 3.400 ;
        RECT 103.000 3.100 103.400 3.500 ;
        RECT 98.200 2.800 99.200 3.100 ;
        RECT 98.800 1.100 99.200 2.800 ;
        RECT 101.000 1.100 101.400 3.100 ;
        RECT 103.100 1.100 103.700 3.100 ;
        RECT 105.400 1.100 105.800 5.400 ;
        RECT 107.000 7.600 107.400 9.900 ;
        RECT 108.600 7.600 109.000 9.900 ;
        RECT 107.000 7.200 109.000 7.600 ;
        RECT 110.200 7.500 110.600 9.900 ;
        RECT 112.400 9.200 112.800 9.900 ;
        RECT 111.800 8.900 112.800 9.200 ;
        RECT 114.600 8.900 115.000 9.900 ;
        RECT 116.700 9.200 117.300 9.900 ;
        RECT 116.600 8.900 117.300 9.200 ;
        RECT 111.800 8.500 112.200 8.900 ;
        RECT 114.600 8.600 114.900 8.900 ;
        RECT 112.600 8.200 113.000 8.600 ;
        RECT 113.500 8.300 114.900 8.600 ;
        RECT 116.600 8.500 117.000 8.900 ;
        RECT 113.500 8.200 113.900 8.300 ;
        RECT 107.000 5.800 107.400 7.200 ;
        RECT 110.600 7.100 111.400 7.200 ;
        RECT 112.700 7.100 113.000 8.200 ;
        RECT 117.500 7.700 117.900 7.800 ;
        RECT 119.000 7.700 119.400 9.900 ;
        RECT 117.500 7.400 119.400 7.700 ;
        RECT 119.800 7.500 120.200 9.900 ;
        RECT 122.000 9.200 122.400 9.900 ;
        RECT 121.400 8.900 122.400 9.200 ;
        RECT 124.200 8.900 124.600 9.900 ;
        RECT 126.300 9.200 126.900 9.900 ;
        RECT 126.200 8.900 126.900 9.200 ;
        RECT 121.400 8.500 121.800 8.900 ;
        RECT 124.200 8.600 124.500 8.900 ;
        RECT 122.200 7.800 122.600 8.600 ;
        RECT 123.100 8.300 124.500 8.600 ;
        RECT 126.200 8.500 126.600 8.900 ;
        RECT 123.100 8.200 123.500 8.300 ;
        RECT 114.200 7.100 114.600 7.200 ;
        RECT 115.500 7.100 115.900 7.200 ;
        RECT 110.600 6.800 116.100 7.100 ;
        RECT 112.100 6.700 112.500 6.800 ;
        RECT 111.300 6.200 111.700 6.300 ;
        RECT 111.300 6.100 113.800 6.200 ;
        RECT 114.200 6.100 114.600 6.200 ;
        RECT 111.300 5.900 114.600 6.100 ;
        RECT 113.400 5.800 114.600 5.900 ;
        RECT 107.000 5.400 109.000 5.800 ;
        RECT 107.000 1.100 107.400 5.400 ;
        RECT 108.600 1.100 109.000 5.400 ;
        RECT 110.200 5.500 113.000 5.600 ;
        RECT 110.200 5.400 113.100 5.500 ;
        RECT 110.200 5.300 115.100 5.400 ;
        RECT 110.200 1.100 110.600 5.300 ;
        RECT 112.700 5.100 115.100 5.300 ;
        RECT 111.800 4.500 114.500 4.800 ;
        RECT 111.800 4.400 112.200 4.500 ;
        RECT 114.100 4.400 114.500 4.500 ;
        RECT 114.800 4.500 115.100 5.100 ;
        RECT 115.800 5.200 116.100 6.800 ;
        RECT 116.600 6.400 117.000 6.500 ;
        RECT 116.600 6.100 118.500 6.400 ;
        RECT 118.100 6.000 118.500 6.100 ;
        RECT 117.300 5.700 117.700 5.800 ;
        RECT 119.000 5.700 119.400 7.400 ;
        RECT 120.200 7.100 121.000 7.200 ;
        RECT 122.300 7.100 122.600 7.800 ;
        RECT 127.100 7.700 127.500 7.800 ;
        RECT 128.600 7.700 129.000 9.900 ;
        RECT 129.400 7.900 129.800 9.900 ;
        RECT 130.200 8.000 130.600 9.900 ;
        RECT 131.800 8.000 132.200 9.900 ;
        RECT 130.200 7.900 132.200 8.000 ;
        RECT 127.100 7.400 129.000 7.700 ;
        RECT 123.800 7.100 124.200 7.200 ;
        RECT 125.100 7.100 125.500 7.200 ;
        RECT 120.200 6.800 125.700 7.100 ;
        RECT 121.700 6.700 122.100 6.800 ;
        RECT 120.900 6.200 121.300 6.300 ;
        RECT 120.900 5.900 123.400 6.200 ;
        RECT 123.000 5.800 123.400 5.900 ;
        RECT 117.300 5.400 119.400 5.700 ;
        RECT 115.800 4.900 117.000 5.200 ;
        RECT 115.500 4.500 115.900 4.600 ;
        RECT 114.800 4.200 115.900 4.500 ;
        RECT 116.700 4.400 117.000 4.900 ;
        RECT 116.700 4.000 117.400 4.400 ;
        RECT 113.500 3.700 113.900 3.800 ;
        RECT 114.900 3.700 115.300 3.800 ;
        RECT 111.800 3.100 112.200 3.500 ;
        RECT 113.500 3.400 115.300 3.700 ;
        RECT 114.600 3.100 114.900 3.400 ;
        RECT 116.600 3.100 117.000 3.500 ;
        RECT 111.800 2.800 112.800 3.100 ;
        RECT 112.400 1.100 112.800 2.800 ;
        RECT 114.600 1.100 115.000 3.100 ;
        RECT 116.700 1.100 117.300 3.100 ;
        RECT 119.000 1.100 119.400 5.400 ;
        RECT 119.800 5.500 122.600 5.600 ;
        RECT 119.800 5.400 122.700 5.500 ;
        RECT 119.800 5.300 124.700 5.400 ;
        RECT 119.800 1.100 120.200 5.300 ;
        RECT 122.300 5.100 124.700 5.300 ;
        RECT 121.400 4.500 124.100 4.800 ;
        RECT 121.400 4.400 121.800 4.500 ;
        RECT 123.700 4.400 124.100 4.500 ;
        RECT 124.400 4.500 124.700 5.100 ;
        RECT 125.400 5.200 125.700 6.800 ;
        RECT 126.200 6.400 126.600 6.500 ;
        RECT 126.200 6.100 128.100 6.400 ;
        RECT 127.700 6.000 128.100 6.100 ;
        RECT 126.900 5.700 127.300 5.800 ;
        RECT 128.600 5.700 129.000 7.400 ;
        RECT 129.500 7.200 129.800 7.900 ;
        RECT 130.300 7.700 132.100 7.900 ;
        RECT 132.600 7.700 133.000 9.900 ;
        RECT 134.700 9.200 135.300 9.900 ;
        RECT 134.700 8.900 135.400 9.200 ;
        RECT 137.000 8.900 137.400 9.900 ;
        RECT 139.200 9.200 139.600 9.900 ;
        RECT 139.200 8.900 140.200 9.200 ;
        RECT 135.000 8.500 135.400 8.900 ;
        RECT 137.100 8.600 137.400 8.900 ;
        RECT 137.100 8.300 138.500 8.600 ;
        RECT 138.100 8.200 138.500 8.300 ;
        RECT 139.000 8.200 139.400 8.600 ;
        RECT 139.800 8.500 140.200 8.900 ;
        RECT 134.100 7.700 134.500 7.800 ;
        RECT 132.600 7.400 134.500 7.700 ;
        RECT 131.400 7.200 131.800 7.400 ;
        RECT 129.400 6.800 130.700 7.200 ;
        RECT 131.400 6.900 132.200 7.200 ;
        RECT 131.800 6.800 132.200 6.900 ;
        RECT 126.900 5.400 129.000 5.700 ;
        RECT 125.400 4.900 126.600 5.200 ;
        RECT 125.100 4.500 125.500 4.600 ;
        RECT 124.400 4.200 125.500 4.500 ;
        RECT 126.300 4.400 126.600 4.900 ;
        RECT 126.300 4.000 127.000 4.400 ;
        RECT 123.100 3.700 123.500 3.800 ;
        RECT 124.500 3.700 124.900 3.800 ;
        RECT 121.400 3.100 121.800 3.500 ;
        RECT 123.100 3.400 124.900 3.700 ;
        RECT 124.200 3.100 124.500 3.400 ;
        RECT 126.200 3.100 126.600 3.500 ;
        RECT 121.400 2.800 122.400 3.100 ;
        RECT 122.000 1.100 122.400 2.800 ;
        RECT 124.200 1.100 124.600 3.100 ;
        RECT 126.300 1.100 126.900 3.100 ;
        RECT 128.600 1.100 129.000 5.400 ;
        RECT 129.400 5.100 129.800 5.200 ;
        RECT 130.400 5.100 130.700 6.800 ;
        RECT 131.000 5.800 131.400 6.600 ;
        RECT 132.600 5.700 133.000 7.400 ;
        RECT 136.100 7.100 136.500 7.200 ;
        RECT 137.400 7.100 137.800 7.200 ;
        RECT 139.000 7.100 139.300 8.200 ;
        RECT 141.400 7.500 141.800 9.900 ;
        RECT 143.800 7.700 144.200 9.900 ;
        RECT 145.900 9.200 146.500 9.900 ;
        RECT 145.900 8.900 146.600 9.200 ;
        RECT 148.200 8.900 148.600 9.900 ;
        RECT 150.400 9.200 150.800 9.900 ;
        RECT 150.400 8.900 151.400 9.200 ;
        RECT 146.200 8.500 146.600 8.900 ;
        RECT 148.300 8.600 148.600 8.900 ;
        RECT 148.300 8.300 149.700 8.600 ;
        RECT 149.300 8.200 149.700 8.300 ;
        RECT 150.200 8.200 150.600 8.600 ;
        RECT 151.000 8.500 151.400 8.900 ;
        RECT 145.300 7.700 145.700 7.800 ;
        RECT 143.800 7.400 145.700 7.700 ;
        RECT 140.600 7.100 141.400 7.200 ;
        RECT 135.900 6.800 141.400 7.100 ;
        RECT 135.000 6.400 135.400 6.500 ;
        RECT 133.500 6.100 135.400 6.400 ;
        RECT 133.500 6.000 133.900 6.100 ;
        RECT 134.300 5.700 134.700 5.800 ;
        RECT 132.600 5.400 134.700 5.700 ;
        RECT 129.400 4.800 130.100 5.100 ;
        RECT 130.400 4.800 130.900 5.100 ;
        RECT 129.800 4.200 130.100 4.800 ;
        RECT 129.800 3.800 130.200 4.200 ;
        RECT 130.500 1.100 130.900 4.800 ;
        RECT 132.600 1.100 133.000 5.400 ;
        RECT 135.900 5.200 136.200 6.800 ;
        RECT 139.500 6.700 139.900 6.800 ;
        RECT 139.000 6.200 139.400 6.300 ;
        RECT 140.300 6.200 140.700 6.300 ;
        RECT 138.200 5.900 140.700 6.200 ;
        RECT 138.200 5.800 138.600 5.900 ;
        RECT 143.800 5.700 144.200 7.400 ;
        RECT 147.300 7.100 147.700 7.200 ;
        RECT 149.400 7.100 149.800 7.200 ;
        RECT 150.200 7.100 150.500 8.200 ;
        RECT 152.600 7.500 153.000 9.900 ;
        RECT 154.700 8.200 155.100 9.900 ;
        RECT 154.200 7.900 155.100 8.200 ;
        RECT 155.800 7.900 156.200 9.900 ;
        RECT 156.600 8.000 157.000 9.900 ;
        RECT 158.200 8.000 158.600 9.900 ;
        RECT 156.600 7.900 158.600 8.000 ;
        RECT 159.000 8.000 159.400 9.900 ;
        RECT 160.600 8.000 161.000 9.900 ;
        RECT 159.000 7.900 161.000 8.000 ;
        RECT 161.400 7.900 161.800 9.900 ;
        RECT 162.500 8.200 162.900 9.900 ;
        RECT 162.500 7.900 163.400 8.200 ;
        RECT 151.800 7.100 152.600 7.200 ;
        RECT 147.100 6.800 152.600 7.100 ;
        RECT 153.400 6.800 153.800 7.600 ;
        RECT 146.200 6.400 146.600 6.500 ;
        RECT 144.700 6.100 146.600 6.400 ;
        RECT 144.700 6.000 145.100 6.100 ;
        RECT 145.500 5.700 145.900 5.800 ;
        RECT 139.000 5.500 141.800 5.600 ;
        RECT 138.900 5.400 141.800 5.500 ;
        RECT 135.000 4.900 136.200 5.200 ;
        RECT 136.900 5.300 141.800 5.400 ;
        RECT 136.900 5.100 139.300 5.300 ;
        RECT 135.000 4.400 135.300 4.900 ;
        RECT 134.600 4.000 135.300 4.400 ;
        RECT 136.100 4.500 136.500 4.600 ;
        RECT 136.900 4.500 137.200 5.100 ;
        RECT 136.100 4.200 137.200 4.500 ;
        RECT 137.500 4.500 140.200 4.800 ;
        RECT 137.500 4.400 137.900 4.500 ;
        RECT 139.800 4.400 140.200 4.500 ;
        RECT 136.700 3.700 137.100 3.800 ;
        RECT 138.100 3.700 138.500 3.800 ;
        RECT 135.000 3.100 135.400 3.500 ;
        RECT 136.700 3.400 138.500 3.700 ;
        RECT 137.100 3.100 137.400 3.400 ;
        RECT 139.800 3.100 140.200 3.500 ;
        RECT 134.700 1.100 135.300 3.100 ;
        RECT 137.000 1.100 137.400 3.100 ;
        RECT 139.200 2.800 140.200 3.100 ;
        RECT 139.200 1.100 139.600 2.800 ;
        RECT 141.400 1.100 141.800 5.300 ;
        RECT 143.800 5.400 145.900 5.700 ;
        RECT 143.800 1.100 144.200 5.400 ;
        RECT 147.100 5.200 147.400 6.800 ;
        RECT 150.700 6.700 151.100 6.800 ;
        RECT 150.200 6.200 150.600 6.300 ;
        RECT 151.500 6.200 151.900 6.300 ;
        RECT 149.400 5.900 151.900 6.200 ;
        RECT 154.200 6.100 154.600 7.900 ;
        RECT 155.900 7.200 156.200 7.900 ;
        RECT 156.700 7.700 158.500 7.900 ;
        RECT 159.100 7.700 160.900 7.900 ;
        RECT 157.800 7.200 158.200 7.400 ;
        RECT 159.400 7.200 159.800 7.400 ;
        RECT 161.400 7.200 161.700 7.900 ;
        RECT 155.800 6.800 157.100 7.200 ;
        RECT 157.800 7.100 158.600 7.200 ;
        RECT 159.000 7.100 159.800 7.200 ;
        RECT 157.800 6.900 159.800 7.100 ;
        RECT 158.200 6.800 159.400 6.900 ;
        RECT 160.500 6.800 161.800 7.200 ;
        RECT 149.400 5.800 149.800 5.900 ;
        RECT 154.200 5.800 156.100 6.100 ;
        RECT 150.200 5.500 153.000 5.600 ;
        RECT 150.100 5.400 153.000 5.500 ;
        RECT 146.200 4.900 147.400 5.200 ;
        RECT 148.100 5.300 153.000 5.400 ;
        RECT 148.100 5.100 150.500 5.300 ;
        RECT 146.200 4.400 146.500 4.900 ;
        RECT 145.800 4.000 146.500 4.400 ;
        RECT 147.300 4.500 147.700 4.600 ;
        RECT 148.100 4.500 148.400 5.100 ;
        RECT 147.300 4.200 148.400 4.500 ;
        RECT 148.700 4.500 151.400 4.800 ;
        RECT 148.700 4.400 149.100 4.500 ;
        RECT 151.000 4.400 151.400 4.500 ;
        RECT 147.900 3.700 148.300 3.800 ;
        RECT 149.300 3.700 149.700 3.800 ;
        RECT 146.200 3.100 146.600 3.500 ;
        RECT 147.900 3.400 149.700 3.700 ;
        RECT 148.300 3.100 148.600 3.400 ;
        RECT 151.000 3.100 151.400 3.500 ;
        RECT 145.900 1.100 146.500 3.100 ;
        RECT 148.200 1.100 148.600 3.100 ;
        RECT 150.400 2.800 151.400 3.100 ;
        RECT 150.400 1.100 150.800 2.800 ;
        RECT 152.600 1.100 153.000 5.300 ;
        RECT 154.200 1.100 154.600 5.800 ;
        RECT 155.800 5.200 156.100 5.800 ;
        RECT 155.000 4.400 155.400 5.200 ;
        RECT 155.800 5.100 156.200 5.200 ;
        RECT 156.800 5.100 157.100 6.800 ;
        RECT 157.400 5.800 157.800 6.600 ;
        RECT 158.200 6.100 158.600 6.200 ;
        RECT 159.800 6.100 160.200 6.600 ;
        RECT 158.200 5.800 160.200 6.100 ;
        RECT 160.500 5.100 160.800 6.800 ;
        RECT 163.000 6.100 163.400 7.900 ;
        RECT 164.600 7.700 165.000 9.900 ;
        RECT 166.700 9.200 167.300 9.900 ;
        RECT 166.700 8.900 167.400 9.200 ;
        RECT 169.000 8.900 169.400 9.900 ;
        RECT 171.200 9.200 171.600 9.900 ;
        RECT 171.200 8.900 172.200 9.200 ;
        RECT 167.000 8.500 167.400 8.900 ;
        RECT 169.100 8.600 169.400 8.900 ;
        RECT 169.100 8.300 170.500 8.600 ;
        RECT 170.100 8.200 170.500 8.300 ;
        RECT 171.000 7.800 171.400 8.600 ;
        RECT 171.800 8.500 172.200 8.900 ;
        RECT 166.100 7.700 166.500 7.800 ;
        RECT 163.800 7.100 164.200 7.600 ;
        RECT 164.600 7.400 166.500 7.700 ;
        RECT 164.600 7.100 165.000 7.400 ;
        RECT 168.100 7.100 168.500 7.200 ;
        RECT 171.000 7.100 171.300 7.800 ;
        RECT 173.400 7.500 173.800 9.900 ;
        RECT 175.500 8.200 175.900 9.900 ;
        RECT 177.400 8.800 177.800 9.900 ;
        RECT 175.000 8.100 175.900 8.200 ;
        RECT 176.600 8.100 177.000 8.600 ;
        RECT 175.000 7.800 177.000 8.100 ;
        RECT 172.600 7.100 173.400 7.200 ;
        RECT 163.800 6.800 165.000 7.100 ;
        RECT 161.400 5.800 163.400 6.100 ;
        RECT 161.400 5.200 161.700 5.800 ;
        RECT 161.400 5.100 161.800 5.200 ;
        RECT 155.800 4.800 156.500 5.100 ;
        RECT 156.800 4.800 157.300 5.100 ;
        RECT 156.200 4.200 156.500 4.800 ;
        RECT 156.200 3.800 156.600 4.200 ;
        RECT 156.900 1.100 157.300 4.800 ;
        RECT 160.300 4.800 160.800 5.100 ;
        RECT 161.100 4.800 161.800 5.100 ;
        RECT 160.300 1.100 160.700 4.800 ;
        RECT 161.100 4.200 161.400 4.800 ;
        RECT 162.200 4.400 162.600 5.200 ;
        RECT 161.000 3.800 161.400 4.200 ;
        RECT 163.000 1.100 163.400 5.800 ;
        RECT 164.600 5.700 165.000 6.800 ;
        RECT 167.900 6.800 173.400 7.100 ;
        RECT 167.000 6.400 167.400 6.500 ;
        RECT 165.500 6.100 167.400 6.400 ;
        RECT 165.500 6.000 165.900 6.100 ;
        RECT 166.300 5.700 166.700 5.800 ;
        RECT 164.600 5.400 166.700 5.700 ;
        RECT 164.600 1.100 165.000 5.400 ;
        RECT 167.900 5.200 168.200 6.800 ;
        RECT 171.500 6.700 171.900 6.800 ;
        RECT 172.300 6.200 172.700 6.300 ;
        RECT 170.200 5.900 172.700 6.200 ;
        RECT 170.200 5.800 170.600 5.900 ;
        RECT 171.000 5.500 173.800 5.600 ;
        RECT 170.900 5.400 173.800 5.500 ;
        RECT 167.000 4.900 168.200 5.200 ;
        RECT 168.900 5.300 173.800 5.400 ;
        RECT 168.900 5.100 171.300 5.300 ;
        RECT 167.000 4.400 167.300 4.900 ;
        RECT 166.600 4.000 167.300 4.400 ;
        RECT 168.100 4.500 168.500 4.600 ;
        RECT 168.900 4.500 169.200 5.100 ;
        RECT 168.100 4.200 169.200 4.500 ;
        RECT 169.500 4.500 172.200 4.800 ;
        RECT 169.500 4.400 169.900 4.500 ;
        RECT 171.800 4.400 172.200 4.500 ;
        RECT 168.700 3.700 169.100 3.800 ;
        RECT 170.100 3.700 170.500 3.800 ;
        RECT 167.000 3.100 167.400 3.500 ;
        RECT 168.700 3.400 170.500 3.700 ;
        RECT 169.100 3.100 169.400 3.400 ;
        RECT 171.800 3.100 172.200 3.500 ;
        RECT 166.700 1.100 167.300 3.100 ;
        RECT 169.000 1.100 169.400 3.100 ;
        RECT 171.200 2.800 172.200 3.100 ;
        RECT 171.200 1.100 171.600 2.800 ;
        RECT 173.400 1.100 173.800 5.300 ;
        RECT 175.000 1.100 175.400 7.800 ;
        RECT 177.500 7.200 177.800 8.800 ;
        RECT 179.300 8.200 179.700 9.900 ;
        RECT 179.300 7.900 180.200 8.200 ;
        RECT 177.400 6.800 177.800 7.200 ;
        RECT 177.500 5.100 177.800 6.800 ;
        RECT 178.200 6.100 178.600 6.200 ;
        RECT 179.800 6.100 180.200 7.900 ;
        RECT 183.000 7.900 183.400 9.900 ;
        RECT 185.400 8.800 185.800 9.900 ;
        RECT 183.700 8.200 184.100 8.600 ;
        RECT 182.200 6.400 182.600 7.200 ;
        RECT 178.200 5.800 180.200 6.100 ;
        RECT 183.000 6.100 183.300 7.900 ;
        RECT 183.800 7.800 184.200 8.200 ;
        RECT 185.500 7.200 185.800 8.800 ;
        RECT 188.600 7.900 189.000 9.900 ;
        RECT 191.000 8.900 191.400 9.900 ;
        RECT 189.300 8.200 189.700 8.600 ;
        RECT 185.400 6.800 185.800 7.200 ;
        RECT 183.800 6.100 184.200 6.200 ;
        RECT 183.000 5.800 184.200 6.100 ;
        RECT 178.200 5.400 178.600 5.800 ;
        RECT 177.400 4.700 178.300 5.100 ;
        RECT 177.900 1.100 178.300 4.700 ;
        RECT 179.800 1.100 180.200 5.800 ;
        RECT 183.800 5.100 184.100 5.800 ;
        RECT 185.500 5.100 185.800 6.800 ;
        RECT 187.800 6.400 188.200 7.200 ;
        RECT 188.600 6.100 188.900 7.900 ;
        RECT 189.400 7.800 189.800 8.200 ;
        RECT 189.400 7.100 189.700 7.800 ;
        RECT 191.100 7.200 191.400 8.900 ;
        RECT 195.800 7.900 196.200 9.900 ;
        RECT 198.200 8.900 198.600 9.900 ;
        RECT 196.500 8.200 196.900 8.600 ;
        RECT 191.000 7.100 191.400 7.200 ;
        RECT 189.400 6.800 191.400 7.100 ;
        RECT 193.400 7.100 193.800 7.200 ;
        RECT 195.000 7.100 195.400 7.200 ;
        RECT 193.400 6.800 195.400 7.100 ;
        RECT 189.400 6.100 189.800 6.200 ;
        RECT 188.600 5.800 189.800 6.100 ;
        RECT 189.400 5.200 189.700 5.800 ;
        RECT 181.400 4.800 183.400 5.100 ;
        RECT 181.400 1.100 181.800 4.800 ;
        RECT 183.000 1.100 183.400 4.800 ;
        RECT 183.800 1.100 184.200 5.100 ;
        RECT 185.400 4.700 186.300 5.100 ;
        RECT 185.900 1.100 186.300 4.700 ;
        RECT 187.000 4.800 189.000 5.100 ;
        RECT 187.000 1.100 187.400 4.800 ;
        RECT 188.600 1.100 189.000 4.800 ;
        RECT 189.400 1.100 189.800 5.200 ;
        RECT 191.100 5.100 191.400 6.800 ;
        RECT 195.000 6.400 195.400 6.800 ;
        RECT 195.800 6.100 196.100 7.900 ;
        RECT 196.600 7.800 197.000 8.200 ;
        RECT 196.600 7.100 196.900 7.800 ;
        RECT 198.300 7.200 198.600 8.900 ;
        RECT 199.800 7.500 200.200 9.900 ;
        RECT 202.000 9.200 202.400 9.900 ;
        RECT 201.400 8.900 202.400 9.200 ;
        RECT 204.200 8.900 204.600 9.900 ;
        RECT 206.300 9.200 206.900 9.900 ;
        RECT 206.200 8.900 206.900 9.200 ;
        RECT 201.400 8.500 201.800 8.900 ;
        RECT 204.200 8.600 204.500 8.900 ;
        RECT 202.200 8.200 202.600 8.600 ;
        RECT 203.100 8.300 204.500 8.600 ;
        RECT 206.200 8.500 206.600 8.900 ;
        RECT 203.100 8.200 203.500 8.300 ;
        RECT 198.200 7.100 198.600 7.200 ;
        RECT 196.600 6.800 198.600 7.100 ;
        RECT 200.200 7.100 201.000 7.200 ;
        RECT 202.300 7.100 202.600 8.200 ;
        RECT 207.100 7.700 207.500 7.800 ;
        RECT 208.600 7.700 209.000 9.900 ;
        RECT 207.100 7.400 209.000 7.700 ;
        RECT 205.100 7.100 205.500 7.200 ;
        RECT 200.200 6.800 205.700 7.100 ;
        RECT 196.600 6.100 197.000 6.200 ;
        RECT 195.800 5.800 197.000 6.100 ;
        RECT 196.600 5.100 196.900 5.800 ;
        RECT 198.300 5.100 198.600 6.800 ;
        RECT 201.700 6.700 202.100 6.800 ;
        RECT 200.900 6.200 201.300 6.300 ;
        RECT 202.200 6.200 202.600 6.300 ;
        RECT 205.400 6.200 205.700 6.800 ;
        RECT 206.200 6.400 206.600 6.500 ;
        RECT 200.900 5.900 203.400 6.200 ;
        RECT 203.000 5.800 203.400 5.900 ;
        RECT 205.400 5.800 205.800 6.200 ;
        RECT 206.200 6.100 208.100 6.400 ;
        RECT 207.700 6.000 208.100 6.100 ;
        RECT 199.800 5.500 202.600 5.600 ;
        RECT 199.800 5.400 202.700 5.500 ;
        RECT 199.800 5.300 204.700 5.400 ;
        RECT 191.000 4.700 191.900 5.100 ;
        RECT 191.500 1.100 191.900 4.700 ;
        RECT 194.200 4.800 196.200 5.100 ;
        RECT 194.200 1.100 194.600 4.800 ;
        RECT 195.800 1.100 196.200 4.800 ;
        RECT 196.600 1.100 197.000 5.100 ;
        RECT 198.200 4.700 199.100 5.100 ;
        RECT 198.700 1.100 199.100 4.700 ;
        RECT 199.800 1.100 200.200 5.300 ;
        RECT 202.300 5.100 204.700 5.300 ;
        RECT 201.400 4.500 204.100 4.800 ;
        RECT 201.400 4.400 201.800 4.500 ;
        RECT 203.700 4.400 204.100 4.500 ;
        RECT 204.400 4.500 204.700 5.100 ;
        RECT 205.400 5.200 205.700 5.800 ;
        RECT 206.900 5.700 207.300 5.800 ;
        RECT 208.600 5.700 209.000 7.400 ;
        RECT 206.900 5.400 209.000 5.700 ;
        RECT 205.400 4.900 206.600 5.200 ;
        RECT 205.100 4.500 205.500 4.600 ;
        RECT 204.400 4.200 205.500 4.500 ;
        RECT 206.300 4.400 206.600 4.900 ;
        RECT 206.300 4.000 207.000 4.400 ;
        RECT 203.100 3.700 203.500 3.800 ;
        RECT 204.500 3.700 204.900 3.800 ;
        RECT 201.400 3.100 201.800 3.500 ;
        RECT 203.100 3.400 204.900 3.700 ;
        RECT 204.200 3.100 204.500 3.400 ;
        RECT 206.200 3.100 206.600 3.500 ;
        RECT 201.400 2.800 202.400 3.100 ;
        RECT 202.000 1.100 202.400 2.800 ;
        RECT 204.200 1.100 204.600 3.100 ;
        RECT 206.300 1.100 206.900 3.100 ;
        RECT 208.600 1.100 209.000 5.400 ;
        RECT 209.400 7.700 209.800 9.900 ;
        RECT 211.500 9.200 212.100 9.900 ;
        RECT 211.500 8.900 212.200 9.200 ;
        RECT 213.800 8.900 214.200 9.900 ;
        RECT 216.000 9.200 216.400 9.900 ;
        RECT 216.000 8.900 217.000 9.200 ;
        RECT 211.800 8.500 212.200 8.900 ;
        RECT 213.900 8.600 214.200 8.900 ;
        RECT 213.900 8.300 215.300 8.600 ;
        RECT 214.900 8.200 215.300 8.300 ;
        RECT 215.800 7.800 216.200 8.600 ;
        RECT 216.600 8.500 217.000 8.900 ;
        RECT 210.900 7.700 211.300 7.800 ;
        RECT 209.400 7.400 211.300 7.700 ;
        RECT 209.400 5.700 209.800 7.400 ;
        RECT 212.900 7.100 213.300 7.200 ;
        RECT 215.800 7.100 216.100 7.800 ;
        RECT 218.200 7.500 218.600 9.900 ;
        RECT 219.300 9.200 219.700 9.900 ;
        RECT 219.300 8.800 220.200 9.200 ;
        RECT 219.300 8.200 219.700 8.800 ;
        RECT 219.300 7.900 220.200 8.200 ;
        RECT 217.400 7.100 218.200 7.200 ;
        RECT 212.700 6.800 218.200 7.100 ;
        RECT 211.800 6.400 212.200 6.500 ;
        RECT 210.300 6.100 212.200 6.400 ;
        RECT 210.300 6.000 210.700 6.100 ;
        RECT 211.100 5.700 211.500 5.800 ;
        RECT 209.400 5.400 211.500 5.700 ;
        RECT 209.400 1.100 209.800 5.400 ;
        RECT 212.700 5.200 213.000 6.800 ;
        RECT 216.300 6.700 216.700 6.800 ;
        RECT 217.100 6.200 217.500 6.300 ;
        RECT 213.400 6.100 213.800 6.200 ;
        RECT 215.000 6.100 217.500 6.200 ;
        RECT 213.400 5.900 217.500 6.100 ;
        RECT 213.400 5.800 215.400 5.900 ;
        RECT 215.800 5.500 218.600 5.600 ;
        RECT 215.700 5.400 218.600 5.500 ;
        RECT 211.800 4.900 213.000 5.200 ;
        RECT 213.700 5.300 218.600 5.400 ;
        RECT 213.700 5.100 216.100 5.300 ;
        RECT 211.800 4.400 212.100 4.900 ;
        RECT 211.400 4.000 212.100 4.400 ;
        RECT 212.900 4.500 213.300 4.600 ;
        RECT 213.700 4.500 214.000 5.100 ;
        RECT 212.900 4.200 214.000 4.500 ;
        RECT 214.300 4.500 217.000 4.800 ;
        RECT 214.300 4.400 214.700 4.500 ;
        RECT 216.600 4.400 217.000 4.500 ;
        RECT 213.500 3.700 213.900 3.800 ;
        RECT 214.900 3.700 215.300 3.800 ;
        RECT 211.800 3.100 212.200 3.500 ;
        RECT 213.500 3.400 215.300 3.700 ;
        RECT 213.900 3.100 214.200 3.400 ;
        RECT 216.600 3.100 217.000 3.500 ;
        RECT 211.500 1.100 212.100 3.100 ;
        RECT 213.800 1.100 214.200 3.100 ;
        RECT 216.000 2.800 217.000 3.100 ;
        RECT 216.000 1.100 216.400 2.800 ;
        RECT 218.200 1.100 218.600 5.300 ;
        RECT 219.000 4.400 219.400 5.200 ;
        RECT 219.800 1.100 220.200 7.900 ;
        RECT 221.400 7.700 221.800 9.900 ;
        RECT 223.500 9.200 224.100 9.900 ;
        RECT 223.500 8.900 224.200 9.200 ;
        RECT 225.800 8.900 226.200 9.900 ;
        RECT 228.000 9.200 228.400 9.900 ;
        RECT 228.000 8.900 229.000 9.200 ;
        RECT 223.800 8.500 224.200 8.900 ;
        RECT 225.900 8.600 226.200 8.900 ;
        RECT 225.900 8.300 227.300 8.600 ;
        RECT 226.900 8.200 227.300 8.300 ;
        RECT 227.800 8.200 228.200 8.600 ;
        RECT 228.600 8.500 229.000 8.900 ;
        RECT 222.900 7.700 223.300 7.800 ;
        RECT 220.600 6.800 221.000 7.600 ;
        RECT 221.400 7.400 223.300 7.700 ;
        RECT 221.400 5.700 221.800 7.400 ;
        RECT 224.900 7.100 225.300 7.200 ;
        RECT 227.800 7.100 228.100 8.200 ;
        RECT 230.200 7.500 230.600 9.900 ;
        RECT 229.400 7.100 230.200 7.200 ;
        RECT 224.700 6.800 230.200 7.100 ;
        RECT 223.800 6.400 224.200 6.500 ;
        RECT 222.300 6.100 224.200 6.400 ;
        RECT 224.700 6.200 225.000 6.800 ;
        RECT 228.300 6.700 228.700 6.800 ;
        RECT 229.100 6.200 229.500 6.300 ;
        RECT 222.300 6.000 222.700 6.100 ;
        RECT 224.600 5.800 225.000 6.200 ;
        RECT 227.000 5.900 229.500 6.200 ;
        RECT 227.000 5.800 227.400 5.900 ;
        RECT 223.100 5.700 223.500 5.800 ;
        RECT 221.400 5.400 223.500 5.700 ;
        RECT 221.400 1.100 221.800 5.400 ;
        RECT 224.700 5.200 225.000 5.800 ;
        RECT 227.800 5.500 230.600 5.600 ;
        RECT 227.700 5.400 230.600 5.500 ;
        RECT 223.800 4.900 225.000 5.200 ;
        RECT 225.700 5.300 230.600 5.400 ;
        RECT 225.700 5.100 228.100 5.300 ;
        RECT 223.800 4.400 224.100 4.900 ;
        RECT 223.400 4.000 224.100 4.400 ;
        RECT 224.900 4.500 225.300 4.600 ;
        RECT 225.700 4.500 226.000 5.100 ;
        RECT 224.900 4.200 226.000 4.500 ;
        RECT 226.300 4.500 229.000 4.800 ;
        RECT 226.300 4.400 226.700 4.500 ;
        RECT 228.600 4.400 229.000 4.500 ;
        RECT 225.500 3.700 225.900 3.800 ;
        RECT 226.900 3.700 227.300 3.800 ;
        RECT 223.800 3.100 224.200 3.500 ;
        RECT 225.500 3.400 227.300 3.700 ;
        RECT 225.900 3.100 226.200 3.400 ;
        RECT 228.600 3.100 229.000 3.500 ;
        RECT 223.500 1.100 224.100 3.100 ;
        RECT 225.800 1.100 226.200 3.100 ;
        RECT 228.000 2.800 229.000 3.100 ;
        RECT 228.000 1.100 228.400 2.800 ;
        RECT 230.200 1.100 230.600 5.300 ;
      LAYER via1 ;
        RECT 14.200 206.800 14.600 207.200 ;
        RECT 15.800 206.800 16.200 207.200 ;
        RECT 6.200 201.800 6.600 202.200 ;
        RECT 15.000 205.100 15.400 205.500 ;
        RECT 31.800 206.800 32.200 207.200 ;
        RECT 35.000 206.800 35.400 207.200 ;
        RECT 33.400 205.900 33.800 206.300 ;
        RECT 23.800 201.800 24.200 202.200 ;
        RECT 31.000 205.100 31.400 205.500 ;
        RECT 27.000 203.800 27.400 204.200 ;
        RECT 46.200 206.800 46.600 207.200 ;
        RECT 44.600 205.800 45.000 206.200 ;
        RECT 45.400 205.100 45.800 205.500 ;
        RECT 39.800 202.800 40.200 203.200 ;
        RECT 43.000 203.800 43.400 204.200 ;
        RECT 56.600 206.800 57.000 207.200 ;
        RECT 54.200 203.800 54.600 204.200 ;
        RECT 67.000 206.800 67.400 207.200 ;
        RECT 63.800 205.800 64.200 206.200 ;
        RECT 64.600 205.100 65.000 205.500 ;
        RECT 62.200 201.800 62.600 202.200 ;
        RECT 73.400 201.800 73.800 202.200 ;
        RECT 82.200 206.800 82.600 207.200 ;
        RECT 92.600 206.800 93.000 207.200 ;
        RECT 76.600 206.100 77.000 206.500 ;
        RECT 80.600 205.900 81.000 206.300 ;
        RECT 90.200 205.800 90.600 206.200 ;
        RECT 94.200 205.900 94.600 206.300 ;
        RECT 83.000 205.100 83.400 205.500 ;
        RECT 74.200 201.800 74.600 202.200 ;
        RECT 91.800 205.100 92.200 205.500 ;
        RECT 86.200 203.800 86.600 204.200 ;
        RECT 102.200 206.800 102.600 207.200 ;
        RECT 100.600 202.800 101.000 203.200 ;
        RECT 101.400 205.100 101.800 205.500 ;
        RECT 124.600 206.800 125.000 207.200 ;
        RECT 112.600 205.800 113.000 206.200 ;
        RECT 119.800 205.800 120.200 206.200 ;
        RECT 108.600 203.800 109.000 204.200 ;
        RECT 110.200 203.800 110.600 204.200 ;
        RECT 119.800 204.800 120.200 205.200 ;
        RECT 126.200 205.900 126.600 206.300 ;
        RECT 123.800 205.100 124.200 205.500 ;
        RECT 123.000 203.800 123.400 204.200 ;
        RECT 151.000 208.800 151.400 209.200 ;
        RECT 143.000 206.800 143.400 207.200 ;
        RECT 132.600 203.800 133.000 204.200 ;
        RECT 134.200 201.800 134.600 202.200 ;
        RECT 139.000 201.800 139.400 202.200 ;
        RECT 142.200 205.100 142.600 205.500 ;
        RECT 153.400 205.800 153.800 206.200 ;
        RECT 149.400 203.800 149.800 204.200 ;
        RECT 155.000 204.800 155.400 205.200 ;
        RECT 168.600 206.800 169.000 207.200 ;
        RECT 173.400 206.800 173.800 207.200 ;
        RECT 163.000 206.100 163.400 206.500 ;
        RECT 159.000 201.800 159.400 202.200 ;
        RECT 167.000 205.900 167.400 206.300 ;
        RECT 169.400 205.100 169.800 205.500 ;
        RECT 184.600 208.800 185.000 209.200 ;
        RECT 178.200 205.900 178.600 206.300 ;
        RECT 160.600 201.800 161.000 202.200 ;
        RECT 173.400 204.800 173.800 205.200 ;
        RECT 175.800 205.100 176.200 205.500 ;
        RECT 186.200 201.800 186.600 202.200 ;
        RECT 205.400 206.800 205.800 207.200 ;
        RECT 211.000 208.800 211.400 209.200 ;
        RECT 206.200 204.800 206.600 205.200 ;
        RECT 216.600 206.800 217.000 207.200 ;
        RECT 213.400 206.100 213.800 206.500 ;
        RECT 210.200 204.800 210.600 205.200 ;
        RECT 209.400 201.800 209.800 202.200 ;
        RECT 219.800 205.100 220.200 205.500 ;
        RECT 220.600 204.800 221.000 205.200 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 221.400 201.800 221.800 202.200 ;
        RECT 225.400 204.800 225.800 205.200 ;
        RECT 227.000 201.800 227.400 202.200 ;
        RECT 0.600 197.800 1.000 198.200 ;
        RECT 7.800 196.200 8.200 196.600 ;
        RECT 9.400 195.500 9.800 195.900 ;
        RECT 18.200 198.800 18.600 199.200 ;
        RECT 15.000 196.800 15.400 197.200 ;
        RECT 11.800 194.800 12.200 195.200 ;
        RECT 21.400 196.800 21.800 197.200 ;
        RECT 25.400 196.800 25.800 197.200 ;
        RECT 15.000 194.800 15.400 195.200 ;
        RECT 18.200 194.800 18.600 195.200 ;
        RECT 23.000 194.800 23.400 195.200 ;
        RECT 38.200 196.800 38.600 197.200 ;
        RECT 47.800 196.800 48.200 197.200 ;
        RECT 27.800 194.800 28.200 195.200 ;
        RECT 9.400 193.100 9.800 193.500 ;
        RECT 12.600 193.800 13.000 194.200 ;
        RECT 15.800 193.800 16.200 194.200 ;
        RECT 19.000 193.800 19.400 194.200 ;
        RECT 23.000 193.800 23.400 194.200 ;
        RECT 27.000 193.800 27.400 194.200 ;
        RECT 28.600 193.800 29.000 194.200 ;
        RECT 29.400 193.100 29.800 193.500 ;
        RECT 45.400 194.800 45.800 195.200 ;
        RECT 41.400 193.800 41.800 194.200 ;
        RECT 40.600 193.100 41.000 193.500 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 52.600 193.800 53.000 194.200 ;
        RECT 56.600 194.800 57.000 195.200 ;
        RECT 57.400 194.800 57.800 195.200 ;
        RECT 59.000 194.800 59.400 195.200 ;
        RECT 60.600 193.800 61.000 194.200 ;
        RECT 62.200 193.800 62.600 194.200 ;
        RECT 49.400 191.800 49.800 192.200 ;
        RECT 61.400 193.100 61.800 193.500 ;
        RECT 55.800 191.800 56.200 192.200 ;
        RECT 71.800 194.800 72.200 195.200 ;
        RECT 75.000 194.800 75.400 195.200 ;
        RECT 79.000 194.800 79.400 195.200 ;
        RECT 82.200 194.800 82.600 195.200 ;
        RECT 84.600 194.800 85.000 195.200 ;
        RECT 87.800 194.800 88.200 195.200 ;
        RECT 91.000 195.800 91.400 196.200 ;
        RECT 72.600 193.800 73.000 194.200 ;
        RECT 79.800 193.800 80.200 194.200 ;
        RECT 83.000 193.800 83.400 194.200 ;
        RECT 86.200 193.800 86.600 194.200 ;
        RECT 91.800 193.100 92.200 193.500 ;
        RECT 70.200 191.800 70.600 192.200 ;
        RECT 102.200 194.800 102.600 195.200 ;
        RECT 105.400 194.800 105.800 195.200 ;
        RECT 126.200 196.800 126.600 197.200 ;
        RECT 103.800 193.800 104.200 194.200 ;
        RECT 108.600 193.800 109.000 194.200 ;
        RECT 107.800 193.100 108.200 193.500 ;
        RECT 100.600 191.800 101.000 192.200 ;
        RECT 121.400 194.800 121.800 195.200 ;
        RECT 116.600 191.800 117.000 192.200 ;
        RECT 117.400 193.100 117.800 193.500 ;
        RECT 127.800 194.800 128.200 195.200 ;
        RECT 135.800 196.800 136.200 197.200 ;
        RECT 141.400 196.800 141.800 197.200 ;
        RECT 138.200 195.800 138.600 196.200 ;
        RECT 138.200 194.800 138.600 195.200 ;
        RECT 119.800 192.800 120.200 193.200 ;
        RECT 132.600 193.800 133.000 194.200 ;
        RECT 139.000 193.800 139.400 194.200 ;
        RECT 148.600 196.200 149.000 196.600 ;
        RECT 150.200 195.500 150.600 195.900 ;
        RECT 158.200 196.200 158.600 196.600 ;
        RECT 159.800 195.500 160.200 195.900 ;
        RECT 161.400 194.800 161.800 195.200 ;
        RECT 150.200 193.100 150.600 193.500 ;
        RECT 163.000 193.800 163.400 194.200 ;
        RECT 159.800 193.100 160.200 193.500 ;
        RECT 173.400 196.200 173.800 196.600 ;
        RECT 175.000 195.500 175.400 195.900 ;
        RECT 176.600 194.800 177.000 195.200 ;
        RECT 151.000 191.800 151.400 192.200 ;
        RECT 175.000 193.100 175.400 193.500 ;
        RECT 180.600 193.800 181.000 194.200 ;
        RECT 184.600 194.800 185.000 195.200 ;
        RECT 185.400 194.800 185.800 195.200 ;
        RECT 187.000 194.800 187.400 195.200 ;
        RECT 189.400 193.800 189.800 194.200 ;
        RECT 166.200 191.800 166.600 192.200 ;
        RECT 192.600 193.800 193.000 194.200 ;
        RECT 200.600 196.200 201.000 196.600 ;
        RECT 202.200 195.500 202.600 195.900 ;
        RECT 203.800 194.800 204.200 195.200 ;
        RECT 183.800 191.800 184.200 192.200 ;
        RECT 205.400 193.800 205.800 194.200 ;
        RECT 202.200 193.100 202.600 193.500 ;
        RECT 207.800 193.800 208.200 194.200 ;
        RECT 215.800 196.200 216.200 196.600 ;
        RECT 217.400 195.500 217.800 195.900 ;
        RECT 219.000 194.800 219.400 195.200 ;
        RECT 217.400 193.100 217.800 193.500 ;
        RECT 228.600 196.200 229.000 196.600 ;
        RECT 230.200 195.500 230.600 195.900 ;
        RECT 220.600 191.800 221.000 192.200 ;
        RECT 230.200 193.100 230.600 193.500 ;
        RECT 221.400 191.800 221.800 192.200 ;
        RECT 4.600 185.800 5.000 186.200 ;
        RECT 0.600 185.100 1.000 185.500 ;
        RECT 16.600 185.100 17.000 185.500 ;
        RECT 9.400 183.800 9.800 184.200 ;
        RECT 27.800 186.800 28.200 187.200 ;
        RECT 32.600 186.800 33.000 187.200 ;
        RECT 58.200 188.800 58.600 189.200 ;
        RECT 33.400 185.800 33.800 186.200 ;
        RECT 25.400 183.800 25.800 184.200 ;
        RECT 38.200 185.800 38.600 186.200 ;
        RECT 46.200 186.800 46.600 187.200 ;
        RECT 47.000 185.800 47.400 186.200 ;
        RECT 35.000 183.800 35.400 184.200 ;
        RECT 39.800 181.800 40.200 182.200 ;
        RECT 42.200 185.100 42.600 185.500 ;
        RECT 66.200 188.800 66.600 189.200 ;
        RECT 53.400 185.800 53.800 186.200 ;
        RECT 51.000 181.800 51.400 182.200 ;
        RECT 64.600 185.800 65.000 186.200 ;
        RECT 71.800 186.800 72.200 187.200 ;
        RECT 73.400 185.800 73.800 186.200 ;
        RECT 63.800 181.800 64.200 182.200 ;
        RECT 90.200 186.800 90.600 187.200 ;
        RECT 79.800 186.100 80.200 186.500 ;
        RECT 71.000 181.800 71.400 182.200 ;
        RECT 83.800 185.900 84.200 186.300 ;
        RECT 86.200 185.100 86.600 185.500 ;
        RECT 77.400 183.800 77.800 184.200 ;
        RECT 89.400 185.800 89.800 186.200 ;
        RECT 99.000 186.800 99.400 187.200 ;
        RECT 88.600 183.800 89.000 184.200 ;
        RECT 98.200 185.800 98.600 186.200 ;
        RECT 110.200 187.800 110.600 188.200 ;
        RECT 114.200 188.800 114.600 189.200 ;
        RECT 102.200 182.800 102.600 183.200 ;
        RECT 111.800 185.800 112.200 186.200 ;
        RECT 118.200 184.800 118.600 185.200 ;
        RECT 132.600 188.800 133.000 189.200 ;
        RECT 124.600 186.100 125.000 186.500 ;
        RECT 131.000 185.100 131.400 185.500 ;
        RECT 122.200 183.800 122.600 184.200 ;
        RECT 135.000 185.800 135.400 186.200 ;
        RECT 149.400 186.800 149.800 187.200 ;
        RECT 162.200 188.800 162.600 189.200 ;
        RECT 139.000 185.800 139.400 186.200 ;
        RECT 147.000 185.800 147.400 186.200 ;
        RECT 143.000 183.800 143.400 184.200 ;
        RECT 146.200 184.800 146.600 185.200 ;
        RECT 152.600 185.900 153.000 186.300 ;
        RECT 149.400 184.800 149.800 185.200 ;
        RECT 150.200 185.100 150.600 185.500 ;
        RECT 159.000 183.800 159.400 184.200 ;
        RECT 161.400 184.800 161.800 185.200 ;
        RECT 165.400 181.800 165.800 182.200 ;
        RECT 169.400 186.100 169.800 186.500 ;
        RECT 171.000 185.800 171.400 186.200 ;
        RECT 173.400 185.900 173.800 186.300 ;
        RECT 175.800 185.100 176.200 185.500 ;
        RECT 167.000 181.800 167.400 182.200 ;
        RECT 178.200 184.800 178.600 185.200 ;
        RECT 185.400 186.800 185.800 187.200 ;
        RECT 186.200 185.800 186.600 186.200 ;
        RECT 190.200 185.800 190.600 186.200 ;
        RECT 207.800 188.800 208.200 189.200 ;
        RECT 196.600 185.800 197.000 186.200 ;
        RECT 189.400 181.800 189.800 182.200 ;
        RECT 201.400 185.800 201.800 186.200 ;
        RECT 207.000 185.800 207.400 186.200 ;
        RECT 225.400 188.800 225.800 189.200 ;
        RECT 210.200 186.100 210.600 186.500 ;
        RECT 214.200 185.900 214.600 186.300 ;
        RECT 216.600 185.100 217.000 185.500 ;
        RECT 219.000 184.800 219.400 185.200 ;
        RECT 224.600 184.800 225.000 185.200 ;
        RECT 6.200 178.800 6.600 179.200 ;
        RECT 15.000 176.200 15.400 176.600 ;
        RECT 16.600 175.500 17.000 175.900 ;
        RECT 33.400 178.800 33.800 179.200 ;
        RECT 6.200 171.800 6.600 172.200 ;
        RECT 28.600 174.800 29.000 175.200 ;
        RECT 25.400 173.800 25.800 174.200 ;
        RECT 16.600 173.100 17.000 173.500 ;
        RECT 7.800 171.800 8.200 172.200 ;
        RECT 23.000 171.800 23.400 172.200 ;
        RECT 24.600 173.100 25.000 173.500 ;
        RECT 35.800 174.800 36.200 175.200 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 42.200 174.800 42.600 175.200 ;
        RECT 43.000 174.800 43.400 175.200 ;
        RECT 47.800 174.800 48.200 175.200 ;
        RECT 41.400 171.800 41.800 172.200 ;
        RECT 43.800 173.100 44.200 173.500 ;
        RECT 62.200 178.800 62.600 179.200 ;
        RECT 54.200 174.800 54.600 175.200 ;
        RECT 55.000 174.800 55.400 175.200 ;
        RECT 58.200 174.800 58.600 175.200 ;
        RECT 59.800 174.800 60.200 175.200 ;
        RECT 60.600 174.800 61.000 175.200 ;
        RECT 59.000 173.800 59.400 174.200 ;
        RECT 66.200 174.800 66.600 175.200 ;
        RECT 67.800 174.800 68.200 175.200 ;
        RECT 68.600 174.800 69.000 175.200 ;
        RECT 69.400 174.800 69.800 175.200 ;
        RECT 70.200 174.800 70.600 175.200 ;
        RECT 75.800 178.800 76.200 179.200 ;
        RECT 86.200 176.800 86.600 177.200 ;
        RECT 82.200 174.800 82.600 175.200 ;
        RECT 78.200 173.800 78.600 174.200 ;
        RECT 71.800 171.800 72.200 172.200 ;
        RECT 77.400 173.100 77.800 173.500 ;
        RECT 87.800 174.800 88.200 175.200 ;
        RECT 88.600 174.800 89.000 175.200 ;
        RECT 97.400 178.800 97.800 179.200 ;
        RECT 93.400 174.800 93.800 175.200 ;
        RECT 94.200 173.800 94.600 174.200 ;
        RECT 99.000 173.800 99.400 174.200 ;
        RECT 101.400 173.800 101.800 174.200 ;
        RECT 104.600 174.800 105.000 175.200 ;
        RECT 115.800 176.800 116.200 177.200 ;
        RECT 108.600 174.800 109.000 175.200 ;
        RECT 111.000 174.800 111.400 175.200 ;
        RECT 125.400 176.800 125.800 177.200 ;
        RECT 114.200 174.800 114.600 175.200 ;
        RECT 107.800 173.800 108.200 174.200 ;
        RECT 109.400 173.800 109.800 174.200 ;
        RECT 112.600 173.800 113.000 174.200 ;
        RECT 116.600 173.100 117.000 173.500 ;
        RECT 102.200 171.800 102.600 172.200 ;
        RECT 129.400 174.800 129.800 175.200 ;
        RECT 130.200 174.800 130.600 175.200 ;
        RECT 143.000 178.800 143.400 179.200 ;
        RECT 131.800 173.800 132.200 174.200 ;
        RECT 132.600 173.800 133.000 174.200 ;
        RECT 136.600 174.800 137.000 175.200 ;
        RECT 137.400 174.800 137.800 175.200 ;
        RECT 139.000 174.800 139.400 175.200 ;
        RECT 141.400 175.800 141.800 176.200 ;
        RECT 142.200 174.800 142.600 175.200 ;
        RECT 150.200 176.200 150.600 176.600 ;
        RECT 151.800 175.500 152.200 175.900 ;
        RECT 153.400 174.800 153.800 175.200 ;
        RECT 154.200 173.800 154.600 174.200 ;
        RECT 151.800 173.100 152.200 173.500 ;
        RECT 159.000 174.800 159.400 175.200 ;
        RECT 171.000 176.800 171.400 177.200 ;
        RECT 172.600 176.800 173.000 177.200 ;
        RECT 157.400 173.800 157.800 174.200 ;
        RECT 161.400 173.800 161.800 174.200 ;
        RECT 175.800 178.800 176.200 179.200 ;
        RECT 163.000 173.800 163.400 174.200 ;
        RECT 163.800 173.100 164.200 173.500 ;
        RECT 173.400 174.800 173.800 175.200 ;
        RECT 174.200 174.800 174.600 175.200 ;
        RECT 166.200 172.800 166.600 173.200 ;
        RECT 183.800 173.800 184.200 174.200 ;
        RECT 188.600 174.800 189.000 175.200 ;
        RECT 189.400 174.800 189.800 175.200 ;
        RECT 187.800 173.800 188.200 174.200 ;
        RECT 194.200 174.800 194.600 175.200 ;
        RECT 179.800 171.800 180.200 172.200 ;
        RECT 199.000 174.800 199.400 175.200 ;
        RECT 196.600 173.800 197.000 174.200 ;
        RECT 199.800 173.800 200.200 174.200 ;
        RECT 207.800 176.200 208.200 176.600 ;
        RECT 209.400 175.500 209.800 175.900 ;
        RECT 212.600 173.800 213.000 174.200 ;
        RECT 213.400 173.800 213.800 174.200 ;
        RECT 209.400 173.100 209.800 173.500 ;
        RECT 200.600 171.800 201.000 172.200 ;
        RECT 215.800 177.800 216.200 178.200 ;
        RECT 223.000 176.200 223.400 176.600 ;
        RECT 224.600 175.500 225.000 175.900 ;
        RECT 225.400 173.800 225.800 174.200 ;
        RECT 224.600 173.100 225.000 173.500 ;
        RECT 229.400 174.800 229.800 175.200 ;
        RECT 230.200 173.800 230.600 174.200 ;
        RECT 3.000 165.900 3.400 166.300 ;
        RECT 0.600 165.100 1.000 165.500 ;
        RECT 9.400 161.800 9.800 162.200 ;
        RECT 14.200 168.800 14.600 169.200 ;
        RECT 11.000 161.800 11.400 162.200 ;
        RECT 13.400 164.800 13.800 165.200 ;
        RECT 19.800 166.800 20.200 167.200 ;
        RECT 20.600 165.100 21.000 165.500 ;
        RECT 30.200 163.800 30.600 164.200 ;
        RECT 31.800 164.800 32.200 165.200 ;
        RECT 36.600 165.800 37.000 166.200 ;
        RECT 42.200 165.800 42.600 166.200 ;
        RECT 47.800 165.800 48.200 166.200 ;
        RECT 37.400 165.100 37.800 165.500 ;
        RECT 49.400 161.800 49.800 162.200 ;
        RECT 86.200 168.800 86.600 169.200 ;
        RECT 59.800 164.800 60.200 165.200 ;
        RECT 64.600 165.800 65.000 166.200 ;
        RECT 78.200 166.800 78.600 167.200 ;
        RECT 69.400 165.800 69.800 166.200 ;
        RECT 79.800 165.900 80.200 166.300 ;
        RECT 63.800 161.800 64.200 162.200 ;
        RECT 73.400 164.800 73.800 165.200 ;
        RECT 77.400 165.100 77.800 165.500 ;
        RECT 91.000 166.800 91.400 167.200 ;
        RECT 98.200 165.800 98.600 166.200 ;
        RECT 97.400 164.800 97.800 165.200 ;
        RECT 115.000 168.800 115.400 169.200 ;
        RECT 102.200 164.800 102.600 165.200 ;
        RECT 108.600 165.900 109.000 166.300 ;
        RECT 106.200 165.100 106.600 165.500 ;
        RECT 119.000 165.800 119.400 166.200 ;
        RECT 126.200 165.800 126.600 166.200 ;
        RECT 150.200 168.800 150.600 169.200 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 135.800 165.800 136.200 166.200 ;
        RECT 131.800 164.800 132.200 165.200 ;
        RECT 127.800 161.800 128.200 162.200 ;
        RECT 142.200 166.800 142.600 167.200 ;
        RECT 146.200 166.800 146.600 167.200 ;
        RECT 137.400 161.800 137.800 162.200 ;
        RECT 141.400 165.100 141.800 165.500 ;
        RECT 159.000 166.800 159.400 167.200 ;
        RECT 151.000 161.800 151.400 162.200 ;
        RECT 157.400 164.800 157.800 165.200 ;
        RECT 158.200 165.100 158.600 165.500 ;
        RECT 167.800 163.800 168.200 164.200 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 194.200 168.800 194.600 169.200 ;
        RECT 175.000 165.800 175.400 166.200 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 184.600 166.800 185.000 167.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 175.000 161.800 175.400 162.200 ;
        RECT 178.200 164.800 178.600 165.200 ;
        RECT 187.800 165.900 188.200 166.300 ;
        RECT 180.600 161.800 181.000 162.200 ;
        RECT 184.600 164.800 185.000 165.200 ;
        RECT 185.400 165.100 185.800 165.500 ;
        RECT 199.800 165.800 200.200 166.200 ;
        RECT 199.000 164.800 199.400 165.200 ;
        RECT 211.000 166.800 211.400 167.200 ;
        RECT 208.600 166.100 209.000 166.500 ;
        RECT 212.600 165.900 213.000 166.300 ;
        RECT 215.000 165.100 215.400 165.500 ;
        RECT 217.400 164.800 217.800 165.200 ;
        RECT 223.000 164.800 223.400 165.200 ;
        RECT 222.200 161.800 222.600 162.200 ;
        RECT 229.400 161.800 229.800 162.200 ;
        RECT 2.200 158.800 2.600 159.200 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 3.000 153.800 3.400 154.200 ;
        RECT 5.400 153.800 5.800 154.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 8.600 153.800 9.000 154.200 ;
        RECT 11.800 153.800 12.200 154.200 ;
        RECT 12.600 153.100 13.000 153.500 ;
        RECT 25.400 154.800 25.800 155.200 ;
        RECT 21.400 151.800 21.800 152.200 ;
        RECT 22.200 153.100 22.600 153.500 ;
        RECT 35.800 154.800 36.200 155.200 ;
        RECT 32.600 153.800 33.000 154.200 ;
        RECT 31.000 151.800 31.400 152.200 ;
        RECT 31.800 153.100 32.200 153.500 ;
        RECT 43.800 154.800 44.200 155.200 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 61.400 156.800 61.800 157.200 ;
        RECT 63.000 156.800 63.400 157.200 ;
        RECT 48.600 153.800 49.000 154.200 ;
        RECT 52.600 154.800 53.000 155.200 ;
        RECT 53.400 154.800 53.800 155.200 ;
        RECT 58.200 154.800 58.600 155.200 ;
        RECT 55.000 153.800 55.400 154.200 ;
        RECT 40.600 151.800 41.000 152.200 ;
        RECT 54.200 153.100 54.600 153.500 ;
        RECT 64.600 154.800 65.000 155.200 ;
        RECT 83.000 158.800 83.400 159.200 ;
        RECT 73.400 154.800 73.800 155.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 70.200 151.800 70.600 152.200 ;
        RECT 74.200 153.100 74.600 153.500 ;
        RECT 79.800 153.800 80.200 154.200 ;
        RECT 97.400 158.800 97.800 159.200 ;
        RECT 95.800 156.800 96.200 157.200 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 85.400 154.800 85.800 155.200 ;
        RECT 92.600 154.800 93.000 155.200 ;
        RECT 99.800 156.800 100.200 157.200 ;
        RECT 89.400 153.800 89.800 154.200 ;
        RECT 88.600 153.100 89.000 153.500 ;
        RECT 102.200 154.800 102.600 155.200 ;
        RECT 99.800 153.800 100.200 154.200 ;
        RECT 103.000 153.800 103.400 154.200 ;
        RECT 109.400 154.800 109.800 155.200 ;
        RECT 105.400 153.800 105.800 154.200 ;
        RECT 106.200 153.100 106.600 153.500 ;
        RECT 104.600 151.800 105.000 152.200 ;
        RECT 119.000 154.800 119.400 155.200 ;
        RECT 116.600 153.800 117.000 154.200 ;
        RECT 115.000 151.800 115.400 152.200 ;
        RECT 115.800 153.100 116.200 153.500 ;
        RECT 129.400 158.800 129.800 159.200 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 124.600 151.800 125.000 152.200 ;
        RECT 126.200 151.800 126.600 152.200 ;
        RECT 138.200 156.800 138.600 157.200 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 130.200 153.800 130.600 154.200 ;
        RECT 131.800 153.800 132.200 154.200 ;
        RECT 131.000 153.100 131.400 153.500 ;
        RECT 143.000 152.800 143.400 153.200 ;
        RECT 147.000 154.800 147.400 155.200 ;
        RECT 145.400 153.800 145.800 154.200 ;
        RECT 139.800 151.800 140.200 152.200 ;
        RECT 155.000 154.800 155.400 155.200 ;
        RECT 156.600 154.800 157.000 155.200 ;
        RECT 155.800 153.800 156.200 154.200 ;
        RECT 151.000 151.800 151.400 152.200 ;
        RECT 153.400 151.800 153.800 152.200 ;
        RECT 160.600 156.800 161.000 157.200 ;
        RECT 167.800 156.200 168.200 156.600 ;
        RECT 169.400 155.500 169.800 155.900 ;
        RECT 171.800 155.800 172.200 156.200 ;
        RECT 171.800 154.800 172.200 155.200 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 174.200 154.800 174.600 155.200 ;
        RECT 169.400 153.100 169.800 153.500 ;
        RECT 172.600 153.800 173.000 154.200 ;
        RECT 178.200 154.800 178.600 155.200 ;
        RECT 178.200 153.800 178.600 154.200 ;
        RECT 181.400 154.800 181.800 155.200 ;
        RECT 183.000 153.800 183.400 154.200 ;
        RECT 193.400 156.200 193.800 156.600 ;
        RECT 195.000 155.500 195.400 155.900 ;
        RECT 179.800 151.800 180.200 152.200 ;
        RECT 197.400 153.800 197.800 154.200 ;
        RECT 195.000 153.100 195.400 153.500 ;
        RECT 199.000 156.800 199.400 157.200 ;
        RECT 199.800 154.800 200.200 155.200 ;
        RECT 200.600 154.800 201.000 155.200 ;
        RECT 207.000 154.800 207.400 155.200 ;
        RECT 208.600 154.800 209.000 155.200 ;
        RECT 216.600 158.800 217.000 159.200 ;
        RECT 215.000 154.800 215.400 155.200 ;
        RECT 212.600 153.800 213.000 154.200 ;
        RECT 215.800 153.800 216.200 154.200 ;
        RECT 223.800 156.200 224.200 156.600 ;
        RECT 225.400 155.500 225.800 155.900 ;
        RECT 227.800 154.800 228.200 155.200 ;
        RECT 210.200 151.800 210.600 152.200 ;
        RECT 227.000 153.800 227.400 154.200 ;
        RECT 225.400 153.100 225.800 153.500 ;
        RECT 228.600 153.800 229.000 154.200 ;
        RECT 230.200 153.800 230.600 154.200 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 4.600 146.800 5.000 147.200 ;
        RECT 0.600 145.100 1.000 145.500 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 23.000 148.800 23.400 149.200 ;
        RECT 13.400 144.800 13.800 145.200 ;
        RECT 17.400 145.800 17.800 146.200 ;
        RECT 17.400 144.800 17.800 145.200 ;
        RECT 18.200 144.800 18.600 145.200 ;
        RECT 42.200 148.800 42.600 149.200 ;
        RECT 30.200 146.800 30.600 147.200 ;
        RECT 23.000 144.800 23.400 145.200 ;
        RECT 36.600 146.800 37.000 147.200 ;
        RECT 29.400 143.800 29.800 144.200 ;
        RECT 41.400 144.800 41.800 145.200 ;
        RECT 51.800 145.800 52.200 146.200 ;
        RECT 57.400 146.800 57.800 147.200 ;
        RECT 58.200 146.800 58.600 147.200 ;
        RECT 59.000 145.800 59.400 146.200 ;
        RECT 49.400 141.800 49.800 142.200 ;
        RECT 55.000 145.100 55.400 145.500 ;
        RECT 66.200 145.800 66.600 146.200 ;
        RECT 63.800 143.800 64.200 144.200 ;
        RECT 77.400 146.800 77.800 147.200 ;
        RECT 73.400 144.800 73.800 145.200 ;
        RECT 78.200 145.800 78.600 146.200 ;
        RECT 84.600 148.800 85.000 149.200 ;
        RECT 91.000 148.800 91.400 149.200 ;
        RECT 80.600 145.800 81.000 146.200 ;
        RECT 96.600 148.800 97.000 149.200 ;
        RECT 91.000 145.800 91.400 146.200 ;
        RECT 92.600 144.800 93.000 145.200 ;
        RECT 83.800 143.800 84.200 144.200 ;
        RECT 91.800 143.800 92.200 144.200 ;
        RECT 91.000 141.800 91.400 142.200 ;
        RECT 93.400 141.800 93.800 142.200 ;
        RECT 100.600 148.800 101.000 149.200 ;
        RECT 106.200 148.800 106.600 149.200 ;
        RECT 101.400 145.800 101.800 146.200 ;
        RECT 99.000 144.800 99.400 145.200 ;
        RECT 102.200 144.800 102.600 145.200 ;
        RECT 104.600 144.800 105.000 145.200 ;
        RECT 109.400 145.800 109.800 146.200 ;
        RECT 112.600 145.800 113.000 146.200 ;
        RECT 120.600 148.800 121.000 149.200 ;
        RECT 116.600 146.800 117.000 147.200 ;
        RECT 100.600 141.800 101.000 142.200 ;
        RECT 113.400 144.800 113.800 145.200 ;
        RECT 111.800 142.800 112.200 143.200 ;
        RECT 121.400 144.800 121.800 145.200 ;
        RECT 123.800 144.800 124.200 145.200 ;
        RECT 126.200 144.800 126.600 145.200 ;
        RECT 131.800 145.800 132.200 146.200 ;
        RECT 131.000 144.800 131.400 145.200 ;
        RECT 133.400 148.800 133.800 149.200 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 132.600 141.800 133.000 142.200 ;
        RECT 136.600 144.800 137.000 145.200 ;
        RECT 139.000 146.800 139.400 147.200 ;
        RECT 142.200 146.800 142.600 147.200 ;
        RECT 147.000 146.800 147.400 147.200 ;
        RECT 143.800 144.800 144.200 145.200 ;
        RECT 149.400 145.800 149.800 146.200 ;
        RECT 164.600 148.800 165.000 149.200 ;
        RECT 156.600 145.800 157.000 146.200 ;
        RECT 160.600 145.800 161.000 146.200 ;
        RECT 154.200 143.800 154.600 144.200 ;
        RECT 152.600 141.800 153.000 142.200 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 172.600 146.800 173.000 147.200 ;
        RECT 167.000 146.100 167.400 146.500 ;
        RECT 162.200 141.800 162.600 142.200 ;
        RECT 171.000 145.900 171.400 146.300 ;
        RECT 175.800 145.800 176.200 146.200 ;
        RECT 173.400 145.100 173.800 145.500 ;
        RECT 177.400 144.800 177.800 145.200 ;
        RECT 187.800 146.800 188.200 147.200 ;
        RECT 205.400 148.800 205.800 149.200 ;
        RECT 182.200 146.100 182.600 146.500 ;
        RECT 193.400 145.800 193.800 146.200 ;
        RECT 188.600 145.100 189.000 145.500 ;
        RECT 192.600 144.800 193.000 145.200 ;
        RECT 194.200 144.800 194.600 145.200 ;
        RECT 199.000 145.900 199.400 146.300 ;
        RECT 196.600 145.100 197.000 145.500 ;
        RECT 216.600 148.800 217.000 149.200 ;
        RECT 210.200 145.900 210.600 146.300 ;
        RECT 206.200 141.800 206.600 142.200 ;
        RECT 207.800 145.100 208.200 145.500 ;
        RECT 223.800 146.800 224.200 147.200 ;
        RECT 224.600 146.800 225.000 147.200 ;
        RECT 219.800 145.800 220.200 146.200 ;
        RECT 223.000 145.900 223.400 146.300 ;
        RECT 219.800 144.800 220.200 145.200 ;
        RECT 220.600 145.100 221.000 145.500 ;
        RECT 229.400 141.800 229.800 142.200 ;
        RECT 10.200 136.800 10.600 137.200 ;
        RECT 3.800 134.800 4.200 135.200 ;
        RECT 0.600 133.100 1.000 133.500 ;
        RECT 24.600 138.800 25.000 139.200 ;
        RECT 10.200 133.800 10.600 134.200 ;
        RECT 14.200 134.800 14.600 135.200 ;
        RECT 20.600 134.800 21.000 135.200 ;
        RECT 15.000 133.800 15.400 134.200 ;
        RECT 16.600 133.800 17.000 134.200 ;
        RECT 15.800 133.100 16.200 133.500 ;
        RECT 18.200 132.800 18.600 133.200 ;
        RECT 37.400 137.800 37.800 138.200 ;
        RECT 26.200 134.800 26.600 135.200 ;
        RECT 27.000 134.800 27.400 135.200 ;
        RECT 32.600 134.800 33.000 135.200 ;
        RECT 29.400 133.800 29.800 134.200 ;
        RECT 28.600 133.100 29.000 133.500 ;
        RECT 41.400 134.800 41.800 135.200 ;
        RECT 44.600 134.800 45.000 135.200 ;
        RECT 45.400 133.800 45.800 134.200 ;
        RECT 47.800 133.800 48.200 134.200 ;
        RECT 72.600 138.800 73.000 139.200 ;
        RECT 51.000 134.800 51.400 135.200 ;
        RECT 55.000 134.800 55.400 135.200 ;
        RECT 51.800 133.100 52.200 133.500 ;
        RECT 61.400 133.800 61.800 134.200 ;
        RECT 67.800 134.800 68.200 135.200 ;
        RECT 64.600 133.800 65.000 134.200 ;
        RECT 63.800 133.100 64.200 133.500 ;
        RECT 60.600 131.800 61.000 132.200 ;
        RECT 75.000 134.800 75.400 135.200 ;
        RECT 75.800 133.800 76.200 134.200 ;
        RECT 80.600 136.800 81.000 137.200 ;
        RECT 79.000 135.800 79.400 136.200 ;
        RECT 83.000 134.800 83.400 135.200 ;
        RECT 83.800 134.800 84.200 135.200 ;
        RECT 99.800 138.800 100.200 139.200 ;
        RECT 103.800 136.800 104.200 137.200 ;
        RECT 78.200 133.800 78.600 134.200 ;
        RECT 72.600 131.800 73.000 132.200 ;
        RECT 87.800 133.800 88.200 134.200 ;
        RECT 87.000 133.100 87.400 133.500 ;
        RECT 96.600 132.800 97.000 133.200 ;
        RECT 95.800 131.800 96.200 132.200 ;
        RECT 102.200 135.800 102.600 136.200 ;
        RECT 105.400 135.800 105.800 136.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 117.400 138.800 117.800 139.200 ;
        RECT 120.600 138.800 121.000 139.200 ;
        RECT 112.600 136.800 113.000 137.200 ;
        RECT 116.600 136.800 117.000 137.200 ;
        RECT 119.800 136.800 120.200 137.200 ;
        RECT 123.000 138.800 123.400 139.200 ;
        RECT 122.200 136.800 122.600 137.200 ;
        RECT 125.400 136.800 125.800 137.200 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 115.000 135.800 115.400 136.200 ;
        RECT 119.000 135.800 119.400 136.200 ;
        RECT 113.400 134.800 113.800 135.200 ;
        RECT 104.600 131.800 105.000 132.200 ;
        RECT 107.800 131.800 108.200 132.200 ;
        RECT 123.800 135.800 124.200 136.200 ;
        RECT 123.000 134.800 123.400 135.200 ;
        RECT 127.000 135.800 127.400 136.200 ;
        RECT 126.200 134.800 126.600 135.200 ;
        RECT 131.000 135.800 131.400 136.200 ;
        RECT 127.800 132.800 128.200 133.200 ;
        RECT 126.200 131.800 126.600 132.200 ;
        RECT 132.600 134.800 133.000 135.200 ;
        RECT 133.400 133.800 133.800 134.200 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 143.000 135.800 143.400 136.200 ;
        RECT 138.200 134.800 138.600 135.200 ;
        RECT 143.000 134.800 143.400 135.200 ;
        RECT 145.400 134.800 145.800 135.200 ;
        RECT 148.600 135.800 149.000 136.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 146.200 133.800 146.600 134.200 ;
        RECT 135.000 131.800 135.400 132.200 ;
        RECT 138.200 131.800 138.600 132.200 ;
        RECT 158.200 134.800 158.600 135.200 ;
        RECT 153.400 133.800 153.800 134.200 ;
        RECT 148.600 132.800 149.000 133.200 ;
        RECT 150.200 131.800 150.600 132.200 ;
        RECT 158.200 133.800 158.600 134.200 ;
        RECT 159.000 133.800 159.400 134.200 ;
        RECT 161.400 133.800 161.800 134.200 ;
        RECT 165.400 136.800 165.800 137.200 ;
        RECT 163.800 135.800 164.200 136.200 ;
        RECT 170.200 134.800 170.600 135.200 ;
        RECT 171.000 134.800 171.400 135.200 ;
        RECT 174.200 134.800 174.600 135.200 ;
        RECT 166.200 133.800 166.600 134.200 ;
        RECT 160.600 131.800 161.000 132.200 ;
        RECT 169.400 133.800 169.800 134.200 ;
        RECT 175.800 133.800 176.200 134.200 ;
        RECT 183.000 138.800 183.400 139.200 ;
        RECT 184.600 136.800 185.000 137.200 ;
        RECT 178.200 133.800 178.600 134.200 ;
        RECT 179.000 133.800 179.400 134.200 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 183.000 134.800 183.400 135.200 ;
        RECT 183.800 133.800 184.200 134.200 ;
        RECT 188.600 136.800 189.000 137.200 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 195.800 136.200 196.200 136.600 ;
        RECT 197.400 135.500 197.800 135.900 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 185.400 131.800 185.800 132.200 ;
        RECT 197.400 133.100 197.800 133.500 ;
        RECT 200.600 133.800 201.000 134.200 ;
        RECT 198.200 131.800 198.600 132.200 ;
        RECT 208.600 136.800 209.000 137.200 ;
        RECT 207.000 135.800 207.400 136.200 ;
        RECT 203.000 133.800 203.400 134.200 ;
        RECT 207.000 134.800 207.400 135.200 ;
        RECT 207.800 133.800 208.200 134.200 ;
        RECT 215.800 136.200 216.200 136.600 ;
        RECT 217.400 135.500 217.800 135.900 ;
        RECT 221.400 134.800 221.800 135.200 ;
        RECT 201.400 131.800 201.800 132.200 ;
        RECT 217.400 133.100 217.800 133.500 ;
        RECT 218.200 133.100 218.600 133.500 ;
        RECT 227.000 131.800 227.400 132.200 ;
        RECT 11.800 126.800 12.200 127.200 ;
        RECT 6.200 126.100 6.600 126.500 ;
        RECT 2.200 124.800 2.600 125.200 ;
        RECT 12.600 125.100 13.000 125.500 ;
        RECT 3.800 121.800 4.200 122.200 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 19.000 125.800 19.400 126.200 ;
        RECT 14.200 121.800 14.600 122.200 ;
        RECT 15.000 125.100 15.400 125.500 ;
        RECT 23.800 121.800 24.200 122.200 ;
        RECT 42.200 128.800 42.600 129.200 ;
        RECT 33.400 126.800 33.800 127.200 ;
        RECT 27.800 125.800 28.200 126.200 ;
        RECT 25.400 121.800 25.800 122.200 ;
        RECT 32.600 125.100 33.000 125.500 ;
        RECT 43.800 121.800 44.200 122.200 ;
        RECT 53.400 128.800 53.800 129.200 ;
        RECT 49.400 121.800 49.800 122.200 ;
        RECT 54.200 124.800 54.600 125.200 ;
        RECT 74.200 127.800 74.600 128.200 ;
        RECT 69.400 125.800 69.800 126.200 ;
        RECT 64.600 121.800 65.000 122.200 ;
        RECT 65.400 125.100 65.800 125.500 ;
        RECT 77.400 127.800 77.800 128.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 80.600 126.800 81.000 127.200 ;
        RECT 87.000 126.800 87.400 127.200 ;
        RECT 86.200 125.900 86.600 126.300 ;
        RECT 81.400 124.800 81.800 125.200 ;
        RECT 83.800 125.100 84.200 125.500 ;
        RECT 95.000 124.800 95.400 125.200 ;
        RECT 92.600 121.800 93.000 122.200 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 115.000 128.800 115.400 129.200 ;
        RECT 97.400 125.800 97.800 126.200 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 118.200 126.800 118.600 127.200 ;
        RECT 134.200 128.800 134.600 129.200 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 101.400 121.800 101.800 122.200 ;
        RECT 104.600 121.800 105.000 122.200 ;
        RECT 115.000 125.800 115.400 126.200 ;
        RECT 118.200 125.800 118.600 126.200 ;
        RECT 128.600 126.800 129.000 127.200 ;
        RECT 124.600 125.800 125.000 126.200 ;
        RECT 129.400 125.800 129.800 126.200 ;
        RECT 125.400 125.100 125.800 125.500 ;
        RECT 111.800 121.800 112.200 122.200 ;
        RECT 113.400 121.800 113.800 122.200 ;
        RECT 119.800 121.800 120.200 122.200 ;
        RECT 123.000 121.800 123.400 122.200 ;
        RECT 142.200 125.800 142.600 126.200 ;
        RECT 139.800 124.800 140.200 125.200 ;
        RECT 152.600 128.800 153.000 129.200 ;
        RECT 147.000 124.800 147.400 125.200 ;
        RECT 146.200 121.800 146.600 122.200 ;
        RECT 171.800 128.800 172.200 129.200 ;
        RECT 155.000 126.100 155.400 126.500 ;
        RECT 159.000 125.900 159.400 126.300 ;
        RECT 161.400 125.100 161.800 125.500 ;
        RECT 167.000 125.800 167.400 126.200 ;
        RECT 165.400 121.800 165.800 122.200 ;
        RECT 179.800 128.800 180.200 129.200 ;
        RECT 170.200 124.800 170.600 125.200 ;
        RECT 176.600 126.800 177.000 127.200 ;
        RECT 174.200 125.800 174.600 126.200 ;
        RECT 177.400 124.800 177.800 125.200 ;
        RECT 189.400 128.800 189.800 129.200 ;
        RECT 195.800 128.800 196.200 129.200 ;
        RECT 187.800 126.800 188.200 127.200 ;
        RECT 193.400 126.800 193.800 127.200 ;
        RECT 182.200 126.100 182.600 126.500 ;
        RECT 188.600 125.100 189.000 125.500 ;
        RECT 203.800 128.800 204.200 129.200 ;
        RECT 203.000 126.800 203.400 127.200 ;
        RECT 200.600 125.800 201.000 126.200 ;
        RECT 219.000 128.800 219.400 129.200 ;
        RECT 213.400 126.800 213.800 127.200 ;
        RECT 218.200 125.800 218.600 126.200 ;
        RECT 215.000 124.800 215.400 125.200 ;
        RECT 223.800 126.800 224.200 127.200 ;
        RECT 221.400 126.100 221.800 126.500 ;
        RECT 227.800 125.100 228.200 125.500 ;
        RECT 1.400 118.800 1.800 119.200 ;
        RECT 13.400 116.800 13.800 117.200 ;
        RECT 7.800 114.800 8.200 115.200 ;
        RECT 4.600 113.100 5.000 113.500 ;
        RECT 15.000 114.800 15.400 115.200 ;
        RECT 15.800 114.800 16.200 115.200 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 19.800 113.800 20.200 114.200 ;
        RECT 20.600 112.800 21.000 113.200 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 24.600 114.800 25.000 115.200 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 25.400 113.800 25.800 114.200 ;
        RECT 21.400 111.800 21.800 112.200 ;
        RECT 23.000 111.800 23.400 112.200 ;
        RECT 27.000 111.800 27.400 112.200 ;
        RECT 35.000 114.800 35.400 115.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 44.600 118.800 45.000 119.200 ;
        RECT 40.600 114.800 41.000 115.200 ;
        RECT 31.000 112.800 31.400 113.200 ;
        RECT 32.600 112.800 33.000 113.200 ;
        RECT 47.000 114.800 47.400 115.200 ;
        RECT 51.000 114.800 51.400 115.200 ;
        RECT 37.400 111.800 37.800 112.200 ;
        RECT 51.800 113.800 52.200 114.200 ;
        RECT 59.800 116.200 60.200 116.600 ;
        RECT 61.400 115.500 61.800 115.900 ;
        RECT 61.400 113.100 61.800 113.500 ;
        RECT 52.600 111.800 53.000 112.200 ;
        RECT 63.800 113.800 64.200 114.200 ;
        RECT 69.400 114.800 69.800 115.200 ;
        RECT 73.400 114.800 73.800 115.200 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 77.400 114.800 77.800 115.200 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 64.600 112.800 65.000 113.200 ;
        RECT 74.200 113.800 74.600 114.200 ;
        RECT 67.000 111.800 67.400 112.200 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 81.400 118.800 81.800 119.200 ;
        RECT 80.600 113.800 81.000 114.200 ;
        RECT 79.800 112.800 80.200 113.200 ;
        RECT 83.000 116.800 83.400 117.200 ;
        RECT 90.200 116.200 90.600 116.600 ;
        RECT 91.800 115.500 92.200 115.900 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 91.800 113.100 92.200 113.500 ;
        RECT 98.200 114.800 98.600 115.200 ;
        RECT 99.000 113.800 99.400 114.200 ;
        RECT 99.800 113.800 100.200 114.200 ;
        RECT 102.200 116.800 102.600 117.200 ;
        RECT 105.400 114.800 105.800 115.200 ;
        RECT 103.800 113.800 104.200 114.200 ;
        RECT 110.200 118.800 110.600 119.200 ;
        RECT 109.400 113.800 109.800 114.200 ;
        RECT 101.400 111.800 101.800 112.200 ;
        RECT 107.000 111.800 107.400 112.200 ;
        RECT 111.000 112.800 111.400 113.200 ;
        RECT 117.400 116.800 117.800 117.200 ;
        RECT 124.600 118.800 125.000 119.200 ;
        RECT 123.800 116.800 124.200 117.200 ;
        RECT 119.000 115.800 119.400 116.200 ;
        RECT 118.200 114.800 118.600 115.200 ;
        RECT 123.000 115.800 123.400 116.200 ;
        RECT 113.400 113.800 113.800 114.200 ;
        RECT 115.800 112.800 116.200 113.200 ;
        RECT 118.200 111.800 118.600 112.200 ;
        RECT 131.000 116.800 131.400 117.200 ;
        RECT 127.000 113.800 127.400 114.200 ;
        RECT 126.200 111.800 126.600 112.200 ;
        RECT 138.200 116.200 138.600 116.600 ;
        RECT 139.800 115.500 140.200 115.900 ;
        RECT 129.400 111.800 129.800 112.200 ;
        RECT 142.200 113.800 142.600 114.200 ;
        RECT 139.800 113.100 140.200 113.500 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 147.800 112.800 148.200 113.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 153.400 113.800 153.800 114.200 ;
        RECT 157.400 114.800 157.800 115.200 ;
        RECT 155.000 113.800 155.400 114.200 ;
        RECT 156.600 113.800 157.000 114.200 ;
        RECT 158.200 113.800 158.600 114.200 ;
        RECT 159.000 113.800 159.400 114.200 ;
        RECT 162.200 118.800 162.600 119.200 ;
        RECT 175.000 115.800 175.400 116.200 ;
        RECT 173.400 114.800 173.800 115.200 ;
        RECT 151.800 111.800 152.200 112.200 ;
        RECT 154.200 111.800 154.600 112.200 ;
        RECT 160.600 111.800 161.000 112.200 ;
        RECT 168.600 111.800 169.000 112.200 ;
        RECT 171.000 111.800 171.400 112.200 ;
        RECT 175.800 113.800 176.200 114.200 ;
        RECT 179.800 114.800 180.200 115.200 ;
        RECT 180.600 114.800 181.000 115.200 ;
        RECT 202.200 116.800 202.600 117.200 ;
        RECT 184.600 113.800 185.000 114.200 ;
        RECT 188.600 114.800 189.000 115.200 ;
        RECT 192.600 114.800 193.000 115.200 ;
        RECT 191.800 113.800 192.200 114.200 ;
        RECT 193.400 113.100 193.800 113.500 ;
        RECT 206.200 114.800 206.600 115.200 ;
        RECT 207.000 114.800 207.400 115.200 ;
        RECT 207.800 113.800 208.200 114.200 ;
        RECT 210.200 118.800 210.600 119.200 ;
        RECT 217.400 116.200 217.800 116.600 ;
        RECT 219.000 115.500 219.400 115.900 ;
        RECT 223.000 114.800 223.400 115.200 ;
        RECT 216.600 112.800 217.000 113.200 ;
        RECT 219.000 113.100 219.400 113.500 ;
        RECT 219.800 113.100 220.200 113.500 ;
        RECT 222.200 112.800 222.600 113.200 ;
        RECT 228.600 111.800 229.000 112.200 ;
        RECT 1.400 108.800 1.800 109.200 ;
        RECT 0.600 104.800 1.000 105.200 ;
        RECT 19.000 108.800 19.400 109.200 ;
        RECT 11.000 106.800 11.400 107.200 ;
        RECT 29.400 108.800 29.800 109.200 ;
        RECT 9.400 105.800 9.800 106.200 ;
        RECT 15.000 105.800 15.400 106.200 ;
        RECT 6.200 104.800 6.600 105.200 ;
        RECT 8.600 104.800 9.000 105.200 ;
        RECT 10.200 105.100 10.600 105.500 ;
        RECT 21.400 105.800 21.800 106.200 ;
        RECT 23.000 104.800 23.400 105.200 ;
        RECT 27.800 104.800 28.200 105.200 ;
        RECT 37.400 105.900 37.800 106.300 ;
        RECT 35.000 105.100 35.400 105.500 ;
        RECT 33.400 101.800 33.800 102.200 ;
        RECT 56.600 108.800 57.000 109.200 ;
        RECT 48.600 106.800 49.000 107.200 ;
        RECT 52.600 105.800 53.000 106.200 ;
        RECT 43.800 101.800 44.200 102.200 ;
        RECT 47.800 105.100 48.200 105.500 ;
        RECT 46.200 101.800 46.600 102.200 ;
        RECT 65.400 106.800 65.800 107.200 ;
        RECT 70.200 106.800 70.600 107.200 ;
        RECT 59.000 103.800 59.400 104.200 ;
        RECT 60.600 104.800 61.000 105.200 ;
        RECT 64.600 105.100 65.000 105.500 ;
        RECT 97.400 108.800 97.800 109.200 ;
        RECT 78.200 105.800 78.600 106.200 ;
        RECT 79.000 105.800 79.400 106.200 ;
        RECT 73.400 103.800 73.800 104.200 ;
        RECT 79.800 103.800 80.200 104.200 ;
        RECT 83.000 104.800 83.400 105.200 ;
        RECT 88.600 105.100 89.000 105.500 ;
        RECT 112.600 108.800 113.000 109.200 ;
        RECT 114.200 108.800 114.600 109.200 ;
        RECT 106.200 106.800 106.600 107.200 ;
        RECT 101.400 104.800 101.800 105.200 ;
        RECT 103.800 105.100 104.200 105.500 ;
        RECT 119.000 108.800 119.400 109.200 ;
        RECT 115.800 105.800 116.200 106.200 ;
        RECT 120.600 105.800 121.000 106.200 ;
        RECT 123.800 106.800 124.200 107.200 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 114.200 101.800 114.600 102.200 ;
        RECT 126.200 104.800 126.600 105.200 ;
        RECT 127.800 105.100 128.200 105.500 ;
        RECT 139.000 106.800 139.400 107.200 ;
        RECT 136.600 103.800 137.000 104.200 ;
        RECT 142.200 104.800 142.600 105.200 ;
        RECT 155.000 107.800 155.400 108.200 ;
        RECT 146.200 105.800 146.600 106.200 ;
        RECT 147.800 104.800 148.200 105.200 ;
        RECT 151.800 104.800 152.200 105.200 ;
        RECT 155.000 105.800 155.400 106.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 154.200 104.800 154.600 105.200 ;
        RECT 167.000 108.800 167.400 109.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 159.000 104.800 159.400 105.200 ;
        RECT 165.400 101.800 165.800 102.200 ;
        RECT 175.000 106.800 175.400 107.200 ;
        RECT 171.000 106.100 171.400 106.500 ;
        RECT 177.400 105.100 177.800 105.500 ;
        RECT 179.800 104.800 180.200 105.200 ;
        RECT 188.600 106.800 189.000 107.200 ;
        RECT 185.400 104.800 185.800 105.200 ;
        RECT 210.200 108.800 210.600 109.200 ;
        RECT 189.400 104.800 189.800 105.200 ;
        RECT 201.400 106.800 201.800 107.200 ;
        RECT 195.800 106.100 196.200 106.500 ;
        RECT 209.400 105.800 209.800 106.200 ;
        RECT 202.200 105.100 202.600 105.500 ;
        RECT 228.600 108.800 229.000 109.200 ;
        RECT 220.600 106.800 221.000 107.200 ;
        RECT 212.600 106.100 213.000 106.500 ;
        RECT 209.400 104.800 209.800 105.200 ;
        RECT 219.000 105.100 219.400 105.500 ;
        RECT 219.800 105.100 220.200 105.500 ;
        RECT 0.600 98.800 1.000 99.200 ;
        RECT 7.800 96.200 8.200 96.600 ;
        RECT 9.400 95.500 9.800 95.900 ;
        RECT 4.600 93.800 5.000 94.200 ;
        RECT 10.200 93.800 10.600 94.200 ;
        RECT 9.400 93.100 9.800 93.500 ;
        RECT 14.200 94.800 14.600 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 30.200 96.800 30.600 97.200 ;
        RECT 15.000 93.800 15.400 94.200 ;
        RECT 19.000 93.800 19.400 94.200 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 21.400 93.100 21.800 93.500 ;
        RECT 32.600 93.800 33.000 94.200 ;
        RECT 31.000 92.800 31.400 93.200 ;
        RECT 31.800 92.800 32.200 93.200 ;
        RECT 39.000 94.800 39.400 95.200 ;
        RECT 50.200 96.800 50.600 97.200 ;
        RECT 45.400 95.800 45.800 96.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 35.000 92.800 35.400 93.200 ;
        RECT 41.400 92.800 41.800 93.200 ;
        RECT 52.600 96.800 53.000 97.200 ;
        RECT 55.800 94.800 56.200 95.200 ;
        RECT 65.400 96.800 65.800 97.200 ;
        RECT 67.800 96.800 68.200 97.200 ;
        RECT 61.400 94.800 61.800 95.200 ;
        RECT 54.200 93.800 54.600 94.200 ;
        RECT 51.800 91.800 52.200 92.200 ;
        RECT 57.400 92.800 57.800 93.200 ;
        RECT 58.200 93.100 58.600 93.500 ;
        RECT 74.200 98.800 74.600 99.200 ;
        RECT 79.800 98.800 80.200 99.200 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 71.800 94.800 72.200 95.200 ;
        RECT 72.600 93.800 73.000 94.200 ;
        RECT 75.800 94.800 76.200 95.200 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 79.000 94.800 79.400 95.200 ;
        RECT 87.000 96.200 87.400 96.600 ;
        RECT 88.600 95.500 89.000 95.900 ;
        RECT 88.600 93.100 89.000 93.500 ;
        RECT 79.800 91.800 80.200 92.200 ;
        RECT 95.000 98.800 95.400 99.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 94.200 96.800 94.600 97.200 ;
        RECT 95.800 95.800 96.200 96.200 ;
        RECT 95.000 94.800 95.400 95.200 ;
        RECT 92.600 91.800 93.000 92.200 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 99.000 93.800 99.400 94.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 108.600 93.800 109.000 94.200 ;
        RECT 112.600 94.800 113.000 95.200 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 100.600 91.800 101.000 92.200 ;
        RECT 120.600 98.800 121.000 99.200 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 119.800 94.800 120.200 95.200 ;
        RECT 115.000 91.800 115.400 92.200 ;
        RECT 117.400 91.800 117.800 92.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 120.600 91.800 121.000 92.200 ;
        RECT 129.400 98.800 129.800 99.200 ;
        RECT 125.400 93.800 125.800 94.200 ;
        RECT 123.800 91.800 124.200 92.200 ;
        RECT 127.000 91.800 127.400 92.200 ;
        RECT 130.200 92.800 130.600 93.200 ;
        RECT 152.600 98.800 153.000 99.200 ;
        RECT 135.800 94.800 136.200 95.200 ;
        RECT 142.200 94.800 142.600 95.200 ;
        RECT 132.600 93.800 133.000 94.200 ;
        RECT 135.800 93.800 136.200 94.200 ;
        RECT 138.200 93.100 138.600 93.500 ;
        RECT 159.000 98.800 159.400 99.200 ;
        RECT 149.400 94.800 149.800 95.200 ;
        RECT 152.600 94.800 153.000 95.200 ;
        RECT 150.200 93.800 150.600 94.200 ;
        RECT 154.200 93.800 154.600 94.200 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 155.000 91.800 155.400 92.200 ;
        RECT 160.600 93.100 161.000 93.500 ;
        RECT 174.200 94.800 174.600 95.200 ;
        RECT 169.400 91.800 169.800 92.200 ;
        RECT 170.200 93.100 170.600 93.500 ;
        RECT 184.600 93.800 185.000 94.200 ;
        RECT 179.000 91.800 179.400 92.200 ;
        RECT 187.800 94.800 188.200 95.200 ;
        RECT 188.600 93.800 189.000 94.200 ;
        RECT 186.200 91.800 186.600 92.200 ;
        RECT 191.800 96.800 192.200 97.200 ;
        RECT 195.800 94.800 196.200 95.200 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 214.200 96.800 214.600 97.200 ;
        RECT 202.200 94.800 202.600 95.200 ;
        RECT 222.200 96.800 222.600 97.200 ;
        RECT 223.800 96.800 224.200 97.200 ;
        RECT 203.800 94.800 204.200 95.200 ;
        RECT 204.600 93.800 205.000 94.200 ;
        RECT 206.200 93.800 206.600 94.200 ;
        RECT 205.400 93.100 205.800 93.500 ;
        RECT 215.800 93.800 216.200 94.200 ;
        RECT 215.000 93.100 215.400 93.500 ;
        RECT 227.000 94.800 227.400 95.200 ;
        RECT 9.400 88.800 9.800 89.200 ;
        RECT 38.200 88.800 38.600 89.200 ;
        RECT 4.600 86.800 5.000 87.200 ;
        RECT 4.600 85.800 5.000 86.200 ;
        RECT 0.600 85.100 1.000 85.500 ;
        RECT 16.600 86.800 17.000 87.200 ;
        RECT 30.200 86.800 30.600 87.200 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 31.800 85.900 32.200 86.300 ;
        RECT 19.000 83.800 19.400 84.200 ;
        RECT 21.400 81.800 21.800 82.200 ;
        RECT 25.400 84.800 25.800 85.200 ;
        RECT 28.600 84.800 29.000 85.200 ;
        RECT 29.400 85.100 29.800 85.500 ;
        RECT 51.800 88.800 52.200 89.200 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 48.600 86.800 49.000 87.200 ;
        RECT 42.200 84.800 42.600 85.200 ;
        RECT 43.000 85.100 43.400 85.500 ;
        RECT 54.200 85.800 54.600 86.200 ;
        RECT 55.800 84.800 56.200 85.200 ;
        RECT 63.000 86.800 63.400 87.200 ;
        RECT 69.400 88.800 69.800 89.200 ;
        RECT 64.600 85.800 65.000 86.200 ;
        RECT 59.000 81.800 59.400 82.200 ;
        RECT 62.200 81.800 62.600 82.200 ;
        RECT 79.000 88.800 79.400 89.200 ;
        RECT 107.800 88.800 108.200 89.200 ;
        RECT 67.800 84.800 68.200 85.200 ;
        RECT 69.400 81.800 69.800 82.200 ;
        RECT 81.400 86.100 81.800 86.500 ;
        RECT 85.400 85.900 85.800 86.300 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 87.800 85.100 88.200 85.500 ;
        RECT 79.000 81.800 79.400 82.200 ;
        RECT 92.600 84.800 93.000 85.200 ;
        RECT 95.000 84.800 95.400 85.200 ;
        RECT 101.400 85.900 101.800 86.300 ;
        RECT 98.200 84.800 98.600 85.200 ;
        RECT 99.000 85.100 99.400 85.500 ;
        RECT 112.600 86.800 113.000 87.200 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 130.200 88.800 130.600 89.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 111.000 84.800 111.400 85.200 ;
        RECT 117.400 84.800 117.800 85.200 ;
        RECT 120.600 84.800 121.000 85.200 ;
        RECT 121.400 85.100 121.800 85.500 ;
        RECT 131.000 88.800 131.400 89.200 ;
        RECT 148.600 88.800 149.000 89.200 ;
        RECT 133.400 86.100 133.800 86.500 ;
        RECT 137.400 85.900 137.800 86.300 ;
        RECT 139.800 85.100 140.200 85.500 ;
        RECT 143.800 84.800 144.200 85.200 ;
        RECT 147.800 84.800 148.200 85.200 ;
        RECT 160.600 88.800 161.000 89.200 ;
        RECT 153.400 86.800 153.800 87.200 ;
        RECT 156.600 86.800 157.000 87.200 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 165.400 88.800 165.800 89.200 ;
        RECT 163.000 86.800 163.400 87.200 ;
        RECT 151.000 81.800 151.400 82.200 ;
        RECT 155.000 84.800 155.400 85.200 ;
        RECT 183.000 88.800 183.400 89.200 ;
        RECT 179.000 86.800 179.400 87.200 ;
        RECT 176.600 85.800 177.000 86.200 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 164.600 81.800 165.000 82.200 ;
        RECT 175.800 84.800 176.200 85.200 ;
        RECT 179.800 85.800 180.200 86.200 ;
        RECT 183.000 84.800 183.400 85.200 ;
        RECT 183.800 84.800 184.200 85.200 ;
        RECT 187.000 85.800 187.400 86.200 ;
        RECT 195.800 86.800 196.200 87.200 ;
        RECT 192.600 85.800 193.000 86.200 ;
        RECT 206.200 86.800 206.600 87.200 ;
        RECT 188.600 81.800 189.000 82.200 ;
        RECT 195.800 84.800 196.200 85.200 ;
        RECT 200.600 86.100 201.000 86.500 ;
        RECT 207.000 85.100 207.400 85.500 ;
        RECT 224.600 88.800 225.000 89.200 ;
        RECT 220.600 86.800 221.000 87.200 ;
        RECT 215.000 86.100 215.400 86.500 ;
        RECT 219.000 85.900 219.400 86.300 ;
        RECT 221.400 85.100 221.800 85.500 ;
        RECT 223.800 84.800 224.200 85.200 ;
        RECT 229.400 84.800 229.800 85.200 ;
        RECT 9.400 76.800 9.800 77.200 ;
        RECT 4.600 74.800 5.000 75.200 ;
        RECT 0.600 73.100 1.000 73.500 ;
        RECT 11.000 74.800 11.400 75.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 30.200 78.800 30.600 79.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 21.400 73.100 21.800 73.500 ;
        RECT 31.800 74.800 32.200 75.200 ;
        RECT 33.400 74.800 33.800 75.200 ;
        RECT 32.600 73.800 33.000 74.200 ;
        RECT 35.800 72.800 36.200 73.200 ;
        RECT 36.600 72.800 37.000 73.200 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 47.800 74.800 48.200 75.200 ;
        RECT 41.400 73.800 41.800 74.200 ;
        RECT 43.000 73.800 43.400 74.200 ;
        RECT 58.200 75.800 58.600 76.200 ;
        RECT 55.800 74.800 56.200 75.200 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 38.200 71.800 38.600 72.200 ;
        RECT 49.400 71.800 49.800 72.200 ;
        RECT 55.800 73.800 56.200 74.200 ;
        RECT 59.800 74.800 60.200 75.200 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 58.200 73.800 58.600 74.200 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 78.200 76.200 78.600 76.600 ;
        RECT 79.800 75.500 80.200 75.900 ;
        RECT 83.000 74.800 83.400 75.200 ;
        RECT 83.800 74.800 84.200 75.200 ;
        RECT 53.400 71.800 53.800 72.200 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 79.800 73.100 80.200 73.500 ;
        RECT 71.000 71.800 71.400 72.200 ;
        RECT 80.600 72.800 81.000 73.200 ;
        RECT 86.200 73.800 86.600 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 97.400 76.200 97.800 76.600 ;
        RECT 99.000 75.500 99.400 75.900 ;
        RECT 106.200 76.800 106.600 77.200 ;
        RECT 99.800 74.800 100.200 75.200 ;
        RECT 100.600 74.800 101.000 75.200 ;
        RECT 104.600 75.800 105.000 76.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 99.000 73.100 99.400 73.500 ;
        RECT 114.200 78.800 114.600 79.200 ;
        RECT 117.400 78.800 117.800 79.200 ;
        RECT 115.000 76.800 115.400 77.200 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 113.400 75.800 113.800 76.200 ;
        RECT 109.400 73.800 109.800 74.200 ;
        RECT 119.800 73.800 120.200 74.200 ;
        RECT 117.400 71.800 117.800 72.200 ;
        RECT 124.600 74.800 125.000 75.200 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 126.200 73.800 126.600 74.200 ;
        RECT 121.400 71.800 121.800 72.200 ;
        RECT 125.400 73.100 125.800 73.500 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 143.800 74.800 144.200 75.200 ;
        RECT 139.800 73.800 140.200 74.200 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 148.600 73.800 149.000 74.200 ;
        RECT 134.200 71.800 134.600 72.200 ;
        RECT 147.800 73.100 148.200 73.500 ;
        RECT 156.600 71.800 157.000 72.200 ;
        RECT 159.800 78.800 160.200 79.200 ;
        RECT 170.200 78.800 170.600 79.200 ;
        RECT 164.600 74.800 165.000 75.200 ;
        RECT 178.200 78.800 178.600 79.200 ;
        RECT 181.400 78.800 181.800 79.200 ;
        RECT 180.600 76.800 181.000 77.200 ;
        RECT 160.600 73.800 161.000 74.200 ;
        RECT 158.200 71.800 158.600 72.200 ;
        RECT 161.400 73.100 161.800 73.500 ;
        RECT 175.000 74.800 175.400 75.200 ;
        RECT 175.800 73.800 176.200 74.200 ;
        RECT 182.200 75.800 182.600 76.200 ;
        RECT 193.400 78.800 193.800 79.200 ;
        RECT 181.400 74.800 181.800 75.200 ;
        RECT 183.000 73.800 183.400 74.200 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 186.200 74.800 186.600 75.200 ;
        RECT 193.400 74.800 193.800 75.200 ;
        RECT 199.800 74.800 200.200 75.200 ;
        RECT 200.600 74.800 201.000 75.200 ;
        RECT 206.200 76.800 206.600 77.200 ;
        RECT 204.600 74.800 205.000 75.200 ;
        RECT 205.400 74.800 205.800 75.200 ;
        RECT 195.800 72.800 196.200 73.200 ;
        RECT 213.400 76.200 213.800 76.600 ;
        RECT 215.000 75.500 215.400 75.900 ;
        RECT 215.800 73.800 216.200 74.200 ;
        RECT 215.000 73.100 215.400 73.500 ;
        RECT 227.000 78.800 227.400 79.200 ;
        RECT 219.800 74.800 220.200 75.200 ;
        RECT 220.600 73.800 221.000 74.200 ;
        RECT 228.600 74.800 229.000 75.200 ;
        RECT 13.400 68.800 13.800 69.200 ;
        RECT 5.400 66.800 5.800 67.200 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 3.000 63.800 3.400 64.200 ;
        RECT 4.600 65.100 5.000 65.500 ;
        RECT 31.000 68.800 31.400 69.200 ;
        RECT 13.400 61.800 13.800 62.200 ;
        RECT 21.400 64.800 21.800 65.200 ;
        RECT 22.200 65.100 22.600 65.500 ;
        RECT 35.800 67.800 36.200 68.200 ;
        RECT 39.800 68.800 40.200 69.200 ;
        RECT 34.200 64.800 34.600 65.200 ;
        RECT 50.200 68.800 50.600 69.200 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 59.800 68.800 60.200 69.200 ;
        RECT 44.600 61.800 45.000 62.200 ;
        RECT 48.600 64.800 49.000 65.200 ;
        RECT 47.000 61.800 47.400 62.200 ;
        RECT 67.000 68.800 67.400 69.200 ;
        RECT 53.400 65.900 53.800 66.300 ;
        RECT 51.000 65.100 51.400 65.500 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 61.400 61.800 61.800 62.200 ;
        RECT 64.600 64.800 65.000 65.200 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 87.800 68.800 88.200 69.200 ;
        RECT 82.200 66.800 82.600 67.200 ;
        RECT 80.600 65.900 81.000 66.300 ;
        RECT 75.800 64.800 76.200 65.200 ;
        RECT 70.200 61.800 70.600 62.200 ;
        RECT 78.200 65.100 78.600 65.500 ;
        RECT 95.000 68.800 95.400 69.200 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 91.800 61.800 92.200 62.200 ;
        RECT 100.600 66.800 101.000 67.200 ;
        RECT 108.600 68.800 109.000 69.200 ;
        RECT 103.000 65.800 103.400 66.200 ;
        RECT 98.200 64.800 98.600 65.200 ;
        RECT 108.600 64.800 109.000 65.200 ;
        RECT 109.400 64.800 109.800 65.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 123.800 66.800 124.200 67.200 ;
        RECT 114.200 64.800 114.600 65.200 ;
        RECT 115.800 64.800 116.200 65.200 ;
        RECT 129.400 68.800 129.800 69.200 ;
        RECT 122.200 64.800 122.600 65.200 ;
        RECT 131.800 66.100 132.200 66.500 ;
        RECT 149.400 68.800 149.800 69.200 ;
        RECT 128.600 64.800 129.000 65.200 ;
        RECT 138.200 65.100 138.600 65.500 ;
        RECT 155.800 66.800 156.200 67.200 ;
        RECT 149.400 64.800 149.800 65.200 ;
        RECT 153.400 65.800 153.800 66.200 ;
        RECT 159.000 66.800 159.400 67.200 ;
        RECT 164.600 68.800 165.000 69.200 ;
        RECT 169.400 68.800 169.800 69.200 ;
        RECT 162.200 66.800 162.600 67.200 ;
        RECT 168.600 66.800 169.000 67.200 ;
        RECT 160.600 61.800 161.000 62.200 ;
        RECT 183.000 68.800 183.400 69.200 ;
        RECT 177.400 66.800 177.800 67.200 ;
        RECT 163.800 63.800 164.200 64.200 ;
        RECT 176.600 65.900 177.000 66.300 ;
        RECT 174.200 65.100 174.600 65.500 ;
        RECT 183.800 64.800 184.200 65.200 ;
        RECT 187.800 64.800 188.200 65.200 ;
        RECT 211.800 68.800 212.200 69.200 ;
        RECT 201.400 66.800 201.800 67.200 ;
        RECT 195.800 66.100 196.200 66.500 ;
        RECT 190.200 61.800 190.600 62.200 ;
        RECT 199.800 65.900 200.200 66.300 ;
        RECT 204.600 65.800 205.000 66.200 ;
        RECT 202.200 65.100 202.600 65.500 ;
        RECT 193.400 61.800 193.800 62.200 ;
        RECT 207.800 64.800 208.200 65.200 ;
        RECT 225.400 66.800 225.800 67.200 ;
        RECT 214.200 66.100 214.600 66.500 ;
        RECT 220.600 65.100 221.000 65.500 ;
        RECT 221.400 65.100 221.800 65.500 ;
        RECT 230.200 61.800 230.600 62.200 ;
        RECT 12.600 56.800 13.000 57.200 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 3.800 53.100 4.200 53.500 ;
        RECT 14.200 58.800 14.600 59.200 ;
        RECT 13.400 53.800 13.800 54.200 ;
        RECT 16.600 54.800 17.000 55.200 ;
        RECT 27.000 58.800 27.400 59.200 ;
        RECT 29.400 58.800 29.800 59.200 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 28.600 53.800 29.000 54.200 ;
        RECT 31.800 54.800 32.200 55.200 ;
        RECT 34.200 55.800 34.600 56.200 ;
        RECT 44.600 56.800 45.000 57.200 ;
        RECT 39.800 54.800 40.200 55.200 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 35.800 53.100 36.200 53.500 ;
        RECT 47.000 54.800 47.400 55.200 ;
        RECT 52.600 54.800 53.000 55.200 ;
        RECT 53.400 54.800 53.800 55.200 ;
        RECT 50.200 53.800 50.600 54.200 ;
        RECT 51.000 52.800 51.400 53.200 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 59.800 54.800 60.200 55.200 ;
        RECT 71.000 58.800 71.400 59.200 ;
        RECT 61.400 53.800 61.800 54.200 ;
        RECT 62.200 53.100 62.600 53.500 ;
        RECT 84.600 58.800 85.000 59.200 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 78.200 54.800 78.600 55.200 ;
        RECT 91.000 58.800 91.400 59.200 ;
        RECT 85.400 54.800 85.800 55.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 73.400 51.800 73.800 52.200 ;
        RECT 102.200 56.800 102.600 57.200 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 103.800 58.800 104.200 59.200 ;
        RECT 94.200 53.800 94.600 54.200 ;
        RECT 93.400 53.100 93.800 53.500 ;
        RECT 108.600 58.800 109.000 59.200 ;
        RECT 107.000 56.800 107.400 57.200 ;
        RECT 104.600 53.800 105.000 54.200 ;
        RECT 107.000 53.800 107.400 54.200 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 111.000 58.800 111.400 59.200 ;
        RECT 111.000 54.800 111.400 55.200 ;
        RECT 111.800 53.800 112.200 54.200 ;
        RECT 122.200 58.800 122.600 59.200 ;
        RECT 118.200 56.800 118.600 57.200 ;
        RECT 121.400 56.800 121.800 57.200 ;
        RECT 115.800 54.800 116.200 55.200 ;
        RECT 116.600 54.800 117.000 55.200 ;
        RECT 119.800 54.800 120.200 55.200 ;
        RECT 123.000 55.800 123.400 56.200 ;
        RECT 131.800 58.800 132.200 59.200 ;
        RECT 131.000 56.800 131.400 57.200 ;
        RECT 125.400 55.800 125.800 56.200 ;
        RECT 122.200 54.800 122.600 55.200 ;
        RECT 125.400 53.800 125.800 54.200 ;
        RECT 129.400 55.800 129.800 56.200 ;
        RECT 127.800 51.800 128.200 52.200 ;
        RECT 132.600 53.800 133.000 54.200 ;
        RECT 141.400 58.800 141.800 59.200 ;
        RECT 135.000 54.800 135.400 55.200 ;
        RECT 135.800 54.800 136.200 55.200 ;
        RECT 147.800 58.800 148.200 59.200 ;
        RECT 142.200 52.800 142.600 53.200 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 144.600 53.800 145.000 54.200 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 148.600 53.800 149.000 54.200 ;
        RECT 160.600 58.800 161.000 59.200 ;
        RECT 155.000 54.800 155.400 55.200 ;
        RECT 151.000 53.800 151.400 54.200 ;
        RECT 151.800 53.100 152.200 53.500 ;
        RECT 150.200 51.800 150.600 52.200 ;
        RECT 154.200 52.800 154.600 53.200 ;
        RECT 165.400 56.800 165.800 57.200 ;
        RECT 161.400 53.800 161.800 54.200 ;
        RECT 165.400 54.800 165.800 55.200 ;
        RECT 167.000 54.800 167.400 55.200 ;
        RECT 167.800 54.800 168.200 55.200 ;
        RECT 166.200 53.800 166.600 54.200 ;
        RECT 180.600 57.800 181.000 58.200 ;
        RECT 172.600 53.800 173.000 54.200 ;
        RECT 160.600 51.800 161.000 52.200 ;
        RECT 171.800 53.100 172.200 53.500 ;
        RECT 182.200 53.800 182.600 54.200 ;
        RECT 183.800 54.800 184.200 55.200 ;
        RECT 184.600 54.800 185.000 55.200 ;
        RECT 185.400 54.800 185.800 55.200 ;
        RECT 189.400 54.800 189.800 55.200 ;
        RECT 198.200 58.800 198.600 59.200 ;
        RECT 199.800 58.800 200.200 59.200 ;
        RECT 189.400 53.800 189.800 54.200 ;
        RECT 195.000 54.800 195.400 55.200 ;
        RECT 194.200 53.800 194.600 54.200 ;
        RECT 195.800 53.800 196.200 54.200 ;
        RECT 201.400 54.800 201.800 55.200 ;
        RECT 202.200 54.800 202.600 55.200 ;
        RECT 206.200 54.800 206.600 55.200 ;
        RECT 207.000 54.800 207.400 55.200 ;
        RECT 211.000 54.800 211.400 55.200 ;
        RECT 200.600 52.800 201.000 53.200 ;
        RECT 213.400 54.800 213.800 55.200 ;
        RECT 215.000 54.800 215.400 55.200 ;
        RECT 216.600 54.800 217.000 55.200 ;
        RECT 211.800 51.800 212.200 52.200 ;
        RECT 224.600 56.200 225.000 56.600 ;
        RECT 226.200 55.500 226.600 55.900 ;
        RECT 229.400 53.800 229.800 54.200 ;
        RECT 226.200 53.100 226.600 53.500 ;
        RECT 217.400 51.800 217.800 52.200 ;
        RECT 0.600 45.100 1.000 45.500 ;
        RECT 17.400 48.800 17.800 49.200 ;
        RECT 11.800 44.800 12.200 45.200 ;
        RECT 21.400 46.800 21.800 47.200 ;
        RECT 22.200 45.800 22.600 46.200 ;
        RECT 17.400 44.800 17.800 45.200 ;
        RECT 18.200 45.100 18.600 45.500 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 46.200 48.800 46.600 49.200 ;
        RECT 29.400 44.800 29.800 45.200 ;
        RECT 32.600 45.800 33.000 46.200 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 35.000 44.800 35.400 45.200 ;
        RECT 37.400 45.100 37.800 45.500 ;
        RECT 48.600 45.800 49.000 46.200 ;
        RECT 44.600 43.800 45.000 44.200 ;
        RECT 50.200 44.800 50.600 45.200 ;
        RECT 74.200 48.800 74.600 49.200 ;
        RECT 66.200 46.800 66.600 47.200 ;
        RECT 55.000 46.100 55.400 46.500 ;
        RECT 59.000 45.900 59.400 46.300 ;
        RECT 69.400 45.800 69.800 46.200 ;
        RECT 61.400 45.100 61.800 45.500 ;
        RECT 52.600 41.800 53.000 42.200 ;
        RECT 65.400 45.100 65.800 45.500 ;
        RECT 80.600 46.800 81.000 47.200 ;
        RECT 81.400 44.800 81.800 45.200 ;
        RECT 90.200 46.800 90.600 47.200 ;
        RECT 94.200 46.800 94.600 47.200 ;
        RECT 98.200 46.800 98.600 47.200 ;
        RECT 86.200 46.100 86.600 46.500 ;
        RECT 92.600 45.100 93.000 45.500 ;
        RECT 109.400 48.800 109.800 49.200 ;
        RECT 101.400 46.800 101.800 47.200 ;
        RECT 111.000 48.800 111.400 49.200 ;
        RECT 103.000 45.900 103.400 46.300 ;
        RECT 83.800 41.800 84.200 42.200 ;
        RECT 98.200 44.800 98.600 45.200 ;
        RECT 100.600 45.100 101.000 45.500 ;
        RECT 122.200 48.800 122.600 49.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 119.800 46.800 120.200 47.200 ;
        RECT 114.200 42.800 114.600 43.200 ;
        RECT 120.600 45.800 121.000 46.200 ;
        RECT 121.400 44.800 121.800 45.200 ;
        RECT 138.200 48.800 138.600 49.200 ;
        RECT 143.800 48.800 144.200 49.200 ;
        RECT 134.200 46.800 134.600 47.200 ;
        RECT 128.600 46.100 129.000 46.500 ;
        RECT 135.000 45.100 135.400 45.500 ;
        RECT 126.200 43.800 126.600 44.200 ;
        RECT 137.400 44.800 137.800 45.200 ;
        RECT 146.200 48.800 146.600 49.200 ;
        RECT 159.800 48.800 160.200 49.200 ;
        RECT 145.400 44.800 145.800 45.200 ;
        RECT 151.800 46.800 152.200 47.200 ;
        RECT 154.200 46.800 154.600 47.200 ;
        RECT 149.400 45.800 149.800 46.200 ;
        RECT 153.400 45.900 153.800 46.300 ;
        RECT 150.200 44.800 150.600 45.200 ;
        RECT 151.000 45.100 151.400 45.500 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 179.000 48.800 179.400 49.200 ;
        RECT 186.200 48.800 186.600 49.200 ;
        RECT 166.200 44.800 166.600 45.200 ;
        RECT 171.000 46.100 171.400 46.500 ;
        RECT 172.600 45.800 173.000 46.200 ;
        RECT 177.400 45.100 177.800 45.500 ;
        RECT 180.600 45.800 181.000 46.200 ;
        RECT 184.600 45.800 185.000 46.200 ;
        RECT 191.800 46.800 192.200 47.200 ;
        RECT 201.400 48.800 201.800 49.200 ;
        RECT 188.600 46.100 189.000 46.500 ;
        RECT 192.600 45.900 193.000 46.300 ;
        RECT 195.000 45.100 195.400 45.500 ;
        RECT 215.800 48.800 216.200 49.200 ;
        RECT 219.800 48.800 220.200 49.200 ;
        RECT 203.000 45.800 203.400 46.200 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 199.000 41.800 199.400 42.200 ;
        RECT 210.200 44.800 210.600 45.200 ;
        RECT 219.000 45.800 219.400 46.200 ;
        RECT 215.800 44.800 216.200 45.200 ;
        RECT 225.400 46.800 225.800 47.200 ;
        RECT 222.200 46.100 222.600 46.500 ;
        RECT 219.000 44.800 219.400 45.200 ;
        RECT 228.600 45.100 229.000 45.500 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 3.000 32.800 3.400 33.200 ;
        RECT 14.200 38.800 14.600 39.200 ;
        RECT 12.600 34.800 13.000 35.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 19.000 34.800 19.400 35.200 ;
        RECT 7.000 31.800 7.400 32.200 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 15.000 33.800 15.400 34.200 ;
        RECT 15.800 33.100 16.200 33.500 ;
        RECT 26.200 38.800 26.600 39.200 ;
        RECT 24.600 31.800 25.000 32.200 ;
        RECT 29.400 38.800 29.800 39.200 ;
        RECT 27.800 34.800 28.200 35.200 ;
        RECT 39.800 36.800 40.200 37.200 ;
        RECT 41.400 36.800 41.800 37.200 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 33.400 33.800 33.800 34.200 ;
        RECT 31.800 32.800 32.200 33.200 ;
        RECT 32.600 33.100 33.000 33.500 ;
        RECT 56.600 38.800 57.000 39.200 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 59.800 38.800 60.200 39.200 ;
        RECT 57.400 34.800 57.800 35.200 ;
        RECT 58.200 34.800 58.600 35.200 ;
        RECT 59.000 33.800 59.400 34.200 ;
        RECT 62.200 34.800 62.600 35.200 ;
        RECT 69.400 38.800 69.800 39.200 ;
        RECT 67.800 34.800 68.200 35.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 72.600 34.800 73.000 35.200 ;
        RECT 76.600 36.800 77.000 37.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 63.800 31.800 64.200 32.200 ;
        RECT 78.200 34.800 78.600 35.200 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 89.400 36.800 89.800 37.200 ;
        RECT 82.200 33.800 82.600 34.200 ;
        RECT 86.200 34.800 86.600 35.200 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 79.800 31.800 80.200 32.200 ;
        RECT 96.600 36.200 97.000 36.600 ;
        RECT 98.200 35.500 98.600 35.900 ;
        RECT 103.000 36.800 103.400 37.200 ;
        RECT 99.000 33.800 99.400 34.200 ;
        RECT 98.200 33.100 98.600 33.500 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 103.800 33.800 104.200 34.200 ;
        RECT 109.400 38.800 109.800 39.200 ;
        RECT 107.000 34.800 107.400 35.200 ;
        RECT 107.800 34.800 108.200 35.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 123.000 38.800 123.400 39.200 ;
        RECT 115.800 34.800 116.200 35.200 ;
        RECT 118.200 34.800 118.600 35.200 ;
        RECT 132.600 38.800 133.000 39.200 ;
        RECT 116.600 33.800 117.000 34.200 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 124.600 34.800 125.000 35.200 ;
        RECT 125.400 34.800 125.800 35.200 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 129.400 34.800 129.800 35.200 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 131.000 34.800 131.400 35.200 ;
        RECT 105.400 31.800 105.800 32.200 ;
        RECT 114.200 31.800 114.600 32.200 ;
        RECT 128.600 33.800 129.000 34.200 ;
        RECT 142.200 36.800 142.600 37.200 ;
        RECT 139.000 35.800 139.400 36.200 ;
        RECT 135.000 33.800 135.400 34.200 ;
        RECT 139.000 34.800 139.400 35.200 ;
        RECT 139.800 33.800 140.200 34.200 ;
        RECT 149.400 36.200 149.800 36.600 ;
        RECT 153.400 38.800 153.800 39.200 ;
        RECT 151.000 35.500 151.400 35.900 ;
        RECT 152.600 34.800 153.000 35.200 ;
        RECT 154.200 34.800 154.600 35.200 ;
        RECT 159.000 34.800 159.400 35.200 ;
        RECT 160.600 34.800 161.000 35.200 ;
        RECT 151.000 33.100 151.400 33.500 ;
        RECT 160.600 33.800 161.000 34.200 ;
        RECT 163.000 33.800 163.400 34.200 ;
        RECT 168.600 38.800 169.000 39.200 ;
        RECT 167.800 32.800 168.200 33.200 ;
        RECT 171.000 33.800 171.400 34.200 ;
        RECT 169.400 32.800 169.800 33.200 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 173.400 33.800 173.800 34.200 ;
        RECT 183.800 38.800 184.200 39.200 ;
        RECT 177.400 34.800 177.800 35.200 ;
        RECT 179.000 34.800 179.400 35.200 ;
        RECT 179.800 34.800 180.200 35.200 ;
        RECT 178.200 33.800 178.600 34.200 ;
        RECT 183.000 34.800 183.400 35.200 ;
        RECT 182.200 33.800 182.600 34.200 ;
        RECT 175.800 31.800 176.200 32.200 ;
        RECT 192.600 36.200 193.000 36.600 ;
        RECT 194.200 35.500 194.600 35.900 ;
        RECT 197.400 34.800 197.800 35.200 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 200.600 34.800 201.000 35.200 ;
        RECT 184.600 32.800 185.000 33.200 ;
        RECT 194.200 33.100 194.600 33.500 ;
        RECT 205.400 38.800 205.800 39.200 ;
        RECT 204.600 33.800 205.000 34.200 ;
        RECT 212.600 36.200 213.000 36.600 ;
        RECT 214.200 35.500 214.600 35.900 ;
        RECT 215.800 34.800 216.200 35.200 ;
        RECT 185.400 31.800 185.800 32.200 ;
        RECT 202.200 31.800 202.600 32.200 ;
        RECT 218.200 33.800 218.600 34.200 ;
        RECT 214.200 33.100 214.600 33.500 ;
        RECT 219.800 33.800 220.200 34.200 ;
        RECT 227.800 36.200 228.200 36.600 ;
        RECT 229.400 35.500 229.800 35.900 ;
        RECT 224.600 34.800 225.000 35.200 ;
        RECT 229.400 33.100 229.800 33.500 ;
        RECT 3.800 28.800 4.200 29.200 ;
        RECT 13.400 28.800 13.800 29.200 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 6.200 26.100 6.600 26.500 ;
        RECT 2.200 24.800 2.600 25.200 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 23.800 28.800 24.200 29.200 ;
        RECT 21.400 26.800 21.800 27.200 ;
        RECT 15.800 26.100 16.200 26.500 ;
        RECT 12.600 25.100 13.000 25.500 ;
        RECT 22.200 25.100 22.600 25.500 ;
        RECT 27.000 28.800 27.400 29.200 ;
        RECT 39.000 28.800 39.400 29.200 ;
        RECT 26.200 24.800 26.600 25.200 ;
        RECT 68.600 28.800 69.000 29.200 ;
        RECT 47.000 26.800 47.400 27.200 ;
        RECT 50.200 26.800 50.600 27.200 ;
        RECT 41.400 26.100 41.800 26.500 ;
        RECT 45.400 25.900 45.800 26.300 ;
        RECT 47.800 25.100 48.200 25.500 ;
        RECT 60.600 26.800 61.000 27.200 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 55.800 24.800 56.200 25.200 ;
        RECT 59.800 25.100 60.200 25.500 ;
        RECT 69.400 28.800 69.800 29.200 ;
        RECT 86.200 28.800 86.600 29.200 ;
        RECT 71.800 26.100 72.200 26.500 ;
        RECT 75.800 25.900 76.200 26.300 ;
        RECT 78.200 25.100 78.600 25.500 ;
        RECT 80.600 24.800 81.000 25.200 ;
        RECT 84.600 25.800 85.000 26.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 97.400 28.800 97.800 29.200 ;
        RECT 99.800 28.800 100.200 29.200 ;
        RECT 115.000 28.800 115.400 29.200 ;
        RECT 88.600 26.100 89.000 26.500 ;
        RECT 95.000 25.100 95.400 25.500 ;
        RECT 97.400 24.800 97.800 25.200 ;
        RECT 107.000 26.800 107.400 27.200 ;
        RECT 104.600 25.800 105.000 26.200 ;
        RECT 108.600 25.900 109.000 26.300 ;
        RECT 105.400 24.800 105.800 25.200 ;
        RECT 106.200 25.100 106.600 25.500 ;
        RECT 115.800 28.800 116.200 29.200 ;
        RECT 122.200 26.800 122.600 27.200 ;
        RECT 118.200 26.100 118.600 26.500 ;
        RECT 124.600 25.100 125.000 25.500 ;
        RECT 125.400 24.800 125.800 25.200 ;
        RECT 149.400 28.800 149.800 29.200 ;
        RECT 134.200 26.800 134.600 27.200 ;
        RECT 140.600 21.800 141.000 22.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 160.600 26.800 161.000 27.200 ;
        RECT 164.600 26.800 165.000 27.200 ;
        RECT 151.800 26.100 152.200 26.500 ;
        RECT 153.400 25.800 153.800 26.200 ;
        RECT 145.400 24.800 145.800 25.200 ;
        RECT 147.800 24.800 148.200 25.200 ;
        RECT 158.200 25.100 158.600 25.500 ;
        RECT 161.400 24.800 161.800 25.200 ;
        RECT 165.400 24.800 165.800 25.200 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 170.200 26.100 170.600 26.500 ;
        RECT 199.000 28.800 199.400 29.200 ;
        RECT 179.800 26.100 180.200 26.500 ;
        RECT 191.000 25.900 191.400 26.300 ;
        RECT 176.600 25.100 177.000 25.500 ;
        RECT 186.200 25.100 186.600 25.500 ;
        RECT 188.600 25.100 189.000 25.500 ;
        RECT 198.200 24.800 198.600 25.200 ;
        RECT 197.400 23.800 197.800 24.200 ;
        RECT 202.200 28.800 202.600 29.200 ;
        RECT 209.400 28.800 209.800 29.200 ;
        RECT 207.000 26.800 207.400 27.200 ;
        RECT 221.400 28.800 221.800 29.200 ;
        RECT 207.000 24.800 207.400 25.200 ;
        RECT 213.400 26.800 213.800 27.200 ;
        RECT 215.800 26.800 216.200 27.200 ;
        RECT 211.800 26.100 212.200 26.500 ;
        RECT 218.200 25.100 218.600 25.500 ;
        RECT 219.000 24.800 219.400 25.200 ;
        RECT 223.800 26.100 224.200 26.500 ;
        RECT 230.200 25.100 230.600 25.500 ;
        RECT 9.400 18.800 9.800 19.200 ;
        RECT 0.600 13.100 1.000 13.500 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 12.600 13.800 13.000 14.200 ;
        RECT 13.400 13.100 13.800 13.500 ;
        RECT 23.800 18.800 24.200 19.200 ;
        RECT 28.600 14.800 29.000 15.200 ;
        RECT 24.600 13.100 25.000 13.500 ;
        RECT 37.400 14.800 37.800 15.200 ;
        RECT 36.600 13.800 37.000 14.200 ;
        RECT 42.200 14.800 42.600 15.200 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 55.800 18.800 56.200 19.200 ;
        RECT 51.800 14.800 52.200 15.200 ;
        RECT 47.800 13.800 48.200 14.200 ;
        RECT 33.400 11.800 33.800 12.200 ;
        RECT 47.000 13.100 47.400 13.500 ;
        RECT 57.400 14.800 57.800 15.200 ;
        RECT 63.000 18.800 63.400 19.200 ;
        RECT 59.000 11.800 59.400 12.200 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 78.200 18.800 78.600 19.200 ;
        RECT 67.000 13.800 67.400 14.200 ;
        RECT 68.600 13.800 69.000 14.200 ;
        RECT 69.400 13.100 69.800 13.500 ;
        RECT 76.600 13.800 77.000 14.200 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 71.800 12.800 72.200 13.200 ;
        RECT 81.400 18.800 81.800 19.200 ;
        RECT 80.600 13.800 81.000 14.200 ;
        RECT 79.800 11.800 80.200 12.200 ;
        RECT 83.000 14.800 83.400 15.200 ;
        RECT 98.200 16.800 98.600 17.200 ;
        RECT 85.400 13.800 85.800 14.200 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 88.600 13.800 89.000 14.200 ;
        RECT 81.400 11.800 81.800 12.200 ;
        RECT 89.400 13.100 89.800 13.500 ;
        RECT 99.800 18.800 100.200 19.200 ;
        RECT 99.000 12.800 99.400 13.200 ;
        RECT 109.400 18.800 109.800 19.200 ;
        RECT 103.800 14.800 104.200 15.200 ;
        RECT 100.600 13.100 101.000 13.500 ;
        RECT 118.200 18.800 118.600 19.200 ;
        RECT 115.800 14.800 116.200 15.200 ;
        RECT 116.600 14.800 117.000 15.200 ;
        RECT 115.000 13.800 115.400 14.200 ;
        RECT 121.400 14.800 121.800 15.200 ;
        RECT 127.800 18.800 128.200 19.200 ;
        RECT 125.400 13.800 125.800 14.200 ;
        RECT 123.000 11.800 123.400 12.200 ;
        RECT 129.400 13.800 129.800 14.200 ;
        RECT 134.200 18.800 134.600 19.200 ;
        RECT 135.000 14.800 135.400 15.200 ;
        RECT 135.800 14.800 136.200 15.200 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 127.800 11.800 128.200 12.200 ;
        RECT 142.200 14.800 142.600 15.200 ;
        RECT 157.400 18.800 157.800 19.200 ;
        RECT 143.000 13.800 143.400 14.200 ;
        RECT 147.000 14.800 147.400 15.200 ;
        RECT 147.800 14.800 148.200 15.200 ;
        RECT 152.600 14.800 153.000 15.200 ;
        RECT 167.800 16.800 168.200 17.200 ;
        RECT 149.400 13.800 149.800 14.200 ;
        RECT 140.600 11.800 141.000 12.200 ;
        RECT 148.600 13.100 149.000 13.500 ;
        RECT 161.400 14.800 161.800 15.200 ;
        RECT 158.200 13.100 158.600 13.500 ;
        RECT 180.600 16.800 181.000 17.200 ;
        RECT 167.800 13.800 168.200 14.200 ;
        RECT 172.600 14.800 173.000 15.200 ;
        RECT 176.600 14.800 177.000 15.200 ;
        RECT 172.600 13.800 173.000 14.200 ;
        RECT 174.200 13.800 174.600 14.200 ;
        RECT 173.400 13.100 173.800 13.500 ;
        RECT 182.200 11.800 182.600 12.200 ;
        RECT 187.000 18.800 187.400 19.200 ;
        RECT 185.400 12.800 185.800 13.200 ;
        RECT 183.800 11.800 184.200 12.200 ;
        RECT 199.000 16.200 199.400 16.600 ;
        RECT 200.600 15.500 201.000 15.900 ;
        RECT 203.800 18.800 204.200 19.200 ;
        RECT 201.400 14.800 201.800 15.200 ;
        RECT 202.200 14.800 202.600 15.200 ;
        RECT 188.600 11.800 189.000 12.200 ;
        RECT 206.200 13.800 206.600 14.200 ;
        RECT 198.200 12.800 198.600 13.200 ;
        RECT 200.600 13.100 201.000 13.500 ;
        RECT 210.200 14.800 210.600 15.200 ;
        RECT 212.600 14.800 213.000 15.200 ;
        RECT 211.000 13.800 211.400 14.200 ;
        RECT 216.600 13.800 217.000 14.200 ;
        RECT 228.600 18.800 229.000 19.200 ;
        RECT 224.600 13.800 225.000 14.200 ;
        RECT 208.600 11.800 209.000 12.200 ;
        RECT 214.200 11.800 214.600 12.200 ;
        RECT 228.600 14.800 229.000 15.200 ;
        RECT 229.400 13.800 229.800 14.200 ;
        RECT 223.000 11.800 223.400 12.200 ;
        RECT 0.600 8.800 1.000 9.200 ;
        RECT 3.800 6.800 4.200 7.200 ;
        RECT 11.800 8.800 12.200 9.200 ;
        RECT 14.200 8.800 14.600 9.200 ;
        RECT 5.400 5.800 5.800 6.200 ;
        RECT 3.800 4.800 4.200 5.200 ;
        RECT 13.400 4.800 13.800 5.200 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 21.400 8.800 21.800 9.200 ;
        RECT 39.000 8.800 39.400 9.200 ;
        RECT 29.400 6.800 29.800 7.200 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 35.800 6.800 36.200 7.200 ;
        RECT 35.000 5.800 35.400 6.200 ;
        RECT 30.200 5.100 30.600 5.500 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 45.400 4.800 45.800 5.200 ;
        RECT 67.800 8.800 68.200 9.200 ;
        RECT 77.400 8.800 77.800 9.200 ;
        RECT 51.800 6.100 52.200 6.500 ;
        RECT 55.800 5.900 56.200 6.300 ;
        RECT 58.200 5.100 58.600 5.500 ;
        RECT 59.000 5.100 59.400 5.500 ;
        RECT 69.400 6.800 69.800 7.200 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 72.600 5.800 73.000 6.200 ;
        RECT 68.600 5.100 69.000 5.500 ;
        RECT 79.800 6.800 80.200 7.200 ;
        RECT 82.200 6.800 82.600 7.200 ;
        RECT 93.400 6.800 93.800 7.200 ;
        RECT 78.200 4.800 78.600 5.200 ;
        RECT 105.400 8.800 105.800 9.200 ;
        RECT 100.600 6.800 101.000 7.200 ;
        RECT 99.000 5.900 99.400 6.300 ;
        RECT 94.200 4.800 94.600 5.200 ;
        RECT 96.600 5.100 97.000 5.500 ;
        RECT 108.600 8.800 109.000 9.200 ;
        RECT 119.000 8.800 119.400 9.200 ;
        RECT 128.600 8.800 129.000 9.200 ;
        RECT 114.200 6.800 114.600 7.200 ;
        RECT 114.200 5.800 114.600 6.200 ;
        RECT 110.200 5.100 110.600 5.500 ;
        RECT 132.600 8.800 133.000 9.200 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 119.800 5.100 120.200 5.500 ;
        RECT 137.400 6.800 137.800 7.200 ;
        RECT 143.800 8.800 144.200 9.200 ;
        RECT 135.000 6.100 135.400 6.500 ;
        RECT 139.000 5.900 139.400 6.300 ;
        RECT 149.400 6.800 149.800 7.200 ;
        RECT 164.600 8.800 165.000 9.200 ;
        RECT 146.200 6.100 146.600 6.500 ;
        RECT 141.400 5.100 141.800 5.500 ;
        RECT 150.200 5.900 150.600 6.300 ;
        RECT 159.000 6.800 159.400 7.200 ;
        RECT 161.400 6.800 161.800 7.200 ;
        RECT 152.600 5.100 153.000 5.500 ;
        RECT 155.000 4.800 155.400 5.200 ;
        RECT 162.200 4.800 162.600 5.200 ;
        RECT 167.000 6.100 167.400 6.500 ;
        RECT 173.400 5.100 173.800 5.500 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 182.200 6.800 182.600 7.200 ;
        RECT 187.800 6.800 188.200 7.200 ;
        RECT 195.800 8.800 196.200 9.200 ;
        RECT 189.400 4.800 189.800 5.200 ;
        RECT 208.600 8.800 209.000 9.200 ;
        RECT 202.200 5.900 202.600 6.300 ;
        RECT 199.800 5.100 200.200 5.500 ;
        RECT 209.400 8.800 209.800 9.200 ;
        RECT 219.800 8.800 220.200 9.200 ;
        RECT 221.400 8.800 221.800 9.200 ;
        RECT 217.400 6.800 217.800 7.200 ;
        RECT 211.800 6.100 212.200 6.500 ;
        RECT 218.200 5.100 218.600 5.500 ;
        RECT 219.000 4.800 219.400 5.200 ;
        RECT 223.800 6.100 224.200 6.500 ;
        RECT 230.200 5.100 230.600 5.500 ;
      LAYER metal2 ;
        RECT 14.200 206.800 14.600 207.200 ;
        RECT 14.200 206.200 14.500 206.800 ;
        RECT 14.200 205.800 14.600 206.200 ;
        RECT 15.000 205.100 15.400 207.900 ;
        RECT 15.800 206.800 16.200 207.200 ;
        RECT 15.800 206.200 16.100 206.800 ;
        RECT 15.800 205.800 16.200 206.200 ;
        RECT 16.600 203.100 17.000 208.900 ;
        RECT 18.200 205.800 18.600 206.200 ;
        RECT 6.200 201.800 6.600 202.200 ;
        RECT 0.600 198.100 1.000 198.200 ;
        RECT 1.400 198.100 1.800 198.200 ;
        RECT 0.600 197.800 1.800 198.100 ;
        RECT 3.000 192.100 3.400 197.900 ;
        RECT 6.200 194.200 6.500 201.800 ;
        RECT 18.200 199.200 18.500 205.800 ;
        RECT 21.400 203.100 21.800 208.900 ;
        RECT 24.600 208.800 25.000 209.200 ;
        RECT 24.600 207.200 24.900 208.800 ;
        RECT 24.600 206.800 25.000 207.200 ;
        RECT 30.200 206.800 30.600 207.200 ;
        RECT 23.000 203.800 23.400 204.200 ;
        RECT 19.800 201.800 20.200 202.200 ;
        RECT 18.200 198.800 18.600 199.200 ;
        RECT 7.000 195.800 7.400 196.200 ;
        RECT 7.000 195.100 7.300 195.800 ;
        RECT 7.000 194.700 7.400 195.100 ;
        RECT 6.200 193.800 6.600 194.200 ;
        RECT 6.200 193.200 6.500 193.800 ;
        RECT 6.200 192.800 6.600 193.200 ;
        RECT 7.800 192.100 8.200 197.900 ;
        RECT 13.400 197.800 13.800 198.200 ;
        RECT 13.400 197.200 13.700 197.800 ;
        RECT 19.800 197.200 20.100 201.800 ;
        RECT 10.200 196.800 10.600 197.200 ;
        RECT 13.400 196.800 13.800 197.200 ;
        RECT 15.000 197.100 15.400 197.200 ;
        RECT 15.800 197.100 16.200 197.200 ;
        RECT 15.000 196.800 16.200 197.100 ;
        RECT 16.600 196.800 17.000 197.200 ;
        RECT 19.800 196.800 20.200 197.200 ;
        RECT 21.400 197.100 21.800 197.200 ;
        RECT 22.200 197.100 22.600 197.200 ;
        RECT 21.400 196.800 22.600 197.100 ;
        RECT 10.200 196.200 10.500 196.800 ;
        RECT 9.400 193.100 9.800 195.900 ;
        RECT 10.200 195.800 10.600 196.200 ;
        RECT 12.600 195.800 13.000 196.200 ;
        RECT 10.200 195.100 10.600 195.200 ;
        RECT 11.000 195.100 11.400 195.200 ;
        RECT 10.200 194.800 11.400 195.100 ;
        RECT 11.800 194.800 12.200 195.200 ;
        RECT 11.800 192.200 12.100 194.800 ;
        RECT 12.600 194.200 12.900 195.800 ;
        RECT 12.600 193.800 13.000 194.200 ;
        RECT 11.800 191.800 12.200 192.200 ;
        RECT 0.600 185.100 1.000 187.900 ;
        RECT 2.200 183.100 2.600 188.900 ;
        RECT 4.600 186.100 5.000 186.200 ;
        RECT 5.400 186.100 5.800 186.200 ;
        RECT 4.600 185.800 5.800 186.100 ;
        RECT 6.200 185.800 6.600 186.200 ;
        RECT 6.200 179.200 6.500 185.800 ;
        RECT 7.000 183.100 7.400 188.900 ;
        RECT 12.600 187.200 12.900 193.800 ;
        RECT 13.400 187.200 13.700 196.800 ;
        RECT 16.600 196.200 16.900 196.800 ;
        RECT 16.600 195.800 17.000 196.200 ;
        RECT 23.000 195.200 23.300 203.800 ;
        RECT 23.800 201.800 24.200 202.200 ;
        RECT 23.800 201.200 24.100 201.800 ;
        RECT 23.800 200.800 24.200 201.200 ;
        RECT 15.000 195.100 15.400 195.200 ;
        RECT 15.800 195.100 16.200 195.200 ;
        RECT 15.000 194.800 16.200 195.100 ;
        RECT 18.200 194.800 18.600 195.200 ;
        RECT 23.000 194.800 23.400 195.200 ;
        RECT 10.200 186.800 10.600 187.200 ;
        RECT 12.600 186.800 13.000 187.200 ;
        RECT 13.400 186.800 13.800 187.200 ;
        RECT 10.200 186.200 10.500 186.800 ;
        RECT 15.000 186.200 15.300 194.800 ;
        RECT 15.800 194.100 16.200 194.200 ;
        RECT 16.600 194.100 17.000 194.200 ;
        RECT 15.800 193.800 17.000 194.100 ;
        RECT 15.800 187.200 16.100 193.800 ;
        RECT 18.200 192.200 18.500 194.800 ;
        RECT 19.000 193.800 19.400 194.200 ;
        RECT 23.000 193.800 23.400 194.200 ;
        RECT 18.200 191.800 18.600 192.200 ;
        RECT 19.000 191.200 19.300 193.800 ;
        RECT 19.000 190.800 19.400 191.200 ;
        RECT 23.000 190.200 23.300 193.800 ;
        RECT 23.000 189.800 23.400 190.200 ;
        RECT 15.800 186.800 16.200 187.200 ;
        RECT 10.200 185.800 10.600 186.200 ;
        RECT 11.000 186.100 11.400 186.200 ;
        RECT 11.800 186.100 12.200 186.200 ;
        RECT 11.000 185.800 12.200 186.100 ;
        RECT 12.600 185.800 13.000 186.200 ;
        RECT 15.000 185.800 15.400 186.200 ;
        RECT 12.600 185.200 12.900 185.800 ;
        RECT 10.200 185.100 10.600 185.200 ;
        RECT 11.000 185.100 11.400 185.200 ;
        RECT 10.200 184.800 11.400 185.100 ;
        RECT 12.600 184.800 13.000 185.200 ;
        RECT 13.400 184.800 13.800 185.200 ;
        RECT 16.600 185.100 17.000 187.900 ;
        RECT 13.400 184.200 13.700 184.800 ;
        RECT 9.400 184.100 9.800 184.200 ;
        RECT 10.200 184.100 10.600 184.200 ;
        RECT 9.400 183.800 10.600 184.100 ;
        RECT 13.400 183.800 13.800 184.200 ;
        RECT 6.200 178.800 6.600 179.200 ;
        RECT 13.400 178.200 13.700 183.800 ;
        RECT 18.200 183.100 18.600 188.900 ;
        RECT 19.800 187.800 20.200 188.200 ;
        RECT 19.800 186.200 20.100 187.800 ;
        RECT 19.800 185.800 20.200 186.200 ;
        RECT 22.200 185.800 22.600 186.200 ;
        RECT 6.200 174.800 6.600 175.200 ;
        RECT 6.200 172.200 6.500 174.800 ;
        RECT 6.200 171.800 6.600 172.200 ;
        RECT 7.800 171.800 8.200 172.200 ;
        RECT 10.200 172.100 10.600 177.900 ;
        RECT 13.400 177.800 13.800 178.200 ;
        RECT 11.000 174.800 11.400 175.200 ;
        RECT 11.000 174.200 11.300 174.800 ;
        RECT 14.200 174.700 14.600 175.100 ;
        RECT 11.000 173.800 11.400 174.200 ;
        RECT 0.600 165.100 1.000 167.900 ;
        RECT 2.200 163.100 2.600 168.900 ;
        RECT 3.000 165.900 3.400 166.300 ;
        RECT 6.200 166.200 6.500 171.800 ;
        RECT 3.000 162.100 3.300 165.900 ;
        RECT 6.200 165.800 6.600 166.200 ;
        RECT 7.000 163.100 7.400 168.900 ;
        RECT 7.800 167.200 8.100 171.800 ;
        RECT 14.200 169.200 14.500 174.700 ;
        RECT 15.000 172.100 15.400 177.900 ;
        RECT 16.600 173.100 17.000 175.900 ;
        RECT 22.200 174.200 22.500 185.800 ;
        RECT 23.000 183.100 23.400 188.900 ;
        RECT 23.800 186.200 24.100 200.800 ;
        RECT 24.600 194.200 24.900 206.800 ;
        RECT 30.200 206.200 30.500 206.800 ;
        RECT 25.400 205.800 25.800 206.200 ;
        RECT 27.800 206.100 28.200 206.200 ;
        RECT 28.600 206.100 29.000 206.200 ;
        RECT 27.800 205.800 29.000 206.100 ;
        RECT 29.400 205.800 29.800 206.200 ;
        RECT 30.200 205.800 30.600 206.200 ;
        RECT 25.400 204.200 25.700 205.800 ;
        RECT 29.400 205.200 29.700 205.800 ;
        RECT 29.400 204.800 29.800 205.200 ;
        RECT 31.000 205.100 31.400 207.900 ;
        RECT 31.800 207.800 32.200 208.200 ;
        RECT 31.800 207.200 32.100 207.800 ;
        RECT 31.800 206.800 32.200 207.200 ;
        RECT 25.400 203.800 25.800 204.200 ;
        RECT 27.000 203.800 27.400 204.200 ;
        RECT 27.000 203.200 27.300 203.800 ;
        RECT 27.000 202.800 27.400 203.200 ;
        RECT 32.600 203.100 33.000 208.900 ;
        RECT 35.000 206.800 35.400 207.200 ;
        RECT 33.400 205.900 33.800 206.300 ;
        RECT 33.400 205.200 33.700 205.900 ;
        RECT 33.400 204.800 33.800 205.200 ;
        RECT 33.400 203.800 33.800 204.200 ;
        RECT 25.400 197.100 25.800 197.200 ;
        RECT 26.200 197.100 26.600 197.200 ;
        RECT 25.400 196.800 26.600 197.100 ;
        RECT 27.800 195.100 28.200 195.200 ;
        RECT 28.600 195.100 29.000 195.200 ;
        RECT 27.800 194.800 29.000 195.100 ;
        RECT 24.600 193.800 25.000 194.200 ;
        RECT 26.200 194.100 26.600 194.200 ;
        RECT 27.000 194.100 27.400 194.200 ;
        RECT 26.200 193.800 27.400 194.100 ;
        RECT 28.600 193.800 29.000 194.200 ;
        RECT 27.000 191.800 27.400 192.200 ;
        RECT 26.200 190.800 26.600 191.200 ;
        RECT 26.200 187.200 26.500 190.800 ;
        RECT 26.200 186.800 26.600 187.200 ;
        RECT 27.000 186.200 27.300 191.800 ;
        RECT 28.600 191.200 28.900 193.800 ;
        RECT 29.400 193.100 29.800 195.900 ;
        RECT 31.000 192.100 31.400 197.900 ;
        RECT 31.800 194.700 32.200 195.100 ;
        RECT 31.800 194.200 32.100 194.700 ;
        RECT 31.800 193.800 32.200 194.200 ;
        RECT 28.600 190.800 29.000 191.200 ;
        RECT 32.600 189.800 33.000 190.200 ;
        RECT 27.800 187.800 28.200 188.200 ;
        RECT 27.800 187.200 28.100 187.800 ;
        RECT 32.600 187.200 32.900 189.800 ;
        RECT 27.800 186.800 28.200 187.200 ;
        RECT 32.600 186.800 33.000 187.200 ;
        RECT 33.400 186.200 33.700 203.800 ;
        RECT 35.000 195.200 35.300 206.800 ;
        RECT 37.400 203.100 37.800 208.900 ;
        RECT 44.600 205.800 45.000 206.200 ;
        RECT 44.600 205.200 44.900 205.800 ;
        RECT 43.000 204.800 43.400 205.200 ;
        RECT 44.600 204.800 45.000 205.200 ;
        RECT 45.400 205.100 45.800 207.900 ;
        RECT 46.200 207.800 46.600 208.200 ;
        RECT 46.200 207.200 46.500 207.800 ;
        RECT 46.200 206.800 46.600 207.200 ;
        RECT 43.000 204.200 43.300 204.800 ;
        RECT 43.000 203.800 43.400 204.200 ;
        RECT 39.000 203.100 39.400 203.200 ;
        RECT 39.800 203.100 40.200 203.200 ;
        RECT 39.000 202.800 40.200 203.100 ;
        RECT 35.000 194.800 35.400 195.200 ;
        RECT 35.800 192.100 36.200 197.900 ;
        RECT 37.400 197.100 37.800 197.200 ;
        RECT 38.200 197.100 38.600 197.200 ;
        RECT 37.400 196.800 38.600 197.100 ;
        RECT 40.600 193.100 41.000 195.900 ;
        RECT 41.400 193.800 41.800 194.200 ;
        RECT 41.400 193.200 41.700 193.800 ;
        RECT 41.400 192.800 41.800 193.200 ;
        RECT 42.200 192.100 42.600 197.900 ;
        RECT 45.400 194.800 45.800 195.200 ;
        RECT 45.400 194.200 45.700 194.800 ;
        RECT 45.400 193.800 45.800 194.200 ;
        RECT 46.200 192.200 46.500 206.800 ;
        RECT 47.000 203.100 47.400 208.900 ;
        RECT 48.600 206.800 49.000 207.200 ;
        RECT 48.600 206.200 48.900 206.800 ;
        RECT 48.600 205.800 49.000 206.200 ;
        RECT 51.800 203.100 52.200 208.900 ;
        RECT 60.600 208.800 61.000 209.200 ;
        RECT 60.600 207.200 60.900 208.800 ;
        RECT 55.000 206.800 55.400 207.200 ;
        RECT 56.600 207.100 57.000 207.200 ;
        RECT 57.400 207.100 57.800 207.200 ;
        RECT 56.600 206.800 57.800 207.100 ;
        RECT 60.600 206.800 61.000 207.200 ;
        RECT 55.000 205.200 55.300 206.800 ;
        RECT 55.800 205.800 56.200 206.200 ;
        RECT 63.800 205.800 64.200 206.200 ;
        RECT 55.000 204.800 55.400 205.200 ;
        RECT 54.200 204.100 54.600 204.200 ;
        RECT 55.000 204.100 55.400 204.200 ;
        RECT 54.200 203.800 55.400 204.100 ;
        RECT 47.800 201.800 48.200 202.200 ;
        RECT 46.200 191.800 46.600 192.200 ;
        RECT 47.000 192.100 47.400 197.900 ;
        RECT 47.800 197.200 48.100 201.800 ;
        RECT 47.800 196.800 48.200 197.200 ;
        RECT 49.400 196.100 49.800 196.200 ;
        RECT 50.200 196.100 50.600 196.200 ;
        RECT 49.400 195.800 50.600 196.100 ;
        RECT 54.200 195.200 54.500 203.800 ;
        RECT 55.800 195.200 56.100 205.800 ;
        RECT 58.200 204.800 58.600 205.200 ;
        RECT 58.200 204.200 58.500 204.800 ;
        RECT 58.200 203.800 58.600 204.200 ;
        RECT 62.200 201.800 62.600 202.200 ;
        RECT 56.600 196.800 57.000 197.200 ;
        RECT 56.600 195.200 56.900 196.800 ;
        RECT 59.800 196.100 60.200 196.200 ;
        RECT 60.600 196.100 61.000 196.200 ;
        RECT 59.800 195.800 61.000 196.100 ;
        RECT 51.000 195.100 51.400 195.200 ;
        RECT 51.800 195.100 52.200 195.200 ;
        RECT 51.000 194.800 52.200 195.100 ;
        RECT 54.200 194.800 54.600 195.200 ;
        RECT 55.800 194.800 56.200 195.200 ;
        RECT 56.600 194.800 57.000 195.200 ;
        RECT 57.400 195.100 57.800 195.200 ;
        RECT 58.200 195.100 58.600 195.200 ;
        RECT 57.400 194.800 58.600 195.100 ;
        RECT 59.000 194.800 59.400 195.200 ;
        RECT 59.000 194.200 59.300 194.800 ;
        RECT 50.200 194.100 50.600 194.200 ;
        RECT 51.000 194.100 51.400 194.200 ;
        RECT 52.600 194.100 53.000 194.200 ;
        RECT 50.200 193.800 51.400 194.100 ;
        RECT 51.800 193.800 53.000 194.100 ;
        RECT 57.400 194.100 57.800 194.200 ;
        RECT 58.200 194.100 58.600 194.200 ;
        RECT 57.400 193.800 58.600 194.100 ;
        RECT 59.000 193.800 59.400 194.200 ;
        RECT 59.800 194.100 60.200 194.200 ;
        RECT 60.600 194.100 61.000 194.200 ;
        RECT 59.800 193.800 61.000 194.100 ;
        RECT 49.400 191.800 49.800 192.200 ;
        RECT 36.600 190.800 37.000 191.200 ;
        RECT 23.800 185.800 24.200 186.200 ;
        RECT 27.000 185.800 27.400 186.200 ;
        RECT 33.400 185.800 33.800 186.200 ;
        RECT 25.400 184.100 25.800 184.200 ;
        RECT 26.200 184.100 26.600 184.200 ;
        RECT 25.400 183.800 26.600 184.100 ;
        RECT 22.200 173.800 22.600 174.200 ;
        RECT 19.800 172.800 20.200 173.200 ;
        RECT 24.600 173.100 25.000 175.900 ;
        RECT 25.400 174.800 25.800 175.200 ;
        RECT 25.400 174.200 25.700 174.800 ;
        RECT 25.400 173.800 25.800 174.200 ;
        RECT 14.200 168.800 14.600 169.200 ;
        RECT 10.200 167.800 10.600 168.200 ;
        RECT 10.200 167.200 10.500 167.800 ;
        RECT 19.800 167.200 20.100 172.800 ;
        RECT 23.000 171.800 23.400 172.200 ;
        RECT 7.800 166.800 8.200 167.200 ;
        RECT 10.200 166.800 10.600 167.200 ;
        RECT 11.000 167.100 11.400 167.200 ;
        RECT 11.800 167.100 12.200 167.200 ;
        RECT 11.000 166.800 12.200 167.100 ;
        RECT 16.600 167.100 17.000 167.200 ;
        RECT 17.400 167.100 17.800 167.200 ;
        RECT 16.600 166.800 17.800 167.100 ;
        RECT 19.000 167.100 19.400 167.200 ;
        RECT 19.800 167.100 20.200 167.200 ;
        RECT 19.000 166.800 20.200 167.100 ;
        RECT 15.800 165.800 16.200 166.200 ;
        RECT 17.400 166.100 17.800 166.200 ;
        RECT 18.200 166.100 18.600 166.200 ;
        RECT 17.400 165.800 18.600 166.100 ;
        RECT 15.800 165.200 16.100 165.800 ;
        RECT 12.600 165.100 13.000 165.200 ;
        RECT 13.400 165.100 13.800 165.200 ;
        RECT 12.600 164.800 13.800 165.100 ;
        RECT 15.800 164.800 16.200 165.200 ;
        RECT 2.200 161.800 3.300 162.100 ;
        RECT 5.400 161.800 5.800 162.200 ;
        RECT 8.600 162.100 9.000 162.200 ;
        RECT 9.400 162.100 9.800 162.200 ;
        RECT 8.600 161.800 9.800 162.100 ;
        RECT 11.000 161.800 11.400 162.200 ;
        RECT 2.200 159.200 2.500 161.800 ;
        RECT 2.200 158.800 2.600 159.200 ;
        RECT 1.400 156.800 1.800 157.200 ;
        RECT 0.600 155.800 1.000 156.200 ;
        RECT 0.600 153.200 0.900 155.800 ;
        RECT 0.600 152.800 1.000 153.200 ;
        RECT 0.600 145.100 1.000 147.900 ;
        RECT 0.600 133.100 1.000 135.900 ;
        RECT 0.600 124.800 1.000 125.200 ;
        RECT 0.600 118.100 0.900 124.800 ;
        RECT 1.400 119.200 1.700 156.800 ;
        RECT 3.800 155.800 4.200 156.200 ;
        RECT 3.800 155.200 4.100 155.800 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 5.400 154.200 5.700 161.800 ;
        RECT 6.200 156.800 6.600 157.200 ;
        RECT 6.200 155.200 6.500 156.800 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 10.200 154.200 10.500 154.800 ;
        RECT 3.000 154.100 3.400 154.200 ;
        RECT 3.800 154.100 4.200 154.200 ;
        RECT 3.000 153.800 4.200 154.100 ;
        RECT 5.400 153.800 5.800 154.200 ;
        RECT 7.800 154.100 8.200 154.200 ;
        RECT 8.600 154.100 9.000 154.200 ;
        RECT 7.800 153.800 9.000 154.100 ;
        RECT 9.400 153.800 9.800 154.200 ;
        RECT 10.200 153.800 10.600 154.200 ;
        RECT 3.800 153.100 4.200 153.200 ;
        RECT 4.600 153.100 5.000 153.200 ;
        RECT 3.800 152.800 5.000 153.100 ;
        RECT 5.400 150.200 5.700 153.800 ;
        RECT 5.400 149.800 5.800 150.200 ;
        RECT 2.200 143.100 2.600 148.900 ;
        RECT 3.800 146.800 4.200 147.200 ;
        RECT 4.600 146.800 5.000 147.200 ;
        RECT 3.800 146.200 4.100 146.800 ;
        RECT 3.800 145.800 4.200 146.200 ;
        RECT 2.200 132.100 2.600 137.900 ;
        RECT 3.800 134.800 4.200 135.200 ;
        RECT 3.800 134.200 4.100 134.800 ;
        RECT 4.600 134.200 4.900 146.800 ;
        RECT 7.000 143.100 7.400 148.900 ;
        RECT 8.600 148.200 8.900 153.800 ;
        RECT 9.400 152.200 9.700 153.800 ;
        RECT 9.400 151.800 9.800 152.200 ;
        RECT 9.400 149.100 9.800 149.200 ;
        RECT 10.200 149.100 10.600 149.200 ;
        RECT 9.400 148.800 10.600 149.100 ;
        RECT 8.600 147.800 9.000 148.200 ;
        RECT 10.200 147.800 10.600 148.200 ;
        RECT 3.800 133.800 4.200 134.200 ;
        RECT 4.600 133.800 5.000 134.200 ;
        RECT 3.000 129.800 3.400 130.200 ;
        RECT 3.000 127.200 3.300 129.800 ;
        RECT 4.600 128.200 4.900 133.800 ;
        RECT 7.000 132.100 7.400 137.900 ;
        RECT 4.600 127.800 5.000 128.200 ;
        RECT 3.000 126.800 3.400 127.200 ;
        RECT 2.200 126.100 2.600 126.200 ;
        RECT 3.000 126.100 3.400 126.200 ;
        RECT 2.200 125.800 3.400 126.100 ;
        RECT 2.200 124.800 2.600 125.200 ;
        RECT 2.200 124.200 2.500 124.800 ;
        RECT 2.200 123.800 2.600 124.200 ;
        RECT 1.400 118.800 1.800 119.200 ;
        RECT 0.600 117.800 1.700 118.100 ;
        RECT 1.400 109.200 1.700 117.800 ;
        RECT 3.000 109.200 3.300 125.800 ;
        RECT 6.200 123.100 6.600 128.900 ;
        RECT 3.800 121.800 4.200 122.200 ;
        RECT 0.600 108.800 1.000 109.200 ;
        RECT 1.400 108.800 1.800 109.200 ;
        RECT 3.000 108.800 3.400 109.200 ;
        RECT 0.600 105.200 0.900 108.800 ;
        RECT 1.400 107.800 1.800 108.200 ;
        RECT 2.200 108.100 2.600 108.200 ;
        RECT 3.000 108.100 3.400 108.200 ;
        RECT 2.200 107.800 3.400 108.100 ;
        RECT 0.600 104.800 1.000 105.200 ;
        RECT 0.600 104.200 0.900 104.800 ;
        RECT 0.600 103.800 1.000 104.200 ;
        RECT 0.600 99.100 1.000 99.200 ;
        RECT 1.400 99.100 1.700 107.800 ;
        RECT 3.800 107.200 4.100 121.800 ;
        RECT 4.600 113.100 5.000 115.900 ;
        RECT 6.200 112.100 6.600 117.900 ;
        RECT 7.800 115.800 8.200 116.200 ;
        RECT 7.800 115.200 8.100 115.800 ;
        RECT 7.800 114.800 8.200 115.200 ;
        RECT 8.600 108.200 8.900 147.800 ;
        RECT 10.200 147.200 10.500 147.800 ;
        RECT 11.000 147.200 11.300 161.800 ;
        RECT 11.800 155.800 12.200 156.200 ;
        RECT 11.800 155.200 12.100 155.800 ;
        RECT 11.800 154.800 12.200 155.200 ;
        RECT 11.800 153.800 12.200 154.200 ;
        RECT 11.800 153.200 12.100 153.800 ;
        RECT 11.800 152.800 12.200 153.200 ;
        RECT 12.600 153.100 13.000 155.900 ;
        RECT 14.200 152.100 14.600 157.900 ;
        RECT 17.400 157.200 17.700 165.800 ;
        RECT 20.600 165.100 21.000 167.900 ;
        RECT 22.200 163.100 22.600 168.900 ;
        RECT 23.000 162.200 23.300 171.800 ;
        RECT 23.800 167.800 24.200 168.200 ;
        RECT 23.800 166.200 24.100 167.800 ;
        RECT 25.400 166.200 25.700 173.800 ;
        RECT 26.200 172.100 26.600 177.900 ;
        RECT 27.000 173.200 27.300 185.800 ;
        RECT 29.400 184.800 29.800 185.200 ;
        RECT 29.400 184.200 29.700 184.800 ;
        RECT 29.400 183.800 29.800 184.200 ;
        RECT 35.000 183.800 35.400 184.200 ;
        RECT 33.400 181.800 33.800 182.200 ;
        RECT 33.400 180.200 33.700 181.800 ;
        RECT 33.400 179.800 33.800 180.200 ;
        RECT 35.000 179.200 35.300 183.800 ;
        RECT 35.800 182.800 36.200 183.200 ;
        RECT 33.400 179.100 33.800 179.200 ;
        RECT 34.200 179.100 34.600 179.200 ;
        RECT 33.400 178.800 34.600 179.100 ;
        RECT 35.000 178.800 35.400 179.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 29.400 175.100 29.800 175.200 ;
        RECT 28.600 174.800 29.800 175.100 ;
        RECT 27.000 172.800 27.400 173.200 ;
        RECT 31.000 172.100 31.400 177.900 ;
        RECT 35.800 177.200 36.100 182.800 ;
        RECT 35.800 176.800 36.200 177.200 ;
        RECT 33.400 176.100 33.800 176.200 ;
        RECT 34.200 176.100 34.600 176.200 ;
        RECT 33.400 175.800 34.600 176.100 ;
        RECT 35.800 175.200 36.100 176.800 ;
        RECT 34.200 175.100 34.600 175.200 ;
        RECT 35.000 175.100 35.400 175.200 ;
        RECT 34.200 174.800 35.400 175.100 ;
        RECT 35.800 174.800 36.200 175.200 ;
        RECT 36.600 174.200 36.900 190.800 ;
        RECT 38.200 186.800 38.600 187.200 ;
        RECT 38.200 186.200 38.500 186.800 ;
        RECT 38.200 185.800 38.600 186.200 ;
        RECT 39.800 186.100 40.200 186.200 ;
        RECT 40.600 186.100 41.000 186.200 ;
        RECT 39.800 185.800 41.000 186.100 ;
        RECT 41.400 185.800 41.800 186.200 ;
        RECT 41.400 182.200 41.700 185.800 ;
        RECT 42.200 185.100 42.600 187.900 ;
        RECT 43.800 183.100 44.200 188.900 ;
        RECT 46.200 187.200 46.500 191.800 ;
        RECT 46.200 186.800 46.600 187.200 ;
        RECT 39.800 181.800 40.200 182.200 ;
        RECT 41.400 181.800 41.800 182.200 ;
        RECT 43.000 181.800 43.400 182.200 ;
        RECT 39.800 179.100 40.100 181.800 ;
        RECT 39.800 178.800 40.900 179.100 ;
        RECT 39.800 177.800 40.200 178.200 ;
        RECT 39.800 175.200 40.100 177.800 ;
        RECT 39.800 174.800 40.200 175.200 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 40.600 169.200 40.900 178.800 ;
        RECT 42.200 178.800 42.600 179.200 ;
        RECT 42.200 175.200 42.500 178.800 ;
        RECT 43.000 175.200 43.300 181.800 ;
        RECT 42.200 174.800 42.600 175.200 ;
        RECT 43.000 174.800 43.400 175.200 ;
        RECT 43.800 173.100 44.200 175.900 ;
        RECT 41.400 171.800 41.800 172.200 ;
        RECT 45.400 172.100 45.800 177.900 ;
        RECT 46.200 174.200 46.500 186.800 ;
        RECT 47.000 186.100 47.400 186.200 ;
        RECT 47.800 186.100 48.200 186.200 ;
        RECT 47.000 185.800 48.200 186.100 ;
        RECT 48.600 183.100 49.000 188.900 ;
        RECT 49.400 185.200 49.700 191.800 ;
        RECT 51.800 187.200 52.100 193.800 ;
        RECT 58.200 192.800 58.600 193.200 ;
        RECT 61.400 193.100 61.800 195.900 ;
        RECT 62.200 195.200 62.500 201.800 ;
        RECT 62.200 194.800 62.600 195.200 ;
        RECT 62.200 193.800 62.600 194.200 ;
        RECT 55.800 191.800 56.200 192.200 ;
        RECT 51.800 186.800 52.200 187.200 ;
        RECT 49.400 184.800 49.800 185.200 ;
        RECT 51.000 181.800 51.400 182.200 ;
        RECT 51.000 180.200 51.300 181.800 ;
        RECT 51.800 181.200 52.100 186.800 ;
        RECT 55.800 186.200 56.100 191.800 ;
        RECT 58.200 189.200 58.500 192.800 ;
        RECT 62.200 192.200 62.500 193.800 ;
        RECT 62.200 191.800 62.600 192.200 ;
        RECT 63.000 192.100 63.400 197.900 ;
        RECT 63.800 197.200 64.100 205.800 ;
        RECT 64.600 205.100 65.000 207.900 ;
        RECT 65.400 202.800 65.800 203.200 ;
        RECT 66.200 203.100 66.600 208.900 ;
        RECT 67.000 206.800 67.400 207.200 ;
        RECT 63.800 196.800 64.200 197.200 ;
        RECT 63.800 194.700 64.200 195.100 ;
        RECT 63.800 194.200 64.100 194.700 ;
        RECT 63.800 193.800 64.200 194.200 ;
        RECT 58.200 188.800 58.600 189.200 ;
        RECT 57.400 187.100 57.800 187.200 ;
        RECT 58.200 187.100 58.600 187.200 ;
        RECT 57.400 186.800 58.600 187.100 ;
        RECT 60.600 187.100 61.000 187.200 ;
        RECT 61.400 187.100 61.800 187.200 ;
        RECT 60.600 186.800 61.800 187.100 ;
        RECT 52.600 185.800 53.000 186.200 ;
        RECT 53.400 186.100 53.800 186.200 ;
        RECT 54.200 186.100 54.600 186.200 ;
        RECT 53.400 185.800 54.600 186.100 ;
        RECT 55.800 185.800 56.200 186.200 ;
        RECT 56.600 185.800 57.000 186.200 ;
        RECT 52.600 183.200 52.900 185.800 ;
        RECT 55.000 184.800 55.400 185.200 ;
        RECT 52.600 182.800 53.000 183.200 ;
        RECT 51.800 180.800 52.200 181.200 ;
        RECT 55.000 180.200 55.300 184.800 ;
        RECT 56.600 183.200 56.900 185.800 ;
        RECT 56.600 182.800 57.000 183.200 ;
        RECT 51.000 179.800 51.400 180.200 ;
        RECT 55.000 179.800 55.400 180.200 ;
        RECT 47.800 175.100 48.200 175.200 ;
        RECT 48.600 175.100 49.000 175.200 ;
        RECT 47.800 174.800 49.000 175.100 ;
        RECT 46.200 173.800 46.600 174.200 ;
        RECT 23.800 165.800 24.200 166.200 ;
        RECT 25.400 165.800 25.800 166.200 ;
        RECT 23.000 161.800 23.400 162.200 ;
        RECT 25.400 158.200 25.700 165.800 ;
        RECT 27.000 163.100 27.400 168.900 ;
        RECT 32.600 168.800 33.000 169.200 ;
        RECT 32.600 168.200 32.900 168.800 ;
        RECT 32.600 167.800 33.000 168.200 ;
        RECT 27.800 166.800 28.200 167.200 ;
        RECT 30.200 166.800 30.600 167.200 ;
        RECT 35.000 166.800 35.400 167.200 ;
        RECT 18.200 157.800 18.600 158.200 ;
        RECT 17.400 156.800 17.800 157.200 ;
        RECT 17.400 155.800 17.800 156.200 ;
        RECT 15.000 154.700 15.400 155.100 ;
        RECT 15.000 154.200 15.300 154.700 ;
        RECT 15.000 153.800 15.400 154.200 ;
        RECT 16.600 153.800 17.000 154.200 ;
        RECT 17.400 154.100 17.700 155.800 ;
        RECT 18.200 155.200 18.500 157.800 ;
        RECT 18.200 154.800 18.600 155.200 ;
        RECT 17.400 153.800 18.500 154.100 ;
        RECT 15.000 148.800 15.400 149.200 ;
        RECT 15.000 147.200 15.300 148.800 ;
        RECT 10.200 146.800 10.600 147.200 ;
        RECT 11.000 146.800 11.400 147.200 ;
        RECT 15.000 146.800 15.400 147.200 ;
        RECT 11.000 145.800 11.400 146.200 ;
        RECT 11.800 146.100 12.200 146.200 ;
        RECT 12.600 146.100 13.000 146.200 ;
        RECT 11.800 145.800 13.000 146.100 ;
        RECT 11.000 144.200 11.300 145.800 ;
        RECT 13.400 144.800 13.800 145.200 ;
        RECT 13.400 144.200 13.700 144.800 ;
        RECT 11.000 143.800 11.400 144.200 ;
        RECT 13.400 143.800 13.800 144.200 ;
        RECT 10.200 136.800 10.600 137.200 ;
        RECT 10.200 134.200 10.500 136.800 ;
        RECT 11.800 135.800 12.200 136.200 ;
        RECT 11.800 135.200 12.100 135.800 ;
        RECT 11.800 134.800 12.200 135.200 ;
        RECT 10.200 133.800 10.600 134.200 ;
        RECT 11.800 134.100 12.200 134.200 ;
        RECT 12.600 134.100 13.000 134.200 ;
        RECT 11.800 133.800 13.000 134.100 ;
        RECT 10.200 129.200 10.500 133.800 ;
        RECT 13.400 132.200 13.700 143.800 ;
        RECT 14.200 135.100 14.600 135.200 ;
        RECT 15.000 135.100 15.400 135.200 ;
        RECT 14.200 134.800 15.400 135.100 ;
        RECT 15.000 133.800 15.400 134.200 ;
        RECT 13.400 131.800 13.800 132.200 ;
        RECT 15.000 131.200 15.300 133.800 ;
        RECT 15.800 133.100 16.200 135.900 ;
        RECT 16.600 134.200 16.900 153.800 ;
        RECT 18.200 149.200 18.500 153.800 ;
        RECT 19.000 152.100 19.400 157.900 ;
        RECT 22.200 153.100 22.600 155.900 ;
        RECT 19.800 151.800 20.200 152.200 ;
        RECT 20.600 152.100 21.000 152.200 ;
        RECT 21.400 152.100 21.800 152.200 ;
        RECT 23.800 152.100 24.200 157.900 ;
        RECT 25.400 157.800 25.800 158.200 ;
        RECT 25.400 156.800 25.800 157.200 ;
        RECT 25.400 155.200 25.700 156.800 ;
        RECT 27.800 155.200 28.100 166.800 ;
        RECT 30.200 164.200 30.500 166.800 ;
        RECT 35.000 166.200 35.300 166.800 ;
        RECT 35.000 165.800 35.400 166.200 ;
        RECT 36.600 165.800 37.000 166.200 ;
        RECT 36.600 165.200 36.900 165.800 ;
        RECT 31.800 165.100 32.200 165.200 ;
        RECT 32.600 165.100 33.000 165.200 ;
        RECT 31.800 164.800 33.000 165.100 ;
        RECT 36.600 164.800 37.000 165.200 ;
        RECT 37.400 165.100 37.800 167.900 ;
        RECT 30.200 163.800 30.600 164.200 ;
        RECT 25.400 154.800 25.800 155.200 ;
        RECT 27.800 154.800 28.200 155.200 ;
        RECT 28.600 152.100 29.000 157.900 ;
        RECT 30.200 156.200 30.500 163.800 ;
        RECT 32.600 157.800 33.000 158.200 ;
        RECT 30.200 155.800 30.600 156.200 ;
        RECT 31.800 153.100 32.200 155.900 ;
        RECT 32.600 154.200 32.900 157.800 ;
        RECT 32.600 153.800 33.000 154.200 ;
        RECT 31.000 152.100 31.400 152.200 ;
        RECT 31.800 152.100 32.200 152.200 ;
        RECT 33.400 152.100 33.800 157.900 ;
        RECT 35.800 154.800 36.200 155.200 ;
        RECT 35.800 153.200 36.100 154.800 ;
        RECT 35.800 152.800 36.200 153.200 ;
        RECT 20.600 151.800 21.800 152.100 ;
        RECT 31.000 151.800 32.200 152.100 ;
        RECT 18.200 148.800 18.600 149.200 ;
        RECT 19.800 147.200 20.100 151.800 ;
        RECT 36.600 150.200 36.900 164.800 ;
        RECT 39.000 163.100 39.400 168.900 ;
        RECT 40.600 168.800 41.000 169.200 ;
        RECT 38.200 152.100 38.600 157.900 ;
        RECT 41.400 155.200 41.700 171.800 ;
        RECT 42.200 167.800 42.600 168.200 ;
        RECT 42.200 166.200 42.500 167.800 ;
        RECT 43.000 166.800 43.400 167.200 ;
        RECT 43.000 166.200 43.300 166.800 ;
        RECT 42.200 165.800 42.600 166.200 ;
        RECT 43.000 165.800 43.400 166.200 ;
        RECT 43.800 163.100 44.200 168.900 ;
        RECT 46.200 166.200 46.500 173.800 ;
        RECT 50.200 172.100 50.600 177.900 ;
        RECT 51.000 171.100 51.300 179.800 ;
        RECT 57.400 177.200 57.700 186.800 ;
        RECT 59.800 185.800 60.200 186.200 ;
        RECT 61.400 185.800 61.800 186.200 ;
        RECT 62.200 186.100 62.600 186.200 ;
        RECT 63.000 186.100 63.400 186.200 ;
        RECT 62.200 185.800 63.400 186.100 ;
        RECT 64.600 185.800 65.000 186.200 ;
        RECT 58.200 185.100 58.600 185.200 ;
        RECT 59.000 185.100 59.400 185.200 ;
        RECT 58.200 184.800 59.400 185.100 ;
        RECT 59.800 183.200 60.100 185.800 ;
        RECT 60.600 184.800 61.000 185.200 ;
        RECT 59.800 182.800 60.200 183.200 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 57.400 176.800 57.800 177.200 ;
        RECT 59.000 176.800 59.400 177.200 ;
        RECT 52.600 176.200 52.900 176.800 ;
        RECT 52.600 175.800 53.000 176.200 ;
        RECT 56.600 176.100 57.000 176.200 ;
        RECT 57.400 176.100 57.800 176.200 ;
        RECT 56.600 175.800 57.800 176.100 ;
        RECT 54.200 174.800 54.600 175.200 ;
        RECT 55.000 175.100 55.400 175.200 ;
        RECT 55.800 175.100 56.200 175.200 ;
        RECT 55.000 174.800 56.200 175.100 ;
        RECT 58.200 174.800 58.600 175.200 ;
        RECT 54.200 174.200 54.500 174.800 ;
        RECT 53.400 173.800 53.800 174.200 ;
        RECT 54.200 173.800 54.600 174.200 ;
        RECT 53.400 172.200 53.700 173.800 ;
        RECT 50.200 170.800 51.300 171.100 ;
        RECT 51.800 171.800 52.200 172.200 ;
        RECT 53.400 171.800 53.800 172.200 ;
        RECT 50.200 166.200 50.500 170.800 ;
        RECT 51.800 167.200 52.100 171.800 ;
        RECT 58.200 171.200 58.500 174.800 ;
        RECT 59.000 174.200 59.300 176.800 ;
        RECT 60.600 175.200 60.900 184.800 ;
        RECT 61.400 180.200 61.700 185.800 ;
        RECT 64.600 185.200 64.900 185.800 ;
        RECT 62.200 184.800 62.600 185.200 ;
        RECT 64.600 184.800 65.000 185.200 ;
        RECT 61.400 179.800 61.800 180.200 ;
        RECT 59.800 174.800 60.200 175.200 ;
        RECT 60.600 174.800 61.000 175.200 ;
        RECT 59.800 174.200 60.100 174.800 ;
        RECT 59.000 173.800 59.400 174.200 ;
        RECT 59.800 173.800 60.200 174.200 ;
        RECT 56.600 170.800 57.000 171.200 ;
        RECT 58.200 170.800 58.600 171.200 ;
        RECT 53.400 168.100 53.800 168.200 ;
        RECT 54.200 168.100 54.600 168.200 ;
        RECT 53.400 167.800 54.600 168.100 ;
        RECT 51.800 166.800 52.200 167.200 ;
        RECT 52.600 166.800 53.000 167.200 ;
        RECT 52.600 166.200 52.900 166.800 ;
        RECT 56.600 166.200 56.900 170.800 ;
        RECT 59.000 167.200 59.300 173.800 ;
        RECT 57.400 167.100 57.800 167.200 ;
        RECT 58.200 167.100 58.600 167.200 ;
        RECT 57.400 166.800 58.600 167.100 ;
        RECT 59.000 166.800 59.400 167.200 ;
        RECT 61.400 166.200 61.700 179.800 ;
        RECT 62.200 179.200 62.500 184.800 ;
        RECT 63.800 181.800 64.200 182.200 ;
        RECT 62.200 178.800 62.600 179.200 ;
        RECT 63.000 175.800 63.400 176.200 ;
        RECT 63.000 175.200 63.300 175.800 ;
        RECT 63.000 174.800 63.400 175.200 ;
        RECT 62.200 168.800 62.600 169.200 ;
        RECT 62.200 166.200 62.500 168.800 ;
        RECT 46.200 165.800 46.600 166.200 ;
        RECT 47.800 165.800 48.200 166.200 ;
        RECT 50.200 165.800 50.600 166.200 ;
        RECT 51.000 166.100 51.400 166.200 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 51.000 165.800 52.200 166.100 ;
        RECT 52.600 165.800 53.000 166.200 ;
        RECT 56.600 165.800 57.000 166.200 ;
        RECT 57.400 165.800 57.800 166.200 ;
        RECT 61.400 165.800 61.800 166.200 ;
        RECT 62.200 165.800 62.600 166.200 ;
        RECT 42.200 160.800 42.600 161.200 ;
        RECT 41.400 154.800 41.800 155.200 ;
        RECT 42.200 154.100 42.500 160.800 ;
        RECT 46.200 157.200 46.500 165.800 ;
        RECT 47.800 165.200 48.100 165.800 ;
        RECT 56.600 165.200 56.900 165.800 ;
        RECT 47.800 164.800 48.200 165.200 ;
        RECT 54.200 165.100 54.600 165.200 ;
        RECT 55.000 165.100 55.400 165.200 ;
        RECT 54.200 164.800 55.400 165.100 ;
        RECT 56.600 164.800 57.000 165.200 ;
        RECT 49.400 161.800 49.800 162.200 ;
        RECT 43.800 157.100 44.200 157.200 ;
        RECT 44.600 157.100 45.000 157.200 ;
        RECT 43.800 156.800 45.000 157.100 ;
        RECT 46.200 156.800 46.600 157.200 ;
        RECT 46.200 155.800 46.600 156.200 ;
        RECT 43.800 155.100 44.200 155.200 ;
        RECT 43.800 154.800 44.900 155.100 ;
        RECT 41.400 153.800 42.500 154.100 ;
        RECT 43.000 154.100 43.400 154.200 ;
        RECT 43.800 154.100 44.200 154.200 ;
        RECT 43.000 153.800 44.200 154.100 ;
        RECT 40.600 151.800 41.000 152.200 ;
        RECT 40.600 151.200 40.900 151.800 ;
        RECT 40.600 150.800 41.000 151.200 ;
        RECT 23.800 149.800 24.200 150.200 ;
        RECT 36.600 149.800 37.000 150.200 ;
        RECT 23.000 148.800 23.400 149.200 ;
        RECT 23.000 148.200 23.300 148.800 ;
        RECT 23.800 148.200 24.100 149.800 ;
        RECT 39.000 148.800 39.400 149.200 ;
        RECT 20.600 147.800 21.000 148.200 ;
        RECT 23.000 147.800 23.400 148.200 ;
        RECT 23.800 147.800 24.200 148.200 ;
        RECT 25.400 147.800 25.800 148.200 ;
        RECT 36.600 147.800 37.000 148.200 ;
        RECT 20.600 147.200 20.900 147.800 ;
        RECT 19.800 146.800 20.200 147.200 ;
        RECT 20.600 146.800 21.000 147.200 ;
        RECT 25.400 147.100 25.700 147.800 ;
        RECT 36.600 147.200 36.900 147.800 ;
        RECT 39.000 147.200 39.300 148.800 ;
        RECT 30.200 147.100 30.600 147.200 ;
        RECT 31.000 147.100 31.400 147.200 ;
        RECT 25.400 146.800 26.500 147.100 ;
        RECT 30.200 146.800 31.400 147.100 ;
        RECT 33.400 147.100 33.800 147.200 ;
        RECT 34.200 147.100 34.600 147.200 ;
        RECT 33.400 146.800 34.600 147.100 ;
        RECT 35.800 147.100 36.200 147.200 ;
        RECT 36.600 147.100 37.000 147.200 ;
        RECT 35.800 146.800 37.000 147.100 ;
        RECT 39.000 146.800 39.400 147.200 ;
        RECT 17.400 146.100 17.800 146.200 ;
        RECT 18.200 146.100 18.600 146.200 ;
        RECT 17.400 145.800 18.600 146.100 ;
        RECT 17.400 144.800 17.800 145.200 ;
        RECT 18.200 144.800 18.600 145.200 ;
        RECT 17.400 144.200 17.700 144.800 ;
        RECT 18.200 144.200 18.500 144.800 ;
        RECT 17.400 143.800 17.800 144.200 ;
        RECT 18.200 143.800 18.600 144.200 ;
        RECT 16.600 133.800 17.000 134.200 ;
        RECT 17.400 132.100 17.800 137.900 ;
        RECT 18.200 132.800 18.600 133.200 ;
        RECT 15.000 130.800 15.400 131.200 ;
        RECT 10.200 128.800 10.600 129.200 ;
        RECT 9.400 125.800 9.800 126.200 ;
        RECT 9.400 125.200 9.700 125.800 ;
        RECT 9.400 124.800 9.800 125.200 ;
        RECT 11.000 123.100 11.400 128.900 ;
        RECT 13.400 128.800 13.800 129.200 ;
        RECT 13.400 128.200 13.700 128.800 ;
        RECT 11.800 127.800 12.200 128.200 ;
        RECT 11.800 127.200 12.100 127.800 ;
        RECT 11.800 126.800 12.200 127.200 ;
        RECT 12.600 125.100 13.000 127.900 ;
        RECT 13.400 127.800 13.800 128.200 ;
        RECT 15.000 125.100 15.400 127.900 ;
        RECT 16.600 123.100 17.000 128.900 ;
        RECT 18.200 127.200 18.500 132.800 ;
        RECT 19.800 128.200 20.100 146.800 ;
        RECT 20.600 146.100 21.000 146.200 ;
        RECT 21.400 146.100 21.800 146.200 ;
        RECT 20.600 145.800 21.800 146.100 ;
        RECT 25.400 145.800 25.800 146.200 ;
        RECT 25.400 145.200 25.700 145.800 ;
        RECT 26.200 145.200 26.500 146.800 ;
        RECT 27.800 145.800 28.200 146.200 ;
        RECT 28.600 146.100 29.000 146.200 ;
        RECT 29.400 146.100 29.800 146.200 ;
        RECT 28.600 145.800 29.800 146.100 ;
        RECT 31.800 145.800 32.200 146.200 ;
        RECT 32.600 145.800 33.000 146.200 ;
        RECT 34.200 145.800 34.600 146.200 ;
        RECT 39.800 145.800 40.200 146.200 ;
        RECT 22.200 145.100 22.600 145.200 ;
        RECT 23.000 145.100 23.400 145.200 ;
        RECT 22.200 144.800 23.400 145.100 ;
        RECT 24.600 144.800 25.000 145.200 ;
        RECT 25.400 144.800 25.800 145.200 ;
        RECT 26.200 144.800 26.600 145.200 ;
        RECT 24.600 139.200 24.900 144.800 ;
        RECT 27.800 144.200 28.100 145.800 ;
        RECT 30.200 145.100 30.600 145.200 ;
        RECT 31.000 145.100 31.400 145.200 ;
        RECT 30.200 144.800 31.400 145.100 ;
        RECT 27.800 143.800 28.200 144.200 ;
        RECT 28.600 144.100 29.000 144.200 ;
        RECT 29.400 144.100 29.800 144.200 ;
        RECT 28.600 143.800 29.800 144.100 ;
        RECT 24.600 138.800 25.000 139.200 ;
        RECT 26.200 138.800 26.600 139.200 ;
        RECT 20.600 135.800 21.000 136.200 ;
        RECT 20.600 135.200 20.900 135.800 ;
        RECT 20.600 134.800 21.000 135.200 ;
        RECT 21.400 133.800 21.800 134.200 ;
        RECT 21.400 133.200 21.700 133.800 ;
        RECT 21.400 132.800 21.800 133.200 ;
        RECT 22.200 132.100 22.600 137.900 ;
        RECT 26.200 135.200 26.500 138.800 ;
        RECT 27.800 136.800 28.200 137.200 ;
        RECT 27.800 136.200 28.100 136.800 ;
        RECT 27.000 135.800 27.400 136.200 ;
        RECT 27.800 135.800 28.200 136.200 ;
        RECT 27.000 135.200 27.300 135.800 ;
        RECT 25.400 134.800 25.800 135.200 ;
        RECT 26.200 134.800 26.600 135.200 ;
        RECT 27.000 134.800 27.400 135.200 ;
        RECT 25.400 134.200 25.700 134.800 ;
        RECT 25.400 133.800 25.800 134.200 ;
        RECT 25.400 133.200 25.700 133.800 ;
        RECT 25.400 132.800 25.800 133.200 ;
        RECT 19.800 127.800 20.200 128.200 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 19.000 126.100 19.400 126.200 ;
        RECT 19.800 126.100 20.200 126.200 ;
        RECT 19.000 125.800 20.200 126.100 ;
        RECT 21.400 123.100 21.800 128.900 ;
        RECT 23.800 128.100 24.200 128.200 ;
        RECT 24.600 128.100 25.000 128.200 ;
        RECT 23.800 127.800 25.000 128.100 ;
        RECT 26.200 128.100 26.500 134.800 ;
        RECT 28.600 133.100 29.000 135.900 ;
        RECT 29.400 134.800 29.800 135.200 ;
        RECT 29.400 134.200 29.700 134.800 ;
        RECT 29.400 133.800 29.800 134.200 ;
        RECT 30.200 132.100 30.600 137.900 ;
        RECT 31.000 137.800 31.400 138.200 ;
        RECT 26.200 127.800 27.300 128.100 ;
        RECT 26.200 126.800 26.600 127.200 ;
        RECT 26.200 125.200 26.500 126.800 ;
        RECT 27.000 126.200 27.300 127.800 ;
        RECT 31.000 126.200 31.300 137.800 ;
        RECT 31.800 136.200 32.100 145.800 ;
        RECT 32.600 138.200 32.900 145.800 ;
        RECT 32.600 137.800 33.000 138.200 ;
        RECT 34.200 137.200 34.500 145.800 ;
        RECT 39.800 144.200 40.100 145.800 ;
        RECT 41.400 145.200 41.700 153.800 ;
        RECT 42.200 152.800 42.600 153.200 ;
        RECT 42.200 149.200 42.500 152.800 ;
        RECT 44.600 149.200 44.900 154.800 ;
        RECT 46.200 153.200 46.500 155.800 ;
        RECT 49.400 155.200 49.700 161.800 ;
        RECT 53.400 158.800 53.800 159.200 ;
        RECT 53.400 155.200 53.700 158.800 ;
        RECT 55.000 156.800 55.400 157.200 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 49.400 154.800 49.800 155.200 ;
        RECT 51.800 155.100 52.200 155.200 ;
        RECT 52.600 155.100 53.000 155.200 ;
        RECT 51.800 154.800 53.000 155.100 ;
        RECT 53.400 154.800 53.800 155.200 ;
        RECT 47.800 154.200 48.100 154.800 ;
        RECT 47.800 153.800 48.200 154.200 ;
        RECT 48.600 153.800 49.000 154.200 ;
        RECT 46.200 152.800 46.600 153.200 ;
        RECT 46.200 152.200 46.500 152.800 ;
        RECT 46.200 151.800 46.600 152.200 ;
        RECT 42.200 148.800 42.600 149.200 ;
        RECT 44.600 148.800 45.000 149.200 ;
        RECT 47.800 148.100 48.200 148.200 ;
        RECT 48.600 148.100 48.900 153.800 ;
        RECT 54.200 153.100 54.600 155.900 ;
        RECT 55.000 154.200 55.300 156.800 ;
        RECT 55.000 153.800 55.400 154.200 ;
        RECT 47.800 147.800 48.900 148.100 ;
        RECT 51.000 151.800 51.400 152.200 ;
        RECT 51.800 151.800 52.200 152.200 ;
        RECT 55.800 152.100 56.200 157.900 ;
        RECT 57.400 152.200 57.700 165.800 ;
        RECT 59.800 165.100 60.200 165.200 ;
        RECT 60.600 165.100 61.000 165.200 ;
        RECT 59.800 164.800 61.000 165.100 ;
        RECT 61.400 159.200 61.700 165.800 ;
        RECT 63.800 163.200 64.100 181.800 ;
        RECT 65.400 175.200 65.700 202.800 ;
        RECT 67.000 202.200 67.300 206.800 ;
        RECT 67.800 206.100 68.200 206.200 ;
        RECT 68.600 206.100 69.000 206.200 ;
        RECT 67.800 205.800 69.000 206.100 ;
        RECT 71.000 203.100 71.400 208.900 ;
        RECT 75.000 205.800 75.400 206.200 ;
        RECT 67.000 201.800 67.400 202.200 ;
        RECT 73.400 201.800 73.800 202.200 ;
        RECT 74.200 201.800 74.600 202.200 ;
        RECT 73.400 201.200 73.700 201.800 ;
        RECT 73.400 200.800 73.800 201.200 ;
        RECT 74.200 200.100 74.500 201.800 ;
        RECT 73.400 199.800 74.500 200.100 ;
        RECT 66.200 195.800 66.600 196.200 ;
        RECT 66.200 189.200 66.500 195.800 ;
        RECT 67.800 192.100 68.200 197.900 ;
        RECT 73.400 196.200 73.700 199.800 ;
        RECT 75.000 199.200 75.300 205.800 ;
        RECT 76.600 203.100 77.000 208.900 ;
        RECT 77.400 205.800 77.800 206.200 ;
        RECT 80.600 205.900 81.000 206.300 ;
        RECT 77.400 202.200 77.700 205.800 ;
        RECT 77.400 201.800 77.800 202.200 ;
        RECT 77.400 200.800 77.800 201.200 ;
        RECT 75.000 198.800 75.400 199.200 ;
        RECT 77.400 197.200 77.700 200.800 ;
        RECT 77.400 196.800 77.800 197.200 ;
        RECT 80.600 197.100 80.900 205.900 ;
        RECT 81.400 203.100 81.800 208.900 ;
        RECT 83.800 208.800 84.200 209.200 ;
        RECT 151.000 209.100 151.400 209.200 ;
        RECT 151.800 209.100 152.200 209.200 ;
        RECT 82.200 207.800 82.600 208.200 ;
        RECT 82.200 207.200 82.500 207.800 ;
        RECT 82.200 206.800 82.600 207.200 ;
        RECT 83.000 205.100 83.400 207.900 ;
        RECT 83.800 207.200 84.100 208.800 ;
        RECT 83.800 206.800 84.200 207.200 ;
        RECT 89.400 206.800 89.800 207.200 ;
        RECT 84.600 205.800 85.000 206.200 ;
        RECT 87.800 206.100 88.200 206.200 ;
        RECT 88.600 206.100 89.000 206.200 ;
        RECT 87.800 205.800 89.000 206.100 ;
        RECT 83.800 201.800 84.200 202.200 ;
        RECT 82.200 198.800 82.600 199.200 ;
        RECT 80.600 196.800 81.700 197.100 ;
        RECT 73.400 195.800 73.800 196.200 ;
        RECT 79.000 195.800 79.400 196.200 ;
        RECT 80.600 195.800 81.000 196.200 ;
        RECT 71.000 194.800 71.400 195.200 ;
        RECT 71.800 194.800 72.200 195.200 ;
        RECT 72.600 194.800 73.000 195.200 ;
        RECT 71.000 194.200 71.300 194.800 ;
        RECT 71.800 194.200 72.100 194.800 ;
        RECT 72.600 194.200 72.900 194.800 ;
        RECT 71.000 193.800 71.400 194.200 ;
        RECT 71.800 193.800 72.200 194.200 ;
        RECT 72.600 193.800 73.000 194.200 ;
        RECT 70.200 191.800 70.600 192.200 ;
        RECT 66.200 188.800 66.600 189.200 ;
        RECT 70.200 188.200 70.500 191.800 ;
        RECT 66.200 187.800 66.600 188.200 ;
        RECT 70.200 187.800 70.600 188.200 ;
        RECT 66.200 185.200 66.500 187.800 ;
        RECT 68.600 187.100 69.000 187.200 ;
        RECT 69.400 187.100 69.800 187.200 ;
        RECT 68.600 186.800 69.800 187.100 ;
        RECT 71.000 187.100 71.400 187.200 ;
        RECT 71.800 187.100 72.200 187.200 ;
        RECT 71.000 186.800 72.200 187.100 ;
        RECT 72.600 186.800 73.000 187.200 ;
        RECT 67.800 185.800 68.200 186.200 ;
        RECT 68.600 185.800 69.000 186.200 ;
        RECT 66.200 184.800 66.600 185.200 ;
        RECT 66.200 178.200 66.500 184.800 ;
        RECT 67.000 183.800 67.400 184.200 ;
        RECT 66.200 177.800 66.600 178.200 ;
        RECT 66.200 175.800 66.600 176.200 ;
        RECT 66.200 175.200 66.500 175.800 ;
        RECT 65.400 174.800 65.800 175.200 ;
        RECT 66.200 174.800 66.600 175.200 ;
        RECT 67.000 175.100 67.300 183.800 ;
        RECT 67.800 183.200 68.100 185.800 ;
        RECT 67.800 182.800 68.200 183.200 ;
        RECT 68.600 179.200 68.900 185.800 ;
        RECT 71.000 181.800 71.400 182.200 ;
        RECT 69.400 179.800 69.800 180.200 ;
        RECT 68.600 178.800 69.000 179.200 ;
        RECT 69.400 178.200 69.700 179.800 ;
        RECT 69.400 177.800 69.800 178.200 ;
        RECT 69.400 175.200 69.700 177.800 ;
        RECT 70.200 175.800 70.600 176.200 ;
        RECT 70.200 175.200 70.500 175.800 ;
        RECT 67.800 175.100 68.200 175.200 ;
        RECT 67.000 174.800 68.200 175.100 ;
        RECT 68.600 174.800 69.000 175.200 ;
        RECT 69.400 174.800 69.800 175.200 ;
        RECT 70.200 174.800 70.600 175.200 ;
        RECT 68.600 174.200 68.900 174.800 ;
        RECT 67.000 173.800 67.400 174.200 ;
        RECT 68.600 173.800 69.000 174.200 ;
        RECT 64.600 167.800 65.000 168.200 ;
        RECT 64.600 166.200 64.900 167.800 ;
        RECT 66.200 166.800 66.600 167.200 ;
        RECT 66.200 166.200 66.500 166.800 ;
        RECT 67.000 166.200 67.300 173.800 ;
        RECT 67.800 168.100 68.200 168.200 ;
        RECT 68.600 168.100 69.000 168.200 ;
        RECT 67.800 167.800 69.000 168.100 ;
        RECT 71.000 167.200 71.300 181.800 ;
        RECT 72.600 175.200 72.900 186.800 ;
        RECT 73.400 186.200 73.700 195.800 ;
        RECT 79.000 195.200 79.300 195.800 ;
        RECT 75.000 195.100 75.400 195.200 ;
        RECT 75.800 195.100 76.200 195.200 ;
        RECT 75.000 194.800 76.200 195.100 ;
        RECT 79.000 194.800 79.400 195.200 ;
        RECT 80.600 194.200 80.900 195.800 ;
        RECT 81.400 195.200 81.700 196.800 ;
        RECT 82.200 195.200 82.500 198.800 ;
        RECT 81.400 194.800 81.800 195.200 ;
        RECT 82.200 194.800 82.600 195.200 ;
        RECT 74.200 193.800 74.600 194.200 ;
        RECT 79.800 193.800 80.200 194.200 ;
        RECT 80.600 193.800 81.000 194.200 ;
        RECT 74.200 191.200 74.500 193.800 ;
        RECT 79.800 193.100 80.100 193.800 ;
        RECT 79.800 192.800 80.900 193.100 ;
        RECT 74.200 190.800 74.600 191.200 ;
        RECT 74.200 187.200 74.500 190.800 ;
        RECT 80.600 190.200 80.900 192.800 ;
        RECT 80.600 189.800 81.000 190.200 ;
        RECT 80.600 189.200 80.900 189.800 ;
        RECT 74.200 186.800 74.600 187.200 ;
        RECT 73.400 185.800 73.800 186.200 ;
        RECT 75.000 186.100 75.400 186.200 ;
        RECT 75.800 186.100 76.200 186.200 ;
        RECT 75.000 185.800 76.200 186.100 ;
        RECT 76.600 185.800 77.000 186.200 ;
        RECT 77.400 185.800 77.800 186.200 ;
        RECT 76.600 185.200 76.900 185.800 ;
        RECT 76.600 184.800 77.000 185.200 ;
        RECT 77.400 184.200 77.700 185.800 ;
        RECT 75.800 183.800 76.200 184.200 ;
        RECT 77.400 183.800 77.800 184.200 ;
        RECT 75.800 179.200 76.100 183.800 ;
        RECT 79.800 183.100 80.200 188.900 ;
        RECT 80.600 188.800 81.000 189.200 ;
        RECT 82.200 184.200 82.500 194.800 ;
        RECT 83.000 193.800 83.400 194.200 ;
        RECT 82.200 183.800 82.600 184.200 ;
        RECT 82.200 180.200 82.500 183.800 ;
        RECT 82.200 179.800 82.600 180.200 ;
        RECT 75.800 178.800 76.200 179.200 ;
        RECT 72.600 174.800 73.000 175.200 ;
        RECT 73.400 174.800 73.800 175.200 ;
        RECT 73.400 173.200 73.700 174.800 ;
        RECT 73.400 172.800 73.800 173.200 ;
        RECT 77.400 173.100 77.800 175.900 ;
        RECT 78.200 173.800 78.600 174.200 ;
        RECT 71.800 171.800 72.200 172.200 ;
        RECT 76.600 171.800 77.000 172.200 ;
        RECT 71.000 166.800 71.400 167.200 ;
        RECT 64.600 165.800 65.000 166.200 ;
        RECT 66.200 165.800 66.600 166.200 ;
        RECT 67.000 165.800 67.400 166.200 ;
        RECT 68.600 166.100 69.000 166.200 ;
        RECT 69.400 166.100 69.800 166.200 ;
        RECT 68.600 165.800 69.800 166.100 ;
        RECT 70.200 165.800 70.600 166.200 ;
        RECT 70.200 165.200 70.500 165.800 ;
        RECT 70.200 164.800 70.600 165.200 ;
        RECT 63.800 162.800 64.200 163.200 ;
        RECT 63.800 161.800 64.200 162.200 ;
        RECT 63.800 159.200 64.100 161.800 ;
        RECT 61.400 158.800 61.800 159.200 ;
        RECT 63.800 158.800 64.200 159.200 ;
        RECT 58.200 155.800 58.600 156.200 ;
        RECT 58.200 155.200 58.500 155.800 ;
        RECT 58.200 154.800 58.600 155.200 ;
        RECT 58.200 153.800 58.600 154.200 ;
        RECT 57.400 151.800 57.800 152.200 ;
        RECT 47.800 147.200 48.100 147.800 ;
        RECT 44.600 147.100 45.000 147.200 ;
        RECT 45.400 147.100 45.800 147.200 ;
        RECT 44.600 146.800 45.800 147.100 ;
        RECT 47.800 146.800 48.200 147.200 ;
        RECT 43.800 145.800 44.200 146.200 ;
        RECT 44.600 145.800 45.000 146.200 ;
        RECT 47.000 146.100 47.400 146.200 ;
        RECT 47.800 146.100 48.200 146.200 ;
        RECT 47.000 145.800 48.200 146.100 ;
        RECT 41.400 144.800 41.800 145.200 ;
        RECT 42.200 145.100 42.600 145.200 ;
        RECT 43.000 145.100 43.400 145.200 ;
        RECT 42.200 144.800 43.400 145.100 ;
        RECT 39.800 143.800 40.200 144.200 ;
        RECT 43.800 143.200 44.100 145.800 ;
        RECT 44.600 145.200 44.900 145.800 ;
        RECT 44.600 144.800 45.000 145.200 ;
        RECT 45.400 145.100 45.800 145.200 ;
        RECT 46.200 145.100 46.600 145.200 ;
        RECT 45.400 144.800 46.600 145.100 ;
        RECT 43.800 142.800 44.200 143.200 ;
        RECT 39.800 141.800 40.200 142.200 ;
        RECT 39.800 140.200 40.100 141.800 ;
        RECT 39.800 139.800 40.200 140.200 ;
        RECT 39.800 138.800 40.200 139.200 ;
        RECT 37.400 138.100 37.800 138.200 ;
        RECT 38.200 138.100 38.600 138.200 ;
        RECT 34.200 136.800 34.600 137.200 ;
        RECT 31.800 135.800 32.200 136.200 ;
        RECT 32.600 135.100 33.000 135.200 ;
        RECT 33.400 135.100 33.800 135.200 ;
        RECT 32.600 134.800 33.800 135.100 ;
        RECT 33.400 133.800 33.800 134.200 ;
        RECT 31.800 126.800 32.200 127.200 ;
        RECT 31.800 126.200 32.100 126.800 ;
        RECT 27.000 125.800 27.400 126.200 ;
        RECT 27.800 126.100 28.200 126.200 ;
        RECT 28.600 126.100 29.000 126.200 ;
        RECT 27.800 125.800 29.000 126.100 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 31.800 125.800 32.200 126.200 ;
        RECT 26.200 124.800 26.600 125.200 ;
        RECT 14.200 121.800 14.600 122.200 ;
        RECT 23.800 122.100 24.200 122.200 ;
        RECT 24.600 122.100 25.000 122.200 ;
        RECT 23.800 121.800 25.000 122.100 ;
        RECT 25.400 121.800 25.800 122.200 ;
        RECT 14.200 118.200 14.500 121.800 ;
        RECT 10.200 114.800 10.600 115.200 ;
        RECT 10.200 111.100 10.500 114.800 ;
        RECT 11.000 112.100 11.400 117.900 ;
        RECT 14.200 117.800 14.600 118.200 ;
        RECT 23.000 117.800 23.400 118.200 ;
        RECT 13.400 117.100 13.800 117.200 ;
        RECT 14.200 117.100 14.600 117.200 ;
        RECT 13.400 116.800 14.600 117.100 ;
        RECT 17.400 116.800 17.800 117.200 ;
        RECT 17.400 116.200 17.700 116.800 ;
        RECT 17.400 115.800 17.800 116.200 ;
        RECT 20.600 115.800 21.000 116.200 ;
        RECT 15.000 114.800 15.400 115.200 ;
        RECT 15.800 115.100 16.200 115.200 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 15.800 114.800 17.000 115.100 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 15.000 114.200 15.300 114.800 ;
        RECT 19.000 114.200 19.300 114.800 ;
        RECT 14.200 113.800 14.600 114.200 ;
        RECT 15.000 113.800 15.400 114.200 ;
        RECT 17.400 113.800 17.800 114.200 ;
        RECT 19.000 113.800 19.400 114.200 ;
        RECT 19.800 113.800 20.200 114.200 ;
        RECT 10.200 110.800 11.300 111.100 ;
        RECT 8.600 107.800 9.000 108.200 ;
        RECT 3.000 106.800 3.400 107.200 ;
        RECT 3.800 107.100 4.200 107.200 ;
        RECT 4.600 107.100 5.000 107.200 ;
        RECT 3.800 106.800 5.000 107.100 ;
        RECT 8.600 107.100 9.000 107.200 ;
        RECT 9.400 107.100 9.800 107.200 ;
        RECT 8.600 106.800 9.800 107.100 ;
        RECT 3.000 106.200 3.300 106.800 ;
        RECT 3.000 105.800 3.400 106.200 ;
        RECT 4.600 105.800 5.000 106.200 ;
        RECT 9.400 105.800 9.800 106.200 ;
        RECT 4.600 105.200 4.900 105.800 ;
        RECT 4.600 104.800 5.000 105.200 ;
        RECT 6.200 104.800 6.600 105.200 ;
        RECT 7.800 105.100 8.200 105.200 ;
        RECT 8.600 105.100 9.000 105.200 ;
        RECT 7.800 104.800 9.000 105.100 ;
        RECT 6.200 101.200 6.500 104.800 ;
        RECT 9.400 102.200 9.700 105.800 ;
        RECT 10.200 105.100 10.600 107.900 ;
        RECT 11.000 107.200 11.300 110.800 ;
        RECT 11.000 106.800 11.400 107.200 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 6.200 100.800 6.600 101.200 ;
        RECT 0.600 98.800 1.700 99.100 ;
        RECT 1.400 96.200 1.700 98.800 ;
        RECT 1.400 95.800 1.800 96.200 ;
        RECT 3.000 92.100 3.400 97.900 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 6.200 94.800 7.400 95.100 ;
        RECT 7.000 94.700 7.400 94.800 ;
        RECT 4.600 93.800 5.000 94.200 ;
        RECT 0.600 85.100 1.000 87.900 ;
        RECT 2.200 83.100 2.600 88.900 ;
        RECT 4.600 87.200 4.900 93.800 ;
        RECT 7.800 92.100 8.200 97.900 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 8.600 93.200 8.900 93.800 ;
        RECT 8.600 92.800 9.000 93.200 ;
        RECT 9.400 93.100 9.800 95.900 ;
        RECT 10.200 95.800 10.600 96.200 ;
        RECT 10.200 94.200 10.500 95.800 ;
        RECT 11.000 94.200 11.300 106.800 ;
        RECT 11.800 103.100 12.200 108.900 ;
        RECT 14.200 103.200 14.500 113.800 ;
        RECT 15.800 107.800 16.200 108.200 ;
        RECT 15.000 106.800 15.400 107.200 ;
        RECT 15.000 106.200 15.300 106.800 ;
        RECT 15.000 105.800 15.400 106.200 ;
        RECT 14.200 102.800 14.600 103.200 ;
        RECT 11.800 96.100 12.200 96.200 ;
        RECT 12.600 96.100 13.000 96.200 ;
        RECT 11.800 95.800 13.000 96.100 ;
        RECT 12.600 95.100 13.000 95.200 ;
        RECT 13.400 95.100 13.800 95.200 ;
        RECT 12.600 94.800 13.800 95.100 ;
        RECT 14.200 95.100 14.600 95.200 ;
        RECT 15.000 95.100 15.400 95.200 ;
        RECT 14.200 94.800 15.400 95.100 ;
        RECT 15.800 94.200 16.100 107.800 ;
        RECT 16.600 103.100 17.000 108.900 ;
        RECT 16.600 95.800 17.000 96.200 ;
        RECT 16.600 95.200 16.900 95.800 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 10.200 93.800 10.600 94.200 ;
        RECT 11.000 93.800 11.400 94.200 ;
        RECT 15.000 93.800 15.400 94.200 ;
        RECT 15.800 93.800 16.200 94.200 ;
        RECT 14.200 93.100 14.600 93.200 ;
        RECT 15.000 93.100 15.300 93.800 ;
        RECT 14.200 92.800 15.300 93.100 ;
        RECT 12.600 90.800 13.000 91.200 ;
        RECT 4.600 86.800 5.000 87.200 ;
        RECT 4.600 86.100 5.000 86.200 ;
        RECT 5.400 86.100 5.800 86.200 ;
        RECT 4.600 85.800 5.800 86.100 ;
        RECT 6.200 85.800 6.600 86.200 ;
        RECT 0.600 73.100 1.000 75.900 ;
        RECT 2.200 72.100 2.600 77.900 ;
        RECT 4.600 76.800 5.000 77.200 ;
        RECT 4.600 75.200 4.900 76.800 ;
        RECT 6.200 75.200 6.500 85.800 ;
        RECT 7.000 83.100 7.400 88.900 ;
        RECT 9.400 88.800 9.800 89.200 ;
        RECT 11.800 88.800 12.200 89.200 ;
        RECT 9.400 88.200 9.700 88.800 ;
        RECT 9.400 87.800 9.800 88.200 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 11.000 86.100 11.400 86.200 ;
        RECT 10.200 85.800 11.400 86.100 ;
        RECT 10.200 85.100 10.600 85.200 ;
        RECT 11.000 85.100 11.400 85.200 ;
        RECT 10.200 84.800 11.400 85.100 ;
        RECT 10.200 83.800 10.600 84.200 ;
        RECT 4.600 74.800 5.000 75.200 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 5.400 73.800 5.800 74.200 ;
        RECT 4.600 65.100 5.000 67.900 ;
        RECT 5.400 67.200 5.700 73.800 ;
        RECT 7.000 72.100 7.400 77.900 ;
        RECT 9.400 76.800 9.800 77.200 ;
        RECT 9.400 76.200 9.700 76.800 ;
        RECT 9.400 75.800 9.800 76.200 ;
        RECT 10.200 74.200 10.500 83.800 ;
        RECT 11.000 77.800 11.400 78.200 ;
        RECT 11.000 77.200 11.300 77.800 ;
        RECT 11.000 76.800 11.400 77.200 ;
        RECT 11.000 74.800 11.400 75.200 ;
        RECT 10.200 73.800 10.600 74.200 ;
        RECT 5.400 66.800 5.800 67.200 ;
        RECT 0.600 63.800 1.000 64.200 ;
        RECT 3.000 64.100 3.400 64.200 ;
        RECT 3.800 64.100 4.200 64.200 ;
        RECT 3.000 63.800 4.200 64.100 ;
        RECT 0.600 55.200 0.900 63.800 ;
        RECT 6.200 63.100 6.600 68.900 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 0.600 54.800 1.000 55.200 ;
        RECT 3.000 54.800 3.400 55.200 ;
        RECT 3.000 54.200 3.300 54.800 ;
        RECT 3.000 53.800 3.400 54.200 ;
        RECT 3.800 53.100 4.200 55.900 ;
        RECT 5.400 52.100 5.800 57.900 ;
        RECT 7.000 56.800 7.400 57.200 ;
        RECT 7.000 55.200 7.300 56.800 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 7.800 54.200 8.100 66.800 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 9.400 66.100 9.800 66.200 ;
        RECT 8.600 65.800 9.800 66.100 ;
        RECT 10.200 65.100 10.500 73.800 ;
        RECT 11.000 72.200 11.300 74.800 ;
        RECT 11.000 71.800 11.400 72.200 ;
        RECT 9.400 64.800 10.500 65.100 ;
        RECT 8.600 54.800 9.000 55.200 ;
        RECT 7.800 53.800 8.200 54.200 ;
        RECT 0.600 45.100 1.000 47.900 ;
        RECT 2.200 43.100 2.600 48.900 ;
        RECT 3.800 47.800 4.200 48.200 ;
        RECT 3.800 46.200 4.100 47.800 ;
        RECT 3.800 45.800 4.200 46.200 ;
        RECT 6.200 45.800 6.600 46.200 ;
        RECT 6.200 42.200 6.500 45.800 ;
        RECT 7.000 43.100 7.400 48.900 ;
        RECT 6.200 41.800 6.600 42.200 ;
        RECT 0.600 36.100 1.000 36.200 ;
        RECT 1.400 36.100 1.800 36.200 ;
        RECT 0.600 35.800 1.800 36.100 ;
        RECT 2.200 35.800 2.600 36.200 ;
        RECT 7.800 36.100 8.200 36.200 ;
        RECT 8.600 36.100 8.900 54.800 ;
        RECT 9.400 54.200 9.700 64.800 ;
        RECT 11.000 63.100 11.400 68.900 ;
        RECT 9.400 53.800 9.800 54.200 ;
        RECT 10.200 52.100 10.600 57.900 ;
        RECT 10.200 46.800 10.600 47.200 ;
        RECT 10.200 46.200 10.500 46.800 ;
        RECT 11.800 46.200 12.100 88.800 ;
        RECT 12.600 87.200 12.900 90.800 ;
        RECT 13.400 89.800 13.800 90.200 ;
        RECT 13.400 88.200 13.700 89.800 ;
        RECT 13.400 87.800 13.800 88.200 ;
        RECT 12.600 86.800 13.000 87.200 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 12.600 71.200 12.900 85.800 ;
        RECT 13.400 85.200 13.700 87.800 ;
        RECT 14.200 85.800 14.600 86.200 ;
        RECT 14.200 85.200 14.500 85.800 ;
        RECT 13.400 84.800 13.800 85.200 ;
        RECT 14.200 84.800 14.600 85.200 ;
        RECT 15.000 84.200 15.300 92.800 ;
        RECT 15.800 85.200 16.100 93.800 ;
        RECT 16.600 89.200 16.900 94.800 ;
        RECT 17.400 89.200 17.700 113.800 ;
        RECT 19.800 113.200 20.100 113.800 ;
        RECT 20.600 113.200 20.900 115.800 ;
        RECT 23.000 115.200 23.300 117.800 ;
        RECT 25.400 116.100 25.700 121.800 ;
        RECT 27.000 116.200 27.300 125.800 ;
        RECT 29.400 124.800 29.800 125.200 ;
        RECT 29.400 122.200 29.700 124.800 ;
        RECT 31.000 123.200 31.300 125.800 ;
        RECT 32.600 125.100 33.000 127.900 ;
        RECT 33.400 127.200 33.700 133.800 ;
        RECT 34.200 130.100 34.500 136.800 ;
        RECT 35.000 132.100 35.400 137.900 ;
        RECT 37.400 137.800 38.600 138.100 ;
        RECT 39.800 136.200 40.100 138.800 ;
        RECT 43.000 137.800 43.400 138.200 ;
        RECT 43.000 136.200 43.300 137.800 ;
        RECT 43.800 136.200 44.100 142.800 ;
        RECT 49.400 141.800 49.800 142.200 ;
        RECT 39.800 135.800 40.200 136.200 ;
        RECT 43.000 135.800 43.400 136.200 ;
        RECT 43.800 135.800 44.200 136.200 ;
        RECT 46.200 136.100 46.600 136.200 ;
        RECT 46.200 135.800 47.300 136.100 ;
        RECT 39.800 135.200 40.100 135.800 ;
        RECT 39.800 134.800 40.200 135.200 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 41.400 135.100 41.800 135.200 ;
        RECT 40.600 134.800 41.800 135.100 ;
        RECT 43.000 134.200 43.300 135.800 ;
        RECT 44.600 135.100 45.000 135.200 ;
        RECT 45.400 135.100 45.800 135.200 ;
        RECT 44.600 134.800 45.800 135.100 ;
        RECT 39.000 134.100 39.400 134.200 ;
        RECT 39.800 134.100 40.200 134.200 ;
        RECT 39.000 133.800 40.200 134.100 ;
        RECT 43.000 133.800 43.400 134.200 ;
        RECT 44.600 133.800 45.000 134.200 ;
        RECT 45.400 134.100 45.800 134.200 ;
        RECT 46.200 134.100 46.600 134.200 ;
        RECT 45.400 133.800 46.600 134.100 ;
        RECT 34.200 129.800 35.300 130.100 ;
        RECT 33.400 126.800 33.800 127.200 ;
        RECT 31.000 122.800 31.400 123.200 ;
        RECT 34.200 123.100 34.600 128.900 ;
        RECT 29.400 121.800 29.800 122.200 ;
        RECT 29.400 117.200 29.700 121.800 ;
        RECT 29.400 116.800 29.800 117.200 ;
        RECT 31.000 116.800 31.400 117.200 ;
        RECT 25.400 115.800 26.500 116.100 ;
        RECT 27.000 115.800 27.400 116.200 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 24.600 115.100 25.000 115.200 ;
        RECT 25.400 115.100 25.800 115.200 ;
        RECT 24.600 114.800 25.800 115.100 ;
        RECT 26.200 115.100 26.500 115.800 ;
        RECT 27.000 115.100 27.400 115.200 ;
        RECT 26.200 114.800 27.400 115.100 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 22.200 114.100 22.600 114.200 ;
        RECT 23.000 114.100 23.400 114.200 ;
        RECT 22.200 113.800 23.400 114.100 ;
        RECT 25.400 113.800 25.800 114.200 ;
        RECT 26.200 114.100 26.600 114.200 ;
        RECT 27.000 114.100 27.400 114.200 ;
        RECT 26.200 113.800 27.400 114.100 ;
        RECT 19.800 112.800 20.200 113.200 ;
        RECT 20.600 112.800 21.000 113.200 ;
        RECT 25.400 112.200 25.700 113.800 ;
        RECT 21.400 112.100 21.800 112.200 ;
        RECT 22.200 112.100 22.600 112.200 ;
        RECT 21.400 111.800 22.600 112.100 ;
        RECT 23.000 111.800 23.400 112.200 ;
        RECT 25.400 111.800 25.800 112.200 ;
        RECT 27.000 111.800 27.400 112.200 ;
        RECT 23.000 109.200 23.300 111.800 ;
        RECT 19.000 108.800 19.400 109.200 ;
        RECT 23.000 108.800 23.400 109.200 ;
        RECT 26.200 108.800 26.600 109.200 ;
        RECT 19.000 107.200 19.300 108.800 ;
        RECT 19.800 107.800 20.200 108.200 ;
        RECT 19.800 107.200 20.100 107.800 ;
        RECT 19.000 106.800 19.400 107.200 ;
        RECT 19.800 106.800 20.200 107.200 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 23.800 106.800 25.000 107.100 ;
        RECT 25.400 106.800 25.800 107.200 ;
        RECT 25.400 106.200 25.700 106.800 ;
        RECT 26.200 106.200 26.500 108.800 ;
        RECT 20.600 105.800 21.000 106.200 ;
        RECT 21.400 106.100 21.800 106.200 ;
        RECT 22.200 106.100 22.600 106.200 ;
        RECT 21.400 105.800 22.600 106.100 ;
        RECT 25.400 105.800 25.800 106.200 ;
        RECT 26.200 105.800 26.600 106.200 ;
        RECT 20.600 105.200 20.900 105.800 ;
        RECT 20.600 104.800 21.000 105.200 ;
        RECT 23.000 104.800 23.400 105.200 ;
        RECT 23.000 104.200 23.300 104.800 ;
        RECT 19.000 103.800 19.400 104.200 ;
        RECT 23.000 103.800 23.400 104.200 ;
        RECT 19.000 96.200 19.300 103.800 ;
        RECT 19.800 101.800 20.200 102.200 ;
        RECT 26.200 101.800 26.600 102.200 ;
        RECT 19.000 95.800 19.400 96.200 ;
        RECT 19.000 94.800 19.400 95.200 ;
        RECT 19.000 94.200 19.300 94.800 ;
        RECT 19.000 93.800 19.400 94.200 ;
        RECT 16.600 88.800 17.000 89.200 ;
        RECT 17.400 88.800 17.800 89.200 ;
        RECT 16.600 87.800 17.000 88.200 ;
        RECT 16.600 87.200 16.900 87.800 ;
        RECT 16.600 86.800 17.000 87.200 ;
        RECT 17.400 86.200 17.700 88.800 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 15.800 84.800 16.200 85.200 ;
        RECT 15.000 83.800 15.400 84.200 ;
        RECT 13.400 75.800 13.800 76.200 ;
        RECT 15.000 75.800 15.400 76.200 ;
        RECT 13.400 72.200 13.700 75.800 ;
        RECT 15.000 74.200 15.300 75.800 ;
        RECT 15.800 74.200 16.100 84.800 ;
        RECT 19.000 83.800 19.400 84.200 ;
        RECT 19.000 78.200 19.300 83.800 ;
        RECT 19.000 77.800 19.400 78.200 ;
        RECT 16.600 76.800 17.000 77.200 ;
        RECT 19.000 76.800 19.400 77.200 ;
        RECT 16.600 75.200 16.900 76.800 ;
        RECT 19.000 76.200 19.300 76.800 ;
        RECT 19.000 75.800 19.400 76.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 18.200 74.800 18.600 75.200 ;
        RECT 15.000 73.800 15.400 74.200 ;
        RECT 15.800 73.800 16.200 74.200 ;
        RECT 13.400 71.800 13.800 72.200 ;
        RECT 12.600 70.800 13.000 71.200 ;
        RECT 13.400 68.800 13.800 69.200 ;
        RECT 13.400 68.200 13.700 68.800 ;
        RECT 13.400 67.800 13.800 68.200 ;
        RECT 16.600 68.100 16.900 74.800 ;
        RECT 18.200 74.200 18.500 74.800 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 15.800 67.800 16.900 68.100 ;
        RECT 17.400 67.800 17.800 68.200 ;
        RECT 15.800 66.200 16.100 67.800 ;
        RECT 17.400 67.200 17.700 67.800 ;
        RECT 16.600 66.800 17.000 67.200 ;
        RECT 17.400 66.800 17.800 67.200 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 13.400 65.800 14.600 66.100 ;
        RECT 15.800 65.800 16.200 66.200 ;
        RECT 14.200 64.800 14.600 65.200 ;
        RECT 13.400 61.800 13.800 62.200 ;
        RECT 12.600 56.800 13.000 57.200 ;
        RECT 12.600 56.200 12.900 56.800 ;
        RECT 12.600 55.800 13.000 56.200 ;
        RECT 13.400 54.200 13.700 61.800 ;
        RECT 14.200 59.200 14.500 64.800 ;
        RECT 14.200 58.800 14.600 59.200 ;
        RECT 15.000 56.100 15.400 56.200 ;
        RECT 15.800 56.100 16.100 65.800 ;
        RECT 16.600 60.200 16.900 66.800 ;
        RECT 19.800 66.200 20.100 101.800 ;
        RECT 20.600 96.800 21.000 97.200 ;
        RECT 20.600 94.200 20.900 96.800 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 21.400 93.100 21.800 95.900 ;
        RECT 23.000 92.100 23.400 97.900 ;
        RECT 23.800 95.000 24.200 95.100 ;
        RECT 24.600 95.000 25.000 95.100 ;
        RECT 23.800 94.700 25.000 95.000 ;
        RECT 24.600 93.800 25.000 94.200 ;
        RECT 21.400 87.100 21.800 87.200 ;
        RECT 22.200 87.100 22.600 87.200 ;
        RECT 21.400 86.800 22.600 87.100 ;
        RECT 20.600 86.100 21.000 86.200 ;
        RECT 21.400 86.100 21.800 86.200 ;
        RECT 20.600 85.800 21.800 86.100 ;
        RECT 23.800 85.800 24.200 86.200 ;
        RECT 23.800 85.200 24.100 85.800 ;
        RECT 23.800 84.800 24.200 85.200 ;
        RECT 24.600 83.200 24.900 93.800 ;
        RECT 26.200 92.200 26.500 101.800 ;
        RECT 26.200 91.800 26.600 92.200 ;
        RECT 27.000 90.100 27.300 111.800 ;
        RECT 27.800 104.800 28.200 105.200 ;
        RECT 27.800 104.200 28.100 104.800 ;
        RECT 27.800 103.800 28.200 104.200 ;
        RECT 28.600 99.200 28.900 114.800 ;
        RECT 31.000 113.200 31.300 116.800 ;
        RECT 35.000 115.200 35.300 129.800 ;
        RECT 42.200 129.100 42.600 129.200 ;
        RECT 43.000 129.100 43.400 129.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 36.600 126.100 37.000 126.200 ;
        RECT 35.800 125.800 37.000 126.100 ;
        RECT 39.000 123.100 39.400 128.900 ;
        RECT 42.200 128.800 43.400 129.100 ;
        RECT 44.600 128.200 44.900 133.800 ;
        RECT 47.000 132.200 47.300 135.800 ;
        RECT 49.400 135.200 49.700 141.800 ;
        RECT 51.000 138.200 51.300 151.800 ;
        RECT 51.800 146.200 52.100 151.800 ;
        RECT 54.200 149.800 54.600 150.200 ;
        RECT 53.400 146.800 53.800 147.200 ;
        RECT 53.400 146.200 53.700 146.800 ;
        RECT 51.800 145.800 52.200 146.200 ;
        RECT 53.400 145.800 53.800 146.200 ;
        RECT 54.200 141.200 54.500 149.800 ;
        RECT 55.000 145.100 55.400 147.900 ;
        RECT 56.600 143.100 57.000 148.900 ;
        RECT 58.200 147.200 58.500 153.800 ;
        RECT 60.600 152.100 61.000 157.900 ;
        RECT 61.400 157.800 61.800 158.200 ;
        RECT 61.400 157.200 61.700 157.800 ;
        RECT 71.800 157.200 72.100 171.800 ;
        RECT 76.600 170.200 76.900 171.800 ;
        RECT 76.600 169.800 77.000 170.200 ;
        RECT 73.400 168.800 73.800 169.200 ;
        RECT 73.400 166.200 73.700 168.800 ;
        RECT 76.600 167.200 76.900 169.800 ;
        RECT 75.000 166.800 75.400 167.200 ;
        RECT 76.600 166.800 77.000 167.200 ;
        RECT 75.000 166.200 75.300 166.800 ;
        RECT 73.400 165.800 73.800 166.200 ;
        RECT 75.000 165.800 75.400 166.200 ;
        RECT 75.800 165.800 76.200 166.200 ;
        RECT 73.400 165.200 73.700 165.800 ;
        RECT 73.400 164.800 73.800 165.200 ;
        RECT 75.800 164.200 76.100 165.800 ;
        RECT 75.800 163.800 76.200 164.200 ;
        RECT 75.000 161.800 75.400 162.200 ;
        RECT 73.400 159.800 73.800 160.200 ;
        RECT 61.400 156.800 61.800 157.200 ;
        RECT 63.000 157.100 63.400 157.200 ;
        RECT 63.800 157.100 64.200 157.200 ;
        RECT 63.000 156.800 64.200 157.100 ;
        RECT 68.600 156.800 69.000 157.200 ;
        RECT 71.800 156.800 72.200 157.200 ;
        RECT 64.600 156.100 65.000 156.200 ;
        RECT 65.400 156.100 65.800 156.200 ;
        RECT 64.600 155.800 65.800 156.100 ;
        RECT 67.000 156.100 67.400 156.200 ;
        RECT 67.800 156.100 68.200 156.200 ;
        RECT 67.000 155.800 68.200 156.100 ;
        RECT 64.600 155.100 65.000 155.200 ;
        RECT 65.400 155.100 65.800 155.200 ;
        RECT 64.600 154.800 65.800 155.100 ;
        RECT 68.600 154.200 68.900 156.800 ;
        RECT 73.400 155.200 73.700 159.800 ;
        RECT 71.000 154.800 71.400 155.200 ;
        RECT 73.400 154.800 73.800 155.200 ;
        RECT 71.000 154.200 71.300 154.800 ;
        RECT 63.800 153.800 64.200 154.200 ;
        RECT 68.600 153.800 69.000 154.200 ;
        RECT 71.000 153.800 71.400 154.200 ;
        RECT 63.800 149.100 64.100 153.800 ;
        RECT 70.200 151.800 70.600 152.200 ;
        RECT 70.200 150.200 70.500 151.800 ;
        RECT 73.400 151.200 73.700 154.800 ;
        RECT 74.200 153.100 74.600 155.900 ;
        RECT 75.000 154.200 75.300 161.800 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 75.000 152.800 75.400 153.200 ;
        RECT 73.400 150.800 73.800 151.200 ;
        RECT 70.200 149.800 70.600 150.200 ;
        RECT 64.600 149.100 65.000 149.200 ;
        RECT 57.400 146.800 57.800 147.200 ;
        RECT 58.200 146.800 58.600 147.200 ;
        RECT 54.200 140.800 54.600 141.200 ;
        RECT 51.000 137.800 51.400 138.200 ;
        RECT 51.000 136.800 51.400 137.200 ;
        RECT 51.000 135.200 51.300 136.800 ;
        RECT 48.600 134.800 49.000 135.200 ;
        RECT 49.400 134.800 49.800 135.200 ;
        RECT 51.000 134.800 51.400 135.200 ;
        RECT 48.600 134.200 48.900 134.800 ;
        RECT 47.800 133.800 48.200 134.200 ;
        RECT 48.600 133.800 49.000 134.200 ;
        RECT 46.200 131.800 46.600 132.200 ;
        RECT 47.000 131.800 47.400 132.200 ;
        RECT 44.600 127.800 45.000 128.200 ;
        RECT 44.600 126.100 45.000 126.200 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 44.600 125.800 45.800 126.100 ;
        RECT 44.600 124.800 45.000 125.200 ;
        RECT 45.400 125.100 45.800 125.200 ;
        RECT 46.200 125.100 46.500 131.800 ;
        RECT 47.000 126.200 47.300 131.800 ;
        RECT 47.800 131.200 48.100 133.800 ;
        RECT 47.800 130.800 48.200 131.200 ;
        RECT 47.800 129.200 48.100 130.800 ;
        RECT 47.800 128.800 48.200 129.200 ;
        RECT 47.800 127.800 48.200 128.200 ;
        RECT 47.800 127.200 48.100 127.800 ;
        RECT 48.600 127.200 48.900 133.800 ;
        RECT 47.800 126.800 48.200 127.200 ;
        RECT 48.600 126.800 49.000 127.200 ;
        RECT 47.000 126.100 47.400 126.200 ;
        RECT 47.000 125.800 48.100 126.100 ;
        RECT 45.400 124.800 46.500 125.100 ;
        RECT 43.800 121.800 44.200 122.200 ;
        RECT 40.600 117.800 41.000 118.200 ;
        RECT 40.600 117.200 40.900 117.800 ;
        RECT 37.400 116.800 37.800 117.200 ;
        RECT 40.600 116.800 41.000 117.200 ;
        RECT 37.400 116.200 37.700 116.800 ;
        RECT 35.800 115.800 36.200 116.200 ;
        RECT 37.400 115.800 37.800 116.200 ;
        RECT 42.200 115.800 42.600 116.200 ;
        RECT 35.800 115.200 36.100 115.800 ;
        RECT 35.000 114.800 35.400 115.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 40.600 115.100 41.000 115.200 ;
        RECT 41.400 115.100 41.800 115.200 ;
        RECT 40.600 114.800 41.800 115.100 ;
        RECT 32.600 113.800 33.000 114.200 ;
        RECT 35.000 113.800 35.400 114.200 ;
        RECT 39.800 114.100 40.200 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 39.800 113.800 41.000 114.100 ;
        RECT 32.600 113.200 32.900 113.800 ;
        RECT 35.000 113.200 35.300 113.800 ;
        RECT 31.000 112.800 31.400 113.200 ;
        RECT 32.600 112.800 33.000 113.200 ;
        RECT 35.000 112.800 35.400 113.200 ;
        RECT 37.400 111.800 37.800 112.200 ;
        RECT 29.400 109.800 29.800 110.200 ;
        RECT 29.400 109.200 29.700 109.800 ;
        RECT 29.400 108.800 29.800 109.200 ;
        RECT 31.000 108.100 31.400 108.200 ;
        RECT 31.800 108.100 32.200 108.200 ;
        RECT 31.000 107.800 32.200 108.100 ;
        RECT 31.800 106.800 32.200 107.200 ;
        RECT 31.800 106.200 32.100 106.800 ;
        RECT 31.800 105.800 32.200 106.200 ;
        RECT 35.000 105.100 35.400 107.900 ;
        RECT 36.600 103.100 37.000 108.900 ;
        RECT 37.400 106.300 37.700 111.800 ;
        RECT 40.600 106.800 41.000 107.200 ;
        RECT 37.400 105.900 37.800 106.300 ;
        RECT 40.600 106.200 40.900 106.800 ;
        RECT 37.400 105.800 37.700 105.900 ;
        RECT 40.600 105.800 41.000 106.200 ;
        RECT 41.400 103.100 41.800 108.900 ;
        RECT 42.200 108.200 42.500 115.800 ;
        RECT 43.000 114.800 43.400 115.200 ;
        RECT 43.000 112.200 43.300 114.800 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 42.200 107.800 42.600 108.200 ;
        RECT 43.800 107.100 44.100 121.800 ;
        RECT 44.600 119.200 44.900 124.800 ;
        RECT 47.000 122.800 47.400 123.200 ;
        RECT 44.600 118.800 45.000 119.200 ;
        RECT 46.200 117.800 46.600 118.200 ;
        RECT 46.200 114.200 46.500 117.800 ;
        RECT 47.000 115.200 47.300 122.800 ;
        RECT 47.000 114.800 47.400 115.200 ;
        RECT 46.200 113.800 46.600 114.200 ;
        RECT 47.800 111.200 48.100 125.800 ;
        RECT 48.600 118.200 48.900 126.800 ;
        RECT 49.400 123.200 49.700 134.800 ;
        RECT 51.000 130.200 51.300 134.800 ;
        RECT 51.800 133.100 52.200 135.900 ;
        RECT 53.400 132.100 53.800 137.900 ;
        RECT 51.000 129.800 51.400 130.200 ;
        RECT 53.400 128.800 53.800 129.200 ;
        RECT 53.400 128.200 53.700 128.800 ;
        RECT 53.400 127.800 53.800 128.200 ;
        RECT 50.200 126.800 50.600 127.200 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 49.400 122.800 49.800 123.200 ;
        RECT 49.400 121.800 49.800 122.200 ;
        RECT 48.600 117.800 49.000 118.200 ;
        RECT 48.600 115.800 49.000 116.200 ;
        RECT 48.600 112.200 48.900 115.800 ;
        RECT 49.400 113.100 49.700 121.800 ;
        RECT 50.200 118.200 50.500 126.800 ;
        RECT 51.000 125.100 51.300 126.800 ;
        RECT 54.200 126.200 54.500 140.800 ;
        RECT 57.400 135.200 57.700 146.800 ;
        RECT 59.000 146.100 59.400 146.200 ;
        RECT 59.800 146.100 60.200 146.200 ;
        RECT 59.000 145.800 60.200 146.100 ;
        RECT 61.400 143.100 61.800 148.900 ;
        RECT 63.800 148.800 65.000 149.100 ;
        RECT 64.600 147.200 64.900 148.800 ;
        RECT 70.200 147.800 70.600 148.200 ;
        RECT 70.200 147.200 70.500 147.800 ;
        RECT 64.600 146.800 65.000 147.200 ;
        RECT 69.400 146.800 69.800 147.200 ;
        RECT 70.200 146.800 70.600 147.200 ;
        RECT 69.400 146.200 69.700 146.800 ;
        RECT 75.000 146.200 75.300 152.800 ;
        RECT 75.800 152.100 76.200 157.900 ;
        RECT 76.600 154.200 76.900 166.800 ;
        RECT 77.400 165.100 77.800 167.900 ;
        RECT 78.200 167.200 78.500 173.800 ;
        RECT 79.000 172.100 79.400 177.900 ;
        RECT 82.200 176.800 82.600 177.200 ;
        RECT 82.200 175.200 82.500 176.800 ;
        RECT 82.200 174.800 82.600 175.200 ;
        RECT 83.000 170.200 83.300 193.800 ;
        RECT 83.800 188.200 84.100 201.800 ;
        RECT 84.600 196.200 84.900 205.800 ;
        RECT 89.400 204.200 89.700 206.800 ;
        RECT 90.200 205.800 90.600 206.200 ;
        RECT 90.200 205.200 90.500 205.800 ;
        RECT 90.200 204.800 90.600 205.200 ;
        RECT 91.800 205.100 92.200 207.900 ;
        RECT 92.600 207.800 93.000 208.200 ;
        RECT 92.600 207.200 92.900 207.800 ;
        RECT 92.600 206.800 93.000 207.200 ;
        RECT 86.200 203.800 86.600 204.200 ;
        RECT 89.400 203.800 89.800 204.200 ;
        RECT 86.200 203.200 86.500 203.800 ;
        RECT 86.200 202.800 86.600 203.200 ;
        RECT 93.400 203.100 93.800 208.900 ;
        RECT 97.400 206.800 97.800 207.200 ;
        RECT 94.200 206.200 94.600 206.300 ;
        RECT 95.000 206.200 95.400 206.300 ;
        RECT 94.200 205.900 95.400 206.200 ;
        RECT 97.400 206.200 97.700 206.800 ;
        RECT 97.400 205.800 97.800 206.200 ;
        RECT 95.800 200.800 96.200 201.200 ;
        RECT 87.800 197.800 88.200 198.200 ;
        RECT 87.800 197.200 88.100 197.800 ;
        RECT 86.200 196.800 86.600 197.200 ;
        RECT 87.800 196.800 88.200 197.200 ;
        RECT 86.200 196.200 86.500 196.800 ;
        RECT 84.600 195.800 85.000 196.200 ;
        RECT 86.200 195.800 86.600 196.200 ;
        RECT 87.000 195.800 87.400 196.200 ;
        RECT 90.200 195.800 90.600 196.200 ;
        RECT 91.000 195.800 91.400 196.200 ;
        RECT 84.600 195.100 85.000 195.200 ;
        RECT 85.400 195.100 85.800 195.200 ;
        RECT 84.600 194.800 85.800 195.100 ;
        RECT 87.000 194.200 87.300 195.800 ;
        RECT 87.800 194.800 88.200 195.200 ;
        RECT 85.400 194.100 85.800 194.200 ;
        RECT 86.200 194.100 86.600 194.200 ;
        RECT 85.400 193.800 86.600 194.100 ;
        RECT 87.000 193.800 87.400 194.200 ;
        RECT 87.800 192.200 88.100 194.800 ;
        RECT 87.800 191.800 88.200 192.200 ;
        RECT 83.800 187.800 84.200 188.200 ;
        RECT 83.800 185.900 84.200 186.300 ;
        RECT 83.800 184.200 84.100 185.900 ;
        RECT 83.800 183.800 84.200 184.200 ;
        RECT 84.600 183.100 85.000 188.900 ;
        RECT 86.200 185.100 86.600 187.900 ;
        RECT 90.200 187.200 90.500 195.800 ;
        RECT 91.000 190.200 91.300 195.800 ;
        RECT 91.800 193.100 92.200 195.900 ;
        RECT 93.400 192.100 93.800 197.900 ;
        RECT 94.200 194.700 94.600 195.100 ;
        RECT 94.200 194.200 94.500 194.700 ;
        RECT 94.200 193.800 94.600 194.200 ;
        RECT 91.000 189.800 91.400 190.200 ;
        RECT 90.200 186.800 90.600 187.200 ;
        RECT 91.800 186.800 92.200 187.200 ;
        RECT 94.200 186.800 94.600 187.200 ;
        RECT 91.800 186.200 92.100 186.800 ;
        RECT 94.200 186.200 94.500 186.800 ;
        RECT 95.800 186.200 96.100 200.800 ;
        RECT 97.400 195.200 97.700 205.800 ;
        RECT 98.200 203.100 98.600 208.900 ;
        RECT 101.400 205.100 101.800 207.900 ;
        RECT 102.200 206.800 102.600 207.200 ;
        RECT 102.200 206.200 102.500 206.800 ;
        RECT 102.200 205.800 102.600 206.200 ;
        RECT 99.800 203.100 100.200 203.200 ;
        RECT 100.600 203.100 101.000 203.200 ;
        RECT 103.000 203.100 103.400 208.900 ;
        RECT 104.600 206.100 105.000 206.200 ;
        RECT 105.400 206.100 105.800 206.200 ;
        RECT 104.600 205.800 105.800 206.100 ;
        RECT 107.800 203.100 108.200 208.900 ;
        RECT 116.600 207.800 117.000 208.200 ;
        RECT 120.600 207.800 121.000 208.200 ;
        RECT 116.600 207.200 116.900 207.800 ;
        RECT 120.600 207.200 120.900 207.800 ;
        RECT 111.000 206.800 111.400 207.200 ;
        RECT 116.600 206.800 117.000 207.200 ;
        RECT 117.400 206.800 117.800 207.200 ;
        RECT 120.600 206.800 121.000 207.200 ;
        RECT 110.200 204.800 110.600 205.200 ;
        RECT 110.200 204.200 110.500 204.800 ;
        RECT 111.000 204.200 111.300 206.800 ;
        RECT 111.800 205.800 112.200 206.200 ;
        RECT 112.600 206.100 113.000 206.200 ;
        RECT 113.400 206.100 113.800 206.200 ;
        RECT 112.600 205.800 113.800 206.100 ;
        RECT 115.800 205.800 116.200 206.200 ;
        RECT 108.600 203.800 109.000 204.200 ;
        RECT 110.200 203.800 110.600 204.200 ;
        RECT 111.000 203.800 111.400 204.200 ;
        RECT 99.800 202.800 101.000 203.100 ;
        RECT 97.400 194.800 97.800 195.200 ;
        RECT 98.200 192.100 98.600 197.900 ;
        RECT 99.800 191.200 100.100 202.800 ;
        RECT 108.600 201.200 108.900 203.800 ;
        RECT 108.600 200.800 109.000 201.200 ;
        RECT 103.800 196.800 104.200 197.200 ;
        RECT 105.400 197.100 105.800 197.200 ;
        RECT 106.200 197.100 106.600 197.200 ;
        RECT 105.400 196.800 106.600 197.100 ;
        RECT 103.800 196.200 104.100 196.800 ;
        RECT 102.200 195.800 102.600 196.200 ;
        RECT 103.800 195.800 104.200 196.200 ;
        RECT 107.000 195.800 107.400 196.200 ;
        RECT 102.200 195.200 102.500 195.800 ;
        RECT 102.200 194.800 102.600 195.200 ;
        RECT 105.400 194.800 105.800 195.200 ;
        RECT 101.400 194.100 101.800 194.200 ;
        RECT 102.200 194.100 102.600 194.200 ;
        RECT 101.400 193.800 102.600 194.100 ;
        RECT 103.800 193.800 104.200 194.200 ;
        RECT 104.600 193.800 105.000 194.200 ;
        RECT 103.800 193.200 104.100 193.800 ;
        RECT 104.600 193.200 104.900 193.800 ;
        RECT 103.800 192.800 104.200 193.200 ;
        RECT 104.600 192.800 105.000 193.200 ;
        RECT 105.400 192.200 105.700 194.800 ;
        RECT 107.000 192.200 107.300 195.800 ;
        RECT 107.800 193.100 108.200 195.900 ;
        RECT 108.600 194.200 108.900 200.800 ;
        RECT 108.600 193.800 109.000 194.200 ;
        RECT 100.600 191.800 101.000 192.200 ;
        RECT 105.400 191.800 105.800 192.200 ;
        RECT 107.000 191.800 107.400 192.200 ;
        RECT 109.400 192.100 109.800 197.900 ;
        RECT 110.200 194.700 110.600 195.100 ;
        RECT 110.200 194.200 110.500 194.700 ;
        RECT 110.200 193.800 110.600 194.200 ;
        RECT 98.200 190.800 98.600 191.200 ;
        RECT 99.800 190.800 100.200 191.200 ;
        RECT 98.200 186.200 98.500 190.800 ;
        RECT 100.600 190.200 100.900 191.800 ;
        RECT 100.600 189.800 101.000 190.200 ;
        RECT 104.600 189.800 105.000 190.200 ;
        RECT 103.800 187.800 104.200 188.200 ;
        RECT 99.000 186.800 99.400 187.200 ;
        RECT 99.000 186.200 99.300 186.800 ;
        RECT 87.000 185.800 87.400 186.200 ;
        RECT 89.400 185.800 89.800 186.200 ;
        RECT 91.800 185.800 92.200 186.200 ;
        RECT 93.400 185.800 93.800 186.200 ;
        RECT 94.200 185.800 94.600 186.200 ;
        RECT 95.000 185.800 95.400 186.200 ;
        RECT 95.800 185.800 96.200 186.200 ;
        RECT 98.200 185.800 98.600 186.200 ;
        RECT 99.000 185.800 99.400 186.200 ;
        RECT 99.800 185.800 100.200 186.200 ;
        RECT 100.600 186.100 101.000 186.200 ;
        RECT 101.400 186.100 101.800 186.200 ;
        RECT 100.600 185.800 101.800 186.100 ;
        RECT 87.000 185.200 87.300 185.800 ;
        RECT 87.000 184.800 87.400 185.200 ;
        RECT 88.600 183.800 89.000 184.200 ;
        RECT 88.600 183.200 88.900 183.800 ;
        RECT 88.600 182.800 89.000 183.200 ;
        RECT 87.000 180.800 87.400 181.200 ;
        RECT 83.800 172.100 84.200 177.900 ;
        RECT 86.200 176.800 86.600 177.200 ;
        RECT 86.200 176.200 86.500 176.800 ;
        RECT 86.200 175.800 86.600 176.200 ;
        RECT 87.000 174.200 87.300 180.800 ;
        RECT 88.600 176.800 89.000 177.200 ;
        RECT 88.600 175.200 88.900 176.800 ;
        RECT 87.800 174.800 88.200 175.200 ;
        RECT 88.600 174.800 89.000 175.200 ;
        RECT 87.800 174.200 88.100 174.800 ;
        RECT 89.400 174.200 89.700 185.800 ;
        RECT 91.800 184.800 92.200 185.200 ;
        RECT 91.800 184.200 92.100 184.800 ;
        RECT 91.800 183.800 92.200 184.200 ;
        RECT 93.400 180.200 93.700 185.800 ;
        RECT 95.000 184.200 95.300 185.800 ;
        RECT 95.000 183.800 95.400 184.200 ;
        RECT 93.400 179.800 93.800 180.200 ;
        RECT 97.400 179.100 97.800 179.200 ;
        RECT 98.200 179.100 98.600 179.200 ;
        RECT 97.400 178.800 98.600 179.100 ;
        RECT 99.800 178.200 100.100 185.800 ;
        RECT 101.400 183.100 101.800 183.200 ;
        RECT 102.200 183.100 102.600 183.200 ;
        RECT 101.400 182.800 102.600 183.100 ;
        RECT 99.800 177.800 100.200 178.200 ;
        RECT 91.800 176.100 92.200 176.200 ;
        RECT 92.600 176.100 93.000 176.200 ;
        RECT 91.800 175.800 93.000 176.100 ;
        RECT 95.800 175.800 96.200 176.200 ;
        RECT 100.600 176.100 101.000 176.200 ;
        RECT 100.600 175.800 101.700 176.100 ;
        RECT 93.400 174.800 93.800 175.200 ;
        RECT 93.400 174.200 93.700 174.800 ;
        RECT 87.000 173.800 87.400 174.200 ;
        RECT 87.800 173.800 88.200 174.200 ;
        RECT 89.400 173.800 89.800 174.200 ;
        RECT 93.400 173.800 93.800 174.200 ;
        RECT 94.200 173.800 94.600 174.200 ;
        RECT 87.000 172.200 87.300 173.800 ;
        RECT 87.000 171.800 87.400 172.200 ;
        RECT 83.000 169.800 83.400 170.200 ;
        RECT 93.400 169.800 93.800 170.200 ;
        RECT 85.400 169.100 85.800 169.200 ;
        RECT 86.200 169.100 86.600 169.200 ;
        RECT 78.200 166.800 78.600 167.200 ;
        RECT 78.200 158.200 78.500 166.800 ;
        RECT 79.000 163.100 79.400 168.900 ;
        RECT 79.800 166.100 80.200 166.300 ;
        RECT 80.600 166.100 81.000 166.200 ;
        RECT 79.800 165.800 81.000 166.100 ;
        RECT 83.000 163.800 83.400 164.200 ;
        RECT 83.000 159.200 83.300 163.800 ;
        RECT 83.800 163.100 84.200 168.900 ;
        RECT 85.400 168.800 86.600 169.100 ;
        RECT 91.000 166.800 91.400 167.200 ;
        RECT 91.000 166.200 91.300 166.800 ;
        RECT 93.400 166.200 93.700 169.800 ;
        RECT 94.200 167.200 94.500 173.800 ;
        RECT 94.200 167.100 94.600 167.200 ;
        RECT 95.000 167.100 95.400 167.200 ;
        RECT 94.200 166.800 95.400 167.100 ;
        RECT 95.800 166.200 96.100 175.800 ;
        RECT 100.600 174.800 101.000 175.200 ;
        RECT 100.600 174.200 100.900 174.800 ;
        RECT 101.400 174.200 101.700 175.800 ;
        RECT 103.800 174.200 104.100 187.800 ;
        RECT 104.600 186.200 104.900 189.800 ;
        RECT 104.600 185.800 105.000 186.200 ;
        RECT 105.400 185.100 105.700 191.800 ;
        RECT 109.400 188.100 109.800 188.200 ;
        RECT 110.200 188.100 110.600 188.200 ;
        RECT 109.400 187.800 110.600 188.100 ;
        RECT 111.000 187.100 111.300 203.800 ;
        RECT 111.800 198.200 112.100 205.800 ;
        RECT 115.800 205.200 116.100 205.800 ;
        RECT 114.200 204.800 114.600 205.200 ;
        RECT 115.800 204.800 116.200 205.200 ;
        RECT 114.200 204.200 114.500 204.800 ;
        RECT 114.200 203.800 114.600 204.200 ;
        RECT 114.200 200.200 114.500 203.800 ;
        RECT 114.200 199.800 114.600 200.200 ;
        RECT 111.800 197.800 112.200 198.200 ;
        RECT 114.200 192.100 114.600 197.900 ;
        RECT 115.800 193.200 116.100 204.800 ;
        RECT 116.600 194.200 116.900 206.800 ;
        RECT 117.400 206.200 117.700 206.800 ;
        RECT 117.400 205.800 117.800 206.200 ;
        RECT 118.200 205.800 118.600 206.200 ;
        RECT 119.800 206.100 120.200 206.200 ;
        RECT 120.600 206.100 121.000 206.200 ;
        RECT 119.800 205.800 121.000 206.100 ;
        RECT 121.400 205.800 121.800 206.200 ;
        RECT 116.600 193.800 117.000 194.200 ;
        RECT 115.800 192.800 116.200 193.200 ;
        RECT 117.400 193.100 117.800 195.900 ;
        RECT 118.200 194.200 118.500 205.800 ;
        RECT 121.400 205.200 121.700 205.800 ;
        RECT 119.800 204.800 120.200 205.200 ;
        RECT 121.400 204.800 121.800 205.200 ;
        RECT 123.000 204.800 123.400 205.200 ;
        RECT 123.800 205.100 124.200 207.900 ;
        RECT 124.600 206.800 125.000 207.200 ;
        RECT 119.800 204.200 120.100 204.800 ;
        RECT 123.000 204.200 123.300 204.800 ;
        RECT 119.800 203.800 120.200 204.200 ;
        RECT 121.400 203.800 121.800 204.200 ;
        RECT 123.000 203.800 123.400 204.200 ;
        RECT 121.400 203.200 121.700 203.800 ;
        RECT 121.400 202.800 121.800 203.200 ;
        RECT 124.600 201.200 124.900 206.800 ;
        RECT 125.400 203.100 125.800 208.900 ;
        RECT 129.400 207.800 129.800 208.200 ;
        RECT 129.400 207.200 129.700 207.800 ;
        RECT 126.200 206.800 126.600 207.200 ;
        RECT 129.400 206.800 129.800 207.200 ;
        RECT 126.200 206.300 126.500 206.800 ;
        RECT 126.200 205.900 126.600 206.300 ;
        RECT 130.200 203.100 130.600 208.900 ;
        RECT 142.200 205.100 142.600 207.900 ;
        RECT 143.000 206.800 143.400 207.200 ;
        RECT 143.000 206.200 143.300 206.800 ;
        RECT 143.000 205.800 143.400 206.200 ;
        RECT 131.800 204.100 132.200 204.200 ;
        RECT 132.600 204.100 133.000 204.200 ;
        RECT 131.800 203.800 133.000 204.100 ;
        RECT 133.400 203.800 133.800 204.200 ;
        RECT 124.600 200.800 125.000 201.200 ;
        RECT 128.600 200.800 129.000 201.200 ;
        RECT 118.200 193.800 118.600 194.200 ;
        RECT 115.800 191.200 116.100 192.800 ;
        RECT 116.600 192.100 117.000 192.200 ;
        RECT 116.600 191.800 117.700 192.100 ;
        RECT 114.200 190.800 114.600 191.200 ;
        RECT 115.800 190.800 116.200 191.200 ;
        RECT 114.200 189.200 114.500 190.800 ;
        RECT 114.200 188.800 114.600 189.200 ;
        RECT 110.200 186.800 111.300 187.100 ;
        RECT 115.800 187.800 116.200 188.200 ;
        RECT 115.800 187.200 116.100 187.800 ;
        RECT 115.800 186.800 116.200 187.200 ;
        RECT 104.600 184.800 105.700 185.100 ;
        RECT 107.800 185.800 108.200 186.200 ;
        RECT 108.600 185.800 109.000 186.200 ;
        RECT 107.800 185.200 108.100 185.800 ;
        RECT 107.800 184.800 108.200 185.200 ;
        RECT 104.600 175.200 104.900 184.800 ;
        RECT 108.600 182.200 108.900 185.800 ;
        RECT 108.600 181.800 109.000 182.200 ;
        RECT 107.000 177.800 107.400 178.200 ;
        RECT 108.600 177.800 109.000 178.200 ;
        RECT 106.200 175.800 106.600 176.200 ;
        RECT 104.600 174.800 105.000 175.200 ;
        RECT 99.000 173.800 99.400 174.200 ;
        RECT 100.600 173.800 101.000 174.200 ;
        RECT 101.400 173.800 101.800 174.200 ;
        RECT 103.800 173.800 104.200 174.200 ;
        RECT 87.000 165.800 87.400 166.200 ;
        RECT 89.400 165.800 89.800 166.200 ;
        RECT 91.000 165.800 91.400 166.200 ;
        RECT 92.600 166.100 93.000 166.200 ;
        RECT 93.400 166.100 93.800 166.200 ;
        RECT 92.600 165.800 93.800 166.100 ;
        RECT 95.000 165.800 95.400 166.200 ;
        RECT 95.800 165.800 96.200 166.200 ;
        RECT 97.400 165.800 97.800 166.200 ;
        RECT 98.200 165.800 98.600 166.200 ;
        RECT 83.000 158.800 83.400 159.200 ;
        RECT 78.200 157.800 78.600 158.200 ;
        RECT 79.000 155.800 79.400 156.200 ;
        RECT 79.000 155.200 79.300 155.800 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 76.600 153.800 77.000 154.200 ;
        RECT 79.800 153.800 80.200 154.200 ;
        RECT 79.800 153.200 80.100 153.800 ;
        RECT 79.800 152.800 80.200 153.200 ;
        RECT 80.600 152.100 81.000 157.900 ;
        RECT 85.400 155.800 85.800 156.200 ;
        RECT 86.200 155.800 86.600 156.200 ;
        RECT 85.400 155.200 85.700 155.800 ;
        RECT 86.200 155.200 86.500 155.800 ;
        RECT 83.800 155.100 84.200 155.200 ;
        RECT 84.600 155.100 85.000 155.200 ;
        RECT 83.800 154.800 85.000 155.100 ;
        RECT 85.400 154.800 85.800 155.200 ;
        RECT 86.200 154.800 86.600 155.200 ;
        RECT 83.800 154.100 84.200 154.200 ;
        RECT 84.600 154.100 85.000 154.200 ;
        RECT 83.800 153.800 85.000 154.100 ;
        RECT 87.000 152.200 87.300 165.800 ;
        RECT 89.400 156.200 89.700 165.800 ;
        RECT 91.800 164.800 92.200 165.200 ;
        RECT 91.800 164.200 92.100 164.800 ;
        RECT 91.800 163.800 92.200 164.200 ;
        RECT 95.000 161.200 95.300 165.800 ;
        RECT 97.400 165.200 97.700 165.800 ;
        RECT 97.400 164.800 97.800 165.200 ;
        RECT 98.200 164.200 98.500 165.800 ;
        RECT 98.200 163.800 98.600 164.200 ;
        RECT 97.400 161.800 97.800 162.200 ;
        RECT 95.000 160.800 95.400 161.200 ;
        RECT 97.400 159.200 97.700 161.800 ;
        RECT 97.400 158.800 97.800 159.200 ;
        RECT 99.000 158.200 99.300 173.800 ;
        RECT 101.400 173.200 101.700 173.800 ;
        RECT 103.800 173.200 104.100 173.800 ;
        RECT 101.400 172.800 101.800 173.200 ;
        RECT 103.800 172.800 104.200 173.200 ;
        RECT 102.200 171.800 102.600 172.200 ;
        RECT 103.000 171.800 103.400 172.200 ;
        RECT 102.200 171.200 102.500 171.800 ;
        RECT 102.200 170.800 102.600 171.200 ;
        RECT 99.800 167.100 100.200 167.200 ;
        RECT 100.600 167.100 101.000 167.200 ;
        RECT 99.800 166.800 101.000 167.100 ;
        RECT 99.800 166.100 100.200 166.200 ;
        RECT 100.600 166.100 101.000 166.200 ;
        RECT 102.200 166.100 102.600 166.200 ;
        RECT 99.800 165.800 101.000 166.100 ;
        RECT 101.400 165.800 102.600 166.100 ;
        RECT 99.800 161.800 100.200 162.200 ;
        RECT 100.600 161.800 101.000 162.200 ;
        RECT 88.600 153.100 89.000 155.900 ;
        RECT 89.400 155.800 89.800 156.200 ;
        RECT 89.400 153.800 89.800 154.200 ;
        RECT 89.400 153.200 89.700 153.800 ;
        RECT 89.400 152.800 89.800 153.200 ;
        RECT 84.600 151.800 85.000 152.200 ;
        RECT 87.000 151.800 87.400 152.200 ;
        RECT 90.200 152.100 90.600 157.900 ;
        RECT 92.600 155.100 93.000 155.200 ;
        RECT 93.400 155.100 93.800 155.200 ;
        RECT 92.600 154.800 93.800 155.100 ;
        RECT 94.200 152.800 94.600 153.200 ;
        RECT 91.000 151.800 91.400 152.200 ;
        RECT 84.600 149.200 84.900 151.800 ;
        RECT 91.000 149.200 91.300 151.800 ;
        RECT 84.600 148.800 85.000 149.200 ;
        RECT 91.000 148.800 91.400 149.200 ;
        RECT 77.400 147.800 77.800 148.200 ;
        RECT 80.600 148.100 81.000 148.200 ;
        RECT 81.400 148.100 81.800 148.200 ;
        RECT 80.600 147.800 81.800 148.100 ;
        RECT 77.400 147.200 77.700 147.800 ;
        RECT 77.400 146.800 77.800 147.200 ;
        RECT 78.200 146.800 78.600 147.200 ;
        RECT 79.000 146.800 79.400 147.200 ;
        RECT 82.200 146.800 82.600 147.200 ;
        RECT 87.000 146.800 87.400 147.200 ;
        RECT 78.200 146.200 78.500 146.800 ;
        RECT 79.000 146.200 79.300 146.800 ;
        RECT 65.400 145.800 65.800 146.200 ;
        RECT 66.200 146.100 66.600 146.200 ;
        RECT 67.000 146.100 67.400 146.200 ;
        RECT 66.200 145.800 67.400 146.100 ;
        RECT 69.400 145.800 69.800 146.200 ;
        RECT 74.200 145.800 74.600 146.200 ;
        RECT 75.000 145.800 75.400 146.200 ;
        RECT 78.200 145.800 78.600 146.200 ;
        RECT 79.000 145.800 79.400 146.200 ;
        RECT 80.600 145.800 81.000 146.200 ;
        RECT 63.800 144.100 64.200 144.200 ;
        RECT 64.600 144.100 65.000 144.200 ;
        RECT 63.800 143.800 65.000 144.100 ;
        RECT 65.400 143.200 65.700 145.800 ;
        RECT 67.800 144.800 68.200 145.200 ;
        RECT 73.400 145.100 73.800 145.200 ;
        RECT 72.600 144.800 73.800 145.100 ;
        RECT 67.800 144.200 68.100 144.800 ;
        RECT 67.800 143.800 68.200 144.200 ;
        RECT 65.400 142.800 65.800 143.200 ;
        RECT 71.800 141.800 72.200 142.200 ;
        RECT 55.000 134.800 55.400 135.200 ;
        RECT 57.400 134.800 57.800 135.200 ;
        RECT 55.000 129.200 55.300 134.800 ;
        RECT 57.400 134.200 57.700 134.800 ;
        RECT 57.400 133.800 57.800 134.200 ;
        RECT 56.600 131.800 57.000 132.200 ;
        RECT 58.200 132.100 58.600 137.900 ;
        RECT 61.400 136.100 61.800 136.200 ;
        RECT 62.200 136.100 62.600 136.200 ;
        RECT 61.400 135.800 62.600 136.100 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 63.000 135.200 63.300 135.800 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 61.400 133.800 61.800 134.200 ;
        RECT 59.800 132.100 60.200 132.200 ;
        RECT 60.600 132.100 61.000 132.200 ;
        RECT 59.800 131.800 61.000 132.100 ;
        RECT 55.000 128.800 55.400 129.200 ;
        RECT 56.600 128.200 56.900 131.800 ;
        RECT 61.400 131.200 61.700 133.800 ;
        RECT 63.800 133.100 64.200 135.900 ;
        RECT 64.600 134.800 65.000 135.200 ;
        RECT 64.600 134.200 64.900 134.800 ;
        RECT 64.600 133.800 65.000 134.200 ;
        RECT 65.400 132.100 65.800 137.900 ;
        RECT 67.800 135.100 68.200 135.200 ;
        RECT 68.600 135.100 69.000 135.200 ;
        RECT 67.800 134.800 69.000 135.100 ;
        RECT 70.200 132.100 70.600 137.900 ;
        RECT 71.800 136.200 72.100 141.800 ;
        RECT 72.600 139.200 72.900 144.800 ;
        RECT 74.200 144.200 74.500 145.800 ;
        RECT 74.200 143.800 74.600 144.200 ;
        RECT 75.000 142.800 75.400 143.200 ;
        RECT 72.600 138.800 73.000 139.200 ;
        RECT 71.800 135.800 72.200 136.200 ;
        RECT 72.600 136.100 73.000 136.200 ;
        RECT 73.400 136.100 73.800 136.200 ;
        RECT 72.600 135.800 73.800 136.100 ;
        RECT 75.000 135.200 75.300 142.800 ;
        RECT 75.800 141.800 76.200 142.200 ;
        RECT 72.600 135.100 73.000 135.200 ;
        RECT 73.400 135.100 73.800 135.200 ;
        RECT 72.600 134.800 73.800 135.100 ;
        RECT 75.000 134.800 75.400 135.200 ;
        RECT 75.000 134.200 75.300 134.800 ;
        RECT 75.800 134.200 76.100 141.800 ;
        RECT 76.600 139.800 77.000 140.200 ;
        RECT 79.000 139.800 79.400 140.200 ;
        RECT 76.600 136.200 76.900 139.800 ;
        RECT 79.000 136.200 79.300 139.800 ;
        RECT 80.600 137.200 80.900 145.800 ;
        RECT 82.200 142.200 82.500 146.800 ;
        RECT 87.000 146.200 87.300 146.800 ;
        RECT 85.400 146.100 85.800 146.200 ;
        RECT 86.200 146.100 86.600 146.200 ;
        RECT 85.400 145.800 86.600 146.100 ;
        RECT 87.000 145.800 87.400 146.200 ;
        RECT 91.000 145.800 91.400 146.200 ;
        RECT 93.400 145.800 93.800 146.200 ;
        RECT 91.000 145.200 91.300 145.800 ;
        RECT 93.400 145.200 93.700 145.800 ;
        RECT 83.800 145.100 84.200 145.200 ;
        RECT 84.600 145.100 85.000 145.200 ;
        RECT 83.800 144.800 85.000 145.100 ;
        RECT 91.000 144.800 91.400 145.200 ;
        RECT 92.600 144.800 93.000 145.200 ;
        RECT 93.400 144.800 93.800 145.200 ;
        RECT 83.800 143.800 84.200 144.200 ;
        RECT 91.800 143.800 92.200 144.200 ;
        RECT 83.800 143.200 84.100 143.800 ;
        RECT 83.800 142.800 84.200 143.200 ;
        RECT 82.200 141.800 82.600 142.200 ;
        RECT 91.000 141.800 91.400 142.200 ;
        RECT 80.600 137.100 81.000 137.200 ;
        RECT 81.400 137.100 81.800 137.200 ;
        RECT 80.600 136.800 81.800 137.100 ;
        RECT 76.600 135.800 77.000 136.200 ;
        RECT 79.000 135.800 79.400 136.200 ;
        RECT 84.600 136.100 85.000 136.200 ;
        RECT 85.400 136.100 85.800 136.200 ;
        RECT 84.600 135.800 85.800 136.100 ;
        RECT 78.200 134.800 78.600 135.200 ;
        RECT 79.800 135.100 80.200 135.200 ;
        RECT 80.600 135.100 81.000 135.200 ;
        RECT 79.800 134.800 81.000 135.100 ;
        RECT 83.000 134.800 83.400 135.200 ;
        RECT 83.800 135.100 84.200 135.200 ;
        RECT 84.600 135.100 85.000 135.200 ;
        RECT 83.800 134.800 85.000 135.100 ;
        RECT 78.200 134.200 78.500 134.800 ;
        RECT 83.000 134.200 83.300 134.800 ;
        RECT 75.000 133.800 75.400 134.200 ;
        RECT 75.800 133.800 76.200 134.200 ;
        RECT 78.200 133.800 78.600 134.200 ;
        RECT 79.800 133.800 80.200 134.200 ;
        RECT 82.200 133.800 82.600 134.200 ;
        RECT 83.000 133.800 83.400 134.200 ;
        RECT 79.800 133.200 80.100 133.800 ;
        RECT 82.200 133.200 82.500 133.800 ;
        RECT 78.200 132.800 78.600 133.200 ;
        RECT 79.800 132.800 80.200 133.200 ;
        RECT 82.200 132.800 82.600 133.200 ;
        RECT 87.000 133.100 87.400 135.900 ;
        RECT 87.800 133.800 88.200 134.200 ;
        RECT 72.600 132.100 73.000 132.200 ;
        RECT 73.400 132.100 73.800 132.200 ;
        RECT 72.600 131.800 73.800 132.100 ;
        RECT 75.000 131.800 75.400 132.200 ;
        RECT 76.600 131.800 77.000 132.200 ;
        RECT 61.400 130.800 61.800 131.200 ;
        RECT 66.200 129.800 66.600 130.200 ;
        RECT 56.600 127.800 57.000 128.200 ;
        RECT 63.000 128.100 63.400 128.200 ;
        RECT 63.800 128.100 64.200 128.200 ;
        RECT 63.000 127.800 64.200 128.100 ;
        RECT 63.000 127.100 63.400 127.200 ;
        RECT 63.800 127.100 64.200 127.200 ;
        RECT 63.000 126.800 64.200 127.100 ;
        RECT 51.800 126.100 52.200 126.200 ;
        RECT 52.600 126.100 53.000 126.200 ;
        RECT 51.800 125.800 53.000 126.100 ;
        RECT 54.200 125.800 54.600 126.200 ;
        RECT 55.800 125.800 56.200 126.200 ;
        RECT 59.000 126.100 59.400 126.200 ;
        RECT 59.800 126.100 60.200 126.200 ;
        RECT 59.000 125.800 60.200 126.100 ;
        RECT 54.200 125.200 54.500 125.800 ;
        RECT 51.000 124.800 52.100 125.100 ;
        RECT 50.200 117.800 50.600 118.200 ;
        RECT 51.000 115.800 51.400 116.200 ;
        RECT 51.000 115.200 51.300 115.800 ;
        RECT 50.200 114.800 50.600 115.200 ;
        RECT 51.000 114.800 51.400 115.200 ;
        RECT 50.200 114.200 50.500 114.800 ;
        RECT 51.800 114.200 52.100 124.800 ;
        RECT 54.200 124.800 54.600 125.200 ;
        RECT 50.200 113.800 50.600 114.200 ;
        RECT 51.800 113.800 52.200 114.200 ;
        RECT 49.400 112.800 50.500 113.100 ;
        RECT 48.600 111.800 49.000 112.200 ;
        RECT 47.800 110.800 48.200 111.200 ;
        RECT 43.000 106.800 44.100 107.100 ;
        RECT 33.400 101.800 33.800 102.200 ;
        RECT 28.600 98.800 29.000 99.200 ;
        RECT 33.400 98.200 33.700 101.800 ;
        RECT 34.200 100.800 34.600 101.200 ;
        RECT 39.800 100.800 40.200 101.200 ;
        RECT 27.800 92.100 28.200 97.900 ;
        RECT 33.400 97.800 33.800 98.200 ;
        RECT 29.400 97.100 29.800 97.200 ;
        RECT 30.200 97.100 30.600 97.200 ;
        RECT 29.400 96.800 30.600 97.100 ;
        RECT 32.600 97.100 33.000 97.200 ;
        RECT 33.400 97.100 33.800 97.200 ;
        RECT 32.600 96.800 33.800 97.100 ;
        RECT 30.200 94.200 30.500 96.800 ;
        RECT 34.200 96.200 34.500 100.800 ;
        RECT 34.200 96.100 34.600 96.200 ;
        RECT 35.000 96.100 35.400 96.200 ;
        RECT 34.200 95.800 35.400 96.100 ;
        RECT 39.000 94.800 39.400 95.200 ;
        RECT 30.200 93.800 30.600 94.200 ;
        RECT 31.800 94.100 32.200 94.200 ;
        RECT 32.600 94.100 33.000 94.200 ;
        RECT 31.800 93.800 33.000 94.100 ;
        RECT 31.000 92.800 31.400 93.200 ;
        RECT 31.800 93.100 32.200 93.200 ;
        RECT 32.600 93.100 33.000 93.200 ;
        RECT 31.800 92.800 33.000 93.100 ;
        RECT 35.000 92.800 35.400 93.200 ;
        RECT 31.000 90.200 31.300 92.800 ;
        RECT 27.000 89.800 28.100 90.100 ;
        RECT 31.000 89.800 31.400 90.200 ;
        RECT 26.200 87.800 26.600 88.200 ;
        RECT 27.000 87.800 27.400 88.200 ;
        RECT 26.200 87.200 26.500 87.800 ;
        RECT 26.200 86.800 26.600 87.200 ;
        RECT 27.000 86.200 27.300 87.800 ;
        RECT 25.400 86.100 25.800 86.200 ;
        RECT 26.200 86.100 26.600 86.200 ;
        RECT 25.400 85.800 26.600 86.100 ;
        RECT 27.000 85.800 27.400 86.200 ;
        RECT 25.400 85.100 25.800 85.200 ;
        RECT 26.200 85.100 26.600 85.200 ;
        RECT 25.400 84.800 26.600 85.100 ;
        RECT 27.000 84.800 27.400 85.200 ;
        RECT 27.000 84.200 27.300 84.800 ;
        RECT 27.800 84.200 28.100 89.800 ;
        RECT 28.600 88.800 29.000 89.200 ;
        RECT 28.600 85.200 28.900 88.800 ;
        RECT 28.600 84.800 29.000 85.200 ;
        RECT 29.400 85.100 29.800 87.900 ;
        RECT 30.200 86.800 30.600 87.200 ;
        RECT 27.000 83.800 27.400 84.200 ;
        RECT 27.800 83.800 28.200 84.200 ;
        RECT 30.200 83.200 30.500 86.800 ;
        RECT 24.600 82.800 25.000 83.200 ;
        RECT 27.000 82.800 27.400 83.200 ;
        RECT 30.200 82.800 30.600 83.200 ;
        RECT 31.000 83.100 31.400 88.900 ;
        RECT 31.800 86.200 32.200 86.300 ;
        RECT 32.600 86.200 33.000 86.300 ;
        RECT 31.800 85.900 33.000 86.200 ;
        RECT 21.400 81.800 21.800 82.200 ;
        RECT 20.600 78.800 21.000 79.200 ;
        RECT 20.600 74.200 20.900 78.800 ;
        RECT 21.400 77.200 21.700 81.800 ;
        RECT 21.400 76.800 21.800 77.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 21.400 73.100 21.800 75.900 ;
        RECT 23.000 72.100 23.400 77.900 ;
        RECT 25.400 76.800 25.800 77.200 ;
        RECT 24.600 75.100 25.000 75.200 ;
        RECT 23.800 74.800 25.000 75.100 ;
        RECT 23.800 74.700 24.200 74.800 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 21.400 66.200 21.700 66.800 ;
        RECT 19.800 65.800 20.200 66.200 ;
        RECT 21.400 65.800 21.800 66.200 ;
        RECT 17.400 64.800 17.800 65.200 ;
        RECT 16.600 59.800 17.000 60.200 ;
        RECT 16.600 57.800 17.000 58.200 ;
        RECT 16.600 57.200 16.900 57.800 ;
        RECT 16.600 56.800 17.000 57.200 ;
        RECT 15.000 55.800 16.100 56.100 ;
        RECT 15.000 55.200 15.300 55.800 ;
        RECT 15.000 54.800 15.400 55.200 ;
        RECT 15.800 55.100 16.200 55.200 ;
        RECT 16.600 55.100 17.000 55.200 ;
        RECT 15.800 54.800 17.000 55.100 ;
        RECT 13.400 53.800 13.800 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 15.800 54.100 16.200 54.200 ;
        RECT 15.000 53.800 16.200 54.100 ;
        RECT 15.000 50.800 15.400 51.200 ;
        RECT 12.600 48.800 13.000 49.200 ;
        RECT 12.600 48.200 12.900 48.800 ;
        RECT 12.600 47.800 13.000 48.200 ;
        RECT 15.000 47.200 15.300 50.800 ;
        RECT 17.400 49.200 17.700 64.800 ;
        RECT 19.000 56.800 19.400 57.200 ;
        RECT 19.000 56.200 19.300 56.800 ;
        RECT 19.000 55.800 19.400 56.200 ;
        RECT 19.000 55.200 19.300 55.800 ;
        RECT 19.000 54.800 19.400 55.200 ;
        RECT 19.800 53.200 20.100 65.800 ;
        RECT 20.600 65.100 21.000 65.200 ;
        RECT 21.400 65.100 21.800 65.200 ;
        RECT 22.200 65.100 22.600 67.900 ;
        RECT 20.600 64.800 21.800 65.100 ;
        RECT 23.800 63.100 24.200 68.900 ;
        RECT 25.400 66.200 25.700 76.800 ;
        RECT 27.000 75.200 27.300 82.800 ;
        RECT 35.000 79.200 35.300 92.800 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 38.200 89.100 38.600 89.200 ;
        RECT 35.800 83.100 36.200 88.900 ;
        RECT 37.400 88.800 38.600 89.100 ;
        RECT 39.000 85.200 39.300 94.800 ;
        RECT 39.800 88.200 40.100 100.800 ;
        RECT 40.600 96.800 41.000 97.200 ;
        RECT 40.600 96.200 40.900 96.800 ;
        RECT 40.600 95.800 41.000 96.200 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 41.400 94.200 41.700 94.800 ;
        RECT 41.400 93.800 41.800 94.200 ;
        RECT 41.400 92.800 41.800 93.200 ;
        RECT 40.600 91.800 41.000 92.200 ;
        RECT 39.800 87.800 40.200 88.200 ;
        RECT 40.600 87.200 40.900 91.800 ;
        RECT 41.400 89.200 41.700 92.800 ;
        RECT 43.000 89.200 43.300 106.800 ;
        RECT 43.800 106.100 44.200 106.200 ;
        RECT 44.600 106.100 45.000 106.200 ;
        RECT 43.800 105.800 45.000 106.100 ;
        RECT 47.800 105.100 48.200 107.900 ;
        RECT 48.600 106.800 49.000 107.200 ;
        RECT 43.800 101.800 44.200 102.200 ;
        RECT 46.200 102.100 46.600 102.200 ;
        RECT 47.000 102.100 47.400 102.200 ;
        RECT 46.200 101.800 47.400 102.100 ;
        RECT 43.800 100.200 44.100 101.800 ;
        RECT 43.800 99.800 44.200 100.200 ;
        RECT 43.800 98.800 44.200 99.200 ;
        RECT 43.800 95.200 44.100 98.800 ;
        RECT 44.600 97.800 45.000 98.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 44.600 95.100 44.900 97.800 ;
        RECT 45.400 96.100 45.800 96.200 ;
        RECT 45.400 95.800 48.100 96.100 ;
        RECT 47.800 95.200 48.100 95.800 ;
        RECT 45.400 95.100 45.800 95.200 ;
        RECT 44.600 94.800 45.800 95.100 ;
        RECT 47.000 94.800 47.400 95.200 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 43.800 90.200 44.100 94.800 ;
        RECT 47.000 94.200 47.300 94.800 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 47.000 93.800 47.400 94.200 ;
        RECT 46.200 91.200 46.500 93.800 ;
        RECT 46.200 90.800 46.600 91.200 ;
        RECT 43.800 89.800 44.200 90.200 ;
        RECT 41.400 88.800 41.800 89.200 ;
        RECT 43.000 88.800 43.400 89.200 ;
        RECT 42.200 87.800 42.600 88.200 ;
        RECT 42.200 87.200 42.500 87.800 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 42.200 86.800 42.600 87.200 ;
        RECT 39.000 84.800 39.400 85.200 ;
        RECT 42.200 84.800 42.600 85.200 ;
        RECT 43.000 85.100 43.400 87.900 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 42.200 82.200 42.500 84.800 ;
        RECT 43.800 83.200 44.100 86.800 ;
        RECT 43.800 82.800 44.200 83.200 ;
        RECT 44.600 83.100 45.000 88.900 ;
        RECT 48.600 87.200 48.900 106.800 ;
        RECT 49.400 103.100 49.800 108.900 ;
        RECT 50.200 104.200 50.500 112.800 ;
        RECT 51.800 110.200 52.100 113.800 ;
        RECT 52.600 112.100 53.000 112.200 ;
        RECT 53.400 112.100 53.800 112.200 ;
        RECT 52.600 111.800 53.800 112.100 ;
        RECT 51.800 109.800 52.200 110.200 ;
        RECT 54.200 110.100 54.500 124.800 ;
        RECT 55.000 112.100 55.400 117.900 ;
        RECT 53.400 109.800 54.500 110.100 ;
        RECT 52.600 106.800 53.000 107.200 ;
        RECT 52.600 106.200 52.900 106.800 ;
        RECT 52.600 105.800 53.000 106.200 ;
        RECT 50.200 103.800 50.600 104.200 ;
        RECT 50.200 97.200 50.500 103.800 ;
        RECT 52.600 99.800 53.000 100.200 ;
        RECT 52.600 97.200 52.900 99.800 ;
        RECT 50.200 96.800 50.600 97.200 ;
        RECT 51.800 96.800 52.200 97.200 ;
        RECT 52.600 96.800 53.000 97.200 ;
        RECT 51.800 96.200 52.100 96.800 ;
        RECT 49.400 95.800 49.800 96.200 ;
        RECT 51.800 95.800 52.200 96.200 ;
        RECT 49.400 92.200 49.700 95.800 ;
        RECT 49.400 91.800 49.800 92.200 ;
        RECT 51.800 91.800 52.200 92.200 ;
        RECT 51.800 91.200 52.100 91.800 ;
        RECT 51.800 90.800 52.200 91.200 ;
        RECT 51.800 89.100 52.200 89.200 ;
        RECT 52.600 89.100 53.000 89.200 ;
        RECT 48.600 86.800 49.000 87.200 ;
        RECT 46.200 86.100 46.600 86.200 ;
        RECT 47.000 86.100 47.400 86.200 ;
        RECT 46.200 85.800 47.400 86.100 ;
        RECT 47.800 83.800 48.200 84.200 ;
        RECT 42.200 81.800 42.600 82.200 ;
        RECT 44.600 81.800 45.000 82.200 ;
        RECT 44.600 79.200 44.900 81.800 ;
        RECT 30.200 79.100 30.600 79.200 ;
        RECT 31.000 79.100 31.400 79.200 ;
        RECT 30.200 78.800 31.400 79.100 ;
        RECT 35.000 78.800 35.400 79.200 ;
        RECT 44.600 78.800 45.000 79.200 ;
        RECT 46.200 78.800 46.600 79.200 ;
        RECT 26.200 74.800 26.600 75.200 ;
        RECT 27.000 74.800 27.400 75.200 ;
        RECT 25.400 65.800 25.800 66.200 ;
        RECT 20.600 55.800 21.000 56.200 ;
        RECT 20.600 55.200 20.900 55.800 ;
        RECT 20.600 54.800 21.000 55.200 ;
        RECT 20.600 54.200 20.900 54.800 ;
        RECT 20.600 53.800 21.000 54.200 ;
        RECT 19.800 52.800 20.200 53.200 ;
        RECT 17.400 48.800 17.800 49.200 ;
        RECT 15.800 47.800 16.200 48.200 ;
        RECT 15.800 47.200 16.100 47.800 ;
        RECT 14.200 46.800 14.600 47.200 ;
        RECT 15.000 46.800 15.400 47.200 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 14.200 46.200 14.500 46.800 ;
        RECT 10.200 45.800 10.600 46.200 ;
        RECT 11.800 45.800 12.200 46.200 ;
        RECT 13.400 46.100 13.800 46.200 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 13.400 45.800 14.600 46.100 ;
        RECT 11.800 45.200 12.100 45.800 ;
        RECT 11.800 44.800 12.200 45.200 ;
        RECT 16.600 45.100 17.000 45.200 ;
        RECT 17.400 45.100 17.800 45.200 ;
        RECT 18.200 45.100 18.600 47.900 ;
        RECT 16.600 44.800 17.800 45.100 ;
        RECT 14.200 43.800 14.600 44.200 ;
        RECT 14.200 39.200 14.500 43.800 ;
        RECT 19.800 43.100 20.200 48.900 ;
        RECT 22.200 47.800 22.600 48.200 ;
        RECT 21.400 46.800 21.800 47.200 ;
        RECT 21.400 42.200 21.700 46.800 ;
        RECT 22.200 46.200 22.500 47.800 ;
        RECT 22.200 45.800 22.600 46.200 ;
        RECT 24.600 43.100 25.000 48.900 ;
        RECT 21.400 41.800 21.800 42.200 ;
        RECT 14.200 38.800 14.600 39.200 ;
        RECT 7.800 35.800 8.900 36.100 ;
        RECT 0.600 31.800 1.000 32.200 ;
        RECT 0.600 25.200 0.900 31.800 ;
        RECT 2.200 26.200 2.500 35.800 ;
        RECT 7.800 35.200 8.100 35.800 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 5.400 35.100 5.800 35.200 ;
        RECT 6.200 35.100 6.600 35.200 ;
        RECT 5.400 34.800 6.600 35.100 ;
        RECT 7.800 34.800 8.200 35.200 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 13.400 35.100 13.800 35.200 ;
        RECT 12.600 34.800 13.800 35.100 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 3.800 34.200 4.100 34.800 ;
        RECT 14.200 34.200 14.500 34.800 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 4.600 33.800 5.000 34.200 ;
        RECT 14.200 33.800 14.600 34.200 ;
        RECT 15.000 33.800 15.400 34.200 ;
        RECT 3.000 32.800 3.400 33.200 ;
        RECT 3.000 29.100 3.300 32.800 ;
        RECT 3.800 29.100 4.200 29.200 ;
        RECT 3.000 28.800 4.200 29.100 ;
        RECT 4.600 27.200 4.900 33.800 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 7.000 31.800 7.400 32.200 ;
        RECT 7.000 31.200 7.300 31.800 ;
        RECT 7.000 30.800 7.400 31.200 ;
        RECT 10.200 29.200 10.500 32.800 ;
        RECT 15.000 32.200 15.300 33.800 ;
        RECT 15.800 33.100 16.200 35.900 ;
        RECT 15.000 31.800 15.400 32.200 ;
        RECT 17.400 32.100 17.800 37.900 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 17.400 30.800 17.800 31.200 ;
        RECT 3.000 27.100 3.400 27.200 ;
        RECT 3.800 27.100 4.200 27.200 ;
        RECT 3.000 26.800 4.200 27.100 ;
        RECT 4.600 26.800 5.000 27.200 ;
        RECT 2.200 26.100 2.600 26.200 ;
        RECT 3.000 26.100 3.400 26.200 ;
        RECT 2.200 25.800 3.400 26.100 ;
        RECT 0.600 24.800 1.000 25.200 ;
        RECT 2.200 24.800 2.600 25.200 ;
        RECT 2.200 24.200 2.500 24.800 ;
        RECT 2.200 23.800 2.600 24.200 ;
        RECT 0.600 13.100 1.000 15.900 ;
        RECT 2.200 12.100 2.600 17.900 ;
        RECT 3.000 14.700 3.400 15.100 ;
        RECT 3.000 9.200 3.300 14.700 ;
        RECT 4.600 11.200 4.900 26.800 ;
        RECT 5.400 23.800 5.800 24.200 ;
        RECT 5.400 15.200 5.700 23.800 ;
        RECT 6.200 23.100 6.600 28.900 ;
        RECT 10.200 28.800 10.600 29.200 ;
        RECT 12.600 29.100 13.000 29.200 ;
        RECT 13.400 29.100 13.800 29.200 ;
        RECT 9.400 25.800 9.800 26.200 ;
        RECT 9.400 25.200 9.700 25.800 ;
        RECT 9.400 24.800 9.800 25.200 ;
        RECT 11.000 23.100 11.400 28.900 ;
        RECT 12.600 28.800 13.800 29.100 ;
        RECT 11.800 27.800 12.200 28.200 ;
        RECT 11.800 27.200 12.100 27.800 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 12.600 25.100 13.000 27.900 ;
        RECT 15.800 23.100 16.200 28.900 ;
        RECT 17.400 26.200 17.700 30.800 ;
        RECT 17.400 25.800 17.800 26.200 ;
        RECT 9.400 19.100 9.800 19.200 ;
        RECT 10.200 19.100 10.600 19.200 ;
        RECT 9.400 18.800 10.600 19.100 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 6.200 12.800 6.600 13.200 ;
        RECT 4.600 10.800 5.000 11.200 ;
        RECT 0.600 9.100 1.000 9.200 ;
        RECT 1.400 9.100 1.800 9.200 ;
        RECT 0.600 8.800 1.800 9.100 ;
        RECT 3.000 8.800 3.400 9.200 ;
        RECT 4.600 7.200 4.900 10.800 ;
        RECT 6.200 8.100 6.500 12.800 ;
        RECT 7.000 12.100 7.400 17.900 ;
        RECT 11.000 16.800 11.400 17.200 ;
        RECT 11.000 15.200 11.300 16.800 ;
        RECT 11.800 16.100 12.200 16.200 ;
        RECT 12.600 16.100 13.000 16.200 ;
        RECT 11.800 15.800 13.000 16.100 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 10.200 13.800 10.600 14.200 ;
        RECT 10.200 13.200 10.500 13.800 ;
        RECT 10.200 12.800 10.600 13.200 ;
        RECT 5.400 7.800 6.500 8.100 ;
        RECT 5.400 7.200 5.700 7.800 ;
        RECT 3.800 7.100 4.200 7.200 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 3.800 6.800 5.000 7.100 ;
        RECT 5.400 6.800 5.800 7.200 ;
        RECT 6.200 6.800 6.600 7.200 ;
        RECT 6.200 6.200 6.500 6.800 ;
        RECT 0.600 5.800 1.000 6.200 ;
        RECT 4.600 6.100 5.000 6.200 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 4.600 5.800 5.800 6.100 ;
        RECT 6.200 5.800 6.600 6.200 ;
        RECT 0.600 5.200 0.900 5.800 ;
        RECT 11.000 5.200 11.300 14.800 ;
        RECT 12.600 14.200 12.900 14.800 ;
        RECT 12.600 13.800 13.000 14.200 ;
        RECT 13.400 13.100 13.800 15.900 ;
        RECT 14.200 15.800 14.600 16.200 ;
        RECT 14.200 9.200 14.500 15.800 ;
        RECT 15.000 12.100 15.400 17.900 ;
        RECT 15.800 14.700 16.200 15.100 ;
        RECT 15.800 14.200 16.100 14.700 ;
        RECT 15.800 13.800 16.200 14.200 ;
        RECT 18.200 9.200 18.500 35.800 ;
        RECT 21.400 35.200 21.700 41.800 ;
        RECT 26.200 39.200 26.500 74.800 ;
        RECT 27.000 66.200 27.300 74.800 ;
        RECT 27.800 72.100 28.200 77.900 ;
        RECT 35.800 77.800 36.200 78.200 ;
        RECT 31.000 75.100 31.400 75.200 ;
        RECT 31.800 75.100 32.200 75.200 ;
        RECT 31.000 74.800 32.200 75.100 ;
        RECT 33.400 75.100 33.800 75.200 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 33.400 74.800 34.600 75.100 ;
        RECT 30.200 74.100 30.600 74.200 ;
        RECT 31.000 74.100 31.400 74.200 ;
        RECT 30.200 73.800 31.400 74.100 ;
        RECT 32.600 73.800 33.000 74.200 ;
        RECT 31.000 69.100 31.400 69.200 ;
        RECT 31.800 69.100 32.200 69.200 ;
        RECT 27.000 65.800 27.400 66.200 ;
        RECT 27.000 59.200 27.300 65.800 ;
        RECT 28.600 63.100 29.000 68.900 ;
        RECT 31.000 68.800 32.200 69.100 ;
        RECT 31.000 67.100 31.400 67.200 ;
        RECT 31.800 67.100 32.200 67.200 ;
        RECT 31.000 66.800 32.200 67.100 ;
        RECT 32.600 66.200 32.900 73.800 ;
        RECT 35.800 73.200 36.100 77.800 ;
        RECT 46.200 76.200 46.500 78.800 ;
        RECT 36.600 75.800 37.000 76.200 ;
        RECT 42.200 75.800 42.600 76.200 ;
        RECT 46.200 75.800 46.600 76.200 ;
        RECT 36.600 73.200 36.900 75.800 ;
        RECT 42.200 75.200 42.500 75.800 ;
        RECT 47.800 75.200 48.100 83.800 ;
        RECT 49.400 83.100 49.800 88.900 ;
        RECT 51.800 88.800 53.000 89.100 ;
        RECT 53.400 88.200 53.700 109.800 ;
        RECT 54.200 103.100 54.600 108.900 ;
        RECT 54.200 96.800 54.600 97.200 ;
        RECT 54.200 96.200 54.500 96.800 ;
        RECT 54.200 95.800 54.600 96.200 ;
        RECT 55.800 95.200 56.100 125.800 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 65.400 125.100 65.800 127.900 ;
        RECT 61.400 123.800 61.800 124.200 ;
        RECT 59.000 121.800 59.400 122.200 ;
        RECT 59.000 118.200 59.300 121.800 ;
        RECT 59.000 117.800 59.400 118.200 ;
        RECT 59.000 116.800 59.400 117.200 ;
        RECT 56.600 115.100 57.000 115.200 ;
        RECT 57.400 115.100 57.800 115.200 ;
        RECT 56.600 114.800 57.800 115.100 ;
        RECT 57.400 111.800 57.800 112.200 ;
        RECT 56.600 109.800 57.000 110.200 ;
        RECT 56.600 109.200 56.900 109.800 ;
        RECT 56.600 108.800 57.000 109.200 ;
        RECT 57.400 108.200 57.700 111.800 ;
        RECT 59.000 109.200 59.300 116.800 ;
        RECT 59.800 112.100 60.200 117.900 ;
        RECT 61.400 117.200 61.700 123.800 ;
        RECT 61.400 116.800 61.800 117.200 ;
        RECT 60.600 113.800 61.000 114.200 ;
        RECT 60.600 110.200 60.900 113.800 ;
        RECT 61.400 113.100 61.800 115.900 ;
        RECT 62.200 113.800 62.600 114.200 ;
        RECT 62.200 113.200 62.500 113.800 ;
        RECT 62.200 112.800 62.600 113.200 ;
        RECT 60.600 109.800 61.000 110.200 ;
        RECT 59.000 108.800 59.400 109.200 ;
        RECT 57.400 107.800 57.800 108.200 ;
        RECT 59.000 107.200 59.300 108.800 ;
        RECT 59.000 106.800 59.400 107.200 ;
        RECT 60.600 107.100 61.000 107.200 ;
        RECT 61.400 107.100 61.800 107.200 ;
        RECT 60.600 106.800 61.800 107.100 ;
        RECT 63.000 106.200 63.300 124.800 ;
        RECT 64.600 121.800 65.000 122.200 ;
        RECT 64.600 115.200 64.900 121.800 ;
        RECT 64.600 114.800 65.000 115.200 ;
        RECT 65.400 115.100 65.800 115.200 ;
        RECT 66.200 115.100 66.500 129.800 ;
        RECT 67.000 123.100 67.400 128.900 ;
        RECT 69.400 125.800 69.800 126.200 ;
        RECT 70.200 125.800 70.600 126.200 ;
        RECT 69.400 119.200 69.700 125.800 ;
        RECT 69.400 118.800 69.800 119.200 ;
        RECT 65.400 114.800 66.500 115.100 ;
        RECT 68.600 115.100 69.000 115.200 ;
        RECT 69.400 115.100 69.800 115.200 ;
        RECT 68.600 114.800 69.800 115.100 ;
        RECT 63.800 113.800 64.200 114.200 ;
        RECT 68.600 113.800 69.000 114.200 ;
        RECT 63.800 113.200 64.100 113.800 ;
        RECT 68.600 113.200 68.900 113.800 ;
        RECT 63.800 112.800 64.200 113.200 ;
        RECT 64.600 112.800 65.000 113.200 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 68.600 112.800 69.000 113.200 ;
        RECT 64.600 112.200 64.900 112.800 ;
        RECT 67.000 112.200 67.300 112.800 ;
        RECT 64.600 111.800 65.000 112.200 ;
        RECT 67.000 111.800 67.400 112.200 ;
        RECT 65.400 109.800 65.800 110.200 ;
        RECT 63.800 106.800 64.200 107.200 ;
        RECT 63.000 105.800 63.400 106.200 ;
        RECT 63.000 105.200 63.300 105.800 ;
        RECT 60.600 105.100 61.000 105.200 ;
        RECT 61.400 105.100 61.800 105.200 ;
        RECT 60.600 104.800 61.800 105.100 ;
        RECT 63.000 104.800 63.400 105.200 ;
        RECT 59.000 103.800 59.400 104.200 ;
        RECT 60.600 103.800 61.000 104.200 ;
        RECT 57.400 96.800 57.800 97.200 ;
        RECT 57.400 96.200 57.700 96.800 ;
        RECT 57.400 95.800 57.800 96.200 ;
        RECT 54.200 94.800 54.600 95.200 ;
        RECT 55.800 94.800 56.200 95.200 ;
        RECT 54.200 94.200 54.500 94.800 ;
        RECT 54.200 93.800 54.600 94.200 ;
        RECT 55.000 93.800 55.400 94.200 ;
        RECT 55.000 93.200 55.300 93.800 ;
        RECT 55.000 92.800 55.400 93.200 ;
        RECT 55.000 91.800 55.400 92.200 ;
        RECT 53.400 87.800 53.800 88.200 ;
        RECT 52.600 86.800 53.000 87.200 ;
        RECT 49.400 77.800 49.800 78.200 ;
        RECT 49.400 76.200 49.700 77.800 ;
        RECT 51.000 76.800 51.400 77.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 50.200 75.800 50.600 76.200 ;
        RECT 50.200 75.200 50.500 75.800 ;
        RECT 40.600 74.800 41.000 75.200 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 47.800 74.800 48.200 75.200 ;
        RECT 50.200 74.800 50.600 75.200 ;
        RECT 38.200 74.100 38.600 74.200 ;
        RECT 39.000 74.100 39.400 74.200 ;
        RECT 38.200 73.800 39.400 74.100 ;
        RECT 35.800 72.800 36.200 73.200 ;
        RECT 36.600 72.800 37.000 73.200 ;
        RECT 39.800 72.800 40.200 73.200 ;
        RECT 35.800 69.200 36.100 72.800 ;
        RECT 38.200 72.100 38.600 72.200 ;
        RECT 39.000 72.100 39.400 72.200 ;
        RECT 38.200 71.800 39.400 72.100 ;
        RECT 39.800 69.200 40.100 72.800 ;
        RECT 40.600 72.200 40.900 74.800 ;
        RECT 43.000 74.200 43.300 74.800 ;
        RECT 44.600 74.200 44.900 74.800 ;
        RECT 41.400 74.100 41.800 74.200 ;
        RECT 42.200 74.100 42.600 74.200 ;
        RECT 41.400 73.800 42.600 74.100 ;
        RECT 43.000 73.800 43.400 74.200 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 44.600 73.800 45.000 74.200 ;
        RECT 47.000 73.800 47.400 74.200 ;
        RECT 48.600 73.800 49.000 74.200 ;
        RECT 51.000 74.100 51.300 76.800 ;
        RECT 50.200 73.800 51.300 74.100 ;
        RECT 52.600 74.200 52.900 86.800 ;
        RECT 53.400 86.200 53.700 87.800 ;
        RECT 53.400 85.800 53.800 86.200 ;
        RECT 54.200 85.800 54.600 86.200 ;
        RECT 54.200 85.200 54.500 85.800 ;
        RECT 54.200 84.800 54.600 85.200 ;
        RECT 53.400 76.100 53.800 76.200 ;
        RECT 54.200 76.100 54.600 76.200 ;
        RECT 53.400 75.800 54.600 76.100 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 43.800 73.200 44.100 73.800 ;
        RECT 43.800 72.800 44.200 73.200 ;
        RECT 40.600 71.800 41.000 72.200 ;
        RECT 42.200 72.100 42.600 72.200 ;
        RECT 41.400 71.800 42.600 72.100 ;
        RECT 35.800 68.800 36.200 69.200 ;
        RECT 39.800 68.800 40.200 69.200 ;
        RECT 35.800 68.100 36.200 68.200 ;
        RECT 36.600 68.100 37.000 68.200 ;
        RECT 35.800 67.800 37.000 68.100 ;
        RECT 35.000 66.800 35.400 67.200 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 41.400 66.200 41.700 71.800 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 45.400 67.100 45.800 67.200 ;
        RECT 46.200 67.100 46.600 67.200 ;
        RECT 45.400 66.800 46.600 67.100 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 32.600 65.800 33.000 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 29.400 62.800 29.800 63.200 ;
        RECT 29.400 59.200 29.700 62.800 ;
        RECT 31.800 59.200 32.100 65.800 ;
        RECT 34.200 64.800 34.600 65.200 ;
        RECT 27.000 58.800 27.400 59.200 ;
        RECT 29.400 58.800 29.800 59.200 ;
        RECT 31.800 58.800 32.200 59.200 ;
        RECT 34.200 58.200 34.500 64.800 ;
        RECT 37.400 64.200 37.700 65.800 ;
        RECT 39.800 64.800 40.200 65.200 ;
        RECT 37.400 63.800 37.800 64.200 ;
        RECT 39.800 63.200 40.100 64.800 ;
        RECT 39.800 62.800 40.200 63.200 ;
        RECT 34.200 57.800 34.600 58.200 ;
        RECT 29.400 56.800 29.800 57.200 ;
        RECT 30.200 56.800 30.600 57.200 ;
        RECT 35.000 56.800 35.400 57.200 ;
        RECT 27.000 55.100 27.400 55.200 ;
        RECT 27.800 55.100 28.200 55.200 ;
        RECT 27.000 54.800 28.200 55.100 ;
        RECT 27.800 54.100 28.200 54.200 ;
        RECT 28.600 54.100 29.000 54.200 ;
        RECT 27.800 53.800 29.000 54.100 ;
        RECT 28.600 52.800 29.000 53.200 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 27.000 46.100 27.400 46.200 ;
        RECT 27.800 46.100 28.100 46.800 ;
        RECT 27.000 45.800 28.100 46.100 ;
        RECT 26.200 38.800 26.600 39.200 ;
        RECT 19.000 34.800 19.400 35.200 ;
        RECT 21.400 34.800 21.800 35.200 ;
        RECT 19.000 33.200 19.300 34.800 ;
        RECT 19.000 32.800 19.400 33.200 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 19.000 15.200 19.300 26.800 ;
        RECT 20.600 23.100 21.000 28.900 ;
        RECT 21.400 28.200 21.700 34.800 ;
        RECT 22.200 32.100 22.600 37.900 ;
        RECT 28.600 35.200 28.900 52.800 ;
        RECT 29.400 46.200 29.700 56.800 ;
        RECT 30.200 56.200 30.500 56.800 ;
        RECT 30.200 55.800 30.600 56.200 ;
        RECT 34.200 55.800 34.600 56.200 ;
        RECT 31.800 54.800 32.200 55.200 ;
        RECT 31.000 53.800 31.400 54.200 ;
        RECT 30.200 48.800 30.600 49.200 ;
        RECT 30.200 48.200 30.500 48.800 ;
        RECT 30.200 47.800 30.600 48.200 ;
        RECT 29.400 45.800 29.800 46.200 ;
        RECT 29.400 45.200 29.700 45.800 ;
        RECT 29.400 44.800 29.800 45.200 ;
        RECT 29.400 41.800 29.800 42.200 ;
        RECT 29.400 39.200 29.700 41.800 ;
        RECT 29.400 38.800 29.800 39.200 ;
        RECT 27.800 35.100 28.200 35.200 ;
        RECT 28.600 35.100 29.000 35.200 ;
        RECT 27.800 34.800 29.000 35.100 ;
        RECT 23.800 33.800 24.200 34.200 ;
        RECT 26.200 34.100 26.600 34.200 ;
        RECT 27.000 34.100 27.400 34.200 ;
        RECT 26.200 33.800 27.400 34.100 ;
        RECT 29.400 34.100 29.800 34.200 ;
        RECT 30.200 34.100 30.600 34.200 ;
        RECT 29.400 33.800 30.600 34.100 ;
        RECT 23.800 29.200 24.100 33.800 ;
        RECT 27.000 32.800 27.400 33.200 ;
        RECT 24.600 31.800 25.000 32.200 ;
        RECT 23.800 28.800 24.200 29.200 ;
        RECT 21.400 27.800 21.800 28.200 ;
        RECT 21.400 27.200 21.700 27.800 ;
        RECT 21.400 26.800 21.800 27.200 ;
        RECT 22.200 25.100 22.600 27.900 ;
        RECT 23.000 27.800 23.400 28.200 ;
        RECT 23.800 27.800 24.200 28.200 ;
        RECT 23.000 19.200 23.300 27.800 ;
        RECT 23.800 19.200 24.100 27.800 ;
        RECT 24.600 27.200 24.900 31.800 ;
        RECT 27.000 29.200 27.300 32.800 ;
        RECT 29.400 32.200 29.700 33.800 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 28.600 30.800 29.000 31.200 ;
        RECT 27.000 28.800 27.400 29.200 ;
        RECT 24.600 26.800 25.000 27.200 ;
        RECT 28.600 26.200 28.900 30.800 ;
        RECT 31.000 28.200 31.300 53.800 ;
        RECT 31.800 53.200 32.100 54.800 ;
        RECT 32.600 53.800 33.000 54.200 ;
        RECT 31.800 52.800 32.200 53.200 ;
        RECT 32.600 51.200 32.900 53.800 ;
        RECT 32.600 50.800 33.000 51.200 ;
        RECT 32.600 47.200 32.900 50.800 ;
        RECT 34.200 49.200 34.500 55.800 ;
        RECT 34.200 48.800 34.600 49.200 ;
        RECT 32.600 46.800 33.000 47.200 ;
        RECT 33.400 46.800 33.800 47.200 ;
        RECT 33.400 46.200 33.700 46.800 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 31.800 45.800 33.000 46.100 ;
        RECT 33.400 45.800 33.800 46.200 ;
        RECT 35.000 45.200 35.300 56.800 ;
        RECT 35.800 53.100 36.200 55.900 ;
        RECT 36.600 54.800 37.000 55.200 ;
        RECT 36.600 54.200 36.900 54.800 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 37.400 52.100 37.800 57.900 ;
        RECT 39.800 55.100 40.200 55.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 39.800 54.800 41.000 55.100 ;
        RECT 41.400 53.200 41.700 65.800 ;
        RECT 42.200 65.200 42.500 66.800 ;
        RECT 47.000 66.200 47.300 73.800 ;
        RECT 48.600 67.200 48.900 73.800 ;
        RECT 49.400 71.800 49.800 72.200 ;
        RECT 48.600 66.800 49.000 67.200 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 47.000 65.800 47.400 66.200 ;
        RECT 42.200 64.800 42.600 65.200 ;
        RECT 43.000 64.200 43.300 65.800 ;
        RECT 48.600 65.100 49.000 65.200 ;
        RECT 49.400 65.100 49.700 71.800 ;
        RECT 50.200 69.200 50.500 73.800 ;
        RECT 52.600 70.200 52.900 73.800 ;
        RECT 53.400 71.800 53.800 72.200 ;
        RECT 52.600 69.800 53.000 70.200 ;
        RECT 50.200 68.800 50.600 69.200 ;
        RECT 51.000 65.100 51.400 67.900 ;
        RECT 48.600 64.800 49.700 65.100 ;
        RECT 43.000 63.800 43.400 64.200 ;
        RECT 50.200 63.800 50.600 64.200 ;
        RECT 43.000 59.200 43.300 63.800 ;
        RECT 47.000 62.800 47.400 63.200 ;
        RECT 47.000 62.200 47.300 62.800 ;
        RECT 44.600 61.800 45.000 62.200 ;
        RECT 47.000 61.800 47.400 62.200 ;
        RECT 44.600 60.200 44.900 61.800 ;
        RECT 44.600 59.800 45.000 60.200 ;
        RECT 43.000 58.800 43.400 59.200 ;
        RECT 41.400 52.800 41.800 53.200 ;
        RECT 42.200 52.100 42.600 57.900 ;
        RECT 50.200 57.200 50.500 63.800 ;
        RECT 52.600 63.100 53.000 68.900 ;
        RECT 53.400 66.300 53.700 71.800 ;
        RECT 53.400 65.900 53.800 66.300 ;
        RECT 53.400 64.800 53.800 65.200 ;
        RECT 53.400 59.200 53.700 64.800 ;
        RECT 53.400 58.800 53.800 59.200 ;
        RECT 55.000 58.200 55.300 91.800 ;
        RECT 55.800 89.100 56.100 94.800 ;
        RECT 57.400 93.800 57.800 94.200 ;
        RECT 57.400 93.200 57.700 93.800 ;
        RECT 57.400 92.800 57.800 93.200 ;
        RECT 58.200 93.100 58.600 95.900 ;
        RECT 55.800 88.800 56.900 89.100 ;
        RECT 55.800 87.800 56.200 88.200 ;
        RECT 55.800 85.200 56.100 87.800 ;
        RECT 55.800 84.800 56.200 85.200 ;
        RECT 55.800 75.200 56.100 84.800 ;
        RECT 56.600 84.200 56.900 88.800 ;
        RECT 57.400 88.800 57.800 89.200 ;
        RECT 57.400 87.200 57.700 88.800 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 59.000 87.100 59.300 103.800 ;
        RECT 59.800 92.100 60.200 97.900 ;
        RECT 60.600 90.200 60.900 103.800 ;
        RECT 61.400 95.100 61.800 95.200 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 61.400 94.800 62.600 95.100 ;
        RECT 60.600 89.800 61.000 90.200 ;
        RECT 59.800 87.100 60.200 87.200 ;
        RECT 59.000 86.800 60.200 87.100 ;
        RECT 60.600 86.200 60.900 89.800 ;
        RECT 63.000 89.200 63.300 104.800 ;
        RECT 63.800 102.200 64.100 106.800 ;
        RECT 64.600 105.100 65.000 107.900 ;
        RECT 65.400 107.200 65.700 109.800 ;
        RECT 65.400 106.800 65.800 107.200 ;
        RECT 63.800 101.800 64.200 102.200 ;
        RECT 63.800 97.200 64.100 101.800 ;
        RECT 63.800 96.800 64.200 97.200 ;
        RECT 63.800 94.800 64.200 95.200 ;
        RECT 63.800 93.200 64.100 94.800 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 64.600 92.100 65.000 97.900 ;
        RECT 65.400 97.200 65.700 106.800 ;
        RECT 66.200 103.100 66.600 108.900 ;
        RECT 67.000 106.100 67.400 106.200 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 67.000 105.800 68.200 106.100 ;
        RECT 68.600 103.200 68.900 112.800 ;
        RECT 69.400 110.800 69.800 111.200 ;
        RECT 68.600 102.800 69.000 103.200 ;
        RECT 68.600 102.200 68.900 102.800 ;
        RECT 68.600 101.800 69.000 102.200 ;
        RECT 69.400 98.200 69.700 110.800 ;
        RECT 70.200 107.200 70.500 125.800 ;
        RECT 71.800 123.100 72.200 128.900 ;
        RECT 74.200 128.800 74.600 129.200 ;
        RECT 74.200 128.200 74.500 128.800 ;
        RECT 75.000 128.200 75.300 131.800 ;
        RECT 76.600 130.200 76.900 131.800 ;
        RECT 76.600 129.800 77.000 130.200 ;
        RECT 74.200 127.800 74.600 128.200 ;
        RECT 75.000 127.800 75.400 128.200 ;
        RECT 75.800 128.100 76.200 128.200 ;
        RECT 76.600 128.100 77.000 128.200 ;
        RECT 75.800 127.800 77.000 128.100 ;
        RECT 77.400 127.800 77.800 128.200 ;
        RECT 77.400 127.200 77.700 127.800 ;
        RECT 78.200 127.200 78.500 132.800 ;
        RECT 79.000 131.800 79.400 132.200 ;
        RECT 87.800 132.100 88.100 133.800 ;
        RECT 88.600 132.100 89.000 137.900 ;
        RECT 90.200 135.100 90.600 135.200 ;
        RECT 89.400 134.800 90.600 135.100 ;
        RECT 89.400 134.700 89.800 134.800 ;
        RECT 87.000 131.800 88.100 132.100 ;
        RECT 77.400 126.800 77.800 127.200 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 79.000 126.200 79.300 131.800 ;
        RECT 80.600 127.100 81.000 127.200 ;
        RECT 81.400 127.100 81.800 127.200 ;
        RECT 80.600 126.800 81.800 127.100 ;
        RECT 83.000 126.800 83.400 127.200 ;
        RECT 79.000 125.800 79.400 126.200 ;
        RECT 79.000 125.200 79.300 125.800 ;
        RECT 79.000 124.800 79.400 125.200 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 81.400 124.800 82.600 125.100 ;
        RECT 75.000 123.800 75.400 124.200 ;
        RECT 81.400 123.800 81.800 124.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 74.200 117.200 74.500 121.800 ;
        RECT 71.800 116.800 72.200 117.200 ;
        RECT 74.200 116.800 74.600 117.200 ;
        RECT 71.800 116.200 72.100 116.800 ;
        RECT 71.800 115.800 72.200 116.200 ;
        RECT 73.400 114.800 73.800 115.200 ;
        RECT 70.200 106.800 70.600 107.200 ;
        RECT 71.000 103.100 71.400 108.900 ;
        RECT 73.400 107.200 73.700 114.800 ;
        RECT 75.000 114.200 75.300 123.800 ;
        RECT 81.400 119.200 81.700 123.800 ;
        RECT 83.000 120.200 83.300 126.800 ;
        RECT 83.800 125.100 84.200 127.900 ;
        RECT 85.400 123.100 85.800 128.900 ;
        RECT 87.000 127.200 87.300 131.800 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 87.000 126.800 87.400 127.200 ;
        RECT 86.200 126.300 86.500 126.800 ;
        RECT 86.200 125.900 86.600 126.300 ;
        RECT 86.200 125.800 86.500 125.900 ;
        RECT 83.000 119.800 83.400 120.200 ;
        RECT 81.400 118.800 81.800 119.200 ;
        RECT 83.000 116.800 83.400 117.200 ;
        RECT 83.000 116.200 83.300 116.800 ;
        RECT 79.000 115.800 79.400 116.200 ;
        RECT 79.800 115.800 80.200 116.200 ;
        RECT 83.000 115.800 83.400 116.200 ;
        RECT 79.000 115.200 79.300 115.800 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 77.400 115.100 77.800 115.200 ;
        RECT 78.200 115.100 78.600 115.200 ;
        RECT 77.400 114.800 78.600 115.100 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 74.200 113.800 74.600 114.200 ;
        RECT 75.000 113.800 75.400 114.200 ;
        RECT 74.200 112.200 74.500 113.800 ;
        RECT 74.200 111.800 74.600 112.200 ;
        RECT 74.200 110.800 74.600 111.200 ;
        RECT 73.400 106.800 73.800 107.200 ;
        RECT 74.200 106.200 74.500 110.800 ;
        RECT 74.200 106.100 74.600 106.200 ;
        RECT 74.200 105.800 75.300 106.100 ;
        RECT 73.400 104.800 73.800 105.200 ;
        RECT 73.400 104.200 73.700 104.800 ;
        RECT 73.400 103.800 73.800 104.200 ;
        RECT 75.000 101.200 75.300 105.800 ;
        RECT 75.800 104.200 76.100 114.800 ;
        RECT 78.200 113.800 78.600 114.200 ;
        RECT 78.200 113.200 78.500 113.800 ;
        RECT 79.800 113.200 80.100 115.800 ;
        RECT 80.600 114.100 81.000 114.200 ;
        RECT 80.600 113.800 81.700 114.100 ;
        RECT 76.600 113.100 77.000 113.200 ;
        RECT 77.400 113.100 77.800 113.200 ;
        RECT 76.600 112.800 77.800 113.100 ;
        RECT 78.200 112.800 78.600 113.200 ;
        RECT 79.800 112.800 80.200 113.200 ;
        RECT 77.400 111.800 77.800 112.200 ;
        RECT 80.600 111.800 81.000 112.200 ;
        RECT 77.400 107.200 77.700 111.800 ;
        RECT 80.600 107.200 80.900 111.800 ;
        RECT 81.400 107.200 81.700 113.800 ;
        RECT 85.400 112.100 85.800 117.900 ;
        RECT 87.000 115.200 87.300 126.800 ;
        RECT 90.200 123.100 90.600 128.900 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 88.600 115.000 89.000 115.100 ;
        RECT 89.400 115.000 89.800 115.100 ;
        RECT 85.400 107.800 85.800 108.200 ;
        RECT 77.400 106.800 77.800 107.200 ;
        RECT 78.200 106.800 78.600 107.200 ;
        RECT 80.600 106.800 81.000 107.200 ;
        RECT 81.400 106.800 81.800 107.200 ;
        RECT 83.800 106.800 84.200 107.200 ;
        RECT 78.200 106.200 78.500 106.800 ;
        RECT 81.400 106.200 81.700 106.800 ;
        RECT 83.800 106.200 84.100 106.800 ;
        RECT 85.400 106.200 85.700 107.800 ;
        RECT 86.200 106.800 86.600 107.200 ;
        RECT 87.000 107.100 87.300 114.800 ;
        RECT 88.600 114.700 89.800 115.000 ;
        RECT 90.200 112.100 90.600 117.900 ;
        RECT 87.800 107.100 88.200 107.200 ;
        RECT 87.000 106.800 88.200 107.100 ;
        RECT 78.200 105.800 78.600 106.200 ;
        RECT 79.000 105.800 79.400 106.200 ;
        RECT 81.400 105.800 81.800 106.200 ;
        RECT 83.800 105.800 84.200 106.200 ;
        RECT 85.400 105.800 85.800 106.200 ;
        RECT 75.800 103.800 76.200 104.200 ;
        RECT 74.200 100.800 74.600 101.200 ;
        RECT 75.000 100.800 75.400 101.200 ;
        RECT 74.200 99.200 74.500 100.800 ;
        RECT 74.200 98.800 74.600 99.200 ;
        RECT 75.000 99.100 75.300 100.800 ;
        RECT 75.800 100.200 76.100 103.800 ;
        RECT 76.600 101.800 77.000 102.200 ;
        RECT 75.800 99.800 76.200 100.200 ;
        RECT 75.000 98.800 76.100 99.100 ;
        RECT 69.400 97.800 69.800 98.200 ;
        RECT 71.800 97.800 72.200 98.200 ;
        RECT 65.400 96.800 65.800 97.200 ;
        RECT 67.800 96.800 68.200 97.200 ;
        RECT 67.800 94.200 68.100 96.800 ;
        RECT 69.400 96.200 69.700 97.800 ;
        RECT 69.400 95.800 69.800 96.200 ;
        RECT 71.800 95.200 72.100 97.800 ;
        RECT 72.600 96.800 73.000 97.200 ;
        RECT 69.400 94.800 69.800 95.200 ;
        RECT 71.800 94.800 72.200 95.200 ;
        RECT 69.400 94.200 69.700 94.800 ;
        RECT 72.600 94.200 72.900 96.800 ;
        RECT 75.800 95.200 76.100 98.800 ;
        RECT 75.800 94.800 76.200 95.200 ;
        RECT 76.600 94.200 76.900 101.800 ;
        RECT 77.400 98.800 77.800 99.200 ;
        RECT 77.400 97.200 77.700 98.800 ;
        RECT 77.400 96.800 77.800 97.200 ;
        RECT 77.400 95.200 77.700 96.800 ;
        RECT 79.000 96.200 79.300 105.800 ;
        RECT 83.000 104.800 83.400 105.200 ;
        RECT 83.000 104.200 83.300 104.800 ;
        RECT 79.800 103.800 80.200 104.200 ;
        RECT 83.000 103.800 83.400 104.200 ;
        RECT 79.800 99.200 80.100 103.800 ;
        RECT 86.200 102.200 86.500 106.800 ;
        RECT 86.200 101.800 86.600 102.200 ;
        RECT 79.800 98.800 80.200 99.200 ;
        RECT 79.000 95.800 79.400 96.200 ;
        RECT 80.600 95.800 81.000 96.200 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 78.200 94.800 79.400 95.100 ;
        RECT 80.600 94.200 80.900 95.800 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 69.400 93.800 69.800 94.200 ;
        RECT 72.600 93.800 73.000 94.200 ;
        RECT 76.600 93.800 77.000 94.200 ;
        RECT 80.600 93.800 81.000 94.200 ;
        RECT 65.400 92.800 65.800 93.200 ;
        RECT 69.400 92.800 69.800 93.200 ;
        RECT 75.800 92.800 76.200 93.200 ;
        RECT 63.000 88.800 63.400 89.200 ;
        RECT 63.000 87.800 63.400 88.200 ;
        RECT 64.600 88.100 65.000 88.200 ;
        RECT 65.400 88.100 65.700 92.800 ;
        RECT 69.400 89.200 69.700 92.800 ;
        RECT 64.600 87.800 65.700 88.100 ;
        RECT 68.600 88.800 69.000 89.200 ;
        RECT 69.400 88.800 69.800 89.200 ;
        RECT 63.000 87.200 63.300 87.800 ;
        RECT 63.000 86.800 63.400 87.200 ;
        RECT 64.600 87.100 65.000 87.200 ;
        RECT 65.400 87.100 65.800 87.200 ;
        RECT 64.600 86.800 65.800 87.100 ;
        RECT 67.800 86.800 68.200 87.200 ;
        RECT 67.800 86.200 68.100 86.800 ;
        RECT 60.600 85.800 61.000 86.200 ;
        RECT 62.200 86.100 62.600 86.200 ;
        RECT 63.000 86.100 63.400 86.200 ;
        RECT 62.200 85.800 63.400 86.100 ;
        RECT 63.800 86.100 64.200 86.200 ;
        RECT 64.600 86.100 65.000 86.200 ;
        RECT 63.800 85.800 65.000 86.100 ;
        RECT 66.200 86.100 66.600 86.200 ;
        RECT 67.000 86.100 67.400 86.200 ;
        RECT 66.200 85.800 67.400 86.100 ;
        RECT 67.800 85.800 68.200 86.200 ;
        RECT 56.600 83.800 57.000 84.200 ;
        RECT 59.800 83.800 60.200 84.200 ;
        RECT 59.000 81.800 59.400 82.200 ;
        RECT 57.400 76.100 57.800 76.200 ;
        RECT 58.200 76.100 58.600 76.200 ;
        RECT 57.400 75.800 58.600 76.100 ;
        RECT 55.800 74.800 56.200 75.200 ;
        RECT 59.000 74.200 59.300 81.800 ;
        RECT 59.800 78.200 60.100 83.800 ;
        RECT 61.400 82.100 61.800 82.200 ;
        RECT 62.200 82.100 62.600 82.200 ;
        RECT 61.400 81.800 62.600 82.100 ;
        RECT 63.800 81.800 64.200 82.200 ;
        RECT 59.800 77.800 60.200 78.200 ;
        RECT 59.800 75.200 60.100 77.800 ;
        RECT 61.400 76.800 61.800 77.200 ;
        RECT 61.400 76.200 61.700 76.800 ;
        RECT 60.600 75.800 61.000 76.200 ;
        RECT 61.400 75.800 61.800 76.200 ;
        RECT 62.200 75.800 62.600 76.200 ;
        RECT 59.800 74.800 60.200 75.200 ;
        RECT 55.800 73.800 56.200 74.200 ;
        RECT 58.200 73.800 58.600 74.200 ;
        RECT 59.000 73.800 59.400 74.200 ;
        RECT 55.800 73.200 56.100 73.800 ;
        RECT 55.800 72.800 56.200 73.200 ;
        RECT 55.800 71.200 56.100 72.800 ;
        RECT 55.800 70.800 56.200 71.200 ;
        RECT 58.200 69.200 58.500 73.800 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 55.800 65.800 57.000 66.100 ;
        RECT 57.400 63.100 57.800 68.900 ;
        RECT 58.200 68.800 58.600 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 59.800 69.100 60.200 69.200 ;
        RECT 59.000 68.800 60.200 69.100 ;
        RECT 60.600 65.200 60.900 75.800 ;
        RECT 62.200 75.200 62.500 75.800 ;
        RECT 63.800 75.200 64.100 81.800 ;
        RECT 66.200 79.200 66.500 85.800 ;
        RECT 67.800 85.100 68.200 85.200 ;
        RECT 67.000 84.800 68.200 85.100 ;
        RECT 66.200 78.800 66.600 79.200 ;
        RECT 66.200 75.800 66.600 76.200 ;
        RECT 66.200 75.200 66.500 75.800 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 62.200 74.800 62.600 75.200 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 61.400 74.200 61.700 74.800 ;
        RECT 61.400 73.800 61.800 74.200 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 65.400 73.800 66.600 74.100 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 62.200 70.200 62.500 71.800 ;
        RECT 62.200 69.800 62.600 70.200 ;
        RECT 63.800 69.800 64.200 70.200 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 63.000 66.800 63.400 67.200 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 58.200 62.800 58.600 63.200 ;
        RECT 55.000 57.800 55.400 58.200 ;
        RECT 56.600 57.800 57.000 58.200 ;
        RECT 43.000 56.800 43.400 57.200 ;
        RECT 44.600 57.100 45.000 57.200 ;
        RECT 45.400 57.100 45.800 57.200 ;
        RECT 44.600 56.800 45.800 57.100 ;
        RECT 50.200 56.800 50.600 57.200 ;
        RECT 53.400 56.800 53.800 57.200 ;
        RECT 35.000 44.800 35.400 45.200 ;
        RECT 37.400 45.100 37.800 47.900 ;
        RECT 39.000 43.100 39.400 48.900 ;
        RECT 39.800 46.800 40.200 47.200 ;
        RECT 31.800 32.800 32.200 33.200 ;
        RECT 32.600 33.100 33.000 35.900 ;
        RECT 33.400 33.800 33.800 34.200 ;
        RECT 31.800 29.200 32.100 32.800 ;
        RECT 31.800 28.800 32.200 29.200 ;
        RECT 31.000 27.800 31.400 28.200 ;
        RECT 33.400 27.200 33.700 33.800 ;
        RECT 34.200 32.100 34.600 37.900 ;
        RECT 37.400 34.800 37.800 35.200 ;
        RECT 37.400 34.200 37.700 34.800 ;
        RECT 37.400 33.800 37.800 34.200 ;
        RECT 39.000 32.100 39.400 37.900 ;
        RECT 39.800 37.200 40.100 46.800 ;
        RECT 40.600 46.100 41.000 46.200 ;
        RECT 41.400 46.100 41.800 46.200 ;
        RECT 40.600 45.800 41.800 46.100 ;
        RECT 43.000 39.200 43.300 56.800 ;
        RECT 45.400 55.800 45.800 56.200 ;
        RECT 48.600 56.100 49.000 56.200 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 48.600 55.800 49.800 56.100 ;
        RECT 45.400 55.200 45.700 55.800 ;
        RECT 45.400 54.800 45.800 55.200 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 46.200 54.800 47.400 55.100 ;
        RECT 50.200 54.200 50.500 56.800 ;
        RECT 53.400 55.200 53.700 56.800 ;
        RECT 55.000 56.200 55.300 57.800 ;
        RECT 56.600 57.200 56.900 57.800 ;
        RECT 56.600 56.800 57.000 57.200 ;
        RECT 58.200 56.200 58.500 62.800 ;
        RECT 59.000 59.800 59.400 60.200 ;
        RECT 55.000 55.800 55.400 56.200 ;
        RECT 58.200 55.800 58.600 56.200 ;
        RECT 51.800 55.100 52.200 55.200 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 51.800 54.800 53.000 55.100 ;
        RECT 53.400 54.800 53.800 55.200 ;
        RECT 55.800 55.100 56.200 55.200 ;
        RECT 56.600 55.100 57.000 55.200 ;
        RECT 55.800 54.800 57.000 55.100 ;
        RECT 59.000 54.200 59.300 59.800 ;
        RECT 59.800 55.800 60.200 56.200 ;
        RECT 59.800 55.200 60.100 55.800 ;
        RECT 59.800 55.100 60.200 55.200 ;
        RECT 60.600 55.100 60.900 64.800 ;
        RECT 62.200 64.200 62.500 66.800 ;
        RECT 63.000 65.200 63.300 66.800 ;
        RECT 63.000 64.800 63.400 65.200 ;
        RECT 63.800 65.100 64.100 69.800 ;
        RECT 64.600 68.200 64.900 73.800 ;
        RECT 67.000 69.200 67.300 84.800 ;
        RECT 68.600 76.200 68.900 88.800 ;
        RECT 75.800 85.200 76.100 92.800 ;
        RECT 79.800 91.800 80.200 92.200 ;
        RECT 79.800 91.200 80.100 91.800 ;
        RECT 77.400 90.800 77.800 91.200 ;
        RECT 79.800 90.800 80.200 91.200 ;
        RECT 76.600 85.800 77.000 86.200 ;
        RECT 76.600 85.200 76.900 85.800 ;
        RECT 75.800 84.800 76.200 85.200 ;
        RECT 76.600 84.800 77.000 85.200 ;
        RECT 69.400 81.800 69.800 82.200 ;
        RECT 68.600 75.800 69.000 76.200 ;
        RECT 68.600 75.200 68.900 75.800 ;
        RECT 69.400 75.200 69.700 81.800 ;
        RECT 68.600 74.800 69.000 75.200 ;
        RECT 69.400 74.800 69.800 75.200 ;
        RECT 67.800 74.100 68.200 74.200 ;
        RECT 68.600 74.100 69.000 74.200 ;
        RECT 67.800 73.800 69.000 74.100 ;
        RECT 72.600 72.800 73.000 73.200 ;
        RECT 67.800 71.800 68.200 72.200 ;
        RECT 71.000 71.800 71.400 72.200 ;
        RECT 67.000 68.800 67.400 69.200 ;
        RECT 64.600 67.800 65.000 68.200 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 64.600 66.200 64.900 66.800 ;
        RECT 64.600 65.800 65.000 66.200 ;
        RECT 64.600 65.100 65.000 65.200 ;
        RECT 63.800 64.800 65.000 65.100 ;
        RECT 62.200 63.800 62.600 64.200 ;
        RECT 61.400 61.800 61.800 62.200 ;
        RECT 61.400 56.200 61.700 61.800 ;
        RECT 61.400 55.800 61.800 56.200 ;
        RECT 59.800 54.800 60.900 55.100 ;
        RECT 61.400 54.800 61.800 55.200 ;
        RECT 61.400 54.200 61.700 54.800 ;
        RECT 45.400 54.100 45.800 54.200 ;
        RECT 46.200 54.100 46.600 54.200 ;
        RECT 45.400 53.800 46.600 54.100 ;
        RECT 50.200 53.800 50.600 54.200 ;
        RECT 52.600 53.800 53.000 54.200 ;
        RECT 55.800 54.100 56.200 54.200 ;
        RECT 56.600 54.100 57.000 54.200 ;
        RECT 55.800 53.800 57.000 54.100 ;
        RECT 59.000 53.800 59.400 54.200 ;
        RECT 61.400 53.800 61.800 54.200 ;
        RECT 51.000 53.100 51.400 53.200 ;
        RECT 51.000 52.800 52.100 53.100 ;
        RECT 51.800 49.200 52.100 52.800 ;
        RECT 46.200 49.100 46.600 49.200 ;
        RECT 47.000 49.100 47.400 49.200 ;
        RECT 43.800 43.100 44.200 48.900 ;
        RECT 46.200 48.800 47.400 49.100 ;
        RECT 51.800 48.800 52.200 49.200 ;
        RECT 51.800 47.200 52.100 48.800 ;
        RECT 47.000 46.800 47.400 47.200 ;
        RECT 47.800 46.800 48.200 47.200 ;
        RECT 50.200 46.800 50.600 47.200 ;
        RECT 51.800 46.800 52.200 47.200 ;
        RECT 44.600 44.800 45.000 45.200 ;
        RECT 44.600 44.200 44.900 44.800 ;
        RECT 44.600 43.800 45.000 44.200 ;
        RECT 40.600 38.800 41.000 39.200 ;
        RECT 43.000 38.800 43.400 39.200 ;
        RECT 39.800 36.800 40.200 37.200 ;
        RECT 39.000 29.100 39.400 29.200 ;
        RECT 39.800 29.100 40.200 29.200 ;
        RECT 39.000 28.800 40.200 29.100 ;
        RECT 29.400 26.800 29.800 27.200 ;
        RECT 30.200 26.800 30.600 27.200 ;
        RECT 33.400 26.800 33.800 27.200 ;
        RECT 26.200 25.800 26.600 26.200 ;
        RECT 28.600 25.800 29.000 26.200 ;
        RECT 26.200 25.200 26.500 25.800 ;
        RECT 28.600 25.200 28.900 25.800 ;
        RECT 26.200 25.100 26.600 25.200 ;
        RECT 27.000 25.100 27.400 25.200 ;
        RECT 26.200 24.800 27.400 25.100 ;
        RECT 28.600 24.800 29.000 25.200 ;
        RECT 23.000 18.800 23.400 19.200 ;
        RECT 23.800 18.800 24.200 19.200 ;
        RECT 29.400 18.200 29.700 26.800 ;
        RECT 30.200 26.200 30.500 26.800 ;
        RECT 30.200 25.800 30.600 26.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 19.000 12.800 19.400 13.200 ;
        RECT 11.800 9.100 12.200 9.200 ;
        RECT 12.600 9.100 13.000 9.200 ;
        RECT 11.800 8.800 13.000 9.100 ;
        RECT 14.200 8.800 14.600 9.200 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 15.000 7.800 15.400 8.200 ;
        RECT 15.000 7.200 15.300 7.800 ;
        RECT 15.000 6.800 15.400 7.200 ;
        RECT 18.200 6.100 18.500 8.800 ;
        RECT 19.000 7.200 19.300 12.800 ;
        RECT 19.800 12.100 20.200 17.900 ;
        RECT 21.400 15.800 21.800 16.200 ;
        RECT 21.400 13.200 21.700 15.800 ;
        RECT 21.400 12.800 21.800 13.200 ;
        RECT 24.600 13.100 25.000 15.900 ;
        RECT 21.400 9.200 21.700 12.800 ;
        RECT 26.200 12.100 26.600 17.900 ;
        RECT 29.400 17.800 29.800 18.200 ;
        RECT 29.400 16.200 29.700 17.800 ;
        RECT 29.400 15.800 29.800 16.200 ;
        RECT 30.200 15.200 30.500 25.800 ;
        RECT 40.600 19.200 40.900 38.800 ;
        RECT 47.000 38.200 47.300 46.800 ;
        RECT 47.800 46.200 48.100 46.800 ;
        RECT 47.800 45.800 48.200 46.200 ;
        RECT 48.600 46.100 49.000 46.200 ;
        RECT 49.400 46.100 49.800 46.200 ;
        RECT 48.600 45.800 49.800 46.100 ;
        RECT 50.200 45.200 50.500 46.800 ;
        RECT 50.200 44.800 50.600 45.200 ;
        RECT 52.600 44.200 52.900 53.800 ;
        RECT 62.200 53.100 62.600 55.900 ;
        RECT 56.600 51.800 57.000 52.200 ;
        RECT 63.800 52.100 64.200 57.900 ;
        RECT 65.400 57.200 65.700 66.800 ;
        RECT 67.800 66.200 68.100 71.800 ;
        RECT 68.600 68.800 69.000 69.200 ;
        RECT 68.600 66.200 68.900 68.800 ;
        RECT 71.000 66.200 71.300 71.800 ;
        RECT 72.600 67.200 72.900 72.800 ;
        RECT 73.400 72.100 73.800 77.900 ;
        RECT 74.200 75.800 74.600 76.200 ;
        RECT 74.200 75.200 74.500 75.800 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 75.000 74.800 75.400 75.200 ;
        RECT 75.000 74.200 75.300 74.800 ;
        RECT 75.800 74.200 76.100 84.800 ;
        RECT 77.400 84.200 77.700 90.800 ;
        RECT 79.000 89.100 79.400 89.200 ;
        RECT 79.800 89.100 80.200 89.200 ;
        RECT 79.000 88.800 80.200 89.100 ;
        RECT 77.400 83.800 77.800 84.200 ;
        RECT 76.600 81.800 77.000 82.200 ;
        RECT 79.000 81.800 79.400 82.200 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 75.800 73.800 76.200 74.200 ;
        RECT 72.600 66.800 73.000 67.200 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 68.600 65.800 69.000 66.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 65.400 56.800 65.800 57.200 ;
        RECT 64.600 54.700 65.000 55.100 ;
        RECT 64.600 54.200 64.900 54.700 ;
        RECT 66.200 54.200 66.500 65.800 ;
        RECT 67.000 64.800 67.400 65.200 ;
        RECT 67.000 64.200 67.300 64.800 ;
        RECT 67.000 63.800 67.400 64.200 ;
        RECT 71.000 63.800 71.400 64.200 ;
        RECT 70.200 61.800 70.600 62.200 ;
        RECT 70.200 61.200 70.500 61.800 ;
        RECT 70.200 60.800 70.600 61.200 ;
        RECT 71.000 59.200 71.300 63.800 ;
        RECT 72.600 60.200 72.900 66.800 ;
        RECT 75.000 66.200 75.300 66.800 ;
        RECT 73.400 65.800 73.800 66.200 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 73.400 65.200 73.700 65.800 ;
        RECT 73.400 64.800 73.800 65.200 ;
        RECT 75.000 65.100 75.400 65.200 ;
        RECT 75.800 65.100 76.200 65.200 ;
        RECT 75.000 64.800 76.200 65.100 ;
        RECT 76.600 63.200 76.900 81.800 ;
        RECT 78.200 72.100 78.600 77.900 ;
        RECT 77.400 67.800 77.800 68.200 ;
        RECT 77.400 67.200 77.700 67.800 ;
        RECT 77.400 66.800 77.800 67.200 ;
        RECT 78.200 65.100 78.600 67.900 ;
        RECT 76.600 62.800 77.000 63.200 ;
        RECT 79.000 60.200 79.300 81.800 ;
        RECT 79.800 73.100 80.200 75.900 ;
        RECT 80.600 75.200 80.900 93.800 ;
        RECT 82.200 92.100 82.600 97.900 ;
        RECT 83.800 96.800 84.200 97.200 ;
        RECT 81.400 83.100 81.800 88.900 ;
        RECT 83.000 87.800 83.400 88.200 ;
        RECT 83.000 86.200 83.300 87.800 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 83.000 85.800 83.400 86.200 ;
        RECT 82.200 77.200 82.500 85.800 ;
        RECT 82.200 76.800 82.600 77.200 ;
        RECT 82.200 76.200 82.500 76.800 ;
        RECT 82.200 75.800 82.600 76.200 ;
        RECT 83.000 75.200 83.300 85.800 ;
        RECT 83.800 76.200 84.100 96.800 ;
        RECT 85.400 95.800 85.800 96.200 ;
        RECT 85.400 95.200 85.700 95.800 ;
        RECT 85.400 94.800 85.800 95.200 ;
        RECT 85.400 93.800 85.800 94.200 ;
        RECT 85.400 88.200 85.700 93.800 ;
        RECT 87.000 92.100 87.400 97.900 ;
        RECT 87.800 94.200 88.100 106.800 ;
        RECT 88.600 105.100 89.000 107.900 ;
        RECT 90.200 103.100 90.600 108.900 ;
        RECT 90.200 98.800 90.600 99.200 ;
        RECT 87.800 93.800 88.200 94.200 ;
        RECT 88.600 93.100 89.000 95.900 ;
        RECT 89.400 94.800 89.800 95.200 ;
        RECT 89.400 94.200 89.700 94.800 ;
        RECT 89.400 93.800 89.800 94.200 ;
        RECT 85.400 87.800 85.800 88.200 ;
        RECT 85.400 85.900 85.800 86.300 ;
        RECT 85.400 85.200 85.700 85.900 ;
        RECT 85.400 84.800 85.800 85.200 ;
        RECT 86.200 83.100 86.600 88.900 ;
        RECT 87.800 85.100 88.200 87.900 ;
        RECT 90.200 87.200 90.500 98.800 ;
        RECT 91.000 97.200 91.300 141.800 ;
        RECT 91.800 124.200 92.100 143.800 ;
        RECT 92.600 143.200 92.900 144.800 ;
        RECT 94.200 144.200 94.500 152.800 ;
        RECT 95.000 152.100 95.400 157.900 ;
        RECT 98.200 157.800 98.600 158.200 ;
        RECT 99.000 157.800 99.400 158.200 ;
        RECT 95.800 156.800 96.200 157.200 ;
        RECT 95.800 156.200 96.100 156.800 ;
        RECT 98.200 156.200 98.500 157.800 ;
        RECT 99.800 157.200 100.100 161.800 ;
        RECT 99.800 156.800 100.200 157.200 ;
        RECT 100.600 156.200 100.900 161.800 ;
        RECT 101.400 160.200 101.700 165.800 ;
        RECT 102.200 164.800 102.600 165.200 ;
        RECT 102.200 164.200 102.500 164.800 ;
        RECT 102.200 163.800 102.600 164.200 ;
        RECT 103.000 160.200 103.300 171.800 ;
        RECT 103.800 167.200 104.100 172.800 ;
        RECT 104.600 170.200 104.900 174.800 ;
        RECT 104.600 169.800 105.000 170.200 ;
        RECT 106.200 169.200 106.500 175.800 ;
        RECT 106.200 168.800 106.600 169.200 ;
        RECT 103.800 166.800 104.200 167.200 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 104.600 166.200 104.900 166.800 ;
        RECT 104.600 165.800 105.000 166.200 ;
        RECT 106.200 165.100 106.600 167.900 ;
        RECT 101.400 159.800 101.800 160.200 ;
        RECT 103.000 159.800 103.400 160.200 ;
        RECT 95.800 155.800 96.200 156.200 ;
        RECT 98.200 155.800 98.600 156.200 ;
        RECT 100.600 155.800 101.000 156.200 ;
        RECT 98.200 154.800 98.600 155.200 ;
        RECT 100.600 155.100 101.000 155.200 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 100.600 154.800 101.800 155.100 ;
        RECT 102.200 154.800 102.600 155.200 ;
        RECT 98.200 154.200 98.500 154.800 ;
        RECT 102.200 154.200 102.500 154.800 ;
        RECT 103.000 154.200 103.300 159.800 ;
        RECT 103.800 156.800 104.200 157.200 ;
        RECT 103.800 156.200 104.100 156.800 ;
        RECT 103.800 155.800 104.200 156.200 ;
        RECT 98.200 153.800 98.600 154.200 ;
        RECT 99.800 153.800 100.200 154.200 ;
        RECT 102.200 153.800 102.600 154.200 ;
        RECT 103.000 153.800 103.400 154.200 ;
        RECT 105.400 153.800 105.800 154.200 ;
        RECT 99.800 153.200 100.100 153.800 ;
        RECT 105.400 153.200 105.700 153.800 ;
        RECT 99.800 152.800 100.200 153.200 ;
        RECT 100.600 152.800 101.000 153.200 ;
        RECT 105.400 152.800 105.800 153.200 ;
        RECT 106.200 153.100 106.600 155.900 ;
        RECT 96.600 149.800 97.000 150.200 ;
        RECT 96.600 149.200 96.900 149.800 ;
        RECT 100.600 149.200 100.900 152.800 ;
        RECT 104.600 151.800 105.000 152.200 ;
        RECT 104.600 149.200 104.900 151.800 ;
        RECT 106.200 150.800 106.600 151.200 ;
        RECT 106.200 149.200 106.500 150.800 ;
        RECT 96.600 148.800 97.000 149.200 ;
        RECT 100.600 148.800 101.000 149.200 ;
        RECT 104.600 148.800 105.000 149.200 ;
        RECT 106.200 148.800 106.600 149.200 ;
        RECT 103.000 147.800 103.400 148.200 ;
        RECT 103.000 147.200 103.300 147.800 ;
        RECT 107.000 147.200 107.300 177.800 ;
        RECT 108.600 175.200 108.900 177.800 ;
        RECT 110.200 175.200 110.500 186.800 ;
        RECT 111.800 185.800 112.200 186.200 ;
        RECT 116.600 185.800 117.000 186.200 ;
        RECT 111.800 179.200 112.100 185.800 ;
        RECT 116.600 180.200 116.900 185.800 ;
        RECT 116.600 179.800 117.000 180.200 ;
        RECT 111.800 178.800 112.200 179.200 ;
        RECT 115.800 176.800 116.200 177.200 ;
        RECT 115.800 176.200 116.100 176.800 ;
        RECT 112.600 176.100 113.000 176.200 ;
        RECT 113.400 176.100 113.800 176.200 ;
        RECT 112.600 175.800 113.800 176.100 ;
        RECT 114.200 176.100 114.600 176.200 ;
        RECT 115.000 176.100 115.400 176.200 ;
        RECT 114.200 175.800 115.400 176.100 ;
        RECT 115.800 175.800 116.200 176.200 ;
        RECT 108.600 174.800 109.000 175.200 ;
        RECT 110.200 174.800 110.600 175.200 ;
        RECT 111.000 174.800 111.400 175.200 ;
        RECT 112.600 174.800 113.000 175.200 ;
        RECT 114.200 174.800 114.600 175.200 ;
        RECT 110.200 174.200 110.500 174.800 ;
        RECT 107.800 174.100 108.200 174.200 ;
        RECT 107.800 173.800 108.900 174.100 ;
        RECT 107.800 163.100 108.200 168.900 ;
        RECT 108.600 166.300 108.900 173.800 ;
        RECT 109.400 173.800 109.800 174.200 ;
        RECT 110.200 173.800 110.600 174.200 ;
        RECT 108.600 165.900 109.000 166.300 ;
        RECT 108.600 165.800 108.900 165.900 ;
        RECT 109.400 162.200 109.700 173.800 ;
        RECT 111.000 170.200 111.300 174.800 ;
        RECT 112.600 174.200 112.900 174.800 ;
        RECT 112.600 173.800 113.000 174.200 ;
        RECT 113.400 173.800 113.800 174.200 ;
        RECT 113.400 171.200 113.700 173.800 ;
        RECT 114.200 173.200 114.500 174.800 ;
        RECT 114.200 172.800 114.600 173.200 ;
        RECT 116.600 173.100 117.000 175.900 ;
        RECT 117.400 173.200 117.700 191.800 ;
        RECT 118.200 190.200 118.500 193.800 ;
        RECT 119.000 192.100 119.400 197.900 ;
        RECT 121.400 196.800 121.800 197.200 ;
        RECT 121.400 195.200 121.700 196.800 ;
        RECT 120.600 194.800 121.000 195.200 ;
        RECT 121.400 194.800 121.800 195.200 ;
        RECT 119.800 192.800 120.200 193.200 ;
        RECT 118.200 189.800 118.600 190.200 ;
        RECT 119.000 186.800 119.400 187.200 ;
        RECT 119.000 186.200 119.300 186.800 ;
        RECT 118.200 185.800 118.600 186.200 ;
        RECT 119.000 185.800 119.400 186.200 ;
        RECT 118.200 185.200 118.500 185.800 ;
        RECT 118.200 184.800 118.600 185.200 ;
        RECT 117.400 172.800 117.800 173.200 ;
        RECT 118.200 172.100 118.600 177.900 ;
        RECT 119.000 174.700 119.400 175.100 ;
        RECT 119.000 174.200 119.300 174.700 ;
        RECT 119.800 174.200 120.100 192.800 ;
        RECT 120.600 186.200 120.900 194.800 ;
        RECT 123.800 192.100 124.200 197.900 ;
        RECT 126.200 196.800 126.600 197.200 ;
        RECT 127.000 197.100 127.400 197.200 ;
        RECT 127.800 197.100 128.200 197.200 ;
        RECT 127.000 196.800 128.200 197.100 ;
        RECT 126.200 196.200 126.500 196.800 ;
        RECT 126.200 195.800 126.600 196.200 ;
        RECT 127.000 195.100 127.400 195.200 ;
        RECT 127.800 195.100 128.200 195.200 ;
        RECT 127.000 194.800 128.200 195.100 ;
        RECT 127.000 193.800 127.400 194.200 ;
        RECT 127.000 193.200 127.300 193.800 ;
        RECT 127.000 192.800 127.400 193.200 ;
        RECT 121.400 189.800 121.800 190.200 ;
        RECT 121.400 187.200 121.700 189.800 ;
        RECT 121.400 186.800 121.800 187.200 ;
        RECT 120.600 185.800 121.000 186.200 ;
        RECT 119.000 173.800 119.400 174.200 ;
        RECT 119.800 173.800 120.200 174.200 ;
        RECT 119.000 172.800 119.400 173.200 ;
        RECT 113.400 170.800 113.800 171.200 ;
        RECT 111.000 169.800 111.400 170.200 ;
        RECT 109.400 161.800 109.800 162.200 ;
        RECT 107.800 152.100 108.200 157.900 ;
        RECT 108.600 155.800 109.000 156.200 ;
        RECT 109.400 155.800 109.800 156.200 ;
        RECT 108.600 154.200 108.900 155.800 ;
        RECT 109.400 155.200 109.700 155.800 ;
        RECT 109.400 154.800 109.800 155.200 ;
        RECT 111.000 154.200 111.300 169.800 ;
        RECT 115.000 169.100 115.400 169.200 ;
        RECT 115.800 169.100 116.200 169.200 ;
        RECT 111.800 165.800 112.200 166.200 ;
        RECT 111.800 155.200 112.100 165.800 ;
        RECT 112.600 163.100 113.000 168.900 ;
        RECT 115.000 168.800 116.200 169.100 ;
        RECT 113.400 167.800 113.800 168.200 ;
        RECT 111.800 154.800 112.200 155.200 ;
        RECT 111.800 154.200 112.100 154.800 ;
        RECT 108.600 153.800 109.000 154.200 ;
        RECT 111.000 153.800 111.400 154.200 ;
        RECT 111.800 153.800 112.200 154.200 ;
        RECT 112.600 152.100 113.000 157.900 ;
        RECT 113.400 149.200 113.700 167.800 ;
        RECT 119.000 166.200 119.300 172.800 ;
        RECT 114.200 165.800 114.600 166.200 ;
        RECT 115.000 166.100 115.400 166.200 ;
        RECT 115.800 166.100 116.200 166.200 ;
        RECT 115.000 165.800 116.200 166.100 ;
        RECT 116.600 165.800 117.000 166.200 ;
        RECT 119.000 165.800 119.400 166.200 ;
        RECT 114.200 149.200 114.500 165.800 ;
        RECT 116.600 165.200 116.900 165.800 ;
        RECT 116.600 164.800 117.000 165.200 ;
        RECT 115.800 153.100 116.200 155.900 ;
        RECT 116.600 154.800 117.000 155.200 ;
        RECT 116.600 154.200 116.900 154.800 ;
        RECT 116.600 153.800 117.000 154.200 ;
        RECT 115.000 152.100 115.400 152.200 ;
        RECT 115.800 152.100 116.200 152.200 ;
        RECT 117.400 152.100 117.800 157.900 ;
        RECT 119.000 154.800 119.400 155.200 ;
        RECT 119.000 154.200 119.300 154.800 ;
        RECT 119.800 154.200 120.100 173.800 ;
        RECT 120.600 171.200 120.900 185.800 ;
        RECT 120.600 170.800 121.000 171.200 ;
        RECT 121.400 165.200 121.700 186.800 ;
        RECT 122.200 184.800 122.600 185.200 ;
        RECT 122.200 184.200 122.500 184.800 ;
        RECT 122.200 183.800 122.600 184.200 ;
        RECT 124.600 183.100 125.000 188.900 ;
        RECT 127.000 187.200 127.300 192.800 ;
        RECT 128.600 188.200 128.900 200.800 ;
        RECT 130.200 196.800 130.600 197.200 ;
        RECT 130.200 196.200 130.500 196.800 ;
        RECT 130.200 195.800 130.600 196.200 ;
        RECT 128.600 187.800 129.000 188.200 ;
        RECT 127.000 186.800 127.400 187.200 ;
        RECT 126.200 186.100 126.600 186.200 ;
        RECT 127.000 186.100 127.400 186.200 ;
        RECT 126.200 185.800 127.400 186.100 ;
        RECT 129.400 183.100 129.800 188.900 ;
        RECT 123.000 172.100 123.400 177.900 ;
        RECT 124.600 177.100 125.000 177.200 ;
        RECT 125.400 177.100 125.800 177.200 ;
        RECT 124.600 176.800 125.800 177.100 ;
        RECT 130.200 176.100 130.500 195.800 ;
        RECT 131.800 194.800 132.200 195.200 ;
        RECT 131.800 191.200 132.100 194.800 ;
        RECT 132.600 193.800 133.000 194.200 ;
        RECT 131.800 190.800 132.200 191.200 ;
        RECT 132.600 189.200 132.900 193.800 ;
        RECT 132.600 188.800 133.000 189.200 ;
        RECT 131.000 185.100 131.400 187.900 ;
        RECT 131.800 186.800 132.200 187.200 ;
        RECT 131.800 184.100 132.100 186.800 ;
        RECT 129.400 175.800 130.500 176.100 ;
        RECT 131.000 183.800 132.100 184.100 ;
        RECT 131.000 176.200 131.300 183.800 ;
        RECT 131.000 175.800 131.400 176.200 ;
        RECT 129.400 175.200 129.700 175.800 ;
        RECT 129.400 174.800 129.800 175.200 ;
        RECT 130.200 174.800 130.600 175.200 ;
        RECT 130.200 174.200 130.500 174.800 ;
        RECT 130.200 173.800 130.600 174.200 ;
        RECT 127.800 171.800 128.200 172.200 ;
        RECT 127.800 167.200 128.100 171.800 ;
        RECT 128.600 169.800 129.000 170.200 ;
        RECT 123.800 166.800 124.200 167.200 ;
        RECT 127.800 166.800 128.200 167.200 ;
        RECT 123.800 166.200 124.100 166.800 ;
        RECT 128.600 166.200 128.900 169.800 ;
        RECT 130.200 168.800 130.600 169.200 ;
        RECT 129.400 166.800 129.800 167.200 ;
        RECT 129.400 166.200 129.700 166.800 ;
        RECT 130.200 166.200 130.500 168.800 ;
        RECT 131.000 168.200 131.300 175.800 ;
        RECT 133.400 175.200 133.700 203.800 ;
        RECT 139.000 202.800 139.400 203.200 ;
        RECT 143.800 203.100 144.200 208.900 ;
        RECT 145.400 206.100 145.800 206.200 ;
        RECT 146.200 206.100 146.600 206.200 ;
        RECT 145.400 205.800 146.600 206.100 ;
        RECT 148.600 203.100 149.000 208.900 ;
        RECT 151.000 208.800 152.200 209.100 ;
        RECT 156.600 208.800 157.000 209.200 ;
        RECT 156.600 207.200 156.900 208.800 ;
        RECT 151.800 206.800 152.200 207.200 ;
        RECT 153.400 206.800 153.800 207.200 ;
        RECT 156.600 206.800 157.000 207.200 ;
        RECT 149.400 203.800 149.800 204.200 ;
        RECT 139.000 202.200 139.300 202.800 ;
        RECT 134.200 201.800 134.600 202.200 ;
        RECT 139.000 202.100 139.400 202.200 ;
        RECT 139.800 202.100 140.200 202.200 ;
        RECT 139.000 201.800 140.200 202.100 ;
        RECT 134.200 198.200 134.500 201.800 ;
        RECT 135.000 199.800 135.400 200.200 ;
        RECT 134.200 197.800 134.600 198.200 ;
        RECT 134.200 195.200 134.500 197.800 ;
        RECT 134.200 194.800 134.600 195.200 ;
        RECT 135.000 186.200 135.300 199.800 ;
        RECT 135.800 196.800 136.200 197.200 ;
        RECT 137.400 196.800 137.800 197.200 ;
        RECT 140.600 197.100 141.000 197.200 ;
        RECT 141.400 197.100 141.800 197.200 ;
        RECT 140.600 196.800 141.800 197.100 ;
        RECT 135.800 196.200 136.100 196.800 ;
        RECT 135.800 195.800 136.200 196.200 ;
        RECT 137.400 186.200 137.700 196.800 ;
        RECT 138.200 196.100 138.600 196.200 ;
        RECT 139.000 196.100 139.400 196.200 ;
        RECT 138.200 195.800 139.400 196.100 ;
        RECT 138.200 195.100 138.600 195.200 ;
        RECT 139.000 195.100 139.400 195.200 ;
        RECT 138.200 194.800 139.400 195.100 ;
        RECT 139.000 193.800 139.400 194.200 ;
        RECT 139.000 193.200 139.300 193.800 ;
        RECT 139.000 192.800 139.400 193.200 ;
        RECT 139.000 189.100 139.300 192.800 ;
        RECT 143.800 192.100 144.200 197.900 ;
        RECT 147.000 195.800 147.400 196.200 ;
        RECT 147.000 195.200 147.300 195.800 ;
        RECT 147.000 194.800 147.400 195.200 ;
        RECT 147.800 194.800 148.200 195.200 ;
        RECT 138.200 188.800 139.300 189.100 ;
        RECT 141.400 190.800 141.800 191.200 ;
        RECT 143.800 190.800 144.200 191.200 ;
        RECT 135.000 185.800 135.400 186.200 ;
        RECT 137.400 185.800 137.800 186.200 ;
        RECT 134.200 184.800 134.600 185.200 ;
        RECT 133.400 174.800 133.800 175.200 ;
        RECT 131.800 173.800 132.200 174.200 ;
        RECT 132.600 173.800 133.000 174.200 ;
        RECT 134.200 174.100 134.500 184.800 ;
        RECT 133.400 173.800 134.500 174.100 ;
        RECT 135.800 181.800 136.200 182.200 ;
        RECT 131.800 173.200 132.100 173.800 ;
        RECT 131.800 172.800 132.200 173.200 ;
        RECT 131.000 167.800 131.400 168.200 ;
        RECT 123.800 165.800 124.200 166.200 ;
        RECT 124.600 165.800 125.000 166.200 ;
        RECT 126.200 165.800 126.600 166.200 ;
        RECT 128.600 165.800 129.000 166.200 ;
        RECT 129.400 165.800 129.800 166.200 ;
        RECT 130.200 165.800 130.600 166.200 ;
        RECT 124.600 165.200 124.900 165.800 ;
        RECT 126.200 165.200 126.500 165.800 ;
        RECT 121.400 164.800 121.800 165.200 ;
        RECT 123.800 164.800 124.200 165.200 ;
        RECT 124.600 164.800 125.000 165.200 ;
        RECT 126.200 164.800 126.600 165.200 ;
        RECT 131.800 164.800 132.200 165.200 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 120.600 155.800 121.000 156.200 ;
        RECT 121.400 155.800 121.800 156.200 ;
        RECT 119.000 153.800 119.400 154.200 ;
        RECT 119.800 153.800 120.200 154.200 ;
        RECT 115.000 151.800 116.200 152.100 ;
        RECT 120.600 149.200 120.900 155.800 ;
        RECT 121.400 155.200 121.700 155.800 ;
        RECT 121.400 154.800 121.800 155.200 ;
        RECT 122.200 152.100 122.600 157.900 ;
        RECT 123.000 155.200 123.300 161.800 ;
        RECT 123.800 160.200 124.100 164.800 ;
        RECT 131.800 164.200 132.100 164.800 ;
        RECT 131.800 163.800 132.200 164.200 ;
        RECT 129.400 162.800 129.800 163.200 ;
        RECT 127.800 161.800 128.200 162.200 ;
        RECT 127.000 160.800 127.400 161.200 ;
        RECT 123.800 159.800 124.200 160.200 ;
        RECT 123.000 154.800 123.400 155.200 ;
        RECT 123.000 151.800 123.400 152.200 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 114.200 148.800 114.600 149.200 ;
        RECT 120.600 148.800 121.000 149.200 ;
        RECT 114.200 148.200 114.500 148.800 ;
        RECT 110.200 147.800 110.600 148.200 ;
        RECT 114.200 147.800 114.600 148.200 ;
        RECT 117.400 147.800 117.800 148.200 ;
        RECT 118.200 147.800 118.600 148.200 ;
        RECT 95.800 147.100 96.200 147.200 ;
        RECT 96.600 147.100 97.000 147.200 ;
        RECT 95.800 146.800 97.000 147.100 ;
        RECT 103.000 146.800 103.400 147.200 ;
        RECT 107.000 146.800 107.400 147.200 ;
        RECT 99.000 146.100 99.400 146.200 ;
        RECT 99.000 145.800 100.100 146.100 ;
        RECT 99.800 145.200 100.100 145.800 ;
        RECT 101.400 145.800 101.800 146.200 ;
        RECT 102.200 145.800 102.600 146.200 ;
        RECT 99.000 144.800 99.400 145.200 ;
        RECT 99.800 144.800 100.200 145.200 ;
        RECT 94.200 143.800 94.600 144.200 ;
        RECT 92.600 142.800 93.000 143.200 ;
        RECT 92.600 140.200 92.900 142.800 ;
        RECT 93.400 141.800 93.800 142.200 ;
        RECT 92.600 139.800 93.000 140.200 ;
        RECT 93.400 139.200 93.700 141.800 ;
        RECT 94.200 139.200 94.500 143.800 ;
        RECT 99.000 143.200 99.300 144.800 ;
        RECT 99.800 143.800 100.200 144.200 ;
        RECT 99.800 143.200 100.100 143.800 ;
        RECT 99.000 142.800 99.400 143.200 ;
        RECT 99.800 142.800 100.200 143.200 ;
        RECT 97.400 141.800 97.800 142.200 ;
        RECT 99.000 142.100 99.300 142.800 ;
        RECT 99.000 141.800 100.100 142.100 ;
        RECT 93.400 138.800 93.800 139.200 ;
        RECT 94.200 138.800 94.600 139.200 ;
        RECT 93.400 132.100 93.800 137.900 ;
        RECT 94.200 137.200 94.500 138.800 ;
        RECT 94.200 136.800 94.600 137.200 ;
        RECT 94.200 135.800 94.600 136.200 ;
        RECT 94.200 129.200 94.500 135.800 ;
        RECT 96.600 134.800 97.000 135.200 ;
        RECT 96.600 134.200 96.900 134.800 ;
        RECT 95.000 133.800 95.400 134.200 ;
        RECT 96.600 133.800 97.000 134.200 ;
        RECT 95.000 131.200 95.300 133.800 ;
        RECT 97.400 133.200 97.700 141.800 ;
        RECT 99.800 139.200 100.100 141.800 ;
        RECT 100.600 141.800 101.000 142.200 ;
        RECT 99.800 138.800 100.200 139.200 ;
        RECT 98.200 135.100 98.600 135.200 ;
        RECT 99.000 135.100 99.400 135.200 ;
        RECT 98.200 134.800 99.400 135.100 ;
        RECT 96.600 133.100 97.000 133.200 ;
        RECT 97.400 133.100 97.800 133.200 ;
        RECT 96.600 132.800 97.800 133.100 ;
        RECT 95.800 131.800 96.200 132.200 ;
        RECT 95.000 130.800 95.400 131.200 ;
        RECT 94.200 128.800 94.600 129.200 ;
        RECT 95.000 125.200 95.300 130.800 ;
        RECT 95.000 124.800 95.400 125.200 ;
        RECT 95.800 125.100 96.100 131.800 ;
        RECT 99.000 128.800 99.400 129.200 ;
        RECT 99.000 128.200 99.300 128.800 ;
        RECT 99.000 127.800 99.400 128.200 ;
        RECT 96.600 126.800 97.000 127.200 ;
        RECT 98.200 127.100 98.600 127.200 ;
        RECT 99.000 127.100 99.400 127.200 ;
        RECT 98.200 126.800 99.400 127.100 ;
        RECT 96.600 125.200 96.900 126.800 ;
        RECT 100.600 126.200 100.900 141.800 ;
        RECT 101.400 137.200 101.700 145.800 ;
        RECT 102.200 145.200 102.500 145.800 ;
        RECT 102.200 144.800 102.600 145.200 ;
        RECT 103.000 144.200 103.300 146.800 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 104.600 146.100 105.000 146.200 ;
        RECT 103.800 145.800 105.000 146.100 ;
        RECT 109.400 145.800 109.800 146.200 ;
        RECT 109.400 145.200 109.700 145.800 ;
        RECT 104.600 144.800 105.000 145.200 ;
        RECT 109.400 144.800 109.800 145.200 ;
        RECT 103.000 143.800 103.400 144.200 ;
        RECT 103.800 142.800 104.200 143.200 ;
        RECT 103.800 137.200 104.100 142.800 ;
        RECT 101.400 136.800 101.800 137.200 ;
        RECT 103.800 136.800 104.200 137.200 ;
        RECT 102.200 135.800 102.600 136.200 ;
        RECT 103.000 135.800 103.400 136.200 ;
        RECT 102.200 135.200 102.500 135.800 ;
        RECT 103.000 135.200 103.300 135.800 ;
        RECT 104.600 135.200 104.900 144.800 ;
        RECT 105.400 143.800 105.800 144.200 ;
        RECT 109.400 143.800 109.800 144.200 ;
        RECT 105.400 142.200 105.700 143.800 ;
        RECT 105.400 141.800 105.800 142.200 ;
        RECT 105.400 137.200 105.700 141.800 ;
        RECT 105.400 136.800 105.800 137.200 ;
        RECT 105.400 135.800 105.800 136.200 ;
        RECT 106.200 135.800 106.600 136.200 ;
        RECT 105.400 135.200 105.700 135.800 ;
        RECT 106.200 135.200 106.500 135.800 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 102.200 134.800 102.600 135.200 ;
        RECT 103.000 134.800 103.400 135.200 ;
        RECT 104.600 134.800 105.000 135.200 ;
        RECT 105.400 134.800 105.800 135.200 ;
        RECT 106.200 134.800 106.600 135.200 ;
        RECT 108.600 134.800 109.000 135.200 ;
        RECT 101.400 134.200 101.700 134.800 ;
        RECT 101.400 133.800 101.800 134.200 ;
        RECT 101.400 126.800 101.800 127.200 ;
        RECT 101.400 126.200 101.700 126.800 ;
        RECT 97.400 125.800 97.800 126.200 ;
        RECT 100.600 125.800 101.000 126.200 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 96.600 125.100 97.000 125.200 ;
        RECT 95.800 124.800 97.000 125.100 ;
        RECT 91.800 123.800 92.200 124.200 ;
        RECT 92.600 121.800 93.000 122.200 ;
        RECT 92.600 120.200 92.900 121.800 ;
        RECT 97.400 121.200 97.700 125.800 ;
        RECT 102.200 125.200 102.500 134.800 ;
        RECT 103.000 127.200 103.300 134.800 ;
        RECT 104.600 131.800 105.000 132.200 ;
        RECT 103.000 126.800 103.400 127.200 ;
        RECT 103.800 126.800 104.200 127.200 ;
        RECT 103.800 126.200 104.100 126.800 ;
        RECT 103.800 125.800 104.200 126.200 ;
        RECT 99.800 124.800 100.200 125.200 ;
        RECT 100.600 124.800 101.000 125.200 ;
        RECT 102.200 124.800 102.600 125.200 ;
        RECT 103.800 124.800 104.200 125.200 ;
        RECT 97.400 120.800 97.800 121.200 ;
        RECT 92.600 119.800 93.000 120.200 ;
        RECT 91.800 113.100 92.200 115.900 ;
        RECT 92.600 115.800 93.000 116.200 ;
        RECT 95.800 115.800 96.200 116.200 ;
        RECT 92.600 114.200 92.900 115.800 ;
        RECT 92.600 113.800 93.000 114.200 ;
        RECT 95.800 113.200 96.100 115.800 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 98.200 114.800 98.600 115.200 ;
        RECT 96.600 114.200 96.900 114.800 ;
        RECT 96.600 113.800 97.000 114.200 ;
        RECT 98.200 113.200 98.500 114.800 ;
        RECT 99.800 114.200 100.100 124.800 ;
        RECT 100.600 124.200 100.900 124.800 ;
        RECT 103.800 124.200 104.100 124.800 ;
        RECT 104.600 124.200 104.900 131.800 ;
        RECT 105.400 125.200 105.700 134.800 ;
        RECT 108.600 134.200 108.900 134.800 ;
        RECT 108.600 133.800 109.000 134.200 ;
        RECT 107.000 132.800 107.400 133.200 ;
        RECT 106.200 127.800 106.600 128.200 ;
        RECT 106.200 127.200 106.500 127.800 ;
        RECT 106.200 126.800 106.600 127.200 ;
        RECT 107.000 126.200 107.300 132.800 ;
        RECT 107.800 131.800 108.200 132.200 ;
        RECT 107.000 125.800 107.400 126.200 ;
        RECT 105.400 124.800 105.800 125.200 ;
        RECT 100.600 123.800 101.000 124.200 ;
        RECT 103.000 124.100 103.400 124.200 ;
        RECT 103.800 124.100 104.200 124.200 ;
        RECT 103.000 123.800 104.200 124.100 ;
        RECT 104.600 123.800 105.000 124.200 ;
        RECT 101.400 121.800 101.800 122.200 ;
        RECT 104.600 121.800 105.000 122.200 ;
        RECT 101.400 118.200 101.700 121.800 ;
        RECT 102.200 119.800 102.600 120.200 ;
        RECT 101.400 117.800 101.800 118.200 ;
        RECT 102.200 117.200 102.500 119.800 ;
        RECT 102.200 116.800 102.600 117.200 ;
        RECT 103.800 116.800 104.200 117.200 ;
        RECT 103.800 116.200 104.100 116.800 ;
        RECT 104.600 116.200 104.900 121.800 ;
        RECT 101.400 116.100 101.800 116.200 ;
        RECT 102.200 116.100 102.600 116.200 ;
        RECT 101.400 115.800 102.600 116.100 ;
        RECT 103.800 115.800 104.200 116.200 ;
        RECT 104.600 115.800 105.000 116.200 ;
        RECT 105.400 115.800 105.800 116.200 ;
        RECT 105.400 115.200 105.700 115.800 ;
        RECT 103.000 115.100 103.400 115.200 ;
        RECT 103.800 115.100 104.200 115.200 ;
        RECT 103.000 114.800 104.200 115.100 ;
        RECT 105.400 114.800 105.800 115.200 ;
        RECT 99.000 113.800 99.400 114.200 ;
        RECT 99.800 113.800 100.200 114.200 ;
        RECT 103.800 114.100 104.200 114.200 ;
        RECT 103.800 113.800 104.900 114.100 ;
        RECT 95.800 112.800 96.200 113.200 ;
        RECT 98.200 112.800 98.600 113.200 ;
        RECT 94.200 107.800 94.600 108.200 ;
        RECT 94.200 107.200 94.500 107.800 ;
        RECT 94.200 106.800 94.600 107.200 ;
        RECT 91.800 105.800 92.200 106.200 ;
        RECT 91.800 105.200 92.100 105.800 ;
        RECT 91.800 104.800 92.200 105.200 ;
        RECT 94.200 102.800 94.600 103.200 ;
        RECT 95.000 103.100 95.400 108.900 ;
        RECT 94.200 97.200 94.500 102.800 ;
        RECT 95.000 101.800 95.400 102.200 ;
        RECT 95.000 99.200 95.300 101.800 ;
        RECT 95.000 98.800 95.400 99.200 ;
        RECT 95.800 98.200 96.100 112.800 ;
        RECT 99.000 111.200 99.300 113.800 ;
        RECT 100.600 112.100 101.000 112.200 ;
        RECT 101.400 112.100 101.800 112.200 ;
        RECT 100.600 111.800 101.800 112.100 ;
        RECT 99.000 110.800 99.400 111.200 ;
        RECT 97.400 109.100 97.800 109.200 ;
        RECT 98.200 109.100 98.600 109.200 ;
        RECT 97.400 108.800 98.600 109.100 ;
        RECT 99.000 108.200 99.300 110.800 ;
        RECT 103.000 108.800 103.400 109.200 ;
        RECT 99.000 107.800 99.400 108.200 ;
        RECT 103.000 107.200 103.300 108.800 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 103.000 106.800 103.400 107.200 ;
        RECT 98.200 106.200 98.500 106.800 ;
        RECT 98.200 105.800 98.600 106.200 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 99.800 106.100 100.200 106.200 ;
        RECT 99.000 105.800 100.200 106.100 ;
        RECT 99.000 105.100 99.400 105.200 ;
        RECT 99.800 105.100 100.200 105.200 ;
        RECT 99.000 104.800 100.200 105.100 ;
        RECT 101.400 105.100 101.800 105.200 ;
        RECT 102.200 105.100 102.600 105.200 ;
        RECT 103.800 105.100 104.200 107.900 ;
        RECT 101.400 104.800 102.600 105.100 ;
        RECT 100.600 101.800 101.000 102.200 ;
        RECT 97.400 99.800 97.800 100.200 ;
        RECT 97.400 99.200 97.700 99.800 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 95.800 97.800 96.200 98.200 ;
        RECT 100.600 97.200 100.900 101.800 ;
        RECT 104.600 99.200 104.900 113.800 ;
        RECT 105.400 110.200 105.700 114.800 ;
        RECT 106.200 112.800 106.600 113.200 ;
        RECT 107.000 113.100 107.300 125.800 ;
        RECT 107.800 121.200 108.100 131.800 ;
        RECT 109.400 128.200 109.700 143.800 ;
        RECT 108.600 127.800 109.000 128.200 ;
        RECT 109.400 127.800 109.800 128.200 ;
        RECT 108.600 127.200 108.900 127.800 ;
        RECT 109.400 127.200 109.700 127.800 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 108.600 125.800 109.000 126.200 ;
        RECT 108.600 122.200 108.900 125.800 ;
        RECT 110.200 124.200 110.500 147.800 ;
        RECT 117.400 147.200 117.700 147.800 ;
        RECT 118.200 147.200 118.500 147.800 ;
        RECT 123.000 147.200 123.300 151.800 ;
        RECT 123.800 149.200 124.100 159.800 ;
        RECT 124.600 152.100 125.000 152.200 ;
        RECT 125.400 152.100 125.800 152.200 ;
        RECT 124.600 151.800 125.800 152.100 ;
        RECT 126.200 151.800 126.600 152.200 ;
        RECT 123.800 148.800 124.200 149.200 ;
        RECT 126.200 147.200 126.500 151.800 ;
        RECT 116.600 146.800 117.000 147.200 ;
        RECT 117.400 146.800 117.800 147.200 ;
        RECT 118.200 147.100 118.600 147.200 ;
        RECT 119.000 147.100 119.400 147.200 ;
        RECT 118.200 146.800 119.400 147.100 ;
        RECT 123.000 146.800 123.400 147.200 ;
        RECT 125.400 146.800 125.800 147.200 ;
        RECT 126.200 146.800 126.600 147.200 ;
        RECT 127.000 147.100 127.300 160.800 ;
        RECT 127.800 156.100 128.100 161.800 ;
        RECT 129.400 159.200 129.700 162.800 ;
        RECT 132.600 162.200 132.900 173.800 ;
        RECT 133.400 166.200 133.700 173.800 ;
        RECT 135.000 171.800 135.400 172.200 ;
        RECT 135.000 170.200 135.300 171.800 ;
        RECT 135.000 169.800 135.400 170.200 ;
        RECT 135.800 167.200 136.100 181.800 ;
        RECT 136.600 177.800 137.000 178.200 ;
        RECT 136.600 175.200 136.900 177.800 ;
        RECT 138.200 175.200 138.500 188.800 ;
        RECT 140.600 187.800 141.000 188.200 ;
        RECT 140.600 187.200 140.900 187.800 ;
        RECT 140.600 186.800 141.000 187.200 ;
        RECT 141.400 186.200 141.700 190.800 ;
        RECT 143.800 187.200 144.100 190.800 ;
        RECT 147.000 189.800 147.400 190.200 ;
        RECT 147.000 187.200 147.300 189.800 ;
        RECT 143.800 186.800 144.200 187.200 ;
        RECT 147.000 186.800 147.400 187.200 ;
        RECT 147.800 186.200 148.100 194.800 ;
        RECT 148.600 192.100 149.000 197.900 ;
        RECT 149.400 194.200 149.700 203.800 ;
        RECT 151.800 196.200 152.100 206.800 ;
        RECT 153.400 206.200 153.700 206.800 ;
        RECT 152.600 205.800 153.000 206.200 ;
        RECT 153.400 205.800 153.800 206.200 ;
        RECT 152.600 205.200 152.900 205.800 ;
        RECT 152.600 204.800 153.000 205.200 ;
        RECT 155.000 204.800 155.400 205.200 ;
        RECT 149.400 193.800 149.800 194.200 ;
        RECT 149.400 188.200 149.700 193.800 ;
        RECT 150.200 193.100 150.600 195.900 ;
        RECT 151.800 195.800 152.200 196.200 ;
        RECT 151.800 195.200 152.100 195.800 ;
        RECT 151.800 194.800 152.200 195.200 ;
        RECT 151.000 191.800 151.400 192.200 ;
        RECT 153.400 192.100 153.800 197.900 ;
        RECT 149.400 187.800 149.800 188.200 ;
        RECT 149.400 186.800 149.800 187.200 ;
        RECT 149.400 186.200 149.700 186.800 ;
        RECT 139.000 186.100 139.400 186.200 ;
        RECT 139.800 186.100 140.200 186.200 ;
        RECT 139.000 185.800 140.200 186.100 ;
        RECT 141.400 185.800 141.800 186.200 ;
        RECT 144.600 185.800 145.000 186.200 ;
        RECT 147.000 185.800 147.400 186.200 ;
        RECT 147.800 185.800 148.200 186.200 ;
        RECT 149.400 185.800 149.800 186.200 ;
        RECT 143.000 183.800 143.400 184.200 ;
        RECT 141.400 181.800 141.800 182.200 ;
        RECT 141.400 176.200 141.700 181.800 ;
        RECT 143.000 179.200 143.300 183.800 ;
        RECT 144.600 179.200 144.900 185.800 ;
        RECT 147.000 185.200 147.300 185.800 ;
        RECT 145.400 185.100 145.800 185.200 ;
        RECT 146.200 185.100 146.600 185.200 ;
        RECT 145.400 184.800 146.600 185.100 ;
        RECT 147.000 184.800 147.400 185.200 ;
        RECT 148.600 185.100 149.000 185.200 ;
        RECT 149.400 185.100 149.800 185.200 ;
        RECT 150.200 185.100 150.600 187.900 ;
        RECT 151.000 186.200 151.300 191.800 ;
        RECT 151.000 185.800 151.400 186.200 ;
        RECT 148.600 184.800 149.800 185.100 ;
        RECT 146.200 184.200 146.500 184.800 ;
        RECT 146.200 183.800 146.600 184.200 ;
        RECT 143.000 178.800 143.400 179.200 ;
        RECT 144.600 178.800 145.000 179.200 ;
        RECT 143.000 178.200 143.300 178.800 ;
        RECT 143.000 177.800 143.400 178.200 ;
        RECT 141.400 175.800 141.800 176.200 ;
        RECT 142.200 175.800 142.600 176.200 ;
        RECT 142.200 175.200 142.500 175.800 ;
        RECT 136.600 174.800 137.000 175.200 ;
        RECT 137.400 174.800 137.800 175.200 ;
        RECT 138.200 174.800 138.600 175.200 ;
        RECT 139.000 174.800 139.400 175.200 ;
        RECT 142.200 174.800 142.600 175.200 ;
        RECT 135.800 166.800 136.200 167.200 ;
        RECT 133.400 165.800 133.800 166.200 ;
        RECT 134.200 165.800 134.600 166.200 ;
        RECT 135.800 165.800 136.200 166.200 ;
        RECT 132.600 161.800 133.000 162.200 ;
        RECT 129.400 158.800 129.800 159.200 ;
        RECT 128.600 156.100 129.000 156.200 ;
        RECT 127.800 155.800 129.000 156.100 ;
        RECT 127.800 155.100 128.200 155.200 ;
        RECT 128.600 155.100 129.000 155.200 ;
        RECT 127.800 154.800 129.000 155.100 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 130.200 154.200 130.500 154.800 ;
        RECT 130.200 153.800 130.600 154.200 ;
        RECT 130.200 153.200 130.500 153.800 ;
        RECT 130.200 152.800 130.600 153.200 ;
        RECT 131.000 153.100 131.400 155.900 ;
        RECT 131.800 155.800 132.200 156.200 ;
        RECT 131.800 154.200 132.100 155.800 ;
        RECT 131.800 153.800 132.200 154.200 ;
        RECT 132.600 152.100 133.000 157.900 ;
        RECT 134.200 154.200 134.500 165.800 ;
        RECT 135.800 165.200 136.100 165.800 ;
        RECT 137.400 165.200 137.700 174.800 ;
        RECT 138.200 174.200 138.500 174.800 ;
        RECT 139.000 174.200 139.300 174.800 ;
        RECT 138.200 173.800 138.600 174.200 ;
        RECT 139.000 173.800 139.400 174.200 ;
        RECT 145.400 172.100 145.800 177.900 ;
        RECT 147.800 175.800 148.200 176.200 ;
        RECT 147.800 175.200 148.100 175.800 ;
        RECT 146.200 174.800 146.600 175.200 ;
        RECT 147.800 174.800 148.200 175.200 ;
        RECT 138.200 166.800 138.600 167.200 ;
        RECT 138.200 166.200 138.500 166.800 ;
        RECT 138.200 165.800 138.600 166.200 ;
        RECT 139.000 166.100 139.400 166.200 ;
        RECT 139.800 166.100 140.200 166.200 ;
        RECT 139.000 165.800 140.200 166.100 ;
        RECT 135.800 164.800 136.200 165.200 ;
        RECT 137.400 164.800 137.800 165.200 ;
        RECT 141.400 165.100 141.800 167.900 ;
        RECT 142.200 166.800 142.600 167.200 ;
        RECT 136.600 162.100 137.000 162.200 ;
        RECT 137.400 162.100 137.800 162.200 ;
        RECT 136.600 161.800 137.800 162.100 ;
        RECT 142.200 158.200 142.500 166.800 ;
        RECT 143.000 163.100 143.400 168.900 ;
        RECT 146.200 168.200 146.500 174.800 ;
        RECT 150.200 172.100 150.600 177.900 ;
        RECT 151.000 172.100 151.300 185.800 ;
        RECT 151.800 183.100 152.200 188.900 ;
        RECT 152.600 188.800 153.000 189.200 ;
        RECT 152.600 188.200 152.900 188.800 ;
        RECT 152.600 187.800 153.000 188.200 ;
        RECT 152.600 186.800 153.000 187.200 ;
        RECT 152.600 186.300 152.900 186.800 ;
        RECT 152.600 185.900 153.000 186.300 ;
        RECT 152.600 185.800 152.900 185.900 ;
        RECT 155.000 181.200 155.300 204.800 ;
        RECT 156.600 201.200 156.900 206.800 ;
        RECT 157.400 205.800 157.800 206.200 ;
        RECT 156.600 200.800 157.000 201.200 ;
        RECT 157.400 200.200 157.700 205.800 ;
        RECT 163.000 203.100 163.400 208.900 ;
        RECT 167.000 205.900 167.400 206.300 ;
        RECT 167.000 204.200 167.300 205.900 ;
        RECT 167.000 203.800 167.400 204.200 ;
        RECT 167.800 203.100 168.200 208.900 ;
        RECT 168.600 206.800 169.000 207.200 ;
        RECT 168.600 206.200 168.900 206.800 ;
        RECT 168.600 205.800 169.000 206.200 ;
        RECT 169.400 205.100 169.800 207.900 ;
        RECT 175.000 207.800 175.400 208.200 ;
        RECT 175.000 207.200 175.300 207.800 ;
        RECT 170.200 206.800 170.600 207.200 ;
        RECT 173.400 206.800 173.800 207.200 ;
        RECT 175.000 206.800 175.400 207.200 ;
        RECT 159.000 201.800 159.400 202.200 ;
        RECT 160.600 201.800 161.000 202.200 ;
        RECT 157.400 199.800 157.800 200.200 ;
        RECT 157.400 194.700 157.800 195.100 ;
        RECT 155.800 192.800 156.200 193.200 ;
        RECT 155.000 180.800 155.400 181.200 ;
        RECT 155.000 179.800 155.400 180.200 ;
        RECT 151.800 173.100 152.200 175.900 ;
        RECT 153.400 175.100 153.800 175.200 ;
        RECT 154.200 175.100 154.600 175.200 ;
        RECT 153.400 174.800 154.600 175.100 ;
        RECT 152.600 174.100 153.000 174.200 ;
        RECT 153.400 174.100 153.800 174.200 ;
        RECT 152.600 173.800 153.800 174.100 ;
        RECT 154.200 173.800 154.600 174.200 ;
        RECT 151.000 171.800 152.100 172.100 ;
        RECT 150.200 169.800 150.600 170.200 ;
        RECT 150.200 169.200 150.500 169.800 ;
        RECT 146.200 167.800 146.600 168.200 ;
        RECT 146.200 167.200 146.500 167.800 ;
        RECT 144.600 166.800 145.000 167.200 ;
        RECT 146.200 166.800 146.600 167.200 ;
        RECT 144.600 166.200 144.900 166.800 ;
        RECT 144.600 165.800 145.000 166.200 ;
        RECT 147.800 163.100 148.200 168.900 ;
        RECT 150.200 168.800 150.600 169.200 ;
        RECT 151.800 168.200 152.100 171.800 ;
        RECT 151.800 167.800 152.200 168.200 ;
        RECT 154.200 167.200 154.500 173.800 ;
        RECT 155.000 167.200 155.300 179.800 ;
        RECT 155.800 176.200 156.100 192.800 ;
        RECT 157.400 189.200 157.700 194.700 ;
        RECT 158.200 192.100 158.600 197.900 ;
        RECT 159.000 197.200 159.300 201.800 ;
        RECT 160.600 198.200 160.900 201.800 ;
        RECT 170.200 199.200 170.500 206.800 ;
        RECT 173.400 206.200 173.700 206.800 ;
        RECT 171.000 205.800 171.400 206.200 ;
        RECT 173.400 205.800 173.800 206.200 ;
        RECT 171.000 205.200 171.300 205.800 ;
        RECT 171.000 204.800 171.400 205.200 ;
        RECT 172.600 205.100 173.000 205.200 ;
        RECT 173.400 205.100 173.800 205.200 ;
        RECT 175.800 205.100 176.200 207.900 ;
        RECT 172.600 204.800 173.800 205.100 ;
        RECT 176.600 203.800 177.000 204.200 ;
        RECT 176.600 199.200 176.900 203.800 ;
        RECT 177.400 203.100 177.800 208.900 ;
        RECT 181.400 206.800 181.800 207.200 ;
        RECT 178.200 205.900 178.600 206.300 ;
        RECT 181.400 206.200 181.700 206.800 ;
        RECT 178.200 205.200 178.500 205.900 ;
        RECT 181.400 205.800 181.800 206.200 ;
        RECT 178.200 204.800 178.600 205.200 ;
        RECT 182.200 203.100 182.600 208.900 ;
        RECT 184.600 208.800 185.000 209.200 ;
        RECT 211.000 208.800 211.400 209.200 ;
        RECT 184.600 208.200 184.900 208.800 ;
        RECT 184.600 207.800 185.000 208.200 ;
        RECT 203.000 206.800 203.400 207.200 ;
        RECT 205.400 207.100 205.800 207.200 ;
        RECT 206.200 207.100 206.600 207.200 ;
        RECT 205.400 206.800 206.600 207.100 ;
        RECT 207.800 206.800 208.200 207.200 ;
        RECT 208.600 206.800 209.000 207.200 ;
        RECT 190.200 206.100 190.600 206.200 ;
        RECT 191.000 206.100 191.400 206.200 ;
        RECT 190.200 205.800 191.400 206.100 ;
        RECT 196.600 205.800 197.000 206.200 ;
        RECT 198.200 206.100 198.600 206.200 ;
        RECT 199.000 206.100 199.400 206.200 ;
        RECT 198.200 205.800 199.400 206.100 ;
        RECT 201.400 205.800 201.800 206.200 ;
        RECT 202.200 205.800 202.600 206.200 ;
        RECT 183.000 204.800 183.400 205.200 ;
        RECT 177.400 201.800 177.800 202.200 ;
        RECT 170.200 198.800 170.600 199.200 ;
        RECT 175.800 198.800 176.200 199.200 ;
        RECT 176.600 198.800 177.000 199.200 ;
        RECT 160.600 197.800 161.000 198.200 ;
        RECT 159.000 196.800 159.400 197.200 ;
        RECT 159.000 194.800 159.400 195.200 ;
        RECT 159.000 194.200 159.300 194.800 ;
        RECT 159.000 193.800 159.400 194.200 ;
        RECT 159.800 193.100 160.200 195.900 ;
        RECT 160.600 195.800 161.000 196.200 ;
        RECT 161.400 195.800 161.800 196.200 ;
        RECT 163.800 196.100 164.200 196.200 ;
        RECT 164.600 196.100 165.000 196.200 ;
        RECT 163.800 195.800 165.000 196.100 ;
        RECT 160.600 194.200 160.900 195.800 ;
        RECT 161.400 195.200 161.700 195.800 ;
        RECT 161.400 194.800 161.800 195.200 ;
        RECT 163.000 194.800 163.400 195.200 ;
        RECT 163.000 194.200 163.300 194.800 ;
        RECT 160.600 193.800 161.000 194.200 ;
        RECT 163.000 193.800 163.400 194.200 ;
        RECT 166.200 191.800 166.600 192.200 ;
        RECT 168.600 192.100 169.000 197.900 ;
        RECT 170.200 195.100 170.600 195.200 ;
        RECT 171.000 195.100 171.400 195.200 ;
        RECT 170.200 194.800 171.400 195.100 ;
        RECT 171.000 193.800 171.400 194.200 ;
        RECT 156.600 183.100 157.000 188.900 ;
        RECT 157.400 188.800 157.800 189.200 ;
        RECT 161.400 189.100 161.800 189.200 ;
        RECT 162.200 189.100 162.600 189.200 ;
        RECT 161.400 188.800 162.600 189.100 ;
        RECT 166.200 188.200 166.500 191.800 ;
        RECT 166.200 187.800 166.600 188.200 ;
        RECT 159.800 186.800 160.200 187.200 ;
        RECT 163.800 187.100 164.200 187.200 ;
        RECT 164.600 187.100 165.000 187.200 ;
        RECT 163.800 186.800 165.000 187.100 ;
        RECT 167.800 187.100 168.200 187.200 ;
        RECT 168.600 187.100 169.000 187.200 ;
        RECT 167.800 186.800 169.000 187.100 ;
        RECT 159.800 186.200 160.100 186.800 ;
        RECT 159.800 185.800 160.200 186.200 ;
        RECT 161.400 185.800 161.800 186.200 ;
        RECT 163.000 186.100 163.400 186.200 ;
        RECT 163.800 186.100 164.200 186.200 ;
        RECT 163.000 185.800 164.200 186.100 ;
        RECT 161.400 185.200 161.700 185.800 ;
        RECT 161.400 184.800 161.800 185.200 ;
        RECT 158.200 184.100 158.600 184.200 ;
        RECT 159.000 184.100 159.400 184.200 ;
        RECT 158.200 183.800 159.400 184.100 ;
        RECT 159.000 180.800 159.400 181.200 ;
        RECT 155.800 175.800 156.200 176.200 ;
        RECT 155.800 175.200 156.100 175.800 ;
        RECT 159.000 175.200 159.300 180.800 ;
        RECT 161.400 179.200 161.700 184.800 ;
        RECT 169.400 183.100 169.800 188.900 ;
        RECT 171.000 186.200 171.300 193.800 ;
        RECT 173.400 192.100 173.800 197.900 ;
        RECT 175.000 193.100 175.400 195.900 ;
        RECT 175.800 194.200 176.100 198.800 ;
        RECT 176.600 194.800 177.000 195.200 ;
        RECT 175.800 193.800 176.200 194.200 ;
        RECT 176.600 193.200 176.900 194.800 ;
        RECT 176.600 192.800 177.000 193.200 ;
        RECT 173.400 187.800 173.800 188.200 ;
        RECT 173.400 186.300 173.700 187.800 ;
        RECT 171.000 185.800 171.400 186.200 ;
        RECT 173.400 185.900 173.800 186.300 ;
        RECT 173.400 185.800 173.700 185.900 ;
        RECT 165.400 181.800 165.800 182.200 ;
        RECT 167.000 181.800 167.400 182.200 ;
        RECT 165.400 180.200 165.700 181.800 ;
        RECT 165.400 179.800 165.800 180.200 ;
        RECT 161.400 178.800 161.800 179.200 ;
        RECT 163.000 176.800 163.400 177.200 ;
        RECT 161.400 175.800 161.800 176.200 ;
        RECT 161.400 175.200 161.700 175.800 ;
        RECT 155.800 174.800 156.200 175.200 ;
        RECT 158.200 174.800 158.600 175.200 ;
        RECT 159.000 174.800 159.400 175.200 ;
        RECT 161.400 174.800 161.800 175.200 ;
        RECT 158.200 174.200 158.500 174.800 ;
        RECT 157.400 173.800 157.800 174.200 ;
        RECT 158.200 173.800 158.600 174.200 ;
        RECT 157.400 170.200 157.700 173.800 ;
        RECT 159.000 172.200 159.300 174.800 ;
        RECT 163.000 174.200 163.300 176.800 ;
        RECT 160.600 174.100 161.000 174.200 ;
        RECT 161.400 174.100 161.800 174.200 ;
        RECT 160.600 173.800 161.800 174.100 ;
        RECT 163.000 173.800 163.400 174.200 ;
        RECT 163.800 173.100 164.200 175.900 ;
        RECT 159.000 171.800 159.400 172.200 ;
        RECT 165.400 172.100 165.800 177.900 ;
        RECT 166.200 174.700 166.600 175.100 ;
        RECT 166.200 174.200 166.500 174.700 ;
        RECT 166.200 173.800 166.600 174.200 ;
        RECT 166.200 172.800 166.600 173.200 ;
        RECT 157.400 169.800 157.800 170.200 ;
        RECT 154.200 166.800 154.600 167.200 ;
        RECT 155.000 166.800 155.400 167.200 ;
        RECT 155.800 167.100 156.200 167.200 ;
        RECT 156.600 167.100 157.000 167.200 ;
        RECT 155.800 166.800 157.000 167.100 ;
        RECT 152.600 165.800 153.000 166.200 ;
        RECT 153.400 165.800 153.800 166.200 ;
        RECT 154.200 165.800 154.600 166.200 ;
        RECT 155.000 166.100 155.400 166.200 ;
        RECT 155.800 166.100 156.200 166.200 ;
        RECT 155.000 165.800 156.200 166.100 ;
        RECT 157.400 165.800 157.800 166.200 ;
        RECT 152.600 165.200 152.900 165.800 ;
        RECT 152.600 164.800 153.000 165.200 ;
        RECT 143.800 161.800 144.200 162.200 ;
        RECT 151.000 161.800 151.400 162.200 ;
        RECT 135.800 155.800 136.200 156.200 ;
        RECT 135.800 155.200 136.100 155.800 ;
        RECT 135.800 154.800 136.200 155.200 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 134.200 153.800 134.600 154.200 ;
        RECT 133.400 149.200 133.700 153.800 ;
        RECT 137.400 152.100 137.800 157.900 ;
        RECT 138.200 157.800 138.600 158.200 ;
        RECT 142.200 157.800 142.600 158.200 ;
        RECT 138.200 157.200 138.500 157.800 ;
        RECT 138.200 156.800 138.600 157.200 ;
        RECT 143.800 156.200 144.100 161.800 ;
        RECT 151.000 157.200 151.300 161.800 ;
        RECT 145.400 156.800 145.800 157.200 ;
        RECT 151.000 156.800 151.400 157.200 ;
        RECT 145.400 156.200 145.700 156.800 ;
        RECT 142.200 155.800 142.600 156.200 ;
        RECT 143.800 155.800 144.200 156.200 ;
        RECT 145.400 155.800 145.800 156.200 ;
        RECT 148.600 155.800 149.000 156.200 ;
        RECT 139.000 152.800 139.400 153.200 ;
        RECT 139.800 153.100 140.200 153.200 ;
        RECT 140.600 153.100 141.000 153.200 ;
        RECT 139.800 152.800 141.000 153.100 ;
        RECT 139.000 152.200 139.300 152.800 ;
        RECT 139.000 151.800 139.400 152.200 ;
        RECT 139.800 151.800 140.200 152.200 ;
        RECT 133.400 148.800 133.800 149.200 ;
        RECT 128.600 147.800 129.000 148.200 ;
        RECT 131.800 147.800 132.200 148.200 ;
        RECT 133.400 147.800 133.800 148.200 ;
        RECT 136.600 147.800 137.000 148.200 ;
        RECT 128.600 147.200 128.900 147.800 ;
        RECT 131.800 147.200 132.100 147.800 ;
        RECT 127.800 147.100 128.200 147.200 ;
        RECT 127.000 146.800 128.200 147.100 ;
        RECT 128.600 146.800 129.000 147.200 ;
        RECT 131.800 146.800 132.200 147.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 114.200 146.100 114.600 146.200 ;
        RECT 112.600 145.800 114.600 146.100 ;
        RECT 113.400 144.800 113.800 145.200 ;
        RECT 111.000 143.100 111.400 143.200 ;
        RECT 111.800 143.100 112.200 143.200 ;
        RECT 111.000 142.800 112.200 143.100 ;
        RECT 112.600 142.800 113.000 143.200 ;
        RECT 112.600 137.200 112.900 142.800 ;
        RECT 113.400 142.200 113.700 144.800 ;
        RECT 116.600 144.200 116.900 146.800 ;
        RECT 119.000 145.800 119.400 146.200 ;
        RECT 121.400 145.800 121.800 146.200 ;
        RECT 119.000 145.200 119.300 145.800 ;
        RECT 121.400 145.200 121.700 145.800 ;
        RECT 123.000 145.200 123.300 146.800 ;
        RECT 123.800 145.800 124.200 146.200 ;
        RECT 123.800 145.200 124.100 145.800 ;
        RECT 119.000 144.800 119.400 145.200 ;
        RECT 121.400 144.800 121.800 145.200 ;
        RECT 123.000 144.800 123.400 145.200 ;
        RECT 123.800 144.800 124.200 145.200 ;
        RECT 116.600 143.800 117.000 144.200 ;
        RECT 120.600 142.800 121.000 143.200 ;
        RECT 113.400 141.800 113.800 142.200 ;
        RECT 117.400 141.800 117.800 142.200 ;
        RECT 113.400 138.200 113.700 141.800 ;
        RECT 117.400 139.200 117.700 141.800 ;
        RECT 120.600 141.200 120.900 142.800 ;
        RECT 120.600 140.800 121.000 141.200 ;
        RECT 120.600 139.200 120.900 140.800 ;
        RECT 117.400 138.800 117.800 139.200 ;
        RECT 120.600 138.800 121.000 139.200 ;
        RECT 123.000 138.800 123.400 139.200 ;
        RECT 123.000 138.200 123.300 138.800 ;
        RECT 113.400 137.800 113.800 138.200 ;
        RECT 119.800 137.800 120.200 138.200 ;
        RECT 123.000 137.800 123.400 138.200 ;
        RECT 119.800 137.200 120.100 137.800 ;
        RECT 125.400 137.200 125.700 146.800 ;
        RECT 126.200 145.800 126.600 146.200 ;
        RECT 126.200 145.200 126.500 145.800 ;
        RECT 126.200 144.800 126.600 145.200 ;
        RECT 127.000 138.200 127.300 146.800 ;
        RECT 127.800 145.800 128.200 146.200 ;
        RECT 129.400 146.100 129.800 146.200 ;
        RECT 130.200 146.100 130.600 146.200 ;
        RECT 129.400 145.800 130.600 146.100 ;
        RECT 131.800 145.800 132.200 146.200 ;
        RECT 127.800 145.200 128.100 145.800 ;
        RECT 131.800 145.200 132.100 145.800 ;
        RECT 133.400 145.200 133.700 147.800 ;
        RECT 136.600 147.200 136.900 147.800 ;
        RECT 139.000 147.200 139.300 151.800 ;
        RECT 139.800 151.200 140.100 151.800 ;
        RECT 139.800 150.800 140.200 151.200 ;
        RECT 142.200 147.200 142.500 155.800 ;
        RECT 148.600 155.200 148.900 155.800 ;
        RECT 145.400 154.800 145.800 155.200 ;
        RECT 147.000 155.100 147.400 155.200 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 147.000 154.800 148.200 155.100 ;
        RECT 148.600 154.800 149.000 155.200 ;
        RECT 149.400 154.800 149.800 155.200 ;
        RECT 145.400 154.200 145.700 154.800 ;
        RECT 145.400 153.800 145.800 154.200 ;
        RECT 146.200 153.800 146.600 154.200 ;
        RECT 146.200 153.200 146.500 153.800 ;
        RECT 143.000 152.800 143.400 153.200 ;
        RECT 146.200 152.800 146.600 153.200 ;
        RECT 148.600 152.800 149.000 153.200 ;
        RECT 143.000 152.200 143.300 152.800 ;
        RECT 143.000 151.800 143.400 152.200 ;
        RECT 144.600 151.800 145.000 152.200 ;
        RECT 135.000 147.100 135.400 147.200 ;
        RECT 135.800 147.100 136.200 147.200 ;
        RECT 135.000 146.800 136.200 147.100 ;
        RECT 136.600 146.800 137.000 147.200 ;
        RECT 139.000 146.800 139.400 147.200 ;
        RECT 139.800 147.100 140.200 147.200 ;
        RECT 140.600 147.100 141.000 147.200 ;
        RECT 139.800 146.800 141.000 147.100 ;
        RECT 142.200 146.800 142.600 147.200 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 141.400 145.800 141.800 146.200 ;
        RECT 135.800 145.200 136.100 145.800 ;
        RECT 127.800 144.800 128.200 145.200 ;
        RECT 130.200 145.100 130.600 145.200 ;
        RECT 131.000 145.100 131.400 145.200 ;
        RECT 130.200 144.800 131.400 145.100 ;
        RECT 131.800 144.800 132.200 145.200 ;
        RECT 133.400 144.800 133.800 145.200 ;
        RECT 135.800 145.100 136.200 145.200 ;
        RECT 136.600 145.100 137.000 145.200 ;
        RECT 135.800 144.800 137.000 145.100 ;
        RECT 137.400 143.800 137.800 144.200 ;
        RECT 132.600 141.800 133.000 142.200 ;
        RECT 127.000 137.800 127.400 138.200 ;
        RECT 129.400 137.800 129.800 138.200 ;
        RECT 112.600 136.800 113.000 137.200 ;
        RECT 116.600 136.800 117.000 137.200 ;
        RECT 119.800 136.800 120.200 137.200 ;
        RECT 121.400 137.100 121.800 137.200 ;
        RECT 122.200 137.100 122.600 137.200 ;
        RECT 121.400 136.800 122.600 137.100 ;
        RECT 125.400 136.800 125.800 137.200 ;
        RECT 116.600 136.200 116.900 136.800 ;
        RECT 115.000 135.800 115.400 136.200 ;
        RECT 116.600 135.800 117.000 136.200 ;
        RECT 119.000 136.100 119.400 136.200 ;
        RECT 119.800 136.100 120.200 136.200 ;
        RECT 119.000 135.800 120.200 136.100 ;
        RECT 123.800 136.100 124.200 136.200 ;
        RECT 124.600 136.100 125.000 136.200 ;
        RECT 123.800 135.800 125.000 136.100 ;
        RECT 115.000 135.200 115.300 135.800 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 113.400 134.800 113.800 135.200 ;
        RECT 115.000 134.800 115.400 135.200 ;
        RECT 115.800 134.800 116.200 135.200 ;
        RECT 119.000 134.800 119.400 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 123.800 135.100 124.200 135.200 ;
        RECT 123.000 134.800 124.200 135.100 ;
        RECT 111.000 134.200 111.300 134.800 ;
        RECT 113.400 134.200 113.700 134.800 ;
        RECT 115.800 134.200 116.100 134.800 ;
        RECT 119.000 134.200 119.300 134.800 ;
        RECT 125.400 134.200 125.700 136.800 ;
        RECT 127.000 136.100 127.400 136.200 ;
        RECT 127.800 136.100 128.200 136.200 ;
        RECT 127.000 135.800 128.200 136.100 ;
        RECT 129.400 135.200 129.700 137.800 ;
        RECT 132.600 137.200 132.900 141.800 ;
        RECT 131.000 136.800 131.400 137.200 ;
        RECT 132.600 136.800 133.000 137.200 ;
        RECT 135.800 136.800 136.200 137.200 ;
        RECT 131.000 136.200 131.300 136.800 ;
        RECT 131.000 135.800 131.400 136.200 ;
        RECT 135.000 135.800 135.400 136.200 ;
        RECT 135.000 135.200 135.300 135.800 ;
        RECT 126.200 135.100 126.600 135.200 ;
        RECT 127.000 135.100 127.400 135.200 ;
        RECT 126.200 134.800 127.400 135.100 ;
        RECT 127.800 134.800 128.200 135.200 ;
        RECT 129.400 134.800 129.800 135.200 ;
        RECT 132.600 134.800 133.000 135.200 ;
        RECT 135.000 134.800 135.400 135.200 ;
        RECT 127.800 134.200 128.100 134.800 ;
        RECT 111.000 133.800 111.400 134.200 ;
        RECT 113.400 133.800 113.800 134.200 ;
        RECT 115.800 133.800 116.200 134.200 ;
        RECT 119.000 133.800 119.400 134.200 ;
        RECT 123.800 133.800 124.200 134.200 ;
        RECT 125.400 133.800 125.800 134.200 ;
        RECT 127.800 133.800 128.200 134.200 ;
        RECT 111.800 132.100 112.200 132.200 ;
        RECT 112.600 132.100 113.000 132.200 ;
        RECT 111.800 131.800 113.000 132.100 ;
        RECT 113.400 130.200 113.700 133.800 ;
        RECT 115.800 131.800 116.200 132.200 ;
        RECT 115.800 131.200 116.100 131.800 ;
        RECT 115.800 130.800 116.200 131.200 ;
        RECT 116.600 130.800 117.000 131.200 ;
        RECT 111.800 129.800 112.200 130.200 ;
        RECT 113.400 129.800 113.800 130.200 ;
        RECT 115.000 129.800 115.400 130.200 ;
        RECT 111.800 126.200 112.100 129.800 ;
        RECT 115.000 129.200 115.300 129.800 ;
        RECT 115.000 128.800 115.400 129.200 ;
        RECT 116.600 128.200 116.900 130.800 ;
        RECT 116.600 127.800 117.000 128.200 ;
        RECT 121.400 127.800 121.800 128.200 ;
        RECT 116.600 127.200 116.900 127.800 ;
        RECT 115.000 126.800 115.400 127.200 ;
        RECT 116.600 126.800 117.000 127.200 ;
        RECT 117.400 127.100 117.800 127.200 ;
        RECT 118.200 127.100 118.600 127.200 ;
        RECT 117.400 126.800 118.600 127.100 ;
        RECT 119.800 126.800 120.200 127.200 ;
        RECT 115.000 126.200 115.300 126.800 ;
        RECT 119.800 126.200 120.100 126.800 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 115.000 125.800 115.400 126.200 ;
        RECT 118.200 125.800 118.600 126.200 ;
        RECT 119.800 125.800 120.200 126.200 ;
        RECT 120.600 125.800 121.000 126.200 ;
        RECT 111.800 125.200 112.100 125.800 ;
        RECT 118.200 125.200 118.500 125.800 ;
        RECT 111.000 124.800 111.400 125.200 ;
        RECT 111.800 124.800 112.200 125.200 ;
        RECT 112.600 124.800 113.000 125.200 ;
        RECT 114.200 124.800 114.600 125.200 ;
        RECT 115.000 124.800 115.400 125.200 ;
        RECT 115.800 124.800 116.200 125.200 ;
        RECT 117.400 124.800 117.800 125.200 ;
        RECT 118.200 124.800 118.600 125.200 ;
        RECT 119.000 124.800 119.400 125.200 ;
        RECT 111.000 124.200 111.300 124.800 ;
        RECT 110.200 123.800 110.600 124.200 ;
        RECT 111.000 123.800 111.400 124.200 ;
        RECT 112.600 122.200 112.900 124.800 ;
        RECT 108.600 121.800 109.000 122.200 ;
        RECT 110.200 121.800 110.600 122.200 ;
        RECT 111.800 121.800 112.200 122.200 ;
        RECT 112.600 121.800 113.000 122.200 ;
        RECT 113.400 121.800 113.800 122.200 ;
        RECT 107.800 120.800 108.200 121.200 ;
        RECT 110.200 119.200 110.500 121.800 ;
        RECT 110.200 118.800 110.600 119.200 ;
        RECT 111.800 118.200 112.100 121.800 ;
        RECT 113.400 120.200 113.700 121.800 ;
        RECT 113.400 119.800 113.800 120.200 ;
        RECT 114.200 119.200 114.500 124.800 ;
        RECT 115.000 124.200 115.300 124.800 ;
        RECT 115.000 123.800 115.400 124.200 ;
        RECT 115.800 122.200 116.100 124.800 ;
        RECT 115.800 121.800 116.200 122.200 ;
        RECT 114.200 118.800 114.600 119.200 ;
        RECT 111.800 117.800 112.200 118.200 ;
        RECT 113.400 117.800 113.800 118.200 ;
        RECT 111.800 116.800 112.200 117.200 ;
        RECT 111.800 116.200 112.100 116.800 ;
        RECT 107.800 116.100 108.200 116.200 ;
        RECT 108.600 116.100 109.000 116.200 ;
        RECT 107.800 115.800 109.000 116.100 ;
        RECT 111.800 115.800 112.200 116.200 ;
        RECT 113.400 114.200 113.700 117.800 ;
        RECT 115.800 117.200 116.100 121.800 ;
        RECT 117.400 117.200 117.700 124.800 ;
        RECT 119.000 117.200 119.300 124.800 ;
        RECT 120.600 124.200 120.900 125.800 ;
        RECT 121.400 125.200 121.700 127.800 ;
        RECT 123.800 126.200 124.100 133.800 ;
        RECT 124.600 132.800 125.000 133.200 ;
        RECT 127.800 133.100 128.200 133.200 ;
        RECT 128.600 133.100 129.000 133.200 ;
        RECT 127.800 132.800 129.000 133.100 ;
        RECT 124.600 132.200 124.900 132.800 ;
        RECT 124.600 131.800 125.000 132.200 ;
        RECT 126.200 131.800 126.600 132.200 ;
        RECT 124.600 126.200 124.900 131.800 ;
        RECT 123.800 125.800 124.200 126.200 ;
        RECT 124.600 125.800 125.000 126.200 ;
        RECT 121.400 124.800 121.800 125.200 ;
        RECT 120.600 123.800 121.000 124.200 ;
        RECT 119.800 121.800 120.200 122.200 ;
        RECT 115.800 116.800 116.200 117.200 ;
        RECT 117.400 116.800 117.800 117.200 ;
        RECT 119.000 116.800 119.400 117.200 ;
        RECT 119.000 116.200 119.300 116.800 ;
        RECT 119.800 116.200 120.100 121.800 ;
        RECT 119.000 115.800 119.400 116.200 ;
        RECT 119.800 115.800 120.200 116.200 ;
        RECT 121.400 115.200 121.700 124.800 ;
        RECT 123.000 121.800 123.400 122.200 ;
        RECT 123.000 117.200 123.300 121.800 ;
        RECT 123.800 117.200 124.100 125.800 ;
        RECT 124.600 124.800 125.000 125.200 ;
        RECT 125.400 125.100 125.800 127.900 ;
        RECT 124.600 123.200 124.900 124.800 ;
        RECT 126.200 123.200 126.500 131.800 ;
        RECT 127.800 129.200 128.100 132.800 ;
        RECT 124.600 122.800 125.000 123.200 ;
        RECT 126.200 122.800 126.600 123.200 ;
        RECT 127.000 123.100 127.400 128.900 ;
        RECT 127.800 128.800 128.200 129.200 ;
        RECT 129.400 128.200 129.700 134.800 ;
        RECT 132.600 132.200 132.900 134.800 ;
        RECT 135.800 134.200 136.100 136.800 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 133.400 133.800 133.800 134.200 ;
        RECT 135.800 133.800 136.200 134.200 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 132.600 131.800 133.000 132.200 ;
        RECT 133.400 129.100 133.700 133.800 ;
        RECT 135.000 131.800 135.400 132.200 ;
        RECT 134.200 129.100 134.600 129.200 ;
        RECT 129.400 127.800 129.800 128.200 ;
        RECT 128.600 126.800 129.000 127.200 ;
        RECT 124.600 119.200 124.900 122.800 ;
        RECT 126.200 119.200 126.500 122.800 ;
        RECT 124.600 118.800 125.000 119.200 ;
        RECT 126.200 118.800 126.600 119.200 ;
        RECT 127.000 117.800 127.400 118.200 ;
        RECT 123.000 116.800 123.400 117.200 ;
        RECT 123.800 116.800 124.200 117.200 ;
        RECT 125.400 116.800 125.800 117.200 ;
        RECT 123.000 116.200 123.300 116.800 ;
        RECT 125.400 116.200 125.700 116.800 ;
        RECT 123.000 115.800 123.400 116.200 ;
        RECT 125.400 115.800 125.800 116.200 ;
        RECT 114.200 115.100 114.600 115.200 ;
        RECT 114.200 114.800 115.300 115.100 ;
        RECT 109.400 113.800 109.800 114.200 ;
        RECT 113.400 114.100 113.800 114.200 ;
        RECT 113.400 113.800 114.500 114.100 ;
        RECT 109.400 113.200 109.700 113.800 ;
        RECT 107.000 112.800 108.100 113.100 ;
        RECT 109.400 112.800 109.800 113.200 ;
        RECT 110.200 113.100 110.600 113.200 ;
        RECT 111.000 113.100 111.400 113.200 ;
        RECT 110.200 112.800 111.400 113.100 ;
        RECT 112.600 112.800 113.000 113.200 ;
        RECT 106.200 110.200 106.500 112.800 ;
        RECT 107.000 111.800 107.400 112.200 ;
        RECT 105.400 109.800 105.800 110.200 ;
        RECT 106.200 109.800 106.600 110.200 ;
        RECT 105.400 103.100 105.800 108.900 ;
        RECT 106.200 107.800 106.600 108.200 ;
        RECT 106.200 107.200 106.500 107.800 ;
        RECT 106.200 106.800 106.600 107.200 ;
        RECT 107.000 106.200 107.300 111.800 ;
        RECT 107.000 105.800 107.400 106.200 ;
        RECT 107.000 100.800 107.400 101.200 ;
        RECT 102.200 98.800 102.600 99.200 ;
        RECT 104.600 98.800 105.000 99.200 ;
        RECT 101.400 97.800 101.800 98.200 ;
        RECT 91.000 96.800 91.400 97.200 ;
        RECT 92.600 96.800 93.000 97.200 ;
        RECT 94.200 96.800 94.600 97.200 ;
        RECT 100.600 96.800 101.000 97.200 ;
        RECT 92.600 96.200 92.900 96.800 ;
        RECT 100.600 96.200 100.900 96.800 ;
        RECT 101.400 96.200 101.700 97.800 ;
        RECT 92.600 95.800 93.000 96.200 ;
        RECT 95.000 95.800 95.400 96.200 ;
        RECT 95.800 95.800 96.200 96.200 ;
        RECT 96.600 95.800 97.000 96.200 ;
        RECT 100.600 95.800 101.000 96.200 ;
        RECT 101.400 95.800 101.800 96.200 ;
        RECT 92.600 95.200 92.900 95.800 ;
        RECT 95.000 95.200 95.300 95.800 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 92.600 94.800 93.000 95.200 ;
        RECT 95.000 94.800 95.400 95.200 ;
        RECT 90.200 86.800 90.600 87.200 ;
        RECT 91.000 86.200 91.300 94.800 ;
        RECT 92.600 91.800 93.000 92.200 ;
        RECT 91.000 85.800 91.400 86.200 ;
        RECT 92.600 85.200 92.900 91.800 ;
        RECT 93.400 88.800 93.800 89.200 ;
        RECT 93.400 87.200 93.700 88.800 ;
        RECT 95.000 88.200 95.300 94.800 ;
        RECT 95.800 93.200 96.100 95.800 ;
        RECT 96.600 95.200 96.900 95.800 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 99.000 94.800 99.400 95.200 ;
        RECT 99.000 94.200 99.300 94.800 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 99.000 93.800 99.400 94.200 ;
        RECT 98.200 93.200 98.500 93.800 ;
        RECT 95.800 92.800 96.200 93.200 ;
        RECT 98.200 92.800 98.600 93.200 ;
        RECT 101.400 92.200 101.700 95.800 ;
        RECT 102.200 95.200 102.500 98.800 ;
        RECT 104.600 96.800 105.000 97.200 ;
        RECT 104.600 96.200 104.900 96.800 ;
        RECT 107.000 96.200 107.300 100.800 ;
        RECT 107.800 100.200 108.100 112.800 ;
        RECT 111.800 111.800 112.200 112.200 ;
        RECT 109.400 108.800 109.800 109.200 ;
        RECT 107.800 99.800 108.200 100.200 ;
        RECT 108.600 97.800 109.000 98.200 ;
        RECT 104.600 95.800 105.000 96.200 ;
        RECT 107.000 95.800 107.400 96.200 ;
        RECT 102.200 94.800 102.600 95.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 103.000 94.200 103.300 94.800 ;
        RECT 108.600 94.200 108.900 97.800 ;
        RECT 109.400 95.200 109.700 108.800 ;
        RECT 110.200 103.100 110.600 108.900 ;
        RECT 111.800 101.200 112.100 111.800 ;
        RECT 112.600 109.200 112.900 112.800 ;
        RECT 114.200 109.200 114.500 113.800 ;
        RECT 115.000 112.200 115.300 114.800 ;
        RECT 118.200 114.800 118.600 115.200 ;
        RECT 121.400 114.800 121.800 115.200 ;
        RECT 123.000 114.800 123.400 115.200 ;
        RECT 118.200 114.200 118.500 114.800 ;
        RECT 123.000 114.200 123.300 114.800 ;
        RECT 127.000 114.200 127.300 117.800 ;
        RECT 127.800 115.800 128.200 116.200 ;
        RECT 127.800 115.200 128.100 115.800 ;
        RECT 127.800 114.800 128.200 115.200 ;
        RECT 118.200 113.800 118.600 114.200 ;
        RECT 119.800 113.800 120.200 114.200 ;
        RECT 121.400 113.800 121.800 114.200 ;
        RECT 123.000 113.800 123.400 114.200 ;
        RECT 127.000 113.800 127.400 114.200 ;
        RECT 119.800 113.200 120.100 113.800 ;
        RECT 121.400 113.200 121.700 113.800 ;
        RECT 115.800 113.100 116.200 113.200 ;
        RECT 116.600 113.100 117.000 113.200 ;
        RECT 115.800 112.800 117.000 113.100 ;
        RECT 119.800 112.800 120.200 113.200 ;
        RECT 121.400 112.800 121.800 113.200 ;
        RECT 115.000 111.800 115.400 112.200 ;
        RECT 118.200 111.800 118.600 112.200 ;
        RECT 119.000 111.800 119.400 112.200 ;
        RECT 126.200 111.800 126.600 112.200 ;
        RECT 118.200 110.200 118.500 111.800 ;
        RECT 118.200 109.800 118.600 110.200 ;
        RECT 112.600 108.800 113.000 109.200 ;
        RECT 114.200 108.800 114.600 109.200 ;
        RECT 117.400 107.800 117.800 108.200 ;
        RECT 117.400 107.200 117.700 107.800 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 117.400 106.800 117.800 107.200 ;
        RECT 111.800 100.800 112.200 101.200 ;
        RECT 113.400 100.200 113.700 106.800 ;
        RECT 115.800 105.800 116.200 106.200 ;
        RECT 115.800 104.200 116.100 105.800 ;
        RECT 115.800 103.800 116.200 104.200 ;
        RECT 114.200 101.800 114.600 102.200 ;
        RECT 115.800 102.100 116.200 102.200 ;
        RECT 116.600 102.100 117.000 102.200 ;
        RECT 115.800 101.800 117.000 102.100 ;
        RECT 113.400 99.800 113.800 100.200 ;
        RECT 111.800 98.800 112.200 99.200 ;
        RECT 113.400 98.800 113.800 99.200 ;
        RECT 109.400 94.800 109.800 95.200 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 103.800 93.800 104.200 94.200 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 108.600 93.800 109.000 94.200 ;
        RECT 109.400 93.800 109.800 94.200 ;
        RECT 110.200 93.800 110.600 94.200 ;
        RECT 103.800 92.200 104.100 93.800 ;
        RECT 107.000 93.100 107.300 93.800 ;
        RECT 107.800 93.100 108.200 93.200 ;
        RECT 107.000 92.800 108.200 93.100 ;
        RECT 100.600 91.800 101.000 92.200 ;
        RECT 101.400 91.800 101.800 92.200 ;
        RECT 103.800 91.800 104.200 92.200 ;
        RECT 104.600 91.800 105.000 92.200 ;
        RECT 107.000 91.800 107.400 92.200 ;
        RECT 99.800 91.100 100.200 91.200 ;
        RECT 100.600 91.100 100.900 91.800 ;
        RECT 99.800 90.800 100.900 91.100 ;
        RECT 95.000 87.800 95.400 88.200 ;
        RECT 93.400 86.800 93.800 87.200 ;
        RECT 95.000 87.100 95.400 87.200 ;
        RECT 95.800 87.100 96.200 87.200 ;
        RECT 95.000 86.800 96.200 87.100 ;
        RECT 98.200 86.800 98.600 87.200 ;
        RECT 98.200 86.200 98.500 86.800 ;
        RECT 96.600 86.100 97.000 86.200 ;
        RECT 97.400 86.100 97.800 86.200 ;
        RECT 96.600 85.800 97.800 86.100 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 91.000 85.100 91.400 85.200 ;
        RECT 91.800 85.100 92.200 85.200 ;
        RECT 91.000 84.800 92.200 85.100 ;
        RECT 92.600 84.800 93.000 85.200 ;
        RECT 95.000 85.100 95.400 85.200 ;
        RECT 95.800 85.100 96.200 85.200 ;
        RECT 95.000 84.800 96.200 85.100 ;
        RECT 97.400 85.100 97.800 85.200 ;
        RECT 98.200 85.100 98.600 85.200 ;
        RECT 99.000 85.100 99.400 87.900 ;
        RECT 97.400 84.800 98.600 85.100 ;
        RECT 93.400 84.100 93.800 84.200 ;
        RECT 94.200 84.100 94.600 84.200 ;
        RECT 93.400 83.800 94.600 84.100 ;
        RECT 100.600 83.100 101.000 88.900 ;
        RECT 104.600 88.200 104.900 91.800 ;
        RECT 104.600 87.800 105.000 88.200 ;
        RECT 101.400 86.800 101.800 87.200 ;
        RECT 104.600 86.800 105.000 87.200 ;
        RECT 101.400 86.300 101.700 86.800 ;
        RECT 101.400 85.900 101.800 86.300 ;
        RECT 104.600 86.200 104.900 86.800 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 105.400 83.100 105.800 88.900 ;
        RECT 98.200 78.800 98.600 79.200 ;
        RECT 99.800 78.800 100.200 79.200 ;
        RECT 83.800 75.800 84.200 76.200 ;
        RECT 85.400 76.100 85.800 76.200 ;
        RECT 86.200 76.100 86.600 76.200 ;
        RECT 85.400 75.800 86.600 76.100 ;
        RECT 83.800 75.200 84.100 75.800 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 83.000 74.800 83.400 75.200 ;
        RECT 83.800 74.800 84.200 75.200 ;
        RECT 86.200 74.800 86.600 75.200 ;
        RECT 86.200 74.200 86.500 74.800 ;
        RECT 80.600 73.800 81.000 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 86.200 73.800 86.600 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 80.600 73.200 80.900 73.800 ;
        RECT 83.000 73.200 83.300 73.800 ;
        RECT 80.600 72.800 81.000 73.200 ;
        RECT 83.000 72.800 83.400 73.200 ;
        RECT 89.400 72.200 89.700 73.800 ;
        RECT 91.800 72.800 92.200 73.200 ;
        RECT 87.000 71.800 87.400 72.200 ;
        RECT 89.400 71.800 89.800 72.200 ;
        RECT 79.800 63.100 80.200 68.900 ;
        RECT 82.200 66.800 82.600 67.200 ;
        RECT 80.600 66.100 81.000 66.300 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 80.600 65.800 81.800 66.100 ;
        RECT 72.600 59.800 73.000 60.200 ;
        RECT 79.000 59.800 79.400 60.200 ;
        RECT 80.600 59.800 81.000 60.200 ;
        RECT 71.000 58.800 71.400 59.200 ;
        RECT 71.800 58.800 72.200 59.200 ;
        RECT 79.000 58.800 79.400 59.200 ;
        RECT 64.600 53.800 65.000 54.200 ;
        RECT 66.200 53.800 66.600 54.200 ;
        RECT 52.600 43.800 53.000 44.200 ;
        RECT 53.400 42.800 53.800 43.200 ;
        RECT 55.000 43.100 55.400 48.900 ;
        RECT 55.800 45.800 56.200 46.200 ;
        RECT 55.800 45.200 56.100 45.800 ;
        RECT 55.800 44.800 56.200 45.200 ;
        RECT 52.600 41.800 53.000 42.200 ;
        RECT 47.000 37.800 47.400 38.200 ;
        RECT 41.400 37.100 41.800 37.200 ;
        RECT 42.200 37.100 42.600 37.200 ;
        RECT 41.400 36.800 42.600 37.100 ;
        RECT 44.600 36.800 45.000 37.200 ;
        RECT 44.600 34.200 44.900 36.800 ;
        RECT 47.000 35.800 47.400 36.200 ;
        RECT 51.000 35.800 51.400 36.200 ;
        RECT 47.000 35.200 47.300 35.800 ;
        RECT 51.000 35.200 51.300 35.800 ;
        RECT 52.600 35.200 52.900 41.800 ;
        RECT 47.000 34.800 47.400 35.200 ;
        RECT 49.400 35.100 49.800 35.200 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 49.400 34.800 50.600 35.100 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 52.600 34.800 53.000 35.200 ;
        RECT 44.600 33.800 45.000 34.200 ;
        RECT 47.000 34.100 47.400 34.200 ;
        RECT 47.800 34.100 48.200 34.200 ;
        RECT 47.000 33.800 48.200 34.100 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 51.800 34.100 52.200 34.200 ;
        RECT 52.600 34.100 53.000 34.200 ;
        RECT 51.800 33.800 53.000 34.100 ;
        RECT 50.200 33.200 50.500 33.800 ;
        RECT 50.200 32.800 50.600 33.200 ;
        RECT 41.400 23.100 41.800 28.900 ;
        RECT 42.200 26.800 42.600 27.200 ;
        RECT 45.400 26.800 45.800 27.200 ;
        RECT 42.200 26.200 42.500 26.800 ;
        RECT 45.400 26.300 45.700 26.800 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 45.400 25.900 45.800 26.300 ;
        RECT 46.200 23.100 46.600 28.900 ;
        RECT 51.800 28.800 52.200 29.200 ;
        RECT 47.000 26.800 47.400 27.200 ;
        RECT 47.000 22.200 47.300 26.800 ;
        RECT 47.800 25.100 48.200 27.900 ;
        RECT 51.800 27.200 52.100 28.800 ;
        RECT 48.600 26.800 49.000 27.200 ;
        RECT 50.200 27.100 50.600 27.200 ;
        RECT 51.000 27.100 51.400 27.200 ;
        RECT 50.200 26.800 51.400 27.100 ;
        RECT 51.800 26.800 52.200 27.200 ;
        RECT 48.600 26.200 48.900 26.800 ;
        RECT 53.400 26.200 53.700 42.800 ;
        RECT 56.600 39.200 56.900 51.800 ;
        RECT 58.200 46.100 58.600 46.200 ;
        RECT 59.000 46.100 59.400 46.300 ;
        RECT 58.200 45.900 59.400 46.100 ;
        RECT 58.200 45.800 59.300 45.900 ;
        RECT 59.800 43.100 60.200 48.900 ;
        RECT 61.400 45.100 61.800 47.900 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 62.200 45.800 63.400 46.100 ;
        RECT 63.800 45.800 64.200 46.200 ;
        RECT 62.200 44.800 62.600 45.200 ;
        RECT 62.200 42.200 62.500 44.800 ;
        RECT 59.800 41.800 60.200 42.200 ;
        RECT 62.200 41.800 62.600 42.200 ;
        RECT 59.800 39.200 60.100 41.800 ;
        RECT 56.600 38.800 57.000 39.200 ;
        RECT 59.800 38.800 60.200 39.200 ;
        RECT 59.800 37.800 60.200 38.200 ;
        RECT 54.200 34.800 54.600 35.200 ;
        RECT 56.600 35.100 57.000 35.200 ;
        RECT 57.400 35.100 57.800 35.200 ;
        RECT 56.600 34.800 57.800 35.100 ;
        RECT 58.200 34.800 58.600 35.200 ;
        RECT 59.000 34.800 59.400 35.200 ;
        RECT 54.200 27.200 54.500 34.800 ;
        RECT 58.200 34.200 58.500 34.800 ;
        RECT 59.000 34.200 59.300 34.800 ;
        RECT 58.200 33.800 58.600 34.200 ;
        RECT 59.000 33.800 59.400 34.200 ;
        RECT 59.800 33.100 60.100 37.800 ;
        RECT 60.600 35.800 61.000 36.200 ;
        RECT 61.400 35.800 61.800 36.200 ;
        RECT 62.200 35.800 62.600 36.200 ;
        RECT 60.600 35.200 60.900 35.800 ;
        RECT 60.600 34.800 61.000 35.200 ;
        RECT 59.000 32.800 60.100 33.100 ;
        RECT 61.400 34.200 61.700 35.800 ;
        RECT 62.200 35.200 62.500 35.800 ;
        RECT 63.800 35.200 64.100 45.800 ;
        RECT 64.600 45.200 64.900 46.800 ;
        RECT 64.600 44.800 65.000 45.200 ;
        RECT 65.400 45.100 65.800 47.900 ;
        RECT 66.200 47.200 66.500 53.800 ;
        RECT 68.600 52.100 69.000 57.900 ;
        RECT 71.800 55.200 72.100 58.800 ;
        RECT 72.600 57.800 73.000 58.200 ;
        RECT 71.800 54.800 72.200 55.200 ;
        RECT 66.200 46.800 66.600 47.200 ;
        RECT 64.600 38.200 64.900 44.800 ;
        RECT 67.000 43.100 67.400 48.900 ;
        RECT 69.400 46.100 69.800 46.200 ;
        RECT 70.200 46.100 70.600 46.200 ;
        RECT 69.400 45.800 70.600 46.100 ;
        RECT 71.000 45.800 71.400 46.200 ;
        RECT 71.000 44.200 71.300 45.800 ;
        RECT 71.000 43.800 71.400 44.200 ;
        RECT 71.800 43.100 72.200 48.900 ;
        RECT 69.400 40.800 69.800 41.200 ;
        RECT 69.400 39.200 69.700 40.800 ;
        RECT 72.600 39.200 72.900 57.800 ;
        RECT 76.600 55.800 77.000 56.200 ;
        RECT 77.400 55.800 77.800 56.200 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 73.400 51.800 73.800 52.200 ;
        RECT 73.400 48.200 73.700 51.800 ;
        RECT 74.200 49.200 74.500 53.800 ;
        RECT 76.600 53.200 76.900 55.800 ;
        RECT 77.400 55.200 77.700 55.800 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 78.200 54.800 78.600 55.200 ;
        RECT 78.200 54.200 78.500 54.800 ;
        RECT 78.200 53.800 78.600 54.200 ;
        RECT 76.600 52.800 77.000 53.200 ;
        RECT 75.800 51.800 76.200 52.200 ;
        RECT 74.200 48.800 74.600 49.200 ;
        RECT 73.400 47.800 73.800 48.200 ;
        RECT 75.000 46.800 75.400 47.200 ;
        RECT 75.000 46.200 75.300 46.800 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 75.000 45.100 75.400 45.200 ;
        RECT 75.800 45.100 76.100 51.800 ;
        RECT 76.600 46.200 76.900 52.800 ;
        RECT 77.400 46.800 77.800 47.200 ;
        RECT 76.600 45.800 77.000 46.200 ;
        RECT 75.000 44.800 76.100 45.100 ;
        RECT 77.400 45.200 77.700 46.800 ;
        RECT 79.000 46.200 79.300 58.800 ;
        RECT 80.600 55.200 80.900 59.800 ;
        RECT 80.600 54.800 81.000 55.200 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 81.400 54.200 81.700 54.800 ;
        RECT 81.400 53.800 81.800 54.200 ;
        RECT 80.600 47.100 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 80.600 46.800 81.800 47.100 ;
        RECT 79.000 45.800 79.400 46.200 ;
        RECT 79.000 45.200 79.300 45.800 ;
        RECT 77.400 44.800 77.800 45.200 ;
        RECT 79.000 44.800 79.400 45.200 ;
        RECT 80.600 45.100 81.000 45.200 ;
        RECT 81.400 45.100 81.800 45.200 ;
        RECT 80.600 44.800 81.800 45.100 ;
        RECT 82.200 44.200 82.500 66.800 ;
        RECT 84.600 63.100 85.000 68.900 ;
        RECT 84.600 59.800 85.000 60.200 ;
        RECT 84.600 59.200 84.900 59.800 ;
        RECT 84.600 58.800 85.000 59.200 ;
        RECT 83.000 54.800 83.400 55.200 ;
        RECT 85.400 54.800 85.800 55.200 ;
        RECT 82.200 43.800 82.600 44.200 ;
        RECT 80.600 41.800 81.000 42.200 ;
        RECT 76.600 39.800 77.000 40.200 ;
        RECT 69.400 38.800 69.800 39.200 ;
        RECT 72.600 38.800 73.000 39.200 ;
        RECT 64.600 37.800 65.000 38.200 ;
        RECT 76.600 37.200 76.900 39.800 ;
        RECT 72.600 36.800 73.000 37.200 ;
        RECT 76.600 36.800 77.000 37.200 ;
        RECT 64.600 36.100 65.000 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 64.600 35.800 65.800 36.100 ;
        RECT 72.600 35.200 72.900 36.800 ;
        RECT 80.600 36.200 80.900 41.800 ;
        RECT 83.000 39.200 83.300 54.800 ;
        RECT 85.400 54.200 85.700 54.800 ;
        RECT 85.400 53.800 85.800 54.200 ;
        RECT 84.600 52.800 85.000 53.200 ;
        RECT 83.800 41.800 84.200 42.200 ;
        RECT 83.800 40.200 84.100 41.800 ;
        RECT 83.800 39.800 84.200 40.200 ;
        RECT 83.000 38.800 83.400 39.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 80.600 35.200 80.900 35.800 ;
        RECT 62.200 34.800 62.600 35.200 ;
        RECT 63.800 34.800 64.200 35.200 ;
        RECT 67.800 34.800 68.200 35.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 72.600 34.800 73.000 35.200 ;
        RECT 78.200 35.100 78.600 35.200 ;
        RECT 79.000 35.100 79.400 35.200 ;
        RECT 78.200 34.800 79.400 35.100 ;
        RECT 80.600 34.800 81.000 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 83.000 34.800 83.400 35.200 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 61.400 33.200 61.700 33.800 ;
        RECT 61.400 32.800 61.800 33.200 ;
        RECT 63.000 32.800 63.400 33.200 ;
        RECT 59.000 27.200 59.300 32.800 ;
        RECT 61.400 30.200 61.700 32.800 ;
        RECT 61.400 29.800 61.800 30.200 ;
        RECT 54.200 26.800 54.600 27.200 ;
        RECT 59.000 26.800 59.400 27.200 ;
        RECT 48.600 25.800 49.000 26.200 ;
        RECT 49.400 26.100 49.800 26.200 ;
        RECT 50.200 26.100 50.600 26.200 ;
        RECT 49.400 25.800 50.600 26.100 ;
        RECT 53.400 25.800 53.800 26.200 ;
        RECT 53.400 25.200 53.700 25.800 ;
        RECT 51.800 24.800 52.200 25.200 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 47.000 21.800 47.400 22.200 ;
        RECT 40.600 18.800 41.000 19.200 ;
        RECT 43.800 18.800 44.200 19.200 ;
        RECT 28.600 15.100 29.000 15.200 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 28.600 14.800 29.800 15.100 ;
        RECT 30.200 14.800 30.600 15.200 ;
        RECT 31.000 12.100 31.400 17.900 ;
        RECT 34.200 16.100 34.600 16.200 ;
        RECT 35.000 16.100 35.400 16.200 ;
        RECT 34.200 15.800 35.400 16.100 ;
        RECT 39.800 15.800 40.200 16.200 ;
        RECT 43.000 15.800 43.400 16.200 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 35.000 15.100 35.400 15.200 ;
        RECT 34.200 14.800 35.400 15.100 ;
        RECT 37.400 14.800 37.800 15.200 ;
        RECT 39.000 14.800 39.400 15.200 ;
        RECT 36.600 13.800 37.000 14.200 ;
        RECT 33.400 12.100 33.800 12.200 ;
        RECT 34.200 12.100 34.600 12.200 ;
        RECT 33.400 11.800 34.600 12.100 ;
        RECT 36.600 11.200 36.900 13.800 ;
        RECT 36.600 10.800 37.000 11.200 ;
        RECT 21.400 8.800 21.800 9.200 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 29.400 6.800 29.800 7.200 ;
        RECT 29.400 6.200 29.700 6.800 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 18.200 5.800 19.400 6.100 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 0.600 4.800 1.000 5.200 ;
        RECT 3.800 5.100 4.200 5.200 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 3.800 4.800 5.000 5.100 ;
        RECT 11.000 4.800 11.400 5.200 ;
        RECT 13.400 5.100 13.800 5.200 ;
        RECT 14.200 5.100 14.600 5.200 ;
        RECT 30.200 5.100 30.600 7.900 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 31.000 6.200 31.300 6.800 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 13.400 4.800 14.600 5.100 ;
        RECT 31.800 3.100 32.200 8.900 ;
        RECT 35.800 8.800 36.200 9.200 ;
        RECT 35.800 7.200 36.100 8.800 ;
        RECT 35.000 6.800 35.400 7.200 ;
        RECT 35.800 6.800 36.200 7.200 ;
        RECT 35.000 6.200 35.300 6.800 ;
        RECT 35.000 5.800 35.400 6.200 ;
        RECT 36.600 3.100 37.000 8.900 ;
        RECT 37.400 6.200 37.700 14.800 ;
        RECT 39.000 9.200 39.300 14.800 ;
        RECT 39.800 9.200 40.100 15.800 ;
        RECT 43.000 15.200 43.300 15.800 ;
        RECT 43.800 15.200 44.100 18.800 ;
        RECT 47.000 17.100 47.300 21.800 ;
        RECT 47.000 16.800 48.100 17.100 ;
        RECT 42.200 14.800 42.600 15.200 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 46.200 14.800 46.600 15.200 ;
        RECT 42.200 14.100 42.500 14.800 ;
        RECT 46.200 14.200 46.500 14.800 ;
        RECT 42.200 13.800 43.300 14.100 ;
        RECT 46.200 13.800 46.600 14.200 ;
        RECT 43.000 12.200 43.300 13.800 ;
        RECT 47.000 13.100 47.400 15.900 ;
        RECT 47.800 14.200 48.100 16.800 ;
        RECT 47.800 13.800 48.200 14.200 ;
        RECT 43.000 11.800 43.400 12.200 ;
        RECT 48.600 12.100 49.000 17.900 ;
        RECT 51.800 15.200 52.100 24.800 ;
        RECT 54.200 19.200 54.500 26.800 ;
        RECT 57.400 25.800 57.800 26.200 ;
        RECT 58.200 25.800 58.600 26.200 ;
        RECT 57.400 25.200 57.700 25.800 ;
        RECT 55.800 24.800 56.200 25.200 ;
        RECT 57.400 24.800 57.800 25.200 ;
        RECT 55.800 24.200 56.100 24.800 ;
        RECT 58.200 24.200 58.500 25.800 ;
        RECT 55.800 23.800 56.200 24.200 ;
        RECT 58.200 23.800 58.600 24.200 ;
        RECT 54.200 18.800 54.600 19.200 ;
        RECT 55.000 19.100 55.400 19.200 ;
        RECT 55.800 19.100 56.200 19.200 ;
        RECT 55.000 18.800 56.200 19.100 ;
        RECT 51.800 14.800 52.200 15.200 ;
        RECT 53.400 12.100 53.800 17.900 ;
        RECT 57.400 15.100 57.800 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 57.400 14.800 58.600 15.100 ;
        RECT 59.000 14.200 59.300 26.800 ;
        RECT 59.800 25.100 60.200 27.900 ;
        RECT 60.600 26.800 61.000 27.200 ;
        RECT 60.600 22.200 60.900 26.800 ;
        RECT 61.400 23.100 61.800 28.900 ;
        RECT 60.600 21.800 61.000 22.200 ;
        RECT 63.000 19.200 63.300 32.800 ;
        RECT 63.800 31.800 64.200 32.200 ;
        RECT 63.800 26.200 64.100 31.800 ;
        RECT 67.800 29.100 68.100 34.800 ;
        RECT 70.200 29.200 70.500 34.800 ;
        RECT 71.000 34.200 71.300 34.800 ;
        RECT 82.200 34.200 82.500 34.800 ;
        RECT 71.000 33.800 71.400 34.200 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 82.200 33.800 82.600 34.200 ;
        RECT 71.800 33.200 72.100 33.800 ;
        RECT 75.000 33.200 75.300 33.800 ;
        RECT 71.800 32.800 72.200 33.200 ;
        RECT 75.000 32.800 75.400 33.200 ;
        RECT 68.600 29.100 69.000 29.200 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 66.200 23.100 66.600 28.900 ;
        RECT 67.800 28.800 69.000 29.100 ;
        RECT 69.400 29.100 69.800 29.200 ;
        RECT 70.200 29.100 70.600 29.200 ;
        RECT 69.400 28.800 70.600 29.100 ;
        RECT 67.000 23.800 67.400 24.200 ;
        RECT 63.000 18.800 63.400 19.200 ;
        RECT 63.800 17.800 64.200 18.200 ;
        RECT 59.800 15.800 60.200 16.200 ;
        RECT 59.800 15.200 60.100 15.800 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 63.800 14.200 64.100 17.800 ;
        RECT 67.000 16.200 67.300 23.800 ;
        RECT 71.800 23.100 72.200 28.900 ;
        RECT 75.800 26.800 76.200 27.200 ;
        RECT 75.800 26.300 76.100 26.800 ;
        RECT 72.600 25.800 73.000 26.200 ;
        RECT 75.800 25.900 76.200 26.300 ;
        RECT 64.600 15.800 65.000 16.200 ;
        RECT 67.000 15.800 67.400 16.200 ;
        RECT 67.800 15.800 68.200 16.200 ;
        RECT 64.600 15.200 64.900 15.800 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 55.800 14.100 56.200 14.200 ;
        RECT 56.600 14.100 57.000 14.200 ;
        RECT 55.800 13.800 57.000 14.100 ;
        RECT 59.000 13.800 59.400 14.200 ;
        RECT 61.400 13.800 61.800 14.200 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 67.000 14.100 67.400 14.200 ;
        RECT 67.800 14.100 68.100 15.800 ;
        RECT 67.000 13.800 68.100 14.100 ;
        RECT 68.600 13.800 69.000 14.200 ;
        RECT 59.000 11.800 59.400 12.200 ;
        RECT 39.000 8.800 39.400 9.200 ;
        RECT 39.800 8.800 40.200 9.200 ;
        RECT 39.000 7.200 39.300 8.800 ;
        RECT 43.000 7.200 43.300 11.800 ;
        RECT 47.800 10.800 48.200 11.200 ;
        RECT 43.800 7.800 44.200 8.200 ;
        RECT 43.800 7.200 44.100 7.800 ;
        RECT 39.000 6.800 39.400 7.200 ;
        RECT 43.000 6.800 43.400 7.200 ;
        RECT 43.800 6.800 44.200 7.200 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 45.400 6.800 46.600 7.100 ;
        RECT 47.800 6.200 48.100 10.800 ;
        RECT 48.600 9.800 49.000 10.200 ;
        RECT 49.400 9.800 49.800 10.200 ;
        RECT 48.600 7.200 48.900 9.800 ;
        RECT 49.400 9.200 49.700 9.800 ;
        RECT 59.000 9.200 59.300 11.800 ;
        RECT 61.400 10.200 61.700 13.800 ;
        RECT 68.600 13.200 68.900 13.800 ;
        RECT 68.600 12.800 69.000 13.200 ;
        RECT 69.400 13.100 69.800 15.900 ;
        RECT 71.000 12.100 71.400 17.900 ;
        RECT 71.800 15.800 72.200 16.200 ;
        RECT 71.800 15.100 72.100 15.800 ;
        RECT 71.800 14.700 72.200 15.100 ;
        RECT 72.600 14.200 72.900 25.800 ;
        RECT 76.600 23.100 77.000 28.900 ;
        RECT 77.400 18.200 77.700 33.800 ;
        RECT 79.800 32.100 80.200 32.200 ;
        RECT 80.600 32.100 81.000 32.200 ;
        RECT 79.800 31.800 81.000 32.100 ;
        RECT 79.000 28.800 79.400 29.200 ;
        RECT 78.200 25.100 78.600 27.900 ;
        RECT 79.000 27.200 79.300 28.800 ;
        RECT 79.000 26.800 79.400 27.200 ;
        RECT 80.600 27.100 81.000 27.200 ;
        RECT 81.400 27.100 81.800 27.200 ;
        RECT 80.600 26.800 81.800 27.100 ;
        RECT 80.600 25.100 81.000 25.200 ;
        RECT 81.400 25.100 81.800 25.200 ;
        RECT 80.600 24.800 81.800 25.100 ;
        RECT 83.000 24.200 83.300 34.800 ;
        RECT 83.800 29.800 84.200 30.200 ;
        RECT 83.800 27.200 84.100 29.800 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 84.600 26.200 84.900 52.800 ;
        RECT 86.200 43.100 86.600 48.900 ;
        RECT 85.400 39.800 85.800 40.200 ;
        RECT 85.400 39.200 85.700 39.800 ;
        RECT 85.400 38.800 85.800 39.200 ;
        RECT 87.000 35.200 87.300 71.800 ;
        RECT 87.800 68.800 88.200 69.200 ;
        RECT 87.800 67.200 88.100 68.800 ;
        RECT 87.800 66.800 88.200 67.200 ;
        RECT 87.800 66.200 88.100 66.800 ;
        RECT 87.800 65.800 88.200 66.200 ;
        RECT 88.600 65.800 89.000 66.200 ;
        RECT 91.800 66.100 92.100 72.800 ;
        RECT 92.600 72.100 93.000 77.900 ;
        RECT 93.400 76.800 93.800 77.200 ;
        RECT 93.400 75.200 93.700 76.800 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 95.000 75.100 95.400 75.200 ;
        RECT 95.800 75.100 96.200 75.200 ;
        RECT 95.000 74.800 96.200 75.100 ;
        RECT 95.000 72.800 95.400 73.200 ;
        RECT 95.000 69.200 95.300 72.800 ;
        RECT 97.400 72.100 97.800 77.900 ;
        RECT 95.000 68.800 95.400 69.200 ;
        RECT 95.800 67.800 96.200 68.200 ;
        RECT 95.800 67.200 96.100 67.800 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 98.200 66.200 98.500 78.800 ;
        RECT 99.000 73.100 99.400 75.900 ;
        RECT 99.800 75.200 100.100 78.800 ;
        RECT 106.200 77.100 106.600 77.200 ;
        RECT 107.000 77.100 107.300 91.800 ;
        RECT 107.800 89.200 108.100 92.800 ;
        RECT 108.600 91.800 109.000 92.200 ;
        RECT 107.800 88.800 108.200 89.200 ;
        RECT 108.600 87.200 108.900 91.800 ;
        RECT 109.400 90.200 109.700 93.800 ;
        RECT 109.400 89.800 109.800 90.200 ;
        RECT 108.600 86.800 109.000 87.200 ;
        RECT 109.400 86.200 109.700 89.800 ;
        RECT 109.400 85.800 109.800 86.200 ;
        RECT 109.400 79.200 109.700 85.800 ;
        RECT 109.400 78.800 109.800 79.200 ;
        RECT 106.200 76.800 107.300 77.100 ;
        RECT 110.200 76.200 110.500 93.800 ;
        RECT 111.000 84.800 111.400 85.200 ;
        RECT 111.000 79.200 111.300 84.800 ;
        RECT 111.000 78.800 111.400 79.200 ;
        RECT 103.000 75.800 103.400 76.200 ;
        RECT 104.600 75.800 105.000 76.200 ;
        RECT 107.800 75.800 108.200 76.200 ;
        RECT 110.200 75.800 110.600 76.200 ;
        RECT 103.000 75.200 103.300 75.800 ;
        RECT 99.800 74.800 100.200 75.200 ;
        RECT 100.600 74.800 101.000 75.200 ;
        RECT 103.000 74.800 103.400 75.200 ;
        RECT 103.800 74.800 104.200 75.200 ;
        RECT 100.600 74.200 100.900 74.800 ;
        RECT 103.800 74.200 104.100 74.800 ;
        RECT 100.600 73.800 101.000 74.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 104.600 73.200 104.900 75.800 ;
        RECT 107.800 75.200 108.100 75.800 ;
        RECT 111.800 75.200 112.100 98.800 ;
        RECT 113.400 95.200 113.700 98.800 ;
        RECT 114.200 98.200 114.500 101.800 ;
        RECT 118.200 98.200 118.500 109.800 ;
        RECT 119.000 109.200 119.300 111.800 ;
        RECT 126.200 109.200 126.500 111.800 ;
        RECT 119.000 108.800 119.400 109.200 ;
        RECT 124.600 108.800 125.000 109.200 ;
        RECT 126.200 108.800 126.600 109.200 ;
        RECT 123.000 107.100 123.400 107.200 ;
        RECT 123.800 107.100 124.200 107.200 ;
        RECT 123.000 106.800 124.200 107.100 ;
        RECT 120.600 105.800 121.000 106.200 ;
        RECT 121.400 105.800 121.800 106.200 ;
        RECT 122.200 105.800 122.600 106.200 ;
        RECT 120.600 105.200 120.900 105.800 ;
        RECT 120.600 104.800 121.000 105.200 ;
        RECT 120.600 103.800 121.000 104.200 ;
        RECT 120.600 99.200 120.900 103.800 ;
        RECT 120.600 98.800 121.000 99.200 ;
        RECT 114.200 97.800 114.600 98.200 ;
        RECT 115.800 97.800 116.200 98.200 ;
        RECT 118.200 97.800 118.600 98.200 ;
        RECT 119.000 97.800 119.400 98.200 ;
        RECT 114.200 96.800 114.600 97.200 ;
        RECT 114.200 96.200 114.500 96.800 ;
        RECT 115.800 96.200 116.100 97.800 ;
        RECT 114.200 95.800 114.600 96.200 ;
        RECT 115.800 95.800 116.200 96.200 ;
        RECT 112.600 94.800 113.000 95.200 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 112.600 93.200 112.900 94.800 ;
        RECT 112.600 92.800 113.000 93.200 ;
        RECT 112.600 86.800 113.000 87.200 ;
        RECT 112.600 84.200 112.900 86.800 ;
        RECT 112.600 83.800 113.000 84.200 ;
        RECT 113.400 81.200 113.700 94.800 ;
        RECT 115.800 94.200 116.100 95.800 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 115.000 91.800 115.400 92.200 ;
        RECT 115.800 91.800 116.200 92.200 ;
        RECT 117.400 91.800 117.800 92.200 ;
        RECT 114.200 88.800 114.600 89.200 ;
        RECT 114.200 88.200 114.500 88.800 ;
        RECT 114.200 87.800 114.600 88.200 ;
        RECT 114.200 86.800 114.600 87.200 ;
        RECT 113.400 80.800 113.800 81.200 ;
        RECT 114.200 79.200 114.500 86.800 ;
        RECT 114.200 78.800 114.600 79.200 ;
        RECT 115.000 77.200 115.300 91.800 ;
        RECT 115.000 76.800 115.400 77.200 ;
        RECT 112.600 75.800 113.000 76.200 ;
        RECT 113.400 75.800 113.800 76.200 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 107.800 74.800 108.200 75.200 ;
        RECT 111.000 75.100 111.400 75.200 ;
        RECT 111.800 75.100 112.200 75.200 ;
        RECT 111.000 74.800 112.200 75.100 ;
        RECT 105.400 74.200 105.700 74.800 ;
        RECT 105.400 73.800 105.800 74.200 ;
        RECT 107.800 74.100 108.200 74.200 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 107.800 73.800 109.000 74.100 ;
        RECT 109.400 73.800 109.800 74.200 ;
        RECT 110.200 73.800 110.600 74.200 ;
        RECT 109.400 73.200 109.700 73.800 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 109.400 72.800 109.800 73.200 ;
        RECT 106.200 71.800 106.600 72.200 ;
        RECT 109.400 71.800 109.800 72.200 ;
        RECT 105.400 70.800 105.800 71.200 ;
        RECT 104.600 68.800 105.000 69.200 ;
        RECT 102.200 68.100 102.600 68.200 ;
        RECT 103.000 68.100 103.400 68.200 ;
        RECT 102.200 67.800 103.400 68.100 ;
        RECT 99.000 67.100 99.400 67.200 ;
        RECT 99.800 67.100 100.200 67.200 ;
        RECT 99.000 66.800 100.200 67.100 ;
        RECT 100.600 67.100 101.000 67.200 ;
        RECT 101.400 67.100 101.800 67.200 ;
        RECT 100.600 66.800 101.800 67.100 ;
        RECT 102.200 66.800 102.600 67.200 ;
        RECT 92.600 66.100 93.000 66.200 ;
        RECT 91.800 65.800 93.000 66.100 ;
        RECT 93.400 65.800 93.800 66.200 ;
        RECT 98.200 65.800 98.600 66.200 ;
        RECT 99.000 65.800 99.400 66.200 ;
        RECT 88.600 55.200 88.900 65.800 ;
        RECT 93.400 65.200 93.700 65.800 ;
        RECT 93.400 64.800 93.800 65.200 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 95.800 64.800 96.200 65.200 ;
        RECT 98.200 65.100 98.600 65.200 ;
        RECT 99.000 65.100 99.300 65.800 ;
        RECT 98.200 64.800 99.300 65.100 ;
        RECT 91.000 62.800 91.400 63.200 ;
        RECT 91.000 59.200 91.300 62.800 ;
        RECT 91.800 61.800 92.200 62.200 ;
        RECT 91.000 58.800 91.400 59.200 ;
        RECT 91.800 55.200 92.100 61.800 ;
        RECT 94.200 60.200 94.500 64.800 ;
        RECT 94.200 59.800 94.600 60.200 ;
        RECT 95.800 58.200 96.100 64.800 ;
        RECT 102.200 58.200 102.500 66.800 ;
        RECT 104.600 66.200 104.900 68.800 ;
        RECT 105.400 67.200 105.700 70.800 ;
        RECT 106.200 67.200 106.500 71.800 ;
        RECT 109.400 69.200 109.700 71.800 ;
        RECT 108.600 68.800 109.000 69.200 ;
        RECT 109.400 68.800 109.800 69.200 ;
        RECT 108.600 68.200 108.900 68.800 ;
        RECT 108.600 67.800 109.000 68.200 ;
        RECT 105.400 66.800 105.800 67.200 ;
        RECT 106.200 66.800 106.600 67.200 ;
        RECT 103.000 66.100 103.400 66.200 ;
        RECT 103.800 66.100 104.200 66.200 ;
        RECT 103.000 65.800 104.200 66.100 ;
        RECT 104.600 66.100 105.000 66.200 ;
        RECT 106.200 66.100 106.600 66.200 ;
        RECT 107.000 66.100 107.400 66.200 ;
        RECT 104.600 65.800 105.700 66.100 ;
        RECT 106.200 65.800 107.400 66.100 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 103.000 64.800 104.100 65.100 ;
        RECT 103.800 59.200 104.100 64.800 ;
        RECT 103.800 58.800 104.200 59.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 91.800 54.800 92.200 55.200 ;
        RECT 89.400 54.200 89.700 54.800 ;
        RECT 89.400 53.800 89.800 54.200 ;
        RECT 93.400 53.100 93.800 55.900 ;
        RECT 94.200 53.800 94.600 54.200 ;
        RECT 94.200 50.200 94.500 53.800 ;
        RECT 95.000 52.100 95.400 57.900 ;
        RECT 95.800 57.800 96.200 58.200 ;
        RECT 96.600 57.800 97.000 58.200 ;
        RECT 96.600 55.200 96.900 57.800 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 99.800 52.100 100.200 57.900 ;
        RECT 102.200 57.800 102.600 58.200 ;
        RECT 102.200 57.100 102.600 57.200 ;
        RECT 103.000 57.100 103.400 57.200 ;
        RECT 102.200 56.800 103.400 57.100 ;
        RECT 104.600 56.800 105.000 57.200 ;
        RECT 104.600 56.200 104.900 56.800 ;
        RECT 105.400 56.200 105.700 65.800 ;
        RECT 107.800 65.100 108.200 65.200 ;
        RECT 108.600 65.100 109.000 65.200 ;
        RECT 107.800 64.800 109.000 65.100 ;
        RECT 109.400 64.800 109.800 65.200 ;
        RECT 108.600 63.800 109.000 64.200 ;
        RECT 108.600 59.200 108.900 63.800 ;
        RECT 109.400 63.200 109.700 64.800 ;
        RECT 110.200 64.200 110.500 73.800 ;
        RECT 111.000 69.800 111.400 70.200 ;
        RECT 111.000 67.200 111.300 69.800 ;
        RECT 112.600 69.200 112.900 75.800 ;
        RECT 113.400 72.200 113.700 75.800 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 115.000 75.100 115.400 75.200 ;
        RECT 114.200 74.800 115.400 75.100 ;
        RECT 113.400 71.800 113.800 72.200 ;
        RECT 113.400 69.800 113.800 70.200 ;
        RECT 114.200 69.800 114.600 70.200 ;
        RECT 112.600 68.800 113.000 69.200 ;
        RECT 111.000 66.800 111.400 67.200 ;
        RECT 111.800 67.100 112.200 67.200 ;
        RECT 112.600 67.100 113.000 67.200 ;
        RECT 111.800 66.800 113.000 67.100 ;
        RECT 110.200 63.800 110.600 64.200 ;
        RECT 109.400 62.800 109.800 63.200 ;
        RECT 111.000 60.800 111.400 61.200 ;
        RECT 111.000 59.200 111.300 60.800 ;
        RECT 108.600 58.800 109.000 59.200 ;
        RECT 111.000 58.800 111.400 59.200 ;
        RECT 107.000 57.100 107.400 57.200 ;
        RECT 107.800 57.100 108.200 57.200 ;
        RECT 107.000 56.800 108.200 57.100 ;
        RECT 109.400 56.800 109.800 57.200 ;
        RECT 109.400 56.200 109.700 56.800 ;
        RECT 111.800 56.200 112.100 66.800 ;
        RECT 112.600 65.800 113.000 66.200 ;
        RECT 103.000 56.100 103.400 56.200 ;
        RECT 103.800 56.100 104.200 56.200 ;
        RECT 103.000 55.800 104.200 56.100 ;
        RECT 104.600 55.800 105.000 56.200 ;
        RECT 105.400 55.800 105.800 56.200 ;
        RECT 107.000 55.800 107.400 56.200 ;
        RECT 109.400 55.800 109.800 56.200 ;
        RECT 111.800 55.800 112.200 56.200 ;
        RECT 95.000 50.800 95.400 51.200 ;
        RECT 94.200 49.800 94.600 50.200 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 90.200 46.800 90.600 47.200 ;
        RECT 87.800 46.200 88.100 46.800 ;
        RECT 87.800 45.800 88.200 46.200 ;
        RECT 90.200 44.200 90.500 46.800 ;
        RECT 90.200 43.800 90.600 44.200 ;
        RECT 89.400 36.800 89.800 37.200 ;
        RECT 89.400 35.200 89.700 36.800 ;
        RECT 86.200 34.800 86.600 35.200 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 86.200 29.200 86.500 34.800 ;
        RECT 87.000 34.200 87.300 34.800 ;
        RECT 87.000 33.800 87.400 34.200 ;
        RECT 86.200 28.800 86.600 29.200 ;
        RECT 84.600 25.800 85.000 26.200 ;
        RECT 84.600 25.200 84.900 25.800 ;
        RECT 84.600 24.800 85.000 25.200 ;
        RECT 78.200 23.800 78.600 24.200 ;
        RECT 83.000 23.800 83.400 24.200 ;
        RECT 78.200 19.200 78.500 23.800 ;
        RECT 88.600 23.100 89.000 28.900 ;
        RECT 90.200 26.200 90.500 43.800 ;
        RECT 91.000 43.100 91.400 48.900 ;
        RECT 92.600 45.100 93.000 47.900 ;
        RECT 94.200 47.200 94.500 49.800 ;
        RECT 95.000 48.200 95.300 50.800 ;
        RECT 101.400 49.800 101.800 50.200 ;
        RECT 99.800 48.800 100.200 49.200 ;
        RECT 95.000 47.800 95.400 48.200 ;
        RECT 95.000 47.200 95.300 47.800 ;
        RECT 99.800 47.200 100.100 48.800 ;
        RECT 94.200 46.800 94.600 47.200 ;
        RECT 95.000 46.800 95.400 47.200 ;
        RECT 97.400 47.100 97.800 47.200 ;
        RECT 98.200 47.100 98.600 47.200 ;
        RECT 97.400 46.800 98.600 47.100 ;
        RECT 99.800 46.800 100.200 47.200 ;
        RECT 95.800 46.100 96.200 46.200 ;
        RECT 96.600 46.100 97.000 46.200 ;
        RECT 95.800 45.800 97.000 46.100 ;
        RECT 98.200 45.800 98.600 46.200 ;
        RECT 98.200 45.200 98.500 45.800 ;
        RECT 98.200 44.800 98.600 45.200 ;
        RECT 100.600 45.100 101.000 47.900 ;
        RECT 101.400 47.200 101.700 49.800 ;
        RECT 101.400 46.800 101.800 47.200 ;
        RECT 98.200 39.200 98.500 44.800 ;
        RECT 99.000 43.800 99.400 44.200 ;
        RECT 98.200 38.800 98.600 39.200 ;
        RECT 91.000 31.800 91.400 32.200 ;
        RECT 91.800 32.100 92.200 37.900 ;
        RECT 95.800 36.800 96.200 37.200 ;
        RECT 95.800 35.100 96.100 36.800 ;
        RECT 95.800 34.700 96.200 35.100 ;
        RECT 96.600 32.100 97.000 37.900 ;
        RECT 97.400 33.800 97.800 34.200 ;
        RECT 97.400 32.200 97.700 33.800 ;
        RECT 98.200 33.100 98.600 35.900 ;
        RECT 99.000 35.200 99.300 43.800 ;
        RECT 102.200 43.100 102.600 48.900 ;
        RECT 103.000 46.800 103.400 47.200 ;
        RECT 103.000 46.300 103.300 46.800 ;
        RECT 103.000 45.900 103.400 46.300 ;
        RECT 103.800 43.200 104.100 55.800 ;
        RECT 104.600 54.200 104.900 55.800 ;
        RECT 107.000 54.200 107.300 55.800 ;
        RECT 112.600 55.200 112.900 65.800 ;
        RECT 111.000 55.100 111.400 55.200 ;
        RECT 111.800 55.100 112.200 55.200 ;
        RECT 111.000 54.800 112.200 55.100 ;
        RECT 112.600 54.800 113.000 55.200 ;
        RECT 104.600 53.800 105.000 54.200 ;
        RECT 107.000 53.800 107.400 54.200 ;
        RECT 111.800 54.100 112.200 54.200 ;
        RECT 111.000 53.800 112.200 54.100 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 107.800 49.200 108.100 52.800 ;
        RECT 111.000 49.200 111.300 53.800 ;
        RECT 106.200 45.800 106.600 46.200 ;
        RECT 103.800 42.800 104.200 43.200 ;
        RECT 104.600 38.800 105.000 39.200 ;
        RECT 103.000 37.800 103.400 38.200 ;
        RECT 103.000 37.200 103.300 37.800 ;
        RECT 103.000 36.800 103.400 37.200 ;
        RECT 104.600 36.200 104.900 38.800 ;
        RECT 100.600 36.100 101.000 36.200 ;
        RECT 101.400 36.100 101.800 36.200 ;
        RECT 100.600 35.800 101.800 36.100 ;
        RECT 103.800 35.800 104.200 36.200 ;
        RECT 104.600 35.800 105.000 36.200 ;
        RECT 99.000 34.800 99.400 35.200 ;
        RECT 99.000 34.200 99.300 34.800 ;
        RECT 99.000 33.800 99.400 34.200 ;
        RECT 100.600 33.200 100.900 35.800 ;
        RECT 103.800 35.200 104.100 35.800 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 103.000 34.100 103.400 34.200 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 103.000 33.800 104.200 34.100 ;
        RECT 100.600 32.800 101.000 33.200 ;
        RECT 97.400 31.800 97.800 32.200 ;
        RECT 91.000 26.200 91.300 31.800 ;
        RECT 97.400 30.800 97.800 31.200 ;
        RECT 97.400 29.200 97.700 30.800 ;
        RECT 99.800 29.800 100.200 30.200 ;
        RECT 99.800 29.200 100.100 29.800 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 90.200 26.100 90.600 26.200 ;
        RECT 89.400 25.800 90.600 26.100 ;
        RECT 91.000 25.800 91.400 26.200 ;
        RECT 81.400 21.800 81.800 22.200 ;
        RECT 79.800 20.800 80.200 21.200 ;
        RECT 79.800 19.200 80.100 20.800 ;
        RECT 81.400 19.200 81.700 21.800 ;
        RECT 78.200 18.800 78.600 19.200 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 81.400 18.800 81.800 19.200 ;
        RECT 72.600 13.800 73.000 14.200 ;
        RECT 71.800 12.800 72.200 13.200 ;
        RECT 61.400 9.800 61.800 10.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 48.600 6.800 49.000 7.200 ;
        RECT 37.400 5.800 37.800 6.200 ;
        RECT 41.400 5.800 41.800 6.200 ;
        RECT 47.800 5.800 48.200 6.200 ;
        RECT 41.400 5.200 41.700 5.800 ;
        RECT 47.800 5.200 48.100 5.800 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 45.400 5.100 45.800 5.200 ;
        RECT 46.200 5.100 46.600 5.200 ;
        RECT 45.400 4.800 46.600 5.100 ;
        RECT 47.800 4.800 48.200 5.200 ;
        RECT 51.800 3.100 52.200 8.900 ;
        RECT 52.600 8.800 53.000 9.200 ;
        RECT 55.800 8.800 56.200 9.200 ;
        RECT 52.600 6.200 52.900 8.800 ;
        RECT 55.800 6.300 56.100 8.800 ;
        RECT 52.600 5.800 53.000 6.200 ;
        RECT 55.800 5.900 56.200 6.300 ;
        RECT 56.600 3.100 57.000 8.900 ;
        RECT 59.000 8.800 59.400 9.200 ;
        RECT 67.800 9.100 68.200 9.200 ;
        RECT 68.600 9.100 69.000 9.200 ;
        RECT 58.200 5.100 58.600 7.900 ;
        RECT 59.000 5.100 59.400 7.900 ;
        RECT 60.600 3.100 61.000 8.900 ;
        RECT 64.600 7.800 65.000 8.200 ;
        RECT 64.600 7.200 64.900 7.800 ;
        RECT 64.600 6.800 65.000 7.200 ;
        RECT 62.200 5.800 62.600 6.200 ;
        RECT 62.200 5.200 62.500 5.800 ;
        RECT 62.200 4.800 62.600 5.200 ;
        RECT 65.400 3.100 65.800 8.900 ;
        RECT 67.800 8.800 69.000 9.100 ;
        RECT 68.600 5.100 69.000 7.900 ;
        RECT 69.400 7.800 69.800 8.200 ;
        RECT 69.400 7.200 69.700 7.800 ;
        RECT 69.400 6.800 69.800 7.200 ;
        RECT 70.200 3.100 70.600 8.900 ;
        RECT 71.800 7.200 72.100 12.800 ;
        RECT 75.800 12.100 76.200 17.900 ;
        RECT 77.400 17.800 77.800 18.200 ;
        RECT 82.200 17.800 82.600 18.200 ;
        RECT 90.200 17.800 90.600 18.200 ;
        RECT 82.200 14.200 82.500 17.800 ;
        RECT 83.000 16.800 83.400 17.200 ;
        RECT 85.400 16.800 85.800 17.200 ;
        RECT 83.000 15.200 83.300 16.800 ;
        RECT 85.400 16.200 85.700 16.800 ;
        RECT 85.400 15.800 85.800 16.200 ;
        RECT 83.000 14.800 83.400 15.200 ;
        RECT 85.400 14.800 85.800 15.200 ;
        RECT 85.400 14.200 85.700 14.800 ;
        RECT 76.600 14.100 77.000 14.200 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 76.600 13.800 77.800 14.100 ;
        RECT 79.000 14.100 79.400 14.200 ;
        RECT 79.800 14.100 80.200 14.200 ;
        RECT 79.000 13.800 80.200 14.100 ;
        RECT 80.600 14.100 81.000 14.200 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 80.600 13.800 81.800 14.100 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 85.400 13.800 85.800 14.200 ;
        RECT 88.600 13.800 89.000 14.200 ;
        RECT 77.400 9.800 77.800 10.200 ;
        RECT 77.400 9.200 77.700 9.800 ;
        RECT 79.000 9.200 79.300 13.800 ;
        RECT 79.800 11.800 80.200 12.200 ;
        RECT 72.600 7.800 73.000 8.200 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 72.600 6.200 72.900 7.800 ;
        RECT 72.600 5.800 73.000 6.200 ;
        RECT 75.000 3.100 75.400 8.900 ;
        RECT 77.400 8.800 77.800 9.200 ;
        RECT 79.000 8.800 79.400 9.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 78.200 7.200 78.500 7.800 ;
        RECT 79.800 7.200 80.100 11.800 ;
        RECT 80.600 10.200 80.900 13.800 ;
        RECT 88.600 13.200 88.900 13.800 ;
        RECT 88.600 12.800 89.000 13.200 ;
        RECT 89.400 13.100 89.800 15.900 ;
        RECT 81.400 12.100 81.800 12.200 ;
        RECT 81.400 11.800 82.500 12.100 ;
        RECT 80.600 9.800 81.000 10.200 ;
        RECT 82.200 7.200 82.500 11.800 ;
        RECT 90.200 7.200 90.500 17.800 ;
        RECT 91.000 12.100 91.400 17.900 ;
        RECT 91.800 14.200 92.100 26.800 ;
        RECT 93.400 23.100 93.800 28.900 ;
        RECT 97.400 28.800 97.800 29.200 ;
        RECT 99.800 28.800 100.200 29.200 ;
        RECT 100.600 29.100 101.000 29.200 ;
        RECT 101.400 29.100 101.800 29.200 ;
        RECT 100.600 28.800 101.800 29.100 ;
        RECT 95.000 25.100 95.400 27.900 ;
        RECT 95.800 27.800 96.200 28.200 ;
        RECT 104.600 28.100 104.900 35.800 ;
        RECT 106.200 34.200 106.500 45.800 ;
        RECT 107.000 43.100 107.400 48.900 ;
        RECT 107.800 48.800 108.200 49.200 ;
        RECT 108.600 49.100 109.000 49.200 ;
        RECT 109.400 49.100 109.800 49.200 ;
        RECT 108.600 48.800 109.800 49.100 ;
        RECT 111.000 48.800 111.400 49.200 ;
        RECT 113.400 48.200 113.700 69.800 ;
        RECT 114.200 67.200 114.500 69.800 ;
        RECT 115.800 68.200 116.100 91.800 ;
        RECT 117.400 90.200 117.700 91.800 ;
        RECT 117.400 89.800 117.800 90.200 ;
        RECT 117.400 88.800 117.800 89.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 116.600 85.200 116.900 85.800 ;
        RECT 117.400 85.200 117.700 88.800 ;
        RECT 118.200 86.800 118.600 87.200 ;
        RECT 116.600 84.800 117.000 85.200 ;
        RECT 117.400 84.800 117.800 85.200 ;
        RECT 118.200 84.100 118.500 86.800 ;
        RECT 119.000 86.200 119.300 97.800 ;
        RECT 119.800 94.800 120.200 95.200 ;
        RECT 119.800 94.200 120.100 94.800 ;
        RECT 121.400 94.200 121.700 105.800 ;
        RECT 122.200 97.200 122.500 105.800 ;
        RECT 124.600 105.200 124.900 108.800 ;
        RECT 128.600 108.200 128.900 126.800 ;
        RECT 129.400 126.100 129.800 126.200 ;
        RECT 130.200 126.100 130.600 126.200 ;
        RECT 129.400 125.800 130.600 126.100 ;
        RECT 131.800 123.100 132.200 128.900 ;
        RECT 133.400 128.800 134.600 129.100 ;
        RECT 134.200 128.200 134.500 128.800 ;
        RECT 134.200 127.800 134.600 128.200 ;
        RECT 135.000 125.200 135.300 131.800 ;
        RECT 137.400 127.200 137.700 143.800 ;
        RECT 141.400 142.200 141.700 145.800 ;
        RECT 143.800 144.800 144.200 145.200 ;
        RECT 143.800 142.200 144.100 144.800 ;
        RECT 141.400 141.800 141.800 142.200 ;
        RECT 143.800 141.800 144.200 142.200 ;
        RECT 143.000 136.800 143.400 137.200 ;
        RECT 143.000 136.200 143.300 136.800 ;
        RECT 140.600 136.100 141.000 136.200 ;
        RECT 141.400 136.100 141.800 136.200 ;
        RECT 140.600 135.800 141.800 136.100 ;
        RECT 143.000 135.800 143.400 136.200 ;
        RECT 143.800 135.200 144.100 141.800 ;
        RECT 144.600 138.200 144.900 151.800 ;
        RECT 145.400 150.800 145.800 151.200 ;
        RECT 145.400 147.200 145.700 150.800 ;
        RECT 147.800 147.800 148.200 148.200 ;
        RECT 147.800 147.200 148.100 147.800 ;
        RECT 148.600 147.200 148.900 152.800 ;
        RECT 149.400 150.200 149.700 154.800 ;
        RECT 153.400 153.200 153.700 165.800 ;
        RECT 154.200 162.200 154.500 165.800 ;
        RECT 157.400 165.200 157.700 165.800 ;
        RECT 155.000 164.800 155.400 165.200 ;
        RECT 157.400 164.800 157.800 165.200 ;
        RECT 158.200 165.100 158.600 167.900 ;
        RECT 159.000 167.800 159.400 168.200 ;
        RECT 159.000 167.200 159.300 167.800 ;
        RECT 159.000 166.800 159.400 167.200 ;
        RECT 154.200 161.800 154.600 162.200 ;
        RECT 155.000 155.200 155.300 164.800 ;
        RECT 155.800 163.800 156.200 164.200 ;
        RECT 155.000 154.800 155.400 155.200 ;
        RECT 155.800 154.200 156.100 163.800 ;
        RECT 159.800 163.100 160.200 168.900 ;
        RECT 161.400 166.800 161.800 167.200 ;
        RECT 161.400 166.200 161.700 166.800 ;
        RECT 161.400 165.800 161.800 166.200 ;
        RECT 164.600 163.100 165.000 168.900 ;
        RECT 166.200 168.200 166.500 172.800 ;
        RECT 166.200 167.800 166.600 168.200 ;
        RECT 167.000 166.200 167.300 181.800 ;
        RECT 170.200 172.100 170.600 177.900 ;
        RECT 171.000 177.200 171.300 185.800 ;
        RECT 174.200 183.100 174.600 188.900 ;
        RECT 175.800 185.100 176.200 187.900 ;
        RECT 176.600 187.800 177.000 188.200 ;
        RECT 176.600 187.200 176.900 187.800 ;
        RECT 176.600 186.800 177.000 187.200 ;
        RECT 175.800 180.800 176.200 181.200 ;
        RECT 175.800 179.200 176.100 180.800 ;
        RECT 175.800 178.800 176.200 179.200 ;
        RECT 171.000 176.800 171.400 177.200 ;
        RECT 171.800 177.100 172.200 177.200 ;
        RECT 172.600 177.100 173.000 177.200 ;
        RECT 171.800 176.800 173.000 177.100 ;
        RECT 176.600 176.800 177.000 177.200 ;
        RECT 176.600 175.200 176.900 176.800 ;
        RECT 173.400 174.800 173.800 175.200 ;
        RECT 174.200 174.800 174.600 175.200 ;
        RECT 176.600 174.800 177.000 175.200 ;
        RECT 177.400 175.100 177.700 201.800 ;
        RECT 182.200 200.800 182.600 201.200 ;
        RECT 180.600 197.800 181.000 198.200 ;
        RECT 179.000 195.800 179.400 196.200 ;
        RECT 179.000 195.200 179.300 195.800 ;
        RECT 179.000 194.800 179.400 195.200 ;
        RECT 179.000 193.200 179.300 194.800 ;
        RECT 180.600 194.200 180.900 197.800 ;
        RECT 182.200 195.200 182.500 200.800 ;
        RECT 182.200 194.800 182.600 195.200 ;
        RECT 180.600 193.800 181.000 194.200 ;
        RECT 179.000 192.800 179.400 193.200 ;
        RECT 178.200 188.100 178.600 188.200 ;
        RECT 179.000 188.100 179.400 188.200 ;
        RECT 178.200 187.800 179.400 188.100 ;
        RECT 180.600 187.200 180.900 193.800 ;
        RECT 181.400 191.800 181.800 192.200 ;
        RECT 181.400 187.200 181.700 191.800 ;
        RECT 183.000 190.200 183.300 204.800 ;
        RECT 186.200 201.800 186.600 202.200 ;
        RECT 186.200 200.200 186.500 201.800 ;
        RECT 186.200 199.800 186.600 200.200 ;
        RECT 192.600 196.800 193.000 197.200 ;
        RECT 192.600 196.200 192.900 196.800 ;
        RECT 184.600 195.800 185.000 196.200 ;
        RECT 189.400 195.800 189.800 196.200 ;
        RECT 192.600 195.800 193.000 196.200 ;
        RECT 184.600 195.200 184.900 195.800 ;
        RECT 189.400 195.200 189.700 195.800 ;
        RECT 184.600 194.800 185.000 195.200 ;
        RECT 185.400 194.800 185.800 195.200 ;
        RECT 186.200 195.100 186.600 195.200 ;
        RECT 187.000 195.100 187.400 195.200 ;
        RECT 186.200 194.800 187.400 195.100 ;
        RECT 189.400 194.800 189.800 195.200 ;
        RECT 185.400 194.200 185.700 194.800 ;
        RECT 192.600 194.200 192.900 195.800 ;
        RECT 185.400 193.800 185.800 194.200 ;
        RECT 186.200 193.800 186.600 194.200 ;
        RECT 188.600 194.100 189.000 194.200 ;
        RECT 189.400 194.100 189.800 194.200 ;
        RECT 188.600 193.800 189.800 194.100 ;
        RECT 192.600 193.800 193.000 194.200 ;
        RECT 186.200 192.200 186.500 193.800 ;
        RECT 183.800 191.800 184.200 192.200 ;
        RECT 186.200 191.800 186.600 192.200 ;
        RECT 195.800 192.100 196.200 197.900 ;
        RECT 196.600 196.200 196.900 205.800 ;
        RECT 199.800 201.800 200.200 202.200 ;
        RECT 196.600 195.800 197.000 196.200 ;
        RECT 196.600 195.200 196.900 195.800 ;
        RECT 196.600 194.800 197.000 195.200 ;
        RECT 199.000 194.800 199.400 195.200 ;
        RECT 199.000 194.200 199.300 194.800 ;
        RECT 199.000 193.800 199.400 194.200 ;
        RECT 183.000 189.800 183.400 190.200 ;
        RECT 183.800 188.200 184.100 191.800 ;
        RECT 186.200 189.800 186.600 190.200 ;
        RECT 183.800 187.800 184.200 188.200 ;
        RECT 180.600 186.800 181.000 187.200 ;
        RECT 181.400 186.800 181.800 187.200 ;
        RECT 183.000 186.800 183.400 187.200 ;
        RECT 184.600 187.100 185.000 187.200 ;
        RECT 185.400 187.100 185.800 187.200 ;
        RECT 184.600 186.800 185.800 187.100 ;
        RECT 178.200 185.800 178.600 186.200 ;
        RECT 179.800 186.100 180.200 186.200 ;
        RECT 180.600 186.100 181.000 186.200 ;
        RECT 179.800 185.800 181.000 186.100 ;
        RECT 178.200 185.200 178.500 185.800 ;
        RECT 178.200 184.800 178.600 185.200 ;
        RECT 178.200 175.100 178.600 175.200 ;
        RECT 177.400 174.800 178.600 175.100 ;
        RECT 172.600 167.800 173.000 168.200 ;
        RECT 172.600 167.200 172.900 167.800 ;
        RECT 167.800 166.800 168.200 167.200 ;
        RECT 169.400 167.100 169.800 167.200 ;
        RECT 170.200 167.100 170.600 167.200 ;
        RECT 169.400 166.800 170.600 167.100 ;
        RECT 172.600 166.800 173.000 167.200 ;
        RECT 167.000 165.800 167.400 166.200 ;
        RECT 167.800 164.200 168.100 166.800 ;
        RECT 171.800 165.800 172.200 166.200 ;
        RECT 171.800 165.200 172.100 165.800 ;
        RECT 168.600 165.100 169.000 165.200 ;
        RECT 169.400 165.100 169.800 165.200 ;
        RECT 168.600 164.800 169.800 165.100 ;
        RECT 171.800 164.800 172.200 165.200 ;
        RECT 167.800 163.800 168.200 164.200 ;
        RECT 167.800 160.200 168.100 163.800 ;
        RECT 167.800 159.800 168.200 160.200 ;
        RECT 158.200 157.100 158.600 157.200 ;
        RECT 159.000 157.100 159.400 157.200 ;
        RECT 158.200 156.800 159.400 157.100 ;
        RECT 160.600 156.800 161.000 157.200 ;
        RECT 160.600 156.200 160.900 156.800 ;
        RECT 156.600 155.800 157.000 156.200 ;
        RECT 157.400 155.800 157.800 156.200 ;
        RECT 159.800 155.800 160.200 156.200 ;
        RECT 160.600 155.800 161.000 156.200 ;
        RECT 156.600 155.200 156.900 155.800 ;
        RECT 156.600 154.800 157.000 155.200 ;
        RECT 157.400 154.200 157.700 155.800 ;
        RECT 159.800 155.200 160.100 155.800 ;
        RECT 159.800 154.800 160.200 155.200 ;
        RECT 155.000 154.100 155.400 154.200 ;
        RECT 155.800 154.100 156.200 154.200 ;
        RECT 155.000 153.800 156.200 154.100 ;
        RECT 157.400 153.800 157.800 154.200 ;
        RECT 151.800 152.800 152.200 153.200 ;
        RECT 153.400 152.800 153.800 153.200 ;
        RECT 151.800 152.200 152.100 152.800 ;
        RECT 151.000 151.800 151.400 152.200 ;
        RECT 151.800 151.800 152.200 152.200 ;
        RECT 153.400 151.800 153.800 152.200 ;
        RECT 149.400 149.800 149.800 150.200 ;
        RECT 149.400 148.200 149.700 149.800 ;
        RECT 149.400 147.800 149.800 148.200 ;
        RECT 145.400 146.800 145.800 147.200 ;
        RECT 146.200 147.100 146.600 147.200 ;
        RECT 147.000 147.100 147.400 147.200 ;
        RECT 146.200 146.800 147.400 147.100 ;
        RECT 147.800 146.800 148.200 147.200 ;
        RECT 148.600 146.800 149.000 147.200 ;
        RECT 151.000 147.100 151.300 151.800 ;
        RECT 153.400 149.200 153.700 151.800 ;
        RECT 155.000 150.800 155.400 151.200 ;
        RECT 157.400 150.800 157.800 151.200 ;
        RECT 153.400 148.800 153.800 149.200 ;
        RECT 154.200 148.800 154.600 149.200 ;
        RECT 154.200 148.200 154.500 148.800 ;
        RECT 154.200 147.800 154.600 148.200 ;
        RECT 151.000 146.800 152.100 147.100 ;
        RECT 145.400 145.800 145.800 146.200 ;
        RECT 148.600 146.100 149.000 146.200 ;
        RECT 149.400 146.100 149.800 146.200 ;
        RECT 148.600 145.800 149.800 146.100 ;
        RECT 150.200 146.100 150.600 146.200 ;
        RECT 151.000 146.100 151.400 146.200 ;
        RECT 150.200 145.800 151.400 146.100 ;
        RECT 145.400 145.200 145.700 145.800 ;
        RECT 145.400 144.800 145.800 145.200 ;
        RECT 149.400 145.100 149.800 145.200 ;
        RECT 150.200 145.100 150.600 145.200 ;
        RECT 149.400 144.800 150.600 145.100 ;
        RECT 151.800 144.200 152.100 146.800 ;
        RECT 155.000 146.200 155.300 150.800 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 156.600 145.800 157.000 146.200 ;
        RECT 156.600 145.200 156.900 145.800 ;
        RECT 156.600 144.800 157.000 145.200 ;
        RECT 151.800 143.800 152.200 144.200 ;
        RECT 154.200 143.800 154.600 144.200 ;
        RECT 152.600 142.100 153.000 142.200 ;
        RECT 153.400 142.100 153.800 142.200 ;
        RECT 152.600 141.800 153.800 142.100 ;
        RECT 147.000 140.800 147.400 141.200 ;
        RECT 144.600 137.800 145.000 138.200 ;
        RECT 147.000 136.200 147.300 140.800 ;
        RECT 153.400 139.800 153.800 140.200 ;
        RECT 153.400 139.200 153.700 139.800 ;
        RECT 153.400 138.800 153.800 139.200 ;
        RECT 144.600 135.800 145.000 136.200 ;
        RECT 147.000 135.800 147.400 136.200 ;
        RECT 147.800 136.100 148.200 136.200 ;
        RECT 148.600 136.100 149.000 136.200 ;
        RECT 147.800 135.800 149.000 136.100 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 139.000 135.100 139.400 135.200 ;
        RECT 138.200 134.800 139.400 135.100 ;
        RECT 143.000 134.800 143.400 135.200 ;
        RECT 143.800 134.800 144.200 135.200 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 139.000 134.100 139.400 134.200 ;
        RECT 138.200 133.800 139.400 134.100 ;
        RECT 143.000 133.200 143.300 134.800 ;
        RECT 144.600 134.200 144.900 135.800 ;
        RECT 145.400 134.800 145.800 135.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 144.600 133.800 145.000 134.200 ;
        RECT 143.800 133.200 144.100 133.800 ;
        RECT 143.000 132.800 143.400 133.200 ;
        RECT 143.800 132.800 144.200 133.200 ;
        RECT 138.200 131.800 138.600 132.200 ;
        RECT 138.200 131.200 138.500 131.800 ;
        RECT 138.200 130.800 138.600 131.200 ;
        RECT 141.400 129.100 141.800 129.200 ;
        RECT 142.200 129.100 142.600 129.200 ;
        RECT 141.400 128.800 142.600 129.100 ;
        RECT 138.200 127.800 138.600 128.200 ;
        RECT 138.200 127.200 138.500 127.800 ;
        RECT 135.800 126.800 136.200 127.200 ;
        RECT 137.400 126.800 137.800 127.200 ;
        RECT 138.200 126.800 138.600 127.200 ;
        RECT 135.800 126.200 136.100 126.800 ;
        RECT 135.800 125.800 136.200 126.200 ;
        RECT 136.600 125.800 137.000 126.200 ;
        RECT 136.600 125.200 136.900 125.800 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 136.600 124.800 137.000 125.200 ;
        RECT 135.000 119.800 135.400 120.200 ;
        RECT 131.000 116.800 131.400 117.200 ;
        RECT 131.000 115.200 131.300 116.800 ;
        RECT 131.000 114.800 131.400 115.200 ;
        RECT 129.400 111.800 129.800 112.200 ;
        RECT 133.400 112.100 133.800 117.900 ;
        RECT 129.400 110.200 129.700 111.800 ;
        RECT 129.400 109.800 129.800 110.200 ;
        RECT 126.200 106.800 126.600 107.200 ;
        RECT 127.000 106.800 127.400 107.200 ;
        RECT 126.200 106.200 126.500 106.800 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 124.600 104.800 125.000 105.200 ;
        RECT 126.200 104.800 126.600 105.200 ;
        RECT 126.200 104.200 126.500 104.800 ;
        RECT 126.200 103.800 126.600 104.200 ;
        RECT 127.000 101.200 127.300 106.800 ;
        RECT 127.800 105.100 128.200 107.900 ;
        RECT 128.600 107.800 129.000 108.200 ;
        RECT 128.600 107.200 128.900 107.800 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 129.400 103.100 129.800 108.900 ;
        RECT 131.000 107.800 131.400 108.200 ;
        RECT 131.000 106.200 131.300 107.800 ;
        RECT 131.000 105.800 131.400 106.200 ;
        RECT 134.200 103.100 134.600 108.900 ;
        RECT 127.000 100.800 127.400 101.200 ;
        RECT 129.400 100.800 129.800 101.200 ;
        RECT 129.400 99.200 129.700 100.800 ;
        RECT 129.400 98.800 129.800 99.200 ;
        RECT 123.000 97.800 123.400 98.200 ;
        RECT 122.200 96.800 122.600 97.200 ;
        RECT 122.200 95.200 122.500 96.800 ;
        RECT 123.000 96.200 123.300 97.800 ;
        RECT 123.000 95.800 123.400 96.200 ;
        RECT 124.600 95.800 125.000 96.200 ;
        RECT 128.600 95.800 129.000 96.200 ;
        RECT 131.000 95.800 131.400 96.200 ;
        RECT 132.600 95.800 133.000 96.200 ;
        RECT 124.600 95.200 124.900 95.800 ;
        RECT 128.600 95.200 128.900 95.800 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 124.600 94.800 125.000 95.200 ;
        RECT 127.800 94.800 128.200 95.200 ;
        RECT 128.600 94.800 129.000 95.200 ;
        RECT 127.800 94.200 128.100 94.800 ;
        RECT 119.800 93.800 120.200 94.200 ;
        RECT 121.400 93.800 121.800 94.200 ;
        RECT 125.400 93.800 125.800 94.200 ;
        RECT 126.200 93.800 126.600 94.200 ;
        RECT 127.800 93.800 128.200 94.200 ;
        RECT 120.600 92.800 121.000 93.200 ;
        RECT 120.600 92.200 120.900 92.800 ;
        RECT 120.600 91.800 121.000 92.200 ;
        RECT 123.800 91.800 124.200 92.200 ;
        RECT 120.600 89.100 121.000 89.200 ;
        RECT 121.400 89.100 121.800 89.200 ;
        RECT 120.600 88.800 121.800 89.100 ;
        RECT 120.600 87.800 121.000 88.200 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 120.600 85.200 120.900 87.800 ;
        RECT 120.600 84.800 121.000 85.200 ;
        RECT 121.400 85.100 121.800 87.900 ;
        RECT 117.400 83.800 118.500 84.100 ;
        RECT 117.400 79.200 117.700 83.800 ;
        RECT 123.000 83.100 123.400 88.900 ;
        RECT 123.800 88.200 124.100 91.800 ;
        RECT 125.400 89.200 125.700 93.800 ;
        RECT 126.200 93.200 126.500 93.800 ;
        RECT 126.200 92.800 126.600 93.200 ;
        RECT 130.200 92.800 130.600 93.200 ;
        RECT 130.200 92.200 130.500 92.800 ;
        RECT 127.000 91.800 127.400 92.200 ;
        RECT 130.200 91.800 130.600 92.200 ;
        RECT 124.600 88.800 125.000 89.200 ;
        RECT 125.400 88.800 125.800 89.200 ;
        RECT 123.800 87.800 124.200 88.200 ;
        RECT 124.600 86.200 124.900 88.800 ;
        RECT 126.200 86.800 126.600 87.200 ;
        RECT 126.200 86.200 126.500 86.800 ;
        RECT 124.600 85.800 125.000 86.200 ;
        RECT 126.200 85.800 126.600 86.200 ;
        RECT 117.400 78.800 117.800 79.200 ;
        RECT 118.200 76.800 118.600 77.200 ;
        RECT 117.400 72.800 117.800 73.200 ;
        RECT 117.400 72.200 117.700 72.800 ;
        RECT 117.400 71.800 117.800 72.200 ;
        RECT 115.800 67.800 116.200 68.200 ;
        RECT 114.200 66.800 114.600 67.200 ;
        RECT 116.600 67.100 117.000 67.200 ;
        RECT 117.400 67.100 117.800 67.200 ;
        RECT 116.600 66.800 117.800 67.100 ;
        RECT 114.200 65.200 114.500 66.800 ;
        RECT 118.200 66.200 118.500 76.800 ;
        RECT 119.800 75.800 120.200 76.200 ;
        RECT 120.600 76.100 121.000 76.200 ;
        RECT 121.400 76.100 121.800 76.200 ;
        RECT 120.600 75.800 121.800 76.100 ;
        RECT 119.800 75.200 120.100 75.800 ;
        RECT 119.800 74.800 120.200 75.200 ;
        RECT 123.800 75.100 124.200 75.200 ;
        RECT 124.600 75.100 125.000 75.200 ;
        RECT 123.800 74.800 125.000 75.100 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 119.000 73.800 120.200 74.100 ;
        RECT 122.200 74.100 122.600 74.200 ;
        RECT 123.000 74.100 123.400 74.200 ;
        RECT 122.200 73.800 123.400 74.100 ;
        RECT 125.400 73.100 125.800 75.900 ;
        RECT 126.200 74.200 126.500 85.800 ;
        RECT 127.000 79.200 127.300 91.800 ;
        RECT 131.000 91.100 131.300 95.800 ;
        RECT 132.600 95.200 132.900 95.800 ;
        RECT 132.600 94.800 133.000 95.200 ;
        RECT 132.600 93.800 133.000 94.200 ;
        RECT 132.600 93.200 132.900 93.800 ;
        RECT 132.600 92.800 133.000 93.200 ;
        RECT 130.200 90.800 131.300 91.100 ;
        RECT 131.800 91.800 132.200 92.200 ;
        RECT 130.200 89.200 130.500 90.800 ;
        RECT 131.800 89.200 132.100 91.800 ;
        RECT 129.400 89.100 129.800 89.200 ;
        RECT 130.200 89.100 130.600 89.200 ;
        RECT 127.800 83.100 128.200 88.900 ;
        RECT 129.400 88.800 130.600 89.100 ;
        RECT 131.000 89.100 131.400 89.200 ;
        RECT 131.800 89.100 132.200 89.200 ;
        RECT 131.000 88.800 132.200 89.100 ;
        RECT 133.400 83.100 133.800 88.900 ;
        RECT 134.200 86.800 134.600 87.200 ;
        RECT 134.200 86.200 134.500 86.800 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 127.000 78.800 127.400 79.200 ;
        RECT 126.200 73.800 126.600 74.200 ;
        RECT 121.400 71.800 121.800 72.200 ;
        RECT 127.000 72.100 127.400 77.900 ;
        RECT 130.200 75.800 130.600 76.200 ;
        RECT 130.200 75.200 130.500 75.800 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 131.000 74.800 131.400 75.200 ;
        RECT 119.800 67.800 120.200 68.200 ;
        RECT 119.800 67.200 120.100 67.800 ;
        RECT 121.400 67.200 121.700 71.800 ;
        RECT 125.400 70.800 125.800 71.200 ;
        RECT 125.400 68.200 125.700 70.800 ;
        RECT 129.400 69.800 129.800 70.200 ;
        RECT 129.400 69.200 129.700 69.800 ;
        RECT 129.400 68.800 129.800 69.200 ;
        RECT 125.400 67.800 125.800 68.200 ;
        RECT 127.800 67.800 128.200 68.200 ;
        RECT 119.000 66.800 119.400 67.200 ;
        RECT 119.800 66.800 120.200 67.200 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 123.000 67.100 123.400 67.200 ;
        RECT 123.800 67.100 124.200 67.200 ;
        RECT 123.000 66.800 124.200 67.100 ;
        RECT 126.200 66.800 126.600 67.200 ;
        RECT 115.800 65.800 116.200 66.200 ;
        RECT 118.200 65.800 118.600 66.200 ;
        RECT 115.800 65.200 116.100 65.800 ;
        RECT 114.200 64.800 114.600 65.200 ;
        RECT 115.800 64.800 116.200 65.200 ;
        RECT 115.800 59.200 116.100 64.800 ;
        RECT 116.600 59.800 117.000 60.200 ;
        RECT 115.800 58.800 116.200 59.200 ;
        RECT 115.800 57.800 116.200 58.200 ;
        RECT 115.800 55.200 116.100 57.800 ;
        RECT 116.600 55.200 116.900 59.800 ;
        RECT 117.400 57.100 117.800 57.200 ;
        RECT 118.200 57.100 118.600 57.200 ;
        RECT 117.400 56.800 118.600 57.100 ;
        RECT 115.800 54.800 116.200 55.200 ;
        RECT 116.600 54.800 117.000 55.200 ;
        RECT 110.200 47.800 110.600 48.200 ;
        RECT 113.400 47.800 113.800 48.200 ;
        RECT 109.400 44.800 109.800 45.200 ;
        RECT 109.400 39.200 109.700 44.800 ;
        RECT 110.200 44.200 110.500 47.800 ;
        RECT 115.800 46.200 116.100 54.800 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 115.000 45.800 115.400 46.200 ;
        RECT 115.800 45.800 116.200 46.200 ;
        RECT 116.600 45.800 117.000 46.200 ;
        RECT 117.400 45.800 117.800 46.200 ;
        RECT 112.600 45.200 112.900 45.800 ;
        RECT 112.600 44.800 113.000 45.200 ;
        RECT 110.200 43.800 110.600 44.200 ;
        RECT 113.400 43.100 113.800 43.200 ;
        RECT 114.200 43.100 114.600 43.200 ;
        RECT 113.400 42.800 114.600 43.100 ;
        RECT 115.000 40.200 115.300 45.800 ;
        RECT 115.000 39.800 115.400 40.200 ;
        RECT 116.600 39.200 116.900 45.800 ;
        RECT 117.400 45.200 117.700 45.800 ;
        RECT 117.400 44.800 117.800 45.200 ;
        RECT 118.200 39.200 118.500 53.800 ;
        RECT 119.000 51.200 119.300 66.800 ;
        RECT 120.600 65.800 121.000 66.200 ;
        RECT 120.600 58.200 120.900 65.800 ;
        RECT 122.200 64.800 122.600 65.200 ;
        RECT 122.200 64.200 122.500 64.800 ;
        RECT 122.200 63.800 122.600 64.200 ;
        RECT 126.200 63.200 126.500 66.800 ;
        RECT 127.800 65.200 128.100 67.800 ;
        RECT 128.600 66.800 129.000 67.200 ;
        RECT 128.600 66.200 128.900 66.800 ;
        RECT 128.600 65.800 129.000 66.200 ;
        RECT 127.800 65.100 128.200 65.200 ;
        RECT 128.600 65.100 129.000 65.200 ;
        RECT 127.800 64.800 129.000 65.100 ;
        RECT 131.000 64.200 131.300 74.800 ;
        RECT 131.800 72.100 132.200 77.900 ;
        RECT 135.000 75.200 135.300 119.800 ;
        RECT 135.800 106.800 136.200 107.200 ;
        RECT 135.800 103.200 136.100 106.800 ;
        RECT 136.600 106.100 136.900 124.800 ;
        RECT 137.400 121.200 137.700 126.800 ;
        RECT 143.000 126.200 143.300 132.800 ;
        RECT 145.400 131.200 145.700 134.800 ;
        RECT 146.200 133.800 146.600 134.200 ;
        RECT 145.400 130.800 145.800 131.200 ;
        RECT 145.400 128.800 145.800 129.200 ;
        RECT 144.600 127.800 145.000 128.200 ;
        RECT 144.600 127.200 144.900 127.800 ;
        RECT 145.400 127.200 145.700 128.800 ;
        RECT 143.800 126.800 144.200 127.200 ;
        RECT 144.600 126.800 145.000 127.200 ;
        RECT 145.400 126.800 145.800 127.200 ;
        RECT 143.800 126.200 144.100 126.800 ;
        RECT 142.200 125.800 142.600 126.200 ;
        RECT 143.000 125.800 143.400 126.200 ;
        RECT 143.800 125.800 144.200 126.200 ;
        RECT 139.000 125.100 139.400 125.200 ;
        RECT 139.800 125.100 140.200 125.200 ;
        RECT 139.000 124.800 140.200 125.100 ;
        RECT 141.400 124.800 141.800 125.200 ;
        RECT 141.400 124.200 141.700 124.800 ;
        RECT 142.200 124.200 142.500 125.800 ;
        RECT 146.200 125.100 146.500 133.800 ;
        RECT 147.000 133.200 147.300 135.800 ;
        RECT 153.400 134.800 153.800 135.200 ;
        RECT 153.400 134.200 153.700 134.800 ;
        RECT 153.400 133.800 153.800 134.200 ;
        RECT 147.000 132.800 147.400 133.200 ;
        RECT 148.600 132.800 149.000 133.200 ;
        RECT 148.600 130.200 148.900 132.800 ;
        RECT 149.400 132.100 149.800 132.200 ;
        RECT 150.200 132.100 150.600 132.200 ;
        RECT 149.400 131.800 150.600 132.100 ;
        RECT 148.600 129.800 149.000 130.200 ;
        RECT 152.600 129.800 153.000 130.200 ;
        RECT 152.600 129.200 152.900 129.800 ;
        RECT 152.600 128.800 153.000 129.200 ;
        RECT 151.800 127.800 152.200 128.200 ;
        RECT 151.800 127.200 152.100 127.800 ;
        RECT 147.000 126.800 147.400 127.200 ;
        RECT 151.800 126.800 152.200 127.200 ;
        RECT 147.000 126.200 147.300 126.800 ;
        RECT 147.000 125.800 147.400 126.200 ;
        RECT 149.400 125.800 149.800 126.200 ;
        RECT 147.000 125.100 147.400 125.200 ;
        RECT 146.200 124.800 147.400 125.100 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 147.800 124.200 148.100 124.800 ;
        RECT 141.400 123.800 141.800 124.200 ;
        RECT 142.200 123.800 142.600 124.200 ;
        RECT 147.800 123.800 148.200 124.200 ;
        RECT 137.400 120.800 137.800 121.200 ;
        RECT 137.400 116.800 137.800 117.200 ;
        RECT 137.400 115.100 137.700 116.800 ;
        RECT 137.400 114.700 137.800 115.100 ;
        RECT 138.200 112.100 138.600 117.900 ;
        RECT 139.000 113.800 139.400 114.200 ;
        RECT 139.000 113.200 139.300 113.800 ;
        RECT 139.000 112.800 139.400 113.200 ;
        RECT 139.800 113.100 140.200 115.900 ;
        RECT 137.400 109.800 137.800 110.200 ;
        RECT 137.400 107.200 137.700 109.800 ;
        RECT 141.400 109.200 141.700 123.800 ;
        RECT 143.800 121.800 144.200 122.200 ;
        RECT 146.200 121.800 146.600 122.200 ;
        RECT 143.800 116.200 144.100 121.800 ;
        RECT 146.200 119.200 146.500 121.800 ;
        RECT 146.200 118.800 146.600 119.200 ;
        RECT 144.600 116.800 145.000 117.200 ;
        RECT 143.800 115.800 144.200 116.200 ;
        RECT 142.200 114.800 142.600 115.200 ;
        RECT 142.200 114.200 142.500 114.800 ;
        RECT 144.600 114.200 144.900 116.800 ;
        RECT 146.200 115.800 146.600 116.200 ;
        RECT 146.200 115.200 146.500 115.800 ;
        RECT 149.400 115.200 149.700 125.800 ;
        RECT 153.400 120.200 153.700 133.800 ;
        RECT 153.400 119.800 153.800 120.200 ;
        RECT 152.600 116.100 153.000 116.200 ;
        RECT 153.400 116.100 153.800 116.200 ;
        RECT 152.600 115.800 153.800 116.100 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 147.800 114.800 148.200 115.200 ;
        RECT 149.400 114.800 149.800 115.200 ;
        RECT 151.000 115.100 151.400 115.200 ;
        RECT 151.800 115.100 152.200 115.200 ;
        RECT 151.000 114.800 152.200 115.100 ;
        RECT 142.200 113.800 142.600 114.200 ;
        RECT 144.600 113.800 145.000 114.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 147.000 110.200 147.300 113.800 ;
        RECT 147.800 113.200 148.100 114.800 ;
        RECT 148.600 114.100 149.000 114.200 ;
        RECT 149.400 114.100 149.800 114.200 ;
        RECT 148.600 113.800 149.800 114.100 ;
        RECT 153.400 114.100 153.800 114.200 ;
        RECT 154.200 114.100 154.500 143.800 ;
        RECT 155.800 136.800 156.200 137.200 ;
        RECT 155.800 136.200 156.100 136.800 ;
        RECT 155.800 135.800 156.200 136.200 ;
        RECT 155.000 123.100 155.400 128.900 ;
        RECT 155.800 125.800 156.200 126.200 ;
        RECT 155.800 121.200 156.100 125.800 ;
        RECT 155.800 120.800 156.200 121.200 ;
        RECT 153.400 113.800 154.500 114.100 ;
        RECT 155.000 117.800 155.400 118.200 ;
        RECT 155.000 114.200 155.300 117.800 ;
        RECT 155.800 116.800 156.200 117.200 ;
        RECT 155.800 116.200 156.100 116.800 ;
        RECT 155.800 115.800 156.200 116.200 ;
        RECT 157.400 115.200 157.700 150.800 ;
        RECT 159.000 146.800 159.400 147.200 ;
        RECT 159.000 146.200 159.300 146.800 ;
        RECT 158.200 145.800 158.600 146.200 ;
        RECT 159.000 145.800 159.400 146.200 ;
        RECT 158.200 144.200 158.500 145.800 ;
        RECT 158.200 143.800 158.600 144.200 ;
        RECT 158.200 135.800 158.600 136.200 ;
        RECT 159.800 136.100 160.100 154.800 ;
        RECT 163.000 152.100 163.400 157.900 ;
        RECT 167.000 155.800 167.400 156.200 ;
        RECT 167.000 155.100 167.300 155.800 ;
        RECT 167.000 154.700 167.400 155.100 ;
        RECT 163.800 151.800 164.200 152.200 ;
        RECT 167.800 152.100 168.200 157.900 ;
        RECT 170.200 156.800 170.600 157.200 ;
        RECT 171.800 156.800 172.200 157.200 ;
        RECT 170.200 156.200 170.500 156.800 ;
        RECT 171.800 156.200 172.100 156.800 ;
        RECT 168.600 153.800 169.000 154.200 ;
        RECT 163.800 150.100 164.100 151.800 ;
        RECT 163.000 149.800 164.100 150.100 ;
        RECT 164.600 149.800 165.000 150.200 ;
        RECT 163.000 146.200 163.300 149.800 ;
        RECT 164.600 149.200 164.900 149.800 ;
        RECT 163.800 149.100 164.200 149.200 ;
        RECT 164.600 149.100 165.000 149.200 ;
        RECT 163.800 148.800 165.000 149.100 ;
        RECT 163.800 146.800 164.200 147.200 ;
        RECT 163.800 146.200 164.100 146.800 ;
        RECT 160.600 145.800 161.000 146.200 ;
        RECT 163.000 145.800 163.400 146.200 ;
        RECT 163.800 145.800 164.200 146.200 ;
        RECT 160.600 145.200 160.900 145.800 ;
        RECT 160.600 144.800 161.000 145.200 ;
        RECT 167.000 143.100 167.400 148.900 ;
        RECT 168.600 147.200 168.900 153.800 ;
        RECT 169.400 153.100 169.800 155.900 ;
        RECT 170.200 155.800 170.600 156.200 ;
        RECT 171.800 155.800 172.200 156.200 ;
        RECT 171.000 155.100 171.400 155.200 ;
        RECT 171.800 155.100 172.200 155.200 ;
        RECT 171.000 154.800 172.200 155.100 ;
        RECT 172.600 154.200 172.900 166.800 ;
        RECT 173.400 164.200 173.700 174.800 ;
        RECT 174.200 170.200 174.500 174.800 ;
        RECT 174.200 169.800 174.600 170.200 ;
        RECT 175.800 167.800 176.200 168.200 ;
        RECT 175.000 165.800 175.400 166.200 ;
        RECT 175.000 165.200 175.300 165.800 ;
        RECT 175.800 165.200 176.100 167.800 ;
        RECT 176.600 166.800 177.000 167.200 ;
        RECT 175.000 164.800 175.400 165.200 ;
        RECT 175.800 164.800 176.200 165.200 ;
        RECT 173.400 163.800 173.800 164.200 ;
        RECT 174.200 163.800 174.600 164.200 ;
        RECT 174.200 163.200 174.500 163.800 ;
        RECT 174.200 162.800 174.600 163.200 ;
        RECT 175.000 161.800 175.400 162.200 ;
        RECT 174.200 159.800 174.600 160.200 ;
        RECT 174.200 155.200 174.500 159.800 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 174.200 154.800 174.600 155.200 ;
        RECT 172.600 153.800 173.000 154.200 ;
        RECT 173.400 151.200 173.700 154.800 ;
        RECT 175.000 153.200 175.300 161.800 ;
        RECT 176.600 153.200 176.900 166.800 ;
        RECT 178.200 166.200 178.500 174.800 ;
        RECT 180.600 173.800 181.000 174.200 ;
        RECT 179.800 171.800 180.200 172.200 ;
        RECT 179.800 167.200 180.100 171.800 ;
        RECT 179.800 166.800 180.200 167.200 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 178.200 165.800 178.600 166.200 ;
        RECT 177.400 165.200 177.700 165.800 ;
        RECT 177.400 164.800 177.800 165.200 ;
        RECT 178.200 165.100 178.600 165.200 ;
        RECT 179.000 165.100 179.400 165.200 ;
        RECT 178.200 164.800 179.400 165.100 ;
        RECT 180.600 164.200 180.900 173.800 ;
        RECT 181.400 167.200 181.700 186.800 ;
        RECT 183.000 186.200 183.300 186.800 ;
        RECT 186.200 186.200 186.500 189.800 ;
        RECT 187.800 187.800 188.200 188.200 ;
        RECT 187.800 186.200 188.100 187.800 ;
        RECT 199.800 187.200 200.100 201.800 ;
        RECT 201.400 198.200 201.700 205.800 ;
        RECT 202.200 205.200 202.500 205.800 ;
        RECT 202.200 204.800 202.600 205.200 ;
        RECT 203.000 199.200 203.300 206.800 ;
        RECT 207.800 206.200 208.100 206.800 ;
        RECT 203.800 205.800 204.200 206.200 ;
        RECT 207.800 205.800 208.200 206.200 ;
        RECT 203.800 205.200 204.100 205.800 ;
        RECT 203.800 204.800 204.200 205.200 ;
        RECT 206.200 205.100 206.600 205.200 ;
        RECT 207.000 205.100 207.400 205.200 ;
        RECT 206.200 204.800 207.400 205.100 ;
        RECT 203.000 198.800 203.400 199.200 ;
        RECT 200.600 192.100 201.000 197.900 ;
        RECT 201.400 197.800 201.800 198.200 ;
        RECT 202.200 193.100 202.600 195.900 ;
        RECT 203.000 194.200 203.300 198.800 ;
        RECT 207.800 197.800 208.200 198.200 ;
        RECT 207.800 197.200 208.100 197.800 ;
        RECT 207.800 196.800 208.200 197.200 ;
        RECT 206.200 195.800 206.600 196.200 ;
        RECT 206.200 195.200 206.500 195.800 ;
        RECT 203.800 195.100 204.200 195.200 ;
        RECT 204.600 195.100 205.000 195.200 ;
        RECT 203.800 194.800 205.000 195.100 ;
        RECT 206.200 194.800 206.600 195.200 ;
        RECT 203.000 193.800 203.400 194.200 ;
        RECT 204.600 194.100 205.000 194.200 ;
        RECT 205.400 194.100 205.800 194.200 ;
        RECT 204.600 193.800 205.800 194.100 ;
        RECT 203.800 187.800 204.200 188.200 ;
        RECT 204.600 187.800 205.000 188.200 ;
        RECT 194.200 186.800 194.600 187.200 ;
        RECT 196.600 186.800 197.000 187.200 ;
        RECT 199.800 186.800 200.200 187.200 ;
        RECT 201.400 186.800 201.800 187.200 ;
        RECT 194.200 186.200 194.500 186.800 ;
        RECT 196.600 186.200 196.900 186.800 ;
        RECT 201.400 186.200 201.700 186.800 ;
        RECT 203.800 186.200 204.100 187.800 ;
        RECT 204.600 187.200 204.900 187.800 ;
        RECT 204.600 186.800 205.000 187.200 ;
        RECT 182.200 185.800 182.600 186.200 ;
        RECT 183.000 185.800 183.400 186.200 ;
        RECT 186.200 185.800 186.600 186.200 ;
        RECT 187.000 185.800 187.400 186.200 ;
        RECT 187.800 185.800 188.200 186.200 ;
        RECT 190.200 185.800 190.600 186.200 ;
        RECT 193.400 185.800 193.800 186.200 ;
        RECT 194.200 185.800 194.600 186.200 ;
        RECT 196.600 185.800 197.000 186.200 ;
        RECT 198.200 185.800 198.600 186.200 ;
        RECT 199.000 185.800 199.400 186.200 ;
        RECT 201.400 185.800 201.800 186.200 ;
        RECT 202.200 186.100 202.600 186.200 ;
        RECT 203.000 186.100 203.400 186.200 ;
        RECT 202.200 185.800 203.400 186.100 ;
        RECT 203.800 185.800 204.200 186.200 ;
        RECT 182.200 182.200 182.500 185.800 ;
        RECT 187.000 185.200 187.300 185.800 ;
        RECT 187.000 184.800 187.400 185.200 ;
        RECT 186.200 183.800 186.600 184.200 ;
        RECT 182.200 181.800 182.600 182.200 ;
        RECT 183.000 178.800 183.400 179.200 ;
        RECT 183.000 176.200 183.300 178.800 ;
        RECT 185.400 176.800 185.800 177.200 ;
        RECT 185.400 176.200 185.700 176.800 ;
        RECT 186.200 176.200 186.500 183.800 ;
        RECT 188.600 181.800 189.000 182.200 ;
        RECT 189.400 181.800 189.800 182.200 ;
        RECT 183.000 175.800 183.400 176.200 ;
        RECT 185.400 175.800 185.800 176.200 ;
        RECT 186.200 175.800 186.600 176.200 ;
        RECT 186.200 175.200 186.500 175.800 ;
        RECT 188.600 175.200 188.900 181.800 ;
        RECT 189.400 176.200 189.700 181.800 ;
        RECT 190.200 179.200 190.500 185.800 ;
        RECT 193.400 185.200 193.700 185.800 ;
        RECT 198.200 185.200 198.500 185.800 ;
        RECT 193.400 184.800 193.800 185.200 ;
        RECT 198.200 184.800 198.600 185.200 ;
        RECT 190.200 178.800 190.600 179.200 ;
        RECT 189.400 175.800 189.800 176.200 ;
        RECT 183.000 174.800 183.400 175.200 ;
        RECT 186.200 174.800 186.600 175.200 ;
        RECT 187.800 174.800 188.200 175.200 ;
        RECT 188.600 174.800 189.000 175.200 ;
        RECT 189.400 174.800 189.800 175.200 ;
        RECT 182.200 171.800 182.600 172.200 ;
        RECT 182.200 168.200 182.500 171.800 ;
        RECT 182.200 167.800 182.600 168.200 ;
        RECT 181.400 167.100 181.800 167.200 ;
        RECT 182.200 167.100 182.600 167.200 ;
        RECT 181.400 166.800 182.600 167.100 ;
        RECT 183.000 166.200 183.300 174.800 ;
        RECT 187.800 174.200 188.100 174.800 ;
        RECT 183.800 173.800 184.200 174.200 ;
        RECT 187.800 173.800 188.200 174.200 ;
        RECT 183.800 173.200 184.100 173.800 ;
        RECT 183.800 172.800 184.200 173.200 ;
        RECT 184.600 171.800 185.000 172.200 ;
        RECT 186.200 171.800 186.600 172.200 ;
        RECT 184.600 171.200 184.900 171.800 ;
        RECT 184.600 170.800 185.000 171.200 ;
        RECT 184.600 166.800 185.000 167.200 ;
        RECT 184.600 166.200 184.900 166.800 ;
        RECT 183.000 165.800 183.400 166.200 ;
        RECT 184.600 165.800 185.000 166.200 ;
        RECT 177.400 163.800 177.800 164.200 ;
        RECT 180.600 163.800 181.000 164.200 ;
        RECT 177.400 154.100 177.700 163.800 ;
        RECT 180.600 161.800 181.000 162.200 ;
        RECT 180.600 158.200 180.900 161.800 ;
        RECT 183.000 159.200 183.300 165.800 ;
        RECT 183.800 165.100 184.200 165.200 ;
        RECT 184.600 165.100 185.000 165.200 ;
        RECT 185.400 165.100 185.800 167.900 ;
        RECT 186.200 165.200 186.500 171.800 ;
        RECT 188.600 170.200 188.900 174.800 ;
        RECT 189.400 174.200 189.700 174.800 ;
        RECT 189.400 173.800 189.800 174.200 ;
        RECT 189.400 172.800 189.800 173.200 ;
        RECT 188.600 169.800 189.000 170.200 ;
        RECT 183.800 164.800 185.000 165.100 ;
        RECT 186.200 164.800 186.600 165.200 ;
        RECT 183.800 163.800 184.200 164.200 ;
        RECT 183.000 158.800 183.400 159.200 ;
        RECT 180.600 157.800 181.000 158.200 ;
        RECT 178.200 156.800 178.600 157.200 ;
        RECT 178.200 155.200 178.500 156.800 ;
        RECT 183.800 156.200 184.100 163.800 ;
        RECT 187.000 163.100 187.400 168.900 ;
        RECT 189.400 167.200 189.700 172.800 ;
        RECT 193.400 172.200 193.700 184.800 ;
        RECT 195.000 181.800 195.400 182.200 ;
        RECT 194.200 177.800 194.600 178.200 ;
        RECT 194.200 175.200 194.500 177.800 ;
        RECT 195.000 177.200 195.300 181.800 ;
        RECT 199.000 181.200 199.300 185.800 ;
        RECT 206.200 184.200 206.500 194.800 ;
        RECT 207.800 194.200 208.100 196.800 ;
        RECT 207.800 193.800 208.200 194.200 ;
        RECT 207.000 189.800 207.400 190.200 ;
        RECT 207.000 186.200 207.300 189.800 ;
        RECT 207.800 188.800 208.200 189.200 ;
        RECT 207.800 188.200 208.100 188.800 ;
        RECT 207.800 187.800 208.200 188.200 ;
        RECT 207.000 185.800 207.400 186.200 ;
        RECT 206.200 183.800 206.600 184.200 ;
        RECT 199.800 181.800 200.200 182.200 ;
        RECT 199.000 180.800 199.400 181.200 ;
        RECT 199.800 179.200 200.100 181.800 ;
        RECT 199.800 178.800 200.200 179.200 ;
        RECT 195.000 176.800 195.400 177.200 ;
        RECT 198.200 176.800 198.600 177.200 ;
        RECT 195.000 175.800 195.400 176.200 ;
        RECT 195.000 175.200 195.300 175.800 ;
        RECT 198.200 175.200 198.500 176.800 ;
        RECT 199.000 175.800 199.400 176.200 ;
        RECT 199.000 175.200 199.300 175.800 ;
        RECT 194.200 174.800 194.600 175.200 ;
        RECT 195.000 174.800 195.400 175.200 ;
        RECT 198.200 174.800 198.600 175.200 ;
        RECT 199.000 174.800 199.400 175.200 ;
        RECT 194.200 173.800 194.600 174.200 ;
        RECT 193.400 171.800 193.800 172.200 ;
        RECT 194.200 169.200 194.500 173.800 ;
        RECT 187.800 166.800 188.200 167.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 187.800 166.300 188.100 166.800 ;
        RECT 187.800 165.900 188.200 166.300 ;
        RECT 186.200 161.800 186.600 162.200 ;
        RECT 184.600 157.100 185.000 157.200 ;
        RECT 185.400 157.100 185.800 157.200 ;
        RECT 184.600 156.800 185.800 157.100 ;
        RECT 179.800 156.100 180.200 156.200 ;
        RECT 180.600 156.100 181.000 156.200 ;
        RECT 179.800 155.800 181.000 156.100 ;
        RECT 183.800 155.800 184.200 156.200 ;
        RECT 183.800 155.200 184.100 155.800 ;
        RECT 178.200 154.800 178.600 155.200 ;
        RECT 181.400 154.800 181.800 155.200 ;
        RECT 183.800 154.800 184.200 155.200 ;
        RECT 181.400 154.200 181.700 154.800 ;
        RECT 178.200 154.100 178.600 154.200 ;
        RECT 177.400 153.800 178.600 154.100 ;
        RECT 179.000 154.100 179.400 154.200 ;
        RECT 179.800 154.100 180.200 154.200 ;
        RECT 179.000 153.800 180.200 154.100 ;
        RECT 181.400 153.800 181.800 154.200 ;
        RECT 183.000 154.100 183.400 154.200 ;
        RECT 183.800 154.100 184.200 154.200 ;
        RECT 183.000 153.800 184.200 154.100 ;
        RECT 175.000 152.800 175.400 153.200 ;
        RECT 176.600 152.800 177.000 153.200 ;
        RECT 175.000 152.100 175.400 152.200 ;
        RECT 175.800 152.100 176.200 152.200 ;
        RECT 175.000 151.800 176.200 152.100 ;
        RECT 173.400 150.800 173.800 151.200 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 170.200 146.100 170.600 146.200 ;
        RECT 171.000 146.100 171.400 146.300 ;
        RECT 170.200 145.900 171.400 146.100 ;
        RECT 170.200 145.800 171.300 145.900 ;
        RECT 171.800 143.100 172.200 148.900 ;
        RECT 172.600 148.800 173.000 149.200 ;
        RECT 172.600 147.200 172.900 148.800 ;
        RECT 178.200 148.200 178.500 153.800 ;
        RECT 179.800 151.800 180.200 152.200 ;
        RECT 179.000 149.800 179.400 150.200 ;
        RECT 172.600 146.800 173.000 147.200 ;
        RECT 173.400 145.100 173.800 147.900 ;
        RECT 178.200 147.800 178.600 148.200 ;
        RECT 179.000 147.200 179.300 149.800 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 179.000 146.800 179.400 147.200 ;
        RECT 174.200 142.200 174.500 146.800 ;
        RECT 175.000 145.800 175.400 146.200 ;
        RECT 175.800 146.100 176.200 146.200 ;
        RECT 176.600 146.100 177.000 146.200 ;
        RECT 175.800 145.800 177.000 146.100 ;
        RECT 175.000 145.200 175.300 145.800 ;
        RECT 175.000 144.800 175.400 145.200 ;
        RECT 176.600 145.100 177.000 145.200 ;
        RECT 177.400 145.100 177.800 145.200 ;
        RECT 176.600 144.800 177.800 145.100 ;
        RECT 162.200 141.800 162.600 142.200 ;
        RECT 167.000 141.800 167.400 142.200 ;
        RECT 171.800 141.800 172.200 142.200 ;
        RECT 174.200 141.800 174.600 142.200 ;
        RECT 160.600 136.100 161.000 136.200 ;
        RECT 159.800 135.800 161.000 136.100 ;
        RECT 162.200 136.100 162.500 141.800 ;
        RECT 163.800 137.800 164.200 138.200 ;
        RECT 163.800 136.200 164.100 137.800 ;
        RECT 165.400 136.800 165.800 137.200 ;
        RECT 163.000 136.100 163.400 136.200 ;
        RECT 162.200 135.800 163.400 136.100 ;
        RECT 163.800 135.800 164.200 136.200 ;
        RECT 158.200 135.200 158.500 135.800 ;
        RECT 158.200 134.800 158.600 135.200 ;
        RECT 158.200 133.800 158.600 134.200 ;
        RECT 159.000 133.800 159.400 134.200 ;
        RECT 158.200 133.200 158.500 133.800 ;
        RECT 158.200 132.800 158.600 133.200 ;
        RECT 159.000 130.200 159.300 133.800 ;
        RECT 159.800 131.200 160.100 135.800 ;
        RECT 163.000 134.800 163.400 135.200 ;
        RECT 164.600 134.800 165.000 135.200 ;
        RECT 163.000 134.200 163.300 134.800 ;
        RECT 164.600 134.200 164.900 134.800 ;
        RECT 160.600 134.100 161.000 134.200 ;
        RECT 161.400 134.100 161.800 134.200 ;
        RECT 160.600 133.800 161.800 134.100 ;
        RECT 163.000 133.800 163.400 134.200 ;
        RECT 164.600 133.800 165.000 134.200 ;
        RECT 160.600 131.800 161.000 132.200 ;
        RECT 159.800 130.800 160.200 131.200 ;
        RECT 159.000 129.800 159.400 130.200 ;
        RECT 159.000 126.800 159.400 127.200 ;
        RECT 159.000 126.300 159.300 126.800 ;
        RECT 159.000 125.900 159.400 126.300 ;
        RECT 159.800 123.100 160.200 128.900 ;
        RECT 160.600 125.200 160.900 131.800 ;
        RECT 163.800 130.800 164.200 131.200 ;
        RECT 160.600 124.800 161.000 125.200 ;
        RECT 161.400 125.100 161.800 127.900 ;
        RECT 162.200 127.100 162.600 127.200 ;
        RECT 163.000 127.100 163.400 127.200 ;
        RECT 162.200 126.800 163.400 127.100 ;
        RECT 163.800 126.200 164.100 130.800 ;
        RECT 165.400 130.200 165.700 136.800 ;
        RECT 167.000 136.200 167.300 141.800 ;
        RECT 167.000 135.800 167.400 136.200 ;
        RECT 171.000 136.100 171.400 136.200 ;
        RECT 170.200 135.800 171.400 136.100 ;
        RECT 170.200 135.200 170.500 135.800 ;
        RECT 170.200 134.800 170.600 135.200 ;
        RECT 171.000 134.800 171.400 135.200 ;
        RECT 166.200 134.100 166.600 134.200 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 166.200 133.800 167.400 134.100 ;
        RECT 168.600 134.100 169.000 134.200 ;
        RECT 169.400 134.100 169.800 134.200 ;
        RECT 168.600 133.800 169.800 134.100 ;
        RECT 170.200 133.800 170.600 134.200 ;
        RECT 170.200 133.200 170.500 133.800 ;
        RECT 170.200 132.800 170.600 133.200 ;
        RECT 171.000 132.200 171.300 134.800 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 171.000 131.800 171.400 132.200 ;
        RECT 167.000 131.200 167.300 131.800 ;
        RECT 167.000 130.800 167.400 131.200 ;
        RECT 165.400 129.800 165.800 130.200 ;
        RECT 169.400 129.800 169.800 130.200 ;
        RECT 169.400 129.200 169.700 129.800 ;
        RECT 171.800 129.200 172.100 141.800 ;
        RECT 172.600 136.800 173.000 137.200 ;
        RECT 172.600 136.200 172.900 136.800 ;
        RECT 172.600 135.800 173.000 136.200 ;
        RECT 173.400 135.100 173.800 135.200 ;
        RECT 174.200 135.100 174.600 135.200 ;
        RECT 173.400 134.800 174.600 135.100 ;
        RECT 173.400 133.800 173.800 134.200 ;
        RECT 173.400 133.200 173.700 133.800 ;
        RECT 173.400 132.800 173.800 133.200 ;
        RECT 174.200 132.800 174.600 133.200 ;
        RECT 169.400 128.800 169.800 129.200 ;
        RECT 171.800 128.800 172.200 129.200 ;
        RECT 174.200 127.200 174.500 132.800 ;
        RECT 164.600 127.100 165.000 127.200 ;
        RECT 165.400 127.100 165.800 127.200 ;
        RECT 164.600 126.800 165.800 127.100 ;
        RECT 168.600 126.800 169.000 127.200 ;
        RECT 174.200 126.800 174.600 127.200 ;
        RECT 168.600 126.200 168.900 126.800 ;
        RECT 175.000 126.200 175.300 144.800 ;
        RECT 179.000 143.800 179.400 144.200 ;
        RECT 176.600 135.800 177.000 136.200 ;
        RECT 178.200 135.800 178.600 136.200 ;
        RECT 176.600 135.200 176.900 135.800 ;
        RECT 176.600 134.800 177.000 135.200 ;
        RECT 178.200 134.200 178.500 135.800 ;
        RECT 179.000 134.200 179.300 143.800 ;
        RECT 179.800 137.200 180.100 151.800 ;
        RECT 179.800 136.800 180.200 137.200 ;
        RECT 180.600 135.800 181.000 136.200 ;
        RECT 180.600 135.200 180.900 135.800 ;
        RECT 180.600 134.800 181.000 135.200 ;
        RECT 175.800 134.100 176.200 134.200 ;
        RECT 176.600 134.100 177.000 134.200 ;
        RECT 175.800 133.800 177.000 134.100 ;
        RECT 178.200 133.800 178.600 134.200 ;
        RECT 179.000 133.800 179.400 134.200 ;
        RECT 179.800 128.800 180.200 129.200 ;
        RECT 179.000 128.100 179.400 128.200 ;
        RECT 179.800 128.100 180.100 128.800 ;
        RECT 179.000 127.800 180.100 128.100 ;
        RECT 179.000 127.200 179.300 127.800 ;
        RECT 176.600 127.100 177.000 127.200 ;
        RECT 177.400 127.100 177.800 127.200 ;
        RECT 176.600 126.800 177.800 127.100 ;
        RECT 179.000 126.800 179.400 127.200 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 167.000 125.800 167.400 126.200 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 174.200 125.800 174.600 126.200 ;
        RECT 175.000 125.800 175.400 126.200 ;
        RECT 162.200 125.200 162.500 125.800 ;
        RECT 162.200 124.800 162.600 125.200 ;
        RECT 167.000 124.200 167.300 125.800 ;
        RECT 167.800 125.100 168.200 125.200 ;
        RECT 168.600 125.100 169.000 125.200 ;
        RECT 167.800 124.800 169.000 125.100 ;
        RECT 170.200 125.100 170.600 125.200 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 170.200 124.800 171.400 125.100 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 166.200 124.100 166.600 124.200 ;
        RECT 165.400 123.800 166.600 124.100 ;
        RECT 167.000 123.800 167.400 124.200 ;
        RECT 165.400 121.800 165.800 122.200 ;
        RECT 162.200 119.800 162.600 120.200 ;
        RECT 162.200 119.200 162.500 119.800 ;
        RECT 162.200 118.800 162.600 119.200 ;
        RECT 164.600 118.800 165.000 119.200 ;
        RECT 159.800 116.100 160.200 116.200 ;
        RECT 160.600 116.100 161.000 116.200 ;
        RECT 159.800 115.800 161.000 116.100 ;
        RECT 163.000 116.100 163.400 116.200 ;
        RECT 163.800 116.100 164.200 116.200 ;
        RECT 163.000 115.800 164.200 116.100 ;
        RECT 157.400 114.800 157.800 115.200 ;
        RECT 159.000 114.800 159.400 115.200 ;
        RECT 163.800 114.800 164.200 115.200 ;
        RECT 155.000 113.800 155.400 114.200 ;
        RECT 155.800 114.100 156.200 114.200 ;
        RECT 156.600 114.100 157.000 114.200 ;
        RECT 155.800 113.800 157.000 114.100 ;
        RECT 157.400 113.200 157.700 114.800 ;
        RECT 159.000 114.200 159.300 114.800 ;
        RECT 163.800 114.200 164.100 114.800 ;
        RECT 164.600 114.200 164.900 118.800 ;
        RECT 165.400 115.200 165.700 121.800 ;
        RECT 166.200 116.100 166.600 116.200 ;
        RECT 167.000 116.100 167.400 116.200 ;
        RECT 173.400 116.100 173.800 116.200 ;
        RECT 166.200 115.800 167.400 116.100 ;
        RECT 172.600 115.800 173.800 116.100 ;
        RECT 165.400 114.800 165.800 115.200 ;
        RECT 167.000 114.800 167.400 115.200 ;
        RECT 167.000 114.200 167.300 114.800 ;
        RECT 158.200 113.800 158.600 114.200 ;
        RECT 159.000 113.800 159.400 114.200 ;
        RECT 163.800 113.800 164.200 114.200 ;
        RECT 164.600 113.800 165.000 114.200 ;
        RECT 167.000 113.800 167.400 114.200 ;
        RECT 167.800 113.800 168.200 114.200 ;
        RECT 147.800 112.800 148.200 113.200 ;
        RECT 157.400 112.800 157.800 113.200 ;
        RECT 148.600 111.800 149.000 112.200 ;
        RECT 151.800 111.800 152.200 112.200 ;
        RECT 154.200 111.800 154.600 112.200 ;
        RECT 155.000 111.800 155.400 112.200 ;
        RECT 147.000 109.800 147.400 110.200 ;
        RECT 141.400 108.800 141.800 109.200 ;
        RECT 148.600 108.200 148.900 111.800 ;
        RECT 151.800 111.200 152.100 111.800 ;
        RECT 154.200 111.200 154.500 111.800 ;
        RECT 149.400 110.800 149.800 111.200 ;
        RECT 151.800 110.800 152.200 111.200 ;
        RECT 154.200 110.800 154.600 111.200 ;
        RECT 139.000 107.800 139.400 108.200 ;
        RECT 148.600 107.800 149.000 108.200 ;
        RECT 139.000 107.200 139.300 107.800 ;
        RECT 148.600 107.200 148.900 107.800 ;
        RECT 149.400 107.200 149.700 110.800 ;
        RECT 150.200 109.800 150.600 110.200 ;
        RECT 137.400 106.800 137.800 107.200 ;
        RECT 139.000 106.800 139.400 107.200 ;
        RECT 143.800 106.800 144.200 107.200 ;
        RECT 148.600 106.800 149.000 107.200 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 137.400 106.100 137.800 106.200 ;
        RECT 136.600 105.800 137.800 106.100 ;
        RECT 137.400 105.200 137.700 105.800 ;
        RECT 137.400 104.800 137.800 105.200 ;
        RECT 141.400 105.100 141.800 105.200 ;
        RECT 142.200 105.100 142.600 105.200 ;
        RECT 141.400 104.800 142.600 105.100 ;
        RECT 136.600 104.100 137.000 104.200 ;
        RECT 137.400 104.100 137.800 104.200 ;
        RECT 136.600 103.800 137.800 104.100 ;
        RECT 135.800 102.800 136.200 103.200 ;
        RECT 135.800 95.200 136.100 102.800 ;
        RECT 135.800 94.800 136.200 95.200 ;
        RECT 135.800 93.800 136.200 94.200 ;
        RECT 135.800 92.200 136.100 93.800 ;
        RECT 138.200 93.100 138.600 95.900 ;
        RECT 135.800 91.800 136.200 92.200 ;
        RECT 139.800 92.100 140.200 97.900 ;
        RECT 142.200 96.200 142.500 104.800 ;
        RECT 143.800 104.200 144.100 106.800 ;
        RECT 145.400 106.100 145.800 106.200 ;
        RECT 146.200 106.100 146.600 106.200 ;
        RECT 145.400 105.800 146.600 106.100 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 147.800 106.100 148.200 106.200 ;
        RECT 147.000 105.800 148.200 106.100 ;
        RECT 148.600 105.800 149.000 106.200 ;
        RECT 145.400 105.100 145.800 105.200 ;
        RECT 146.200 105.100 146.600 105.200 ;
        RECT 145.400 104.800 146.600 105.100 ;
        RECT 147.800 105.100 148.200 105.200 ;
        RECT 148.600 105.100 148.900 105.800 ;
        RECT 147.800 104.800 148.900 105.100 ;
        RECT 143.800 103.800 144.200 104.200 ;
        RECT 149.400 100.800 149.800 101.200 ;
        RECT 143.800 97.800 144.200 98.200 ;
        RECT 142.200 95.800 142.600 96.200 ;
        RECT 143.800 95.200 144.100 97.800 ;
        RECT 142.200 95.100 142.600 95.200 ;
        RECT 143.000 95.100 143.400 95.200 ;
        RECT 142.200 94.800 143.400 95.100 ;
        RECT 143.800 94.800 144.200 95.200 ;
        RECT 144.600 92.100 145.000 97.900 ;
        RECT 147.800 96.100 148.200 96.200 ;
        RECT 147.800 95.800 148.900 96.100 ;
        RECT 147.000 95.100 147.400 95.200 ;
        RECT 147.800 95.100 148.200 95.200 ;
        RECT 147.000 94.800 148.200 95.100 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 147.000 89.200 147.300 91.800 ;
        RECT 147.800 89.800 148.200 90.200 ;
        RECT 137.400 86.800 137.800 87.200 ;
        RECT 137.400 86.300 137.700 86.800 ;
        RECT 137.400 85.900 137.800 86.300 ;
        RECT 138.200 83.100 138.600 88.900 ;
        RECT 140.600 88.800 141.000 89.200 ;
        RECT 147.000 88.800 147.400 89.200 ;
        RECT 139.800 85.100 140.200 87.900 ;
        RECT 140.600 87.200 140.900 88.800 ;
        RECT 147.000 87.800 147.400 88.200 ;
        RECT 147.000 87.200 147.300 87.800 ;
        RECT 140.600 86.800 141.000 87.200 ;
        RECT 143.800 87.100 144.200 87.200 ;
        RECT 144.600 87.100 145.000 87.200 ;
        RECT 143.800 86.800 145.000 87.100 ;
        RECT 147.000 86.800 147.400 87.200 ;
        RECT 143.800 85.800 144.200 86.200 ;
        RECT 145.400 86.100 145.800 86.200 ;
        RECT 146.200 86.100 146.600 86.200 ;
        RECT 145.400 85.800 146.600 86.100 ;
        RECT 143.800 85.200 144.100 85.800 ;
        RECT 147.800 85.200 148.100 89.800 ;
        RECT 148.600 89.200 148.900 95.800 ;
        RECT 149.400 95.200 149.700 100.800 ;
        RECT 149.400 94.800 149.800 95.200 ;
        RECT 149.400 90.200 149.700 94.800 ;
        RECT 150.200 94.200 150.500 109.800 ;
        RECT 151.800 108.800 152.200 109.200 ;
        RECT 151.800 105.200 152.100 108.800 ;
        RECT 155.000 108.200 155.300 111.800 ;
        RECT 158.200 109.200 158.500 113.800 ;
        RECT 160.600 111.800 161.000 112.200 ;
        RECT 158.200 108.800 158.600 109.200 ;
        RECT 155.000 107.800 155.400 108.200 ;
        RECT 156.600 107.800 157.000 108.200 ;
        RECT 156.600 107.200 156.900 107.800 ;
        RECT 160.600 107.200 160.900 111.800 ;
        RECT 162.200 108.100 162.600 108.200 ;
        RECT 163.000 108.100 163.400 108.200 ;
        RECT 162.200 107.800 163.400 108.100 ;
        RECT 163.800 107.200 164.100 113.800 ;
        RECT 167.800 112.200 168.100 113.800 ;
        RECT 167.800 111.800 168.200 112.200 ;
        RECT 168.600 111.800 169.000 112.200 ;
        RECT 171.000 111.800 171.400 112.200 ;
        RECT 167.000 109.100 167.400 109.200 ;
        RECT 167.800 109.100 168.200 109.200 ;
        RECT 167.000 108.800 168.200 109.100 ;
        RECT 167.800 107.800 168.200 108.200 ;
        RECT 167.800 107.200 168.100 107.800 ;
        RECT 156.600 106.800 157.000 107.200 ;
        RECT 159.000 107.100 159.400 107.200 ;
        RECT 159.800 107.100 160.200 107.200 ;
        RECT 159.000 106.800 160.200 107.100 ;
        RECT 160.600 106.800 161.000 107.200 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 166.200 107.100 166.600 107.200 ;
        RECT 167.000 107.100 167.400 107.200 ;
        RECT 166.200 106.800 167.400 107.100 ;
        RECT 167.800 106.800 168.200 107.200 ;
        RECT 155.000 105.800 155.400 106.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 159.000 106.100 159.400 106.200 ;
        RECT 158.200 105.800 159.400 106.100 ;
        RECT 159.800 105.800 160.200 106.200 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 163.800 106.100 164.200 106.200 ;
        RECT 163.000 105.800 164.200 106.100 ;
        RECT 164.600 106.100 165.000 106.200 ;
        RECT 165.400 106.100 165.800 106.200 ;
        RECT 164.600 105.800 165.800 106.100 ;
        RECT 151.800 104.800 152.200 105.200 ;
        RECT 152.600 104.800 153.000 105.200 ;
        RECT 153.400 105.100 153.800 105.200 ;
        RECT 154.200 105.100 154.600 105.200 ;
        RECT 153.400 104.800 154.600 105.100 ;
        RECT 151.800 103.200 152.100 104.800 ;
        RECT 151.800 102.800 152.200 103.200 ;
        RECT 152.600 99.200 152.900 104.800 ;
        RECT 151.000 98.800 151.400 99.200 ;
        RECT 152.600 98.800 153.000 99.200 ;
        RECT 151.000 96.200 151.300 98.800 ;
        RECT 155.000 97.200 155.300 105.800 ;
        RECT 155.000 96.800 155.400 97.200 ;
        RECT 156.600 96.200 156.900 105.800 ;
        RECT 157.400 104.800 157.800 105.200 ;
        RECT 159.000 105.100 159.400 105.200 ;
        RECT 159.800 105.100 160.100 105.800 ;
        RECT 159.000 104.800 160.100 105.100 ;
        RECT 163.800 104.800 164.200 105.200 ;
        RECT 157.400 104.200 157.700 104.800 ;
        RECT 157.400 103.800 157.800 104.200 ;
        RECT 159.000 103.800 159.400 104.200 ;
        RECT 159.000 99.200 159.300 103.800 ;
        RECT 159.000 98.800 159.400 99.200 ;
        RECT 151.000 95.800 151.400 96.200 ;
        RECT 156.600 95.800 157.000 96.200 ;
        RECT 156.600 95.200 156.900 95.800 ;
        RECT 151.800 95.100 152.200 95.200 ;
        RECT 152.600 95.100 153.000 95.200 ;
        RECT 151.800 94.800 153.000 95.100 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 150.200 93.800 150.600 94.200 ;
        RECT 154.200 93.800 154.600 94.200 ;
        RECT 151.800 90.800 152.200 91.200 ;
        RECT 149.400 89.800 149.800 90.200 ;
        RECT 148.600 88.800 149.000 89.200 ;
        RECT 149.400 88.800 149.800 89.200 ;
        RECT 149.400 87.200 149.700 88.800 ;
        RECT 151.800 87.200 152.100 90.800 ;
        RECT 153.400 88.800 153.800 89.200 ;
        RECT 153.400 87.200 153.700 88.800 ;
        RECT 149.400 86.800 149.800 87.200 ;
        RECT 151.800 86.800 152.200 87.200 ;
        RECT 152.600 86.800 153.000 87.200 ;
        RECT 153.400 86.800 153.800 87.200 ;
        RECT 149.400 85.200 149.700 86.800 ;
        RECT 143.800 84.800 144.200 85.200 ;
        RECT 147.800 84.800 148.200 85.200 ;
        RECT 149.400 84.800 149.800 85.200 ;
        RECT 144.600 78.800 145.000 79.200 ;
        RECT 143.000 77.800 143.400 78.200 ;
        RECT 136.600 75.800 137.000 76.200 ;
        RECT 138.200 75.800 138.600 76.200 ;
        RECT 136.600 75.200 136.900 75.800 ;
        RECT 138.200 75.200 138.500 75.800 ;
        RECT 143.000 75.200 143.300 77.800 ;
        RECT 143.800 75.800 144.200 76.200 ;
        RECT 143.800 75.200 144.100 75.800 ;
        RECT 135.000 74.800 135.400 75.200 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 138.200 74.800 138.600 75.200 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 143.800 74.800 144.200 75.200 ;
        RECT 134.200 74.100 134.600 74.200 ;
        RECT 135.000 74.100 135.400 74.200 ;
        RECT 134.200 73.800 135.400 74.100 ;
        RECT 139.800 73.800 140.200 74.200 ;
        RECT 141.400 74.100 141.800 74.200 ;
        RECT 142.200 74.100 142.600 74.200 ;
        RECT 141.400 73.800 142.600 74.100 ;
        RECT 139.800 72.200 140.100 73.800 ;
        RECT 134.200 72.100 134.600 72.200 ;
        RECT 135.000 72.100 135.400 72.200 ;
        RECT 134.200 71.800 135.400 72.100 ;
        RECT 139.800 71.800 140.200 72.200 ;
        RECT 143.000 70.800 143.400 71.200 ;
        RECT 131.000 63.800 131.400 64.200 ;
        RECT 122.200 62.800 122.600 63.200 ;
        RECT 126.200 62.800 126.600 63.200 ;
        RECT 131.800 63.100 132.200 68.900 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 133.400 66.100 133.800 66.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 133.400 65.800 134.600 66.100 ;
        RECT 132.600 63.100 132.900 65.800 ;
        RECT 136.600 63.100 137.000 68.900 ;
        RECT 143.000 68.200 143.300 70.800 ;
        RECT 142.200 68.100 142.600 68.200 ;
        RECT 143.000 68.100 143.400 68.200 ;
        RECT 138.200 65.100 138.600 67.900 ;
        RECT 142.200 67.800 143.400 68.100 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 139.000 64.100 139.300 66.800 ;
        RECT 144.600 66.200 144.900 78.800 ;
        RECT 145.400 77.800 145.800 78.200 ;
        RECT 145.400 76.200 145.700 77.800 ;
        RECT 147.800 77.200 148.100 84.800 ;
        RECT 151.000 81.800 151.400 82.200 ;
        RECT 147.800 76.800 148.200 77.200 ;
        RECT 145.400 75.800 145.800 76.200 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 147.000 73.200 147.300 73.800 ;
        RECT 147.000 72.800 147.400 73.200 ;
        RECT 147.800 73.100 148.200 75.900 ;
        RECT 148.600 75.800 149.000 76.200 ;
        RECT 148.600 74.200 148.900 75.800 ;
        RECT 148.600 73.800 149.000 74.200 ;
        RECT 149.400 72.100 149.800 77.900 ;
        RECT 151.000 76.200 151.300 81.800 ;
        RECT 151.000 75.800 151.400 76.200 ;
        RECT 151.800 75.200 152.100 86.800 ;
        RECT 152.600 86.200 152.900 86.800 ;
        RECT 152.600 85.800 153.000 86.200 ;
        RECT 154.200 86.100 154.500 93.800 ;
        RECT 160.600 93.100 161.000 95.900 ;
        RECT 155.000 91.800 155.400 92.200 ;
        RECT 160.600 91.800 161.000 92.200 ;
        RECT 162.200 92.100 162.600 97.900 ;
        RECT 163.000 94.700 163.400 95.100 ;
        RECT 163.000 92.200 163.300 94.700 ;
        RECT 163.000 91.800 163.400 92.200 ;
        RECT 155.000 89.100 155.300 91.800 ;
        RECT 160.600 89.200 160.900 91.800 ;
        RECT 163.000 90.800 163.400 91.200 ;
        RECT 155.000 88.800 156.100 89.100 ;
        RECT 160.600 88.800 161.000 89.200 ;
        RECT 161.400 88.800 161.800 89.200 ;
        RECT 153.400 85.800 154.500 86.100 ;
        RECT 155.800 87.200 156.100 88.800 ;
        RECT 161.400 88.200 161.700 88.800 ;
        RECT 161.400 87.800 161.800 88.200 ;
        RECT 163.000 87.200 163.300 90.800 ;
        RECT 155.800 86.800 156.200 87.200 ;
        RECT 156.600 87.100 157.000 87.200 ;
        RECT 157.400 87.100 157.800 87.200 ;
        RECT 156.600 86.800 157.800 87.100 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 163.000 86.800 163.400 87.200 ;
        RECT 155.800 86.200 156.100 86.800 ;
        RECT 155.800 85.800 156.200 86.200 ;
        RECT 162.200 85.800 162.600 86.200 ;
        RECT 153.400 85.200 153.700 85.800 ;
        RECT 153.400 84.800 153.800 85.200 ;
        RECT 154.200 85.100 154.600 85.200 ;
        RECT 155.000 85.100 155.400 85.200 ;
        RECT 154.200 84.800 155.400 85.100 ;
        RECT 151.000 75.100 151.400 75.200 ;
        RECT 150.200 74.800 151.400 75.100 ;
        RECT 151.800 74.800 152.200 75.200 ;
        RECT 150.200 74.700 150.600 74.800 ;
        RECT 151.000 71.800 151.400 72.200 ;
        RECT 149.400 69.100 149.800 69.200 ;
        RECT 150.200 69.100 150.600 69.200 ;
        RECT 149.400 68.800 150.600 69.100 ;
        RECT 147.000 66.800 147.400 67.200 ;
        RECT 140.600 66.100 141.000 66.200 ;
        RECT 141.400 66.100 141.800 66.200 ;
        RECT 140.600 65.800 141.800 66.100 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 146.200 65.800 146.600 66.200 ;
        RECT 146.200 65.200 146.500 65.800 ;
        RECT 138.200 63.800 139.300 64.100 ;
        RECT 141.400 64.800 141.800 65.200 ;
        RECT 143.800 65.100 144.200 65.200 ;
        RECT 143.000 64.800 144.200 65.100 ;
        RECT 146.200 64.800 146.600 65.200 ;
        RECT 132.600 62.800 133.700 63.100 ;
        RECT 122.200 59.200 122.500 62.800 ;
        RECT 122.200 58.800 122.600 59.200 ;
        RECT 131.800 59.100 132.200 59.200 ;
        RECT 132.600 59.100 133.000 59.200 ;
        RECT 131.800 58.800 133.000 59.100 ;
        RECT 120.600 57.800 121.000 58.200 ;
        RECT 121.400 57.800 121.800 58.200 ;
        RECT 120.600 56.200 120.900 57.800 ;
        RECT 121.400 57.200 121.700 57.800 ;
        RECT 121.400 56.800 121.800 57.200 ;
        RECT 123.800 56.800 124.200 57.200 ;
        RECT 129.400 56.800 129.800 57.200 ;
        RECT 131.000 57.100 131.400 57.200 ;
        RECT 131.800 57.100 132.200 57.200 ;
        RECT 131.000 56.800 132.200 57.100 ;
        RECT 132.600 56.800 133.000 57.200 ;
        RECT 123.800 56.200 124.100 56.800 ;
        RECT 129.400 56.200 129.700 56.800 ;
        RECT 132.600 56.200 132.900 56.800 ;
        RECT 120.600 55.800 121.000 56.200 ;
        RECT 123.000 55.800 123.400 56.200 ;
        RECT 123.800 55.800 124.200 56.200 ;
        RECT 124.600 55.800 125.000 56.200 ;
        RECT 125.400 56.100 125.800 56.200 ;
        RECT 125.400 55.800 127.300 56.100 ;
        RECT 129.400 55.800 129.800 56.200 ;
        RECT 132.600 55.800 133.000 56.200 ;
        RECT 119.800 54.800 120.200 55.200 ;
        RECT 122.200 54.800 122.600 55.200 ;
        RECT 123.000 55.100 123.300 55.800 ;
        RECT 123.000 54.800 124.100 55.100 ;
        RECT 119.000 50.800 119.400 51.200 ;
        RECT 119.800 47.200 120.100 54.800 ;
        RECT 122.200 49.200 122.500 54.800 ;
        RECT 123.000 51.800 123.400 52.200 ;
        RECT 122.200 48.800 122.600 49.200 ;
        RECT 123.000 47.200 123.300 51.800 ;
        RECT 123.800 49.200 124.100 54.800 ;
        RECT 123.800 48.800 124.200 49.200 ;
        RECT 119.800 46.800 120.200 47.200 ;
        RECT 123.000 46.800 123.400 47.200 ;
        RECT 120.600 45.800 121.000 46.200 ;
        RECT 120.600 44.200 120.900 45.800 ;
        RECT 121.400 44.800 121.800 45.200 ;
        RECT 123.000 44.800 123.400 45.200 ;
        RECT 120.600 43.800 121.000 44.200 ;
        RECT 121.400 43.200 121.700 44.800 ;
        RECT 121.400 42.800 121.800 43.200 ;
        RECT 123.000 39.200 123.300 44.800 ;
        RECT 109.400 38.800 109.800 39.200 ;
        RECT 116.600 38.800 117.000 39.200 ;
        RECT 118.200 38.800 118.600 39.200 ;
        RECT 123.000 38.800 123.400 39.200 ;
        RECT 110.200 37.800 110.600 38.200 ;
        RECT 107.000 35.800 107.400 36.200 ;
        RECT 107.000 35.200 107.300 35.800 ;
        RECT 110.200 35.200 110.500 37.800 ;
        RECT 113.400 36.800 113.800 37.200 ;
        RECT 113.400 36.200 113.700 36.800 ;
        RECT 116.600 36.200 116.900 38.800 ;
        RECT 124.600 37.200 124.900 55.800 ;
        RECT 126.200 54.800 126.600 55.200 ;
        RECT 126.200 54.200 126.500 54.800 ;
        RECT 127.000 54.200 127.300 55.800 ;
        RECT 130.200 54.800 130.600 55.200 ;
        RECT 130.200 54.200 130.500 54.800 ;
        RECT 125.400 53.800 125.800 54.200 ;
        RECT 126.200 53.800 126.600 54.200 ;
        RECT 127.000 53.800 127.400 54.200 ;
        RECT 130.200 53.800 130.600 54.200 ;
        RECT 132.600 53.800 133.000 54.200 ;
        RECT 125.400 53.200 125.700 53.800 ;
        RECT 125.400 52.800 125.800 53.200 ;
        RECT 132.600 52.200 132.900 53.800 ;
        RECT 127.800 51.800 128.200 52.200 ;
        RECT 132.600 51.800 133.000 52.200 ;
        RECT 127.800 50.200 128.100 51.800 ;
        RECT 133.400 51.100 133.700 62.800 ;
        RECT 138.200 61.200 138.500 63.800 ;
        RECT 138.200 60.800 138.600 61.200 ;
        RECT 141.400 59.200 141.700 64.800 ;
        RECT 143.000 59.200 143.300 64.800 ;
        RECT 144.600 63.800 145.000 64.200 ;
        RECT 141.400 58.800 141.800 59.200 ;
        RECT 143.000 58.800 143.400 59.200 ;
        RECT 142.200 57.800 142.600 58.200 ;
        RECT 135.800 56.800 136.200 57.200 ;
        RECT 134.200 55.800 134.600 56.200 ;
        RECT 135.000 55.800 135.400 56.200 ;
        RECT 134.200 54.200 134.500 55.800 ;
        RECT 135.000 55.200 135.300 55.800 ;
        RECT 135.800 55.200 136.100 56.800 ;
        RECT 135.000 54.800 135.400 55.200 ;
        RECT 135.800 54.800 136.200 55.200 ;
        RECT 138.200 54.800 138.600 55.200 ;
        RECT 138.200 54.200 138.500 54.800 ;
        RECT 134.200 53.800 134.600 54.200 ;
        RECT 136.600 53.800 137.000 54.200 ;
        RECT 138.200 53.800 138.600 54.200 ;
        RECT 136.600 53.200 136.900 53.800 ;
        RECT 142.200 53.200 142.500 57.800 ;
        RECT 143.800 55.800 144.200 56.200 ;
        RECT 136.600 52.800 137.000 53.200 ;
        RECT 142.200 52.800 142.600 53.200 ;
        RECT 143.000 52.800 143.400 53.200 ;
        RECT 133.400 50.800 134.500 51.100 ;
        RECT 127.800 49.800 128.200 50.200 ;
        RECT 125.400 47.800 125.800 48.200 ;
        RECT 125.400 47.200 125.700 47.800 ;
        RECT 125.400 46.800 125.800 47.200 ;
        RECT 125.400 44.100 125.800 44.200 ;
        RECT 126.200 44.100 126.600 44.200 ;
        RECT 125.400 43.800 126.600 44.100 ;
        RECT 128.600 43.100 129.000 48.900 ;
        RECT 131.800 48.800 132.200 49.200 ;
        RECT 131.800 46.200 132.100 48.800 ;
        RECT 131.800 45.800 132.200 46.200 ;
        RECT 132.600 44.800 133.000 45.200 ;
        RECT 132.600 39.200 132.900 44.800 ;
        RECT 133.400 43.100 133.800 48.900 ;
        RECT 134.200 47.200 134.500 50.800 ;
        RECT 140.600 49.800 141.000 50.200 ;
        RECT 137.400 49.100 137.800 49.200 ;
        RECT 138.200 49.100 138.600 49.200 ;
        RECT 137.400 48.800 138.600 49.100 ;
        RECT 134.200 46.800 134.600 47.200 ;
        RECT 132.600 38.800 133.000 39.200 ;
        RECT 124.600 36.800 125.000 37.200 ;
        RECT 130.200 36.800 130.600 37.200 ;
        RECT 113.400 35.800 113.800 36.200 ;
        RECT 116.600 35.800 117.000 36.200 ;
        RECT 118.200 35.800 118.600 36.200 ;
        RECT 119.800 36.100 120.200 36.200 ;
        RECT 119.800 35.800 120.900 36.100 ;
        RECT 113.400 35.200 113.700 35.800 ;
        RECT 118.200 35.200 118.500 35.800 ;
        RECT 107.000 34.800 107.400 35.200 ;
        RECT 107.800 35.100 108.200 35.200 ;
        RECT 108.600 35.100 109.000 35.200 ;
        RECT 107.800 34.800 109.000 35.100 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 111.000 34.800 111.400 35.200 ;
        RECT 113.400 34.800 113.800 35.200 ;
        RECT 115.000 35.100 115.400 35.200 ;
        RECT 115.800 35.100 116.200 35.200 ;
        RECT 115.000 34.800 116.200 35.100 ;
        RECT 118.200 34.800 118.600 35.200 ;
        RECT 119.800 34.800 120.200 35.200 ;
        RECT 111.000 34.200 111.300 34.800 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 111.000 33.800 111.400 34.200 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 116.600 34.100 117.000 34.200 ;
        RECT 115.800 33.800 117.000 34.100 ;
        RECT 117.400 33.800 117.800 34.200 ;
        RECT 103.800 27.800 104.900 28.100 ;
        RECT 105.400 31.800 105.800 32.200 ;
        RECT 95.800 27.200 96.100 27.800 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 97.400 26.800 97.800 27.200 ;
        RECT 102.200 26.800 102.600 27.200 ;
        RECT 103.000 26.800 103.400 27.200 ;
        RECT 97.400 25.200 97.700 26.800 ;
        RECT 97.400 24.800 97.800 25.200 ;
        RECT 99.800 24.800 100.200 25.200 ;
        RECT 97.400 21.200 97.700 24.800 ;
        RECT 99.800 22.200 100.100 24.800 ;
        RECT 99.800 21.800 100.200 22.200 ;
        RECT 97.400 20.800 97.800 21.200 ;
        RECT 99.800 20.800 100.200 21.200 ;
        RECT 99.800 19.200 100.100 20.800 ;
        RECT 102.200 19.200 102.500 26.800 ;
        RECT 99.800 18.800 100.200 19.200 ;
        RECT 102.200 18.800 102.600 19.200 ;
        RECT 92.600 15.800 93.000 16.200 ;
        RECT 92.600 15.200 92.900 15.800 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 91.800 13.800 92.200 14.200 ;
        RECT 94.200 11.800 94.600 12.200 ;
        RECT 95.800 12.100 96.200 17.900 ;
        RECT 98.200 16.800 98.600 17.200 ;
        RECT 98.200 13.200 98.500 16.800 ;
        RECT 98.200 13.100 98.600 13.200 ;
        RECT 99.000 13.100 99.400 13.200 ;
        RECT 100.600 13.100 101.000 15.900 ;
        RECT 98.200 12.800 99.400 13.100 ;
        RECT 102.200 12.100 102.600 17.900 ;
        RECT 94.200 9.200 94.500 11.800 ;
        RECT 103.000 10.200 103.300 26.800 ;
        RECT 103.800 26.200 104.100 27.800 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 104.600 26.200 104.900 26.800 ;
        RECT 103.800 25.800 104.200 26.200 ;
        RECT 104.600 25.800 105.000 26.200 ;
        RECT 103.800 17.200 104.100 25.800 ;
        RECT 105.400 25.200 105.700 31.800 ;
        RECT 106.200 29.200 106.500 33.800 ;
        RECT 111.000 32.200 111.300 33.800 ;
        RECT 107.000 31.800 107.400 32.200 ;
        RECT 111.000 31.800 111.400 32.200 ;
        RECT 114.200 31.800 114.600 32.200 ;
        RECT 115.800 31.800 116.200 32.200 ;
        RECT 106.200 28.800 106.600 29.200 ;
        RECT 105.400 24.800 105.800 25.200 ;
        RECT 106.200 25.100 106.600 27.900 ;
        RECT 107.000 27.200 107.300 31.800 ;
        RECT 114.200 30.200 114.500 31.800 ;
        RECT 114.200 29.800 114.600 30.200 ;
        RECT 115.800 29.200 116.100 31.800 ;
        RECT 114.200 29.100 114.600 29.200 ;
        RECT 115.000 29.100 115.400 29.200 ;
        RECT 107.000 26.800 107.400 27.200 ;
        RECT 107.800 23.100 108.200 28.900 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 108.600 26.300 108.900 26.800 ;
        RECT 108.600 25.900 109.000 26.300 ;
        RECT 111.800 25.800 112.200 26.200 ;
        RECT 111.800 25.200 112.100 25.800 ;
        RECT 110.200 24.800 110.600 25.200 ;
        RECT 111.800 24.800 112.200 25.200 ;
        RECT 109.400 19.800 109.800 20.200 ;
        RECT 109.400 19.200 109.700 19.800 ;
        RECT 109.400 18.800 109.800 19.200 ;
        RECT 103.800 16.800 104.200 17.200 ;
        RECT 103.800 15.800 104.200 16.200 ;
        RECT 103.800 15.200 104.100 15.800 ;
        RECT 103.800 14.800 104.200 15.200 ;
        RECT 106.200 14.800 106.600 15.200 ;
        RECT 105.400 13.800 105.800 14.200 ;
        RECT 103.000 9.800 103.400 10.200 ;
        RECT 105.400 9.200 105.700 13.800 ;
        RECT 91.800 8.800 92.200 9.200 ;
        RECT 94.200 8.800 94.600 9.200 ;
        RECT 95.800 8.800 96.200 9.200 ;
        RECT 104.600 9.100 105.000 9.200 ;
        RECT 105.400 9.100 105.800 9.200 ;
        RECT 78.200 6.800 78.600 7.200 ;
        RECT 79.800 6.800 80.200 7.200 ;
        RECT 82.200 6.800 82.600 7.200 ;
        RECT 87.000 6.800 87.400 7.200 ;
        RECT 90.200 6.800 90.600 7.200 ;
        RECT 87.000 6.200 87.300 6.800 ;
        RECT 91.800 6.200 92.100 8.800 ;
        RECT 93.400 6.800 93.800 7.200 ;
        RECT 93.400 6.200 93.700 6.800 ;
        RECT 83.000 5.800 83.400 6.200 ;
        RECT 87.000 5.800 87.400 6.200 ;
        RECT 91.800 5.800 92.200 6.200 ;
        RECT 93.400 5.800 93.800 6.200 ;
        RECT 83.000 5.200 83.300 5.800 ;
        RECT 94.200 5.200 94.500 8.800 ;
        RECT 95.800 7.200 96.100 8.800 ;
        RECT 95.800 6.800 96.200 7.200 ;
        RECT 78.200 4.800 78.600 5.200 ;
        RECT 83.000 4.800 83.400 5.200 ;
        RECT 94.200 4.800 94.600 5.200 ;
        RECT 96.600 5.100 97.000 7.900 ;
        RECT 78.200 4.200 78.500 4.800 ;
        RECT 78.200 3.800 78.600 4.200 ;
        RECT 98.200 3.100 98.600 8.900 ;
        RECT 100.600 7.800 101.000 8.200 ;
        RECT 100.600 7.200 100.900 7.800 ;
        RECT 100.600 6.800 101.000 7.200 ;
        RECT 99.000 5.900 99.400 6.300 ;
        RECT 99.000 5.200 99.300 5.900 ;
        RECT 99.000 4.800 99.400 5.200 ;
        RECT 103.000 3.100 103.400 8.900 ;
        RECT 104.600 8.800 105.800 9.100 ;
        RECT 106.200 8.200 106.500 14.800 ;
        RECT 107.000 12.100 107.400 17.900 ;
        RECT 108.600 17.800 109.000 18.200 ;
        RECT 108.600 9.200 108.900 17.800 ;
        RECT 110.200 15.200 110.500 24.800 ;
        RECT 112.600 23.100 113.000 28.900 ;
        RECT 114.200 28.800 115.400 29.100 ;
        RECT 115.800 28.800 116.200 29.200 ;
        RECT 115.000 18.800 115.400 19.200 ;
        RECT 111.000 16.800 111.400 17.200 ;
        RECT 111.000 16.200 111.300 16.800 ;
        RECT 111.000 15.800 111.400 16.200 ;
        RECT 113.400 15.800 113.800 16.200 ;
        RECT 113.400 15.200 113.700 15.800 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 113.400 14.800 113.800 15.200 ;
        RECT 115.000 14.200 115.300 18.800 ;
        RECT 116.600 16.200 116.900 33.800 ;
        RECT 117.400 21.200 117.700 33.800 ;
        RECT 118.200 23.100 118.600 28.900 ;
        RECT 119.800 22.200 120.100 34.800 ;
        RECT 120.600 34.200 120.900 35.800 ;
        RECT 124.600 35.200 124.900 36.800 ;
        RECT 125.400 35.800 125.800 36.200 ;
        RECT 125.400 35.200 125.700 35.800 ;
        RECT 130.200 35.200 130.500 36.800 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 124.600 34.800 125.000 35.200 ;
        RECT 125.400 34.800 125.800 35.200 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 129.400 34.800 129.800 35.200 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 131.000 34.800 131.400 35.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 120.600 33.800 121.000 34.200 ;
        RECT 121.400 28.800 121.800 29.200 ;
        RECT 121.400 26.200 121.700 28.800 ;
        RECT 122.200 26.800 122.600 27.200 ;
        RECT 121.400 25.800 121.800 26.200 ;
        RECT 121.400 23.800 121.800 24.200 ;
        RECT 118.200 21.800 118.600 22.200 ;
        RECT 119.800 21.800 120.200 22.200 ;
        RECT 117.400 20.800 117.800 21.200 ;
        RECT 118.200 19.200 118.500 21.800 ;
        RECT 118.200 18.800 118.600 19.200 ;
        RECT 121.400 16.200 121.700 23.800 ;
        RECT 115.800 15.800 116.200 16.200 ;
        RECT 116.600 15.800 117.000 16.200 ;
        RECT 120.600 15.800 121.000 16.200 ;
        RECT 121.400 15.800 121.800 16.200 ;
        RECT 115.800 15.200 116.100 15.800 ;
        RECT 115.800 14.800 116.200 15.200 ;
        RECT 116.600 14.800 117.000 15.200 ;
        RECT 119.000 14.800 119.400 15.200 ;
        RECT 116.600 14.200 116.900 14.800 ;
        RECT 119.000 14.200 119.300 14.800 ;
        RECT 120.600 14.200 120.900 15.800 ;
        RECT 121.400 15.200 121.700 15.800 ;
        RECT 121.400 14.800 121.800 15.200 ;
        RECT 110.200 13.800 110.600 14.200 ;
        RECT 115.000 13.800 115.400 14.200 ;
        RECT 116.600 13.800 117.000 14.200 ;
        RECT 119.000 13.800 119.400 14.200 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 110.200 10.200 110.500 13.800 ;
        RECT 110.200 9.800 110.600 10.200 ;
        RECT 119.000 9.200 119.300 13.800 ;
        RECT 120.600 9.200 120.900 13.800 ;
        RECT 108.600 8.800 109.000 9.200 ;
        RECT 106.200 7.800 106.600 8.200 ;
        RECT 110.200 5.100 110.600 7.900 ;
        RECT 111.800 3.100 112.200 8.900 ;
        RECT 114.200 7.800 114.600 8.200 ;
        RECT 114.200 7.200 114.500 7.800 ;
        RECT 114.200 6.800 114.600 7.200 ;
        RECT 114.200 6.100 114.600 6.200 ;
        RECT 115.000 6.100 115.400 6.200 ;
        RECT 114.200 5.800 115.400 6.100 ;
        RECT 116.600 3.100 117.000 8.900 ;
        RECT 119.000 8.800 119.400 9.200 ;
        RECT 120.600 8.800 121.000 9.200 ;
        RECT 119.800 5.100 120.200 7.900 ;
        RECT 121.400 3.100 121.800 8.900 ;
        RECT 122.200 8.200 122.500 26.800 ;
        RECT 123.000 23.100 123.400 28.900 ;
        RECT 123.800 22.200 124.100 34.800 ;
        RECT 125.400 33.800 125.800 34.200 ;
        RECT 125.400 29.200 125.700 33.800 ;
        RECT 125.400 28.800 125.800 29.200 ;
        RECT 124.600 25.100 125.000 27.900 ;
        RECT 125.400 26.800 125.800 27.200 ;
        RECT 125.400 25.200 125.700 26.800 ;
        RECT 125.400 24.800 125.800 25.200 ;
        RECT 123.800 21.800 124.200 22.200 ;
        RECT 126.200 19.200 126.500 34.800 ;
        RECT 128.600 34.200 128.900 34.800 ;
        RECT 128.600 33.800 129.000 34.200 ;
        RECT 127.000 29.800 127.400 30.200 ;
        RECT 127.000 27.200 127.300 29.800 ;
        RECT 129.400 29.200 129.700 34.800 ;
        RECT 131.000 34.200 131.300 34.800 ;
        RECT 131.000 33.800 131.400 34.200 ;
        RECT 133.400 33.200 133.700 34.800 ;
        RECT 134.200 34.200 134.500 46.800 ;
        RECT 135.000 45.100 135.400 47.900 ;
        RECT 140.600 47.200 140.900 49.800 ;
        RECT 143.000 47.200 143.300 52.800 ;
        RECT 143.800 52.200 144.100 55.800 ;
        RECT 144.600 54.200 144.900 63.800 ;
        RECT 147.000 59.200 147.300 66.800 ;
        RECT 151.000 66.200 151.300 71.800 ;
        RECT 151.800 70.200 152.100 74.800 ;
        RECT 153.400 73.800 153.800 74.200 ;
        RECT 153.400 72.200 153.700 73.800 ;
        RECT 153.400 71.800 153.800 72.200 ;
        RECT 154.200 72.100 154.600 77.900 ;
        RECT 155.800 74.200 156.100 85.800 ;
        RECT 162.200 85.200 162.500 85.800 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 163.800 84.200 164.100 104.800 ;
        RECT 167.800 104.200 168.100 106.800 ;
        RECT 167.800 103.800 168.200 104.200 ;
        RECT 165.400 101.800 165.800 102.200 ;
        RECT 165.400 91.200 165.700 101.800 ;
        RECT 166.200 97.800 166.600 98.200 ;
        RECT 166.200 95.200 166.500 97.800 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 167.000 92.100 167.400 97.900 ;
        RECT 168.600 96.200 168.900 111.800 ;
        RECT 171.000 110.200 171.300 111.800 ;
        RECT 171.000 109.800 171.400 110.200 ;
        RECT 171.000 103.100 171.400 108.900 ;
        RECT 172.600 105.200 172.900 115.800 ;
        RECT 173.400 115.100 173.800 115.200 ;
        RECT 174.200 115.100 174.500 125.800 ;
        RECT 175.000 123.200 175.300 125.800 ;
        RECT 177.400 124.800 177.800 125.200 ;
        RECT 177.400 123.200 177.700 124.800 ;
        RECT 175.000 122.800 175.400 123.200 ;
        RECT 177.400 122.800 177.800 123.200 ;
        RECT 173.400 114.800 174.500 115.100 ;
        RECT 175.000 115.800 175.400 116.200 ;
        RECT 180.600 116.100 181.000 116.200 ;
        RECT 179.800 115.800 181.000 116.100 ;
        RECT 172.600 104.800 173.000 105.200 ;
        RECT 173.400 101.200 173.700 114.800 ;
        RECT 175.000 114.200 175.300 115.800 ;
        RECT 179.800 115.200 180.100 115.800 ;
        RECT 175.800 114.800 176.200 115.200 ;
        RECT 179.800 114.800 180.200 115.200 ;
        RECT 180.600 114.800 181.000 115.200 ;
        RECT 175.800 114.200 176.100 114.800 ;
        RECT 175.000 113.800 175.400 114.200 ;
        RECT 175.800 113.800 176.200 114.200 ;
        RECT 178.200 113.800 178.600 114.200 ;
        RECT 179.800 113.800 180.200 114.200 ;
        RECT 176.600 112.800 177.000 113.200 ;
        RECT 175.000 106.800 175.400 107.200 ;
        RECT 174.200 105.800 174.600 106.200 ;
        RECT 174.200 105.200 174.500 105.800 ;
        RECT 174.200 104.800 174.600 105.200 ;
        RECT 173.400 100.800 173.800 101.200 ;
        RECT 175.000 98.100 175.300 106.800 ;
        RECT 175.800 103.100 176.200 108.900 ;
        RECT 176.600 108.200 176.900 112.800 ;
        RECT 178.200 112.200 178.500 113.800 ;
        RECT 179.800 113.200 180.100 113.800 ;
        RECT 179.800 112.800 180.200 113.200 ;
        RECT 178.200 111.800 178.600 112.200 ;
        RECT 180.600 108.200 180.900 114.800 ;
        RECT 176.600 107.800 177.000 108.200 ;
        RECT 176.600 99.100 176.900 107.800 ;
        RECT 177.400 105.100 177.800 107.900 ;
        RECT 180.600 107.800 181.000 108.200 ;
        RECT 181.400 107.200 181.700 153.800 ;
        RECT 182.200 143.100 182.600 148.900 ;
        RECT 183.800 146.100 184.200 146.200 ;
        RECT 183.000 145.800 184.200 146.100 ;
        RECT 183.000 139.200 183.300 145.800 ;
        RECT 183.000 138.800 183.400 139.200 ;
        RECT 184.600 136.800 185.000 137.200 ;
        RECT 184.600 136.200 184.900 136.800 ;
        RECT 184.600 135.800 185.000 136.200 ;
        RECT 182.200 135.100 182.600 135.200 ;
        RECT 183.000 135.100 183.400 135.200 ;
        RECT 182.200 134.800 183.400 135.100 ;
        RECT 186.200 134.200 186.500 161.800 ;
        RECT 188.600 152.100 189.000 157.900 ;
        RECT 189.400 149.200 189.700 166.800 ;
        RECT 191.800 163.100 192.200 168.900 ;
        RECT 194.200 168.800 194.600 169.200 ;
        RECT 195.000 164.200 195.300 174.800 ;
        RECT 196.600 174.100 197.000 174.200 ;
        RECT 199.800 174.100 200.200 174.200 ;
        RECT 200.600 174.100 201.000 174.200 ;
        RECT 196.600 173.800 197.700 174.100 ;
        RECT 199.800 173.800 201.000 174.100 ;
        RECT 197.400 172.200 197.700 173.800 ;
        RECT 196.600 171.800 197.000 172.200 ;
        RECT 197.400 171.800 197.800 172.200 ;
        RECT 200.600 171.800 201.000 172.200 ;
        RECT 203.000 172.100 203.400 177.900 ;
        RECT 204.600 176.800 205.000 177.200 ;
        RECT 204.600 175.200 204.900 176.800 ;
        RECT 204.600 174.800 205.000 175.200 ;
        RECT 207.000 174.800 207.400 175.200 ;
        RECT 196.600 166.200 196.900 171.800 ;
        RECT 197.400 166.800 197.800 167.200 ;
        RECT 197.400 166.200 197.700 166.800 ;
        RECT 196.600 165.800 197.000 166.200 ;
        RECT 197.400 165.800 197.800 166.200 ;
        RECT 199.000 165.800 199.400 166.200 ;
        RECT 199.800 165.800 200.200 166.200 ;
        RECT 195.000 163.800 195.400 164.200 ;
        RECT 190.200 154.800 190.600 155.200 ;
        RECT 190.200 154.200 190.500 154.800 ;
        RECT 190.200 153.800 190.600 154.200 ;
        RECT 193.400 152.100 193.800 157.900 ;
        RECT 196.600 156.200 196.900 165.800 ;
        RECT 199.000 165.200 199.300 165.800 ;
        RECT 199.800 165.200 200.100 165.800 ;
        RECT 199.000 164.800 199.400 165.200 ;
        RECT 199.800 164.800 200.200 165.200 ;
        RECT 200.600 164.200 200.900 171.800 ;
        RECT 201.400 168.800 201.800 169.200 ;
        RECT 201.400 166.200 201.700 168.800 ;
        RECT 203.000 167.800 203.400 168.200 ;
        RECT 203.000 167.200 203.300 167.800 ;
        RECT 203.000 166.800 203.400 167.200 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 202.200 165.800 202.600 166.200 ;
        RECT 201.400 164.800 201.800 165.200 ;
        RECT 199.000 163.800 199.400 164.200 ;
        RECT 200.600 163.800 201.000 164.200 ;
        RECT 199.000 157.200 199.300 163.800 ;
        RECT 201.400 159.200 201.700 164.800 ;
        RECT 201.400 158.800 201.800 159.200 ;
        RECT 202.200 157.200 202.500 165.800 ;
        RECT 199.000 156.800 199.400 157.200 ;
        RECT 202.200 156.800 202.600 157.200 ;
        RECT 194.200 153.800 194.600 154.200 ;
        RECT 194.200 149.200 194.500 153.800 ;
        RECT 195.000 153.100 195.400 155.900 ;
        RECT 196.600 155.800 197.000 156.200 ;
        RECT 207.000 155.200 207.300 174.800 ;
        RECT 207.800 172.100 208.200 177.900 ;
        RECT 208.600 176.200 208.900 206.800 ;
        RECT 211.000 206.200 211.300 208.800 ;
        RECT 211.000 205.800 211.400 206.200 ;
        RECT 210.200 204.800 210.600 205.200 ;
        RECT 210.200 202.200 210.500 204.800 ;
        RECT 213.400 203.100 213.800 208.900 ;
        RECT 215.000 206.800 215.400 207.200 ;
        RECT 216.600 206.800 217.000 207.200 ;
        RECT 215.000 206.200 215.300 206.800 ;
        RECT 215.000 205.800 215.400 206.200 ;
        RECT 209.400 201.800 209.800 202.200 ;
        RECT 210.200 201.800 210.600 202.200 ;
        RECT 209.400 177.100 209.700 201.800 ;
        RECT 211.000 192.100 211.400 197.900 ;
        RECT 211.800 195.800 212.200 196.200 ;
        RECT 211.800 195.200 212.100 195.800 ;
        RECT 211.800 194.800 212.200 195.200 ;
        RECT 214.200 194.800 214.600 195.200 ;
        RECT 210.200 183.100 210.600 188.900 ;
        RECT 211.000 186.100 211.400 186.200 ;
        RECT 211.800 186.100 212.100 194.800 ;
        RECT 214.200 194.200 214.500 194.800 ;
        RECT 214.200 193.800 214.600 194.200 ;
        RECT 215.800 192.100 216.200 197.900 ;
        RECT 216.600 195.200 216.900 206.800 ;
        RECT 218.200 203.100 218.600 208.900 ;
        RECT 219.800 205.100 220.200 207.900 ;
        RECT 221.400 207.100 221.800 207.200 ;
        RECT 222.200 207.100 222.600 207.200 ;
        RECT 221.400 206.800 222.600 207.100 ;
        RECT 223.000 207.100 223.400 207.200 ;
        RECT 223.800 207.100 224.200 207.200 ;
        RECT 223.000 206.800 224.200 207.100 ;
        RECT 223.800 205.800 224.200 206.200 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 223.800 205.200 224.100 205.800 ;
        RECT 224.600 205.200 224.900 205.800 ;
        RECT 220.600 204.800 221.000 205.200 ;
        RECT 223.800 204.800 224.200 205.200 ;
        RECT 224.600 204.800 225.000 205.200 ;
        RECT 225.400 205.100 225.800 205.200 ;
        RECT 226.200 205.100 226.600 205.200 ;
        RECT 225.400 204.800 226.600 205.100 ;
        RECT 220.600 204.100 220.900 204.800 ;
        RECT 219.800 203.800 220.900 204.100 ;
        RECT 216.600 194.800 217.000 195.200 ;
        RECT 216.600 194.200 216.900 194.800 ;
        RECT 216.600 193.800 217.000 194.200 ;
        RECT 217.400 193.100 217.800 195.900 ;
        RECT 219.000 195.100 219.400 195.200 ;
        RECT 219.800 195.100 220.100 203.800 ;
        RECT 221.400 201.800 221.800 202.200 ;
        RECT 226.200 202.100 226.600 202.200 ;
        RECT 227.000 202.100 227.400 202.200 ;
        RECT 226.200 201.800 227.400 202.100 ;
        RECT 220.600 196.100 221.000 196.200 ;
        RECT 221.400 196.100 221.700 201.800 ;
        RECT 220.600 195.800 221.700 196.100 ;
        RECT 219.000 194.800 220.100 195.100 ;
        RECT 218.200 193.800 218.600 194.200 ;
        RECT 211.000 185.800 212.100 186.100 ;
        RECT 214.200 186.800 214.600 187.200 ;
        RECT 214.200 186.300 214.500 186.800 ;
        RECT 214.200 185.900 214.600 186.300 ;
        RECT 210.200 177.100 210.600 177.200 ;
        RECT 209.400 176.800 210.600 177.100 ;
        RECT 208.600 175.800 209.000 176.200 ;
        RECT 208.600 173.800 209.000 174.200 ;
        RECT 208.600 173.200 208.900 173.800 ;
        RECT 208.600 172.800 209.000 173.200 ;
        RECT 209.400 173.100 209.800 175.900 ;
        RECT 210.200 175.800 210.600 176.200 ;
        RECT 210.200 175.200 210.500 175.800 ;
        RECT 210.200 174.800 210.600 175.200 ;
        RECT 211.000 173.200 211.300 185.800 ;
        RECT 215.000 183.100 215.400 188.900 ;
        RECT 217.400 188.800 217.800 189.200 ;
        RECT 216.600 185.100 217.000 187.900 ;
        RECT 217.400 187.200 217.700 188.800 ;
        RECT 217.400 186.800 217.800 187.200 ;
        RECT 218.200 182.200 218.500 193.800 ;
        RECT 219.000 186.800 219.400 187.200 ;
        RECT 219.000 186.200 219.300 186.800 ;
        RECT 219.000 185.800 219.400 186.200 ;
        RECT 219.000 184.800 219.400 185.200 ;
        RECT 219.000 184.200 219.300 184.800 ;
        RECT 219.000 183.800 219.400 184.200 ;
        RECT 218.200 181.800 218.600 182.200 ;
        RECT 215.000 178.100 215.400 178.200 ;
        RECT 215.800 178.100 216.200 178.200 ;
        RECT 215.000 177.800 216.200 178.100 ;
        RECT 215.000 175.800 215.400 176.200 ;
        RECT 215.000 175.200 215.300 175.800 ;
        RECT 215.000 174.800 215.400 175.200 ;
        RECT 211.800 174.100 212.200 174.200 ;
        RECT 212.600 174.100 213.000 174.200 ;
        RECT 211.800 173.800 213.000 174.100 ;
        RECT 213.400 173.800 213.800 174.200 ;
        RECT 211.000 172.800 211.400 173.200 ;
        RECT 207.800 167.800 208.200 168.200 ;
        RECT 207.800 167.200 208.100 167.800 ;
        RECT 207.800 166.800 208.200 167.200 ;
        RECT 208.600 163.100 209.000 168.900 ;
        RECT 211.000 167.200 211.300 172.800 ;
        RECT 213.400 170.200 213.700 173.800 ;
        RECT 214.200 171.800 214.600 172.200 ;
        RECT 218.200 172.100 218.600 177.900 ;
        RECT 219.000 174.800 219.400 175.200 ;
        RECT 219.000 173.200 219.300 174.800 ;
        RECT 219.000 172.800 219.400 173.200 ;
        RECT 213.400 169.800 213.800 170.200 ;
        RECT 211.000 166.800 211.400 167.200 ;
        RECT 212.600 165.900 213.000 166.300 ;
        RECT 212.600 165.200 212.900 165.900 ;
        RECT 212.600 164.800 213.000 165.200 ;
        RECT 213.400 163.100 213.800 168.900 ;
        RECT 212.600 156.800 213.000 157.200 ;
        RECT 211.000 155.800 211.400 156.200 ;
        RECT 211.000 155.200 211.300 155.800 ;
        RECT 199.000 155.100 199.400 155.200 ;
        RECT 199.800 155.100 200.200 155.200 ;
        RECT 199.000 154.800 200.200 155.100 ;
        RECT 200.600 154.800 201.000 155.200 ;
        RECT 203.000 154.800 203.400 155.200 ;
        RECT 207.000 154.800 207.400 155.200 ;
        RECT 208.600 155.100 209.000 155.200 ;
        RECT 209.400 155.100 209.800 155.200 ;
        RECT 208.600 154.800 209.800 155.100 ;
        RECT 211.000 154.800 211.400 155.200 ;
        RECT 197.400 153.800 197.800 154.200 ;
        RECT 195.800 152.800 196.200 153.200 ;
        RECT 187.000 143.100 187.400 148.900 ;
        RECT 187.800 148.800 188.200 149.200 ;
        RECT 189.400 148.800 189.800 149.200 ;
        RECT 194.200 148.800 194.600 149.200 ;
        RECT 195.000 148.800 195.400 149.200 ;
        RECT 187.800 147.200 188.100 148.800 ;
        RECT 187.800 146.800 188.200 147.200 ;
        RECT 188.600 145.100 189.000 147.900 ;
        RECT 189.400 147.800 189.800 148.200 ;
        RECT 189.400 147.200 189.700 147.800 ;
        RECT 189.400 146.800 189.800 147.200 ;
        RECT 192.600 146.800 193.000 147.200 ;
        RECT 187.800 137.100 188.200 137.200 ;
        RECT 188.600 137.100 189.000 137.200 ;
        RECT 187.800 136.800 189.000 137.100 ;
        RECT 183.000 134.100 183.400 134.200 ;
        RECT 183.800 134.100 184.200 134.200 ;
        RECT 183.000 133.800 184.200 134.100 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 185.400 131.800 185.800 132.200 ;
        RECT 182.200 123.100 182.600 128.900 ;
        RECT 183.000 128.800 183.400 129.200 ;
        RECT 183.000 117.100 183.300 128.800 ;
        RECT 183.800 126.800 184.200 127.200 ;
        RECT 183.800 126.200 184.100 126.800 ;
        RECT 183.800 125.800 184.200 126.200 ;
        RECT 185.400 125.200 185.700 131.800 ;
        RECT 185.400 124.800 185.800 125.200 ;
        RECT 182.200 116.800 183.300 117.100 ;
        RECT 183.800 123.800 184.200 124.200 ;
        RECT 182.200 116.200 182.500 116.800 ;
        RECT 182.200 115.800 182.600 116.200 ;
        RECT 183.000 115.800 183.400 116.200 ;
        RECT 183.000 115.200 183.300 115.800 ;
        RECT 183.000 114.800 183.400 115.200 ;
        RECT 183.800 113.100 184.100 123.800 ;
        RECT 186.200 120.200 186.500 133.800 ;
        RECT 189.400 133.200 189.700 146.800 ;
        RECT 190.200 145.800 190.600 146.200 ;
        RECT 190.200 145.200 190.500 145.800 ;
        RECT 192.600 145.200 192.900 146.800 ;
        RECT 193.400 146.100 193.800 146.200 ;
        RECT 194.200 146.100 194.600 146.200 ;
        RECT 193.400 145.800 194.600 146.100 ;
        RECT 190.200 144.800 190.600 145.200 ;
        RECT 192.600 144.800 193.000 145.200 ;
        RECT 194.200 144.800 194.600 145.200 ;
        RECT 189.400 132.800 189.800 133.200 ;
        RECT 191.000 132.100 191.400 137.900 ;
        RECT 192.600 135.800 193.000 136.200 ;
        RECT 192.600 135.200 192.900 135.800 ;
        RECT 192.600 134.800 193.000 135.200 ;
        RECT 194.200 133.200 194.500 144.800 ;
        RECT 195.000 134.200 195.300 148.800 ;
        RECT 195.800 147.200 196.100 152.800 ;
        RECT 195.800 146.800 196.200 147.200 ;
        RECT 196.600 145.100 197.000 147.900 ;
        RECT 195.000 133.800 195.400 134.200 ;
        RECT 194.200 132.800 194.600 133.200 ;
        RECT 193.400 131.800 193.800 132.200 ;
        RECT 195.800 132.100 196.200 137.900 ;
        RECT 197.400 137.200 197.700 153.800 ;
        RECT 200.600 153.200 200.900 154.800 ;
        RECT 203.000 153.200 203.300 154.800 ;
        RECT 204.600 154.100 205.000 154.200 ;
        RECT 205.400 154.100 205.800 154.200 ;
        RECT 204.600 153.800 205.800 154.100 ;
        RECT 207.000 154.100 207.400 154.200 ;
        RECT 207.800 154.100 208.200 154.200 ;
        RECT 207.000 153.800 208.200 154.100 ;
        RECT 200.600 152.800 201.000 153.200 ;
        RECT 203.000 152.800 203.400 153.200 ;
        RECT 198.200 151.800 198.600 152.200 ;
        RECT 198.200 151.200 198.500 151.800 ;
        RECT 198.200 150.800 198.600 151.200 ;
        RECT 200.600 149.200 200.900 152.800 ;
        RECT 198.200 143.100 198.600 148.900 ;
        RECT 199.000 148.800 199.400 149.200 ;
        RECT 200.600 148.800 201.000 149.200 ;
        RECT 199.000 148.200 199.300 148.800 ;
        RECT 199.000 147.800 199.400 148.200 ;
        RECT 199.000 146.800 199.400 147.200 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 199.000 146.300 199.300 146.800 ;
        RECT 199.000 145.900 199.400 146.300 ;
        RECT 202.200 146.200 202.500 146.800 ;
        RECT 202.200 145.800 202.600 146.200 ;
        RECT 203.000 143.100 203.400 148.900 ;
        RECT 204.600 148.200 204.900 153.800 ;
        RECT 210.200 151.800 210.600 152.200 ;
        RECT 205.400 149.800 205.800 150.200 ;
        RECT 205.400 149.200 205.700 149.800 ;
        RECT 205.400 148.800 205.800 149.200 ;
        RECT 207.000 148.800 207.400 149.200 ;
        RECT 207.000 148.200 207.300 148.800 ;
        RECT 204.600 147.800 205.000 148.200 ;
        RECT 207.000 147.800 207.400 148.200 ;
        RECT 207.000 146.800 207.400 147.200 ;
        RECT 207.000 146.200 207.300 146.800 ;
        RECT 207.000 145.800 207.400 146.200 ;
        RECT 207.800 145.100 208.200 147.900 ;
        RECT 209.400 143.100 209.800 148.900 ;
        RECT 210.200 146.300 210.500 151.800 ;
        RECT 210.200 145.900 210.600 146.300 ;
        RECT 210.200 145.800 210.500 145.900 ;
        RECT 206.200 141.800 206.600 142.200 ;
        RECT 199.800 140.800 200.200 141.200 ;
        RECT 197.400 136.800 197.800 137.200 ;
        RECT 198.200 136.800 198.600 137.200 ;
        RECT 198.200 136.200 198.500 136.800 ;
        RECT 196.600 133.800 197.000 134.200 ;
        RECT 187.000 123.100 187.400 128.900 ;
        RECT 189.400 128.800 189.800 129.200 ;
        RECT 189.400 128.200 189.700 128.800 ;
        RECT 187.800 127.800 188.200 128.200 ;
        RECT 187.800 127.200 188.100 127.800 ;
        RECT 187.800 126.800 188.200 127.200 ;
        RECT 188.600 125.100 189.000 127.900 ;
        RECT 189.400 127.800 189.800 128.200 ;
        RECT 193.400 127.200 193.700 131.800 ;
        RECT 195.800 130.800 196.200 131.200 ;
        RECT 195.800 129.200 196.100 130.800 ;
        RECT 195.800 128.800 196.200 129.200 ;
        RECT 196.600 127.200 196.900 133.800 ;
        RECT 197.400 133.100 197.800 135.900 ;
        RECT 198.200 135.800 198.600 136.200 ;
        RECT 199.800 135.200 200.100 140.800 ;
        RECT 203.000 136.800 203.400 137.200 ;
        RECT 200.600 135.800 201.000 136.200 ;
        RECT 199.800 134.800 200.200 135.200 ;
        RECT 198.200 131.800 198.600 132.200 ;
        RECT 193.400 126.800 193.800 127.200 ;
        RECT 196.600 126.800 197.000 127.200 ;
        RECT 198.200 127.100 198.500 131.800 ;
        RECT 199.800 130.200 200.100 134.800 ;
        RECT 200.600 134.200 200.900 135.800 ;
        RECT 203.000 134.200 203.300 136.800 ;
        RECT 206.200 136.200 206.500 141.800 ;
        RECT 211.000 139.200 211.300 154.800 ;
        RECT 212.600 154.200 212.900 156.800 ;
        RECT 213.400 156.100 213.800 156.200 ;
        RECT 214.200 156.100 214.500 171.800 ;
        RECT 216.600 169.800 217.000 170.200 ;
        RECT 215.000 165.100 215.400 167.900 ;
        RECT 215.800 167.800 216.200 168.200 ;
        RECT 215.800 167.200 216.100 167.800 ;
        RECT 215.800 166.800 216.200 167.200 ;
        RECT 216.600 159.200 216.900 169.800 ;
        RECT 218.200 166.800 218.600 167.200 ;
        RECT 217.400 165.800 217.800 166.200 ;
        RECT 217.400 165.200 217.700 165.800 ;
        RECT 218.200 165.200 218.500 166.800 ;
        RECT 219.800 166.200 220.100 194.800 ;
        RECT 220.600 191.800 221.000 192.200 ;
        RECT 221.400 191.800 221.800 192.200 ;
        RECT 223.800 192.100 224.200 197.900 ;
        RECT 224.600 195.800 225.000 196.200 ;
        RECT 224.600 195.200 224.900 195.800 ;
        RECT 224.600 194.800 225.000 195.200 ;
        RECT 225.400 194.800 225.800 195.200 ;
        RECT 220.600 191.200 220.900 191.800 ;
        RECT 220.600 190.800 221.000 191.200 ;
        RECT 221.400 190.200 221.700 191.800 ;
        RECT 221.400 189.800 221.800 190.200 ;
        RECT 223.000 189.800 223.400 190.200 ;
        RECT 223.000 187.200 223.300 189.800 ;
        RECT 225.400 189.200 225.700 194.800 ;
        RECT 228.600 192.100 229.000 197.900 ;
        RECT 230.200 193.100 230.600 195.900 ;
        RECT 225.400 188.800 225.800 189.200 ;
        RECT 222.200 186.800 222.600 187.200 ;
        RECT 223.000 186.800 223.400 187.200 ;
        RECT 227.000 187.100 227.400 187.200 ;
        RECT 227.800 187.100 228.200 187.200 ;
        RECT 227.000 186.800 228.200 187.100 ;
        RECT 221.400 185.800 221.800 186.200 ;
        RECT 221.400 184.200 221.700 185.800 ;
        RECT 221.400 183.800 221.800 184.200 ;
        RECT 222.200 181.200 222.500 186.800 ;
        RECT 227.000 185.800 227.400 186.200 ;
        RECT 227.000 185.200 227.300 185.800 ;
        RECT 224.600 185.100 225.000 185.200 ;
        RECT 225.400 185.100 225.800 185.200 ;
        RECT 224.600 184.800 225.800 185.100 ;
        RECT 227.000 184.800 227.400 185.200 ;
        RECT 220.600 180.800 221.000 181.200 ;
        RECT 222.200 180.800 222.600 181.200 ;
        RECT 220.600 174.200 220.900 180.800 ;
        RECT 221.400 175.100 221.800 175.200 ;
        RECT 221.400 174.800 222.600 175.100 ;
        RECT 222.200 174.700 222.600 174.800 ;
        RECT 220.600 173.800 221.000 174.200 ;
        RECT 220.600 167.200 220.900 173.800 ;
        RECT 223.000 172.100 223.400 177.900 ;
        RECT 225.400 177.800 225.800 178.200 ;
        RECT 224.600 173.100 225.000 175.900 ;
        RECT 225.400 174.200 225.700 177.800 ;
        RECT 227.000 176.200 227.300 184.800 ;
        RECT 230.200 181.800 230.600 182.200 ;
        RECT 226.200 176.100 226.600 176.200 ;
        RECT 227.000 176.100 227.400 176.200 ;
        RECT 226.200 175.800 227.400 176.100 ;
        RECT 229.400 175.800 229.800 176.200 ;
        RECT 229.400 175.200 229.700 175.800 ;
        RECT 227.800 174.800 228.200 175.200 ;
        RECT 229.400 174.800 229.800 175.200 ;
        RECT 227.800 174.200 228.100 174.800 ;
        RECT 230.200 174.200 230.500 181.800 ;
        RECT 225.400 173.800 225.800 174.200 ;
        RECT 227.800 173.800 228.200 174.200 ;
        RECT 230.200 173.800 230.600 174.200 ;
        RECT 220.600 166.800 221.000 167.200 ;
        RECT 221.400 166.800 221.800 167.200 ;
        RECT 219.800 165.800 220.200 166.200 ;
        RECT 217.400 164.800 217.800 165.200 ;
        RECT 218.200 164.800 218.600 165.200 ;
        RECT 216.600 158.800 217.000 159.200 ;
        RECT 216.600 158.200 216.900 158.800 ;
        RECT 216.600 157.800 217.000 158.200 ;
        RECT 213.400 155.800 214.500 156.100 ;
        RECT 216.600 156.800 217.000 157.200 ;
        RECT 213.400 155.100 213.800 155.200 ;
        RECT 214.200 155.100 214.600 155.200 ;
        RECT 213.400 154.800 214.600 155.100 ;
        RECT 215.000 154.800 215.400 155.200 ;
        RECT 215.800 154.800 216.200 155.200 ;
        RECT 212.600 153.800 213.000 154.200 ;
        RECT 215.000 152.200 215.300 154.800 ;
        RECT 215.800 154.200 216.100 154.800 ;
        RECT 215.800 153.800 216.200 154.200 ;
        RECT 215.000 151.800 215.400 152.200 ;
        RECT 216.600 149.200 216.900 156.800 ;
        RECT 217.400 153.800 217.800 154.200 ;
        RECT 213.400 145.800 213.800 146.200 ;
        RECT 211.000 138.800 211.400 139.200 ;
        RECT 207.800 137.100 208.200 137.200 ;
        RECT 208.600 137.100 209.000 137.200 ;
        RECT 207.800 136.800 209.000 137.100 ;
        RECT 204.600 135.800 205.000 136.200 ;
        RECT 206.200 135.800 206.600 136.200 ;
        RECT 207.000 136.100 207.400 136.200 ;
        RECT 207.800 136.100 208.200 136.200 ;
        RECT 207.000 135.800 208.200 136.100 ;
        RECT 204.600 135.200 204.900 135.800 ;
        RECT 204.600 134.800 205.000 135.200 ;
        RECT 206.200 135.100 206.600 135.200 ;
        RECT 207.000 135.100 207.400 135.200 ;
        RECT 206.200 134.800 207.400 135.100 ;
        RECT 207.800 134.800 208.200 135.200 ;
        RECT 207.800 134.200 208.100 134.800 ;
        RECT 200.600 133.800 201.000 134.200 ;
        RECT 203.000 133.800 203.400 134.200 ;
        RECT 207.800 133.800 208.200 134.200 ;
        RECT 201.400 132.800 201.800 133.200 ;
        RECT 203.800 132.800 204.200 133.200 ;
        RECT 201.400 132.200 201.700 132.800 ;
        RECT 201.400 131.800 201.800 132.200 ;
        RECT 199.800 129.800 200.200 130.200 ;
        RECT 203.800 129.200 204.100 132.800 ;
        RECT 207.000 131.800 207.400 132.200 ;
        RECT 211.000 132.100 211.400 137.900 ;
        RECT 213.400 134.200 213.700 145.800 ;
        RECT 214.200 143.100 214.600 148.900 ;
        RECT 216.600 148.800 217.000 149.200 ;
        RECT 217.400 147.200 217.700 153.800 ;
        RECT 219.000 152.100 219.400 157.900 ;
        RECT 219.800 152.200 220.100 165.800 ;
        RECT 220.600 154.200 220.900 166.800 ;
        RECT 221.400 156.200 221.700 166.800 ;
        RECT 223.000 165.100 223.400 165.200 ;
        RECT 223.800 165.100 224.200 165.200 ;
        RECT 223.000 164.800 224.200 165.100 ;
        RECT 227.800 164.800 228.200 165.200 ;
        RECT 222.200 161.800 222.600 162.200 ;
        RECT 222.200 156.200 222.500 161.800 ;
        RECT 221.400 155.800 221.800 156.200 ;
        RECT 222.200 155.800 222.600 156.200 ;
        RECT 221.400 155.100 221.800 155.200 ;
        RECT 222.200 155.100 222.600 155.200 ;
        RECT 221.400 154.800 222.600 155.100 ;
        RECT 220.600 153.800 221.000 154.200 ;
        RECT 219.800 151.800 220.200 152.200 ;
        RECT 223.800 152.100 224.200 157.900 ;
        RECT 226.200 156.800 226.600 157.200 ;
        RECT 226.200 156.200 226.500 156.800 ;
        RECT 224.600 154.800 225.000 155.200 ;
        RECT 224.600 154.200 224.900 154.800 ;
        RECT 224.600 153.800 225.000 154.200 ;
        RECT 217.400 146.800 217.800 147.200 ;
        RECT 215.000 145.800 215.400 146.200 ;
        RECT 217.400 146.100 217.800 146.200 ;
        RECT 218.200 146.100 218.600 146.200 ;
        RECT 217.400 145.800 218.600 146.100 ;
        RECT 219.000 146.100 219.400 146.200 ;
        RECT 219.800 146.100 220.200 146.200 ;
        RECT 219.000 145.800 220.200 146.100 ;
        RECT 214.200 135.800 214.600 136.200 ;
        RECT 214.200 135.200 214.500 135.800 ;
        RECT 214.200 134.800 214.600 135.200 ;
        RECT 213.400 133.800 213.800 134.200 ;
        RECT 203.000 128.800 203.400 129.200 ;
        RECT 203.800 128.800 204.200 129.200 ;
        RECT 197.400 126.800 198.500 127.100 ;
        RECT 200.600 127.800 201.000 128.200 ;
        RECT 190.200 126.100 190.600 126.200 ;
        RECT 191.000 126.100 191.400 126.200 ;
        RECT 190.200 125.800 191.400 126.100 ;
        RECT 194.200 125.800 194.600 126.200 ;
        RECT 189.400 124.800 189.800 125.200 ;
        RECT 189.400 124.200 189.700 124.800 ;
        RECT 189.400 123.800 189.800 124.200 ;
        RECT 188.600 121.800 189.000 122.200 ;
        RECT 186.200 119.800 186.600 120.200 ;
        RECT 184.600 117.800 185.000 118.200 ;
        RECT 184.600 114.200 184.900 117.800 ;
        RECT 188.600 117.200 188.900 121.800 ;
        RECT 188.600 116.800 189.000 117.200 ;
        RECT 192.600 116.800 193.000 117.200 ;
        RECT 188.600 116.200 188.900 116.800 ;
        RECT 188.600 115.800 189.000 116.200 ;
        RECT 192.600 115.200 192.900 116.800 ;
        RECT 185.400 115.100 185.800 115.200 ;
        RECT 186.200 115.100 186.600 115.200 ;
        RECT 185.400 114.800 186.600 115.100 ;
        RECT 187.800 115.100 188.200 115.200 ;
        RECT 188.600 115.100 189.000 115.200 ;
        RECT 187.800 114.800 189.000 115.100 ;
        RECT 192.600 114.800 193.000 115.200 ;
        RECT 184.600 113.800 185.000 114.200 ;
        RECT 185.400 114.100 185.800 114.200 ;
        RECT 186.200 114.100 186.600 114.200 ;
        RECT 185.400 113.800 186.600 114.100 ;
        RECT 191.800 113.800 192.200 114.200 ;
        RECT 183.800 112.800 184.900 113.100 ;
        RECT 183.000 112.100 183.400 112.200 ;
        RECT 183.800 112.100 184.200 112.200 ;
        RECT 183.000 111.800 184.200 112.100 ;
        RECT 183.800 110.800 184.200 111.200 ;
        RECT 183.800 107.200 184.100 110.800 ;
        RECT 184.600 109.200 184.900 112.800 ;
        RECT 191.800 112.200 192.100 113.800 ;
        RECT 193.400 113.100 193.800 115.900 ;
        RECT 191.800 111.800 192.200 112.200 ;
        RECT 186.200 109.800 186.600 110.200 ;
        RECT 184.600 108.800 185.000 109.200 ;
        RECT 186.200 107.200 186.500 109.800 ;
        RECT 178.200 106.800 178.600 107.200 ;
        RECT 180.600 106.800 181.000 107.200 ;
        RECT 181.400 106.800 181.800 107.200 ;
        RECT 183.000 106.800 183.400 107.200 ;
        RECT 183.800 106.800 184.200 107.200 ;
        RECT 186.200 106.800 186.600 107.200 ;
        RECT 187.000 106.800 187.400 107.200 ;
        RECT 188.600 107.100 189.000 107.200 ;
        RECT 189.400 107.100 189.800 107.200 ;
        RECT 188.600 106.800 189.800 107.100 ;
        RECT 178.200 106.200 178.500 106.800 ;
        RECT 178.200 105.800 178.600 106.200 ;
        RECT 179.800 105.800 180.200 106.200 ;
        RECT 179.800 105.200 180.100 105.800 ;
        RECT 180.600 105.200 180.900 106.800 ;
        RECT 183.000 106.200 183.300 106.800 ;
        RECT 181.400 106.100 181.800 106.200 ;
        RECT 182.200 106.100 182.600 106.200 ;
        RECT 181.400 105.800 182.600 106.100 ;
        RECT 183.000 105.800 183.400 106.200 ;
        RECT 179.800 104.800 180.200 105.200 ;
        RECT 180.600 104.800 181.000 105.200 ;
        RECT 176.600 98.800 177.700 99.100 ;
        RECT 175.800 98.100 176.200 98.200 ;
        RECT 168.600 95.800 169.000 96.200 ;
        RECT 170.200 93.100 170.600 95.900 ;
        RECT 169.400 91.800 169.800 92.200 ;
        RECT 171.800 92.100 172.200 97.900 ;
        RECT 175.000 97.800 176.200 98.100 ;
        RECT 174.200 96.800 174.600 97.200 ;
        RECT 174.200 95.200 174.500 96.800 ;
        RECT 175.800 95.200 176.100 97.800 ;
        RECT 174.200 94.800 174.600 95.200 ;
        RECT 175.800 94.800 176.200 95.200 ;
        RECT 176.600 92.100 177.000 97.900 ;
        RECT 169.400 91.200 169.700 91.800 ;
        RECT 165.400 90.800 165.800 91.200 ;
        RECT 167.000 90.800 167.400 91.200 ;
        RECT 169.400 90.800 169.800 91.200 ;
        RECT 165.400 89.100 165.800 89.200 ;
        RECT 166.200 89.100 166.600 89.200 ;
        RECT 165.400 88.800 166.600 89.100 ;
        RECT 164.600 88.100 165.000 88.200 ;
        RECT 165.400 88.100 165.800 88.200 ;
        RECT 164.600 87.800 165.800 88.100 ;
        RECT 167.000 86.200 167.300 90.800 ;
        RECT 177.400 88.200 177.700 98.800 ;
        RECT 180.600 97.100 181.000 97.200 ;
        RECT 181.400 97.100 181.800 97.200 ;
        RECT 180.600 96.800 181.800 97.100 ;
        RECT 183.000 95.800 183.400 96.200 ;
        RECT 183.000 95.200 183.300 95.800 ;
        RECT 179.800 95.100 180.200 95.200 ;
        RECT 180.600 95.100 181.000 95.200 ;
        RECT 179.800 94.800 181.000 95.100 ;
        RECT 183.000 94.800 183.400 95.200 ;
        RECT 179.000 93.800 179.400 94.200 ;
        RECT 179.800 93.800 180.200 94.200 ;
        RECT 179.000 92.200 179.300 93.800 ;
        RECT 179.000 91.800 179.400 92.200 ;
        RECT 179.800 90.200 180.100 93.800 ;
        RECT 183.000 91.800 183.400 92.200 ;
        RECT 179.800 89.800 180.200 90.200 ;
        RECT 183.000 89.200 183.300 91.800 ;
        RECT 183.800 90.200 184.100 106.800 ;
        RECT 187.000 106.200 187.300 106.800 ;
        RECT 187.000 105.800 187.400 106.200 ;
        RECT 189.400 106.100 189.800 106.200 ;
        RECT 188.600 105.800 189.800 106.100 ;
        RECT 187.000 105.200 187.300 105.800 ;
        RECT 185.400 105.100 185.800 105.200 ;
        RECT 186.200 105.100 186.600 105.200 ;
        RECT 185.400 104.800 186.600 105.100 ;
        RECT 187.000 104.800 187.400 105.200 ;
        RECT 187.000 95.100 187.400 95.200 ;
        RECT 187.800 95.100 188.200 95.200 ;
        RECT 187.000 94.800 188.200 95.100 ;
        RECT 188.600 94.200 188.900 105.800 ;
        RECT 189.400 105.100 189.800 105.200 ;
        RECT 190.200 105.100 190.600 105.200 ;
        RECT 189.400 104.800 190.600 105.100 ;
        RECT 191.800 101.800 192.200 102.200 ;
        RECT 190.200 98.800 190.600 99.200 ;
        RECT 184.600 94.100 185.000 94.200 ;
        RECT 185.400 94.100 185.800 94.200 ;
        RECT 184.600 93.800 185.800 94.100 ;
        RECT 187.000 93.800 187.400 94.200 ;
        RECT 188.600 94.100 189.000 94.200 ;
        RECT 187.800 93.800 189.000 94.100 ;
        RECT 186.200 91.800 186.600 92.200 ;
        RECT 183.800 89.800 184.200 90.200 ;
        RECT 183.000 88.800 183.400 89.200 ;
        RECT 168.600 88.100 169.000 88.200 ;
        RECT 169.400 88.100 169.800 88.200 ;
        RECT 168.600 87.800 169.800 88.100 ;
        RECT 176.600 87.800 177.000 88.200 ;
        RECT 177.400 87.800 177.800 88.200 ;
        RECT 179.000 87.800 179.400 88.200 ;
        RECT 183.800 87.800 184.200 88.200 ;
        RECT 176.600 87.200 176.900 87.800 ;
        RECT 179.000 87.200 179.300 87.800 ;
        RECT 183.800 87.200 184.100 87.800 ;
        RECT 167.800 87.100 168.200 87.200 ;
        RECT 168.600 87.100 169.000 87.200 ;
        RECT 167.800 86.800 169.000 87.100 ;
        RECT 171.000 87.100 171.400 87.200 ;
        RECT 171.800 87.100 172.200 87.200 ;
        RECT 171.000 86.800 172.200 87.100 ;
        RECT 176.600 86.800 177.000 87.200 ;
        RECT 179.000 86.800 179.400 87.200 ;
        RECT 180.600 87.100 181.000 87.200 ;
        RECT 180.600 86.800 182.500 87.100 ;
        RECT 183.800 86.800 184.200 87.200 ;
        RECT 185.400 86.800 185.800 87.200 ;
        RECT 167.000 85.800 167.400 86.200 ;
        RECT 168.600 85.800 169.000 86.200 ;
        RECT 170.200 85.800 170.600 86.200 ;
        RECT 171.800 85.800 172.200 86.200 ;
        RECT 176.600 85.800 177.000 86.200 ;
        RECT 178.200 86.100 178.600 86.200 ;
        RECT 179.000 86.100 179.400 86.200 ;
        RECT 178.200 85.800 179.400 86.100 ;
        RECT 179.800 85.800 180.200 86.200 ;
        RECT 180.600 86.100 181.000 86.200 ;
        RECT 181.400 86.100 181.800 86.200 ;
        RECT 180.600 85.800 181.800 86.100 ;
        RECT 165.400 85.100 165.800 85.200 ;
        RECT 166.200 85.100 166.600 85.200 ;
        RECT 165.400 84.800 166.600 85.100 ;
        RECT 167.000 84.200 167.300 85.800 ;
        RECT 168.600 85.200 168.900 85.800 ;
        RECT 168.600 84.800 169.000 85.200 ;
        RECT 159.800 83.800 160.200 84.200 ;
        RECT 163.800 83.800 164.200 84.200 ;
        RECT 167.000 83.800 167.400 84.200 ;
        RECT 159.800 79.200 160.100 83.800 ;
        RECT 163.800 81.200 164.100 83.800 ;
        RECT 164.600 81.800 165.000 82.200 ;
        RECT 163.800 80.800 164.200 81.200 ;
        RECT 159.800 78.800 160.200 79.200 ;
        RECT 155.800 74.100 156.200 74.200 ;
        RECT 155.000 73.800 156.200 74.100 ;
        RECT 159.800 74.100 160.200 74.200 ;
        RECT 160.600 74.100 161.000 74.200 ;
        RECT 159.800 73.800 161.000 74.100 ;
        RECT 151.800 69.800 152.200 70.200 ;
        RECT 153.400 66.200 153.700 71.800 ;
        RECT 155.000 66.200 155.300 73.800 ;
        RECT 155.800 72.100 156.200 72.200 ;
        RECT 156.600 72.100 157.000 72.200 ;
        RECT 155.800 71.800 157.000 72.100 ;
        RECT 158.200 71.800 158.600 72.200 ;
        RECT 158.200 71.200 158.500 71.800 ;
        RECT 158.200 70.800 158.600 71.200 ;
        RECT 160.600 70.100 160.900 73.800 ;
        RECT 161.400 73.100 161.800 75.900 ;
        RECT 163.000 72.100 163.400 77.900 ;
        RECT 164.600 75.200 164.900 81.800 ;
        RECT 164.600 74.800 165.000 75.200 ;
        RECT 165.400 73.800 165.800 74.200 ;
        RECT 165.400 72.200 165.700 73.800 ;
        RECT 165.400 71.800 165.800 72.200 ;
        RECT 167.800 72.100 168.200 77.900 ;
        RECT 168.600 70.200 168.900 84.800 ;
        RECT 170.200 79.200 170.500 85.800 ;
        RECT 171.800 84.200 172.100 85.800 ;
        RECT 174.200 84.800 174.600 85.200 ;
        RECT 175.000 85.100 175.400 85.200 ;
        RECT 175.800 85.100 176.200 85.200 ;
        RECT 175.000 84.800 176.200 85.100 ;
        RECT 171.800 83.800 172.200 84.200 ;
        RECT 170.200 78.800 170.600 79.200 ;
        RECT 172.600 76.100 173.000 76.200 ;
        RECT 173.400 76.100 173.800 76.200 ;
        RECT 172.600 75.800 173.800 76.100 ;
        RECT 174.200 75.200 174.500 84.800 ;
        RECT 176.600 84.200 176.900 85.800 ;
        RECT 179.800 85.200 180.100 85.800 ;
        RECT 179.800 84.800 180.200 85.200 ;
        RECT 182.200 85.100 182.500 86.800 ;
        RECT 183.800 85.800 184.200 86.200 ;
        RECT 183.800 85.200 184.100 85.800 ;
        RECT 181.400 84.800 182.500 85.100 ;
        RECT 183.000 84.800 183.400 85.200 ;
        RECT 183.800 84.800 184.200 85.200 ;
        RECT 176.600 83.800 177.000 84.200 ;
        RECT 178.200 81.800 178.600 82.200 ;
        RECT 178.200 79.200 178.500 81.800 ;
        RECT 181.400 79.200 181.700 84.800 ;
        RECT 183.000 81.200 183.300 84.800 ;
        RECT 185.400 83.200 185.700 86.800 ;
        RECT 186.200 84.200 186.500 91.800 ;
        RECT 187.000 86.200 187.300 93.800 ;
        RECT 187.000 85.800 187.400 86.200 ;
        RECT 187.000 84.800 187.400 85.200 ;
        RECT 186.200 83.800 186.600 84.200 ;
        RECT 185.400 82.800 185.800 83.200 ;
        RECT 183.000 80.800 183.400 81.200 ;
        RECT 178.200 78.800 178.600 79.200 ;
        RECT 181.400 78.800 181.800 79.200 ;
        RECT 179.800 77.100 180.200 77.200 ;
        RECT 180.600 77.100 181.000 77.200 ;
        RECT 179.800 76.800 181.000 77.100 ;
        RECT 184.600 76.800 185.000 77.200 ;
        RECT 184.600 76.200 184.900 76.800 ;
        RECT 186.200 76.200 186.500 83.800 ;
        RECT 187.000 79.200 187.300 84.800 ;
        RECT 187.800 82.200 188.100 93.800 ;
        RECT 189.400 91.800 189.800 92.200 ;
        RECT 189.400 90.200 189.700 91.800 ;
        RECT 189.400 89.800 189.800 90.200 ;
        RECT 189.400 87.800 189.800 88.200 ;
        RECT 189.400 86.200 189.700 87.800 ;
        RECT 190.200 86.200 190.500 98.800 ;
        RECT 191.800 97.200 192.100 101.800 ;
        RECT 191.800 96.800 192.200 97.200 ;
        RECT 191.800 95.800 192.200 96.200 ;
        RECT 191.800 95.200 192.100 95.800 ;
        RECT 194.200 95.200 194.500 125.800 ;
        RECT 195.000 112.100 195.400 117.900 ;
        RECT 195.800 115.800 196.200 116.200 ;
        RECT 195.800 115.100 196.100 115.800 ;
        RECT 195.800 114.700 196.200 115.100 ;
        RECT 196.600 114.200 196.900 126.800 ;
        RECT 197.400 118.200 197.700 126.800 ;
        RECT 200.600 126.200 200.900 127.800 ;
        RECT 203.000 127.200 203.300 128.800 ;
        RECT 203.000 126.800 203.400 127.200 ;
        RECT 207.000 126.200 207.300 131.800 ;
        RECT 208.600 130.800 209.000 131.200 ;
        RECT 207.800 126.800 208.200 127.200 ;
        RECT 207.800 126.200 208.100 126.800 ;
        RECT 208.600 126.200 208.900 130.800 ;
        RECT 213.400 128.800 213.800 129.200 ;
        RECT 210.200 128.100 210.600 128.200 ;
        RECT 211.000 128.100 211.400 128.200 ;
        RECT 210.200 127.800 211.400 128.100 ;
        RECT 213.400 127.200 213.700 128.800 ;
        RECT 213.400 126.800 213.800 127.200 ;
        RECT 198.200 125.800 198.600 126.200 ;
        RECT 199.000 126.100 199.400 126.200 ;
        RECT 199.800 126.100 200.200 126.200 ;
        RECT 199.000 125.800 200.200 126.100 ;
        RECT 200.600 125.800 201.000 126.200 ;
        RECT 202.200 126.100 202.600 126.200 ;
        RECT 203.000 126.100 203.400 126.200 ;
        RECT 202.200 125.800 203.400 126.100 ;
        RECT 204.600 125.800 205.000 126.200 ;
        RECT 207.000 125.800 207.400 126.200 ;
        RECT 207.800 125.800 208.200 126.200 ;
        RECT 208.600 125.800 209.000 126.200 ;
        RECT 209.400 126.100 209.800 126.200 ;
        RECT 210.200 126.100 210.600 126.200 ;
        RECT 209.400 125.800 210.600 126.100 ;
        RECT 198.200 125.200 198.500 125.800 ;
        RECT 198.200 124.800 198.600 125.200 ;
        RECT 203.000 124.800 203.400 125.200 ;
        RECT 197.400 117.800 197.800 118.200 ;
        RECT 196.600 113.800 197.000 114.200 ;
        RECT 199.800 112.100 200.200 117.900 ;
        RECT 201.400 117.100 201.800 117.200 ;
        RECT 202.200 117.100 202.600 117.200 ;
        RECT 201.400 116.800 202.600 117.100 ;
        RECT 203.000 114.200 203.300 124.800 ;
        RECT 203.800 114.800 204.200 115.200 ;
        RECT 203.000 113.800 203.400 114.200 ;
        RECT 203.800 110.200 204.100 114.800 ;
        RECT 204.600 112.200 204.900 125.800 ;
        RECT 205.400 124.800 205.800 125.200 ;
        RECT 205.400 122.200 205.700 124.800 ;
        RECT 205.400 121.800 205.800 122.200 ;
        RECT 205.400 115.100 205.800 115.200 ;
        RECT 206.200 115.100 206.600 115.200 ;
        RECT 205.400 114.800 206.600 115.100 ;
        RECT 207.000 114.800 207.400 115.200 ;
        RECT 207.800 114.800 208.200 115.200 ;
        RECT 204.600 111.800 205.000 112.200 ;
        RECT 203.800 109.800 204.200 110.200 ;
        RECT 195.800 103.100 196.200 108.900 ;
        RECT 197.400 106.800 197.800 107.200 ;
        RECT 197.400 106.200 197.700 106.800 ;
        RECT 197.400 105.800 197.800 106.200 ;
        RECT 200.600 103.100 201.000 108.900 ;
        RECT 201.400 106.800 201.800 107.200 ;
        RECT 201.400 98.200 201.700 106.800 ;
        RECT 202.200 105.100 202.600 107.900 ;
        RECT 204.600 106.200 204.900 111.800 ;
        RECT 207.000 109.200 207.300 114.800 ;
        RECT 207.800 114.200 208.100 114.800 ;
        RECT 208.600 114.200 208.900 125.800 ;
        RECT 210.200 119.200 210.500 125.800 ;
        RECT 215.000 125.200 215.300 145.800 ;
        RECT 219.800 144.800 220.200 145.200 ;
        RECT 220.600 145.100 221.000 147.900 ;
        RECT 219.800 144.200 220.100 144.800 ;
        RECT 219.800 143.800 220.200 144.200 ;
        RECT 222.200 143.100 222.600 148.900 ;
        RECT 224.600 147.200 224.900 153.800 ;
        RECT 225.400 153.100 225.800 155.900 ;
        RECT 226.200 155.800 226.600 156.200 ;
        RECT 227.800 155.200 228.100 164.800 ;
        RECT 229.400 161.800 229.800 162.200 ;
        RECT 227.800 154.800 228.200 155.200 ;
        RECT 227.000 153.800 227.400 154.200 ;
        RECT 226.200 152.800 226.600 153.200 ;
        RECT 225.400 151.800 225.800 152.200 ;
        RECT 223.000 146.800 223.400 147.200 ;
        RECT 223.800 146.800 224.200 147.200 ;
        RECT 224.600 146.800 225.000 147.200 ;
        RECT 223.000 146.300 223.300 146.800 ;
        RECT 223.000 145.900 223.400 146.300 ;
        RECT 223.000 143.800 223.400 144.200 ;
        RECT 215.800 132.100 216.200 137.900 ;
        RECT 217.400 133.100 217.800 135.900 ;
        RECT 218.200 133.100 218.600 135.900 ;
        RECT 219.800 132.100 220.200 137.900 ;
        RECT 221.400 134.800 221.800 135.200 ;
        RECT 221.400 133.200 221.700 134.800 ;
        RECT 221.400 132.800 221.800 133.200 ;
        RECT 218.200 129.100 218.600 129.200 ;
        RECT 219.000 129.100 219.400 129.200 ;
        RECT 218.200 128.800 219.400 129.100 ;
        RECT 217.400 127.100 217.800 127.200 ;
        RECT 218.200 127.100 218.600 127.200 ;
        RECT 217.400 126.800 218.600 127.100 ;
        RECT 216.600 126.100 217.000 126.200 ;
        RECT 217.400 126.100 217.800 126.200 ;
        RECT 216.600 125.800 217.800 126.100 ;
        RECT 218.200 125.800 218.600 126.200 ;
        RECT 218.200 125.200 218.500 125.800 ;
        RECT 215.000 125.100 215.400 125.200 ;
        RECT 215.800 125.100 216.200 125.200 ;
        RECT 215.000 124.800 216.200 125.100 ;
        RECT 218.200 124.800 218.600 125.200 ;
        RECT 210.200 118.800 210.600 119.200 ;
        RECT 209.400 116.100 209.800 116.200 ;
        RECT 210.200 116.100 210.600 116.200 ;
        RECT 209.400 115.800 210.600 116.100 ;
        RECT 210.200 114.800 210.600 115.200 ;
        RECT 207.800 113.800 208.200 114.200 ;
        RECT 208.600 113.800 209.000 114.200 ;
        RECT 208.600 111.800 209.000 112.200 ;
        RECT 207.000 108.800 207.400 109.200 ;
        RECT 207.000 107.100 207.400 107.200 ;
        RECT 207.800 107.100 208.200 107.200 ;
        RECT 207.000 106.800 208.200 107.100 ;
        RECT 204.600 105.800 205.000 106.200 ;
        RECT 207.800 105.800 208.200 106.200 ;
        RECT 201.400 97.800 201.800 98.200 ;
        RECT 198.200 96.800 198.600 97.200 ;
        RECT 195.800 96.100 196.200 96.200 ;
        RECT 196.600 96.100 197.000 96.200 ;
        RECT 195.800 95.800 197.000 96.100 ;
        RECT 198.200 95.200 198.500 96.800 ;
        RECT 191.800 94.800 192.200 95.200 ;
        RECT 194.200 94.800 194.600 95.200 ;
        RECT 195.000 95.100 195.400 95.200 ;
        RECT 195.800 95.100 196.200 95.200 ;
        RECT 195.000 94.800 196.200 95.100 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 199.000 95.100 199.400 95.200 ;
        RECT 199.800 95.100 200.200 95.200 ;
        RECT 199.000 94.800 200.200 95.100 ;
        RECT 191.800 93.800 192.200 94.200 ;
        RECT 191.800 92.200 192.100 93.800 ;
        RECT 191.800 91.800 192.200 92.200 ;
        RECT 192.600 88.800 193.000 89.200 ;
        RECT 192.600 87.200 192.900 88.800 ;
        RECT 197.400 87.800 197.800 88.200 ;
        RECT 197.400 87.200 197.700 87.800 ;
        RECT 199.000 87.200 199.300 94.800 ;
        RECT 199.800 94.100 200.200 94.200 ;
        RECT 200.600 94.100 201.000 94.200 ;
        RECT 199.800 93.800 201.000 94.100 ;
        RECT 192.600 86.800 193.000 87.200 ;
        RECT 195.800 86.800 196.200 87.200 ;
        RECT 197.400 86.800 197.800 87.200 ;
        RECT 199.000 86.800 199.400 87.200 ;
        RECT 195.800 86.200 196.100 86.800 ;
        RECT 189.400 85.800 189.800 86.200 ;
        RECT 190.200 85.800 190.600 86.200 ;
        RECT 192.600 85.800 193.000 86.200 ;
        RECT 193.400 85.800 193.800 86.200 ;
        RECT 195.800 85.800 196.200 86.200 ;
        RECT 187.800 81.800 188.200 82.200 ;
        RECT 188.600 81.800 189.000 82.200 ;
        RECT 187.000 78.800 187.400 79.200 ;
        RECT 181.400 75.800 181.800 76.200 ;
        RECT 182.200 75.800 182.600 76.200 ;
        RECT 183.000 75.800 183.400 76.200 ;
        RECT 184.600 75.800 185.000 76.200 ;
        RECT 186.200 76.100 186.600 76.200 ;
        RECT 185.400 75.800 186.600 76.100 ;
        RECT 181.400 75.200 181.700 75.800 ;
        RECT 182.200 75.200 182.500 75.800 ;
        RECT 183.000 75.200 183.300 75.800 ;
        RECT 185.400 75.200 185.700 75.800 ;
        RECT 188.600 75.200 188.900 81.800 ;
        RECT 192.600 78.100 192.900 85.800 ;
        RECT 193.400 85.200 193.700 85.800 ;
        RECT 193.400 84.800 193.800 85.200 ;
        RECT 195.800 84.800 196.200 85.200 ;
        RECT 195.800 84.200 196.100 84.800 ;
        RECT 195.800 83.800 196.200 84.200 ;
        RECT 193.400 82.800 193.800 83.200 ;
        RECT 200.600 83.100 201.000 88.900 ;
        RECT 201.400 87.200 201.700 97.800 ;
        RECT 202.200 96.100 202.600 96.200 ;
        RECT 203.000 96.100 203.400 96.200 ;
        RECT 202.200 95.800 203.400 96.100 ;
        RECT 203.800 95.800 204.200 96.200 ;
        RECT 203.800 95.200 204.100 95.800 ;
        RECT 204.600 95.200 204.900 105.800 ;
        RECT 207.800 105.200 208.100 105.800 ;
        RECT 207.800 104.800 208.200 105.200 ;
        RECT 208.600 105.100 208.900 111.800 ;
        RECT 210.200 109.200 210.500 114.800 ;
        RECT 212.600 112.100 213.000 117.900 ;
        RECT 216.600 115.800 217.000 116.200 ;
        RECT 216.600 115.100 216.900 115.800 ;
        RECT 216.600 114.700 217.000 115.100 ;
        RECT 216.600 112.800 217.000 113.200 ;
        RECT 210.200 108.800 210.600 109.200 ;
        RECT 209.400 106.100 209.800 106.200 ;
        RECT 210.200 106.100 210.600 106.200 ;
        RECT 209.400 105.800 210.600 106.100 ;
        RECT 209.400 105.100 209.800 105.200 ;
        RECT 208.600 104.800 209.800 105.100 ;
        RECT 212.600 103.100 213.000 108.900 ;
        RECT 216.600 108.200 216.900 112.800 ;
        RECT 217.400 112.100 217.800 117.900 ;
        RECT 216.600 107.800 217.000 108.200 ;
        RECT 214.200 106.100 214.600 106.200 ;
        RECT 215.000 106.100 215.400 106.200 ;
        RECT 214.200 105.800 215.400 106.100 ;
        RECT 217.400 103.100 217.800 108.900 ;
        RECT 202.200 94.800 202.600 95.200 ;
        RECT 203.800 94.800 204.200 95.200 ;
        RECT 204.600 94.800 205.000 95.200 ;
        RECT 202.200 94.200 202.500 94.800 ;
        RECT 204.600 94.200 204.900 94.800 ;
        RECT 202.200 93.800 202.600 94.200 ;
        RECT 204.600 93.800 205.000 94.200 ;
        RECT 205.400 93.100 205.800 95.900 ;
        RECT 206.200 93.800 206.600 94.200 ;
        RECT 202.200 88.800 202.600 89.200 ;
        RECT 201.400 86.800 201.800 87.200 ;
        RECT 193.400 79.200 193.700 82.800 ;
        RECT 193.400 78.800 193.800 79.200 ;
        RECT 199.800 78.800 200.200 79.200 ;
        RECT 192.600 77.800 193.700 78.100 ;
        RECT 191.800 76.800 192.200 77.200 ;
        RECT 191.800 76.200 192.100 76.800 ;
        RECT 191.800 75.800 192.200 76.200 ;
        RECT 193.400 75.200 193.700 77.800 ;
        RECT 195.800 76.800 196.200 77.200 ;
        RECT 174.200 74.800 174.600 75.200 ;
        RECT 175.000 74.800 175.400 75.200 ;
        RECT 176.600 74.800 177.000 75.200 ;
        RECT 181.400 74.800 181.800 75.200 ;
        RECT 182.200 74.800 182.600 75.200 ;
        RECT 183.000 74.800 183.400 75.200 ;
        RECT 183.800 74.800 184.200 75.200 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 186.200 75.100 186.600 75.200 ;
        RECT 187.000 75.100 187.400 75.200 ;
        RECT 186.200 74.800 187.400 75.100 ;
        RECT 188.600 74.800 189.000 75.200 ;
        RECT 193.400 74.800 193.800 75.200 ;
        RECT 175.000 74.200 175.300 74.800 ;
        RECT 175.000 73.800 175.400 74.200 ;
        RECT 175.800 73.800 176.200 74.200 ;
        RECT 175.800 73.200 176.100 73.800 ;
        RECT 175.800 72.800 176.200 73.200 ;
        RECT 176.600 71.200 176.900 74.800 ;
        RECT 183.000 73.800 183.400 74.200 ;
        RECT 183.000 73.200 183.300 73.800 ;
        RECT 183.000 72.800 183.400 73.200 ;
        RECT 177.400 71.800 177.800 72.200 ;
        RECT 176.600 70.800 177.000 71.200 ;
        RECT 160.600 69.800 161.700 70.100 ;
        RECT 168.600 69.800 169.000 70.200 ;
        RECT 171.000 69.800 171.400 70.200 ;
        RECT 171.800 69.800 172.200 70.200 ;
        RECT 159.000 68.800 159.400 69.200 ;
        RECT 160.600 68.800 161.000 69.200 ;
        RECT 159.000 67.200 159.300 68.800 ;
        RECT 160.600 68.200 160.900 68.800 ;
        RECT 160.600 67.800 161.000 68.200 ;
        RECT 155.800 67.100 156.200 67.200 ;
        RECT 156.600 67.100 157.000 67.200 ;
        RECT 155.800 66.800 157.000 67.100 ;
        RECT 159.000 66.800 159.400 67.200 ;
        RECT 161.400 66.200 161.700 69.800 ;
        RECT 164.600 69.100 165.000 69.200 ;
        RECT 165.400 69.100 165.800 69.200 ;
        RECT 164.600 68.800 165.800 69.100 ;
        RECT 168.600 68.800 169.000 69.200 ;
        RECT 169.400 69.100 169.800 69.200 ;
        RECT 170.200 69.100 170.600 69.200 ;
        RECT 169.400 68.800 170.600 69.100 ;
        RECT 168.600 67.200 168.900 68.800 ;
        RECT 162.200 66.800 162.600 67.200 ;
        RECT 167.000 67.100 167.400 67.200 ;
        RECT 167.800 67.100 168.200 67.200 ;
        RECT 167.000 66.800 168.200 67.100 ;
        RECT 168.600 66.800 169.000 67.200 ;
        RECT 147.800 65.800 148.200 66.200 ;
        RECT 149.400 66.100 149.800 66.200 ;
        RECT 150.200 66.100 150.600 66.200 ;
        RECT 149.400 65.800 150.600 66.100 ;
        RECT 151.000 65.800 151.400 66.200 ;
        RECT 153.400 65.800 153.800 66.200 ;
        RECT 155.000 65.800 155.400 66.200 ;
        RECT 161.400 65.800 161.800 66.200 ;
        RECT 147.800 59.200 148.100 65.800 ;
        RECT 148.600 65.100 149.000 65.200 ;
        RECT 149.400 65.100 149.800 65.200 ;
        RECT 148.600 64.800 149.800 65.100 ;
        RECT 162.200 62.200 162.500 66.800 ;
        RECT 166.200 65.800 166.600 66.200 ;
        RECT 167.800 65.800 168.200 66.200 ;
        RECT 163.800 64.800 164.200 65.200 ;
        RECT 164.600 65.100 165.000 65.200 ;
        RECT 165.400 65.100 165.800 65.200 ;
        RECT 164.600 64.800 165.800 65.100 ;
        RECT 163.800 64.200 164.100 64.800 ;
        RECT 163.800 63.800 164.200 64.200 ;
        RECT 163.000 62.800 163.400 63.200 ;
        RECT 151.800 61.800 152.200 62.200 ;
        RECT 160.600 61.800 161.000 62.200 ;
        RECT 162.200 61.800 162.600 62.200 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 147.800 58.800 148.200 59.200 ;
        RECT 151.800 57.200 152.100 61.800 ;
        RECT 160.600 60.200 160.900 61.800 ;
        RECT 155.000 59.800 155.400 60.200 ;
        RECT 160.600 59.800 161.000 60.200 ;
        RECT 151.800 56.800 152.200 57.200 ;
        RECT 146.200 55.800 146.600 56.200 ;
        RECT 149.400 55.800 149.800 56.200 ;
        RECT 144.600 53.800 145.000 54.200 ;
        RECT 144.600 53.200 144.900 53.800 ;
        RECT 144.600 52.800 145.000 53.200 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 145.400 52.200 145.700 52.800 ;
        RECT 143.800 51.800 144.200 52.200 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 143.800 49.200 144.100 51.800 ;
        RECT 146.200 49.200 146.500 55.800 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 148.600 54.800 149.000 55.200 ;
        RECT 147.800 54.200 148.100 54.800 ;
        RECT 148.600 54.200 148.900 54.800 ;
        RECT 147.800 53.800 148.200 54.200 ;
        RECT 148.600 53.800 149.000 54.200 ;
        RECT 149.400 53.100 149.700 55.800 ;
        RECT 148.600 52.800 149.700 53.100 ;
        RECT 151.000 53.800 151.400 54.200 ;
        RECT 147.800 49.800 148.200 50.200 ;
        RECT 143.800 48.800 144.200 49.200 ;
        RECT 146.200 48.800 146.600 49.200 ;
        RECT 147.000 47.800 147.400 48.200 ;
        RECT 147.000 47.200 147.300 47.800 ;
        RECT 147.800 47.200 148.100 49.800 ;
        RECT 135.800 46.800 136.200 47.200 ;
        RECT 140.600 46.800 141.000 47.200 ;
        RECT 143.000 46.800 143.400 47.200 ;
        RECT 147.000 46.800 147.400 47.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 135.800 44.200 136.100 46.800 ;
        RECT 137.400 45.800 137.800 46.200 ;
        RECT 139.000 46.100 139.400 46.200 ;
        RECT 139.800 46.100 140.200 46.200 ;
        RECT 139.000 45.800 140.200 46.100 ;
        RECT 137.400 45.200 137.700 45.800 ;
        RECT 137.400 44.800 137.800 45.200 ;
        RECT 135.800 43.800 136.200 44.200 ;
        RECT 143.000 37.200 143.300 46.800 ;
        RECT 148.600 46.200 148.900 52.800 ;
        RECT 150.200 51.800 150.600 52.200 ;
        RECT 149.400 46.800 149.800 47.200 ;
        RECT 149.400 46.200 149.700 46.800 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 149.400 45.800 149.800 46.200 ;
        RECT 144.600 45.100 145.000 45.200 ;
        RECT 145.400 45.100 145.800 45.200 ;
        RECT 144.600 44.800 145.800 45.100 ;
        RECT 148.600 42.200 148.900 45.800 ;
        RECT 150.200 45.200 150.500 51.800 ;
        RECT 151.000 49.200 151.300 53.800 ;
        RECT 151.800 53.100 152.200 55.900 ;
        RECT 153.400 52.100 153.800 57.900 ;
        RECT 155.000 55.200 155.300 59.800 ;
        RECT 160.600 59.100 161.000 59.200 ;
        RECT 161.400 59.100 161.800 59.200 ;
        RECT 160.600 58.800 161.800 59.100 ;
        RECT 155.000 54.800 155.400 55.200 ;
        RECT 157.400 53.800 157.800 54.200 ;
        RECT 157.400 53.200 157.700 53.800 ;
        RECT 154.200 52.800 154.600 53.200 ;
        RECT 157.400 52.800 157.800 53.200 ;
        RECT 151.000 48.800 151.400 49.200 ;
        RECT 150.200 44.800 150.600 45.200 ;
        RECT 151.000 45.100 151.400 47.900 ;
        RECT 151.800 46.800 152.200 47.200 ;
        RECT 151.800 43.200 152.100 46.800 ;
        RECT 150.200 42.800 150.600 43.200 ;
        RECT 151.800 42.800 152.200 43.200 ;
        RECT 152.600 43.100 153.000 48.900 ;
        RECT 154.200 47.200 154.500 52.800 ;
        RECT 158.200 52.100 158.600 57.900 ;
        RECT 161.400 57.800 161.800 58.200 ;
        RECT 161.400 54.200 161.700 57.800 ;
        RECT 163.000 56.200 163.300 62.800 ;
        RECT 166.200 59.200 166.500 65.800 ;
        RECT 167.800 64.200 168.100 65.800 ;
        RECT 171.000 65.200 171.300 69.800 ;
        RECT 171.800 66.100 172.100 69.800 ;
        RECT 172.600 67.100 173.000 67.200 ;
        RECT 173.400 67.100 173.800 67.200 ;
        RECT 172.600 66.800 173.800 67.100 ;
        RECT 172.600 66.100 173.000 66.200 ;
        RECT 171.800 65.800 173.000 66.100 ;
        RECT 171.000 64.800 171.400 65.200 ;
        RECT 174.200 65.100 174.600 67.900 ;
        RECT 167.800 63.800 168.200 64.200 ;
        RECT 175.800 63.100 176.200 68.900 ;
        RECT 177.400 67.200 177.700 71.800 ;
        RECT 183.000 69.800 183.400 70.200 ;
        RECT 183.000 69.200 183.300 69.800 ;
        RECT 183.800 69.200 184.100 74.800 ;
        RECT 188.600 70.800 189.000 71.200 ;
        RECT 176.600 66.800 177.000 67.200 ;
        RECT 177.400 66.800 177.800 67.200 ;
        RECT 176.600 66.300 176.900 66.800 ;
        RECT 176.600 65.900 177.000 66.300 ;
        RECT 166.200 58.800 166.600 59.200 ;
        RECT 165.400 57.100 165.800 57.200 ;
        RECT 166.200 57.100 166.600 57.200 ;
        RECT 165.400 56.800 166.600 57.100 ;
        RECT 163.000 55.800 163.400 56.200 ;
        RECT 163.000 55.200 163.300 55.800 ;
        RECT 163.000 54.800 163.400 55.200 ;
        RECT 164.600 55.100 165.000 55.200 ;
        RECT 165.400 55.100 165.800 55.200 ;
        RECT 164.600 54.800 165.800 55.100 ;
        RECT 167.000 54.800 167.400 55.200 ;
        RECT 167.800 54.800 168.200 55.200 ;
        RECT 170.200 54.800 170.600 55.200 ;
        RECT 161.400 53.800 161.800 54.200 ;
        RECT 166.200 53.800 166.600 54.200 ;
        RECT 160.600 51.800 161.000 52.200 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 159.800 49.100 160.200 49.200 ;
        RECT 154.200 46.800 154.600 47.200 ;
        RECT 153.400 45.900 153.800 46.300 ;
        RECT 153.400 45.200 153.700 45.900 ;
        RECT 153.400 44.800 153.800 45.200 ;
        RECT 153.400 42.800 153.800 43.200 ;
        RECT 157.400 43.100 157.800 48.900 ;
        RECT 159.000 48.800 160.200 49.100 ;
        RECT 160.600 46.200 160.900 51.800 ;
        RECT 166.200 50.200 166.500 53.800 ;
        RECT 167.000 53.200 167.300 54.800 ;
        RECT 167.000 52.800 167.400 53.200 ;
        RECT 163.000 49.800 163.400 50.200 ;
        RECT 165.400 49.800 165.800 50.200 ;
        RECT 166.200 49.800 166.600 50.200 ;
        RECT 163.000 47.200 163.300 49.800 ;
        RECT 163.000 46.800 163.400 47.200 ;
        RECT 160.600 45.800 161.000 46.200 ;
        RECT 163.800 45.800 164.200 46.200 ;
        RECT 163.800 45.200 164.100 45.800 ;
        RECT 163.800 44.800 164.200 45.200 ;
        RECT 148.600 41.800 149.000 42.200 ;
        RECT 135.000 36.800 135.400 37.200 ;
        RECT 141.400 37.100 141.800 37.200 ;
        RECT 142.200 37.100 142.600 37.200 ;
        RECT 141.400 36.800 142.600 37.100 ;
        RECT 143.000 36.800 143.400 37.200 ;
        RECT 135.000 34.200 135.300 36.800 ;
        RECT 136.600 35.800 137.000 36.200 ;
        RECT 139.000 36.100 139.400 36.200 ;
        RECT 139.800 36.100 140.200 36.200 ;
        RECT 139.000 35.800 140.200 36.100 ;
        RECT 136.600 35.200 136.900 35.800 ;
        RECT 136.600 34.800 137.000 35.200 ;
        RECT 139.000 35.100 139.400 35.200 ;
        RECT 139.800 35.100 140.200 35.200 ;
        RECT 139.000 34.800 140.200 35.100 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 135.000 33.800 135.400 34.200 ;
        RECT 139.800 33.800 140.200 34.200 ;
        RECT 133.400 32.800 133.800 33.200 ;
        RECT 129.400 28.800 129.800 29.200 ;
        RECT 134.200 27.200 134.500 33.800 ;
        RECT 139.800 28.200 140.100 33.800 ;
        RECT 143.000 31.200 143.300 36.800 ;
        RECT 144.600 32.100 145.000 37.900 ;
        RECT 147.800 35.800 148.200 36.200 ;
        RECT 147.800 35.200 148.100 35.800 ;
        RECT 145.400 34.800 145.800 35.200 ;
        RECT 147.800 34.800 148.200 35.200 ;
        RECT 145.400 34.200 145.700 34.800 ;
        RECT 145.400 33.800 145.800 34.200 ;
        RECT 146.200 32.800 146.600 33.200 ;
        RECT 143.000 30.800 143.400 31.200 ;
        RECT 143.800 28.800 144.200 29.200 ;
        RECT 139.800 27.800 140.200 28.200 ;
        RECT 143.000 27.800 143.400 28.200 ;
        RECT 127.000 26.800 127.400 27.200 ;
        RECT 134.200 26.800 134.600 27.200 ;
        RECT 134.200 25.200 134.500 26.800 ;
        RECT 134.200 24.800 134.600 25.200 ;
        RECT 131.000 22.800 131.400 23.200 ;
        RECT 140.600 22.800 141.000 23.200 ;
        RECT 126.200 18.800 126.600 19.200 ;
        RECT 127.800 18.800 128.200 19.200 ;
        RECT 127.800 18.200 128.100 18.800 ;
        RECT 127.800 17.800 128.200 18.200 ;
        RECT 131.000 16.200 131.300 22.800 ;
        RECT 140.600 22.200 140.900 22.800 ;
        RECT 134.200 21.800 134.600 22.200 ;
        RECT 137.400 21.800 137.800 22.200 ;
        RECT 140.600 21.800 141.000 22.200 ;
        RECT 134.200 19.200 134.500 21.800 ;
        RECT 134.200 18.800 134.600 19.200 ;
        RECT 123.000 16.100 123.400 16.200 ;
        RECT 123.800 16.100 124.200 16.200 ;
        RECT 123.000 15.800 124.200 16.100 ;
        RECT 126.200 15.800 126.600 16.200 ;
        RECT 131.000 15.800 131.400 16.200 ;
        RECT 135.800 15.800 136.200 16.200 ;
        RECT 126.200 15.200 126.500 15.800 ;
        RECT 126.200 14.800 126.600 15.200 ;
        RECT 125.400 13.800 125.800 14.200 ;
        RECT 128.600 14.100 129.000 14.200 ;
        RECT 129.400 14.100 129.800 14.200 ;
        RECT 128.600 13.800 129.800 14.100 ;
        RECT 123.000 11.800 123.400 12.200 ;
        RECT 122.200 7.800 122.600 8.200 ;
        RECT 123.000 6.200 123.300 11.800 ;
        RECT 125.400 11.200 125.700 13.800 ;
        RECT 127.800 11.800 128.200 12.200 ;
        RECT 130.200 11.800 130.600 12.200 ;
        RECT 125.400 10.800 125.800 11.200 ;
        RECT 127.800 10.200 128.100 11.800 ;
        RECT 128.600 10.800 129.000 11.200 ;
        RECT 127.800 9.800 128.200 10.200 ;
        RECT 128.600 9.200 128.900 10.800 ;
        RECT 123.800 7.800 124.200 8.200 ;
        RECT 123.800 7.200 124.100 7.800 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 123.000 5.800 123.400 6.200 ;
        RECT 126.200 3.100 126.600 8.900 ;
        RECT 128.600 8.800 129.000 9.200 ;
        RECT 129.400 6.800 129.800 7.200 ;
        RECT 129.400 6.200 129.700 6.800 ;
        RECT 129.400 5.800 129.800 6.200 ;
        RECT 129.400 5.100 129.800 5.200 ;
        RECT 130.200 5.100 130.500 11.800 ;
        RECT 131.000 6.200 131.300 15.800 ;
        RECT 135.800 15.200 136.100 15.800 ;
        RECT 132.600 14.800 133.000 15.200 ;
        RECT 135.000 14.800 135.400 15.200 ;
        RECT 135.800 14.800 136.200 15.200 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 132.600 11.200 132.900 14.800 ;
        RECT 135.000 14.200 135.300 14.800 ;
        RECT 136.600 14.200 136.900 14.800 ;
        RECT 135.000 13.800 135.400 14.200 ;
        RECT 136.600 13.800 137.000 14.200 ;
        RECT 132.600 10.800 133.000 11.200 ;
        RECT 135.000 10.200 135.300 13.800 ;
        RECT 132.600 9.800 133.000 10.200 ;
        RECT 135.000 9.800 135.400 10.200 ;
        RECT 132.600 9.200 132.900 9.800 ;
        RECT 131.800 8.800 132.200 9.200 ;
        RECT 132.600 8.800 133.000 9.200 ;
        RECT 131.800 7.200 132.100 8.800 ;
        RECT 131.800 6.800 132.200 7.200 ;
        RECT 131.000 5.800 131.400 6.200 ;
        RECT 129.400 4.800 130.500 5.100 ;
        RECT 135.000 3.100 135.400 8.900 ;
        RECT 137.400 8.200 137.700 21.800 ;
        RECT 138.200 15.800 138.600 16.200 ;
        RECT 142.200 15.800 142.600 16.200 ;
        RECT 138.200 15.200 138.500 15.800 ;
        RECT 142.200 15.200 142.500 15.800 ;
        RECT 138.200 14.800 138.600 15.200 ;
        RECT 141.400 15.100 141.800 15.200 ;
        RECT 142.200 15.100 142.600 15.200 ;
        RECT 141.400 14.800 142.600 15.100 ;
        RECT 143.000 14.200 143.300 27.800 ;
        RECT 143.800 27.200 144.100 28.800 ;
        RECT 143.800 26.800 144.200 27.200 ;
        RECT 145.400 25.800 145.800 26.200 ;
        RECT 145.400 25.200 145.700 25.800 ;
        RECT 145.400 24.800 145.800 25.200 ;
        RECT 145.400 24.200 145.700 24.800 ;
        RECT 145.400 23.800 145.800 24.200 ;
        RECT 146.200 19.200 146.500 32.800 ;
        RECT 149.400 32.100 149.800 37.900 ;
        RECT 150.200 34.200 150.500 42.800 ;
        RECT 153.400 39.200 153.700 42.800 ;
        RECT 157.400 41.800 157.800 42.200 ;
        RECT 155.000 39.800 155.400 40.200 ;
        RECT 152.600 38.800 153.000 39.200 ;
        RECT 153.400 38.800 153.800 39.200 ;
        RECT 150.200 33.800 150.600 34.200 ;
        RECT 151.000 33.100 151.400 35.900 ;
        RECT 152.600 35.200 152.900 38.800 ;
        RECT 154.200 36.800 154.600 37.200 ;
        RECT 154.200 35.200 154.500 36.800 ;
        RECT 152.600 34.800 153.000 35.200 ;
        RECT 154.200 34.800 154.600 35.200 ;
        RECT 155.000 34.200 155.300 39.800 ;
        RECT 157.400 39.200 157.700 41.800 ;
        RECT 157.400 38.800 157.800 39.200 ;
        RECT 160.600 37.800 161.000 38.200 ;
        RECT 159.800 35.800 160.200 36.200 ;
        RECT 155.800 34.800 156.200 35.200 ;
        RECT 159.000 34.800 159.400 35.200 ;
        RECT 151.800 34.100 152.200 34.200 ;
        RECT 152.600 34.100 153.000 34.200 ;
        RECT 151.800 33.800 153.000 34.100 ;
        RECT 155.000 33.800 155.400 34.200 ;
        RECT 155.800 30.200 156.100 34.800 ;
        RECT 159.000 33.200 159.300 34.800 ;
        RECT 159.000 32.800 159.400 33.200 ;
        RECT 155.800 29.800 156.200 30.200 ;
        RECT 157.400 29.800 157.800 30.200 ;
        RECT 148.600 29.100 149.000 29.200 ;
        RECT 149.400 29.100 149.800 29.200 ;
        RECT 148.600 28.800 149.800 29.100 ;
        RECT 148.600 26.800 149.000 27.200 ;
        RECT 147.000 26.100 147.400 26.200 ;
        RECT 147.800 26.100 148.200 26.200 ;
        RECT 147.000 25.800 148.200 26.100 ;
        RECT 147.800 24.800 148.200 25.200 ;
        RECT 147.800 24.200 148.100 24.800 ;
        RECT 148.600 24.200 148.900 26.800 ;
        RECT 147.800 23.800 148.200 24.200 ;
        RECT 148.600 23.800 149.000 24.200 ;
        RECT 147.800 22.800 148.200 23.200 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 147.800 15.200 148.100 22.800 ;
        RECT 148.600 19.200 148.900 23.800 ;
        RECT 151.800 23.100 152.200 28.900 ;
        RECT 152.600 26.800 153.000 27.200 ;
        RECT 149.400 21.800 149.800 22.200 ;
        RECT 148.600 18.800 149.000 19.200 ;
        RECT 143.800 14.800 144.200 15.200 ;
        RECT 147.000 14.800 147.400 15.200 ;
        RECT 147.800 14.800 148.200 15.200 ;
        RECT 143.000 13.800 143.400 14.200 ;
        RECT 140.600 11.800 141.000 12.200 ;
        RECT 137.400 7.800 137.800 8.200 ;
        RECT 137.400 7.200 137.700 7.800 ;
        RECT 137.400 6.800 137.800 7.200 ;
        RECT 139.000 5.900 139.400 6.300 ;
        RECT 139.000 5.200 139.300 5.900 ;
        RECT 139.000 4.800 139.400 5.200 ;
        RECT 139.800 3.100 140.200 8.900 ;
        RECT 140.600 5.200 140.900 11.800 ;
        RECT 143.000 9.200 143.300 13.800 ;
        RECT 143.800 9.200 144.100 14.800 ;
        RECT 147.000 10.200 147.300 14.800 ;
        RECT 148.600 13.100 149.000 15.900 ;
        RECT 149.400 14.200 149.700 21.800 ;
        RECT 149.400 13.800 149.800 14.200 ;
        RECT 147.000 9.800 147.400 10.200 ;
        RECT 143.000 8.800 143.400 9.200 ;
        RECT 143.800 8.800 144.200 9.200 ;
        RECT 143.800 8.200 144.100 8.800 ;
        RECT 140.600 4.800 141.000 5.200 ;
        RECT 141.400 5.100 141.800 7.900 ;
        RECT 143.800 7.800 144.200 8.200 ;
        RECT 146.200 3.100 146.600 8.900 ;
        RECT 149.400 7.200 149.700 13.800 ;
        RECT 150.200 12.100 150.600 17.900 ;
        RECT 152.600 15.200 152.900 26.800 ;
        RECT 153.400 25.800 153.800 26.200 ;
        RECT 155.000 25.800 155.400 26.200 ;
        RECT 153.400 22.200 153.700 25.800 ;
        RECT 155.000 25.200 155.300 25.800 ;
        RECT 155.000 24.800 155.400 25.200 ;
        RECT 156.600 23.100 157.000 28.900 ;
        RECT 153.400 21.800 153.800 22.200 ;
        RECT 157.400 19.200 157.700 29.800 ;
        RECT 158.200 25.100 158.600 27.900 ;
        RECT 159.000 26.800 159.400 27.200 ;
        RECT 159.000 24.200 159.300 26.800 ;
        RECT 159.800 26.200 160.100 35.800 ;
        RECT 160.600 35.200 160.900 37.800 ;
        RECT 163.000 37.100 163.400 37.200 ;
        RECT 163.800 37.100 164.200 37.200 ;
        RECT 163.000 36.800 164.200 37.100 ;
        RECT 164.600 36.800 165.000 37.200 ;
        RECT 164.600 36.200 164.900 36.800 ;
        RECT 161.400 36.100 161.800 36.200 ;
        RECT 162.200 36.100 162.600 36.200 ;
        RECT 161.400 35.800 162.600 36.100 ;
        RECT 164.600 35.800 165.000 36.200 ;
        RECT 160.600 35.100 161.000 35.200 ;
        RECT 160.600 34.800 161.700 35.100 ;
        RECT 161.400 34.200 161.700 34.800 ;
        RECT 165.400 34.200 165.700 49.800 ;
        RECT 167.800 49.200 168.100 54.800 ;
        RECT 168.600 52.100 169.000 52.200 ;
        RECT 169.400 52.100 169.800 52.200 ;
        RECT 168.600 51.800 169.800 52.100 ;
        RECT 167.800 48.800 168.200 49.200 ;
        RECT 170.200 48.200 170.500 54.800 ;
        RECT 171.800 53.100 172.200 55.900 ;
        RECT 172.600 54.800 173.000 55.200 ;
        RECT 172.600 54.200 172.900 54.800 ;
        RECT 172.600 53.800 173.000 54.200 ;
        RECT 170.200 47.800 170.600 48.200 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 166.200 46.200 166.500 46.800 ;
        RECT 166.200 45.800 166.600 46.200 ;
        RECT 166.200 45.100 166.600 45.200 ;
        RECT 167.000 45.100 167.400 45.200 ;
        RECT 166.200 44.800 167.400 45.100 ;
        RECT 166.200 35.200 166.500 44.800 ;
        RECT 171.000 43.100 171.400 48.900 ;
        RECT 172.600 46.200 172.900 53.800 ;
        RECT 173.400 52.100 173.800 57.900 ;
        RECT 174.200 56.800 174.600 57.200 ;
        RECT 174.200 55.100 174.500 56.800 ;
        RECT 177.400 55.200 177.700 66.800 ;
        RECT 180.600 63.100 181.000 68.900 ;
        RECT 183.000 68.800 183.400 69.200 ;
        RECT 183.800 68.800 184.200 69.200 ;
        RECT 187.000 69.100 187.400 69.200 ;
        RECT 187.800 69.100 188.200 69.200 ;
        RECT 187.000 68.800 188.200 69.100 ;
        RECT 185.400 67.800 185.800 68.200 ;
        RECT 186.200 67.800 186.600 68.200 ;
        RECT 185.400 67.200 185.700 67.800 ;
        RECT 186.200 67.200 186.500 67.800 ;
        RECT 185.400 66.800 185.800 67.200 ;
        RECT 186.200 66.800 186.600 67.200 ;
        RECT 188.600 66.200 188.900 70.800 ;
        RECT 188.600 65.800 189.000 66.200 ;
        RECT 190.200 65.800 190.600 66.200 ;
        RECT 183.800 65.100 184.200 65.200 ;
        RECT 183.000 64.800 184.200 65.100 ;
        RECT 187.800 64.800 188.200 65.200 ;
        RECT 179.800 58.100 180.200 58.200 ;
        RECT 180.600 58.100 181.000 58.200 ;
        RECT 174.200 54.700 174.600 55.100 ;
        RECT 177.400 54.800 177.800 55.200 ;
        RECT 178.200 52.100 178.600 57.900 ;
        RECT 179.800 57.800 181.000 58.100 ;
        RECT 182.200 54.800 182.600 55.200 ;
        RECT 182.200 54.200 182.500 54.800 ;
        RECT 182.200 53.800 182.600 54.200 ;
        RECT 179.000 52.800 179.400 53.200 ;
        RECT 179.000 49.200 179.300 52.800 ;
        RECT 183.000 49.200 183.300 64.800 ;
        RECT 186.200 63.800 186.600 64.200 ;
        RECT 186.200 59.200 186.500 63.800 ;
        RECT 186.200 58.800 186.600 59.200 ;
        RECT 183.800 57.800 184.200 58.200 ;
        RECT 183.800 55.200 184.100 57.800 ;
        RECT 184.600 55.800 185.000 56.200 ;
        RECT 184.600 55.200 184.900 55.800 ;
        RECT 183.800 54.800 184.200 55.200 ;
        RECT 184.600 54.800 185.000 55.200 ;
        RECT 185.400 54.800 185.800 55.200 ;
        RECT 172.600 45.800 173.000 46.200 ;
        RECT 173.400 46.100 173.800 46.200 ;
        RECT 174.200 46.100 174.600 46.200 ;
        RECT 173.400 45.800 174.600 46.100 ;
        RECT 175.800 43.100 176.200 48.900 ;
        RECT 179.000 48.800 179.400 49.200 ;
        RECT 183.000 48.800 183.400 49.200 ;
        RECT 177.400 45.100 177.800 47.900 ;
        RECT 179.000 46.200 179.300 48.800 ;
        RECT 181.400 47.800 181.800 48.200 ;
        RECT 180.600 46.800 181.000 47.200 ;
        RECT 180.600 46.200 180.900 46.800 ;
        RECT 181.400 46.200 181.700 47.800 ;
        RECT 183.800 47.200 184.100 54.800 ;
        RECT 185.400 54.200 185.700 54.800 ;
        RECT 185.400 53.800 185.800 54.200 ;
        RECT 185.400 49.100 185.700 53.800 ;
        RECT 187.800 53.200 188.100 64.800 ;
        RECT 188.600 58.200 188.900 65.800 ;
        RECT 190.200 62.200 190.500 65.800 ;
        RECT 193.400 64.200 193.700 74.800 ;
        RECT 195.800 73.200 196.100 76.800 ;
        RECT 199.800 75.200 200.100 78.800 ;
        RECT 202.200 77.100 202.500 88.800 ;
        RECT 203.000 86.100 203.400 86.200 ;
        RECT 203.800 86.100 204.200 86.200 ;
        RECT 203.000 85.800 204.200 86.100 ;
        RECT 205.400 83.100 205.800 88.900 ;
        RECT 206.200 87.200 206.500 93.800 ;
        RECT 207.000 92.100 207.400 97.900 ;
        RECT 207.800 95.000 208.200 95.100 ;
        RECT 208.600 95.000 209.000 95.100 ;
        RECT 207.800 94.700 209.000 95.000 ;
        RECT 211.000 94.800 211.400 95.200 ;
        RECT 211.000 94.200 211.300 94.800 ;
        RECT 211.000 93.800 211.400 94.200 ;
        RECT 211.800 92.100 212.200 97.900 ;
        RECT 213.400 97.100 213.800 97.200 ;
        RECT 214.200 97.100 214.600 97.200 ;
        RECT 213.400 96.800 214.600 97.100 ;
        RECT 215.000 93.100 215.400 95.900 ;
        RECT 215.800 93.800 216.200 94.200 ;
        RECT 215.800 93.200 216.100 93.800 ;
        RECT 215.800 92.800 216.200 93.200 ;
        RECT 216.600 92.100 217.000 97.900 ;
        RECT 217.400 94.700 217.800 95.100 ;
        RECT 217.400 94.200 217.700 94.700 ;
        RECT 217.400 93.800 217.800 94.200 ;
        RECT 208.600 89.800 209.000 90.200 ;
        RECT 206.200 86.800 206.600 87.200 ;
        RECT 207.000 85.100 207.400 87.900 ;
        RECT 208.600 86.200 208.900 89.800 ;
        RECT 213.400 87.100 213.800 87.200 ;
        RECT 214.200 87.100 214.600 87.200 ;
        RECT 213.400 86.800 214.600 87.100 ;
        RECT 207.800 85.800 208.200 86.200 ;
        RECT 208.600 85.800 209.000 86.200 ;
        RECT 207.800 85.200 208.100 85.800 ;
        RECT 207.800 84.800 208.200 85.200 ;
        RECT 214.200 83.800 214.600 84.200 ;
        RECT 209.400 81.800 209.800 82.200 ;
        RECT 209.400 79.200 209.700 81.800 ;
        RECT 209.400 78.800 209.800 79.200 ;
        RECT 203.800 77.800 204.200 78.200 ;
        RECT 202.200 76.800 203.300 77.100 ;
        RECT 200.600 75.800 201.000 76.200 ;
        RECT 202.200 75.800 202.600 76.200 ;
        RECT 200.600 75.200 200.900 75.800 ;
        RECT 202.200 75.200 202.500 75.800 ;
        RECT 196.600 74.800 197.000 75.200 ;
        RECT 197.400 74.800 197.800 75.200 ;
        RECT 199.800 74.800 200.200 75.200 ;
        RECT 200.600 74.800 201.000 75.200 ;
        RECT 202.200 74.800 202.600 75.200 ;
        RECT 196.600 73.200 196.900 74.800 ;
        RECT 197.400 74.200 197.700 74.800 ;
        RECT 197.400 73.800 197.800 74.200 ;
        RECT 198.200 73.800 198.600 74.200 ;
        RECT 201.400 73.800 201.800 74.200 ;
        RECT 195.800 72.800 196.200 73.200 ;
        RECT 196.600 72.800 197.000 73.200 ;
        RECT 193.400 63.800 193.800 64.200 ;
        RECT 195.800 63.100 196.200 68.900 ;
        RECT 190.200 61.800 190.600 62.200 ;
        RECT 193.400 61.800 193.800 62.200 ;
        RECT 189.400 59.800 189.800 60.200 ;
        RECT 188.600 57.800 189.000 58.200 ;
        RECT 189.400 55.200 189.700 59.800 ;
        RECT 190.200 56.200 190.500 61.800 ;
        RECT 191.000 60.800 191.400 61.200 ;
        RECT 191.000 56.200 191.300 60.800 ;
        RECT 193.400 60.200 193.700 61.800 ;
        RECT 193.400 59.800 193.800 60.200 ;
        RECT 198.200 59.200 198.500 73.800 ;
        RECT 201.400 73.200 201.700 73.800 ;
        RECT 201.400 72.800 201.800 73.200 ;
        RECT 199.800 65.900 200.200 66.300 ;
        RECT 199.800 65.200 200.100 65.900 ;
        RECT 199.800 64.800 200.200 65.200 ;
        RECT 199.800 62.800 200.200 63.200 ;
        RECT 200.600 63.100 201.000 68.900 ;
        RECT 201.400 66.800 201.800 67.200 ;
        RECT 201.400 64.200 201.700 66.800 ;
        RECT 202.200 65.100 202.600 67.900 ;
        RECT 203.000 67.200 203.300 76.800 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 201.400 63.800 201.800 64.200 ;
        RECT 199.800 59.200 200.100 62.800 ;
        RECT 198.200 58.800 198.600 59.200 ;
        RECT 199.800 58.800 200.200 59.200 ;
        RECT 203.000 57.200 203.300 66.800 ;
        RECT 203.800 66.200 204.100 77.800 ;
        RECT 206.200 77.100 206.600 77.200 ;
        RECT 207.000 77.100 207.400 77.200 ;
        RECT 206.200 76.800 207.400 77.100 ;
        RECT 204.600 74.800 205.000 75.200 ;
        RECT 205.400 74.800 205.800 75.200 ;
        RECT 204.600 70.200 204.900 74.800 ;
        RECT 204.600 69.800 205.000 70.200 ;
        RECT 203.800 65.800 204.200 66.200 ;
        RECT 204.600 65.800 205.000 66.200 ;
        RECT 195.800 56.800 196.200 57.200 ;
        RECT 203.000 56.800 203.400 57.200 ;
        RECT 190.200 55.800 190.600 56.200 ;
        RECT 191.000 55.800 191.400 56.200 ;
        RECT 191.000 55.200 191.300 55.800 ;
        RECT 189.400 54.800 189.800 55.200 ;
        RECT 191.000 54.800 191.400 55.200 ;
        RECT 194.200 55.100 194.600 55.200 ;
        RECT 195.000 55.100 195.400 55.200 ;
        RECT 194.200 54.800 195.400 55.100 ;
        RECT 188.600 54.100 189.000 54.200 ;
        RECT 189.400 54.100 189.800 54.200 ;
        RECT 188.600 53.800 189.800 54.100 ;
        RECT 194.200 53.800 194.600 54.200 ;
        RECT 187.800 52.800 188.200 53.200 ;
        RECT 194.200 49.200 194.500 53.800 ;
        RECT 195.000 50.200 195.300 54.800 ;
        RECT 195.800 54.200 196.100 56.800 ;
        RECT 196.600 54.800 197.000 55.200 ;
        RECT 200.600 55.100 201.000 55.200 ;
        RECT 201.400 55.100 201.800 55.200 ;
        RECT 200.600 54.800 201.800 55.100 ;
        RECT 202.200 55.100 202.600 55.200 ;
        RECT 203.000 55.100 203.400 55.200 ;
        RECT 202.200 54.800 203.400 55.100 ;
        RECT 195.800 53.800 196.200 54.200 ;
        RECT 195.000 49.800 195.400 50.200 ;
        RECT 186.200 49.100 186.600 49.200 ;
        RECT 185.400 48.800 186.600 49.100 ;
        RECT 183.800 46.800 184.200 47.200 ;
        RECT 179.000 45.800 179.400 46.200 ;
        RECT 180.600 45.800 181.000 46.200 ;
        RECT 181.400 45.800 181.800 46.200 ;
        RECT 182.200 45.800 182.600 46.200 ;
        RECT 184.600 45.800 185.000 46.200 ;
        RECT 168.600 39.800 169.000 40.200 ;
        RECT 168.600 39.200 168.900 39.800 ;
        RECT 168.600 38.800 169.000 39.200 ;
        RECT 180.600 37.200 180.900 45.800 ;
        RECT 167.800 36.800 168.200 37.200 ;
        RECT 173.400 36.800 173.800 37.200 ;
        RECT 180.600 36.800 181.000 37.200 ;
        RECT 167.800 36.200 168.100 36.800 ;
        RECT 167.800 35.800 168.200 36.200 ;
        RECT 173.400 35.200 173.700 36.800 ;
        RECT 174.200 36.100 174.600 36.200 ;
        RECT 175.000 36.100 175.400 36.200 ;
        RECT 174.200 35.800 175.400 36.100 ;
        RECT 177.400 35.800 177.800 36.200 ;
        RECT 177.400 35.200 177.700 35.800 ;
        RECT 166.200 34.800 166.600 35.200 ;
        RECT 171.000 34.800 171.400 35.200 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 177.400 34.800 177.800 35.200 ;
        RECT 178.200 35.100 178.600 35.200 ;
        RECT 179.000 35.100 179.400 35.200 ;
        RECT 178.200 34.800 179.400 35.100 ;
        RECT 179.800 34.800 180.200 35.200 ;
        RECT 171.000 34.200 171.300 34.800 ;
        RECT 160.600 33.800 161.000 34.200 ;
        RECT 161.400 33.800 161.800 34.200 ;
        RECT 163.000 33.800 163.400 34.200 ;
        RECT 165.400 33.800 165.800 34.200 ;
        RECT 171.000 33.800 171.400 34.200 ;
        RECT 173.400 33.800 173.800 34.200 ;
        RECT 178.200 33.800 178.600 34.200 ;
        RECT 179.800 34.100 180.100 34.800 ;
        RECT 179.000 33.800 180.100 34.100 ;
        RECT 182.200 34.200 182.500 45.800 ;
        RECT 184.600 44.200 184.900 45.800 ;
        RECT 184.600 43.800 185.000 44.200 ;
        RECT 188.600 43.100 189.000 48.900 ;
        RECT 192.600 48.800 193.000 49.200 ;
        RECT 191.800 46.800 192.200 47.200 ;
        RECT 183.800 38.800 184.200 39.200 ;
        RECT 183.800 38.200 184.100 38.800 ;
        RECT 183.800 37.800 184.200 38.200 ;
        RECT 183.000 34.800 183.400 35.200 ;
        RECT 182.200 33.800 182.600 34.200 ;
        RECT 160.600 30.200 160.900 33.800 ;
        RECT 163.000 33.200 163.300 33.800 ;
        RECT 163.000 32.800 163.400 33.200 ;
        RECT 167.800 33.100 168.200 33.200 ;
        RECT 167.800 32.800 168.900 33.100 ;
        RECT 161.400 31.800 161.800 32.200 ;
        RECT 167.800 31.800 168.200 32.200 ;
        RECT 161.400 30.200 161.700 31.800 ;
        RECT 163.000 30.800 163.400 31.200 ;
        RECT 165.400 30.800 165.800 31.200 ;
        RECT 160.600 29.800 161.000 30.200 ;
        RECT 161.400 29.800 161.800 30.200 ;
        RECT 162.200 27.800 162.600 28.200 ;
        RECT 162.200 27.200 162.500 27.800 ;
        RECT 160.600 27.100 161.000 27.200 ;
        RECT 161.400 27.100 161.800 27.200 ;
        RECT 160.600 26.800 161.800 27.100 ;
        RECT 162.200 26.800 162.600 27.200 ;
        RECT 163.000 26.200 163.300 30.800 ;
        RECT 164.600 26.800 165.000 27.200 ;
        RECT 159.800 25.800 160.200 26.200 ;
        RECT 163.000 25.800 163.400 26.200 ;
        RECT 164.600 25.200 164.900 26.800 ;
        RECT 165.400 25.200 165.700 30.800 ;
        RECT 167.800 29.200 168.100 31.800 ;
        RECT 168.600 31.200 168.900 32.800 ;
        RECT 169.400 32.800 169.800 33.200 ;
        RECT 171.800 32.800 172.200 33.200 ;
        RECT 169.400 32.200 169.700 32.800 ;
        RECT 169.400 31.800 169.800 32.200 ;
        RECT 168.600 30.800 169.000 31.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 166.200 27.100 166.600 27.200 ;
        RECT 167.000 27.100 167.400 27.200 ;
        RECT 166.200 26.800 167.400 27.100 ;
        RECT 160.600 25.100 161.000 25.200 ;
        RECT 161.400 25.100 161.800 25.200 ;
        RECT 160.600 24.800 161.800 25.100 ;
        RECT 164.600 24.800 165.000 25.200 ;
        RECT 165.400 24.800 165.800 25.200 ;
        RECT 159.000 23.800 159.400 24.200 ;
        RECT 167.800 23.800 168.200 24.200 ;
        RECT 157.400 18.800 157.800 19.200 ;
        RECT 152.600 14.800 153.000 15.200 ;
        RECT 155.000 12.100 155.400 17.900 ;
        RECT 157.400 13.800 157.800 14.200 ;
        RECT 149.400 6.800 149.800 7.200 ;
        RECT 150.200 5.900 150.600 6.300 ;
        RECT 150.200 5.200 150.500 5.900 ;
        RECT 150.200 4.800 150.600 5.200 ;
        RECT 151.000 3.100 151.400 8.900 ;
        RECT 152.600 5.100 153.000 7.900 ;
        RECT 153.400 7.800 153.800 8.200 ;
        RECT 153.400 7.200 153.700 7.800 ;
        RECT 153.400 6.800 153.800 7.200 ;
        RECT 155.800 6.800 156.200 7.200 ;
        RECT 155.000 5.800 155.400 6.200 ;
        RECT 155.000 5.200 155.300 5.800 ;
        RECT 155.800 5.200 156.100 6.800 ;
        RECT 157.400 6.200 157.700 13.800 ;
        RECT 158.200 13.100 158.600 15.900 ;
        RECT 158.200 11.800 158.600 12.200 ;
        RECT 158.200 6.200 158.500 11.800 ;
        RECT 159.000 7.200 159.300 23.800 ;
        RECT 160.600 21.800 161.000 22.200 ;
        RECT 159.800 12.100 160.200 17.900 ;
        RECT 160.600 14.200 160.900 21.800 ;
        RECT 161.400 16.800 161.800 17.200 ;
        RECT 161.400 15.200 161.700 16.800 ;
        RECT 161.400 14.800 161.800 15.200 ;
        RECT 162.200 14.800 162.600 15.200 ;
        RECT 160.600 13.800 161.000 14.200 ;
        RECT 159.000 6.800 159.400 7.200 ;
        RECT 161.400 6.800 161.800 7.200 ;
        RECT 161.400 6.200 161.700 6.800 ;
        RECT 156.600 6.100 157.000 6.200 ;
        RECT 157.400 6.100 157.800 6.200 ;
        RECT 156.600 5.800 157.800 6.100 ;
        RECT 158.200 5.800 158.600 6.200 ;
        RECT 161.400 5.800 161.800 6.200 ;
        RECT 158.200 5.200 158.500 5.800 ;
        RECT 162.200 5.200 162.500 14.800 ;
        RECT 164.600 12.100 165.000 17.900 ;
        RECT 167.800 17.200 168.100 23.800 ;
        RECT 170.200 23.100 170.600 28.900 ;
        RECT 171.000 25.800 171.400 26.200 ;
        RECT 171.000 22.200 171.300 25.800 ;
        RECT 171.000 21.800 171.400 22.200 ;
        RECT 167.800 16.800 168.200 17.200 ;
        RECT 168.600 16.800 169.000 17.200 ;
        RECT 167.800 14.200 168.100 16.800 ;
        RECT 168.600 15.100 168.900 16.800 ;
        RECT 169.400 16.100 169.800 16.200 ;
        RECT 170.200 16.100 170.600 16.200 ;
        RECT 169.400 15.800 170.600 16.100 ;
        RECT 168.600 14.800 169.700 15.100 ;
        RECT 169.400 14.200 169.700 14.800 ;
        RECT 167.800 13.800 168.200 14.200 ;
        RECT 169.400 13.800 169.800 14.200 ;
        RECT 171.000 12.200 171.300 21.800 ;
        RECT 171.800 14.100 172.100 32.800 ;
        RECT 173.400 32.200 173.700 33.800 ;
        RECT 178.200 33.200 178.500 33.800 ;
        RECT 178.200 32.800 178.600 33.200 ;
        RECT 173.400 31.800 173.800 32.200 ;
        RECT 175.800 31.800 176.200 32.200 ;
        RECT 177.400 31.800 177.800 32.200 ;
        RECT 175.800 31.200 176.100 31.800 ;
        RECT 172.600 30.800 173.000 31.200 ;
        RECT 175.800 30.800 176.200 31.200 ;
        RECT 172.600 26.200 172.900 30.800 ;
        RECT 177.400 29.200 177.700 31.800 ;
        RECT 172.600 25.800 173.000 26.200 ;
        RECT 175.000 23.100 175.400 28.900 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 176.600 25.100 177.000 27.900 ;
        RECT 179.000 24.200 179.300 33.800 ;
        RECT 183.000 32.200 183.300 34.800 ;
        RECT 184.600 32.800 185.000 33.200 ;
        RECT 183.000 31.800 183.400 32.200 ;
        RECT 181.400 30.800 181.800 31.200 ;
        RECT 184.600 31.100 184.900 32.800 ;
        RECT 185.400 32.100 185.800 32.200 ;
        RECT 186.200 32.100 186.600 32.200 ;
        RECT 187.800 32.100 188.200 37.900 ;
        RECT 191.000 35.800 191.400 36.200 ;
        RECT 191.000 35.200 191.300 35.800 ;
        RECT 191.000 34.800 191.400 35.200 ;
        RECT 191.800 34.200 192.100 46.800 ;
        RECT 192.600 46.300 192.900 48.800 ;
        RECT 192.600 45.900 193.000 46.300 ;
        RECT 192.600 45.800 192.900 45.900 ;
        RECT 193.400 43.100 193.800 48.900 ;
        RECT 194.200 48.800 194.600 49.200 ;
        RECT 195.000 45.100 195.400 47.900 ;
        RECT 196.600 47.200 196.900 54.800 ;
        RECT 200.600 52.800 201.000 53.200 ;
        RECT 202.200 53.100 202.600 53.200 ;
        RECT 203.000 53.100 203.400 53.200 ;
        RECT 202.200 52.800 203.400 53.100 ;
        RECT 200.600 52.200 200.900 52.800 ;
        RECT 200.600 51.800 201.000 52.200 ;
        RECT 201.400 50.800 201.800 51.200 ;
        RECT 201.400 49.200 201.700 50.800 ;
        RECT 203.800 49.200 204.100 65.800 ;
        RECT 204.600 65.200 204.900 65.800 ;
        RECT 204.600 64.800 205.000 65.200 ;
        RECT 204.600 54.800 205.000 55.200 ;
        RECT 201.400 48.800 201.800 49.200 ;
        RECT 203.800 48.800 204.200 49.200 ;
        RECT 204.600 47.200 204.900 54.800 ;
        RECT 205.400 51.200 205.700 74.800 ;
        RECT 208.600 72.100 209.000 77.900 ;
        RECT 211.800 75.800 212.200 76.200 ;
        RECT 212.600 75.800 213.000 76.200 ;
        RECT 211.000 72.800 211.400 73.200 ;
        RECT 210.200 71.800 210.600 72.200 ;
        RECT 206.200 66.800 206.600 67.200 ;
        RECT 206.200 60.200 206.500 66.800 ;
        RECT 210.200 66.200 210.500 71.800 ;
        RECT 211.000 67.200 211.300 72.800 ;
        RECT 211.800 69.200 212.100 75.800 ;
        RECT 212.600 75.100 212.900 75.800 ;
        RECT 212.600 74.700 213.000 75.100 ;
        RECT 213.400 72.100 213.800 77.900 ;
        RECT 214.200 74.200 214.500 83.800 ;
        RECT 215.000 83.100 215.400 88.900 ;
        RECT 217.400 79.800 217.800 80.200 ;
        RECT 215.800 76.800 216.200 77.200 ;
        RECT 214.200 73.800 214.600 74.200 ;
        RECT 215.000 73.100 215.400 75.900 ;
        RECT 215.800 74.200 216.100 76.800 ;
        RECT 217.400 76.200 217.700 79.800 ;
        RECT 217.400 75.800 217.800 76.200 ;
        RECT 217.400 74.800 217.800 75.200 ;
        RECT 217.400 74.200 217.700 74.800 ;
        RECT 215.800 73.800 216.200 74.200 ;
        RECT 217.400 73.800 217.800 74.200 ;
        RECT 218.200 72.200 218.500 124.800 ;
        RECT 220.600 123.800 221.000 124.200 ;
        RECT 219.000 113.100 219.400 115.900 ;
        RECT 219.800 113.100 220.200 115.900 ;
        RECT 219.000 105.100 219.400 107.900 ;
        RECT 219.800 105.100 220.200 107.900 ;
        RECT 220.600 107.200 220.900 123.800 ;
        RECT 221.400 123.100 221.800 128.900 ;
        RECT 221.400 112.100 221.800 117.900 ;
        RECT 223.000 115.200 223.300 143.800 ;
        RECT 223.800 135.200 224.100 146.800 ;
        RECT 223.800 134.800 224.200 135.200 ;
        RECT 223.800 127.200 224.100 134.800 ;
        RECT 224.600 132.100 225.000 137.900 ;
        RECT 223.800 126.800 224.200 127.200 ;
        RECT 223.800 126.100 224.200 126.200 ;
        RECT 224.600 126.100 225.000 126.200 ;
        RECT 223.800 125.800 225.000 126.100 ;
        RECT 223.000 114.800 223.400 115.200 ;
        RECT 223.000 113.800 223.400 114.200 ;
        RECT 222.200 112.800 222.600 113.200 ;
        RECT 220.600 106.800 221.000 107.200 ;
        RECT 221.400 103.100 221.800 108.900 ;
        RECT 220.600 94.800 221.000 95.200 ;
        RECT 219.000 88.800 219.400 89.200 ;
        RECT 219.000 86.300 219.300 88.800 ;
        RECT 219.000 85.900 219.400 86.300 ;
        RECT 219.000 85.800 219.300 85.900 ;
        RECT 219.800 83.100 220.200 88.900 ;
        RECT 220.600 87.200 220.900 94.800 ;
        RECT 221.400 92.100 221.800 97.900 ;
        RECT 222.200 97.200 222.500 112.800 ;
        RECT 223.000 106.200 223.300 113.800 ;
        RECT 223.000 105.800 223.400 106.200 ;
        RECT 222.200 96.800 222.600 97.200 ;
        RECT 223.800 96.800 224.200 97.200 ;
        RECT 223.800 96.200 224.100 96.800 ;
        RECT 223.800 95.800 224.200 96.200 ;
        RECT 223.800 89.100 224.200 89.200 ;
        RECT 224.600 89.100 225.000 89.200 ;
        RECT 223.800 88.800 225.000 89.100 ;
        RECT 220.600 86.800 221.000 87.200 ;
        RECT 220.600 84.200 220.900 86.800 ;
        RECT 221.400 85.100 221.800 87.900 ;
        RECT 222.200 87.800 222.600 88.200 ;
        RECT 222.200 87.200 222.500 87.800 ;
        RECT 222.200 86.800 222.600 87.200 ;
        RECT 225.400 86.200 225.700 151.800 ;
        RECT 226.200 148.200 226.500 152.800 ;
        RECT 227.000 150.200 227.300 153.800 ;
        RECT 227.000 149.800 227.400 150.200 ;
        RECT 226.200 147.800 226.600 148.200 ;
        RECT 227.000 143.100 227.400 148.900 ;
        RECT 227.800 145.200 228.100 154.800 ;
        RECT 229.400 154.200 229.700 161.800 ;
        RECT 230.200 154.200 230.500 173.800 ;
        RECT 228.600 153.800 229.000 154.200 ;
        RECT 229.400 153.800 229.800 154.200 ;
        RECT 230.200 153.800 230.600 154.200 ;
        RECT 227.800 144.800 228.200 145.200 ;
        RECT 228.600 134.200 228.900 153.800 ;
        RECT 229.400 141.800 229.800 142.200 ;
        RECT 228.600 133.800 229.000 134.200 ;
        RECT 226.200 132.100 226.600 132.200 ;
        RECT 227.000 132.100 227.400 132.200 ;
        RECT 226.200 131.800 227.400 132.100 ;
        RECT 226.200 123.100 226.600 128.900 ;
        RECT 227.800 125.100 228.200 127.900 ;
        RECT 228.600 125.800 229.000 126.200 ;
        RECT 226.200 112.100 226.600 117.900 ;
        RECT 228.600 117.200 228.900 125.800 ;
        RECT 229.400 124.200 229.700 141.800 ;
        RECT 229.400 123.800 229.800 124.200 ;
        RECT 228.600 116.800 229.000 117.200 ;
        RECT 227.800 112.100 228.200 112.200 ;
        RECT 228.600 112.100 229.000 112.200 ;
        RECT 227.800 111.800 229.000 112.100 ;
        RECT 228.600 109.800 229.000 110.200 ;
        RECT 228.600 109.200 228.900 109.800 ;
        RECT 226.200 103.100 226.600 108.900 ;
        RECT 228.600 108.800 229.000 109.200 ;
        RECT 229.400 108.100 229.800 108.200 ;
        RECT 228.600 107.800 229.800 108.100 ;
        RECT 227.000 96.800 227.400 97.200 ;
        RECT 227.000 95.200 227.300 96.800 ;
        RECT 227.000 94.800 227.400 95.200 ;
        RECT 227.800 89.800 228.200 90.200 ;
        RECT 227.800 87.200 228.100 89.800 ;
        RECT 228.600 89.200 228.900 107.800 ;
        RECT 228.600 88.800 229.000 89.200 ;
        RECT 227.000 86.800 227.400 87.200 ;
        RECT 227.800 86.800 228.200 87.200 ;
        RECT 223.800 85.800 224.200 86.200 ;
        RECT 225.400 86.100 225.800 86.200 ;
        RECT 226.200 86.100 226.600 86.200 ;
        RECT 225.400 85.800 226.600 86.100 ;
        RECT 223.800 85.200 224.100 85.800 ;
        RECT 227.000 85.200 227.300 86.800 ;
        RECT 223.800 84.800 224.200 85.200 ;
        RECT 227.000 84.800 227.400 85.200 ;
        RECT 229.400 84.800 229.800 85.200 ;
        RECT 220.600 83.800 221.000 84.200 ;
        RECT 219.800 79.800 220.200 80.200 ;
        RECT 219.800 75.200 220.100 79.800 ;
        RECT 223.800 78.200 224.100 84.800 ;
        RECT 227.000 83.800 227.400 84.200 ;
        RECT 227.000 79.200 227.300 83.800 ;
        RECT 227.000 78.800 227.400 79.200 ;
        RECT 223.800 77.800 224.200 78.200 ;
        RECT 219.800 74.800 220.200 75.200 ;
        RECT 228.600 74.800 229.000 75.200 ;
        RECT 220.600 73.800 221.000 74.200 ;
        RECT 220.600 73.200 220.900 73.800 ;
        RECT 220.600 72.800 221.000 73.200 ;
        RECT 218.200 71.800 218.600 72.200 ;
        RECT 227.000 69.800 227.400 70.200 ;
        RECT 211.800 68.800 212.200 69.200 ;
        RECT 211.000 66.800 211.400 67.200 ;
        RECT 207.800 65.800 208.200 66.200 ;
        RECT 208.600 66.100 209.000 66.200 ;
        RECT 209.400 66.100 209.800 66.200 ;
        RECT 208.600 65.800 209.800 66.100 ;
        RECT 210.200 65.800 210.600 66.200 ;
        RECT 207.800 65.200 208.100 65.800 ;
        RECT 207.800 64.800 208.200 65.200 ;
        RECT 208.600 65.100 209.000 65.200 ;
        RECT 209.400 65.100 209.800 65.200 ;
        RECT 208.600 64.800 209.800 65.100 ;
        RECT 210.200 62.800 210.600 63.200 ;
        RECT 206.200 59.800 206.600 60.200 ;
        RECT 206.200 55.800 206.600 56.200 ;
        RECT 206.200 55.200 206.500 55.800 ;
        RECT 206.200 54.800 206.600 55.200 ;
        RECT 207.000 54.800 207.400 55.200 ;
        RECT 208.600 55.100 209.000 55.200 ;
        RECT 209.400 55.100 209.800 55.200 ;
        RECT 208.600 54.800 209.800 55.100 ;
        RECT 205.400 50.800 205.800 51.200 ;
        RECT 207.000 48.200 207.300 54.800 ;
        RECT 210.200 50.200 210.500 62.800 ;
        RECT 211.000 62.200 211.300 66.800 ;
        RECT 212.600 64.100 213.000 64.200 ;
        RECT 213.400 64.100 213.800 64.200 ;
        RECT 212.600 63.800 213.800 64.100 ;
        RECT 214.200 63.100 214.600 68.900 ;
        RECT 216.600 66.100 217.000 66.200 ;
        RECT 217.400 66.100 217.800 66.200 ;
        RECT 216.600 65.800 217.800 66.100 ;
        RECT 219.000 63.100 219.400 68.900 ;
        RECT 220.600 65.100 221.000 67.900 ;
        RECT 221.400 65.100 221.800 67.900 ;
        RECT 223.000 63.100 223.400 68.900 ;
        RECT 227.000 68.200 227.300 69.800 ;
        RECT 228.600 69.200 228.900 74.800 ;
        RECT 227.000 67.800 227.400 68.200 ;
        RECT 225.400 66.800 225.800 67.200 ;
        RECT 224.600 65.800 225.000 66.200 ;
        RECT 224.600 65.200 224.900 65.800 ;
        RECT 224.600 64.800 225.000 65.200 ;
        RECT 211.000 61.800 211.400 62.200 ;
        RECT 214.200 61.800 214.600 62.200 ;
        RECT 213.400 55.800 213.800 56.200 ;
        RECT 213.400 55.200 213.700 55.800 ;
        RECT 211.000 54.800 211.400 55.200 ;
        RECT 213.400 54.800 213.800 55.200 ;
        RECT 211.000 50.200 211.300 54.800 ;
        RECT 214.200 54.200 214.500 61.800 ;
        RECT 215.000 58.800 215.400 59.200 ;
        RECT 215.000 55.200 215.300 58.800 ;
        RECT 216.600 56.100 217.000 56.200 ;
        RECT 215.800 55.800 217.000 56.100 ;
        RECT 215.000 54.800 215.400 55.200 ;
        RECT 214.200 53.800 214.600 54.200 ;
        RECT 214.200 53.200 214.500 53.800 ;
        RECT 214.200 52.800 214.600 53.200 ;
        RECT 211.800 51.800 212.200 52.200 ;
        RECT 214.200 51.800 214.600 52.200 ;
        RECT 210.200 49.800 210.600 50.200 ;
        RECT 211.000 49.800 211.400 50.200 ;
        RECT 205.400 47.800 205.800 48.200 ;
        RECT 207.000 47.800 207.400 48.200 ;
        RECT 208.600 47.800 209.000 48.200 ;
        RECT 196.600 46.800 197.000 47.200 ;
        RECT 203.000 46.800 203.400 47.200 ;
        RECT 203.800 46.800 204.200 47.200 ;
        RECT 204.600 46.800 205.000 47.200 ;
        RECT 196.600 46.200 196.900 46.800 ;
        RECT 203.000 46.200 203.300 46.800 ;
        RECT 196.600 45.800 197.000 46.200 ;
        RECT 203.000 45.800 203.400 46.200 ;
        RECT 199.000 41.800 199.400 42.200 ;
        RECT 191.800 33.800 192.200 34.200 ;
        RECT 192.600 32.100 193.000 37.900 ;
        RECT 199.000 37.200 199.300 41.800 ;
        RECT 199.000 36.800 199.400 37.200 ;
        RECT 201.400 36.800 201.800 37.200 ;
        RECT 203.000 36.800 203.400 37.200 ;
        RECT 193.400 33.800 193.800 34.200 ;
        RECT 185.400 31.800 186.600 32.100 ;
        RECT 184.600 30.800 185.700 31.100 ;
        RECT 179.000 23.800 179.400 24.200 ;
        RECT 179.800 23.100 180.200 28.900 ;
        RECT 181.400 26.200 181.700 30.800 ;
        RECT 185.400 29.200 185.700 30.800 ;
        RECT 180.600 25.800 181.000 26.200 ;
        RECT 181.400 25.800 181.800 26.200 ;
        RECT 172.600 15.800 173.000 16.200 ;
        RECT 172.600 15.200 172.900 15.800 ;
        RECT 172.600 14.800 173.000 15.200 ;
        RECT 172.600 14.100 173.000 14.200 ;
        RECT 171.800 13.800 173.000 14.100 ;
        RECT 173.400 13.100 173.800 15.900 ;
        RECT 174.200 13.800 174.600 14.200 ;
        RECT 174.200 12.200 174.500 13.800 ;
        RECT 171.000 11.800 171.400 12.200 ;
        RECT 174.200 11.800 174.600 12.200 ;
        RECT 175.000 12.100 175.400 17.900 ;
        RECT 177.400 16.800 177.800 17.200 ;
        RECT 176.600 14.800 177.000 15.200 ;
        RECT 164.600 9.800 165.000 10.200 ;
        RECT 164.600 9.200 164.900 9.800 ;
        RECT 164.600 8.800 165.000 9.200 ;
        RECT 155.000 4.800 155.400 5.200 ;
        RECT 155.800 4.800 156.200 5.200 ;
        RECT 158.200 4.800 158.600 5.200 ;
        RECT 161.400 5.100 161.800 5.200 ;
        RECT 162.200 5.100 162.600 5.200 ;
        RECT 161.400 4.800 162.600 5.100 ;
        RECT 167.000 3.100 167.400 8.900 ;
        RECT 171.000 8.200 171.300 11.800 ;
        RECT 176.600 10.200 176.900 14.800 ;
        RECT 176.600 9.800 177.000 10.200 ;
        RECT 177.400 9.200 177.700 16.800 ;
        RECT 179.800 12.100 180.200 17.900 ;
        RECT 180.600 17.200 180.900 25.800 ;
        RECT 184.600 23.100 185.000 28.900 ;
        RECT 185.400 28.800 185.800 29.200 ;
        RECT 186.200 25.100 186.600 27.900 ;
        RECT 187.800 27.800 188.200 28.200 ;
        RECT 186.200 19.100 186.600 19.200 ;
        RECT 187.000 19.100 187.400 19.200 ;
        RECT 186.200 18.800 187.400 19.100 ;
        RECT 180.600 16.800 181.000 17.200 ;
        RECT 187.000 15.800 187.400 16.200 ;
        RECT 187.000 15.200 187.300 15.800 ;
        RECT 187.000 14.800 187.400 15.200 ;
        RECT 185.400 12.800 185.800 13.200 ;
        RECT 185.400 12.200 185.700 12.800 ;
        RECT 182.200 12.100 182.600 12.200 ;
        RECT 183.000 12.100 183.400 12.200 ;
        RECT 182.200 11.800 183.400 12.100 ;
        RECT 183.800 11.800 184.200 12.200 ;
        RECT 185.400 11.800 185.800 12.200 ;
        RECT 183.800 11.200 184.100 11.800 ;
        RECT 182.200 10.800 182.600 11.200 ;
        RECT 183.800 10.800 184.200 11.200 ;
        RECT 171.000 7.800 171.400 8.200 ;
        RECT 169.400 6.100 169.800 6.200 ;
        RECT 170.200 6.100 170.600 6.200 ;
        RECT 169.400 5.800 170.600 6.100 ;
        RECT 171.800 3.100 172.200 8.900 ;
        RECT 177.400 8.800 177.800 9.200 ;
        RECT 173.400 5.100 173.800 7.900 ;
        RECT 182.200 7.200 182.500 10.800 ;
        RECT 183.000 9.800 183.400 10.200 ;
        RECT 183.000 9.200 183.300 9.800 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 183.800 8.800 184.200 9.200 ;
        RECT 185.400 8.800 185.800 9.200 ;
        RECT 183.800 8.200 184.100 8.800 ;
        RECT 185.400 8.200 185.700 8.800 ;
        RECT 183.800 7.800 184.200 8.200 ;
        RECT 185.400 7.800 185.800 8.200 ;
        RECT 187.800 7.200 188.100 27.800 ;
        RECT 188.600 25.100 189.000 27.900 ;
        RECT 190.200 23.100 190.600 28.900 ;
        RECT 191.000 25.900 191.400 26.300 ;
        RECT 191.000 25.200 191.300 25.900 ;
        RECT 191.000 24.800 191.400 25.200 ;
        RECT 193.400 17.200 193.700 33.800 ;
        RECT 194.200 33.100 194.600 35.900 ;
        RECT 198.200 35.800 198.600 36.200 ;
        RECT 199.000 35.800 199.400 36.200 ;
        RECT 200.600 35.800 201.000 36.200 ;
        RECT 198.200 35.200 198.500 35.800 ;
        RECT 197.400 34.800 197.800 35.200 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 196.600 33.800 197.000 34.200 ;
        RECT 196.600 33.200 196.900 33.800 ;
        RECT 196.600 32.800 197.000 33.200 ;
        RECT 196.600 30.200 196.900 32.800 ;
        RECT 196.600 29.800 197.000 30.200 ;
        RECT 195.000 23.100 195.400 28.900 ;
        RECT 196.600 26.800 197.000 27.200 ;
        RECT 196.600 24.100 196.900 26.800 ;
        RECT 197.400 26.200 197.700 34.800 ;
        RECT 199.000 29.200 199.300 35.800 ;
        RECT 200.600 35.200 200.900 35.800 ;
        RECT 199.800 34.800 200.200 35.200 ;
        RECT 200.600 34.800 201.000 35.200 ;
        RECT 199.800 34.200 200.100 34.800 ;
        RECT 199.800 33.800 200.200 34.200 ;
        RECT 199.800 31.800 200.200 32.200 ;
        RECT 199.000 28.800 199.400 29.200 ;
        RECT 199.800 27.200 200.100 31.800 ;
        RECT 199.800 26.800 200.200 27.200 ;
        RECT 200.600 26.800 201.000 27.200 ;
        RECT 200.600 26.200 200.900 26.800 ;
        RECT 197.400 25.800 197.800 26.200 ;
        RECT 198.200 25.800 198.600 26.200 ;
        RECT 200.600 25.800 201.000 26.200 ;
        RECT 198.200 25.200 198.500 25.800 ;
        RECT 198.200 24.800 198.600 25.200 ;
        RECT 197.400 24.100 197.800 24.200 ;
        RECT 196.600 23.800 197.800 24.100 ;
        RECT 201.400 20.200 201.700 36.800 ;
        RECT 203.000 36.200 203.300 36.800 ;
        RECT 203.000 35.800 203.400 36.200 ;
        RECT 202.200 32.800 202.600 33.200 ;
        RECT 202.200 32.200 202.500 32.800 ;
        RECT 202.200 31.800 202.600 32.200 ;
        RECT 202.200 30.800 202.600 31.200 ;
        RECT 202.200 29.200 202.500 30.800 ;
        RECT 202.200 28.800 202.600 29.200 ;
        RECT 201.400 19.800 201.800 20.200 ;
        RECT 193.400 16.800 193.800 17.200 ;
        RECT 189.400 15.800 189.800 16.200 ;
        RECT 189.400 14.200 189.700 15.800 ;
        RECT 189.400 13.800 189.800 14.200 ;
        RECT 188.600 12.800 189.000 13.200 ;
        RECT 188.600 12.200 188.900 12.800 ;
        RECT 188.600 12.100 189.000 12.200 ;
        RECT 189.400 12.100 189.800 12.200 ;
        RECT 188.600 11.800 189.800 12.100 ;
        RECT 193.400 11.800 193.800 12.200 ;
        RECT 194.200 12.100 194.600 17.900 ;
        RECT 195.800 14.800 196.200 15.200 ;
        RECT 193.400 7.200 193.700 11.800 ;
        RECT 195.800 9.200 196.100 14.800 ;
        RECT 198.200 12.800 198.600 13.200 ;
        RECT 195.800 8.800 196.200 9.200 ;
        RECT 182.200 6.800 182.600 7.200 ;
        RECT 187.800 6.800 188.200 7.200 ;
        RECT 193.400 6.800 193.800 7.200 ;
        RECT 198.200 6.200 198.500 12.800 ;
        RECT 199.000 12.100 199.400 17.900 ;
        RECT 200.600 13.100 201.000 15.900 ;
        RECT 201.400 15.200 201.700 19.800 ;
        RECT 201.400 14.800 201.800 15.200 ;
        RECT 202.200 14.800 202.600 15.200 ;
        RECT 202.200 10.200 202.500 14.800 ;
        RECT 202.200 9.800 202.600 10.200 ;
        RECT 198.200 5.800 198.600 6.200 ;
        RECT 189.400 4.800 189.800 5.200 ;
        RECT 199.800 5.100 200.200 7.900 ;
        RECT 189.400 4.200 189.700 4.800 ;
        RECT 189.400 3.800 189.800 4.200 ;
        RECT 201.400 3.100 201.800 8.900 ;
        RECT 202.200 5.900 202.600 6.300 ;
        RECT 202.200 5.200 202.500 5.900 ;
        RECT 203.000 5.200 203.300 35.800 ;
        RECT 203.800 30.200 204.100 46.800 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 204.600 34.200 204.900 45.800 ;
        RECT 205.400 39.200 205.700 47.800 ;
        RECT 208.600 47.200 208.900 47.800 ;
        RECT 208.600 46.800 209.000 47.200 ;
        RECT 210.200 46.200 210.500 49.800 ;
        RECT 211.800 47.200 212.100 51.800 ;
        RECT 214.200 47.200 214.500 51.800 ;
        RECT 211.800 46.800 212.200 47.200 ;
        RECT 213.400 46.800 213.800 47.200 ;
        RECT 214.200 46.800 214.600 47.200 ;
        RECT 213.400 46.200 213.700 46.800 ;
        RECT 207.000 45.800 207.400 46.200 ;
        RECT 207.800 46.100 208.200 46.200 ;
        RECT 208.600 46.100 209.000 46.200 ;
        RECT 207.800 45.800 209.000 46.100 ;
        RECT 210.200 45.800 210.600 46.200 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 212.600 45.800 213.000 46.200 ;
        RECT 213.400 45.800 213.800 46.200 ;
        RECT 207.000 44.200 207.300 45.800 ;
        RECT 210.200 45.200 210.500 45.800 ;
        RECT 210.200 44.800 210.600 45.200 ;
        RECT 207.000 43.800 207.400 44.200 ;
        RECT 205.400 38.800 205.800 39.200 ;
        RECT 204.600 33.800 205.000 34.200 ;
        RECT 204.600 31.200 204.900 33.800 ;
        RECT 207.800 32.100 208.200 37.900 ;
        RECT 211.800 35.100 212.100 45.800 ;
        RECT 212.600 45.200 212.900 45.800 ;
        RECT 212.600 44.800 213.000 45.200 ;
        RECT 215.000 45.100 215.300 54.800 ;
        RECT 215.800 49.200 216.100 55.800 ;
        RECT 216.600 55.100 217.000 55.200 ;
        RECT 217.400 55.100 217.800 55.200 ;
        RECT 216.600 54.800 217.800 55.100 ;
        RECT 216.600 52.100 217.000 52.200 ;
        RECT 217.400 52.100 217.800 52.200 ;
        RECT 219.800 52.100 220.200 57.900 ;
        RECT 221.400 55.100 221.800 55.200 ;
        RECT 222.200 55.100 222.600 55.200 ;
        RECT 221.400 54.800 222.600 55.100 ;
        RECT 224.600 52.100 225.000 57.900 ;
        RECT 225.400 54.200 225.700 66.800 ;
        RECT 227.800 63.100 228.200 68.900 ;
        RECT 228.600 68.800 229.000 69.200 ;
        RECT 229.400 63.200 229.700 84.800 ;
        RECT 229.400 62.800 229.800 63.200 ;
        RECT 230.200 61.800 230.600 62.200 ;
        RECT 225.400 53.800 225.800 54.200 ;
        RECT 216.600 51.800 217.800 52.100 ;
        RECT 219.800 49.800 220.200 50.200 ;
        RECT 219.800 49.200 220.100 49.800 ;
        RECT 215.800 48.800 216.200 49.200 ;
        RECT 217.400 48.800 217.800 49.200 ;
        RECT 219.800 48.800 220.200 49.200 ;
        RECT 216.600 46.800 217.000 47.200 ;
        RECT 215.800 45.100 216.200 45.200 ;
        RECT 215.000 44.800 216.200 45.100 ;
        RECT 215.800 40.800 216.200 41.200 ;
        RECT 211.800 34.700 212.200 35.100 ;
        RECT 212.600 32.100 213.000 37.900 ;
        RECT 215.800 36.200 216.100 40.800 ;
        RECT 213.400 33.800 213.800 34.200 ;
        RECT 204.600 30.800 205.000 31.200 ;
        RECT 203.800 29.800 204.200 30.200 ;
        RECT 211.000 29.800 211.400 30.200 ;
        RECT 203.800 27.200 204.100 29.800 ;
        RECT 209.400 28.800 209.800 29.200 ;
        RECT 209.400 28.200 209.700 28.800 ;
        RECT 209.400 27.800 209.800 28.200 ;
        RECT 203.800 26.800 204.200 27.200 ;
        RECT 206.200 27.100 206.600 27.200 ;
        RECT 207.000 27.100 207.400 27.200 ;
        RECT 206.200 26.800 207.400 27.100 ;
        RECT 203.800 26.100 204.200 26.200 ;
        RECT 204.600 26.100 205.000 26.200 ;
        RECT 203.800 25.800 205.000 26.100 ;
        RECT 207.000 25.800 207.400 26.200 ;
        RECT 207.000 25.200 207.300 25.800 ;
        RECT 207.000 24.800 207.400 25.200 ;
        RECT 203.800 23.800 204.200 24.200 ;
        RECT 203.800 19.200 204.100 23.800 ;
        RECT 203.800 18.800 204.200 19.200 ;
        RECT 207.800 15.800 208.200 16.200 ;
        RECT 207.800 14.200 208.100 15.800 ;
        RECT 210.200 14.800 210.600 15.200 ;
        RECT 210.200 14.200 210.500 14.800 ;
        RECT 211.000 14.200 211.300 29.800 ;
        RECT 211.800 23.100 212.200 28.900 ;
        RECT 213.400 27.200 213.700 33.800 ;
        RECT 214.200 33.100 214.600 35.900 ;
        RECT 215.800 35.800 216.200 36.200 ;
        RECT 215.800 35.200 216.100 35.800 ;
        RECT 216.600 35.200 216.900 46.800 ;
        RECT 217.400 46.200 217.700 48.800 ;
        RECT 220.600 46.800 221.000 47.200 ;
        RECT 217.400 45.800 217.800 46.200 ;
        RECT 219.000 46.100 219.400 46.200 ;
        RECT 219.800 46.100 220.200 46.200 ;
        RECT 219.000 45.800 220.200 46.100 ;
        RECT 219.000 44.800 219.400 45.200 ;
        RECT 217.400 36.100 217.800 36.200 ;
        RECT 218.200 36.100 218.600 36.200 ;
        RECT 217.400 35.800 218.600 36.100 ;
        RECT 215.000 34.800 215.400 35.200 ;
        RECT 215.800 34.800 216.200 35.200 ;
        RECT 216.600 34.800 217.000 35.200 ;
        RECT 218.200 34.800 218.600 35.200 ;
        RECT 215.000 34.200 215.300 34.800 ;
        RECT 218.200 34.200 218.500 34.800 ;
        RECT 215.000 33.800 215.400 34.200 ;
        RECT 218.200 33.800 218.600 34.200 ;
        RECT 219.000 29.200 219.300 44.800 ;
        RECT 219.800 43.800 220.200 44.200 ;
        RECT 219.800 37.200 220.100 43.800 ;
        RECT 219.800 36.800 220.200 37.200 ;
        RECT 219.800 34.200 220.100 36.800 ;
        RECT 219.800 33.800 220.200 34.200 ;
        RECT 219.800 32.800 220.200 33.200 ;
        RECT 213.400 26.800 213.800 27.200 ;
        RECT 215.000 26.800 215.400 27.200 ;
        RECT 215.800 26.800 216.200 27.200 ;
        RECT 215.000 26.200 215.300 26.800 ;
        RECT 215.000 25.800 215.400 26.200 ;
        RECT 215.000 15.800 215.400 16.200 ;
        RECT 215.000 15.200 215.300 15.800 ;
        RECT 211.800 15.100 212.200 15.200 ;
        RECT 212.600 15.100 213.000 15.200 ;
        RECT 211.800 14.800 213.000 15.100 ;
        RECT 215.000 14.800 215.400 15.200 ;
        RECT 206.200 13.800 206.600 14.200 ;
        RECT 207.800 13.800 208.200 14.200 ;
        RECT 210.200 13.800 210.600 14.200 ;
        RECT 211.000 13.800 211.400 14.200 ;
        RECT 206.200 11.200 206.500 13.800 ;
        RECT 208.600 12.100 209.000 12.200 ;
        RECT 209.400 12.100 209.800 12.200 ;
        RECT 208.600 11.800 209.800 12.100 ;
        RECT 213.400 11.800 213.800 12.200 ;
        RECT 214.200 11.800 214.600 12.200 ;
        RECT 206.200 10.800 206.600 11.200 ;
        RECT 209.400 10.800 209.800 11.200 ;
        RECT 209.400 9.200 209.700 10.800 ;
        RECT 207.800 9.100 208.200 9.200 ;
        RECT 208.600 9.100 209.000 9.200 ;
        RECT 204.600 6.100 205.000 6.200 ;
        RECT 205.400 6.100 205.800 6.200 ;
        RECT 204.600 5.800 205.800 6.100 ;
        RECT 202.200 4.800 202.600 5.200 ;
        RECT 203.000 4.800 203.400 5.200 ;
        RECT 206.200 3.100 206.600 8.900 ;
        RECT 207.800 8.800 209.000 9.100 ;
        RECT 209.400 8.800 209.800 9.200 ;
        RECT 211.800 3.100 212.200 8.900 ;
        RECT 213.400 6.200 213.700 11.800 ;
        RECT 214.200 7.200 214.500 11.800 ;
        RECT 215.800 8.200 216.100 26.800 ;
        RECT 216.600 23.100 217.000 28.900 ;
        RECT 219.000 28.800 219.400 29.200 ;
        RECT 218.200 25.100 218.600 27.900 ;
        RECT 219.000 25.800 219.400 26.200 ;
        RECT 219.000 25.200 219.300 25.800 ;
        RECT 219.000 24.800 219.400 25.200 ;
        RECT 216.600 13.800 217.000 14.200 ;
        RECT 216.600 10.200 216.900 13.800 ;
        RECT 216.600 9.800 217.000 10.200 ;
        RECT 219.800 9.200 220.100 32.800 ;
        RECT 220.600 27.200 220.900 46.800 ;
        RECT 222.200 43.100 222.600 48.900 ;
        RECT 225.400 47.200 225.700 53.800 ;
        RECT 226.200 53.100 226.600 55.900 ;
        RECT 227.000 55.800 227.400 56.200 ;
        RECT 227.000 55.200 227.300 55.800 ;
        RECT 227.000 54.800 227.400 55.200 ;
        RECT 228.600 54.100 229.000 54.200 ;
        RECT 229.400 54.100 229.800 54.200 ;
        RECT 228.600 53.800 229.800 54.100 ;
        RECT 225.400 46.800 225.800 47.200 ;
        RECT 223.800 46.100 224.200 46.200 ;
        RECT 224.600 46.100 225.000 46.200 ;
        RECT 223.800 45.800 225.000 46.100 ;
        RECT 223.000 32.100 223.400 37.900 ;
        RECT 224.600 35.100 225.000 35.200 ;
        RECT 225.400 35.100 225.700 46.800 ;
        RECT 227.000 43.100 227.400 48.900 ;
        RECT 228.600 45.100 229.000 47.900 ;
        RECT 224.600 34.800 225.700 35.100 ;
        RECT 226.200 34.800 226.600 35.200 ;
        RECT 221.400 30.800 221.800 31.200 ;
        RECT 221.400 29.200 221.700 30.800 ;
        RECT 221.400 28.800 221.800 29.200 ;
        RECT 220.600 26.800 221.000 27.200 ;
        RECT 220.600 25.800 221.000 26.200 ;
        RECT 215.800 7.800 216.200 8.200 ;
        RECT 214.200 6.800 214.600 7.200 ;
        RECT 213.400 5.800 213.800 6.200 ;
        RECT 216.600 3.100 217.000 8.900 ;
        RECT 219.800 8.800 220.200 9.200 ;
        RECT 217.400 6.800 217.800 7.200 ;
        RECT 217.400 6.200 217.700 6.800 ;
        RECT 217.400 5.800 217.800 6.200 ;
        RECT 218.200 5.100 218.600 7.900 ;
        RECT 220.600 7.200 220.900 25.800 ;
        RECT 223.800 23.100 224.200 28.900 ;
        RECT 224.600 27.200 224.900 34.800 ;
        RECT 226.200 34.200 226.500 34.800 ;
        RECT 226.200 33.800 226.600 34.200 ;
        RECT 225.400 32.800 225.800 33.200 ;
        RECT 224.600 26.800 225.000 27.200 ;
        RECT 224.600 26.200 224.900 26.800 ;
        RECT 224.600 25.800 225.000 26.200 ;
        RECT 225.400 25.100 225.700 32.800 ;
        RECT 227.000 31.800 227.400 32.200 ;
        RECT 227.800 32.100 228.200 37.900 ;
        RECT 229.400 33.100 229.800 35.900 ;
        RECT 230.200 33.200 230.500 61.800 ;
        RECT 230.200 32.800 230.600 33.200 ;
        RECT 227.000 26.200 227.300 31.800 ;
        RECT 227.000 25.800 227.400 26.200 ;
        RECT 224.600 24.800 225.700 25.100 ;
        RECT 224.600 14.200 224.900 24.800 ;
        RECT 228.600 23.100 229.000 28.900 ;
        RECT 229.400 26.800 229.800 27.200 ;
        RECT 228.600 21.800 229.000 22.200 ;
        RECT 228.600 19.200 228.900 21.800 ;
        RECT 228.600 18.800 229.000 19.200 ;
        RECT 225.400 16.100 225.800 16.200 ;
        RECT 226.200 16.100 226.600 16.200 ;
        RECT 225.400 15.800 226.600 16.100 ;
        RECT 228.600 15.800 229.000 16.200 ;
        RECT 228.600 15.200 228.900 15.800 ;
        RECT 228.600 14.800 229.000 15.200 ;
        RECT 229.400 14.200 229.700 26.800 ;
        RECT 230.200 25.100 230.600 27.900 ;
        RECT 224.600 13.800 225.000 14.200 ;
        RECT 229.400 13.800 229.800 14.200 ;
        RECT 223.000 11.800 223.400 12.200 ;
        RECT 221.400 9.800 221.800 10.200 ;
        RECT 221.400 9.200 221.700 9.800 ;
        RECT 221.400 8.800 221.800 9.200 ;
        RECT 220.600 6.800 221.000 7.200 ;
        RECT 223.000 6.200 223.300 11.800 ;
        RECT 223.000 5.800 223.400 6.200 ;
        RECT 219.000 4.800 219.400 5.200 ;
        RECT 219.000 4.200 219.300 4.800 ;
        RECT 219.000 3.800 219.400 4.200 ;
        RECT 223.800 3.100 224.200 8.900 ;
        RECT 227.000 6.800 227.400 7.200 ;
        RECT 227.000 6.200 227.300 6.800 ;
        RECT 224.600 6.100 225.000 6.200 ;
        RECT 225.400 6.100 225.800 6.200 ;
        RECT 224.600 5.800 225.800 6.100 ;
        RECT 227.000 5.800 227.400 6.200 ;
        RECT 228.600 3.100 229.000 8.900 ;
        RECT 230.200 5.100 230.600 7.900 ;
      LAYER via2 ;
        RECT 1.400 197.800 1.800 198.200 ;
        RECT 15.800 196.800 16.200 197.200 ;
        RECT 22.200 196.800 22.600 197.200 ;
        RECT 11.000 194.800 11.400 195.200 ;
        RECT 5.400 185.800 5.800 186.200 ;
        RECT 15.800 194.800 16.200 195.200 ;
        RECT 16.600 193.800 17.000 194.200 ;
        RECT 11.000 184.800 11.400 185.200 ;
        RECT 10.200 183.800 10.600 184.200 ;
        RECT 26.200 196.800 26.600 197.200 ;
        RECT 28.600 194.800 29.000 195.200 ;
        RECT 57.400 206.800 57.800 207.200 ;
        RECT 55.000 203.800 55.400 204.200 ;
        RECT 58.200 194.800 58.600 195.200 ;
        RECT 51.000 193.800 51.400 194.200 ;
        RECT 52.600 193.800 53.000 194.200 ;
        RECT 26.200 183.800 26.600 184.200 ;
        RECT 17.400 166.800 17.800 167.200 ;
        RECT 18.200 165.800 18.600 166.200 ;
        RECT 3.800 153.800 4.200 154.200 ;
        RECT 4.600 152.800 5.000 153.200 ;
        RECT 10.200 148.800 10.600 149.200 ;
        RECT 3.000 125.800 3.400 126.200 ;
        RECT 34.200 178.800 34.600 179.200 ;
        RECT 29.400 174.800 29.800 175.200 ;
        RECT 35.000 174.800 35.400 175.200 ;
        RECT 47.800 185.800 48.200 186.200 ;
        RECT 58.200 186.800 58.600 187.200 ;
        RECT 61.400 186.800 61.800 187.200 ;
        RECT 54.200 185.800 54.600 186.200 ;
        RECT 48.600 174.800 49.000 175.200 ;
        RECT 12.600 145.800 13.000 146.200 ;
        RECT 12.600 133.800 13.000 134.200 ;
        RECT 15.000 134.800 15.400 135.200 ;
        RECT 32.600 164.800 33.000 165.200 ;
        RECT 31.800 151.800 32.200 152.200 ;
        RECT 63.000 185.800 63.400 186.200 ;
        RECT 59.000 184.800 59.400 185.200 ;
        RECT 57.400 175.800 57.800 176.200 ;
        RECT 55.800 174.800 56.200 175.200 ;
        RECT 58.200 166.800 58.600 167.200 ;
        RECT 51.800 165.800 52.200 166.200 ;
        RECT 44.600 156.800 45.000 157.200 ;
        RECT 43.800 153.800 44.200 154.200 ;
        RECT 31.000 146.800 31.400 147.200 ;
        RECT 34.200 146.800 34.600 147.200 ;
        RECT 18.200 145.800 18.600 146.200 ;
        RECT 19.800 125.800 20.200 126.200 ;
        RECT 60.600 164.800 61.000 165.200 ;
        RECT 68.600 205.800 69.000 206.200 ;
        RECT 88.600 205.800 89.000 206.200 ;
        RECT 69.400 186.800 69.800 187.200 ;
        RECT 68.600 167.800 69.000 168.200 ;
        RECT 75.800 194.800 76.200 195.200 ;
        RECT 45.400 146.800 45.800 147.200 ;
        RECT 47.800 145.800 48.200 146.200 ;
        RECT 43.000 144.800 43.400 145.200 ;
        RECT 46.200 144.800 46.600 145.200 ;
        RECT 33.400 134.800 33.800 135.200 ;
        RECT 28.600 125.800 29.000 126.200 ;
        RECT 24.600 121.800 25.000 122.200 ;
        RECT 14.200 116.800 14.600 117.200 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 12.600 95.800 13.000 96.200 ;
        RECT 15.000 94.800 15.400 95.200 ;
        RECT 5.400 85.800 5.800 86.200 ;
        RECT 11.000 85.800 11.400 86.200 ;
        RECT 11.000 84.800 11.400 85.200 ;
        RECT 3.800 63.800 4.200 64.200 ;
        RECT 9.400 65.800 9.800 66.200 ;
        RECT 1.400 35.800 1.800 36.200 ;
        RECT 38.200 137.800 38.600 138.200 ;
        RECT 45.400 134.800 45.800 135.200 ;
        RECT 46.200 133.800 46.600 134.200 ;
        RECT 25.400 114.800 25.800 115.200 ;
        RECT 23.000 113.800 23.400 114.200 ;
        RECT 27.000 113.800 27.400 114.200 ;
        RECT 22.200 111.800 22.600 112.200 ;
        RECT 22.200 105.800 22.600 106.200 ;
        RECT 24.600 94.700 25.000 95.100 ;
        RECT 36.600 125.800 37.000 126.200 ;
        RECT 43.000 128.800 43.400 129.200 ;
        RECT 63.800 156.800 64.200 157.200 ;
        RECT 65.400 155.800 65.800 156.200 ;
        RECT 67.800 155.800 68.200 156.200 ;
        RECT 65.400 154.800 65.800 155.200 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 59.800 145.800 60.200 146.200 ;
        RECT 64.600 148.800 65.000 149.200 ;
        RECT 95.000 205.900 95.400 206.300 ;
        RECT 85.400 194.800 85.800 195.200 ;
        RECT 105.400 205.800 105.800 206.200 ;
        RECT 113.400 205.800 113.800 206.200 ;
        RECT 106.200 196.800 106.600 197.200 ;
        RECT 102.200 193.800 102.600 194.200 ;
        RECT 101.400 185.800 101.800 186.200 ;
        RECT 98.200 178.800 98.600 179.200 ;
        RECT 92.600 175.800 93.000 176.200 ;
        RECT 80.600 165.800 81.000 166.200 ;
        RECT 95.000 166.800 95.400 167.200 ;
        RECT 120.600 205.800 121.000 206.200 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 100.600 166.800 101.000 167.200 ;
        RECT 93.400 154.800 93.800 155.200 ;
        RECT 67.000 145.800 67.400 146.200 ;
        RECT 64.600 143.800 65.000 144.200 ;
        RECT 62.200 135.800 62.600 136.200 ;
        RECT 68.600 134.800 69.000 135.200 ;
        RECT 81.400 136.800 81.800 137.200 ;
        RECT 85.400 135.800 85.800 136.200 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 84.600 134.800 85.000 135.200 ;
        RECT 73.400 131.800 73.800 132.200 ;
        RECT 63.800 126.800 64.200 127.200 ;
        RECT 52.600 125.800 53.000 126.200 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 33.400 96.800 33.800 97.200 ;
        RECT 35.000 95.800 35.400 96.200 ;
        RECT 32.600 92.800 33.000 93.200 ;
        RECT 26.200 85.800 26.600 86.200 ;
        RECT 26.200 84.800 26.600 85.200 ;
        RECT 32.600 85.900 33.000 86.300 ;
        RECT 24.600 74.800 25.000 75.200 ;
        RECT 47.000 101.800 47.400 102.200 ;
        RECT 53.400 111.800 53.800 112.200 ;
        RECT 47.000 85.800 47.400 86.200 ;
        RECT 31.000 78.800 31.400 79.200 ;
        RECT 6.200 34.800 6.600 35.200 ;
        RECT 13.400 34.800 13.800 35.200 ;
        RECT 3.800 26.800 4.200 27.200 ;
        RECT 3.000 25.800 3.400 26.200 ;
        RECT 10.200 18.800 10.600 19.200 ;
        RECT 1.400 8.800 1.800 9.200 ;
        RECT 4.600 6.800 5.000 7.200 ;
        RECT 34.200 74.800 34.600 75.200 ;
        RECT 31.800 68.800 32.200 69.200 ;
        RECT 52.600 88.800 53.000 89.200 ;
        RECT 61.400 104.800 61.800 105.200 ;
        RECT 39.000 71.800 39.400 72.200 ;
        RECT 42.200 73.800 42.600 74.200 ;
        RECT 54.200 75.800 54.600 76.200 ;
        RECT 42.200 71.800 42.600 72.200 ;
        RECT 36.600 67.800 37.000 68.200 ;
        RECT 28.600 34.800 29.000 35.200 ;
        RECT 40.600 54.800 41.000 55.200 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 90.200 134.800 90.600 135.200 ;
        RECT 81.400 126.800 81.800 127.200 ;
        RECT 82.200 124.800 82.600 125.200 ;
        RECT 78.200 114.800 78.600 115.200 ;
        RECT 63.000 85.800 63.400 86.200 ;
        RECT 67.000 85.800 67.400 86.200 ;
        RECT 66.200 73.800 66.600 74.200 ;
        RECT 45.400 56.800 45.800 57.200 ;
        RECT 41.400 45.800 41.800 46.200 ;
        RECT 49.400 55.800 49.800 56.200 ;
        RECT 68.600 73.800 69.000 74.200 ;
        RECT 46.200 53.800 46.600 54.200 ;
        RECT 56.600 53.800 57.000 54.200 ;
        RECT 47.000 48.800 47.400 49.200 ;
        RECT 39.800 28.800 40.200 29.200 ;
        RECT 27.000 24.800 27.400 25.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 49.400 45.800 49.800 46.200 ;
        RECT 79.800 88.800 80.200 89.200 ;
        RECT 113.400 175.800 113.800 176.200 ;
        RECT 115.000 175.800 115.400 176.200 ;
        RECT 115.800 168.800 116.200 169.200 ;
        RECT 115.800 151.800 116.200 152.200 ;
        RECT 146.200 205.800 146.600 206.200 ;
        RECT 151.800 208.800 152.200 209.200 ;
        RECT 139.800 201.800 140.200 202.200 ;
        RECT 139.000 195.800 139.400 196.200 ;
        RECT 139.000 194.800 139.400 195.200 ;
        RECT 96.600 146.800 97.000 147.200 ;
        RECT 99.000 134.800 99.400 135.200 ;
        RECT 97.400 132.800 97.800 133.200 ;
        RECT 99.000 126.800 99.400 127.200 ;
        RECT 96.600 124.800 97.000 125.200 ;
        RECT 102.200 115.800 102.600 116.200 ;
        RECT 98.200 108.800 98.600 109.200 ;
        RECT 99.800 105.800 100.200 106.200 ;
        RECT 99.800 104.800 100.200 105.200 ;
        RECT 102.200 104.800 102.600 105.200 ;
        RECT 125.400 151.800 125.800 152.200 ;
        RECT 119.000 146.800 119.400 147.200 ;
        RECT 139.800 185.800 140.200 186.200 ;
        RECT 128.600 154.800 129.000 155.200 ;
        RECT 139.800 165.800 140.200 166.200 ;
        RECT 154.200 174.800 154.600 175.200 ;
        RECT 153.400 173.800 153.800 174.200 ;
        RECT 206.200 206.800 206.600 207.200 ;
        RECT 191.000 205.800 191.400 206.200 ;
        RECT 199.000 205.800 199.400 206.200 ;
        RECT 164.600 195.800 165.000 196.200 ;
        RECT 156.600 166.800 157.000 167.200 ;
        RECT 130.200 145.800 130.600 146.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 119.800 135.800 120.200 136.200 ;
        RECT 124.600 135.800 125.000 136.200 ;
        RECT 123.800 134.800 124.200 135.200 ;
        RECT 127.800 135.800 128.200 136.200 ;
        RECT 127.000 134.800 127.400 135.200 ;
        RECT 112.600 131.800 113.000 132.200 ;
        RECT 108.600 115.800 109.000 116.200 ;
        RECT 128.600 132.800 129.000 133.200 ;
        RECT 116.600 112.800 117.000 113.200 ;
        RECT 116.600 101.800 117.000 102.200 ;
        RECT 107.800 92.800 108.200 93.200 ;
        RECT 97.400 85.800 97.800 86.200 ;
        RECT 91.800 84.800 92.200 85.200 ;
        RECT 95.800 84.800 96.200 85.200 ;
        RECT 94.200 83.800 94.600 84.200 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 42.200 36.800 42.600 37.200 ;
        RECT 50.200 34.800 50.600 35.200 ;
        RECT 51.000 26.800 51.400 27.200 ;
        RECT 70.200 45.800 70.600 46.200 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 65.400 35.800 65.800 36.200 ;
        RECT 79.000 34.800 79.400 35.200 ;
        RECT 50.200 25.800 50.600 26.200 ;
        RECT 29.400 14.800 29.800 15.200 ;
        RECT 35.000 15.800 35.400 16.200 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 34.200 11.800 34.600 12.200 ;
        RECT 4.600 4.800 5.000 5.200 ;
        RECT 14.200 4.800 14.600 5.200 ;
        RECT 58.200 14.800 58.600 15.200 ;
        RECT 70.200 28.800 70.600 29.200 ;
        RECT 80.600 31.800 81.000 32.200 ;
        RECT 81.400 26.800 81.800 27.200 ;
        RECT 81.400 24.800 81.800 25.200 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 108.600 73.800 109.000 74.200 ;
        RECT 103.000 67.800 103.400 68.200 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 101.400 66.800 101.800 67.200 ;
        RECT 103.800 65.800 104.200 66.200 ;
        RECT 103.000 56.800 103.400 57.200 ;
        RECT 115.000 74.800 115.400 75.200 ;
        RECT 112.600 66.800 113.000 67.200 ;
        RECT 107.800 56.800 108.200 57.200 ;
        RECT 103.800 55.800 104.200 56.200 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 101.400 35.800 101.800 36.200 ;
        RECT 90.200 25.800 90.600 26.200 ;
        RECT 46.200 4.800 46.600 5.200 ;
        RECT 68.600 8.800 69.000 9.200 ;
        RECT 77.400 13.800 77.800 14.200 ;
        RECT 79.800 13.800 80.200 14.200 ;
        RECT 81.400 13.800 81.800 14.200 ;
        RECT 101.400 28.800 101.800 29.200 ;
        RECT 130.200 125.800 130.600 126.200 ;
        RECT 170.200 166.800 170.600 167.200 ;
        RECT 159.000 156.800 159.400 157.200 ;
        RECT 153.400 141.800 153.800 142.200 ;
        RECT 139.000 134.800 139.400 135.200 ;
        RECT 142.200 128.800 142.600 129.200 ;
        RECT 121.400 88.800 121.800 89.200 ;
        RECT 123.000 73.800 123.400 74.200 ;
        RECT 131.800 88.800 132.200 89.200 ;
        RECT 179.000 164.800 179.400 165.200 ;
        RECT 207.000 204.800 207.400 205.200 ;
        RECT 204.600 194.800 205.000 195.200 ;
        RECT 180.600 155.800 181.000 156.200 ;
        RECT 183.800 153.800 184.200 154.200 ;
        RECT 175.800 151.800 176.200 152.200 ;
        RECT 176.600 145.800 177.000 146.200 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 167.000 133.800 167.400 134.200 ;
        RECT 165.400 126.800 165.800 127.200 ;
        RECT 176.600 133.800 177.000 134.200 ;
        RECT 177.400 126.800 177.800 127.200 ;
        RECT 168.600 124.800 169.000 125.200 ;
        RECT 171.000 124.800 171.400 125.200 ;
        RECT 163.800 115.800 164.200 116.200 ;
        RECT 167.000 115.800 167.400 116.200 ;
        RECT 137.400 103.800 137.800 104.200 ;
        RECT 143.000 94.800 143.400 95.200 ;
        RECT 144.600 86.800 145.000 87.200 ;
        RECT 167.800 108.800 168.200 109.200 ;
        RECT 167.000 106.800 167.400 107.200 ;
        RECT 135.000 71.800 135.400 72.200 ;
        RECT 157.400 86.800 157.800 87.200 ;
        RECT 151.000 74.800 151.400 75.200 ;
        RECT 150.200 68.800 150.600 69.200 ;
        RECT 141.400 65.800 141.800 66.200 ;
        RECT 132.600 58.800 133.000 59.200 ;
        RECT 131.800 56.800 132.200 57.200 ;
        RECT 108.600 34.800 109.000 35.200 ;
        RECT 115.000 5.800 115.400 6.200 ;
        RECT 200.600 173.800 201.000 174.200 ;
        RECT 223.800 206.800 224.200 207.200 ;
        RECT 226.200 204.800 226.600 205.200 ;
        RECT 210.200 176.800 210.600 177.200 ;
        RECT 209.400 154.800 209.800 155.200 ;
        RECT 194.200 145.800 194.600 146.200 ;
        RECT 205.400 153.800 205.800 154.200 ;
        RECT 225.400 184.800 225.800 185.200 ;
        RECT 214.200 154.800 214.600 155.200 ;
        RECT 207.800 135.800 208.200 136.200 ;
        RECT 223.800 164.800 224.200 165.200 ;
        RECT 186.200 114.800 186.600 115.200 ;
        RECT 183.800 111.800 184.200 112.200 ;
        RECT 189.400 106.800 189.800 107.200 ;
        RECT 175.800 97.800 176.200 98.200 ;
        RECT 166.200 88.800 166.600 89.200 ;
        RECT 165.400 87.800 165.800 88.200 ;
        RECT 181.400 96.800 181.800 97.200 ;
        RECT 180.600 94.800 181.000 95.200 ;
        RECT 189.400 105.800 189.800 106.200 ;
        RECT 186.200 104.800 186.600 105.200 ;
        RECT 190.200 104.800 190.600 105.200 ;
        RECT 185.400 93.800 185.800 94.200 ;
        RECT 169.400 87.800 169.800 88.200 ;
        RECT 168.600 86.800 169.000 87.200 ;
        RECT 171.800 86.800 172.200 87.200 ;
        RECT 179.000 85.800 179.400 86.200 ;
        RECT 166.200 84.800 166.600 85.200 ;
        RECT 155.800 73.800 156.200 74.200 ;
        RECT 211.000 127.800 211.400 128.200 ;
        RECT 203.000 125.800 203.400 126.200 ;
        RECT 210.200 125.800 210.600 126.200 ;
        RECT 217.400 125.800 217.800 126.200 ;
        RECT 215.800 124.800 216.200 125.200 ;
        RECT 210.200 115.800 210.600 116.200 ;
        RECT 207.800 106.800 208.200 107.200 ;
        RECT 196.600 95.800 197.000 96.200 ;
        RECT 199.800 94.800 200.200 95.200 ;
        RECT 200.600 93.800 201.000 94.200 ;
        RECT 186.200 75.800 186.600 76.200 ;
        RECT 203.000 95.800 203.400 96.200 ;
        RECT 210.200 105.800 210.600 106.200 ;
        RECT 187.000 74.800 187.400 75.200 ;
        RECT 156.600 66.800 157.000 67.200 ;
        RECT 165.400 68.800 165.800 69.200 ;
        RECT 170.200 68.800 170.600 69.200 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 165.400 64.800 165.800 65.200 ;
        RECT 161.400 58.800 161.800 59.200 ;
        RECT 166.200 56.800 166.600 57.200 ;
        RECT 139.800 35.800 140.200 36.200 ;
        RECT 139.800 34.800 140.200 35.200 ;
        RECT 152.600 33.800 153.000 34.200 ;
        RECT 163.800 36.800 164.200 37.200 ;
        RECT 169.400 51.800 169.800 52.200 ;
        RECT 167.000 44.800 167.400 45.200 ;
        RECT 187.800 68.800 188.200 69.200 ;
        RECT 208.600 94.700 209.000 95.100 ;
        RECT 207.000 76.800 207.400 77.200 ;
        RECT 203.000 54.800 203.400 55.200 ;
        RECT 161.400 26.800 161.800 27.200 ;
        RECT 170.200 15.800 170.600 16.200 ;
        RECT 186.200 31.800 186.600 32.200 ;
        RECT 229.400 107.800 229.800 108.200 ;
        RECT 209.400 65.800 209.800 66.200 ;
        RECT 209.400 64.800 209.800 65.200 ;
        RECT 209.400 54.800 209.800 55.200 ;
        RECT 183.000 11.800 183.400 12.200 ;
        RECT 189.400 11.800 189.800 12.200 ;
        RECT 208.600 45.800 209.000 46.200 ;
        RECT 217.400 54.800 217.800 55.200 ;
        RECT 219.800 45.800 220.200 46.200 ;
        RECT 209.400 11.800 209.800 12.200 ;
        RECT 225.400 5.800 225.800 6.200 ;
      LAYER metal3 ;
        RECT 24.600 209.100 25.000 209.200 ;
        RECT 60.600 209.100 61.000 209.200 ;
        RECT 83.800 209.100 84.200 209.200 ;
        RECT 151.800 209.100 152.200 209.200 ;
        RECT 156.600 209.100 157.000 209.200 ;
        RECT 24.600 208.800 116.900 209.100 ;
        RECT 151.800 208.800 157.000 209.100 ;
        RECT 116.600 208.200 116.900 208.800 ;
        RECT 31.800 207.800 32.200 208.200 ;
        RECT 46.200 207.800 46.600 208.200 ;
        RECT 82.200 208.100 82.600 208.200 ;
        RECT 92.600 208.100 93.000 208.200 ;
        RECT 82.200 207.800 93.000 208.100 ;
        RECT 116.600 208.100 117.000 208.200 ;
        RECT 120.600 208.100 121.000 208.200 ;
        RECT 116.600 207.800 121.000 208.100 ;
        RECT 175.000 208.100 175.400 208.200 ;
        RECT 184.600 208.100 185.000 208.200 ;
        RECT 175.000 207.800 185.000 208.100 ;
        RECT 31.800 207.100 32.100 207.800 ;
        RECT 46.200 207.100 46.500 207.800 ;
        RECT 14.200 206.800 46.500 207.100 ;
        RECT 48.600 207.100 49.000 207.200 ;
        RECT 57.400 207.100 57.800 207.200 ;
        RECT 48.600 206.800 57.800 207.100 ;
        RECT 97.400 207.100 97.800 207.200 ;
        RECT 111.000 207.100 111.400 207.200 ;
        RECT 97.400 206.800 102.500 207.100 ;
        RECT 111.000 206.800 117.700 207.100 ;
        RECT 14.200 206.200 14.500 206.800 ;
        RECT 15.800 206.200 16.100 206.800 ;
        RECT 14.200 205.800 14.600 206.200 ;
        RECT 15.800 205.800 16.200 206.200 ;
        RECT 27.800 206.100 28.200 206.200 ;
        RECT 27.800 205.800 28.900 206.100 ;
        RECT 29.400 205.800 29.800 206.200 ;
        RECT 30.200 206.100 30.600 206.200 ;
        RECT 31.000 206.100 31.400 206.200 ;
        RECT 30.200 205.800 31.400 206.100 ;
        RECT 33.400 205.800 33.800 206.200 ;
        RECT 63.800 206.100 64.200 206.200 ;
        RECT 44.600 205.800 64.200 206.100 ;
        RECT 68.600 206.100 69.000 206.200 ;
        RECT 75.000 206.100 75.400 206.200 ;
        RECT 88.600 206.100 89.000 206.200 ;
        RECT 95.000 206.100 95.400 206.300 ;
        RECT 68.600 205.800 75.400 206.100 ;
        RECT 87.800 205.900 95.400 206.100 ;
        RECT 102.200 206.200 102.500 206.800 ;
        RECT 117.400 206.200 117.700 206.800 ;
        RECT 126.200 206.800 126.600 207.200 ;
        RECT 129.400 207.100 129.800 207.200 ;
        RECT 129.400 206.800 143.300 207.100 ;
        RECT 87.800 205.800 95.300 205.900 ;
        RECT 102.200 205.800 102.600 206.200 ;
        RECT 105.400 206.100 105.800 206.200 ;
        RECT 113.400 206.100 113.800 206.200 ;
        RECT 105.400 205.800 113.800 206.100 ;
        RECT 117.400 205.800 117.800 206.200 ;
        RECT 120.600 206.100 121.000 206.200 ;
        RECT 126.200 206.100 126.500 206.800 ;
        RECT 120.600 205.800 126.500 206.100 ;
        RECT 143.000 206.200 143.300 206.800 ;
        RECT 153.400 206.800 153.800 207.200 ;
        RECT 181.400 207.100 181.800 207.200 ;
        RECT 168.600 206.800 181.800 207.100 ;
        RECT 206.200 207.100 206.600 207.200 ;
        RECT 215.000 207.100 215.400 207.200 ;
        RECT 206.200 206.800 215.400 207.100 ;
        RECT 221.400 207.100 221.800 207.200 ;
        RECT 222.200 207.100 222.600 207.200 ;
        RECT 221.400 206.800 222.600 207.100 ;
        RECT 223.000 207.100 223.400 207.200 ;
        RECT 223.800 207.100 224.200 207.200 ;
        RECT 223.000 206.800 224.200 207.100 ;
        RECT 143.000 205.800 143.400 206.200 ;
        RECT 146.200 206.100 146.600 206.200 ;
        RECT 153.400 206.100 153.700 206.800 ;
        RECT 146.200 205.800 153.700 206.100 ;
        RECT 168.600 206.200 168.900 206.800 ;
        RECT 168.600 205.800 169.000 206.200 ;
        RECT 173.400 206.100 173.800 206.200 ;
        RECT 181.400 206.100 181.700 206.800 ;
        RECT 191.000 206.100 191.400 206.200 ;
        RECT 196.600 206.100 197.000 206.200 ;
        RECT 173.400 205.800 178.500 206.100 ;
        RECT 181.400 205.800 197.000 206.100 ;
        RECT 199.000 206.100 199.400 206.200 ;
        RECT 207.800 206.100 208.200 206.200 ;
        RECT 211.000 206.100 211.400 206.200 ;
        RECT 199.000 205.800 211.400 206.100 ;
        RECT 213.400 206.100 213.800 206.200 ;
        RECT 213.400 205.800 224.100 206.100 ;
        RECT 29.400 205.200 29.700 205.800 ;
        RECT 33.400 205.200 33.700 205.800 ;
        RECT 44.600 205.200 44.900 205.800 ;
        RECT 178.200 205.200 178.500 205.800 ;
        RECT 223.800 205.200 224.100 205.800 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 224.600 205.200 224.900 205.800 ;
        RECT 29.400 204.800 29.800 205.200 ;
        RECT 33.400 204.800 33.800 205.200 ;
        RECT 43.000 204.800 43.400 205.200 ;
        RECT 44.600 204.800 45.000 205.200 ;
        RECT 55.000 205.100 55.400 205.200 ;
        RECT 57.400 205.100 57.800 205.200 ;
        RECT 55.000 204.800 57.800 205.100 ;
        RECT 58.200 204.800 58.600 205.200 ;
        RECT 90.200 205.100 90.600 205.200 ;
        RECT 91.000 205.100 91.400 205.200 ;
        RECT 90.200 204.800 91.400 205.100 ;
        RECT 110.200 205.100 110.600 205.200 ;
        RECT 115.800 205.100 116.200 205.200 ;
        RECT 121.400 205.100 121.800 205.200 ;
        RECT 110.200 204.800 114.500 205.100 ;
        RECT 115.800 204.800 121.800 205.100 ;
        RECT 123.000 204.800 123.400 205.200 ;
        RECT 152.600 205.100 153.000 205.200 ;
        RECT 155.000 205.100 155.400 205.200 ;
        RECT 171.000 205.100 171.400 205.200 ;
        RECT 172.600 205.100 173.000 205.200 ;
        RECT 152.600 204.800 173.000 205.100 ;
        RECT 178.200 204.800 178.600 205.200 ;
        RECT 201.400 205.100 201.800 205.200 ;
        RECT 202.200 205.100 202.600 205.200 ;
        RECT 201.400 204.800 202.600 205.100 ;
        RECT 203.800 205.100 204.200 205.200 ;
        RECT 207.000 205.100 207.400 205.200 ;
        RECT 217.400 205.100 217.800 205.200 ;
        RECT 203.800 204.800 217.800 205.100 ;
        RECT 223.800 204.800 224.200 205.200 ;
        RECT 224.600 204.800 225.000 205.200 ;
        RECT 226.200 205.100 226.600 205.200 ;
        RECT 228.600 205.100 229.000 205.200 ;
        RECT 226.200 204.800 229.000 205.100 ;
        RECT 23.000 204.100 23.400 204.200 ;
        RECT 25.400 204.100 25.800 204.200 ;
        RECT 33.400 204.100 33.800 204.200 ;
        RECT 43.000 204.100 43.300 204.800 ;
        RECT 23.000 203.800 43.300 204.100 ;
        RECT 55.000 204.100 55.400 204.200 ;
        RECT 58.200 204.100 58.500 204.800 ;
        RECT 114.200 204.200 114.500 204.800 ;
        RECT 55.000 203.800 58.500 204.100 ;
        RECT 75.800 204.100 76.200 204.200 ;
        RECT 89.400 204.100 89.800 204.200 ;
        RECT 111.000 204.100 111.400 204.200 ;
        RECT 75.800 203.800 111.400 204.100 ;
        RECT 114.200 203.800 114.600 204.200 ;
        RECT 119.800 204.100 120.200 204.200 ;
        RECT 123.000 204.100 123.300 204.800 ;
        RECT 131.800 204.100 132.200 204.200 ;
        RECT 133.400 204.100 133.800 204.200 ;
        RECT 119.800 203.800 121.700 204.100 ;
        RECT 123.000 203.800 133.800 204.100 ;
        RECT 167.000 204.100 167.400 204.200 ;
        RECT 176.600 204.100 177.000 204.200 ;
        RECT 167.000 203.800 177.000 204.100 ;
        RECT 121.400 203.200 121.700 203.800 ;
        RECT 27.000 203.100 27.400 203.200 ;
        RECT 39.000 203.100 39.400 203.200 ;
        RECT 65.400 203.100 65.800 203.200 ;
        RECT 27.000 202.800 65.800 203.100 ;
        RECT 86.200 203.100 86.600 203.200 ;
        RECT 99.800 203.100 100.200 203.200 ;
        RECT 86.200 202.800 100.200 203.100 ;
        RECT 121.400 202.800 121.800 203.200 ;
        RECT 127.800 203.100 128.200 203.200 ;
        RECT 139.000 203.100 139.400 203.200 ;
        RECT 127.800 202.800 139.400 203.100 ;
        RECT 19.800 202.100 20.200 202.200 ;
        RECT 47.800 202.100 48.200 202.200 ;
        RECT 67.000 202.100 67.400 202.200 ;
        RECT 77.400 202.100 77.800 202.200 ;
        RECT 83.800 202.100 84.200 202.200 ;
        RECT 19.800 201.800 24.100 202.100 ;
        RECT 47.800 201.800 84.200 202.100 ;
        RECT 139.800 202.100 140.200 202.200 ;
        RECT 177.400 202.100 177.800 202.200 ;
        RECT 139.800 201.800 177.800 202.100 ;
        RECT 210.200 202.100 210.600 202.200 ;
        RECT 211.000 202.100 211.400 202.200 ;
        RECT 210.200 201.800 211.400 202.100 ;
        RECT 225.400 202.100 225.800 202.200 ;
        RECT 226.200 202.100 226.600 202.200 ;
        RECT 225.400 201.800 226.600 202.100 ;
        RECT 23.800 201.200 24.100 201.800 ;
        RECT 23.800 200.800 24.200 201.200 ;
        RECT 73.400 201.100 73.800 201.200 ;
        RECT 77.400 201.100 77.800 201.200 ;
        RECT 95.800 201.100 96.200 201.200 ;
        RECT 73.400 200.800 96.200 201.100 ;
        RECT 108.600 201.100 109.000 201.200 ;
        RECT 124.600 201.100 125.000 201.200 ;
        RECT 128.600 201.100 129.000 201.200 ;
        RECT 108.600 200.800 129.000 201.100 ;
        RECT 156.600 201.100 157.000 201.200 ;
        RECT 182.200 201.100 182.600 201.200 ;
        RECT 156.600 200.800 182.600 201.100 ;
        RECT 114.200 200.100 114.600 200.200 ;
        RECT 135.000 200.100 135.400 200.200 ;
        RECT 114.200 199.800 135.400 200.100 ;
        RECT 156.600 200.100 157.000 200.200 ;
        RECT 157.400 200.100 157.800 200.200 ;
        RECT 186.200 200.100 186.600 200.200 ;
        RECT 201.400 200.100 201.800 200.200 ;
        RECT 156.600 199.800 201.800 200.100 ;
        RECT 82.200 199.100 82.600 199.200 ;
        RECT 170.200 199.100 170.600 199.200 ;
        RECT 175.800 199.100 176.200 199.200 ;
        RECT 203.000 199.100 203.400 199.200 ;
        RECT 82.200 198.800 203.400 199.100 ;
        RECT 1.400 198.100 1.800 198.200 ;
        RECT 13.400 198.100 13.800 198.200 ;
        RECT 1.400 197.800 13.800 198.100 ;
        RECT 87.800 197.800 88.200 198.200 ;
        RECT 111.000 198.100 111.400 198.200 ;
        RECT 111.800 198.100 112.200 198.200 ;
        RECT 134.200 198.100 134.600 198.200 ;
        RECT 111.000 197.800 134.600 198.100 ;
        RECT 160.600 198.100 161.000 198.200 ;
        RECT 180.600 198.100 181.000 198.200 ;
        RECT 160.600 197.800 181.000 198.100 ;
        RECT 201.400 198.100 201.800 198.200 ;
        RECT 207.800 198.100 208.200 198.200 ;
        RECT 201.400 197.800 208.200 198.100 ;
        RECT 10.200 197.100 10.600 197.200 ;
        RECT 15.800 197.100 16.200 197.200 ;
        RECT 10.200 196.800 16.200 197.100 ;
        RECT 16.600 197.100 17.000 197.200 ;
        RECT 22.200 197.100 22.600 197.200 ;
        RECT 26.200 197.100 26.600 197.200 ;
        RECT 37.400 197.100 37.800 197.200 ;
        RECT 56.600 197.100 57.000 197.200 ;
        RECT 16.600 196.800 22.600 197.100 ;
        RECT 25.400 196.800 57.000 197.100 ;
        RECT 63.800 197.100 64.200 197.200 ;
        RECT 64.600 197.100 65.000 197.200 ;
        RECT 63.800 196.800 65.000 197.100 ;
        RECT 86.200 197.100 86.600 197.200 ;
        RECT 87.800 197.100 88.100 197.800 ;
        RECT 86.200 196.800 88.100 197.100 ;
        RECT 103.800 197.100 104.200 197.200 ;
        RECT 106.200 197.100 106.600 197.200 ;
        RECT 103.800 196.800 106.600 197.100 ;
        RECT 121.400 197.100 121.800 197.200 ;
        RECT 127.000 197.100 127.400 197.200 ;
        RECT 121.400 196.800 128.100 197.100 ;
        RECT 130.200 196.800 130.600 197.200 ;
        RECT 137.400 197.100 137.800 197.200 ;
        RECT 140.600 197.100 141.000 197.200 ;
        RECT 135.800 196.800 141.000 197.100 ;
        RECT 159.000 197.100 159.400 197.200 ;
        RECT 160.600 197.100 161.000 197.200 ;
        RECT 159.000 196.800 161.000 197.100 ;
        RECT 7.000 195.800 7.400 196.200 ;
        RECT 12.600 196.100 13.000 196.200 ;
        RECT 30.200 196.100 30.600 196.200 ;
        RECT 12.600 195.800 30.600 196.100 ;
        RECT 49.400 196.100 49.800 196.200 ;
        RECT 50.200 196.100 50.600 196.200 ;
        RECT 49.400 195.800 50.600 196.100 ;
        RECT 59.800 196.100 60.200 196.200 ;
        RECT 66.200 196.100 66.600 196.200 ;
        RECT 79.000 196.100 79.400 196.200 ;
        RECT 84.600 196.100 85.000 196.200 ;
        RECT 87.000 196.100 87.400 196.200 ;
        RECT 90.200 196.100 90.600 196.200 ;
        RECT 59.800 195.800 66.600 196.100 ;
        RECT 71.000 195.800 90.600 196.100 ;
        RECT 102.200 196.100 102.600 196.200 ;
        RECT 126.200 196.100 126.600 196.200 ;
        RECT 130.200 196.100 130.500 196.800 ;
        RECT 102.200 195.800 122.500 196.100 ;
        RECT 126.200 195.800 130.500 196.100 ;
        RECT 135.800 196.200 136.100 196.800 ;
        RECT 135.800 195.800 136.200 196.200 ;
        RECT 139.000 196.100 139.400 196.200 ;
        RECT 147.000 196.100 147.400 196.200 ;
        RECT 138.200 195.800 147.400 196.100 ;
        RECT 151.800 196.100 152.200 196.200 ;
        RECT 160.600 196.100 161.000 196.200 ;
        RECT 151.800 195.800 161.000 196.100 ;
        RECT 161.400 196.100 161.800 196.200 ;
        RECT 163.800 196.100 164.200 196.200 ;
        RECT 164.600 196.100 165.000 196.200 ;
        RECT 161.400 195.800 165.000 196.100 ;
        RECT 184.600 196.100 185.000 196.200 ;
        RECT 192.600 196.100 193.000 196.200 ;
        RECT 184.600 195.800 193.000 196.100 ;
        RECT 196.600 196.100 197.000 196.200 ;
        RECT 211.800 196.100 212.200 196.200 ;
        RECT 196.600 195.800 212.200 196.100 ;
        RECT 224.600 195.800 225.000 196.200 ;
        RECT 7.000 195.100 7.300 195.800 ;
        RECT 71.000 195.200 71.300 195.800 ;
        RECT 122.200 195.200 122.500 195.800 ;
        RECT 11.000 195.100 11.400 195.200 ;
        RECT 7.000 194.800 11.400 195.100 ;
        RECT 15.800 195.100 16.200 195.200 ;
        RECT 23.000 195.100 23.400 195.200 ;
        RECT 15.800 194.800 23.400 195.100 ;
        RECT 28.600 195.100 29.000 195.200 ;
        RECT 51.000 195.100 51.400 195.200 ;
        RECT 51.800 195.100 52.200 195.200 ;
        RECT 55.800 195.100 56.200 195.200 ;
        RECT 28.600 194.800 56.200 195.100 ;
        RECT 57.400 195.100 57.800 195.200 ;
        RECT 58.200 195.100 58.600 195.200 ;
        RECT 57.400 194.800 58.600 195.100 ;
        RECT 59.000 194.800 59.400 195.200 ;
        RECT 62.200 195.100 62.600 195.200 ;
        RECT 71.000 195.100 71.400 195.200 ;
        RECT 62.200 194.800 71.400 195.100 ;
        RECT 72.600 194.800 73.000 195.200 ;
        RECT 75.800 195.100 76.200 195.200 ;
        RECT 76.600 195.100 77.000 195.200 ;
        RECT 85.400 195.100 85.800 195.200 ;
        RECT 90.200 195.100 90.600 195.200 ;
        RECT 120.600 195.100 121.000 195.200 ;
        RECT 75.800 194.800 121.000 195.100 ;
        RECT 122.200 195.100 122.600 195.200 ;
        RECT 127.000 195.100 127.400 195.200 ;
        RECT 122.200 194.800 127.400 195.100 ;
        RECT 134.200 195.100 134.600 195.200 ;
        RECT 139.000 195.100 139.400 195.200 ;
        RECT 147.800 195.100 148.200 195.200 ;
        RECT 151.800 195.100 152.200 195.200 ;
        RECT 134.200 194.800 152.200 195.100 ;
        RECT 159.000 194.800 159.400 195.200 ;
        RECT 163.000 195.100 163.400 195.200 ;
        RECT 170.200 195.100 170.600 195.200 ;
        RECT 163.000 194.800 170.600 195.100 ;
        RECT 179.000 195.100 179.400 195.200 ;
        RECT 186.200 195.100 186.600 195.200 ;
        RECT 189.400 195.100 189.800 195.200 ;
        RECT 179.000 194.800 189.800 195.100 ;
        RECT 204.600 195.100 205.000 195.200 ;
        RECT 206.200 195.100 206.600 195.200 ;
        RECT 204.600 194.800 206.600 195.100 ;
        RECT 216.600 195.100 217.000 195.200 ;
        RECT 224.600 195.100 224.900 195.800 ;
        RECT 216.600 194.800 224.900 195.100 ;
        RECT 59.000 194.200 59.300 194.800 ;
        RECT 16.600 194.100 17.000 194.200 ;
        RECT 24.600 194.100 25.000 194.200 ;
        RECT 16.600 193.800 25.000 194.100 ;
        RECT 26.200 194.100 26.600 194.200 ;
        RECT 31.800 194.100 32.200 194.200 ;
        RECT 26.200 193.800 32.200 194.100 ;
        RECT 45.400 194.100 45.800 194.200 ;
        RECT 51.000 194.100 51.400 194.200 ;
        RECT 45.400 193.800 51.400 194.100 ;
        RECT 52.600 194.100 53.000 194.200 ;
        RECT 57.400 194.100 57.800 194.200 ;
        RECT 52.600 193.800 57.800 194.100 ;
        RECT 59.000 193.800 59.400 194.200 ;
        RECT 59.800 194.100 60.200 194.200 ;
        RECT 63.800 194.100 64.200 194.200 ;
        RECT 59.800 193.800 64.200 194.100 ;
        RECT 71.000 194.100 71.400 194.200 ;
        RECT 71.800 194.100 72.200 194.200 ;
        RECT 71.000 193.800 72.200 194.100 ;
        RECT 72.600 194.100 72.900 194.800 ;
        RECT 80.600 194.100 81.000 194.200 ;
        RECT 72.600 193.800 81.000 194.100 ;
        RECT 85.400 194.100 85.800 194.200 ;
        RECT 94.200 194.100 94.600 194.200 ;
        RECT 85.400 193.800 94.600 194.100 ;
        RECT 102.200 193.800 102.600 194.200 ;
        RECT 110.200 194.100 110.600 194.200 ;
        RECT 103.800 193.800 110.600 194.100 ;
        RECT 115.800 194.100 116.200 194.200 ;
        RECT 116.600 194.100 117.000 194.200 ;
        RECT 115.800 193.800 117.000 194.100 ;
        RECT 118.200 194.100 118.600 194.200 ;
        RECT 141.400 194.100 141.800 194.200 ;
        RECT 118.200 193.800 141.800 194.100 ;
        RECT 159.000 194.100 159.300 194.800 ;
        RECT 171.000 194.100 171.400 194.200 ;
        RECT 159.000 193.800 171.400 194.100 ;
        RECT 185.400 193.800 185.800 194.200 ;
        RECT 188.600 194.100 189.000 194.200 ;
        RECT 199.000 194.100 199.400 194.200 ;
        RECT 188.600 193.800 199.400 194.100 ;
        RECT 204.600 194.100 205.000 194.200 ;
        RECT 214.200 194.100 214.600 194.200 ;
        RECT 204.600 193.800 214.600 194.100 ;
        RECT 102.200 193.200 102.500 193.800 ;
        RECT 103.800 193.200 104.100 193.800 ;
        RECT 185.400 193.200 185.700 193.800 ;
        RECT 6.200 193.100 6.600 193.200 ;
        RECT 41.400 193.100 41.800 193.200 ;
        RECT 6.200 192.800 41.800 193.100 ;
        RECT 50.200 193.100 50.600 193.200 ;
        RECT 58.200 193.100 58.600 193.200 ;
        RECT 50.200 192.800 58.600 193.100 ;
        RECT 102.200 192.800 102.600 193.200 ;
        RECT 103.800 192.800 104.200 193.200 ;
        RECT 104.600 193.100 105.000 193.200 ;
        RECT 115.800 193.100 116.200 193.200 ;
        RECT 104.600 192.800 116.200 193.100 ;
        RECT 127.000 193.100 127.400 193.200 ;
        RECT 139.000 193.100 139.400 193.200 ;
        RECT 127.000 192.800 139.400 193.100 ;
        RECT 155.800 193.100 156.200 193.200 ;
        RECT 176.600 193.100 177.000 193.200 ;
        RECT 179.000 193.100 179.400 193.200 ;
        RECT 155.800 192.800 179.400 193.100 ;
        RECT 185.400 192.800 185.800 193.200 ;
        RECT 11.800 192.100 12.200 192.200 ;
        RECT 18.200 192.100 18.600 192.200 ;
        RECT 19.000 192.100 19.400 192.200 ;
        RECT 11.800 191.800 19.400 192.100 ;
        RECT 27.000 192.100 27.400 192.200 ;
        RECT 29.400 192.100 29.800 192.200 ;
        RECT 27.000 191.800 29.800 192.100 ;
        RECT 46.200 192.100 46.600 192.200 ;
        RECT 62.200 192.100 62.600 192.200 ;
        RECT 46.200 191.800 62.600 192.100 ;
        RECT 87.800 192.100 88.200 192.200 ;
        RECT 105.400 192.100 105.800 192.200 ;
        RECT 87.800 191.800 105.800 192.100 ;
        RECT 107.000 192.100 107.400 192.200 ;
        RECT 116.600 192.100 117.000 192.200 ;
        RECT 107.000 191.800 117.000 192.100 ;
        RECT 181.400 192.100 181.800 192.200 ;
        RECT 186.200 192.100 186.600 192.200 ;
        RECT 181.400 191.800 186.600 192.100 ;
        RECT 219.000 192.100 219.400 192.200 ;
        RECT 219.000 191.800 220.900 192.100 ;
        RECT 220.600 191.200 220.900 191.800 ;
        RECT 19.000 191.100 19.400 191.200 ;
        RECT 26.200 191.100 26.600 191.200 ;
        RECT 28.600 191.100 29.000 191.200 ;
        RECT 36.600 191.100 37.000 191.200 ;
        RECT 74.200 191.100 74.600 191.200 ;
        RECT 19.000 190.800 74.600 191.100 ;
        RECT 98.200 191.100 98.600 191.200 ;
        RECT 99.800 191.100 100.200 191.200 ;
        RECT 98.200 190.800 100.200 191.100 ;
        RECT 114.200 191.100 114.600 191.200 ;
        RECT 115.800 191.100 116.200 191.200 ;
        RECT 131.800 191.100 132.200 191.200 ;
        RECT 141.400 191.100 141.800 191.200 ;
        RECT 143.800 191.100 144.200 191.200 ;
        RECT 114.200 190.800 144.200 191.100 ;
        RECT 220.600 190.800 221.000 191.200 ;
        RECT 23.000 190.100 23.400 190.200 ;
        RECT 32.600 190.100 33.000 190.200 ;
        RECT 80.600 190.100 81.000 190.200 ;
        RECT 23.000 189.800 81.000 190.100 ;
        RECT 91.000 190.100 91.400 190.200 ;
        RECT 100.600 190.100 101.000 190.200 ;
        RECT 104.600 190.100 105.000 190.200 ;
        RECT 91.000 189.800 105.000 190.100 ;
        RECT 106.200 190.100 106.600 190.200 ;
        RECT 118.200 190.100 118.600 190.200 ;
        RECT 106.200 189.800 118.600 190.100 ;
        RECT 121.400 190.100 121.800 190.200 ;
        RECT 147.000 190.100 147.400 190.200 ;
        RECT 121.400 189.800 147.400 190.100 ;
        RECT 183.000 190.100 183.400 190.200 ;
        RECT 186.200 190.100 186.600 190.200 ;
        RECT 183.000 189.800 186.600 190.100 ;
        RECT 207.000 190.100 207.400 190.200 ;
        RECT 221.400 190.100 221.800 190.200 ;
        RECT 223.000 190.100 223.400 190.200 ;
        RECT 207.000 189.800 223.400 190.100 ;
        RECT 80.600 189.100 81.000 189.200 ;
        RECT 132.600 189.100 133.000 189.200 ;
        RECT 80.600 188.800 133.000 189.100 ;
        RECT 152.600 188.800 153.000 189.200 ;
        RECT 157.400 189.100 157.800 189.200 ;
        RECT 161.400 189.100 161.800 189.200 ;
        RECT 217.400 189.100 217.800 189.200 ;
        RECT 157.400 188.800 161.800 189.100 ;
        RECT 207.800 188.800 217.800 189.100 ;
        RECT 19.800 188.100 20.200 188.200 ;
        RECT 27.800 188.100 28.200 188.200 ;
        RECT 19.800 187.800 28.200 188.100 ;
        RECT 66.200 188.100 66.600 188.200 ;
        RECT 70.200 188.100 70.600 188.200 ;
        RECT 66.200 187.800 70.600 188.100 ;
        RECT 103.800 188.100 104.200 188.200 ;
        RECT 109.400 188.100 109.800 188.200 ;
        RECT 115.800 188.100 116.200 188.200 ;
        RECT 103.800 187.800 116.200 188.100 ;
        RECT 132.600 188.100 132.900 188.800 ;
        RECT 140.600 188.100 141.000 188.200 ;
        RECT 132.600 187.800 141.000 188.100 ;
        RECT 149.400 188.100 149.800 188.200 ;
        RECT 152.600 188.100 152.900 188.800 ;
        RECT 207.800 188.200 208.100 188.800 ;
        RECT 149.400 187.800 152.900 188.100 ;
        RECT 173.400 188.100 173.800 188.200 ;
        RECT 175.000 188.100 175.400 188.200 ;
        RECT 173.400 187.800 175.400 188.100 ;
        RECT 176.600 187.800 177.000 188.200 ;
        RECT 178.200 188.100 178.600 188.200 ;
        RECT 179.000 188.100 179.400 188.200 ;
        RECT 178.200 187.800 179.400 188.100 ;
        RECT 183.800 188.100 184.200 188.200 ;
        RECT 187.800 188.100 188.200 188.200 ;
        RECT 183.800 187.800 188.200 188.100 ;
        RECT 203.800 188.100 204.200 188.200 ;
        RECT 207.800 188.100 208.200 188.200 ;
        RECT 203.800 187.800 208.200 188.100 ;
        RECT 13.400 187.100 13.800 187.200 ;
        RECT 38.200 187.100 38.600 187.200 ;
        RECT 13.400 186.800 38.600 187.100 ;
        RECT 58.200 187.100 58.600 187.200 ;
        RECT 61.400 187.100 61.800 187.200 ;
        RECT 69.400 187.100 69.800 187.200 ;
        RECT 71.000 187.100 71.400 187.200 ;
        RECT 58.200 186.800 71.400 187.100 ;
        RECT 74.200 187.100 74.600 187.200 ;
        RECT 127.000 187.100 127.400 187.200 ;
        RECT 152.600 187.100 153.000 187.200 ;
        RECT 74.200 186.800 127.400 187.100 ;
        RECT 149.400 186.800 153.000 187.100 ;
        RECT 159.000 187.100 159.400 187.200 ;
        RECT 160.600 187.100 161.000 187.200 ;
        RECT 163.800 187.100 164.200 187.200 ;
        RECT 159.000 186.800 164.200 187.100 ;
        RECT 167.800 187.100 168.200 187.200 ;
        RECT 176.600 187.100 176.900 187.800 ;
        RECT 167.800 186.800 176.900 187.100 ;
        RECT 180.600 187.100 181.000 187.200 ;
        RECT 183.000 187.100 183.400 187.200 ;
        RECT 180.600 186.800 183.400 187.100 ;
        RECT 184.600 187.100 185.000 187.200 ;
        RECT 194.200 187.100 194.600 187.200 ;
        RECT 184.600 186.800 194.600 187.100 ;
        RECT 196.600 187.100 197.000 187.200 ;
        RECT 199.800 187.100 200.200 187.200 ;
        RECT 196.600 186.800 200.200 187.100 ;
        RECT 201.400 187.100 201.800 187.200 ;
        RECT 204.600 187.100 205.000 187.200 ;
        RECT 201.400 186.800 205.000 187.100 ;
        RECT 214.200 186.800 214.600 187.200 ;
        RECT 222.200 187.100 222.600 187.200 ;
        RECT 227.000 187.100 227.400 187.200 ;
        RECT 222.200 186.800 227.400 187.100 ;
        RECT 149.400 186.200 149.700 186.800 ;
        RECT 5.400 186.100 5.800 186.200 ;
        RECT 10.200 186.100 10.600 186.200 ;
        RECT 5.400 185.800 10.600 186.100 ;
        RECT 11.000 186.100 11.400 186.200 ;
        RECT 11.800 186.100 12.200 186.200 ;
        RECT 11.000 185.800 12.200 186.100 ;
        RECT 23.800 186.100 24.200 186.200 ;
        RECT 39.800 186.100 40.200 186.200 ;
        RECT 47.800 186.100 48.200 186.200 ;
        RECT 54.200 186.100 54.600 186.200 ;
        RECT 23.800 185.800 40.200 186.100 ;
        RECT 47.000 185.800 54.600 186.100 ;
        RECT 55.800 186.100 56.200 186.200 ;
        RECT 63.000 186.100 63.400 186.200 ;
        RECT 55.800 185.800 63.400 186.100 ;
        RECT 63.800 186.100 64.200 186.200 ;
        RECT 68.600 186.100 69.000 186.200 ;
        RECT 63.800 185.800 69.000 186.100 ;
        RECT 75.000 186.100 75.400 186.200 ;
        RECT 77.400 186.100 77.800 186.200 ;
        RECT 87.000 186.100 87.400 186.200 ;
        RECT 75.000 185.800 87.400 186.100 ;
        RECT 87.800 186.100 88.200 186.200 ;
        RECT 91.800 186.100 92.200 186.200 ;
        RECT 87.800 185.800 92.200 186.100 ;
        RECT 94.200 186.100 94.600 186.200 ;
        RECT 95.000 186.100 95.400 186.200 ;
        RECT 94.200 185.800 95.400 186.100 ;
        RECT 99.000 186.100 99.400 186.200 ;
        RECT 101.400 186.100 101.800 186.200 ;
        RECT 99.000 185.800 101.800 186.100 ;
        RECT 118.200 185.800 118.600 186.200 ;
        RECT 119.000 186.100 119.400 186.200 ;
        RECT 126.200 186.100 126.600 186.200 ;
        RECT 119.000 185.800 126.600 186.100 ;
        RECT 139.800 186.100 140.200 186.200 ;
        RECT 147.000 186.100 147.400 186.200 ;
        RECT 139.800 185.800 147.400 186.100 ;
        RECT 149.400 185.800 149.800 186.200 ;
        RECT 151.000 186.100 151.400 186.200 ;
        RECT 159.800 186.100 160.200 186.200 ;
        RECT 151.000 185.800 160.200 186.100 ;
        RECT 161.400 186.100 161.800 186.200 ;
        RECT 163.000 186.100 163.400 186.200 ;
        RECT 178.200 186.100 178.600 186.200 ;
        RECT 179.800 186.100 180.200 186.200 ;
        RECT 161.400 185.800 180.200 186.100 ;
        RECT 185.400 186.100 185.800 186.200 ;
        RECT 202.200 186.100 202.600 186.200 ;
        RECT 185.400 185.800 202.600 186.100 ;
        RECT 214.200 186.100 214.500 186.800 ;
        RECT 219.000 186.100 219.400 186.200 ;
        RECT 214.200 185.800 219.400 186.100 ;
        RECT 11.000 185.100 11.400 185.200 ;
        RECT 12.600 185.100 13.000 185.200 ;
        RECT 11.000 184.800 13.000 185.100 ;
        RECT 13.400 184.800 13.800 185.200 ;
        RECT 29.400 184.800 29.800 185.200 ;
        RECT 49.400 185.100 49.800 185.200 ;
        RECT 59.000 185.100 59.400 185.200 ;
        RECT 60.600 185.100 61.000 185.200 ;
        RECT 49.400 184.800 61.000 185.100 ;
        RECT 62.200 185.100 62.600 185.200 ;
        RECT 64.600 185.100 65.000 185.200 ;
        RECT 62.200 184.800 65.000 185.100 ;
        RECT 76.600 185.100 77.000 185.200 ;
        RECT 105.400 185.100 105.800 185.200 ;
        RECT 76.600 184.800 105.800 185.100 ;
        RECT 107.800 185.100 108.200 185.200 ;
        RECT 118.200 185.100 118.500 185.800 ;
        RECT 122.200 185.100 122.600 185.200 ;
        RECT 107.800 184.800 122.600 185.100 ;
        RECT 134.200 185.100 134.600 185.200 ;
        RECT 145.400 185.100 145.800 185.200 ;
        RECT 134.200 184.800 145.800 185.100 ;
        RECT 147.000 185.100 147.400 185.200 ;
        RECT 148.600 185.100 149.000 185.200 ;
        RECT 147.000 184.800 149.000 185.100 ;
        RECT 187.000 185.100 187.400 185.200 ;
        RECT 193.400 185.100 193.800 185.200 ;
        RECT 198.200 185.100 198.600 185.200 ;
        RECT 187.000 184.800 198.600 185.100 ;
        RECT 225.400 185.100 225.800 185.200 ;
        RECT 227.000 185.100 227.400 185.200 ;
        RECT 225.400 184.800 227.400 185.100 ;
        RECT 10.200 184.100 10.600 184.200 ;
        RECT 13.400 184.100 13.700 184.800 ;
        RECT 10.200 183.800 13.700 184.100 ;
        RECT 26.200 184.100 26.600 184.200 ;
        RECT 29.400 184.100 29.700 184.800 ;
        RECT 67.000 184.100 67.400 184.200 ;
        RECT 26.200 183.800 67.400 184.100 ;
        RECT 75.800 184.100 76.200 184.200 ;
        RECT 82.200 184.100 82.600 184.200 ;
        RECT 75.800 183.800 82.600 184.100 ;
        RECT 83.800 184.100 84.200 184.200 ;
        RECT 87.800 184.100 88.200 184.200 ;
        RECT 91.800 184.100 92.200 184.200 ;
        RECT 83.800 183.800 88.200 184.100 ;
        RECT 88.600 183.800 92.200 184.100 ;
        RECT 95.000 184.100 95.400 184.200 ;
        RECT 95.800 184.100 96.200 184.200 ;
        RECT 95.000 183.800 96.200 184.100 ;
        RECT 146.200 184.100 146.600 184.200 ;
        RECT 158.200 184.100 158.600 184.200 ;
        RECT 146.200 183.800 158.600 184.100 ;
        RECT 186.200 184.100 186.600 184.200 ;
        RECT 206.200 184.100 206.600 184.200 ;
        RECT 219.000 184.100 219.400 184.200 ;
        RECT 221.400 184.100 221.800 184.200 ;
        RECT 186.200 183.800 221.800 184.100 ;
        RECT 88.600 183.200 88.900 183.800 ;
        RECT 35.800 183.100 36.200 183.200 ;
        RECT 52.600 183.100 53.000 183.200 ;
        RECT 35.800 182.800 53.000 183.100 ;
        RECT 55.800 183.100 56.200 183.200 ;
        RECT 56.600 183.100 57.000 183.200 ;
        RECT 59.800 183.100 60.200 183.200 ;
        RECT 67.800 183.100 68.200 183.200 ;
        RECT 55.800 182.800 68.200 183.100 ;
        RECT 88.600 182.800 89.000 183.200 ;
        RECT 101.400 183.100 101.800 183.200 ;
        RECT 151.800 183.100 152.200 183.200 ;
        RECT 101.400 182.800 152.200 183.100 ;
        RECT 41.400 182.100 41.800 182.200 ;
        RECT 43.000 182.100 43.400 182.200 ;
        RECT 63.800 182.100 64.200 182.200 ;
        RECT 108.600 182.100 109.000 182.200 ;
        RECT 153.400 182.100 153.800 182.200 ;
        RECT 41.400 181.800 153.800 182.100 ;
        RECT 155.000 182.100 155.400 182.200 ;
        RECT 182.200 182.100 182.600 182.200 ;
        RECT 188.600 182.100 189.000 182.200 ;
        RECT 155.000 181.800 189.000 182.100 ;
        RECT 218.200 182.100 218.600 182.200 ;
        RECT 230.200 182.100 230.600 182.200 ;
        RECT 218.200 181.800 230.600 182.100 ;
        RECT 51.800 181.100 52.200 181.200 ;
        RECT 87.000 181.100 87.400 181.200 ;
        RECT 51.800 180.800 87.400 181.100 ;
        RECT 155.000 181.100 155.400 181.200 ;
        RECT 159.000 181.100 159.400 181.200 ;
        RECT 155.000 180.800 159.400 181.100 ;
        RECT 175.800 181.100 176.200 181.200 ;
        RECT 199.000 181.100 199.400 181.200 ;
        RECT 175.800 180.800 199.400 181.100 ;
        RECT 220.600 181.100 221.000 181.200 ;
        RECT 222.200 181.100 222.600 181.200 ;
        RECT 220.600 180.800 222.600 181.100 ;
        RECT 33.400 180.100 33.800 180.200 ;
        RECT 34.200 180.100 34.600 180.200 ;
        RECT 33.400 179.800 34.600 180.100 ;
        RECT 51.000 180.100 51.400 180.200 ;
        RECT 55.000 180.100 55.400 180.200 ;
        RECT 51.000 179.800 55.400 180.100 ;
        RECT 61.400 180.100 61.800 180.200 ;
        RECT 69.400 180.100 69.800 180.200 ;
        RECT 61.400 179.800 69.800 180.100 ;
        RECT 82.200 180.100 82.600 180.200 ;
        RECT 93.400 180.100 93.800 180.200 ;
        RECT 82.200 179.800 93.800 180.100 ;
        RECT 98.200 180.100 98.600 180.200 ;
        RECT 116.600 180.100 117.000 180.200 ;
        RECT 98.200 179.800 117.000 180.100 ;
        RECT 155.000 180.100 155.400 180.200 ;
        RECT 165.400 180.100 165.800 180.200 ;
        RECT 155.000 179.800 165.800 180.100 ;
        RECT 34.200 179.100 34.600 179.200 ;
        RECT 35.000 179.100 35.400 179.200 ;
        RECT 42.200 179.100 42.600 179.200 ;
        RECT 34.200 178.800 42.600 179.100 ;
        RECT 68.600 179.100 69.000 179.200 ;
        RECT 98.200 179.100 98.600 179.200 ;
        RECT 111.800 179.100 112.200 179.200 ;
        RECT 68.600 178.800 112.200 179.100 ;
        RECT 116.600 179.100 116.900 179.800 ;
        RECT 144.600 179.100 145.000 179.200 ;
        RECT 116.600 178.800 145.000 179.100 ;
        RECT 160.600 179.100 161.000 179.200 ;
        RECT 161.400 179.100 161.800 179.200 ;
        RECT 160.600 178.800 161.800 179.100 ;
        RECT 183.000 179.100 183.400 179.200 ;
        RECT 199.800 179.100 200.200 179.200 ;
        RECT 183.000 178.800 200.200 179.100 ;
        RECT 13.400 178.100 13.800 178.200 ;
        RECT 39.800 178.100 40.200 178.200 ;
        RECT 13.400 177.800 40.200 178.100 ;
        RECT 66.200 178.100 66.600 178.200 ;
        RECT 67.000 178.100 67.400 178.200 ;
        RECT 66.200 177.800 67.400 178.100 ;
        RECT 69.400 178.100 69.800 178.200 ;
        RECT 85.400 178.100 85.800 178.200 ;
        RECT 99.800 178.100 100.200 178.200 ;
        RECT 107.000 178.100 107.400 178.200 ;
        RECT 69.400 177.800 107.400 178.100 ;
        RECT 108.600 178.100 109.000 178.200 ;
        RECT 111.000 178.100 111.400 178.200 ;
        RECT 108.600 177.800 111.400 178.100 ;
        RECT 136.600 178.100 137.000 178.200 ;
        RECT 143.000 178.100 143.400 178.200 ;
        RECT 136.600 177.800 143.400 178.100 ;
        RECT 194.200 178.100 194.600 178.200 ;
        RECT 215.000 178.100 215.400 178.200 ;
        RECT 225.400 178.100 225.800 178.200 ;
        RECT 194.200 177.800 225.800 178.100 ;
        RECT 11.800 177.100 12.200 177.200 ;
        RECT 35.800 177.100 36.200 177.200 ;
        RECT 11.800 176.800 36.200 177.100 ;
        RECT 57.400 177.100 57.800 177.200 ;
        RECT 59.000 177.100 59.400 177.200 ;
        RECT 57.400 176.800 59.400 177.100 ;
        RECT 82.200 177.100 82.600 177.200 ;
        RECT 88.600 177.100 89.000 177.200 ;
        RECT 124.600 177.100 125.000 177.200 ;
        RECT 82.200 176.800 89.000 177.100 ;
        RECT 115.800 176.800 125.000 177.100 ;
        RECT 163.000 177.100 163.400 177.200 ;
        RECT 171.800 177.100 172.200 177.200 ;
        RECT 176.600 177.100 177.000 177.200 ;
        RECT 163.000 176.800 177.000 177.100 ;
        RECT 185.400 177.100 185.800 177.200 ;
        RECT 195.000 177.100 195.400 177.200 ;
        RECT 185.400 176.800 195.400 177.100 ;
        RECT 198.200 177.100 198.600 177.200 ;
        RECT 204.600 177.100 205.000 177.200 ;
        RECT 198.200 176.800 205.000 177.100 ;
        RECT 209.400 177.100 209.800 177.200 ;
        RECT 210.200 177.100 210.600 177.200 ;
        RECT 209.400 176.800 210.600 177.100 ;
        RECT 115.800 176.200 116.100 176.800 ;
        RECT 33.400 176.100 33.800 176.200 ;
        RECT 34.200 176.100 34.600 176.200 ;
        RECT 33.400 175.800 34.600 176.100 ;
        RECT 52.600 176.100 53.000 176.200 ;
        RECT 57.400 176.100 57.800 176.200 ;
        RECT 63.000 176.100 63.400 176.200 ;
        RECT 52.600 175.800 63.400 176.100 ;
        RECT 66.200 175.800 66.600 176.200 ;
        RECT 70.200 175.800 70.600 176.200 ;
        RECT 86.200 176.100 86.600 176.200 ;
        RECT 92.600 176.100 93.000 176.200 ;
        RECT 95.800 176.100 96.200 176.200 ;
        RECT 86.200 175.800 96.200 176.100 ;
        RECT 113.400 176.100 113.800 176.200 ;
        RECT 115.000 176.100 115.400 176.200 ;
        RECT 113.400 175.800 115.400 176.100 ;
        RECT 115.800 175.800 116.200 176.200 ;
        RECT 142.200 176.100 142.600 176.200 ;
        RECT 147.800 176.100 148.200 176.200 ;
        RECT 142.200 175.800 148.200 176.100 ;
        RECT 179.800 176.100 180.200 176.200 ;
        RECT 189.400 176.100 189.800 176.200 ;
        RECT 179.800 175.800 189.800 176.100 ;
        RECT 199.000 175.800 199.400 176.200 ;
        RECT 203.000 176.100 203.400 176.200 ;
        RECT 208.600 176.100 209.000 176.200 ;
        RECT 203.000 175.800 209.000 176.100 ;
        RECT 210.200 175.800 210.600 176.200 ;
        RECT 215.000 175.800 215.400 176.200 ;
        RECT 217.400 176.100 217.800 176.200 ;
        RECT 226.200 176.100 226.600 176.200 ;
        RECT 229.400 176.100 229.800 176.200 ;
        RECT 217.400 175.800 229.800 176.100 ;
        RECT 6.200 175.100 6.600 175.200 ;
        RECT 6.200 174.800 11.300 175.100 ;
        RECT 11.000 174.200 11.300 174.800 ;
        RECT 25.400 174.800 25.800 175.200 ;
        RECT 29.400 175.100 29.800 175.200 ;
        RECT 35.000 175.100 35.400 175.200 ;
        RECT 29.400 174.800 35.400 175.100 ;
        RECT 48.600 175.100 49.000 175.200 ;
        RECT 55.800 175.100 56.200 175.200 ;
        RECT 48.600 174.800 56.200 175.100 ;
        RECT 59.800 174.800 60.200 175.200 ;
        RECT 66.200 175.100 66.500 175.800 ;
        RECT 70.200 175.100 70.500 175.800 ;
        RECT 106.200 175.100 106.600 175.200 ;
        RECT 66.200 174.800 70.500 175.100 ;
        RECT 87.800 174.800 106.600 175.100 ;
        RECT 110.200 174.800 110.600 175.200 ;
        RECT 112.600 175.100 113.000 175.200 ;
        RECT 123.000 175.100 123.400 175.200 ;
        RECT 154.200 175.100 154.600 175.200 ;
        RECT 155.800 175.100 156.200 175.200 ;
        RECT 112.600 174.800 119.300 175.100 ;
        RECT 123.000 174.800 156.200 175.100 ;
        RECT 158.200 174.800 158.600 175.200 ;
        RECT 159.000 175.100 159.400 175.200 ;
        RECT 161.400 175.100 161.800 175.200 ;
        RECT 159.000 174.800 161.800 175.100 ;
        RECT 183.000 175.100 183.400 175.200 ;
        RECT 186.200 175.100 186.600 175.200 ;
        RECT 183.000 174.800 186.600 175.100 ;
        RECT 187.800 175.100 188.200 175.200 ;
        RECT 195.000 175.100 195.400 175.200 ;
        RECT 199.000 175.100 199.300 175.800 ;
        RECT 187.800 174.800 189.700 175.100 ;
        RECT 195.000 174.800 199.300 175.100 ;
        RECT 201.400 175.100 201.800 175.200 ;
        RECT 207.000 175.100 207.400 175.200 ;
        RECT 210.200 175.100 210.500 175.800 ;
        RECT 201.400 174.800 210.500 175.100 ;
        RECT 215.000 175.200 215.300 175.800 ;
        RECT 215.000 174.800 215.400 175.200 ;
        RECT 221.400 175.100 221.800 175.200 ;
        RECT 227.800 175.100 228.200 175.200 ;
        RECT 221.400 174.800 228.200 175.100 ;
        RECT 11.000 174.100 11.400 174.200 ;
        RECT 22.200 174.100 22.600 174.200 ;
        RECT 25.400 174.100 25.700 174.800 ;
        RECT 59.800 174.200 60.100 174.800 ;
        RECT 87.800 174.200 88.100 174.800 ;
        RECT 11.000 173.800 25.700 174.100 ;
        RECT 35.800 174.100 36.200 174.200 ;
        RECT 51.800 174.100 52.200 174.200 ;
        RECT 54.200 174.100 54.600 174.200 ;
        RECT 35.800 173.800 54.600 174.100 ;
        RECT 59.800 173.800 60.200 174.200 ;
        RECT 66.200 174.100 66.600 174.200 ;
        RECT 67.000 174.100 67.400 174.200 ;
        RECT 66.200 173.800 67.400 174.100 ;
        RECT 68.600 174.100 69.000 174.200 ;
        RECT 71.000 174.100 71.400 174.200 ;
        RECT 68.600 173.800 71.400 174.100 ;
        RECT 87.800 173.800 88.200 174.200 ;
        RECT 89.400 174.100 89.800 174.200 ;
        RECT 93.400 174.100 93.800 174.200 ;
        RECT 98.200 174.100 98.600 174.200 ;
        RECT 89.400 173.800 98.600 174.100 ;
        RECT 100.600 174.100 101.000 174.200 ;
        RECT 110.200 174.100 110.500 174.800 ;
        RECT 100.600 173.800 110.500 174.100 ;
        RECT 119.000 174.200 119.300 174.800 ;
        RECT 119.000 173.800 119.400 174.200 ;
        RECT 129.400 174.100 129.800 174.200 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 138.200 174.100 138.600 174.200 ;
        RECT 129.400 173.800 130.600 174.100 ;
        RECT 131.800 173.800 138.600 174.100 ;
        RECT 139.000 174.100 139.400 174.200 ;
        RECT 141.400 174.100 141.800 174.200 ;
        RECT 153.400 174.100 153.800 174.200 ;
        RECT 158.200 174.100 158.500 174.800 ;
        RECT 189.400 174.200 189.700 174.800 ;
        RECT 159.000 174.100 159.400 174.200 ;
        RECT 139.000 173.800 159.400 174.100 ;
        RECT 160.600 174.100 161.000 174.200 ;
        RECT 166.200 174.100 166.600 174.200 ;
        RECT 160.600 173.800 166.600 174.100 ;
        RECT 180.600 174.100 181.000 174.200 ;
        RECT 189.400 174.100 189.800 174.200 ;
        RECT 194.200 174.100 194.600 174.200 ;
        RECT 180.600 173.800 184.100 174.100 ;
        RECT 189.400 173.800 194.600 174.100 ;
        RECT 200.600 174.100 201.000 174.200 ;
        RECT 211.800 174.100 212.200 174.200 ;
        RECT 220.600 174.100 221.000 174.200 ;
        RECT 200.600 173.800 221.000 174.100 ;
        RECT 131.800 173.200 132.100 173.800 ;
        RECT 183.800 173.200 184.100 173.800 ;
        RECT 19.800 173.100 20.200 173.200 ;
        RECT 24.600 173.100 25.000 173.200 ;
        RECT 27.000 173.100 27.400 173.200 ;
        RECT 19.800 172.800 27.400 173.100 ;
        RECT 27.800 173.100 28.200 173.200 ;
        RECT 73.400 173.100 73.800 173.200 ;
        RECT 86.200 173.100 86.600 173.200 ;
        RECT 27.800 172.800 86.600 173.100 ;
        RECT 101.400 173.100 101.800 173.200 ;
        RECT 103.000 173.100 103.400 173.200 ;
        RECT 101.400 172.800 103.400 173.100 ;
        RECT 103.800 173.100 104.200 173.200 ;
        RECT 114.200 173.100 114.600 173.200 ;
        RECT 103.800 172.800 114.600 173.100 ;
        RECT 117.400 173.100 117.800 173.200 ;
        RECT 119.000 173.100 119.400 173.200 ;
        RECT 117.400 172.800 119.400 173.100 ;
        RECT 131.800 172.800 132.200 173.200 ;
        RECT 183.800 172.800 184.200 173.200 ;
        RECT 189.400 173.100 189.800 173.200 ;
        RECT 208.600 173.100 209.000 173.200 ;
        RECT 211.000 173.100 211.400 173.200 ;
        RECT 219.000 173.100 219.400 173.200 ;
        RECT 189.400 172.800 219.400 173.100 ;
        RECT 51.800 172.100 52.200 172.200 ;
        RECT 53.400 172.100 53.800 172.200 ;
        RECT 76.600 172.100 77.000 172.200 ;
        RECT 51.800 171.800 77.000 172.100 ;
        RECT 87.000 172.100 87.400 172.200 ;
        RECT 94.200 172.100 94.600 172.200 ;
        RECT 103.000 172.100 103.400 172.200 ;
        RECT 87.000 171.800 103.400 172.100 ;
        RECT 104.600 172.100 105.000 172.200 ;
        RECT 159.000 172.100 159.400 172.200 ;
        RECT 104.600 171.800 159.400 172.100 ;
        RECT 193.400 172.100 193.800 172.200 ;
        RECT 196.600 172.100 197.000 172.200 ;
        RECT 193.400 171.800 197.000 172.100 ;
        RECT 197.400 172.100 197.800 172.200 ;
        RECT 200.600 172.100 201.000 172.200 ;
        RECT 197.400 171.800 201.000 172.100 ;
        RECT 56.600 171.100 57.000 171.200 ;
        RECT 58.200 171.100 58.600 171.200 ;
        RECT 56.600 170.800 58.600 171.100 ;
        RECT 102.200 171.100 102.600 171.200 ;
        RECT 113.400 171.100 113.800 171.200 ;
        RECT 115.800 171.100 116.200 171.200 ;
        RECT 102.200 170.800 116.200 171.100 ;
        RECT 120.600 171.100 121.000 171.200 ;
        RECT 167.800 171.100 168.200 171.200 ;
        RECT 120.600 170.800 168.200 171.100 ;
        RECT 168.600 171.100 169.000 171.200 ;
        RECT 184.600 171.100 185.000 171.200 ;
        RECT 168.600 170.800 185.000 171.100 ;
        RECT 76.600 170.100 77.000 170.200 ;
        RECT 83.000 170.100 83.400 170.200 ;
        RECT 76.600 169.800 83.400 170.100 ;
        RECT 93.400 170.100 93.800 170.200 ;
        RECT 104.600 170.100 105.000 170.200 ;
        RECT 93.400 169.800 105.000 170.100 ;
        RECT 111.000 170.100 111.400 170.200 ;
        RECT 122.200 170.100 122.600 170.200 ;
        RECT 111.000 169.800 122.600 170.100 ;
        RECT 128.600 170.100 129.000 170.200 ;
        RECT 135.000 170.100 135.400 170.200 ;
        RECT 128.600 169.800 135.400 170.100 ;
        RECT 150.200 170.100 150.600 170.200 ;
        RECT 157.400 170.100 157.800 170.200 ;
        RECT 174.200 170.100 174.600 170.200 ;
        RECT 150.200 169.800 174.600 170.100 ;
        RECT 187.800 170.100 188.200 170.200 ;
        RECT 188.600 170.100 189.000 170.200 ;
        RECT 187.800 169.800 189.000 170.100 ;
        RECT 213.400 170.100 213.800 170.200 ;
        RECT 216.600 170.100 217.000 170.200 ;
        RECT 213.400 169.800 217.000 170.100 ;
        RECT 32.600 168.800 33.000 169.200 ;
        RECT 40.600 169.100 41.000 169.200 ;
        RECT 62.200 169.100 62.600 169.200 ;
        RECT 40.600 168.800 62.600 169.100 ;
        RECT 73.400 169.100 73.800 169.200 ;
        RECT 85.400 169.100 85.800 169.200 ;
        RECT 73.400 168.800 85.800 169.100 ;
        RECT 106.200 169.100 106.600 169.200 ;
        RECT 115.800 169.100 116.200 169.200 ;
        RECT 130.200 169.100 130.600 169.200 ;
        RECT 106.200 168.800 130.600 169.100 ;
        RECT 152.600 169.100 153.000 169.200 ;
        RECT 201.400 169.100 201.800 169.200 ;
        RECT 152.600 168.800 201.800 169.100 ;
        RECT 23.800 168.100 24.200 168.200 ;
        RECT 32.600 168.100 32.900 168.800 ;
        RECT 23.800 167.800 32.900 168.100 ;
        RECT 42.200 168.100 42.600 168.200 ;
        RECT 53.400 168.100 53.800 168.200 ;
        RECT 42.200 167.800 53.800 168.100 ;
        RECT 64.600 168.100 65.000 168.200 ;
        RECT 68.600 168.100 69.000 168.200 ;
        RECT 64.600 167.800 69.000 168.100 ;
        RECT 113.400 168.100 113.800 168.200 ;
        RECT 131.000 168.100 131.400 168.200 ;
        RECT 113.400 167.800 131.400 168.100 ;
        RECT 146.200 168.100 146.600 168.200 ;
        RECT 159.000 168.100 159.400 168.200 ;
        RECT 166.200 168.100 166.600 168.200 ;
        RECT 146.200 167.800 166.600 168.100 ;
        RECT 172.600 167.800 173.000 168.200 ;
        RECT 175.800 168.100 176.200 168.200 ;
        RECT 182.200 168.100 182.600 168.200 ;
        RECT 175.800 167.800 182.600 168.100 ;
        RECT 207.800 167.800 208.200 168.200 ;
        RECT 215.800 167.800 216.200 168.200 ;
        RECT 7.800 167.100 8.200 167.200 ;
        RECT 10.200 167.100 10.600 167.200 ;
        RECT 11.000 167.100 11.400 167.200 ;
        RECT 7.800 166.800 11.400 167.100 ;
        RECT 17.400 167.100 17.800 167.200 ;
        RECT 19.000 167.100 19.400 167.200 ;
        RECT 17.400 166.800 19.400 167.100 ;
        RECT 27.800 167.100 28.200 167.200 ;
        RECT 43.000 167.100 43.400 167.200 ;
        RECT 27.800 166.800 43.400 167.100 ;
        RECT 51.800 167.100 52.200 167.200 ;
        RECT 52.600 167.100 53.000 167.200 ;
        RECT 51.800 166.800 53.000 167.100 ;
        RECT 58.200 167.100 58.600 167.200 ;
        RECT 59.000 167.100 59.400 167.200 ;
        RECT 58.200 166.800 59.400 167.100 ;
        RECT 66.200 166.800 66.600 167.200 ;
        RECT 75.000 166.800 75.400 167.200 ;
        RECT 95.000 167.100 95.400 167.200 ;
        RECT 100.600 167.100 101.000 167.200 ;
        RECT 103.800 167.100 104.200 167.200 ;
        RECT 95.000 166.800 104.200 167.100 ;
        RECT 123.800 167.100 124.200 167.200 ;
        RECT 127.800 167.100 128.200 167.200 ;
        RECT 123.800 166.800 128.200 167.100 ;
        RECT 129.400 166.800 129.800 167.200 ;
        RECT 135.800 167.100 136.200 167.200 ;
        RECT 138.200 167.100 138.600 167.200 ;
        RECT 135.800 166.800 138.600 167.100 ;
        RECT 144.600 167.100 145.000 167.200 ;
        RECT 154.200 167.100 154.600 167.200 ;
        RECT 144.600 166.800 154.600 167.100 ;
        RECT 155.800 167.100 156.200 167.200 ;
        RECT 156.600 167.100 157.000 167.200 ;
        RECT 155.800 166.800 157.000 167.100 ;
        RECT 161.400 167.100 161.800 167.200 ;
        RECT 170.200 167.100 170.600 167.200 ;
        RECT 161.400 166.800 170.600 167.100 ;
        RECT 172.600 167.100 172.900 167.800 ;
        RECT 179.800 167.100 180.200 167.200 ;
        RECT 181.400 167.100 181.800 167.200 ;
        RECT 172.600 166.800 181.800 167.100 ;
        RECT 187.800 166.800 188.200 167.200 ;
        RECT 197.400 167.100 197.800 167.200 ;
        RECT 203.000 167.100 203.400 167.200 ;
        RECT 197.400 166.800 203.400 167.100 ;
        RECT 207.800 167.100 208.100 167.800 ;
        RECT 215.800 167.100 216.100 167.800 ;
        RECT 207.800 166.800 216.100 167.100 ;
        RECT 18.200 166.100 18.600 166.200 ;
        RECT 27.800 166.100 28.200 166.200 ;
        RECT 18.200 165.800 28.200 166.100 ;
        RECT 35.000 166.100 35.400 166.200 ;
        RECT 35.800 166.100 36.200 166.200 ;
        RECT 35.000 165.800 36.200 166.100 ;
        RECT 43.000 166.100 43.300 166.800 ;
        RECT 46.200 166.100 46.600 166.200 ;
        RECT 43.000 165.800 46.600 166.100 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 66.200 166.100 66.500 166.800 ;
        RECT 67.000 166.100 67.400 166.200 ;
        RECT 51.800 165.800 67.400 166.100 ;
        RECT 68.600 166.100 69.000 166.200 ;
        RECT 73.400 166.100 73.800 166.200 ;
        RECT 68.600 165.800 73.800 166.100 ;
        RECT 75.000 166.100 75.300 166.800 ;
        RECT 80.600 166.100 81.000 166.200 ;
        RECT 75.000 165.800 81.000 166.100 ;
        RECT 91.000 166.100 91.400 166.200 ;
        RECT 92.600 166.100 93.000 166.200 ;
        RECT 91.000 165.800 93.000 166.100 ;
        RECT 97.400 165.800 97.800 166.200 ;
        RECT 98.200 166.100 98.600 166.200 ;
        RECT 99.800 166.100 100.200 166.200 ;
        RECT 104.600 166.100 105.000 166.200 ;
        RECT 98.200 165.800 105.000 166.100 ;
        RECT 105.400 166.100 105.800 166.200 ;
        RECT 114.200 166.100 114.600 166.200 ;
        RECT 115.000 166.100 115.400 166.200 ;
        RECT 105.400 165.800 115.400 166.100 ;
        RECT 121.400 166.100 121.800 166.200 ;
        RECT 129.400 166.100 129.700 166.800 ;
        RECT 139.800 166.100 140.200 166.200 ;
        RECT 121.400 165.800 140.200 166.100 ;
        RECT 152.600 166.100 153.000 166.200 ;
        RECT 155.000 166.100 155.400 166.200 ;
        RECT 152.600 165.800 155.400 166.100 ;
        RECT 157.400 166.100 157.800 166.200 ;
        RECT 167.000 166.100 167.400 166.200 ;
        RECT 184.600 166.100 185.000 166.200 ;
        RECT 187.800 166.100 188.100 166.800 ;
        RECT 157.400 165.800 167.400 166.100 ;
        RECT 175.000 165.800 177.700 166.100 ;
        RECT 184.600 165.800 188.100 166.100 ;
        RECT 199.000 165.800 199.400 166.200 ;
        RECT 217.400 166.100 217.800 166.200 ;
        RECT 219.800 166.100 220.200 166.200 ;
        RECT 217.400 165.800 220.200 166.100 ;
        RECT 11.000 165.100 11.400 165.200 ;
        RECT 12.600 165.100 13.000 165.200 ;
        RECT 15.800 165.100 16.200 165.200 ;
        RECT 11.000 164.800 16.200 165.100 ;
        RECT 32.600 165.100 33.000 165.200 ;
        RECT 36.600 165.100 37.000 165.200 ;
        RECT 32.600 164.800 37.000 165.100 ;
        RECT 47.800 165.100 48.200 165.200 ;
        RECT 54.200 165.100 54.600 165.200 ;
        RECT 47.800 164.800 54.600 165.100 ;
        RECT 56.600 165.100 57.000 165.200 ;
        RECT 60.600 165.100 61.000 165.200 ;
        RECT 70.200 165.100 70.600 165.200 ;
        RECT 71.800 165.100 72.200 165.200 ;
        RECT 56.600 164.800 72.200 165.100 ;
        RECT 97.400 165.100 97.700 165.800 ;
        RECT 124.600 165.200 124.900 165.800 ;
        RECT 175.000 165.200 175.300 165.800 ;
        RECT 177.400 165.200 177.700 165.800 ;
        RECT 100.600 165.100 101.000 165.200 ;
        RECT 116.600 165.100 117.000 165.200 ;
        RECT 97.400 164.800 101.000 165.100 ;
        RECT 102.200 164.800 117.000 165.100 ;
        RECT 121.400 165.100 121.800 165.200 ;
        RECT 123.800 165.100 124.200 165.200 ;
        RECT 121.400 164.800 124.200 165.100 ;
        RECT 124.600 164.800 125.000 165.200 ;
        RECT 125.400 165.100 125.800 165.200 ;
        RECT 126.200 165.100 126.600 165.200 ;
        RECT 135.800 165.100 136.200 165.200 ;
        RECT 125.400 164.800 126.600 165.100 ;
        RECT 131.800 164.800 136.200 165.100 ;
        RECT 136.600 165.100 137.000 165.200 ;
        RECT 137.400 165.100 137.800 165.200 ;
        RECT 136.600 164.800 137.800 165.100 ;
        RECT 155.000 165.100 155.400 165.200 ;
        RECT 157.400 165.100 157.800 165.200 ;
        RECT 155.000 164.800 157.800 165.100 ;
        RECT 168.600 165.100 169.000 165.200 ;
        RECT 169.400 165.100 169.800 165.200 ;
        RECT 171.800 165.100 172.200 165.200 ;
        RECT 168.600 164.800 172.200 165.100 ;
        RECT 175.000 164.800 175.400 165.200 ;
        RECT 177.400 164.800 177.800 165.200 ;
        RECT 178.200 165.100 178.600 165.200 ;
        RECT 179.000 165.100 179.400 165.200 ;
        RECT 178.200 164.800 179.400 165.100 ;
        RECT 183.800 165.100 184.200 165.200 ;
        RECT 186.200 165.100 186.600 165.200 ;
        RECT 183.800 164.800 186.600 165.100 ;
        RECT 187.000 165.100 187.400 165.200 ;
        RECT 199.000 165.100 199.300 165.800 ;
        RECT 187.000 164.800 199.300 165.100 ;
        RECT 199.800 165.100 200.200 165.200 ;
        RECT 201.400 165.100 201.800 165.200 ;
        RECT 199.800 164.800 201.800 165.100 ;
        RECT 212.600 165.100 213.000 165.200 ;
        RECT 218.200 165.100 218.600 165.200 ;
        RECT 212.600 164.800 218.600 165.100 ;
        RECT 223.800 165.100 224.200 165.200 ;
        RECT 227.800 165.100 228.200 165.200 ;
        RECT 223.800 164.800 228.200 165.100 ;
        RECT 102.200 164.200 102.500 164.800 ;
        RECT 131.800 164.200 132.100 164.800 ;
        RECT 53.400 164.100 53.800 164.200 ;
        RECT 59.000 164.100 59.400 164.200 ;
        RECT 75.800 164.100 76.200 164.200 ;
        RECT 53.400 163.800 76.200 164.100 ;
        RECT 83.000 164.100 83.400 164.200 ;
        RECT 91.800 164.100 92.200 164.200 ;
        RECT 98.200 164.100 98.600 164.200 ;
        RECT 83.000 163.800 98.600 164.100 ;
        RECT 99.000 164.100 99.400 164.200 ;
        RECT 102.200 164.100 102.600 164.200 ;
        RECT 99.000 163.800 102.600 164.100 ;
        RECT 131.800 163.800 132.200 164.200 ;
        RECT 155.800 164.100 156.200 164.200 ;
        RECT 173.400 164.100 173.800 164.200 ;
        RECT 155.800 163.800 173.800 164.100 ;
        RECT 177.400 164.100 177.800 164.200 ;
        RECT 180.600 164.100 181.000 164.200 ;
        RECT 177.400 163.800 181.000 164.100 ;
        RECT 183.800 164.100 184.200 164.200 ;
        RECT 195.000 164.100 195.400 164.200 ;
        RECT 183.800 163.800 195.400 164.100 ;
        RECT 199.000 164.100 199.400 164.200 ;
        RECT 200.600 164.100 201.000 164.200 ;
        RECT 199.000 163.800 201.000 164.100 ;
        RECT 63.800 163.100 64.200 163.200 ;
        RECT 106.200 163.100 106.600 163.200 ;
        RECT 63.800 162.800 106.600 163.100 ;
        RECT 129.400 163.100 129.800 163.200 ;
        RECT 174.200 163.100 174.600 163.200 ;
        RECT 129.400 162.800 174.600 163.100 ;
        RECT 5.400 162.100 5.800 162.200 ;
        RECT 8.600 162.100 9.000 162.200 ;
        RECT 5.400 161.800 9.000 162.100 ;
        RECT 23.000 162.100 23.400 162.200 ;
        RECT 75.000 162.100 75.400 162.200 ;
        RECT 23.000 161.800 75.400 162.100 ;
        RECT 97.400 162.100 97.800 162.200 ;
        RECT 99.000 162.100 99.400 162.200 ;
        RECT 97.400 161.800 99.400 162.100 ;
        RECT 99.800 162.100 100.200 162.200 ;
        RECT 102.200 162.100 102.600 162.200 ;
        RECT 109.400 162.100 109.800 162.200 ;
        RECT 99.800 161.800 109.800 162.100 ;
        RECT 123.800 162.100 124.200 162.200 ;
        RECT 132.600 162.100 133.000 162.200 ;
        RECT 123.800 161.800 133.000 162.100 ;
        RECT 136.600 162.100 137.000 162.200 ;
        RECT 143.800 162.100 144.200 162.200 ;
        RECT 136.600 161.800 144.200 162.100 ;
        RECT 153.400 162.100 153.800 162.200 ;
        RECT 154.200 162.100 154.600 162.200 ;
        RECT 186.200 162.100 186.600 162.200 ;
        RECT 202.200 162.100 202.600 162.200 ;
        RECT 153.400 161.800 202.600 162.100 ;
        RECT 42.200 161.100 42.600 161.200 ;
        RECT 95.000 161.100 95.400 161.200 ;
        RECT 127.000 161.100 127.400 161.200 ;
        RECT 42.200 160.800 127.400 161.100 ;
        RECT 73.400 160.100 73.800 160.200 ;
        RECT 101.400 160.100 101.800 160.200 ;
        RECT 73.400 159.800 101.800 160.100 ;
        RECT 103.000 160.100 103.400 160.200 ;
        RECT 123.800 160.100 124.200 160.200 ;
        RECT 103.000 159.800 124.200 160.100 ;
        RECT 167.800 160.100 168.200 160.200 ;
        RECT 174.200 160.100 174.600 160.200 ;
        RECT 167.800 159.800 174.600 160.100 ;
        RECT 53.400 159.100 53.800 159.200 ;
        RECT 61.400 159.100 61.800 159.200 ;
        RECT 53.400 158.800 61.800 159.100 ;
        RECT 63.800 159.100 64.200 159.200 ;
        RECT 100.600 159.100 101.000 159.200 ;
        RECT 63.800 158.800 101.000 159.100 ;
        RECT 114.200 159.100 114.600 159.200 ;
        RECT 183.000 159.100 183.400 159.200 ;
        RECT 114.200 158.800 183.400 159.100 ;
        RECT 18.200 158.100 18.600 158.200 ;
        RECT 25.400 158.100 25.800 158.200 ;
        RECT 32.600 158.100 33.000 158.200 ;
        RECT 18.200 157.800 33.000 158.100 ;
        RECT 61.400 158.100 61.800 158.200 ;
        RECT 78.200 158.100 78.600 158.200 ;
        RECT 61.400 157.800 78.600 158.100 ;
        RECT 98.200 158.100 98.600 158.200 ;
        RECT 99.000 158.100 99.400 158.200 ;
        RECT 123.800 158.100 124.200 158.200 ;
        RECT 98.200 157.800 124.200 158.100 ;
        RECT 138.200 158.100 138.600 158.200 ;
        RECT 142.200 158.100 142.600 158.200 ;
        RECT 138.200 157.800 142.600 158.100 ;
        RECT 180.600 158.100 181.000 158.200 ;
        RECT 183.800 158.100 184.200 158.200 ;
        RECT 180.600 157.800 184.200 158.100 ;
        RECT 207.000 158.100 207.400 158.200 ;
        RECT 216.600 158.100 217.000 158.200 ;
        RECT 207.000 157.800 217.000 158.100 ;
        RECT 1.400 157.100 1.800 157.200 ;
        RECT 6.200 157.100 6.600 157.200 ;
        RECT 17.400 157.100 17.800 157.200 ;
        RECT 1.400 156.800 17.800 157.100 ;
        RECT 25.400 157.100 25.800 157.200 ;
        RECT 44.600 157.100 45.000 157.200 ;
        RECT 25.400 156.800 45.000 157.100 ;
        RECT 46.200 157.100 46.600 157.200 ;
        RECT 55.000 157.100 55.400 157.200 ;
        RECT 46.200 156.800 55.400 157.100 ;
        RECT 63.800 157.100 64.200 157.200 ;
        RECT 68.600 157.100 69.000 157.200 ;
        RECT 63.800 156.800 69.000 157.100 ;
        RECT 71.800 157.100 72.200 157.200 ;
        RECT 103.800 157.100 104.200 157.200 ;
        RECT 71.800 156.800 104.200 157.100 ;
        RECT 143.800 157.100 144.200 157.200 ;
        RECT 151.000 157.100 151.400 157.200 ;
        RECT 143.800 156.800 151.400 157.100 ;
        RECT 159.000 157.100 159.400 157.200 ;
        RECT 170.200 157.100 170.600 157.200 ;
        RECT 159.000 156.800 170.600 157.100 ;
        RECT 171.800 156.800 172.200 157.200 ;
        RECT 178.200 157.100 178.600 157.200 ;
        RECT 184.600 157.100 185.000 157.200 ;
        RECT 178.200 156.800 185.000 157.100 ;
        RECT 202.200 157.100 202.600 157.200 ;
        RECT 212.600 157.100 213.000 157.200 ;
        RECT 216.600 157.100 217.000 157.200 ;
        RECT 202.200 156.800 217.000 157.100 ;
        RECT 226.200 156.800 226.600 157.200 ;
        RECT 17.400 156.100 17.800 156.200 ;
        RECT 11.800 155.800 17.800 156.100 ;
        RECT 30.200 156.100 30.600 156.200 ;
        RECT 55.800 156.100 56.200 156.200 ;
        RECT 30.200 155.800 56.200 156.100 ;
        RECT 58.200 156.100 58.600 156.200 ;
        RECT 65.400 156.100 65.800 156.200 ;
        RECT 58.200 155.800 65.800 156.100 ;
        RECT 67.000 156.100 67.400 156.200 ;
        RECT 67.800 156.100 68.200 156.200 ;
        RECT 67.000 155.800 68.200 156.100 ;
        RECT 79.000 156.100 79.400 156.200 ;
        RECT 85.400 156.100 85.800 156.200 ;
        RECT 89.400 156.100 89.800 156.200 ;
        RECT 79.000 155.800 85.800 156.100 ;
        RECT 86.200 155.800 89.800 156.100 ;
        RECT 95.800 156.100 96.200 156.200 ;
        RECT 108.600 156.100 109.000 156.200 ;
        RECT 95.800 155.800 109.000 156.100 ;
        RECT 109.400 156.100 109.800 156.200 ;
        RECT 120.600 156.100 121.000 156.200 ;
        RECT 109.400 155.800 121.000 156.100 ;
        RECT 121.400 156.100 121.800 156.200 ;
        RECT 131.800 156.100 132.200 156.200 ;
        RECT 121.400 155.800 132.200 156.100 ;
        RECT 135.800 156.100 136.200 156.200 ;
        RECT 142.200 156.100 142.600 156.200 ;
        RECT 135.800 155.800 142.600 156.100 ;
        RECT 145.400 156.100 145.800 156.200 ;
        RECT 154.200 156.100 154.600 156.200 ;
        RECT 145.400 155.800 154.600 156.100 ;
        RECT 156.600 155.800 157.000 156.200 ;
        RECT 157.400 156.100 157.800 156.200 ;
        RECT 160.600 156.100 161.000 156.200 ;
        RECT 157.400 155.800 161.000 156.100 ;
        RECT 167.000 156.100 167.400 156.200 ;
        RECT 171.800 156.100 172.100 156.800 ;
        RECT 167.000 155.800 172.100 156.100 ;
        RECT 179.800 156.100 180.200 156.200 ;
        RECT 180.600 156.100 181.000 156.200 ;
        RECT 179.800 155.800 181.000 156.100 ;
        RECT 196.600 155.800 197.000 156.200 ;
        RECT 210.200 156.100 210.600 156.200 ;
        RECT 221.400 156.100 221.800 156.200 ;
        RECT 210.200 155.800 221.800 156.100 ;
        RECT 222.200 156.100 222.600 156.200 ;
        RECT 226.200 156.100 226.500 156.800 ;
        RECT 222.200 155.800 226.500 156.100 ;
        RECT 11.800 155.200 12.100 155.800 ;
        RECT 86.200 155.200 86.500 155.800 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 10.200 155.100 10.600 155.200 ;
        RECT 3.800 154.800 10.600 155.100 ;
        RECT 11.800 154.800 12.200 155.200 ;
        RECT 41.400 155.100 41.800 155.200 ;
        RECT 51.800 155.100 52.200 155.200 ;
        RECT 41.400 154.800 52.200 155.100 ;
        RECT 65.400 155.100 65.800 155.200 ;
        RECT 67.000 155.100 67.400 155.200 ;
        RECT 65.400 154.800 67.400 155.100 ;
        RECT 83.800 155.100 84.200 155.200 ;
        RECT 84.600 155.100 85.000 155.200 ;
        RECT 83.800 154.800 85.000 155.100 ;
        RECT 86.200 154.800 86.600 155.200 ;
        RECT 93.400 155.100 93.800 155.200 ;
        RECT 100.600 155.100 101.000 155.200 ;
        RECT 93.400 154.800 101.000 155.100 ;
        RECT 116.600 154.800 117.000 155.200 ;
        RECT 123.000 155.100 123.400 155.200 ;
        RECT 125.400 155.100 125.800 155.200 ;
        RECT 123.000 154.800 125.800 155.100 ;
        RECT 127.800 155.100 128.200 155.200 ;
        RECT 128.600 155.100 129.000 155.200 ;
        RECT 127.800 154.800 129.000 155.100 ;
        RECT 130.200 155.100 130.600 155.200 ;
        RECT 145.400 155.100 145.800 155.200 ;
        RECT 130.200 154.800 145.800 155.100 ;
        RECT 147.000 155.100 147.400 155.200 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 147.000 154.800 148.200 155.100 ;
        RECT 148.600 155.100 149.000 155.200 ;
        RECT 156.600 155.100 156.900 155.800 ;
        RECT 196.600 155.200 196.900 155.800 ;
        RECT 148.600 154.800 156.900 155.100 ;
        RECT 159.800 155.100 160.200 155.200 ;
        RECT 171.000 155.100 171.400 155.200 ;
        RECT 159.800 154.800 171.400 155.100 ;
        RECT 181.400 155.100 181.800 155.200 ;
        RECT 183.800 155.100 184.200 155.200 ;
        RECT 181.400 154.800 184.200 155.100 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 199.000 154.800 199.400 155.200 ;
        RECT 209.400 155.100 209.800 155.200 ;
        RECT 211.000 155.100 211.400 155.200 ;
        RECT 213.400 155.100 213.800 155.200 ;
        RECT 209.400 154.800 213.800 155.100 ;
        RECT 214.200 154.800 214.600 155.200 ;
        RECT 215.800 154.800 216.200 155.200 ;
        RECT 220.600 155.100 221.000 155.200 ;
        RECT 221.400 155.100 221.800 155.200 ;
        RECT 220.600 154.800 221.800 155.100 ;
        RECT 224.600 154.800 225.000 155.200 ;
        RECT 10.200 154.200 10.500 154.800 ;
        RECT 3.800 154.100 4.200 154.200 ;
        RECT 7.800 154.100 8.200 154.200 ;
        RECT 3.800 153.800 8.200 154.100 ;
        RECT 10.200 153.800 10.600 154.200 ;
        RECT 15.000 154.100 15.400 154.200 ;
        RECT 11.800 153.800 15.400 154.100 ;
        RECT 43.800 153.800 44.200 154.200 ;
        RECT 47.800 154.100 48.200 154.200 ;
        RECT 56.600 154.100 57.000 154.200 ;
        RECT 71.000 154.100 71.400 154.200 ;
        RECT 47.800 153.800 71.400 154.100 ;
        RECT 76.600 154.100 77.000 154.200 ;
        RECT 84.600 154.100 85.000 154.200 ;
        RECT 98.200 154.100 98.600 154.200 ;
        RECT 76.600 153.800 98.600 154.100 ;
        RECT 102.200 154.100 102.600 154.200 ;
        RECT 111.000 154.100 111.400 154.200 ;
        RECT 102.200 153.800 111.400 154.100 ;
        RECT 111.800 154.100 112.200 154.200 ;
        RECT 116.600 154.100 116.900 154.800 ;
        RECT 199.000 154.200 199.300 154.800 ;
        RECT 214.200 154.200 214.500 154.800 ;
        RECT 111.800 153.800 116.900 154.100 ;
        RECT 119.000 154.100 119.400 154.200 ;
        RECT 133.400 154.100 133.800 154.200 ;
        RECT 119.000 153.800 133.800 154.100 ;
        RECT 134.200 154.100 134.600 154.200 ;
        RECT 155.000 154.100 155.400 154.200 ;
        RECT 134.200 153.800 155.400 154.100 ;
        RECT 172.600 154.100 173.000 154.200 ;
        RECT 179.000 154.100 179.400 154.200 ;
        RECT 172.600 153.800 179.400 154.100 ;
        RECT 180.600 154.100 181.000 154.200 ;
        RECT 181.400 154.100 181.800 154.200 ;
        RECT 180.600 153.800 181.800 154.100 ;
        RECT 183.800 154.100 184.200 154.200 ;
        RECT 190.200 154.100 190.600 154.200 ;
        RECT 183.800 153.800 190.600 154.100 ;
        RECT 199.000 153.800 199.400 154.200 ;
        RECT 205.400 154.100 205.800 154.200 ;
        RECT 207.000 154.100 207.400 154.200 ;
        RECT 207.800 154.100 208.200 154.200 ;
        RECT 205.400 153.800 208.200 154.100 ;
        RECT 214.200 153.800 214.600 154.200 ;
        RECT 215.800 154.100 216.100 154.800 ;
        RECT 217.400 154.100 217.800 154.200 ;
        RECT 220.600 154.100 221.000 154.200 ;
        RECT 215.800 153.800 221.000 154.100 ;
        RECT 224.600 154.100 224.900 154.800 ;
        RECT 229.400 154.100 229.800 154.200 ;
        RECT 224.600 153.800 229.800 154.100 ;
        RECT 11.800 153.200 12.100 153.800 ;
        RECT 43.800 153.200 44.100 153.800 ;
        RECT 155.000 153.200 155.300 153.800 ;
        RECT 0.600 153.100 1.000 153.200 ;
        RECT 4.600 153.100 5.000 153.200 ;
        RECT 0.600 152.800 5.000 153.100 ;
        RECT 11.800 152.800 12.200 153.200 ;
        RECT 35.800 153.100 36.200 153.200 ;
        RECT 42.200 153.100 42.600 153.200 ;
        RECT 35.800 152.800 42.600 153.100 ;
        RECT 43.800 152.800 44.200 153.200 ;
        RECT 46.200 153.100 46.600 153.200 ;
        RECT 75.000 153.100 75.400 153.200 ;
        RECT 46.200 152.800 75.400 153.100 ;
        RECT 79.800 153.100 80.200 153.200 ;
        RECT 89.400 153.100 89.800 153.200 ;
        RECT 79.800 152.800 89.800 153.100 ;
        RECT 94.200 153.100 94.600 153.200 ;
        RECT 99.800 153.100 100.200 153.200 ;
        RECT 94.200 152.800 100.200 153.100 ;
        RECT 100.600 153.100 101.000 153.200 ;
        RECT 104.600 153.100 105.000 153.200 ;
        RECT 100.600 152.800 105.000 153.100 ;
        RECT 105.400 153.100 105.800 153.200 ;
        RECT 130.200 153.100 130.600 153.200 ;
        RECT 105.400 152.800 130.600 153.100 ;
        RECT 139.000 153.100 139.400 153.200 ;
        RECT 139.800 153.100 140.200 153.200 ;
        RECT 146.200 153.100 146.600 153.200 ;
        RECT 139.000 152.800 140.200 153.100 ;
        RECT 143.000 152.800 146.600 153.100 ;
        RECT 148.600 153.100 149.000 153.200 ;
        RECT 153.400 153.100 153.800 153.200 ;
        RECT 148.600 152.800 153.800 153.100 ;
        RECT 155.000 152.800 155.400 153.200 ;
        RECT 175.000 153.100 175.400 153.200 ;
        RECT 175.800 153.100 176.200 153.200 ;
        RECT 175.000 152.800 176.200 153.100 ;
        RECT 176.600 153.100 177.000 153.200 ;
        RECT 180.600 153.100 181.000 153.200 ;
        RECT 176.600 152.800 181.000 153.100 ;
        RECT 195.800 153.100 196.200 153.200 ;
        RECT 200.600 153.100 201.000 153.200 ;
        RECT 195.800 152.800 201.000 153.100 ;
        RECT 203.000 153.100 203.400 153.200 ;
        RECT 226.200 153.100 226.600 153.200 ;
        RECT 203.000 152.800 226.600 153.100 ;
        RECT 143.000 152.200 143.300 152.800 ;
        RECT 9.400 152.100 9.800 152.200 ;
        RECT 11.800 152.100 12.200 152.200 ;
        RECT 9.400 151.800 12.200 152.100 ;
        RECT 19.800 152.100 20.200 152.200 ;
        RECT 20.600 152.100 21.000 152.200 ;
        RECT 19.800 151.800 21.000 152.100 ;
        RECT 31.800 152.100 32.200 152.200 ;
        RECT 46.200 152.100 46.600 152.200 ;
        RECT 31.800 151.800 46.600 152.100 ;
        RECT 51.800 152.100 52.200 152.200 ;
        RECT 57.400 152.100 57.800 152.200 ;
        RECT 84.600 152.100 85.000 152.200 ;
        RECT 87.000 152.100 87.400 152.200 ;
        RECT 51.800 151.800 87.400 152.100 ;
        RECT 91.000 152.100 91.400 152.200 ;
        RECT 114.200 152.100 114.600 152.200 ;
        RECT 91.000 151.800 114.600 152.100 ;
        RECT 115.800 152.100 116.200 152.200 ;
        RECT 123.000 152.100 123.400 152.200 ;
        RECT 115.800 151.800 123.400 152.100 ;
        RECT 125.400 152.100 125.800 152.200 ;
        RECT 139.000 152.100 139.400 152.200 ;
        RECT 125.400 151.800 139.400 152.100 ;
        RECT 143.000 151.800 143.400 152.200 ;
        RECT 144.600 152.100 145.000 152.200 ;
        RECT 151.800 152.100 152.200 152.200 ;
        RECT 144.600 151.800 152.200 152.100 ;
        RECT 163.800 152.100 164.200 152.200 ;
        RECT 175.800 152.100 176.200 152.200 ;
        RECT 163.800 151.800 176.200 152.100 ;
        RECT 179.800 152.100 180.200 152.200 ;
        RECT 215.000 152.100 215.400 152.200 ;
        RECT 179.800 151.800 215.400 152.100 ;
        RECT 219.800 152.100 220.200 152.200 ;
        RECT 225.400 152.100 225.800 152.200 ;
        RECT 219.800 151.800 225.800 152.100 ;
        RECT 40.600 151.100 41.000 151.200 ;
        RECT 45.400 151.100 45.800 151.200 ;
        RECT 40.600 150.800 45.800 151.100 ;
        RECT 73.400 151.100 73.800 151.200 ;
        RECT 74.200 151.100 74.600 151.200 ;
        RECT 73.400 150.800 74.600 151.100 ;
        RECT 91.000 151.100 91.400 151.200 ;
        RECT 106.200 151.100 106.600 151.200 ;
        RECT 123.000 151.100 123.400 151.200 ;
        RECT 91.000 150.800 123.400 151.100 ;
        RECT 139.800 151.100 140.200 151.200 ;
        RECT 145.400 151.100 145.800 151.200 ;
        RECT 155.000 151.100 155.400 151.200 ;
        RECT 139.800 150.800 155.400 151.100 ;
        RECT 157.400 151.100 157.800 151.200 ;
        RECT 173.400 151.100 173.800 151.200 ;
        RECT 157.400 150.800 173.800 151.100 ;
        RECT 198.200 150.800 198.600 151.200 ;
        RECT 198.200 150.200 198.500 150.800 ;
        RECT 5.400 150.100 5.800 150.200 ;
        RECT 23.800 150.100 24.200 150.200 ;
        RECT 5.400 149.800 24.200 150.100 ;
        RECT 36.600 150.100 37.000 150.200 ;
        RECT 54.200 150.100 54.600 150.200 ;
        RECT 36.600 149.800 54.600 150.100 ;
        RECT 70.200 150.100 70.600 150.200 ;
        RECT 87.000 150.100 87.400 150.200 ;
        RECT 70.200 149.800 87.400 150.100 ;
        RECT 95.800 150.100 96.200 150.200 ;
        RECT 96.600 150.100 97.000 150.200 ;
        RECT 149.400 150.100 149.800 150.200 ;
        RECT 95.800 149.800 149.800 150.100 ;
        RECT 164.600 150.100 165.000 150.200 ;
        RECT 179.000 150.100 179.400 150.200 ;
        RECT 164.600 149.800 179.400 150.100 ;
        RECT 198.200 149.800 198.600 150.200 ;
        RECT 205.400 149.800 205.800 150.200 ;
        RECT 216.600 150.100 217.000 150.200 ;
        RECT 227.000 150.100 227.400 150.200 ;
        RECT 216.600 149.800 227.400 150.100 ;
        RECT 10.200 149.100 10.600 149.200 ;
        RECT 15.000 149.100 15.400 149.200 ;
        RECT 39.000 149.100 39.400 149.200 ;
        RECT 10.200 148.800 15.400 149.100 ;
        RECT 23.000 148.800 39.400 149.100 ;
        RECT 44.600 149.100 45.000 149.200 ;
        RECT 64.600 149.100 65.000 149.200 ;
        RECT 104.600 149.100 105.000 149.200 ;
        RECT 113.400 149.100 113.800 149.200 ;
        RECT 44.600 148.800 81.700 149.100 ;
        RECT 104.600 148.800 113.800 149.100 ;
        RECT 114.200 149.100 114.600 149.200 ;
        RECT 115.800 149.100 116.200 149.200 ;
        RECT 147.000 149.100 147.400 149.200 ;
        RECT 114.200 148.800 147.400 149.100 ;
        RECT 147.800 149.100 148.200 149.200 ;
        RECT 153.400 149.100 153.800 149.200 ;
        RECT 147.800 148.800 153.800 149.100 ;
        RECT 154.200 149.100 154.600 149.200 ;
        RECT 163.800 149.100 164.200 149.200 ;
        RECT 154.200 148.800 164.200 149.100 ;
        RECT 172.600 149.100 173.000 149.200 ;
        RECT 187.800 149.100 188.200 149.200 ;
        RECT 189.400 149.100 189.800 149.200 ;
        RECT 172.600 148.800 189.800 149.100 ;
        RECT 194.200 149.100 194.600 149.200 ;
        RECT 195.000 149.100 195.400 149.200 ;
        RECT 199.000 149.100 199.400 149.200 ;
        RECT 194.200 148.800 199.400 149.100 ;
        RECT 200.600 149.100 201.000 149.200 ;
        RECT 205.400 149.100 205.700 149.800 ;
        RECT 200.600 148.800 205.700 149.100 ;
        RECT 207.000 148.800 207.400 149.200 ;
        RECT 23.000 148.200 23.300 148.800 ;
        RECT 8.600 148.100 9.000 148.200 ;
        RECT 10.200 148.100 10.600 148.200 ;
        RECT 8.600 147.800 10.600 148.100 ;
        RECT 20.600 147.800 21.000 148.200 ;
        RECT 23.000 147.800 23.400 148.200 ;
        RECT 36.600 148.100 37.000 148.200 ;
        RECT 47.800 148.100 48.200 148.200 ;
        RECT 70.200 148.100 70.600 148.200 ;
        RECT 36.600 147.800 70.600 148.100 ;
        RECT 77.400 148.100 77.800 148.200 ;
        RECT 80.600 148.100 81.000 148.200 ;
        RECT 77.400 147.800 81.000 148.100 ;
        RECT 81.400 148.100 81.700 148.800 ;
        RECT 207.000 148.200 207.300 148.800 ;
        RECT 118.200 148.100 118.600 148.200 ;
        RECT 81.400 147.800 118.600 148.100 ;
        RECT 127.800 148.100 128.200 148.200 ;
        RECT 128.600 148.100 129.000 148.200 ;
        RECT 127.800 147.800 129.000 148.100 ;
        RECT 130.200 148.100 130.600 148.200 ;
        RECT 131.800 148.100 132.200 148.200 ;
        RECT 130.200 147.800 132.200 148.100 ;
        RECT 133.400 148.100 133.800 148.200 ;
        RECT 136.600 148.100 137.000 148.200 ;
        RECT 133.400 147.800 137.000 148.100 ;
        RECT 147.800 147.800 148.200 148.200 ;
        RECT 149.400 148.100 149.800 148.200 ;
        RECT 178.200 148.100 178.600 148.200 ;
        RECT 149.400 147.800 178.600 148.100 ;
        RECT 189.400 148.100 189.800 148.200 ;
        RECT 204.600 148.100 205.000 148.200 ;
        RECT 189.400 147.800 205.000 148.100 ;
        RECT 207.000 147.800 207.400 148.200 ;
        RECT 3.800 146.800 4.200 147.200 ;
        RECT 11.000 147.100 11.400 147.200 ;
        RECT 20.600 147.100 20.900 147.800 ;
        RECT 11.000 146.800 20.900 147.100 ;
        RECT 30.200 147.100 30.600 147.200 ;
        RECT 31.000 147.100 31.400 147.200 ;
        RECT 30.200 146.800 31.400 147.100 ;
        RECT 34.200 147.100 34.600 147.200 ;
        RECT 35.800 147.100 36.200 147.200 ;
        RECT 34.200 146.800 36.200 147.100 ;
        RECT 45.400 147.100 45.800 147.200 ;
        RECT 47.800 147.100 48.200 147.200 ;
        RECT 45.400 146.800 48.200 147.100 ;
        RECT 53.400 147.100 53.800 147.200 ;
        RECT 69.400 147.100 69.800 147.200 ;
        RECT 53.400 146.800 69.800 147.100 ;
        RECT 70.200 147.100 70.600 147.200 ;
        RECT 78.200 147.100 78.600 147.200 ;
        RECT 70.200 146.800 78.600 147.100 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 96.600 147.100 97.000 147.200 ;
        RECT 103.000 147.100 103.400 147.200 ;
        RECT 79.800 146.800 103.400 147.100 ;
        RECT 105.400 147.100 105.800 147.200 ;
        RECT 117.400 147.100 117.800 147.200 ;
        RECT 105.400 146.800 117.800 147.100 ;
        RECT 119.000 147.100 119.400 147.200 ;
        RECT 126.200 147.100 126.600 147.200 ;
        RECT 135.000 147.100 135.400 147.200 ;
        RECT 139.800 147.100 140.200 147.200 ;
        RECT 119.000 146.800 140.200 147.100 ;
        RECT 146.200 146.800 146.600 147.200 ;
        RECT 147.800 147.100 148.100 147.800 ;
        RECT 152.600 147.100 153.000 147.200 ;
        RECT 159.000 147.100 159.400 147.200 ;
        RECT 147.800 146.800 151.300 147.100 ;
        RECT 152.600 146.800 159.400 147.100 ;
        RECT 163.800 147.100 164.200 147.200 ;
        RECT 196.600 147.100 197.000 147.200 ;
        RECT 163.800 146.800 197.000 147.100 ;
        RECT 199.000 146.800 199.400 147.200 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 223.000 146.800 223.400 147.200 ;
        RECT 3.800 146.100 4.100 146.800 ;
        RECT 146.200 146.200 146.500 146.800 ;
        RECT 12.600 146.100 13.000 146.200 ;
        RECT 3.800 145.800 13.000 146.100 ;
        RECT 18.200 146.100 18.600 146.200 ;
        RECT 20.600 146.100 21.000 146.200 ;
        RECT 21.400 146.100 21.800 146.200 ;
        RECT 18.200 145.800 20.100 146.100 ;
        RECT 20.600 145.800 21.800 146.100 ;
        RECT 25.400 146.100 25.800 146.200 ;
        RECT 28.600 146.100 29.000 146.200 ;
        RECT 25.400 145.800 29.000 146.100 ;
        RECT 47.800 146.100 48.200 146.200 ;
        RECT 53.400 146.100 53.800 146.200 ;
        RECT 47.800 145.800 53.800 146.100 ;
        RECT 59.800 146.100 60.200 146.200 ;
        RECT 67.000 146.100 67.400 146.200 ;
        RECT 59.800 145.800 67.400 146.100 ;
        RECT 69.400 146.100 69.800 146.200 ;
        RECT 79.000 146.100 79.400 146.200 ;
        RECT 69.400 145.800 79.400 146.100 ;
        RECT 85.400 145.800 85.800 146.200 ;
        RECT 87.000 146.100 87.400 146.200 ;
        RECT 101.400 146.100 101.800 146.200 ;
        RECT 87.000 145.800 101.800 146.100 ;
        RECT 102.200 146.100 102.600 146.200 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 102.200 145.800 104.200 146.100 ;
        RECT 109.400 145.800 113.000 146.100 ;
        RECT 119.000 146.100 119.400 146.200 ;
        RECT 121.400 146.100 121.800 146.200 ;
        RECT 119.000 145.800 121.800 146.100 ;
        RECT 123.800 146.100 124.200 146.200 ;
        RECT 124.600 146.100 125.000 146.200 ;
        RECT 123.800 145.800 125.000 146.100 ;
        RECT 126.200 145.800 126.600 146.200 ;
        RECT 129.400 146.100 129.800 146.200 ;
        RECT 130.200 146.100 130.600 146.200 ;
        RECT 137.400 146.100 137.800 146.200 ;
        RECT 129.400 145.800 137.800 146.100 ;
        RECT 143.000 146.100 143.400 146.200 ;
        RECT 143.000 145.800 145.700 146.100 ;
        RECT 146.200 145.800 146.600 146.200 ;
        RECT 148.600 146.100 149.000 146.200 ;
        RECT 149.400 146.100 149.800 146.200 ;
        RECT 148.600 145.800 149.800 146.100 ;
        RECT 150.200 146.100 150.600 146.200 ;
        RECT 151.000 146.100 151.300 146.800 ;
        RECT 170.200 146.100 170.600 146.200 ;
        RECT 176.600 146.100 177.000 146.200 ;
        RECT 150.200 145.800 151.300 146.100 ;
        RECT 156.600 145.800 160.900 146.100 ;
        RECT 170.200 145.800 177.000 146.100 ;
        RECT 194.200 146.100 194.600 146.200 ;
        RECT 199.000 146.100 199.300 146.800 ;
        RECT 194.200 145.800 199.300 146.100 ;
        RECT 202.200 146.100 202.500 146.800 ;
        RECT 207.000 146.100 207.400 146.200 ;
        RECT 202.200 145.800 207.400 146.100 ;
        RECT 211.000 146.100 211.400 146.200 ;
        RECT 215.000 146.100 215.400 146.200 ;
        RECT 217.400 146.100 217.800 146.200 ;
        RECT 211.000 145.800 217.800 146.100 ;
        RECT 219.000 146.100 219.400 146.200 ;
        RECT 223.000 146.100 223.300 146.800 ;
        RECT 219.000 145.800 223.300 146.100 ;
        RECT 10.200 145.100 10.600 145.200 ;
        RECT 19.800 145.100 20.100 145.800 ;
        RECT 85.400 145.200 85.700 145.800 ;
        RECT 22.200 145.100 22.600 145.200 ;
        RECT 10.200 144.800 18.500 145.100 ;
        RECT 19.800 144.800 22.600 145.100 ;
        RECT 24.600 145.100 25.000 145.200 ;
        RECT 26.200 145.100 26.600 145.200 ;
        RECT 30.200 145.100 30.600 145.200 ;
        RECT 24.600 144.800 30.600 145.100 ;
        RECT 43.000 145.100 43.400 145.200 ;
        RECT 44.600 145.100 45.000 145.200 ;
        RECT 43.000 144.800 45.000 145.100 ;
        RECT 45.400 145.100 45.800 145.200 ;
        RECT 46.200 145.100 46.600 145.200 ;
        RECT 45.400 144.800 46.600 145.100 ;
        RECT 57.400 145.100 57.800 145.200 ;
        RECT 75.000 145.100 75.400 145.200 ;
        RECT 83.800 145.100 84.200 145.200 ;
        RECT 57.400 144.800 84.200 145.100 ;
        RECT 85.400 144.800 85.800 145.200 ;
        RECT 91.000 145.100 91.400 145.200 ;
        RECT 93.400 145.100 93.800 145.200 ;
        RECT 99.800 145.100 100.200 145.200 ;
        RECT 102.200 145.100 102.500 145.800 ;
        RECT 91.000 144.800 102.500 145.100 ;
        RECT 109.400 145.200 109.700 145.800 ;
        RECT 119.000 145.200 119.300 145.800 ;
        RECT 109.400 144.800 109.800 145.200 ;
        RECT 119.000 144.800 119.400 145.200 ;
        RECT 123.000 145.100 123.400 145.200 ;
        RECT 126.200 145.100 126.500 145.800 ;
        RECT 145.400 145.200 145.700 145.800 ;
        RECT 156.600 145.200 156.900 145.800 ;
        RECT 160.600 145.200 160.900 145.800 ;
        RECT 123.000 144.800 126.500 145.100 ;
        RECT 127.800 145.100 128.200 145.200 ;
        RECT 130.200 145.100 130.600 145.200 ;
        RECT 127.800 144.800 130.600 145.100 ;
        RECT 131.800 145.100 132.200 145.200 ;
        RECT 135.000 145.100 135.400 145.200 ;
        RECT 131.800 144.800 135.400 145.100 ;
        RECT 135.800 144.800 136.200 145.200 ;
        RECT 145.400 144.800 145.800 145.200 ;
        RECT 149.400 145.100 149.800 145.200 ;
        RECT 150.200 145.100 150.600 145.200 ;
        RECT 149.400 144.800 150.600 145.100 ;
        RECT 156.600 144.800 157.000 145.200 ;
        RECT 160.600 144.800 161.000 145.200 ;
        RECT 163.800 145.100 164.200 145.200 ;
        RECT 175.000 145.100 175.400 145.200 ;
        RECT 176.600 145.100 177.000 145.200 ;
        RECT 163.800 144.800 177.000 145.100 ;
        RECT 190.200 145.100 190.600 145.200 ;
        RECT 194.200 145.100 194.600 145.200 ;
        RECT 227.800 145.100 228.200 145.200 ;
        RECT 190.200 144.800 228.200 145.100 ;
        RECT 18.200 144.200 18.500 144.800 ;
        RECT 135.800 144.200 136.100 144.800 ;
        RECT 11.000 144.100 11.400 144.200 ;
        RECT 13.400 144.100 13.800 144.200 ;
        RECT 11.000 143.800 13.800 144.100 ;
        RECT 17.400 143.800 17.800 144.200 ;
        RECT 18.200 143.800 18.600 144.200 ;
        RECT 27.800 143.800 28.200 144.200 ;
        RECT 28.600 144.100 29.000 144.200 ;
        RECT 39.800 144.100 40.200 144.200 ;
        RECT 28.600 143.800 40.200 144.100 ;
        RECT 64.600 144.100 65.000 144.200 ;
        RECT 67.800 144.100 68.200 144.200 ;
        RECT 70.200 144.100 70.600 144.200 ;
        RECT 64.600 143.800 70.600 144.100 ;
        RECT 71.000 144.100 71.400 144.200 ;
        RECT 74.200 144.100 74.600 144.200 ;
        RECT 79.000 144.100 79.400 144.200 ;
        RECT 102.200 144.100 102.600 144.200 ;
        RECT 71.000 143.800 79.400 144.100 ;
        RECT 83.800 143.800 102.600 144.100 ;
        RECT 103.000 144.100 103.400 144.200 ;
        RECT 109.400 144.100 109.800 144.200 ;
        RECT 103.000 143.800 109.800 144.100 ;
        RECT 116.600 144.100 117.000 144.200 ;
        RECT 121.400 144.100 121.800 144.200 ;
        RECT 116.600 143.800 121.800 144.100 ;
        RECT 135.800 143.800 136.200 144.200 ;
        RECT 137.400 144.100 137.800 144.200 ;
        RECT 147.800 144.100 148.200 144.200 ;
        RECT 137.400 143.800 148.200 144.100 ;
        RECT 158.200 144.100 158.600 144.200 ;
        RECT 179.000 144.100 179.400 144.200 ;
        RECT 158.200 143.800 179.400 144.100 ;
        RECT 219.800 144.100 220.200 144.200 ;
        RECT 220.600 144.100 221.000 144.200 ;
        RECT 219.800 143.800 221.000 144.100 ;
        RECT 223.000 144.100 223.400 144.200 ;
        RECT 224.600 144.100 225.000 144.200 ;
        RECT 223.000 143.800 225.000 144.100 ;
        RECT 17.400 143.200 17.700 143.800 ;
        RECT 27.800 143.200 28.100 143.800 ;
        RECT 83.800 143.200 84.100 143.800 ;
        RECT 17.400 142.800 17.800 143.200 ;
        RECT 27.800 142.800 28.200 143.200 ;
        RECT 43.800 143.100 44.200 143.200 ;
        RECT 65.400 143.100 65.800 143.200 ;
        RECT 75.000 143.100 75.400 143.200 ;
        RECT 43.800 142.800 75.400 143.100 ;
        RECT 83.800 142.800 84.200 143.200 ;
        RECT 92.600 143.100 93.000 143.200 ;
        RECT 99.000 143.100 99.400 143.200 ;
        RECT 92.600 142.800 99.400 143.100 ;
        RECT 99.800 143.100 100.200 143.200 ;
        RECT 103.000 143.100 103.400 143.200 ;
        RECT 103.800 143.100 104.200 143.200 ;
        RECT 111.000 143.100 111.400 143.200 ;
        RECT 112.600 143.100 113.000 143.200 ;
        RECT 99.800 142.800 113.000 143.100 ;
        RECT 120.600 143.100 121.000 143.200 ;
        RECT 169.400 143.100 169.800 143.200 ;
        RECT 179.800 143.100 180.200 143.200 ;
        RECT 120.600 142.800 180.200 143.100 ;
        RECT 75.800 142.100 76.200 142.200 ;
        RECT 76.600 142.100 77.000 142.200 ;
        RECT 75.800 141.800 77.000 142.100 ;
        RECT 82.200 142.100 82.600 142.200 ;
        RECT 97.400 142.100 97.800 142.200 ;
        RECT 82.200 141.800 97.800 142.100 ;
        RECT 105.400 142.100 105.800 142.200 ;
        RECT 113.400 142.100 113.800 142.200 ;
        RECT 105.400 141.800 113.800 142.100 ;
        RECT 117.400 142.100 117.800 142.200 ;
        RECT 141.400 142.100 141.800 142.200 ;
        RECT 143.800 142.100 144.200 142.200 ;
        RECT 153.400 142.100 153.800 142.200 ;
        RECT 167.000 142.100 167.400 142.200 ;
        RECT 117.400 141.800 144.200 142.100 ;
        RECT 152.600 141.800 167.400 142.100 ;
        RECT 167.800 142.100 168.200 142.200 ;
        RECT 171.800 142.100 172.200 142.200 ;
        RECT 174.200 142.100 174.600 142.200 ;
        RECT 167.800 141.800 174.600 142.100 ;
        RECT 54.200 141.100 54.600 141.200 ;
        RECT 120.600 141.100 121.000 141.200 ;
        RECT 54.200 140.800 121.000 141.100 ;
        RECT 147.000 141.100 147.400 141.200 ;
        RECT 155.800 141.100 156.200 141.200 ;
        RECT 199.800 141.100 200.200 141.200 ;
        RECT 147.000 140.800 200.200 141.100 ;
        RECT 39.800 140.100 40.200 140.200 ;
        RECT 51.800 140.100 52.200 140.200 ;
        RECT 39.800 139.800 52.200 140.100 ;
        RECT 76.600 140.100 77.000 140.200 ;
        RECT 79.000 140.100 79.400 140.200 ;
        RECT 92.600 140.100 93.000 140.200 ;
        RECT 76.600 139.800 93.000 140.100 ;
        RECT 152.600 140.100 153.000 140.200 ;
        RECT 153.400 140.100 153.800 140.200 ;
        RECT 152.600 139.800 153.800 140.100 ;
        RECT 26.200 139.100 26.600 139.200 ;
        RECT 39.800 139.100 40.200 139.200 ;
        RECT 26.200 138.800 40.200 139.100 ;
        RECT 76.600 139.100 77.000 139.200 ;
        RECT 93.400 139.100 93.800 139.200 ;
        RECT 76.600 138.800 93.800 139.100 ;
        RECT 94.200 139.100 94.600 139.200 ;
        RECT 103.000 139.100 103.400 139.200 ;
        RECT 161.400 139.100 161.800 139.200 ;
        RECT 94.200 138.800 103.400 139.100 ;
        RECT 123.000 138.800 161.800 139.100 ;
        RECT 211.000 138.800 211.400 139.200 ;
        RECT 123.000 138.200 123.300 138.800 ;
        RECT 211.000 138.200 211.300 138.800 ;
        RECT 31.000 138.100 31.400 138.200 ;
        RECT 32.600 138.100 33.000 138.200 ;
        RECT 31.000 137.800 33.000 138.100 ;
        RECT 38.200 138.100 38.600 138.200 ;
        RECT 43.000 138.100 43.400 138.200 ;
        RECT 38.200 137.800 43.400 138.100 ;
        RECT 51.000 138.100 51.400 138.200 ;
        RECT 111.800 138.100 112.200 138.200 ;
        RECT 51.000 137.800 112.200 138.100 ;
        RECT 113.400 138.100 113.800 138.200 ;
        RECT 119.800 138.100 120.200 138.200 ;
        RECT 113.400 137.800 120.200 138.100 ;
        RECT 123.000 137.800 123.400 138.200 ;
        RECT 127.000 137.800 127.400 138.200 ;
        RECT 129.400 138.100 129.800 138.200 ;
        RECT 144.600 138.100 145.000 138.200 ;
        RECT 129.400 137.800 145.000 138.100 ;
        RECT 154.200 138.100 154.600 138.200 ;
        RECT 163.800 138.100 164.200 138.200 ;
        RECT 154.200 137.800 164.200 138.100 ;
        RECT 211.000 137.800 211.400 138.200 ;
        RECT 127.000 137.200 127.300 137.800 ;
        RECT 27.800 136.800 28.200 137.200 ;
        RECT 34.200 137.100 34.600 137.200 ;
        RECT 51.000 137.100 51.400 137.200 ;
        RECT 34.200 136.800 51.400 137.100 ;
        RECT 62.200 136.800 62.600 137.200 ;
        RECT 81.400 137.100 81.800 137.200 ;
        RECT 94.200 137.100 94.600 137.200 ;
        RECT 81.400 136.800 94.600 137.100 ;
        RECT 101.400 137.100 101.800 137.200 ;
        RECT 105.400 137.100 105.800 137.200 ;
        RECT 121.400 137.100 121.800 137.200 ;
        RECT 101.400 136.800 105.800 137.100 ;
        RECT 117.400 136.800 121.800 137.100 ;
        RECT 127.000 136.800 127.400 137.200 ;
        RECT 131.000 136.800 131.400 137.200 ;
        RECT 132.600 137.100 133.000 137.200 ;
        RECT 135.800 137.100 136.200 137.200 ;
        RECT 132.600 136.800 136.200 137.100 ;
        RECT 143.000 136.800 143.400 137.200 ;
        RECT 145.400 137.100 145.800 137.200 ;
        RECT 154.200 137.100 154.600 137.200 ;
        RECT 155.800 137.100 156.200 137.200 ;
        RECT 145.400 136.800 156.200 137.100 ;
        RECT 172.600 137.100 173.000 137.200 ;
        RECT 179.800 137.100 180.200 137.200 ;
        RECT 187.800 137.100 188.200 137.200 ;
        RECT 172.600 136.800 180.200 137.100 ;
        RECT 184.600 136.800 188.200 137.100 ;
        RECT 197.400 136.800 197.800 137.200 ;
        RECT 198.200 136.800 198.600 137.200 ;
        RECT 203.000 137.100 203.400 137.200 ;
        RECT 207.800 137.100 208.200 137.200 ;
        RECT 203.000 136.800 208.200 137.100 ;
        RECT 20.600 136.100 21.000 136.200 ;
        RECT 27.000 136.100 27.400 136.200 ;
        RECT 20.600 135.800 27.400 136.100 ;
        RECT 27.800 136.100 28.100 136.800 ;
        RECT 62.200 136.200 62.500 136.800 ;
        RECT 117.400 136.200 117.700 136.800 ;
        RECT 31.800 136.100 32.200 136.200 ;
        RECT 27.800 135.800 32.200 136.100 ;
        RECT 39.800 136.100 40.200 136.200 ;
        RECT 43.800 136.100 44.200 136.200 ;
        RECT 39.800 135.800 44.200 136.100 ;
        RECT 62.200 135.800 62.600 136.200 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 71.800 136.100 72.200 136.200 ;
        RECT 72.600 136.100 73.000 136.200 ;
        RECT 71.800 135.800 73.000 136.100 ;
        RECT 85.400 136.100 85.800 136.200 ;
        RECT 94.200 136.100 94.600 136.200 ;
        RECT 85.400 135.800 94.600 136.100 ;
        RECT 103.000 136.100 103.400 136.200 ;
        RECT 106.200 136.100 106.600 136.200 ;
        RECT 103.000 135.800 106.600 136.100 ;
        RECT 116.600 136.100 117.000 136.200 ;
        RECT 117.400 136.100 117.800 136.200 ;
        RECT 116.600 135.800 117.800 136.100 ;
        RECT 119.800 136.100 120.200 136.200 ;
        RECT 124.600 136.100 125.000 136.200 ;
        RECT 127.800 136.100 128.200 136.200 ;
        RECT 131.000 136.100 131.300 136.800 ;
        RECT 119.800 135.800 131.300 136.100 ;
        RECT 135.000 135.800 135.400 136.200 ;
        RECT 140.600 136.100 141.000 136.200 ;
        RECT 141.400 136.100 141.800 136.200 ;
        RECT 140.600 135.800 141.800 136.100 ;
        RECT 143.000 136.100 143.300 136.800 ;
        RECT 184.600 136.200 184.900 136.800 ;
        RECT 197.400 136.200 197.700 136.800 ;
        RECT 198.200 136.200 198.500 136.800 ;
        RECT 144.600 136.100 145.000 136.200 ;
        RECT 143.000 135.800 145.000 136.100 ;
        RECT 145.400 136.100 145.800 136.200 ;
        RECT 147.800 136.100 148.200 136.200 ;
        RECT 145.400 135.800 148.200 136.100 ;
        RECT 156.600 136.100 157.000 136.200 ;
        RECT 158.200 136.100 158.600 136.200 ;
        RECT 156.600 135.800 158.600 136.100 ;
        RECT 178.200 136.100 178.600 136.200 ;
        RECT 184.600 136.100 185.000 136.200 ;
        RECT 178.200 135.800 185.000 136.100 ;
        RECT 186.200 136.100 186.600 136.200 ;
        RECT 192.600 136.100 193.000 136.200 ;
        RECT 186.200 135.800 193.000 136.100 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 198.200 135.800 198.600 136.200 ;
        RECT 200.600 136.100 201.000 136.200 ;
        RECT 206.200 136.100 206.600 136.200 ;
        RECT 207.800 136.100 208.200 136.200 ;
        RECT 214.200 136.100 214.600 136.200 ;
        RECT 200.600 135.800 206.600 136.100 ;
        RECT 207.000 135.800 214.600 136.100 ;
        RECT 63.000 135.200 63.300 135.800 ;
        RECT 11.800 135.100 12.200 135.200 ;
        RECT 15.000 135.100 15.400 135.200 ;
        RECT 23.000 135.100 23.400 135.200 ;
        RECT 11.800 134.800 23.400 135.100 ;
        RECT 24.600 135.100 25.000 135.200 ;
        RECT 25.400 135.100 25.800 135.200 ;
        RECT 24.600 134.800 25.800 135.100 ;
        RECT 29.400 134.800 29.800 135.200 ;
        RECT 33.400 135.100 33.800 135.200 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 33.400 134.800 41.000 135.100 ;
        RECT 45.400 135.100 45.800 135.200 ;
        RECT 49.400 135.100 49.800 135.200 ;
        RECT 45.400 134.800 49.800 135.100 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 64.600 134.800 65.000 135.200 ;
        RECT 68.600 135.100 69.000 135.200 ;
        RECT 72.600 135.100 73.000 135.200 ;
        RECT 68.600 134.800 73.000 135.100 ;
        RECT 78.200 135.100 78.600 135.200 ;
        RECT 79.800 135.100 80.200 135.200 ;
        RECT 80.600 135.100 81.000 135.200 ;
        RECT 78.200 134.800 81.000 135.100 ;
        RECT 84.600 135.100 85.000 135.200 ;
        RECT 90.200 135.100 90.600 135.200 ;
        RECT 84.600 134.800 90.600 135.100 ;
        RECT 92.600 135.100 93.000 135.200 ;
        RECT 96.600 135.100 97.000 135.200 ;
        RECT 92.600 134.800 97.000 135.100 ;
        RECT 99.000 135.100 99.400 135.200 ;
        RECT 101.400 135.100 101.800 135.200 ;
        RECT 99.000 134.800 101.800 135.100 ;
        RECT 102.200 135.100 102.600 135.200 ;
        RECT 104.600 135.100 105.000 135.200 ;
        RECT 105.400 135.100 105.800 135.200 ;
        RECT 108.600 135.100 109.000 135.200 ;
        RECT 102.200 134.800 109.000 135.100 ;
        RECT 115.000 135.100 115.400 135.200 ;
        RECT 119.800 135.100 120.100 135.800 ;
        RECT 135.000 135.200 135.300 135.800 ;
        RECT 115.000 134.800 120.100 135.100 ;
        RECT 123.800 135.100 124.200 135.200 ;
        RECT 127.000 135.100 127.400 135.200 ;
        RECT 127.800 135.100 128.200 135.200 ;
        RECT 123.800 134.800 128.200 135.100 ;
        RECT 135.000 134.800 135.400 135.200 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 139.000 135.100 139.400 135.200 ;
        RECT 138.200 134.800 139.400 135.100 ;
        RECT 143.800 135.100 144.200 135.200 ;
        RECT 151.000 135.100 151.400 135.200 ;
        RECT 173.400 135.100 173.800 135.200 ;
        RECT 176.600 135.100 177.000 135.200 ;
        RECT 143.800 134.800 177.000 135.100 ;
        RECT 178.200 135.100 178.600 135.200 ;
        RECT 180.600 135.100 181.000 135.200 ;
        RECT 182.200 135.100 182.600 135.200 ;
        RECT 204.600 135.100 205.000 135.200 ;
        RECT 206.200 135.100 206.600 135.200 ;
        RECT 178.200 134.800 206.600 135.100 ;
        RECT 207.000 135.100 207.400 135.200 ;
        RECT 207.800 135.100 208.200 135.200 ;
        RECT 207.000 134.800 208.200 135.100 ;
        RECT 3.800 134.100 4.200 134.200 ;
        RECT 12.600 134.100 13.000 134.200 ;
        RECT 3.800 133.800 13.000 134.100 ;
        RECT 21.400 134.100 21.800 134.200 ;
        RECT 29.400 134.100 29.700 134.800 ;
        RECT 21.400 133.800 29.700 134.100 ;
        RECT 35.800 134.100 36.200 134.200 ;
        RECT 39.000 134.100 39.400 134.200 ;
        RECT 35.800 133.800 39.400 134.100 ;
        RECT 43.000 134.100 43.400 134.200 ;
        RECT 44.600 134.100 45.000 134.200 ;
        RECT 43.000 133.800 45.000 134.100 ;
        RECT 46.200 134.100 46.600 134.200 ;
        RECT 48.600 134.100 49.000 134.200 ;
        RECT 46.200 133.800 49.000 134.100 ;
        RECT 57.400 134.100 57.800 134.200 ;
        RECT 64.600 134.100 64.900 134.800 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 57.400 133.800 64.900 134.100 ;
        RECT 75.000 134.100 75.400 134.200 ;
        RECT 79.800 134.100 80.200 134.200 ;
        RECT 75.000 133.800 80.200 134.100 ;
        RECT 83.000 134.100 83.400 134.200 ;
        RECT 95.000 134.100 95.400 134.200 ;
        RECT 83.000 133.800 95.400 134.100 ;
        RECT 101.400 134.100 101.800 134.200 ;
        RECT 111.000 134.100 111.400 134.200 ;
        RECT 101.400 133.800 111.400 134.100 ;
        RECT 113.400 134.100 113.800 134.200 ;
        RECT 115.800 134.100 116.200 134.200 ;
        RECT 119.000 134.100 119.400 134.200 ;
        RECT 113.400 133.800 119.400 134.100 ;
        RECT 123.800 134.100 124.200 134.200 ;
        RECT 125.400 134.100 125.800 134.200 ;
        RECT 123.800 133.800 125.800 134.100 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 137.400 134.100 137.800 134.200 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 141.400 134.100 141.800 134.200 ;
        RECT 137.400 133.800 141.800 134.100 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 146.200 134.100 146.600 134.200 ;
        RECT 160.600 134.100 161.000 134.200 ;
        RECT 146.200 133.800 161.000 134.100 ;
        RECT 163.000 134.100 163.400 134.200 ;
        RECT 164.600 134.100 165.000 134.200 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 168.600 134.100 169.000 134.200 ;
        RECT 163.000 133.800 165.000 134.100 ;
        RECT 166.200 133.800 169.000 134.100 ;
        RECT 176.600 134.100 177.000 134.200 ;
        RECT 177.400 134.100 177.800 134.200 ;
        RECT 176.600 133.800 177.800 134.100 ;
        RECT 183.000 134.100 183.400 134.200 ;
        RECT 183.800 134.100 184.200 134.200 ;
        RECT 207.000 134.100 207.400 134.200 ;
        RECT 218.200 134.100 218.600 134.200 ;
        RECT 228.600 134.100 229.000 134.200 ;
        RECT 183.000 133.800 229.000 134.100 ;
        RECT 25.400 133.100 25.800 133.200 ;
        RECT 78.200 133.100 78.600 133.200 ;
        RECT 82.200 133.100 82.600 133.200 ;
        RECT 25.400 132.800 82.600 133.100 ;
        RECT 97.400 133.100 97.800 133.200 ;
        RECT 107.000 133.100 107.400 133.200 ;
        RECT 110.200 133.100 110.600 133.200 ;
        RECT 97.400 132.800 110.600 133.100 ;
        RECT 111.000 133.100 111.300 133.800 ;
        RECT 143.800 133.200 144.100 133.800 ;
        RECT 124.600 133.100 125.000 133.200 ;
        RECT 111.000 132.800 125.000 133.100 ;
        RECT 128.600 133.100 129.000 133.200 ;
        RECT 143.000 133.100 143.400 133.200 ;
        RECT 128.600 132.800 143.400 133.100 ;
        RECT 143.800 132.800 144.200 133.200 ;
        RECT 144.600 133.100 145.000 133.200 ;
        RECT 147.000 133.100 147.400 133.200 ;
        RECT 144.600 132.800 147.400 133.100 ;
        RECT 157.400 133.100 157.800 133.200 ;
        RECT 158.200 133.100 158.600 133.200 ;
        RECT 170.200 133.100 170.600 133.200 ;
        RECT 157.400 132.800 170.600 133.100 ;
        RECT 173.400 133.100 173.800 133.200 ;
        RECT 174.200 133.100 174.600 133.200 ;
        RECT 189.400 133.100 189.800 133.200 ;
        RECT 173.400 132.800 189.800 133.100 ;
        RECT 194.200 133.100 194.600 133.200 ;
        RECT 195.800 133.100 196.200 133.200 ;
        RECT 194.200 132.800 196.200 133.100 ;
        RECT 201.400 132.800 201.800 133.200 ;
        RECT 203.800 133.100 204.200 133.200 ;
        RECT 221.400 133.100 221.800 133.200 ;
        RECT 203.800 132.800 221.800 133.100 ;
        RECT 13.400 132.100 13.800 132.200 ;
        RECT 19.000 132.100 19.400 132.200 ;
        RECT 47.000 132.100 47.400 132.200 ;
        RECT 13.400 131.800 47.400 132.100 ;
        RECT 56.600 132.100 57.000 132.200 ;
        RECT 59.800 132.100 60.200 132.200 ;
        RECT 56.600 131.800 60.200 132.100 ;
        RECT 73.400 132.100 73.800 132.200 ;
        RECT 75.000 132.100 75.400 132.200 ;
        RECT 73.400 131.800 75.400 132.100 ;
        RECT 79.000 132.100 79.400 132.200 ;
        RECT 112.600 132.100 113.000 132.200 ;
        RECT 118.200 132.100 118.600 132.200 ;
        RECT 79.000 131.800 118.600 132.100 ;
        RECT 124.600 132.100 125.000 132.200 ;
        RECT 132.600 132.100 133.000 132.200 ;
        RECT 149.400 132.100 149.800 132.200 ;
        RECT 124.600 131.800 149.800 132.100 ;
        RECT 156.600 132.100 157.000 132.200 ;
        RECT 171.000 132.100 171.400 132.200 ;
        RECT 156.600 131.800 171.400 132.100 ;
        RECT 193.400 132.100 193.800 132.200 ;
        RECT 201.400 132.100 201.700 132.800 ;
        RECT 193.400 131.800 201.700 132.100 ;
        RECT 207.000 132.100 207.400 132.200 ;
        RECT 226.200 132.100 226.600 132.200 ;
        RECT 207.000 131.800 226.600 132.100 ;
        RECT 15.000 130.800 15.400 131.200 ;
        RECT 47.800 131.100 48.200 131.200 ;
        RECT 61.400 131.100 61.800 131.200 ;
        RECT 47.800 130.800 61.800 131.100 ;
        RECT 95.000 131.100 95.400 131.200 ;
        RECT 115.800 131.100 116.200 131.200 ;
        RECT 95.000 130.800 116.200 131.100 ;
        RECT 116.600 131.100 117.000 131.200 ;
        RECT 137.400 131.100 137.800 131.200 ;
        RECT 116.600 130.800 137.800 131.100 ;
        RECT 138.200 131.100 138.600 131.200 ;
        RECT 145.400 131.100 145.800 131.200 ;
        RECT 159.800 131.100 160.200 131.200 ;
        RECT 163.800 131.100 164.200 131.200 ;
        RECT 138.200 130.800 145.800 131.100 ;
        RECT 147.800 130.800 164.200 131.100 ;
        RECT 167.000 131.100 167.400 131.200 ;
        RECT 190.200 131.100 190.600 131.200 ;
        RECT 167.000 130.800 190.600 131.100 ;
        RECT 195.800 131.100 196.200 131.200 ;
        RECT 196.600 131.100 197.000 131.200 ;
        RECT 195.800 130.800 197.000 131.100 ;
        RECT 197.400 131.100 197.800 131.200 ;
        RECT 208.600 131.100 209.000 131.200 ;
        RECT 197.400 130.800 209.000 131.100 ;
        RECT 15.000 130.200 15.300 130.800 ;
        RECT 3.000 130.100 3.400 130.200 ;
        RECT 15.000 130.100 15.400 130.200 ;
        RECT 3.000 129.800 15.400 130.100 ;
        RECT 51.000 130.100 51.400 130.200 ;
        RECT 66.200 130.100 66.600 130.200 ;
        RECT 76.600 130.100 77.000 130.200 ;
        RECT 51.000 129.800 77.000 130.100 ;
        RECT 111.800 130.100 112.200 130.200 ;
        RECT 113.400 130.100 113.800 130.200 ;
        RECT 111.800 129.800 113.800 130.100 ;
        RECT 115.000 130.100 115.400 130.200 ;
        RECT 147.800 130.100 148.100 130.800 ;
        RECT 115.000 129.800 148.100 130.100 ;
        RECT 148.600 130.100 149.000 130.200 ;
        RECT 152.600 130.100 153.000 130.200 ;
        RECT 159.000 130.100 159.400 130.200 ;
        RECT 148.600 129.800 159.400 130.100 ;
        RECT 165.400 130.100 165.800 130.200 ;
        RECT 169.400 130.100 169.800 130.200 ;
        RECT 165.400 129.800 169.800 130.100 ;
        RECT 199.800 130.100 200.200 130.200 ;
        RECT 207.800 130.100 208.200 130.200 ;
        RECT 199.800 129.800 208.200 130.100 ;
        RECT 10.200 129.100 10.600 129.200 ;
        RECT 13.400 129.100 13.800 129.200 ;
        RECT 10.200 128.800 13.800 129.100 ;
        RECT 43.000 129.100 43.400 129.200 ;
        RECT 47.800 129.100 48.200 129.200 ;
        RECT 55.000 129.100 55.400 129.200 ;
        RECT 43.000 128.800 48.200 129.100 ;
        RECT 53.400 128.800 55.400 129.100 ;
        RECT 74.200 128.800 74.600 129.200 ;
        RECT 99.000 129.100 99.400 129.200 ;
        RECT 127.800 129.100 128.200 129.200 ;
        RECT 99.000 128.800 128.200 129.100 ;
        RECT 142.200 129.100 142.600 129.200 ;
        RECT 145.400 129.100 145.800 129.200 ;
        RECT 142.200 128.800 145.800 129.100 ;
        RECT 183.000 129.100 183.400 129.200 ;
        RECT 190.200 129.100 190.600 129.200 ;
        RECT 203.000 129.100 203.400 129.200 ;
        RECT 183.000 128.800 189.700 129.100 ;
        RECT 190.200 128.800 203.400 129.100 ;
        RECT 213.400 129.100 213.800 129.200 ;
        RECT 218.200 129.100 218.600 129.200 ;
        RECT 213.400 128.800 218.600 129.100 ;
        RECT 53.400 128.200 53.700 128.800 ;
        RECT 4.600 128.100 5.000 128.200 ;
        RECT 11.800 128.100 12.200 128.200 ;
        RECT 4.600 127.800 12.200 128.100 ;
        RECT 19.800 128.100 20.200 128.200 ;
        RECT 23.800 128.100 24.200 128.200 ;
        RECT 19.800 127.800 24.200 128.100 ;
        RECT 47.800 128.100 48.200 128.200 ;
        RECT 48.600 128.100 49.000 128.200 ;
        RECT 47.800 127.800 49.000 128.100 ;
        RECT 53.400 127.800 53.800 128.200 ;
        RECT 55.800 128.100 56.200 128.200 ;
        RECT 63.000 128.100 63.400 128.200 ;
        RECT 55.800 127.800 63.400 128.100 ;
        RECT 74.200 128.100 74.500 128.800 ;
        RECT 189.400 128.200 189.700 128.800 ;
        RECT 75.800 128.100 76.200 128.200 ;
        RECT 106.200 128.100 106.600 128.200 ;
        RECT 74.200 127.800 76.200 128.100 ;
        RECT 77.400 127.800 106.600 128.100 ;
        RECT 109.400 128.100 109.800 128.200 ;
        RECT 116.600 128.100 117.000 128.200 ;
        RECT 109.400 127.800 117.000 128.100 ;
        RECT 121.400 128.100 121.800 128.200 ;
        RECT 129.400 128.100 129.800 128.200 ;
        RECT 121.400 127.800 129.800 128.100 ;
        RECT 134.200 128.100 134.600 128.200 ;
        RECT 138.200 128.100 138.600 128.200 ;
        RECT 134.200 127.800 138.600 128.100 ;
        RECT 144.600 127.800 145.000 128.200 ;
        RECT 151.800 128.100 152.200 128.200 ;
        RECT 179.000 128.100 179.400 128.200 ;
        RECT 151.800 127.800 179.400 128.100 ;
        RECT 187.800 127.800 188.200 128.200 ;
        RECT 189.400 127.800 189.800 128.200 ;
        RECT 200.600 128.100 201.000 128.200 ;
        RECT 211.000 128.100 211.400 128.200 ;
        RECT 200.600 127.800 211.400 128.100 ;
        RECT 11.800 127.100 12.100 127.800 ;
        RECT 77.400 127.200 77.700 127.800 ;
        RECT 18.200 127.100 18.600 127.200 ;
        RECT 48.600 127.100 49.000 127.200 ;
        RECT 11.800 126.800 18.600 127.100 ;
        RECT 31.800 126.800 49.000 127.100 ;
        RECT 51.000 127.100 51.400 127.200 ;
        RECT 53.400 127.100 53.800 127.200 ;
        RECT 51.000 126.800 53.800 127.100 ;
        RECT 54.200 127.100 54.600 127.200 ;
        RECT 63.800 127.100 64.200 127.200 ;
        RECT 64.600 127.100 65.000 127.200 ;
        RECT 54.200 126.800 65.000 127.100 ;
        RECT 77.400 126.800 77.800 127.200 ;
        RECT 81.400 127.100 81.800 127.200 ;
        RECT 86.200 127.100 86.600 127.200 ;
        RECT 81.400 126.800 86.600 127.100 ;
        RECT 99.000 127.100 99.400 127.200 ;
        RECT 101.400 127.100 101.800 127.200 ;
        RECT 103.000 127.100 103.400 127.200 ;
        RECT 103.800 127.100 104.200 127.200 ;
        RECT 99.000 126.800 104.200 127.100 ;
        RECT 108.600 127.100 109.000 127.200 ;
        RECT 114.200 127.100 114.600 127.200 ;
        RECT 108.600 126.800 114.600 127.100 ;
        RECT 115.000 127.100 115.400 127.200 ;
        RECT 117.400 127.100 117.800 127.200 ;
        RECT 119.800 127.100 120.200 127.200 ;
        RECT 115.000 126.800 120.200 127.100 ;
        RECT 135.800 126.800 136.200 127.200 ;
        RECT 143.000 127.100 143.400 127.200 ;
        RECT 143.800 127.100 144.200 127.200 ;
        RECT 143.000 126.800 144.200 127.100 ;
        RECT 144.600 127.100 144.900 127.800 ;
        RECT 147.000 127.100 147.400 127.200 ;
        RECT 144.600 126.800 147.400 127.100 ;
        RECT 159.000 127.100 159.400 127.200 ;
        RECT 163.000 127.100 163.400 127.200 ;
        RECT 159.000 126.800 163.400 127.100 ;
        RECT 165.400 127.100 165.800 127.200 ;
        RECT 174.200 127.100 174.600 127.200 ;
        RECT 165.400 126.800 174.600 127.100 ;
        RECT 177.400 127.100 177.800 127.200 ;
        RECT 183.800 127.100 184.200 127.200 ;
        RECT 177.400 126.800 184.200 127.100 ;
        RECT 187.800 127.100 188.100 127.800 ;
        RECT 196.600 127.100 197.000 127.200 ;
        RECT 187.800 126.800 197.000 127.100 ;
        RECT 210.200 126.800 210.600 127.200 ;
        RECT 217.400 127.100 217.800 127.200 ;
        RECT 218.200 127.100 218.600 127.200 ;
        RECT 217.400 126.800 218.600 127.100 ;
        RECT 31.800 126.200 32.100 126.800 ;
        RECT 3.000 126.100 3.400 126.200 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 3.000 125.800 13.800 126.100 ;
        RECT 19.800 126.100 20.200 126.200 ;
        RECT 28.600 126.100 29.000 126.200 ;
        RECT 19.800 125.800 29.000 126.100 ;
        RECT 31.800 125.800 32.200 126.200 ;
        RECT 36.600 126.100 37.000 126.200 ;
        RECT 44.600 126.100 45.000 126.200 ;
        RECT 36.600 125.800 45.000 126.100 ;
        RECT 52.600 126.100 53.000 126.200 ;
        RECT 54.200 126.100 54.600 126.200 ;
        RECT 52.600 125.800 54.600 126.100 ;
        RECT 55.800 126.100 56.200 126.200 ;
        RECT 59.800 126.100 60.200 126.200 ;
        RECT 60.600 126.100 61.000 126.200 ;
        RECT 55.800 125.800 61.000 126.100 ;
        RECT 92.600 126.100 93.000 126.200 ;
        RECT 100.600 126.100 101.000 126.200 ;
        RECT 92.600 125.800 101.000 126.100 ;
        RECT 101.400 126.100 101.800 126.200 ;
        RECT 118.200 126.100 118.600 126.200 ;
        RECT 101.400 125.800 118.600 126.100 ;
        RECT 119.800 126.100 120.200 126.200 ;
        RECT 120.600 126.100 121.000 126.200 ;
        RECT 123.800 126.100 124.200 126.200 ;
        RECT 119.800 125.800 124.200 126.100 ;
        RECT 130.200 126.100 130.600 126.200 ;
        RECT 135.800 126.100 136.100 126.800 ;
        RECT 210.200 126.200 210.500 126.800 ;
        RECT 130.200 125.800 136.100 126.100 ;
        RECT 143.000 126.100 143.400 126.200 ;
        RECT 149.400 126.100 149.800 126.200 ;
        RECT 143.000 125.800 149.800 126.100 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 168.600 126.100 169.000 126.200 ;
        RECT 180.600 126.100 181.000 126.200 ;
        RECT 168.600 125.800 181.000 126.100 ;
        RECT 188.600 126.100 189.000 126.200 ;
        RECT 190.200 126.100 190.600 126.200 ;
        RECT 188.600 125.800 190.600 126.100 ;
        RECT 191.000 126.100 191.400 126.200 ;
        RECT 199.000 126.100 199.400 126.200 ;
        RECT 203.000 126.100 203.400 126.200 ;
        RECT 204.600 126.100 205.000 126.200 ;
        RECT 207.800 126.100 208.200 126.200 ;
        RECT 191.000 125.800 200.100 126.100 ;
        RECT 203.000 125.800 208.200 126.100 ;
        RECT 210.200 125.800 210.600 126.200 ;
        RECT 217.400 126.100 217.800 126.200 ;
        RECT 223.800 126.100 224.200 126.200 ;
        RECT 216.600 125.800 224.200 126.100 ;
        RECT 9.400 125.100 9.800 125.200 ;
        RECT 2.200 124.800 9.800 125.100 ;
        RECT 11.800 125.100 12.200 125.200 ;
        RECT 26.200 125.100 26.600 125.200 ;
        RECT 44.600 125.100 45.000 125.200 ;
        RECT 11.800 124.800 45.000 125.100 ;
        RECT 63.000 125.100 63.400 125.200 ;
        RECT 79.000 125.100 79.400 125.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 63.000 124.800 82.600 125.100 ;
        RECT 96.600 125.100 97.000 125.200 ;
        RECT 99.800 125.100 100.200 125.200 ;
        RECT 96.600 124.800 100.200 125.100 ;
        RECT 100.600 125.100 101.000 125.200 ;
        RECT 103.000 125.100 103.400 125.200 ;
        RECT 100.600 124.800 103.400 125.100 ;
        RECT 103.800 125.100 104.200 125.200 ;
        RECT 111.000 125.100 111.400 125.200 ;
        RECT 103.800 124.800 111.400 125.100 ;
        RECT 111.800 125.100 112.200 125.200 ;
        RECT 114.200 125.100 114.600 125.200 ;
        RECT 111.800 124.800 114.600 125.100 ;
        RECT 115.000 125.100 115.400 125.200 ;
        RECT 116.600 125.100 117.000 125.200 ;
        RECT 117.400 125.100 117.800 125.200 ;
        RECT 115.000 124.800 117.800 125.100 ;
        RECT 118.200 125.100 118.600 125.200 ;
        RECT 121.400 125.100 121.800 125.200 ;
        RECT 118.200 124.800 121.800 125.100 ;
        RECT 124.600 125.100 125.000 125.200 ;
        RECT 135.000 125.100 135.400 125.200 ;
        RECT 136.600 125.100 137.000 125.200 ;
        RECT 124.600 124.800 137.000 125.100 ;
        RECT 138.200 125.100 138.600 125.200 ;
        RECT 139.000 125.100 139.400 125.200 ;
        RECT 146.200 125.100 146.600 125.200 ;
        RECT 138.200 124.800 146.600 125.100 ;
        RECT 160.600 125.100 161.000 125.200 ;
        RECT 162.200 125.100 162.500 125.800 ;
        RECT 160.600 124.800 162.500 125.100 ;
        RECT 168.600 125.100 169.000 125.200 ;
        RECT 169.400 125.100 169.800 125.200 ;
        RECT 168.600 124.800 169.800 125.100 ;
        RECT 170.200 125.100 170.600 125.200 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 170.200 124.800 171.400 125.100 ;
        RECT 185.400 125.100 185.800 125.200 ;
        RECT 198.200 125.100 198.600 125.200 ;
        RECT 203.000 125.100 203.400 125.200 ;
        RECT 185.400 124.800 189.700 125.100 ;
        RECT 198.200 124.800 203.400 125.100 ;
        RECT 215.800 125.100 216.200 125.200 ;
        RECT 218.200 125.100 218.600 125.200 ;
        RECT 215.800 124.800 218.600 125.100 ;
        RECT 2.200 124.200 2.500 124.800 ;
        RECT 189.400 124.200 189.700 124.800 ;
        RECT 2.200 123.800 2.600 124.200 ;
        RECT 81.400 124.100 81.800 124.200 ;
        RECT 91.800 124.100 92.200 124.200 ;
        RECT 103.000 124.100 103.400 124.200 ;
        RECT 81.400 123.800 103.400 124.100 ;
        RECT 104.600 124.100 105.000 124.200 ;
        RECT 107.000 124.100 107.400 124.200 ;
        RECT 104.600 123.800 107.400 124.100 ;
        RECT 107.800 124.100 108.200 124.200 ;
        RECT 110.200 124.100 110.600 124.200 ;
        RECT 141.400 124.100 141.800 124.200 ;
        RECT 107.800 123.800 141.800 124.100 ;
        RECT 142.200 124.100 142.600 124.200 ;
        RECT 147.800 124.100 148.200 124.200 ;
        RECT 142.200 123.800 148.200 124.100 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 166.200 124.100 166.600 124.200 ;
        RECT 165.400 123.800 166.600 124.100 ;
        RECT 167.000 124.100 167.400 124.200 ;
        RECT 183.800 124.100 184.200 124.200 ;
        RECT 167.000 123.800 184.200 124.100 ;
        RECT 189.400 123.800 189.800 124.200 ;
        RECT 225.400 124.100 225.800 124.200 ;
        RECT 229.400 124.100 229.800 124.200 ;
        RECT 225.400 123.800 229.800 124.100 ;
        RECT 31.000 123.100 31.400 123.200 ;
        RECT 47.000 123.100 47.400 123.200 ;
        RECT 49.400 123.100 49.800 123.200 ;
        RECT 31.000 122.800 49.800 123.100 ;
        RECT 67.000 123.100 67.400 123.200 ;
        RECT 124.600 123.100 125.000 123.200 ;
        RECT 67.000 122.800 125.000 123.100 ;
        RECT 126.200 123.100 126.600 123.200 ;
        RECT 164.600 123.100 165.000 123.200 ;
        RECT 175.000 123.100 175.400 123.200 ;
        RECT 177.400 123.100 177.800 123.200 ;
        RECT 126.200 122.800 177.800 123.100 ;
        RECT 24.600 122.100 25.000 122.200 ;
        RECT 29.400 122.100 29.800 122.200 ;
        RECT 24.600 121.800 29.800 122.100 ;
        RECT 108.600 122.100 109.000 122.200 ;
        RECT 110.200 122.100 110.600 122.200 ;
        RECT 108.600 121.800 110.600 122.100 ;
        RECT 112.600 122.100 113.000 122.200 ;
        RECT 115.800 122.100 116.200 122.200 ;
        RECT 112.600 121.800 116.200 122.100 ;
        RECT 119.800 122.100 120.200 122.200 ;
        RECT 135.800 122.100 136.200 122.200 ;
        RECT 143.800 122.100 144.200 122.200 ;
        RECT 119.800 121.800 144.200 122.100 ;
        RECT 188.600 122.100 189.000 122.200 ;
        RECT 202.200 122.100 202.600 122.200 ;
        RECT 205.400 122.100 205.800 122.200 ;
        RECT 188.600 121.800 205.800 122.100 ;
        RECT 97.400 121.100 97.800 121.200 ;
        RECT 105.400 121.100 105.800 121.200 ;
        RECT 97.400 120.800 105.800 121.100 ;
        RECT 107.800 121.100 108.200 121.200 ;
        RECT 119.800 121.100 120.200 121.200 ;
        RECT 137.400 121.100 137.800 121.200 ;
        RECT 107.800 120.800 119.300 121.100 ;
        RECT 119.800 120.800 137.800 121.100 ;
        RECT 142.200 121.100 142.600 121.200 ;
        RECT 155.800 121.100 156.200 121.200 ;
        RECT 142.200 120.800 156.200 121.100 ;
        RECT 83.000 120.100 83.400 120.200 ;
        RECT 92.600 120.100 93.000 120.200 ;
        RECT 102.200 120.100 102.600 120.200 ;
        RECT 83.000 119.800 102.600 120.100 ;
        RECT 108.600 120.100 109.000 120.200 ;
        RECT 113.400 120.100 113.800 120.200 ;
        RECT 108.600 119.800 113.800 120.100 ;
        RECT 119.000 120.100 119.300 120.800 ;
        RECT 135.000 120.100 135.400 120.200 ;
        RECT 119.000 119.800 135.400 120.100 ;
        RECT 153.400 120.100 153.800 120.200 ;
        RECT 162.200 120.100 162.600 120.200 ;
        RECT 153.400 119.800 162.600 120.100 ;
        RECT 186.200 120.100 186.600 120.200 ;
        RECT 189.400 120.100 189.800 120.200 ;
        RECT 186.200 119.800 189.800 120.100 ;
        RECT 14.200 119.100 14.600 119.200 ;
        RECT 126.200 119.100 126.600 119.200 ;
        RECT 14.200 118.800 126.600 119.100 ;
        RECT 146.200 119.100 146.600 119.200 ;
        RECT 164.600 119.100 165.000 119.200 ;
        RECT 146.200 118.800 165.000 119.100 ;
        RECT 14.200 118.100 14.600 118.200 ;
        RECT 23.000 118.100 23.400 118.200 ;
        RECT 14.200 117.800 23.400 118.100 ;
        RECT 40.600 117.800 41.000 118.200 ;
        RECT 46.200 118.100 46.600 118.200 ;
        RECT 48.600 118.100 49.000 118.200 ;
        RECT 46.200 117.800 49.000 118.100 ;
        RECT 50.200 117.800 50.600 118.200 ;
        RECT 59.000 118.100 59.400 118.200 ;
        RECT 99.000 118.100 99.400 118.200 ;
        RECT 59.000 117.800 99.400 118.100 ;
        RECT 101.400 117.800 101.800 118.200 ;
        RECT 111.000 118.100 111.400 118.200 ;
        RECT 111.800 118.100 112.200 118.200 ;
        RECT 111.000 117.800 112.200 118.100 ;
        RECT 113.400 118.100 113.800 118.200 ;
        RECT 127.000 118.100 127.400 118.200 ;
        RECT 154.200 118.100 154.600 118.200 ;
        RECT 155.000 118.100 155.400 118.200 ;
        RECT 113.400 117.800 155.400 118.100 ;
        RECT 184.600 118.100 185.000 118.200 ;
        RECT 197.400 118.100 197.800 118.200 ;
        RECT 184.600 117.800 197.800 118.100 ;
        RECT 14.200 117.100 14.600 117.200 ;
        RECT 29.400 117.100 29.800 117.200 ;
        RECT 31.000 117.100 31.400 117.200 ;
        RECT 14.200 116.800 17.700 117.100 ;
        RECT 29.400 116.800 31.400 117.100 ;
        RECT 37.400 117.100 37.800 117.200 ;
        RECT 40.600 117.100 40.900 117.800 ;
        RECT 37.400 116.800 40.900 117.100 ;
        RECT 50.200 117.200 50.500 117.800 ;
        RECT 101.400 117.200 101.700 117.800 ;
        RECT 50.200 116.800 50.600 117.200 ;
        RECT 59.000 117.100 59.400 117.200 ;
        RECT 61.400 117.100 61.800 117.200 ;
        RECT 74.200 117.100 74.600 117.200 ;
        RECT 59.000 116.800 61.800 117.100 ;
        RECT 71.800 116.800 74.600 117.100 ;
        RECT 101.400 116.800 101.800 117.200 ;
        RECT 103.800 117.100 104.200 117.200 ;
        RECT 109.400 117.100 109.800 117.200 ;
        RECT 103.800 116.800 109.800 117.100 ;
        RECT 111.800 117.100 112.200 117.200 ;
        RECT 112.600 117.100 113.000 117.200 ;
        RECT 111.800 116.800 113.000 117.100 ;
        RECT 115.800 117.100 116.200 117.200 ;
        RECT 119.000 117.100 119.400 117.200 ;
        RECT 123.000 117.100 123.400 117.200 ;
        RECT 115.800 116.800 123.400 117.100 ;
        RECT 125.400 116.800 125.800 117.200 ;
        RECT 137.400 117.100 137.800 117.200 ;
        RECT 144.600 117.100 145.000 117.200 ;
        RECT 137.400 116.800 145.000 117.100 ;
        RECT 155.800 116.800 156.200 117.200 ;
        RECT 188.600 117.100 189.000 117.200 ;
        RECT 163.800 116.800 189.000 117.100 ;
        RECT 192.600 117.100 193.000 117.200 ;
        RECT 201.400 117.100 201.800 117.200 ;
        RECT 228.600 117.100 229.000 117.200 ;
        RECT 192.600 116.800 229.000 117.100 ;
        RECT 17.400 116.200 17.700 116.800 ;
        RECT 71.800 116.200 72.100 116.800 ;
        RECT 125.400 116.200 125.700 116.800 ;
        RECT 155.800 116.200 156.100 116.800 ;
        RECT 163.800 116.200 164.100 116.800 ;
        RECT 7.800 115.800 8.200 116.200 ;
        RECT 17.400 116.100 17.800 116.200 ;
        RECT 20.600 116.100 21.000 116.200 ;
        RECT 17.400 115.800 21.000 116.100 ;
        RECT 27.000 116.100 27.400 116.200 ;
        RECT 35.800 116.100 36.200 116.200 ;
        RECT 51.000 116.100 51.400 116.200 ;
        RECT 27.000 115.800 51.400 116.100 ;
        RECT 71.800 115.800 72.200 116.200 ;
        RECT 79.000 115.800 79.400 116.200 ;
        RECT 79.800 116.100 80.200 116.200 ;
        RECT 83.000 116.100 83.400 116.200 ;
        RECT 92.600 116.100 93.000 116.200 ;
        RECT 79.800 115.800 93.000 116.100 ;
        RECT 102.200 115.800 102.600 116.200 ;
        RECT 104.600 115.800 105.000 116.200 ;
        RECT 105.400 116.100 105.800 116.200 ;
        RECT 108.600 116.100 109.000 116.200 ;
        RECT 119.800 116.100 120.200 116.200 ;
        RECT 105.400 115.800 120.200 116.100 ;
        RECT 125.400 115.800 125.800 116.200 ;
        RECT 127.800 115.800 128.200 116.200 ;
        RECT 143.800 116.100 144.200 116.200 ;
        RECT 146.200 116.100 146.600 116.200 ;
        RECT 143.800 115.800 146.600 116.100 ;
        RECT 151.800 116.100 152.200 116.200 ;
        RECT 152.600 116.100 153.000 116.200 ;
        RECT 151.800 115.800 153.000 116.100 ;
        RECT 155.800 115.800 156.200 116.200 ;
        RECT 159.800 116.100 160.200 116.200 ;
        RECT 160.600 116.100 161.000 116.200 ;
        RECT 159.800 115.800 161.000 116.100 ;
        RECT 163.800 115.800 164.200 116.200 ;
        RECT 167.000 116.100 167.400 116.200 ;
        RECT 175.000 116.100 175.400 116.200 ;
        RECT 166.200 115.800 175.400 116.100 ;
        RECT 175.800 115.800 176.200 116.200 ;
        RECT 183.000 115.800 183.400 116.200 ;
        RECT 195.800 115.800 196.200 116.200 ;
        RECT 210.200 116.100 210.600 116.200 ;
        RECT 211.000 116.100 211.400 116.200 ;
        RECT 210.200 115.800 211.400 116.100 ;
        RECT 216.600 115.800 217.000 116.200 ;
        RECT 7.800 115.100 8.100 115.800 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 7.800 114.800 17.000 115.100 ;
        RECT 25.400 115.100 25.800 115.200 ;
        RECT 27.800 115.100 28.200 115.200 ;
        RECT 28.600 115.100 29.000 115.200 ;
        RECT 25.400 114.800 29.000 115.100 ;
        RECT 41.400 115.100 41.800 115.200 ;
        RECT 47.000 115.100 47.400 115.200 ;
        RECT 56.600 115.100 57.000 115.200 ;
        RECT 41.400 114.800 47.400 115.100 ;
        RECT 50.200 114.800 57.000 115.100 ;
        RECT 64.600 115.100 65.000 115.200 ;
        RECT 65.400 115.100 65.800 115.200 ;
        RECT 64.600 114.800 65.800 115.100 ;
        RECT 68.600 115.100 69.000 115.200 ;
        RECT 69.400 115.100 69.800 115.200 ;
        RECT 68.600 114.800 69.800 115.100 ;
        RECT 78.200 115.100 78.600 115.200 ;
        RECT 79.000 115.100 79.300 115.800 ;
        RECT 102.200 115.200 102.500 115.800 ;
        RECT 104.600 115.200 104.900 115.800 ;
        RECT 127.800 115.200 128.100 115.800 ;
        RECT 163.800 115.200 164.100 115.800 ;
        RECT 175.800 115.200 176.100 115.800 ;
        RECT 183.000 115.200 183.300 115.800 ;
        RECT 96.600 115.100 97.000 115.200 ;
        RECT 78.200 114.800 79.300 115.100 ;
        RECT 88.600 114.800 97.000 115.100 ;
        RECT 102.200 114.800 102.600 115.200 ;
        RECT 103.000 115.100 103.400 115.200 ;
        RECT 103.800 115.100 104.200 115.200 ;
        RECT 103.000 114.800 104.200 115.100 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 105.400 115.100 105.800 115.200 ;
        RECT 114.200 115.100 114.600 115.200 ;
        RECT 105.400 114.800 114.600 115.100 ;
        RECT 117.400 115.100 117.800 115.200 ;
        RECT 121.400 115.100 121.800 115.200 ;
        RECT 117.400 114.800 121.800 115.100 ;
        RECT 127.800 114.800 128.200 115.200 ;
        RECT 131.000 115.100 131.400 115.200 ;
        RECT 142.200 115.100 142.600 115.200 ;
        RECT 147.800 115.100 148.200 115.200 ;
        RECT 131.000 114.800 148.200 115.100 ;
        RECT 149.400 115.100 149.800 115.200 ;
        RECT 151.000 115.100 151.400 115.200 ;
        RECT 151.800 115.100 152.200 115.200 ;
        RECT 149.400 114.800 152.200 115.100 ;
        RECT 159.000 114.800 159.400 115.200 ;
        RECT 163.800 114.800 164.200 115.200 ;
        RECT 165.400 115.100 165.800 115.200 ;
        RECT 166.200 115.100 166.600 115.200 ;
        RECT 165.400 114.800 166.600 115.100 ;
        RECT 175.800 114.800 176.200 115.200 ;
        RECT 183.000 114.800 183.400 115.200 ;
        RECT 184.600 115.100 185.000 115.200 ;
        RECT 186.200 115.100 186.600 115.200 ;
        RECT 184.600 114.800 186.600 115.100 ;
        RECT 187.800 115.100 188.200 115.200 ;
        RECT 195.800 115.100 196.100 115.800 ;
        RECT 216.600 115.200 216.900 115.800 ;
        RECT 187.800 114.800 196.100 115.100 ;
        RECT 205.400 115.100 205.800 115.200 ;
        RECT 207.800 115.100 208.200 115.200 ;
        RECT 210.200 115.100 210.600 115.200 ;
        RECT 205.400 114.800 210.600 115.100 ;
        RECT 216.600 114.800 217.000 115.200 ;
        RECT 50.200 114.200 50.500 114.800 ;
        RECT 88.600 114.700 89.000 114.800 ;
        RECT 15.000 113.800 15.400 114.200 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 19.000 114.100 19.400 114.200 ;
        RECT 17.400 113.800 19.400 114.100 ;
        RECT 23.000 114.100 23.400 114.200 ;
        RECT 27.000 114.100 27.400 114.200 ;
        RECT 30.200 114.100 30.600 114.200 ;
        RECT 23.000 113.800 30.600 114.100 ;
        RECT 32.600 113.800 33.000 114.200 ;
        RECT 35.000 113.800 35.400 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 46.200 114.100 46.600 114.200 ;
        RECT 40.600 113.800 46.600 114.100 ;
        RECT 50.200 113.800 50.600 114.200 ;
        RECT 62.200 113.800 68.900 114.100 ;
        RECT 15.000 113.200 15.300 113.800 ;
        RECT 15.000 112.800 15.400 113.200 ;
        RECT 19.800 113.100 20.200 113.200 ;
        RECT 26.200 113.100 26.600 113.200 ;
        RECT 32.600 113.100 32.900 113.800 ;
        RECT 19.800 112.800 32.900 113.100 ;
        RECT 35.000 113.200 35.300 113.800 ;
        RECT 62.200 113.200 62.500 113.800 ;
        RECT 68.600 113.200 68.900 113.800 ;
        RECT 78.200 113.800 78.600 114.200 ;
        RECT 79.000 114.100 79.400 114.200 ;
        RECT 103.800 114.100 104.200 114.200 ;
        RECT 79.000 113.800 104.200 114.100 ;
        RECT 118.200 114.100 118.600 114.200 ;
        RECT 121.400 114.100 121.800 114.200 ;
        RECT 123.000 114.100 123.400 114.200 ;
        RECT 118.200 113.800 123.400 114.100 ;
        RECT 141.400 114.100 141.800 114.200 ;
        RECT 148.600 114.100 149.000 114.200 ;
        RECT 150.200 114.100 150.600 114.200 ;
        RECT 141.400 113.800 150.600 114.100 ;
        RECT 155.800 114.100 156.200 114.200 ;
        RECT 159.000 114.100 159.300 114.800 ;
        RECT 155.800 113.800 159.300 114.100 ;
        RECT 163.800 114.100 164.200 114.200 ;
        RECT 167.000 114.100 167.400 114.200 ;
        RECT 175.000 114.100 175.400 114.200 ;
        RECT 185.400 114.100 185.800 114.200 ;
        RECT 163.800 113.800 174.500 114.100 ;
        RECT 175.000 113.800 185.800 114.100 ;
        RECT 204.600 114.100 205.000 114.200 ;
        RECT 208.600 114.100 209.000 114.200 ;
        RECT 204.600 113.800 209.000 114.100 ;
        RECT 219.000 114.100 219.400 114.200 ;
        RECT 223.000 114.100 223.400 114.200 ;
        RECT 219.000 113.800 223.400 114.100 ;
        RECT 78.200 113.200 78.500 113.800 ;
        RECT 35.000 112.800 35.400 113.200 ;
        RECT 62.200 112.800 62.600 113.200 ;
        RECT 63.800 113.100 64.200 113.200 ;
        RECT 64.600 113.100 65.000 113.200 ;
        RECT 63.800 112.800 65.000 113.100 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 68.600 112.800 69.000 113.200 ;
        RECT 76.600 113.100 77.000 113.200 ;
        RECT 77.400 113.100 77.800 113.200 ;
        RECT 76.600 112.800 77.800 113.100 ;
        RECT 78.200 112.800 78.600 113.200 ;
        RECT 95.800 113.100 96.200 113.200 ;
        RECT 98.200 113.100 98.600 113.200 ;
        RECT 106.200 113.100 106.600 113.200 ;
        RECT 95.800 112.800 106.600 113.100 ;
        RECT 109.400 113.100 109.800 113.200 ;
        RECT 110.200 113.100 110.600 113.200 ;
        RECT 112.600 113.100 113.000 113.200 ;
        RECT 109.400 112.800 113.000 113.100 ;
        RECT 116.600 113.100 117.000 113.200 ;
        RECT 119.800 113.100 120.200 113.200 ;
        RECT 116.600 112.800 120.200 113.100 ;
        RECT 139.000 113.100 139.400 113.200 ;
        RECT 142.200 113.100 142.600 113.200 ;
        RECT 139.000 112.800 142.600 113.100 ;
        RECT 148.600 113.100 149.000 113.200 ;
        RECT 157.400 113.100 157.800 113.200 ;
        RECT 148.600 112.800 157.800 113.100 ;
        RECT 174.200 113.100 174.500 113.800 ;
        RECT 176.600 113.100 177.000 113.200 ;
        RECT 179.800 113.100 180.200 113.200 ;
        RECT 174.200 112.800 180.200 113.100 ;
        RECT 22.200 112.100 22.600 112.200 ;
        RECT 25.400 112.100 25.800 112.200 ;
        RECT 21.400 111.800 25.800 112.100 ;
        RECT 43.000 111.800 43.400 112.200 ;
        RECT 48.600 112.100 49.000 112.200 ;
        RECT 53.400 112.100 53.800 112.200 ;
        RECT 57.400 112.100 57.800 112.200 ;
        RECT 48.600 111.800 57.800 112.100 ;
        RECT 64.600 112.100 65.000 112.200 ;
        RECT 67.000 112.100 67.300 112.800 ;
        RECT 74.200 112.100 74.600 112.200 ;
        RECT 77.400 112.100 77.800 112.200 ;
        RECT 80.600 112.100 81.000 112.200 ;
        RECT 64.600 111.800 81.000 112.100 ;
        RECT 100.600 112.100 101.000 112.200 ;
        RECT 114.200 112.100 114.600 112.200 ;
        RECT 100.600 111.800 114.600 112.100 ;
        RECT 115.000 112.100 115.400 112.200 ;
        RECT 119.000 112.100 119.400 112.200 ;
        RECT 115.000 111.800 119.400 112.100 ;
        RECT 119.800 112.100 120.100 112.800 ;
        RECT 148.600 112.100 149.000 112.200 ;
        RECT 119.800 111.800 149.000 112.100 ;
        RECT 155.000 112.100 155.400 112.200 ;
        RECT 167.800 112.100 168.200 112.200 ;
        RECT 155.000 111.800 168.200 112.100 ;
        RECT 178.200 112.100 178.600 112.200 ;
        RECT 183.800 112.100 184.200 112.200 ;
        RECT 178.200 111.800 184.200 112.100 ;
        RECT 191.800 112.100 192.200 112.200 ;
        RECT 204.600 112.100 205.000 112.200 ;
        RECT 191.800 111.800 205.000 112.100 ;
        RECT 227.800 111.800 228.200 112.200 ;
        RECT 43.000 111.200 43.300 111.800 ;
        RECT 227.800 111.200 228.100 111.800 ;
        RECT 43.000 110.800 43.400 111.200 ;
        RECT 47.800 111.100 48.200 111.200 ;
        RECT 69.400 111.100 69.800 111.200 ;
        RECT 47.800 110.800 69.800 111.100 ;
        RECT 73.400 111.100 73.800 111.200 ;
        RECT 74.200 111.100 74.600 111.200 ;
        RECT 73.400 110.800 74.600 111.100 ;
        RECT 99.000 111.100 99.400 111.200 ;
        RECT 149.400 111.100 149.800 111.200 ;
        RECT 151.800 111.100 152.200 111.200 ;
        RECT 99.000 110.800 137.700 111.100 ;
        RECT 149.400 110.800 152.200 111.100 ;
        RECT 154.200 111.100 154.600 111.200 ;
        RECT 179.000 111.100 179.400 111.200 ;
        RECT 154.200 110.800 179.400 111.100 ;
        RECT 180.600 111.100 181.000 111.200 ;
        RECT 183.800 111.100 184.200 111.200 ;
        RECT 180.600 110.800 184.200 111.100 ;
        RECT 227.800 110.800 228.200 111.200 ;
        RECT 137.400 110.200 137.700 110.800 ;
        RECT 29.400 110.100 29.800 110.200 ;
        RECT 51.800 110.100 52.200 110.200 ;
        RECT 29.400 109.800 52.200 110.100 ;
        RECT 56.600 109.800 57.000 110.200 ;
        RECT 60.600 110.100 61.000 110.200 ;
        RECT 65.400 110.100 65.800 110.200 ;
        RECT 60.600 109.800 65.800 110.100 ;
        RECT 103.800 110.100 104.200 110.200 ;
        RECT 105.400 110.100 105.800 110.200 ;
        RECT 103.800 109.800 105.800 110.100 ;
        RECT 106.200 110.100 106.600 110.200 ;
        RECT 118.200 110.100 118.600 110.200 ;
        RECT 119.000 110.100 119.400 110.200 ;
        RECT 106.200 109.800 119.400 110.100 ;
        RECT 129.400 110.100 129.800 110.200 ;
        RECT 135.000 110.100 135.400 110.200 ;
        RECT 129.400 109.800 135.400 110.100 ;
        RECT 137.400 110.100 137.800 110.200 ;
        RECT 147.000 110.100 147.400 110.200 ;
        RECT 150.200 110.100 150.600 110.200 ;
        RECT 171.000 110.100 171.400 110.200 ;
        RECT 186.200 110.100 186.600 110.200 ;
        RECT 137.400 109.800 186.600 110.100 ;
        RECT 203.800 110.100 204.200 110.200 ;
        RECT 222.200 110.100 222.600 110.200 ;
        RECT 228.600 110.100 229.000 110.200 ;
        RECT 203.800 109.800 229.000 110.100 ;
        RECT 0.600 109.100 1.000 109.200 ;
        RECT 3.000 109.100 3.400 109.200 ;
        RECT 0.600 108.800 3.400 109.100 ;
        RECT 23.000 109.100 23.400 109.200 ;
        RECT 26.200 109.100 26.600 109.200 ;
        RECT 23.000 108.800 26.600 109.100 ;
        RECT 56.600 109.100 56.900 109.800 ;
        RECT 59.000 109.100 59.400 109.200 ;
        RECT 56.600 108.800 59.400 109.100 ;
        RECT 98.200 109.100 98.600 109.200 ;
        RECT 103.000 109.100 103.400 109.200 ;
        RECT 109.400 109.100 109.800 109.200 ;
        RECT 98.200 108.800 109.800 109.100 ;
        RECT 114.200 109.100 114.600 109.200 ;
        RECT 124.600 109.100 125.000 109.200 ;
        RECT 114.200 108.800 125.000 109.100 ;
        RECT 126.200 109.100 126.600 109.200 ;
        RECT 128.600 109.100 129.000 109.200 ;
        RECT 126.200 108.800 129.000 109.100 ;
        RECT 141.400 109.100 141.800 109.200 ;
        RECT 151.800 109.100 152.200 109.200 ;
        RECT 141.400 108.800 152.200 109.100 ;
        RECT 158.200 109.100 158.600 109.200 ;
        RECT 167.800 109.100 168.200 109.200 ;
        RECT 158.200 108.800 168.200 109.100 ;
        RECT 207.000 109.100 207.400 109.200 ;
        RECT 207.800 109.100 208.200 109.200 ;
        RECT 207.000 108.800 208.200 109.100 ;
        RECT 1.400 108.100 1.800 108.200 ;
        RECT 2.200 108.100 2.600 108.200 ;
        RECT 8.600 108.100 9.000 108.200 ;
        RECT 15.800 108.100 16.200 108.200 ;
        RECT 19.800 108.100 20.200 108.200 ;
        RECT 31.000 108.100 31.400 108.200 ;
        RECT 1.400 107.800 3.300 108.100 ;
        RECT 8.600 107.800 20.200 108.100 ;
        RECT 24.600 107.800 31.400 108.100 ;
        RECT 85.400 108.100 85.800 108.200 ;
        RECT 99.000 108.100 99.400 108.200 ;
        RECT 85.400 107.800 99.400 108.100 ;
        RECT 106.200 108.100 106.600 108.200 ;
        RECT 128.600 108.100 129.000 108.200 ;
        RECT 106.200 107.800 129.000 108.100 ;
        RECT 131.000 108.100 131.400 108.200 ;
        RECT 139.000 108.100 139.400 108.200 ;
        RECT 131.000 107.800 139.400 108.100 ;
        RECT 148.600 108.100 149.000 108.200 ;
        RECT 162.200 108.100 162.600 108.200 ;
        RECT 176.600 108.100 177.000 108.200 ;
        RECT 148.600 107.800 177.000 108.100 ;
        RECT 180.600 107.800 181.000 108.200 ;
        RECT 228.600 108.100 229.000 108.200 ;
        RECT 229.400 108.100 229.800 108.200 ;
        RECT 228.600 107.800 229.800 108.100 ;
        RECT 3.000 107.100 3.400 107.200 ;
        RECT 3.800 107.100 4.200 107.200 ;
        RECT 8.600 107.100 9.000 107.200 ;
        RECT 3.000 106.800 4.200 107.100 ;
        RECT 7.800 106.800 9.000 107.100 ;
        RECT 15.000 106.800 15.400 107.200 ;
        RECT 19.000 107.100 19.400 107.200 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 24.600 107.100 24.900 107.800 ;
        RECT 19.000 106.800 24.900 107.100 ;
        RECT 25.400 106.800 25.800 107.200 ;
        RECT 40.600 107.100 41.000 107.200 ;
        RECT 48.600 107.100 49.000 107.200 ;
        RECT 40.600 106.800 49.000 107.100 ;
        RECT 52.600 107.100 53.000 107.200 ;
        RECT 60.600 107.100 61.000 107.200 ;
        RECT 52.600 106.800 61.000 107.100 ;
        RECT 73.400 107.100 73.800 107.200 ;
        RECT 78.200 107.100 78.600 107.200 ;
        RECT 81.400 107.100 81.800 107.200 ;
        RECT 73.400 106.800 81.800 107.100 ;
        RECT 94.200 107.100 94.600 107.200 ;
        RECT 106.200 107.100 106.500 107.800 ;
        RECT 180.600 107.200 180.900 107.800 ;
        RECT 94.200 106.800 106.500 107.100 ;
        RECT 117.400 107.100 117.800 107.200 ;
        RECT 121.400 107.100 121.800 107.200 ;
        RECT 123.000 107.100 123.400 107.200 ;
        RECT 117.400 106.800 123.400 107.100 ;
        RECT 126.200 107.100 126.600 107.200 ;
        RECT 135.800 107.100 136.200 107.200 ;
        RECT 126.200 106.800 136.200 107.100 ;
        RECT 149.400 107.100 149.800 107.200 ;
        RECT 156.600 107.100 157.000 107.200 ;
        RECT 158.200 107.100 158.600 107.200 ;
        RECT 149.400 106.800 158.600 107.100 ;
        RECT 159.000 107.100 159.400 107.200 ;
        RECT 159.800 107.100 160.200 107.200 ;
        RECT 163.800 107.100 164.200 107.200 ;
        RECT 159.000 106.800 164.200 107.100 ;
        RECT 166.200 107.100 166.600 107.200 ;
        RECT 167.000 107.100 167.400 107.200 ;
        RECT 166.200 106.800 167.400 107.100 ;
        RECT 167.800 107.100 168.200 107.200 ;
        RECT 178.200 107.100 178.600 107.200 ;
        RECT 167.800 106.800 178.600 107.100 ;
        RECT 179.800 106.800 180.200 107.200 ;
        RECT 180.600 106.800 181.000 107.200 ;
        RECT 181.400 107.100 181.800 107.200 ;
        RECT 187.000 107.100 187.400 107.200 ;
        RECT 181.400 106.800 187.400 107.100 ;
        RECT 189.400 107.100 189.800 107.200 ;
        RECT 197.400 107.100 197.800 107.200 ;
        RECT 189.400 106.800 197.800 107.100 ;
        RECT 207.000 107.100 207.400 107.200 ;
        RECT 207.800 107.100 208.200 107.200 ;
        RECT 207.000 106.800 208.200 107.100 ;
        RECT 4.600 106.100 5.000 106.200 ;
        RECT 7.800 106.100 8.100 106.800 ;
        RECT 4.600 105.800 8.100 106.100 ;
        RECT 15.000 106.100 15.300 106.800 ;
        RECT 25.400 106.200 25.700 106.800 ;
        RECT 179.800 106.200 180.100 106.800 ;
        RECT 22.200 106.100 22.600 106.200 ;
        RECT 15.000 105.800 22.600 106.100 ;
        RECT 25.400 105.800 25.800 106.200 ;
        RECT 31.800 106.100 32.200 106.200 ;
        RECT 36.600 106.100 37.000 106.200 ;
        RECT 43.800 106.100 44.200 106.200 ;
        RECT 31.800 105.800 44.200 106.100 ;
        RECT 67.000 106.100 67.400 106.200 ;
        RECT 83.800 106.100 84.200 106.200 ;
        RECT 67.000 105.800 84.200 106.100 ;
        RECT 94.200 106.100 94.600 106.200 ;
        RECT 98.200 106.100 98.600 106.200 ;
        RECT 94.200 105.800 98.600 106.100 ;
        RECT 99.800 106.100 100.200 106.200 ;
        RECT 122.200 106.100 122.600 106.200 ;
        RECT 99.800 105.800 101.700 106.100 ;
        RECT 101.400 105.200 101.700 105.800 ;
        RECT 120.600 105.800 122.600 106.100 ;
        RECT 145.400 106.100 145.800 106.200 ;
        RECT 147.000 106.100 147.400 106.200 ;
        RECT 145.400 105.800 147.400 106.100 ;
        RECT 155.000 106.100 155.400 106.200 ;
        RECT 156.600 106.100 157.000 106.200 ;
        RECT 155.000 105.800 157.000 106.100 ;
        RECT 157.400 106.100 157.800 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 157.400 105.800 158.600 106.100 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 164.600 106.100 165.000 106.200 ;
        RECT 163.000 105.800 165.000 106.100 ;
        RECT 179.800 106.100 180.200 106.200 ;
        RECT 181.400 106.100 181.800 106.200 ;
        RECT 179.800 105.800 181.800 106.100 ;
        RECT 183.000 105.800 183.400 106.200 ;
        RECT 188.600 106.100 189.000 106.200 ;
        RECT 189.400 106.100 189.800 106.200 ;
        RECT 188.600 105.800 189.800 106.100 ;
        RECT 210.200 106.100 210.600 106.200 ;
        RECT 214.200 106.100 214.600 106.200 ;
        RECT 210.200 105.800 214.600 106.100 ;
        RECT 120.600 105.200 120.900 105.800 ;
        RECT 183.000 105.200 183.300 105.800 ;
        RECT 7.800 105.100 8.200 105.200 ;
        RECT 19.800 105.100 20.200 105.200 ;
        RECT 7.800 104.800 20.200 105.100 ;
        RECT 20.600 105.100 21.000 105.200 ;
        RECT 23.000 105.100 23.400 105.200 ;
        RECT 20.600 104.800 23.400 105.100 ;
        RECT 61.400 105.100 61.800 105.200 ;
        RECT 63.000 105.100 63.400 105.200 ;
        RECT 61.400 104.800 63.400 105.100 ;
        RECT 73.400 105.100 73.800 105.200 ;
        RECT 91.800 105.100 92.200 105.200 ;
        RECT 99.800 105.100 100.200 105.200 ;
        RECT 73.400 104.800 83.300 105.100 ;
        RECT 91.800 104.800 100.200 105.100 ;
        RECT 101.400 105.100 101.800 105.200 ;
        RECT 102.200 105.100 102.600 105.200 ;
        RECT 101.400 104.800 102.600 105.100 ;
        RECT 120.600 104.800 121.000 105.200 ;
        RECT 135.800 105.100 136.200 105.200 ;
        RECT 126.200 104.800 136.200 105.100 ;
        RECT 137.400 105.100 137.800 105.200 ;
        RECT 141.400 105.100 141.800 105.200 ;
        RECT 137.400 104.800 141.800 105.100 ;
        RECT 145.400 105.100 145.800 105.200 ;
        RECT 146.200 105.100 146.600 105.200 ;
        RECT 145.400 104.800 146.600 105.100 ;
        RECT 152.600 105.100 153.000 105.200 ;
        RECT 153.400 105.100 153.800 105.200 ;
        RECT 152.600 104.800 153.800 105.100 ;
        RECT 157.400 104.800 157.800 105.200 ;
        RECT 163.800 105.100 164.200 105.200 ;
        RECT 172.600 105.100 173.000 105.200 ;
        RECT 163.800 104.800 173.000 105.100 ;
        RECT 174.200 105.100 174.600 105.200 ;
        RECT 180.600 105.100 181.000 105.200 ;
        RECT 174.200 104.800 181.000 105.100 ;
        RECT 183.000 104.800 183.400 105.200 ;
        RECT 186.200 104.800 186.600 105.200 ;
        RECT 187.000 105.100 187.400 105.200 ;
        RECT 190.200 105.100 190.600 105.200 ;
        RECT 187.000 104.800 190.600 105.100 ;
        RECT 207.800 105.100 208.200 105.200 ;
        RECT 211.000 105.100 211.400 105.200 ;
        RECT 207.800 104.800 211.400 105.100 ;
        RECT 23.000 104.200 23.300 104.800 ;
        RECT 83.000 104.200 83.300 104.800 ;
        RECT 126.200 104.200 126.500 104.800 ;
        RECT 157.400 104.200 157.700 104.800 ;
        RECT 186.200 104.200 186.500 104.800 ;
        RECT 0.600 104.100 1.000 104.200 ;
        RECT 19.000 104.100 19.400 104.200 ;
        RECT 0.600 103.800 19.400 104.100 ;
        RECT 23.000 103.800 23.400 104.200 ;
        RECT 27.800 104.100 28.200 104.200 ;
        RECT 50.200 104.100 50.600 104.200 ;
        RECT 27.800 103.800 50.600 104.100 ;
        RECT 60.600 104.100 61.000 104.200 ;
        RECT 75.800 104.100 76.200 104.200 ;
        RECT 60.600 103.800 76.200 104.100 ;
        RECT 83.000 103.800 83.400 104.200 ;
        RECT 115.800 104.100 116.200 104.200 ;
        RECT 120.600 104.100 121.000 104.200 ;
        RECT 115.800 103.800 121.000 104.100 ;
        RECT 126.200 103.800 126.600 104.200 ;
        RECT 137.400 104.100 137.800 104.200 ;
        RECT 143.800 104.100 144.200 104.200 ;
        RECT 137.400 103.800 144.200 104.100 ;
        RECT 157.400 103.800 157.800 104.200 ;
        RECT 159.000 104.100 159.400 104.200 ;
        RECT 159.800 104.100 160.200 104.200 ;
        RECT 159.000 103.800 160.200 104.100 ;
        RECT 186.200 103.800 186.600 104.200 ;
        RECT 11.800 103.100 12.200 103.200 ;
        RECT 14.200 103.100 14.600 103.200 ;
        RECT 43.800 103.100 44.200 103.200 ;
        RECT 68.600 103.100 69.000 103.200 ;
        RECT 11.800 102.800 69.000 103.100 ;
        RECT 83.000 103.100 83.300 103.800 ;
        RECT 94.200 103.100 94.600 103.200 ;
        RECT 83.000 102.800 94.600 103.100 ;
        RECT 135.800 103.100 136.200 103.200 ;
        RECT 144.600 103.100 145.000 103.200 ;
        RECT 135.800 102.800 145.000 103.100 ;
        RECT 151.800 103.100 152.200 103.200 ;
        RECT 163.000 103.100 163.400 103.200 ;
        RECT 151.800 102.800 163.400 103.100 ;
        RECT 9.400 102.100 9.800 102.200 ;
        RECT 19.800 102.100 20.200 102.200 ;
        RECT 21.400 102.100 21.800 102.200 ;
        RECT 47.000 102.100 47.400 102.200 ;
        RECT 63.800 102.100 64.200 102.200 ;
        RECT 9.400 101.800 21.800 102.100 ;
        RECT 46.200 101.800 64.200 102.100 ;
        RECT 68.600 102.100 69.000 102.200 ;
        RECT 76.600 102.100 77.000 102.200 ;
        RECT 86.200 102.100 86.600 102.200 ;
        RECT 68.600 101.800 86.600 102.100 ;
        RECT 95.000 102.100 95.400 102.200 ;
        RECT 99.800 102.100 100.200 102.200 ;
        RECT 95.000 101.800 100.200 102.100 ;
        RECT 100.600 102.100 101.000 102.200 ;
        RECT 116.600 102.100 117.000 102.200 ;
        RECT 121.400 102.100 121.800 102.200 ;
        RECT 160.600 102.100 161.000 102.200 ;
        RECT 100.600 101.800 161.000 102.100 ;
        RECT 6.200 101.100 6.600 101.200 ;
        RECT 17.400 101.100 17.800 101.200 ;
        RECT 34.200 101.100 34.600 101.200 ;
        RECT 6.200 100.800 34.600 101.100 ;
        RECT 39.800 101.100 40.200 101.200 ;
        RECT 63.800 101.100 64.200 101.200 ;
        RECT 74.200 101.100 74.600 101.200 ;
        RECT 39.800 100.800 74.600 101.100 ;
        RECT 75.000 101.100 75.400 101.200 ;
        RECT 95.000 101.100 95.400 101.200 ;
        RECT 75.000 100.800 95.400 101.100 ;
        RECT 100.600 101.100 101.000 101.200 ;
        RECT 107.000 101.100 107.400 101.200 ;
        RECT 100.600 100.800 107.400 101.100 ;
        RECT 111.800 101.100 112.200 101.200 ;
        RECT 120.600 101.100 121.000 101.200 ;
        RECT 111.800 100.800 121.000 101.100 ;
        RECT 127.000 101.100 127.400 101.200 ;
        RECT 129.400 101.100 129.800 101.200 ;
        RECT 127.000 100.800 129.800 101.100 ;
        RECT 149.400 101.100 149.800 101.200 ;
        RECT 151.000 101.100 151.400 101.200 ;
        RECT 149.400 100.800 151.400 101.100 ;
        RECT 173.400 101.100 173.800 101.200 ;
        RECT 207.000 101.100 207.400 101.200 ;
        RECT 226.200 101.100 226.600 101.200 ;
        RECT 173.400 100.800 226.600 101.100 ;
        RECT 43.800 100.100 44.200 100.200 ;
        RECT 52.600 100.100 53.000 100.200 ;
        RECT 43.800 99.800 53.000 100.100 ;
        RECT 75.800 100.100 76.200 100.200 ;
        RECT 97.400 100.100 97.800 100.200 ;
        RECT 107.800 100.100 108.200 100.200 ;
        RECT 113.400 100.100 113.800 100.200 ;
        RECT 75.800 99.800 113.800 100.100 ;
        RECT 28.600 99.100 29.000 99.200 ;
        RECT 43.800 99.100 44.200 99.200 ;
        RECT 28.600 98.800 44.200 99.100 ;
        RECT 77.400 99.100 77.800 99.200 ;
        RECT 90.200 99.100 90.600 99.200 ;
        RECT 94.200 99.100 94.600 99.200 ;
        RECT 77.400 98.800 94.600 99.100 ;
        RECT 95.000 99.100 95.400 99.200 ;
        RECT 102.200 99.100 102.600 99.200 ;
        RECT 95.000 98.800 102.600 99.100 ;
        RECT 104.600 99.100 105.000 99.200 ;
        RECT 111.800 99.100 112.200 99.200 ;
        RECT 104.600 98.800 112.200 99.100 ;
        RECT 113.400 99.100 113.800 99.200 ;
        RECT 127.000 99.100 127.400 99.200 ;
        RECT 148.600 99.100 149.000 99.200 ;
        RECT 113.400 98.800 149.000 99.100 ;
        RECT 151.000 99.100 151.400 99.200 ;
        RECT 185.400 99.100 185.800 99.200 ;
        RECT 190.200 99.100 190.600 99.200 ;
        RECT 151.000 98.800 190.600 99.100 ;
        RECT 33.400 98.100 33.800 98.200 ;
        RECT 44.600 98.100 45.000 98.200 ;
        RECT 33.400 97.800 45.000 98.100 ;
        RECT 69.400 98.100 69.800 98.200 ;
        RECT 71.800 98.100 72.200 98.200 ;
        RECT 95.800 98.100 96.200 98.200 ;
        RECT 69.400 97.800 96.200 98.100 ;
        RECT 101.400 98.100 101.800 98.200 ;
        RECT 107.800 98.100 108.200 98.200 ;
        RECT 101.400 97.800 108.200 98.100 ;
        RECT 108.600 98.100 109.000 98.200 ;
        RECT 114.200 98.100 114.600 98.200 ;
        RECT 115.800 98.100 116.200 98.200 ;
        RECT 108.600 97.800 116.200 98.100 ;
        RECT 118.200 98.100 118.600 98.200 ;
        RECT 119.000 98.100 119.400 98.200 ;
        RECT 123.000 98.100 123.400 98.200 ;
        RECT 118.200 97.800 123.400 98.100 ;
        RECT 142.200 98.100 142.600 98.200 ;
        RECT 143.800 98.100 144.200 98.200 ;
        RECT 148.600 98.100 149.000 98.200 ;
        RECT 166.200 98.100 166.600 98.200 ;
        RECT 175.800 98.100 176.200 98.200 ;
        RECT 201.400 98.100 201.800 98.200 ;
        RECT 142.200 97.800 201.800 98.100 ;
        RECT 20.600 97.100 21.000 97.200 ;
        RECT 29.400 97.100 29.800 97.200 ;
        RECT 20.600 96.800 29.800 97.100 ;
        RECT 33.400 97.100 33.800 97.200 ;
        RECT 40.600 97.100 41.000 97.200 ;
        RECT 33.400 96.800 41.000 97.100 ;
        RECT 51.000 97.100 51.400 97.200 ;
        RECT 51.800 97.100 52.200 97.200 ;
        RECT 51.000 96.800 52.200 97.100 ;
        RECT 54.200 97.100 54.600 97.200 ;
        RECT 57.400 97.100 57.800 97.200 ;
        RECT 54.200 96.800 57.800 97.100 ;
        RECT 63.800 97.100 64.200 97.200 ;
        RECT 72.600 97.100 73.000 97.200 ;
        RECT 77.400 97.100 77.800 97.200 ;
        RECT 63.800 96.800 77.800 97.100 ;
        RECT 83.800 97.100 84.200 97.200 ;
        RECT 91.000 97.100 91.400 97.200 ;
        RECT 83.800 96.800 91.400 97.100 ;
        RECT 92.600 97.100 93.000 97.200 ;
        RECT 93.400 97.100 93.800 97.200 ;
        RECT 92.600 96.800 93.800 97.100 ;
        RECT 95.000 97.100 95.400 97.200 ;
        RECT 100.600 97.100 101.000 97.200 ;
        RECT 95.000 96.800 101.000 97.100 ;
        RECT 104.600 96.800 105.000 97.200 ;
        RECT 114.200 96.800 114.600 97.200 ;
        RECT 122.200 97.100 122.600 97.200 ;
        RECT 147.800 97.100 148.200 97.200 ;
        RECT 155.000 97.100 155.400 97.200 ;
        RECT 122.200 96.800 145.700 97.100 ;
        RECT 147.800 96.800 155.400 97.100 ;
        RECT 174.200 97.100 174.600 97.200 ;
        RECT 181.400 97.100 181.800 97.200 ;
        RECT 174.200 96.800 181.800 97.100 ;
        RECT 198.200 97.100 198.600 97.200 ;
        RECT 213.400 97.100 213.800 97.200 ;
        RECT 227.000 97.100 227.400 97.200 ;
        RECT 198.200 96.800 227.400 97.100 ;
        RECT 104.600 96.200 104.900 96.800 ;
        RECT 1.400 96.100 1.800 96.200 ;
        RECT 10.200 96.100 10.600 96.200 ;
        RECT 1.400 95.800 10.600 96.100 ;
        RECT 12.600 96.100 13.000 96.200 ;
        RECT 14.200 96.100 14.600 96.200 ;
        RECT 12.600 95.800 14.600 96.100 ;
        RECT 16.600 96.100 17.000 96.200 ;
        RECT 19.000 96.100 19.400 96.200 ;
        RECT 16.600 95.800 19.400 96.100 ;
        RECT 31.000 96.100 31.400 96.200 ;
        RECT 35.000 96.100 35.400 96.200 ;
        RECT 63.000 96.100 63.400 96.200 ;
        RECT 80.600 96.100 81.000 96.200 ;
        RECT 85.400 96.100 85.800 96.200 ;
        RECT 31.000 95.800 81.000 96.100 ;
        RECT 82.200 95.800 85.800 96.100 ;
        RECT 95.000 96.100 95.400 96.200 ;
        RECT 95.000 95.800 96.900 96.100 ;
        RECT 104.600 95.800 105.000 96.200 ;
        RECT 106.200 96.100 106.600 96.200 ;
        RECT 114.200 96.100 114.500 96.800 ;
        RECT 106.200 95.800 114.500 96.100 ;
        RECT 115.800 96.100 116.200 96.200 ;
        RECT 124.600 96.100 125.000 96.200 ;
        RECT 115.800 95.800 125.000 96.100 ;
        RECT 128.600 96.100 129.000 96.200 ;
        RECT 132.600 96.100 133.000 96.200 ;
        RECT 128.600 95.800 133.000 96.100 ;
        RECT 142.200 96.100 142.600 96.200 ;
        RECT 144.600 96.100 145.000 96.200 ;
        RECT 142.200 95.800 145.000 96.100 ;
        RECT 145.400 96.100 145.700 96.800 ;
        RECT 156.600 96.100 157.000 96.200 ;
        RECT 145.400 95.800 157.000 96.100 ;
        RECT 168.600 96.100 169.000 96.200 ;
        RECT 191.800 96.100 192.200 96.200 ;
        RECT 168.600 95.800 192.200 96.100 ;
        RECT 196.600 96.100 197.000 96.200 ;
        RECT 202.200 96.100 202.600 96.200 ;
        RECT 203.000 96.100 203.400 96.200 ;
        RECT 196.600 95.800 203.400 96.100 ;
        RECT 203.800 96.100 204.200 96.200 ;
        RECT 223.800 96.100 224.200 96.200 ;
        RECT 203.800 95.800 224.200 96.100 ;
        RECT 6.200 95.100 6.600 95.200 ;
        RECT 12.600 95.100 13.000 95.200 ;
        RECT 6.200 94.800 13.000 95.100 ;
        RECT 14.200 95.100 14.600 95.200 ;
        RECT 15.000 95.100 15.400 95.200 ;
        RECT 14.200 94.800 15.400 95.100 ;
        RECT 19.000 95.100 19.400 95.200 ;
        RECT 19.000 94.800 25.000 95.100 ;
        RECT 24.600 94.700 25.000 94.800 ;
        RECT 47.000 94.800 47.400 95.200 ;
        RECT 54.200 94.800 54.600 95.200 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 69.400 95.100 69.800 95.200 ;
        RECT 62.200 94.800 69.800 95.100 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 82.200 95.100 82.500 95.800 ;
        RECT 96.600 95.200 96.900 95.800 ;
        RECT 78.200 94.800 82.500 95.100 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 89.400 95.100 89.800 95.200 ;
        RECT 83.000 94.800 89.800 95.100 ;
        RECT 91.000 95.100 91.400 95.200 ;
        RECT 92.600 95.100 93.000 95.200 ;
        RECT 91.000 94.800 93.000 95.100 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 98.200 95.100 98.600 95.200 ;
        RECT 99.000 95.100 99.400 95.200 ;
        RECT 124.600 95.100 125.000 95.200 ;
        RECT 127.800 95.100 128.200 95.200 ;
        RECT 138.200 95.100 138.600 95.200 ;
        RECT 98.200 94.800 99.400 95.100 ;
        RECT 102.200 94.800 138.600 95.100 ;
        RECT 143.000 95.100 143.400 95.200 ;
        RECT 147.000 95.100 147.400 95.200 ;
        RECT 143.000 94.800 147.400 95.100 ;
        RECT 151.800 95.100 152.200 95.200 ;
        RECT 152.600 95.100 153.000 95.200 ;
        RECT 151.800 94.800 153.000 95.100 ;
        RECT 171.800 95.100 172.200 95.200 ;
        RECT 180.600 95.100 181.000 95.200 ;
        RECT 183.000 95.100 183.400 95.200 ;
        RECT 185.400 95.100 185.800 95.200 ;
        RECT 171.800 94.800 185.800 95.100 ;
        RECT 187.000 95.100 187.400 95.200 ;
        RECT 187.800 95.100 188.200 95.200 ;
        RECT 194.200 95.100 194.600 95.200 ;
        RECT 187.000 94.800 194.600 95.100 ;
        RECT 195.000 95.100 195.400 95.200 ;
        RECT 197.400 95.100 197.800 95.200 ;
        RECT 195.000 94.800 197.800 95.100 ;
        RECT 199.800 95.100 200.200 95.200 ;
        RECT 204.600 95.100 205.000 95.200 ;
        RECT 199.800 94.800 205.000 95.100 ;
        RECT 206.200 95.100 206.600 95.200 ;
        RECT 206.200 94.800 209.000 95.100 ;
        RECT 11.000 94.100 11.400 94.200 ;
        RECT 24.600 94.100 25.000 94.200 ;
        RECT 8.600 93.800 25.000 94.100 ;
        RECT 30.200 94.100 30.600 94.200 ;
        RECT 31.800 94.100 32.200 94.200 ;
        RECT 30.200 93.800 32.200 94.100 ;
        RECT 41.400 94.100 41.800 94.200 ;
        RECT 47.000 94.100 47.300 94.800 ;
        RECT 54.200 94.200 54.500 94.800 ;
        RECT 41.400 93.800 47.300 94.100 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 54.200 94.100 54.600 94.200 ;
        RECT 48.600 93.800 54.600 94.100 ;
        RECT 57.400 93.800 57.800 94.200 ;
        RECT 80.600 94.100 81.000 94.200 ;
        RECT 102.200 94.100 102.500 94.800 ;
        RECT 208.600 94.700 209.000 94.800 ;
        RECT 210.200 94.800 217.700 95.100 ;
        RECT 80.600 93.800 102.500 94.100 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 109.400 94.100 109.800 94.200 ;
        RECT 103.000 93.800 109.800 94.100 ;
        RECT 113.400 94.100 113.800 94.200 ;
        RECT 119.800 94.100 120.200 94.200 ;
        RECT 121.400 94.100 121.800 94.200 ;
        RECT 154.200 94.100 154.600 94.200 ;
        RECT 113.400 93.800 154.600 94.100 ;
        RECT 179.000 94.100 179.400 94.200 ;
        RECT 185.400 94.100 185.800 94.200 ;
        RECT 187.000 94.100 187.400 94.200 ;
        RECT 179.000 93.800 187.400 94.100 ;
        RECT 199.800 94.100 200.200 94.200 ;
        RECT 200.600 94.100 201.000 94.200 ;
        RECT 199.800 93.800 201.000 94.100 ;
        RECT 202.200 94.100 202.600 94.200 ;
        RECT 210.200 94.100 210.500 94.800 ;
        RECT 217.400 94.200 217.700 94.800 ;
        RECT 202.200 93.800 210.500 94.100 ;
        RECT 211.000 94.100 211.400 94.200 ;
        RECT 211.000 93.800 216.100 94.100 ;
        RECT 217.400 93.800 217.800 94.200 ;
        RECT 8.600 93.200 8.900 93.800 ;
        RECT 8.600 92.800 9.000 93.200 ;
        RECT 14.200 93.100 14.600 93.200 ;
        RECT 15.000 93.100 15.400 93.200 ;
        RECT 32.600 93.100 33.000 93.200 ;
        RECT 55.000 93.100 55.400 93.200 ;
        RECT 14.200 92.800 15.400 93.100 ;
        RECT 31.800 92.800 55.400 93.100 ;
        RECT 57.400 93.100 57.700 93.800 ;
        RECT 215.800 93.200 216.100 93.800 ;
        RECT 62.200 93.100 62.600 93.200 ;
        RECT 57.400 92.800 62.600 93.100 ;
        RECT 63.800 93.100 64.200 93.200 ;
        RECT 69.400 93.100 69.800 93.200 ;
        RECT 63.800 92.800 69.800 93.100 ;
        RECT 75.800 93.100 76.200 93.200 ;
        RECT 95.800 93.100 96.200 93.200 ;
        RECT 98.200 93.100 98.600 93.200 ;
        RECT 75.800 92.800 98.600 93.100 ;
        RECT 107.800 93.100 108.200 93.200 ;
        RECT 112.600 93.100 113.000 93.200 ;
        RECT 107.800 92.800 113.000 93.100 ;
        RECT 120.600 92.800 121.000 93.200 ;
        RECT 125.400 93.100 125.800 93.200 ;
        RECT 126.200 93.100 126.600 93.200 ;
        RECT 125.400 92.800 126.600 93.100 ;
        RECT 129.400 93.100 129.800 93.200 ;
        RECT 132.600 93.100 133.000 93.200 ;
        RECT 204.600 93.100 205.000 93.200 ;
        RECT 129.400 92.800 205.000 93.100 ;
        RECT 215.800 92.800 216.200 93.200 ;
        RECT 26.200 92.100 26.600 92.200 ;
        RECT 40.600 92.100 41.000 92.200 ;
        RECT 26.200 91.800 41.000 92.100 ;
        RECT 49.400 92.100 49.800 92.200 ;
        RECT 55.000 92.100 55.400 92.200 ;
        RECT 101.400 92.100 101.800 92.200 ;
        RECT 49.400 91.800 101.800 92.100 ;
        RECT 103.800 92.100 104.200 92.200 ;
        RECT 108.600 92.100 109.000 92.200 ;
        RECT 115.800 92.100 116.200 92.200 ;
        RECT 120.600 92.100 120.900 92.800 ;
        RECT 103.800 91.800 120.900 92.100 ;
        RECT 130.200 92.100 130.600 92.200 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 130.200 91.800 132.200 92.100 ;
        RECT 135.800 92.100 136.200 92.200 ;
        RECT 136.600 92.100 137.000 92.200 ;
        RECT 135.800 91.800 137.000 92.100 ;
        RECT 160.600 92.100 161.000 92.200 ;
        RECT 163.000 92.100 163.400 92.200 ;
        RECT 160.600 91.800 163.400 92.100 ;
        RECT 183.000 92.100 183.400 92.200 ;
        RECT 191.800 92.100 192.200 92.200 ;
        RECT 183.000 91.800 192.200 92.100 ;
        RECT 11.800 91.100 12.200 91.200 ;
        RECT 12.600 91.100 13.000 91.200 ;
        RECT 11.800 90.800 13.000 91.100 ;
        RECT 30.200 91.100 30.600 91.200 ;
        RECT 46.200 91.100 46.600 91.200 ;
        RECT 30.200 90.800 46.600 91.100 ;
        RECT 51.800 91.100 52.200 91.200 ;
        RECT 75.800 91.100 76.200 91.200 ;
        RECT 51.800 90.800 76.200 91.100 ;
        RECT 77.400 91.100 77.800 91.200 ;
        RECT 79.800 91.100 80.200 91.200 ;
        RECT 77.400 90.800 80.200 91.100 ;
        RECT 99.800 91.100 100.200 91.200 ;
        RECT 100.600 91.100 101.000 91.200 ;
        RECT 99.800 90.800 101.000 91.100 ;
        RECT 151.800 91.100 152.200 91.200 ;
        RECT 155.000 91.100 155.400 91.200 ;
        RECT 151.800 90.800 155.400 91.100 ;
        RECT 163.000 91.100 163.400 91.200 ;
        RECT 165.400 91.100 165.800 91.200 ;
        RECT 163.000 90.800 165.800 91.100 ;
        RECT 167.000 91.100 167.400 91.200 ;
        RECT 169.400 91.100 169.800 91.200 ;
        RECT 167.000 90.800 169.800 91.100 ;
        RECT 13.400 90.100 13.800 90.200 ;
        RECT 31.000 90.100 31.400 90.200 ;
        RECT 13.400 89.800 31.400 90.100 ;
        RECT 42.200 90.100 42.600 90.200 ;
        RECT 43.800 90.100 44.200 90.200 ;
        RECT 60.600 90.100 61.000 90.200 ;
        RECT 42.200 89.800 61.000 90.100 ;
        RECT 109.400 90.100 109.800 90.200 ;
        RECT 117.400 90.100 117.800 90.200 ;
        RECT 109.400 89.800 117.800 90.100 ;
        RECT 147.800 90.100 148.200 90.200 ;
        RECT 149.400 90.100 149.800 90.200 ;
        RECT 147.800 89.800 149.800 90.100 ;
        RECT 154.200 90.100 154.600 90.200 ;
        RECT 179.800 90.100 180.200 90.200 ;
        RECT 154.200 89.800 180.200 90.100 ;
        RECT 183.800 90.100 184.200 90.200 ;
        RECT 184.600 90.100 185.000 90.200 ;
        RECT 183.800 89.800 185.000 90.100 ;
        RECT 189.400 90.100 189.800 90.200 ;
        RECT 190.200 90.100 190.600 90.200 ;
        RECT 189.400 89.800 190.600 90.100 ;
        RECT 208.600 90.100 209.000 90.200 ;
        RECT 227.800 90.100 228.200 90.200 ;
        RECT 208.600 89.800 228.200 90.100 ;
        RECT 11.800 89.100 12.200 89.200 ;
        RECT 16.600 89.100 17.000 89.200 ;
        RECT 11.800 88.800 17.000 89.100 ;
        RECT 17.400 89.100 17.800 89.200 ;
        RECT 28.600 89.100 29.000 89.200 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 41.400 89.100 41.800 89.200 ;
        RECT 17.400 88.800 27.300 89.100 ;
        RECT 28.600 88.800 41.800 89.100 ;
        RECT 43.000 89.100 43.400 89.200 ;
        RECT 43.800 89.100 44.200 89.200 ;
        RECT 43.000 88.800 44.200 89.100 ;
        RECT 52.600 89.100 53.000 89.200 ;
        RECT 57.400 89.100 57.800 89.200 ;
        RECT 52.600 88.800 57.800 89.100 ;
        RECT 63.000 89.100 63.400 89.200 ;
        RECT 68.600 89.100 69.000 89.200 ;
        RECT 63.000 88.800 69.000 89.100 ;
        RECT 79.800 89.100 80.200 89.200 ;
        RECT 83.000 89.100 83.400 89.200 ;
        RECT 79.800 88.800 83.400 89.100 ;
        RECT 89.400 89.100 89.800 89.200 ;
        RECT 93.400 89.100 93.800 89.200 ;
        RECT 89.400 88.800 93.800 89.100 ;
        RECT 114.200 88.800 114.600 89.200 ;
        RECT 117.400 89.100 117.800 89.200 ;
        RECT 118.200 89.100 118.600 89.200 ;
        RECT 121.400 89.100 121.800 89.200 ;
        RECT 124.600 89.100 125.000 89.200 ;
        RECT 117.400 88.800 118.600 89.100 ;
        RECT 120.600 88.800 125.000 89.100 ;
        RECT 125.400 89.100 125.800 89.200 ;
        RECT 129.400 89.100 129.800 89.200 ;
        RECT 125.400 88.800 129.800 89.100 ;
        RECT 131.800 89.100 132.200 89.200 ;
        RECT 140.600 89.100 141.000 89.200 ;
        RECT 131.800 88.800 141.000 89.100 ;
        RECT 147.000 89.100 147.400 89.200 ;
        RECT 149.400 89.100 149.800 89.200 ;
        RECT 147.000 88.800 149.800 89.100 ;
        RECT 152.600 89.100 153.000 89.200 ;
        RECT 153.400 89.100 153.800 89.200 ;
        RECT 152.600 88.800 153.800 89.100 ;
        RECT 161.400 89.100 161.800 89.200 ;
        RECT 166.200 89.100 166.600 89.200 ;
        RECT 161.400 88.800 166.600 89.100 ;
        RECT 176.600 88.800 177.000 89.200 ;
        RECT 179.800 89.100 180.100 89.800 ;
        RECT 183.000 89.100 183.400 89.200 ;
        RECT 192.600 89.100 193.000 89.200 ;
        RECT 202.200 89.100 202.600 89.200 ;
        RECT 179.800 88.800 202.600 89.100 ;
        RECT 219.000 89.100 219.400 89.200 ;
        RECT 223.800 89.100 224.200 89.200 ;
        RECT 219.000 88.800 224.200 89.100 ;
        RECT 27.000 88.200 27.300 88.800 ;
        RECT 9.400 88.100 9.800 88.200 ;
        RECT 13.400 88.100 13.800 88.200 ;
        RECT 9.400 87.800 13.800 88.100 ;
        RECT 16.600 88.100 17.000 88.200 ;
        RECT 26.200 88.100 26.600 88.200 ;
        RECT 16.600 87.800 26.600 88.100 ;
        RECT 27.000 88.100 27.400 88.200 ;
        RECT 39.800 88.100 40.200 88.200 ;
        RECT 27.000 87.800 40.200 88.100 ;
        RECT 42.200 88.100 42.600 88.200 ;
        RECT 51.800 88.100 52.200 88.200 ;
        RECT 42.200 87.800 52.200 88.100 ;
        RECT 53.400 88.100 53.800 88.200 ;
        RECT 55.800 88.100 56.200 88.200 ;
        RECT 53.400 87.800 56.200 88.100 ;
        RECT 56.600 88.100 57.000 88.200 ;
        RECT 63.000 88.100 63.400 88.200 ;
        RECT 78.200 88.100 78.600 88.200 ;
        RECT 56.600 87.800 78.600 88.100 ;
        RECT 83.000 88.100 83.400 88.200 ;
        RECT 94.200 88.100 94.600 88.200 ;
        RECT 95.000 88.100 95.400 88.200 ;
        RECT 83.000 87.800 95.400 88.100 ;
        RECT 98.200 88.100 98.600 88.200 ;
        RECT 104.600 88.100 105.000 88.200 ;
        RECT 98.200 87.800 105.000 88.100 ;
        RECT 114.200 88.100 114.500 88.800 ;
        RECT 176.600 88.200 176.900 88.800 ;
        RECT 116.600 88.100 117.000 88.200 ;
        RECT 114.200 87.800 117.000 88.100 ;
        RECT 120.600 88.100 121.000 88.200 ;
        RECT 123.800 88.100 124.200 88.200 ;
        RECT 120.600 87.800 124.200 88.100 ;
        RECT 135.000 88.100 135.400 88.200 ;
        RECT 147.000 88.100 147.400 88.200 ;
        RECT 154.200 88.100 154.600 88.200 ;
        RECT 135.000 87.800 154.600 88.100 ;
        RECT 165.400 88.100 165.800 88.200 ;
        RECT 169.400 88.100 169.800 88.200 ;
        RECT 165.400 87.800 169.800 88.100 ;
        RECT 176.600 87.800 177.000 88.200 ;
        RECT 179.000 88.100 179.400 88.200 ;
        RECT 183.800 88.100 184.200 88.200 ;
        RECT 179.000 87.800 184.200 88.100 ;
        RECT 189.400 88.100 189.800 88.200 ;
        RECT 197.400 88.100 197.800 88.200 ;
        RECT 189.400 87.800 197.800 88.100 ;
        RECT 222.200 87.800 222.600 88.200 ;
        RECT 26.200 87.200 26.500 87.800 ;
        RECT 12.600 87.100 13.000 87.200 ;
        RECT 21.400 87.100 21.800 87.200 ;
        RECT 12.600 86.800 21.800 87.100 ;
        RECT 26.200 86.800 26.600 87.200 ;
        RECT 64.600 87.100 65.000 87.200 ;
        RECT 65.400 87.100 65.800 87.200 ;
        RECT 64.600 86.800 65.800 87.100 ;
        RECT 67.800 87.100 68.200 87.200 ;
        RECT 89.400 87.100 89.800 87.200 ;
        RECT 67.800 86.800 89.800 87.100 ;
        RECT 90.200 87.100 90.600 87.200 ;
        RECT 95.000 87.100 95.400 87.200 ;
        RECT 90.200 86.800 95.400 87.100 ;
        RECT 98.200 87.100 98.600 87.200 ;
        RECT 101.400 87.100 101.800 87.200 ;
        RECT 98.200 86.800 101.800 87.100 ;
        RECT 104.600 87.100 105.000 87.200 ;
        RECT 126.200 87.100 126.600 87.200 ;
        RECT 134.200 87.100 134.600 87.200 ;
        RECT 104.600 86.800 134.600 87.100 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 144.600 87.100 145.000 87.200 ;
        RECT 137.400 86.800 145.000 87.100 ;
        RECT 152.600 87.100 153.000 87.200 ;
        RECT 155.800 87.100 156.200 87.200 ;
        RECT 152.600 86.800 156.200 87.100 ;
        RECT 156.600 87.100 157.000 87.200 ;
        RECT 157.400 87.100 157.800 87.200 ;
        RECT 156.600 86.800 157.800 87.100 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 168.600 87.100 169.000 87.200 ;
        RECT 171.800 87.100 172.200 87.200 ;
        RECT 174.200 87.100 174.600 87.200 ;
        RECT 199.000 87.100 199.400 87.200 ;
        RECT 168.600 86.800 199.400 87.100 ;
        RECT 213.400 87.100 213.800 87.200 ;
        RECT 222.200 87.100 222.500 87.800 ;
        RECT 213.400 86.800 222.500 87.100 ;
        RECT 5.400 86.100 5.800 86.200 ;
        RECT 11.000 86.100 11.400 86.200 ;
        RECT 5.400 85.800 11.400 86.100 ;
        RECT 17.400 86.100 17.800 86.200 ;
        RECT 20.600 86.100 21.000 86.200 ;
        RECT 17.400 85.800 21.000 86.100 ;
        RECT 26.200 86.100 26.600 86.200 ;
        RECT 32.600 86.100 33.000 86.300 ;
        RECT 26.200 85.900 33.000 86.100 ;
        RECT 47.000 86.100 47.400 86.200 ;
        RECT 63.000 86.100 63.400 86.200 ;
        RECT 63.800 86.100 64.200 86.200 ;
        RECT 26.200 85.800 32.900 85.900 ;
        RECT 47.000 85.800 54.500 86.100 ;
        RECT 63.000 85.800 64.200 86.100 ;
        RECT 67.000 86.100 67.400 86.200 ;
        RECT 73.400 86.100 73.800 86.200 ;
        RECT 83.000 86.100 83.400 86.200 ;
        RECT 67.000 85.800 73.800 86.100 ;
        RECT 76.600 85.800 83.400 86.100 ;
        RECT 90.200 86.100 90.600 86.200 ;
        RECT 91.000 86.100 91.400 86.200 ;
        RECT 90.200 85.800 91.400 86.100 ;
        RECT 97.400 86.100 97.800 86.200 ;
        RECT 104.600 86.100 105.000 86.200 ;
        RECT 110.200 86.100 110.600 86.200 ;
        RECT 97.400 85.800 110.600 86.100 ;
        RECT 111.000 86.100 111.400 86.200 ;
        RECT 143.800 86.100 144.200 86.200 ;
        RECT 145.400 86.100 145.800 86.200 ;
        RECT 178.200 86.100 178.600 86.200 ;
        RECT 111.000 85.800 178.600 86.100 ;
        RECT 179.000 86.100 179.400 86.200 ;
        RECT 180.600 86.100 181.000 86.200 ;
        RECT 179.000 85.800 181.000 86.100 ;
        RECT 183.800 85.800 184.200 86.200 ;
        RECT 195.800 86.100 196.200 86.200 ;
        RECT 203.000 86.100 203.400 86.200 ;
        RECT 195.800 85.800 203.400 86.100 ;
        RECT 207.800 85.800 208.200 86.200 ;
        RECT 223.800 86.100 224.200 86.200 ;
        RECT 225.400 86.100 225.800 86.200 ;
        RECT 223.800 85.800 225.800 86.100 ;
        RECT 54.200 85.200 54.500 85.800 ;
        RECT 76.600 85.200 76.900 85.800 ;
        RECT 11.000 85.100 11.400 85.200 ;
        RECT 14.200 85.100 14.600 85.200 ;
        RECT 11.000 84.800 14.600 85.100 ;
        RECT 15.800 85.100 16.200 85.200 ;
        RECT 23.800 85.100 24.200 85.200 ;
        RECT 15.800 84.800 24.200 85.100 ;
        RECT 26.200 85.100 26.600 85.200 ;
        RECT 39.000 85.100 39.400 85.200 ;
        RECT 41.400 85.100 41.800 85.200 ;
        RECT 26.200 84.800 27.300 85.100 ;
        RECT 39.000 84.800 41.800 85.100 ;
        RECT 54.200 84.800 54.600 85.200 ;
        RECT 76.600 84.800 77.000 85.200 ;
        RECT 85.400 85.100 85.800 85.200 ;
        RECT 91.800 85.100 92.200 85.200 ;
        RECT 85.400 84.800 92.200 85.100 ;
        RECT 95.000 85.100 95.400 85.200 ;
        RECT 95.800 85.100 96.200 85.200 ;
        RECT 95.000 84.800 96.200 85.100 ;
        RECT 97.400 85.100 97.800 85.200 ;
        RECT 98.200 85.100 98.600 85.200 ;
        RECT 97.400 84.800 98.600 85.100 ;
        RECT 116.600 85.100 117.000 85.200 ;
        RECT 152.600 85.100 153.000 85.200 ;
        RECT 116.600 84.800 153.000 85.100 ;
        RECT 153.400 84.800 153.800 85.200 ;
        RECT 154.200 85.100 154.600 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 154.200 84.800 162.600 85.100 ;
        RECT 163.800 85.100 164.200 85.200 ;
        RECT 166.200 85.100 166.600 85.200 ;
        RECT 168.600 85.100 169.000 85.200 ;
        RECT 163.800 84.800 169.000 85.100 ;
        RECT 175.000 85.100 175.400 85.200 ;
        RECT 179.800 85.100 180.200 85.200 ;
        RECT 175.000 84.800 180.200 85.100 ;
        RECT 182.200 85.100 182.600 85.200 ;
        RECT 183.800 85.100 184.100 85.800 ;
        RECT 207.800 85.200 208.100 85.800 ;
        RECT 182.200 84.800 184.100 85.100 ;
        RECT 186.200 85.100 186.600 85.200 ;
        RECT 187.000 85.100 187.400 85.200 ;
        RECT 186.200 84.800 187.400 85.100 ;
        RECT 193.400 85.100 193.800 85.200 ;
        RECT 195.800 85.100 196.200 85.200 ;
        RECT 193.400 84.800 196.200 85.100 ;
        RECT 207.800 84.800 208.200 85.200 ;
        RECT 219.000 85.100 219.400 85.200 ;
        RECT 223.000 85.100 223.400 85.200 ;
        RECT 227.000 85.100 227.400 85.200 ;
        RECT 219.000 84.800 227.400 85.100 ;
        RECT 27.000 84.200 27.300 84.800 ;
        RECT 153.400 84.200 153.700 84.800 ;
        RECT 195.800 84.200 196.100 84.800 ;
        RECT 10.200 84.100 10.600 84.200 ;
        RECT 15.000 84.100 15.400 84.200 ;
        RECT 10.200 83.800 15.400 84.100 ;
        RECT 27.000 83.800 27.400 84.200 ;
        RECT 27.800 84.100 28.200 84.200 ;
        RECT 47.800 84.100 48.200 84.200 ;
        RECT 27.800 83.800 48.200 84.100 ;
        RECT 56.600 84.100 57.000 84.200 ;
        RECT 59.800 84.100 60.200 84.200 ;
        RECT 56.600 83.800 60.200 84.100 ;
        RECT 94.200 84.100 94.600 84.200 ;
        RECT 112.600 84.100 113.000 84.200 ;
        RECT 94.200 83.800 113.000 84.100 ;
        RECT 153.400 83.800 153.800 84.200 ;
        RECT 159.800 84.100 160.200 84.200 ;
        RECT 163.800 84.100 164.200 84.200 ;
        RECT 159.800 83.800 164.200 84.100 ;
        RECT 167.000 84.100 167.400 84.200 ;
        RECT 171.800 84.100 172.200 84.200 ;
        RECT 167.000 83.800 172.200 84.100 ;
        RECT 176.600 84.100 177.000 84.200 ;
        RECT 180.600 84.100 181.000 84.200 ;
        RECT 186.200 84.100 186.600 84.200 ;
        RECT 176.600 83.800 186.600 84.100 ;
        RECT 195.800 83.800 196.200 84.200 ;
        RECT 220.600 84.100 221.000 84.200 ;
        RECT 227.000 84.100 227.400 84.200 ;
        RECT 220.600 83.800 227.400 84.100 ;
        RECT 24.600 83.100 25.000 83.200 ;
        RECT 27.000 83.100 27.400 83.200 ;
        RECT 30.200 83.100 30.600 83.200 ;
        RECT 43.800 83.100 44.200 83.200 ;
        RECT 24.600 82.800 44.200 83.100 ;
        RECT 185.400 83.100 185.800 83.200 ;
        RECT 193.400 83.100 193.800 83.200 ;
        RECT 185.400 82.800 193.800 83.100 ;
        RECT 42.200 82.100 42.600 82.200 ;
        RECT 44.600 82.100 45.000 82.200 ;
        RECT 42.200 81.800 45.000 82.100 ;
        RECT 61.400 82.100 61.800 82.200 ;
        RECT 63.800 82.100 64.200 82.200 ;
        RECT 61.400 81.800 64.200 82.100 ;
        RECT 178.200 82.100 178.600 82.200 ;
        RECT 187.800 82.100 188.200 82.200 ;
        RECT 178.200 81.800 188.200 82.100 ;
        RECT 103.000 81.100 103.400 81.200 ;
        RECT 113.400 81.100 113.800 81.200 ;
        RECT 103.000 80.800 113.800 81.100 ;
        RECT 163.800 81.100 164.200 81.200 ;
        RECT 183.000 81.100 183.400 81.200 ;
        RECT 163.800 80.800 183.400 81.100 ;
        RECT 179.800 80.100 180.200 80.200 ;
        RECT 217.400 80.100 217.800 80.200 ;
        RECT 219.800 80.100 220.200 80.200 ;
        RECT 179.800 79.800 220.200 80.100 ;
        RECT 20.600 79.100 21.000 79.200 ;
        RECT 31.000 79.100 31.400 79.200 ;
        RECT 35.000 79.100 35.400 79.200 ;
        RECT 20.600 78.800 35.400 79.100 ;
        RECT 46.200 79.100 46.600 79.200 ;
        RECT 50.200 79.100 50.600 79.200 ;
        RECT 66.200 79.100 66.600 79.200 ;
        RECT 46.200 78.800 66.600 79.100 ;
        RECT 98.200 79.100 98.600 79.200 ;
        RECT 99.800 79.100 100.200 79.200 ;
        RECT 109.400 79.100 109.800 79.200 ;
        RECT 98.200 78.800 109.800 79.100 ;
        RECT 127.000 79.100 127.400 79.200 ;
        RECT 144.600 79.100 145.000 79.200 ;
        RECT 127.000 78.800 145.000 79.100 ;
        RECT 199.800 79.100 200.200 79.200 ;
        RECT 209.400 79.100 209.800 79.200 ;
        RECT 199.800 78.800 209.800 79.100 ;
        RECT 11.000 77.800 11.400 78.200 ;
        RECT 19.000 78.100 19.400 78.200 ;
        RECT 35.800 78.100 36.200 78.200 ;
        RECT 19.000 77.800 36.200 78.100 ;
        RECT 49.400 78.100 49.800 78.200 ;
        RECT 59.800 78.100 60.200 78.200 ;
        RECT 49.400 77.800 60.200 78.100 ;
        RECT 72.600 78.100 73.000 78.200 ;
        RECT 107.000 78.100 107.400 78.200 ;
        RECT 143.000 78.100 143.400 78.200 ;
        RECT 145.400 78.100 145.800 78.200 ;
        RECT 203.800 78.100 204.200 78.200 ;
        RECT 223.800 78.100 224.200 78.200 ;
        RECT 72.600 77.800 224.200 78.100 ;
        RECT 4.600 77.100 5.000 77.200 ;
        RECT 11.000 77.100 11.300 77.800 ;
        RECT 4.600 76.800 11.300 77.100 ;
        RECT 14.200 77.100 14.600 77.200 ;
        RECT 16.600 77.100 17.000 77.200 ;
        RECT 19.000 77.100 19.400 77.200 ;
        RECT 14.200 76.800 19.400 77.100 ;
        RECT 21.400 77.100 21.800 77.200 ;
        RECT 25.400 77.100 25.800 77.200 ;
        RECT 21.400 76.800 25.800 77.100 ;
        RECT 51.000 77.100 51.400 77.200 ;
        RECT 61.400 77.100 61.800 77.200 ;
        RECT 51.000 76.800 61.800 77.100 ;
        RECT 82.200 77.100 82.600 77.200 ;
        RECT 93.400 77.100 93.800 77.200 ;
        RECT 82.200 76.800 93.800 77.100 ;
        RECT 118.200 77.100 118.600 77.200 ;
        RECT 137.400 77.100 137.800 77.200 ;
        RECT 147.800 77.100 148.200 77.200 ;
        RECT 118.200 76.800 148.200 77.100 ;
        RECT 148.600 76.800 149.000 77.200 ;
        RECT 179.000 77.100 179.400 77.200 ;
        RECT 179.800 77.100 180.200 77.200 ;
        RECT 179.000 76.800 180.200 77.100 ;
        RECT 184.600 77.100 185.000 77.200 ;
        RECT 187.800 77.100 188.200 77.200 ;
        RECT 184.600 76.800 188.200 77.100 ;
        RECT 190.200 77.100 190.600 77.200 ;
        RECT 191.800 77.100 192.200 77.200 ;
        RECT 190.200 76.800 192.200 77.100 ;
        RECT 195.800 77.100 196.200 77.200 ;
        RECT 207.000 77.100 207.400 77.200 ;
        RECT 215.800 77.100 216.200 77.200 ;
        RECT 195.800 76.800 216.200 77.100 ;
        RECT 148.600 76.200 148.900 76.800 ;
        RECT 9.400 76.100 9.800 76.200 ;
        RECT 15.000 76.100 15.400 76.200 ;
        RECT 36.600 76.100 37.000 76.200 ;
        RECT 9.400 75.800 37.000 76.100 ;
        RECT 42.200 75.800 42.600 76.200 ;
        RECT 43.000 76.100 43.400 76.200 ;
        RECT 50.200 76.100 50.600 76.200 ;
        RECT 51.000 76.100 51.400 76.200 ;
        RECT 43.000 75.800 51.400 76.100 ;
        RECT 54.200 76.100 54.600 76.200 ;
        RECT 57.400 76.100 57.800 76.200 ;
        RECT 54.200 75.800 57.800 76.100 ;
        RECT 60.600 76.100 61.000 76.200 ;
        RECT 66.200 76.100 66.600 76.200 ;
        RECT 60.600 75.800 66.600 76.100 ;
        RECT 74.200 76.100 74.600 76.200 ;
        RECT 82.200 76.100 82.600 76.200 ;
        RECT 74.200 75.800 82.600 76.100 ;
        RECT 83.800 76.100 84.200 76.200 ;
        RECT 85.400 76.100 85.800 76.200 ;
        RECT 83.800 75.800 85.800 76.100 ;
        RECT 103.000 76.100 103.400 76.200 ;
        RECT 110.200 76.100 110.600 76.200 ;
        RECT 103.000 75.800 110.600 76.100 ;
        RECT 120.600 76.100 121.000 76.200 ;
        RECT 121.400 76.100 121.800 76.200 ;
        RECT 120.600 75.800 121.800 76.100 ;
        RECT 130.200 76.100 130.600 76.200 ;
        RECT 136.600 76.100 137.000 76.200 ;
        RECT 130.200 75.800 137.000 76.100 ;
        RECT 143.800 75.800 144.200 76.200 ;
        RECT 148.600 75.800 149.000 76.200 ;
        RECT 151.000 76.100 151.400 76.200 ;
        RECT 172.600 76.100 173.000 76.200 ;
        RECT 151.000 75.800 173.000 76.100 ;
        RECT 181.400 76.100 181.800 76.200 ;
        RECT 183.000 76.100 183.400 76.200 ;
        RECT 181.400 75.800 183.400 76.100 ;
        RECT 186.200 76.100 186.600 76.200 ;
        RECT 200.600 76.100 201.000 76.200 ;
        RECT 201.400 76.100 201.800 76.200 ;
        RECT 186.200 75.800 201.800 76.100 ;
        RECT 202.200 76.100 202.600 76.200 ;
        RECT 211.800 76.100 212.200 76.200 ;
        RECT 202.200 75.800 212.200 76.100 ;
        RECT 212.600 75.800 213.000 76.200 ;
        RECT 42.200 75.200 42.500 75.800 ;
        RECT 18.200 75.100 18.600 75.200 ;
        RECT 24.600 75.100 25.000 75.200 ;
        RECT 18.200 74.800 25.000 75.100 ;
        RECT 26.200 75.100 26.600 75.200 ;
        RECT 31.000 75.100 31.400 75.200 ;
        RECT 26.200 74.800 31.400 75.100 ;
        RECT 34.200 75.100 34.600 75.200 ;
        RECT 42.200 75.100 42.600 75.200 ;
        RECT 34.200 74.800 42.600 75.100 ;
        RECT 43.000 75.100 43.400 75.200 ;
        RECT 43.800 75.100 44.200 75.200 ;
        RECT 43.000 74.800 44.200 75.100 ;
        RECT 59.800 75.100 60.200 75.200 ;
        RECT 62.200 75.100 62.600 75.200 ;
        RECT 59.800 74.800 62.600 75.100 ;
        RECT 66.200 75.100 66.500 75.800 ;
        RECT 68.600 75.100 69.000 75.200 ;
        RECT 66.200 74.800 69.000 75.100 ;
        RECT 69.400 75.100 69.800 75.200 ;
        RECT 74.200 75.100 74.500 75.800 ;
        RECT 69.400 74.800 74.500 75.100 ;
        RECT 86.200 75.100 86.600 75.200 ;
        RECT 95.000 75.100 95.400 75.200 ;
        RECT 86.200 74.800 95.400 75.100 ;
        RECT 99.000 75.100 99.400 75.200 ;
        RECT 103.800 75.100 104.200 75.200 ;
        RECT 107.800 75.100 108.200 75.200 ;
        RECT 99.000 74.800 100.900 75.100 ;
        RECT 103.800 74.800 108.200 75.100 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 115.000 75.100 115.400 75.200 ;
        RECT 114.200 74.800 115.400 75.100 ;
        RECT 119.800 75.100 120.200 75.200 ;
        RECT 123.800 75.100 124.200 75.200 ;
        RECT 126.200 75.100 126.600 75.200 ;
        RECT 119.800 74.800 126.600 75.100 ;
        RECT 135.000 75.100 135.400 75.200 ;
        RECT 138.200 75.100 138.600 75.200 ;
        RECT 143.000 75.100 143.400 75.200 ;
        RECT 135.000 74.800 143.400 75.100 ;
        RECT 143.800 75.100 144.100 75.800 ;
        RECT 151.000 75.100 151.400 75.200 ;
        RECT 143.800 74.800 151.400 75.100 ;
        RECT 151.800 75.100 152.200 75.200 ;
        RECT 173.400 75.100 173.800 75.200 ;
        RECT 151.800 74.800 173.800 75.100 ;
        RECT 182.200 75.100 182.600 75.200 ;
        RECT 183.800 75.100 184.200 75.200 ;
        RECT 182.200 74.800 184.200 75.100 ;
        RECT 186.200 75.100 186.600 75.200 ;
        RECT 187.000 75.100 187.400 75.200 ;
        RECT 186.200 74.800 187.400 75.100 ;
        RECT 187.800 75.100 188.200 75.200 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 187.800 74.800 197.800 75.100 ;
        RECT 202.200 75.100 202.500 75.800 ;
        RECT 203.000 75.100 203.400 75.200 ;
        RECT 202.200 74.800 203.400 75.100 ;
        RECT 204.600 75.100 205.000 75.200 ;
        RECT 205.400 75.100 205.800 75.200 ;
        RECT 204.600 74.800 205.800 75.100 ;
        RECT 212.600 75.100 212.900 75.800 ;
        RECT 217.400 75.100 217.800 75.200 ;
        RECT 212.600 74.800 217.800 75.100 ;
        RECT 100.600 74.200 100.900 74.800 ;
        RECT 111.800 74.200 112.100 74.800 ;
        RECT 29.400 74.100 29.800 74.200 ;
        RECT 30.200 74.100 30.600 74.200 ;
        RECT 38.200 74.100 38.600 74.200 ;
        RECT 42.200 74.100 42.600 74.200 ;
        RECT 44.600 74.100 45.000 74.200 ;
        RECT 29.400 73.800 38.600 74.100 ;
        RECT 41.400 73.800 45.000 74.100 ;
        RECT 48.600 74.100 49.000 74.200 ;
        RECT 49.400 74.100 49.800 74.200 ;
        RECT 48.600 73.800 49.800 74.100 ;
        RECT 61.400 74.100 61.800 74.200 ;
        RECT 63.800 74.100 64.200 74.200 ;
        RECT 61.400 73.800 64.200 74.100 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 65.400 73.800 66.600 74.100 ;
        RECT 68.600 74.100 69.000 74.200 ;
        RECT 75.000 74.100 75.400 74.200 ;
        RECT 68.600 73.800 75.400 74.100 ;
        RECT 75.800 74.100 76.200 74.200 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 80.600 74.100 81.000 74.200 ;
        RECT 75.800 73.800 81.000 74.100 ;
        RECT 100.600 73.800 101.000 74.200 ;
        RECT 105.400 74.100 105.800 74.200 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 105.400 73.800 109.000 74.100 ;
        RECT 109.400 73.800 109.800 74.200 ;
        RECT 111.800 73.800 112.200 74.200 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 119.000 73.800 120.200 74.100 ;
        RECT 122.200 74.100 122.600 74.200 ;
        RECT 123.000 74.100 123.400 74.200 ;
        RECT 134.200 74.100 134.600 74.200 ;
        RECT 141.400 74.100 141.800 74.200 ;
        RECT 153.400 74.100 153.800 74.200 ;
        RECT 122.200 73.800 141.800 74.100 ;
        RECT 147.000 73.800 153.800 74.100 ;
        RECT 155.800 74.100 156.200 74.200 ;
        RECT 159.800 74.100 160.200 74.200 ;
        RECT 155.800 73.800 160.200 74.100 ;
        RECT 175.000 74.100 175.400 74.200 ;
        RECT 198.200 74.100 198.600 74.200 ;
        RECT 199.000 74.100 199.400 74.200 ;
        RECT 175.000 73.800 199.400 74.100 ;
        RECT 109.400 73.200 109.700 73.800 ;
        RECT 147.000 73.200 147.300 73.800 ;
        RECT 39.800 73.100 40.200 73.200 ;
        RECT 43.800 73.100 44.200 73.200 ;
        RECT 39.800 72.800 44.200 73.100 ;
        RECT 55.800 73.100 56.200 73.200 ;
        RECT 65.400 73.100 65.800 73.200 ;
        RECT 55.800 72.800 65.800 73.100 ;
        RECT 72.600 73.100 73.000 73.200 ;
        RECT 83.000 73.100 83.400 73.200 ;
        RECT 72.600 72.800 83.400 73.100 ;
        RECT 95.000 73.100 95.400 73.200 ;
        RECT 104.600 73.100 105.000 73.200 ;
        RECT 95.000 72.800 105.000 73.100 ;
        RECT 109.400 72.800 109.800 73.200 ;
        RECT 117.400 72.800 117.800 73.200 ;
        RECT 147.000 72.800 147.400 73.200 ;
        RECT 175.800 73.100 176.200 73.200 ;
        RECT 177.400 73.100 177.800 73.200 ;
        RECT 175.800 72.800 177.800 73.100 ;
        RECT 183.000 73.100 183.400 73.200 ;
        RECT 183.800 73.100 184.200 73.200 ;
        RECT 183.000 72.800 184.200 73.100 ;
        RECT 196.600 73.100 197.000 73.200 ;
        RECT 201.400 73.100 201.800 73.200 ;
        RECT 196.600 72.800 201.800 73.100 ;
        RECT 211.000 73.100 211.400 73.200 ;
        RECT 219.000 73.100 219.400 73.200 ;
        RECT 220.600 73.100 221.000 73.200 ;
        RECT 211.000 72.800 221.000 73.100 ;
        RECT 10.200 72.100 10.600 72.200 ;
        RECT 11.000 72.100 11.400 72.200 ;
        RECT 13.400 72.100 13.800 72.200 ;
        RECT 16.600 72.100 17.000 72.200 ;
        RECT 10.200 71.800 17.000 72.100 ;
        RECT 39.000 72.100 39.400 72.200 ;
        RECT 40.600 72.100 41.000 72.200 ;
        RECT 39.000 71.800 41.000 72.100 ;
        RECT 41.400 72.100 41.800 72.200 ;
        RECT 42.200 72.100 42.600 72.200 ;
        RECT 41.400 71.800 42.600 72.100 ;
        RECT 67.800 72.100 68.200 72.200 ;
        RECT 87.000 72.100 87.400 72.200 ;
        RECT 102.200 72.100 102.600 72.200 ;
        RECT 67.800 71.800 102.600 72.100 ;
        RECT 109.400 72.100 109.800 72.200 ;
        RECT 113.400 72.100 113.800 72.200 ;
        RECT 117.400 72.100 117.700 72.800 ;
        RECT 109.400 71.800 113.800 72.100 ;
        RECT 114.200 71.800 117.700 72.100 ;
        RECT 135.000 72.100 135.400 72.200 ;
        RECT 139.800 72.100 140.200 72.200 ;
        RECT 151.000 72.100 151.400 72.200 ;
        RECT 135.000 71.800 151.400 72.100 ;
        RECT 153.400 72.100 153.800 72.200 ;
        RECT 155.800 72.100 156.200 72.200 ;
        RECT 153.400 71.800 156.200 72.100 ;
        RECT 165.400 72.100 165.800 72.200 ;
        RECT 177.400 72.100 177.800 72.200 ;
        RECT 165.400 71.800 177.800 72.100 ;
        RECT 185.400 72.100 185.800 72.200 ;
        RECT 203.000 72.100 203.400 72.200 ;
        RECT 210.200 72.100 210.600 72.200 ;
        RECT 218.200 72.100 218.600 72.200 ;
        RECT 185.400 71.800 218.600 72.100 ;
        RECT 12.600 71.100 13.000 71.200 ;
        RECT 35.000 71.100 35.400 71.200 ;
        RECT 55.800 71.100 56.200 71.200 ;
        RECT 12.600 70.800 56.200 71.100 ;
        RECT 105.400 71.100 105.800 71.200 ;
        RECT 106.200 71.100 106.600 71.200 ;
        RECT 114.200 71.100 114.500 71.800 ;
        RECT 105.400 70.800 114.500 71.100 ;
        RECT 116.600 71.100 117.000 71.200 ;
        RECT 125.400 71.100 125.800 71.200 ;
        RECT 116.600 70.800 125.800 71.100 ;
        RECT 143.000 71.100 143.400 71.200 ;
        RECT 158.200 71.100 158.600 71.200 ;
        RECT 143.000 70.800 158.600 71.100 ;
        RECT 176.600 71.100 177.000 71.200 ;
        RECT 188.600 71.100 189.000 71.200 ;
        RECT 176.600 70.800 189.000 71.100 ;
        RECT 45.400 70.100 45.800 70.200 ;
        RECT 52.600 70.100 53.000 70.200 ;
        RECT 45.400 69.800 53.000 70.100 ;
        RECT 62.200 70.100 62.600 70.200 ;
        RECT 63.800 70.100 64.200 70.200 ;
        RECT 62.200 69.800 64.200 70.100 ;
        RECT 95.800 70.100 96.200 70.200 ;
        RECT 111.000 70.100 111.400 70.200 ;
        RECT 113.400 70.100 113.800 70.200 ;
        RECT 95.800 69.800 113.800 70.100 ;
        RECT 114.200 70.100 114.600 70.200 ;
        RECT 129.400 70.100 129.800 70.200 ;
        RECT 114.200 69.800 129.800 70.100 ;
        RECT 130.200 70.100 130.600 70.200 ;
        RECT 151.800 70.100 152.200 70.200 ;
        RECT 130.200 69.800 152.200 70.100 ;
        RECT 168.600 70.100 169.000 70.200 ;
        RECT 171.000 70.100 171.400 70.200 ;
        RECT 168.600 69.800 171.400 70.100 ;
        RECT 171.800 70.100 172.200 70.200 ;
        RECT 183.000 70.100 183.400 70.200 ;
        RECT 204.600 70.100 205.000 70.200 ;
        RECT 227.000 70.100 227.400 70.200 ;
        RECT 171.800 69.800 190.500 70.100 ;
        RECT 204.600 69.800 227.400 70.100 ;
        RECT 31.800 69.100 32.200 69.200 ;
        RECT 35.800 69.100 36.200 69.200 ;
        RECT 31.800 68.800 36.200 69.100 ;
        RECT 58.200 69.100 58.600 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 68.600 69.100 69.000 69.200 ;
        RECT 58.200 68.800 69.000 69.100 ;
        RECT 104.600 69.100 105.000 69.200 ;
        RECT 105.400 69.100 105.800 69.200 ;
        RECT 148.600 69.100 149.000 69.200 ;
        RECT 150.200 69.100 150.600 69.200 ;
        RECT 157.400 69.100 157.800 69.200 ;
        RECT 104.600 68.800 105.800 69.100 ;
        RECT 108.600 68.800 149.000 69.100 ;
        RECT 149.400 68.800 157.800 69.100 ;
        RECT 158.200 69.100 158.600 69.200 ;
        RECT 159.000 69.100 159.400 69.200 ;
        RECT 158.200 68.800 159.400 69.100 ;
        RECT 160.600 69.100 161.000 69.200 ;
        RECT 165.400 69.100 165.800 69.200 ;
        RECT 160.600 68.800 165.800 69.100 ;
        RECT 167.800 69.100 168.200 69.200 ;
        RECT 168.600 69.100 169.000 69.200 ;
        RECT 170.200 69.100 170.600 69.200 ;
        RECT 171.000 69.100 171.400 69.200 ;
        RECT 167.800 68.800 169.000 69.100 ;
        RECT 169.400 68.800 171.400 69.100 ;
        RECT 171.800 69.100 172.200 69.200 ;
        RECT 187.800 69.100 188.200 69.200 ;
        RECT 171.800 68.800 188.200 69.100 ;
        RECT 190.200 69.100 190.500 69.800 ;
        RECT 228.600 69.100 229.000 69.200 ;
        RECT 190.200 68.800 229.000 69.100 ;
        RECT 108.600 68.200 108.900 68.800 ;
        RECT 13.400 68.100 13.800 68.200 ;
        RECT 17.400 68.100 17.800 68.200 ;
        RECT 13.400 67.800 17.800 68.100 ;
        RECT 35.800 68.100 36.200 68.200 ;
        RECT 36.600 68.100 37.000 68.200 ;
        RECT 35.800 67.800 37.000 68.100 ;
        RECT 59.000 68.100 59.400 68.200 ;
        RECT 64.600 68.100 65.000 68.200 ;
        RECT 59.000 67.800 65.000 68.100 ;
        RECT 75.800 67.800 76.200 68.200 ;
        RECT 77.400 67.800 77.800 68.200 ;
        RECT 95.800 67.800 96.200 68.200 ;
        RECT 99.800 67.800 100.200 68.200 ;
        RECT 102.200 68.100 102.600 68.200 ;
        RECT 103.000 68.100 103.400 68.200 ;
        RECT 102.200 67.800 103.400 68.100 ;
        RECT 108.600 67.800 109.000 68.200 ;
        RECT 112.600 68.100 113.000 68.200 ;
        RECT 115.800 68.100 116.200 68.200 ;
        RECT 119.800 68.100 120.200 68.200 ;
        RECT 112.600 67.800 120.200 68.100 ;
        RECT 127.800 68.100 128.200 68.200 ;
        RECT 142.200 68.100 142.600 68.200 ;
        RECT 127.800 67.800 142.600 68.100 ;
        RECT 145.400 68.100 145.800 68.200 ;
        RECT 185.400 68.100 185.800 68.200 ;
        RECT 145.400 67.800 185.800 68.100 ;
        RECT 186.200 67.800 186.600 68.200 ;
        RECT 21.400 67.100 21.800 67.200 ;
        RECT 31.000 67.100 31.400 67.200 ;
        RECT 21.400 66.800 31.400 67.100 ;
        RECT 35.000 67.100 35.400 67.200 ;
        RECT 45.400 67.100 45.800 67.200 ;
        RECT 35.000 66.800 45.800 67.100 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 75.800 67.100 76.100 67.800 ;
        RECT 64.600 66.800 76.100 67.100 ;
        RECT 77.400 67.100 77.700 67.800 ;
        RECT 95.800 67.200 96.100 67.800 ;
        RECT 99.800 67.200 100.100 67.800 ;
        RECT 87.800 67.100 88.200 67.200 ;
        RECT 77.400 66.800 88.200 67.100 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 100.600 67.100 101.000 67.200 ;
        RECT 101.400 67.100 101.800 67.200 ;
        RECT 100.600 66.800 101.800 67.100 ;
        RECT 112.600 67.100 113.000 67.200 ;
        RECT 115.800 67.100 116.200 67.200 ;
        RECT 112.600 66.800 116.200 67.100 ;
        RECT 116.600 67.100 117.000 67.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 123.000 67.100 123.400 67.200 ;
        RECT 116.600 66.800 119.300 67.100 ;
        RECT 121.400 66.800 123.400 67.100 ;
        RECT 128.600 67.100 129.000 67.200 ;
        RECT 154.200 67.100 154.600 67.200 ;
        RECT 128.600 66.800 154.600 67.100 ;
        RECT 155.800 67.100 156.200 67.200 ;
        RECT 156.600 67.100 157.000 67.200 ;
        RECT 155.800 66.800 157.000 67.100 ;
        RECT 167.800 67.100 168.200 67.200 ;
        RECT 172.600 67.100 173.000 67.200 ;
        RECT 174.200 67.100 174.600 67.200 ;
        RECT 167.800 66.800 174.600 67.100 ;
        RECT 175.800 67.100 176.200 67.200 ;
        RECT 176.600 67.100 177.000 67.200 ;
        RECT 175.800 66.800 177.000 67.100 ;
        RECT 183.800 67.100 184.200 67.200 ;
        RECT 186.200 67.100 186.500 67.800 ;
        RECT 183.800 66.800 186.500 67.100 ;
        RECT 9.400 66.100 9.800 66.200 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 9.400 65.800 13.800 66.100 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 47.000 66.100 47.400 66.200 ;
        RECT 31.800 65.800 47.400 66.100 ;
        RECT 55.800 66.100 56.200 66.200 ;
        RECT 66.200 66.100 66.600 66.200 ;
        RECT 55.800 65.800 66.600 66.100 ;
        RECT 75.000 66.100 75.400 66.200 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 75.000 65.800 81.800 66.100 ;
        RECT 88.600 66.100 89.000 66.200 ;
        RECT 98.200 66.100 98.600 66.200 ;
        RECT 103.800 66.100 104.200 66.200 ;
        RECT 106.200 66.100 106.600 66.200 ;
        RECT 88.600 65.800 98.600 66.100 ;
        RECT 103.000 65.800 106.600 66.100 ;
        RECT 112.600 66.100 113.000 66.200 ;
        RECT 113.400 66.100 113.800 66.200 ;
        RECT 112.600 65.800 113.800 66.100 ;
        RECT 115.800 66.100 116.200 66.200 ;
        RECT 118.200 66.100 118.600 66.200 ;
        RECT 115.800 65.800 118.600 66.100 ;
        RECT 119.000 66.100 119.300 66.800 ;
        RECT 133.400 66.100 133.800 66.200 ;
        RECT 119.000 65.800 133.800 66.100 ;
        RECT 141.400 66.100 141.800 66.200 ;
        RECT 142.200 66.100 142.600 66.200 ;
        RECT 145.400 66.100 145.800 66.200 ;
        RECT 141.400 65.800 145.800 66.100 ;
        RECT 146.200 65.800 146.600 66.200 ;
        RECT 149.400 66.100 149.800 66.200 ;
        RECT 189.400 66.100 189.800 66.200 ;
        RECT 190.200 66.100 190.600 66.200 ;
        RECT 149.400 65.800 190.600 66.100 ;
        RECT 203.800 66.100 204.200 66.200 ;
        RECT 207.800 66.100 208.200 66.200 ;
        RECT 203.800 65.800 208.200 66.100 ;
        RECT 209.400 66.100 209.800 66.200 ;
        RECT 216.600 66.100 217.000 66.200 ;
        RECT 209.400 65.800 217.000 66.100 ;
        RECT 224.600 65.800 225.000 66.200 ;
        RECT 17.400 65.100 17.800 65.200 ;
        RECT 20.600 65.100 21.000 65.200 ;
        RECT 17.400 64.800 21.000 65.100 ;
        RECT 42.200 65.100 42.600 65.200 ;
        RECT 43.000 65.100 43.400 65.200 ;
        RECT 42.200 64.800 43.400 65.100 ;
        RECT 53.400 65.100 53.800 65.200 ;
        RECT 63.000 65.100 63.400 65.200 ;
        RECT 53.400 64.800 63.400 65.100 ;
        RECT 67.000 64.800 67.400 65.200 ;
        RECT 68.600 65.100 69.000 65.200 ;
        RECT 73.400 65.100 73.800 65.200 ;
        RECT 75.000 65.100 75.400 65.200 ;
        RECT 76.600 65.100 77.000 65.200 ;
        RECT 68.600 64.800 77.000 65.100 ;
        RECT 93.400 65.100 93.800 65.200 ;
        RECT 103.000 65.100 103.400 65.200 ;
        RECT 104.600 65.100 105.000 65.200 ;
        RECT 93.400 64.800 105.000 65.100 ;
        RECT 107.800 65.100 108.200 65.200 ;
        RECT 117.400 65.100 117.800 65.200 ;
        RECT 127.800 65.100 128.200 65.200 ;
        RECT 107.800 64.800 128.200 65.100 ;
        RECT 135.800 65.100 136.200 65.200 ;
        RECT 141.400 65.100 141.800 65.200 ;
        RECT 135.800 64.800 141.800 65.100 ;
        RECT 146.200 65.100 146.500 65.800 ;
        RECT 224.600 65.200 224.900 65.800 ;
        RECT 148.600 65.100 149.000 65.200 ;
        RECT 146.200 64.800 149.000 65.100 ;
        RECT 163.800 64.800 164.200 65.200 ;
        RECT 165.400 65.100 165.800 65.200 ;
        RECT 171.000 65.100 171.400 65.200 ;
        RECT 172.600 65.100 173.000 65.200 ;
        RECT 165.400 64.800 173.000 65.100 ;
        RECT 186.200 64.800 186.600 65.200 ;
        RECT 199.800 65.100 200.200 65.200 ;
        RECT 204.600 65.100 205.000 65.200 ;
        RECT 199.800 64.800 205.000 65.100 ;
        RECT 209.400 65.100 209.800 65.200 ;
        RECT 210.200 65.100 210.600 65.200 ;
        RECT 209.400 64.800 210.600 65.100 ;
        RECT 224.600 64.800 225.000 65.200 ;
        RECT 0.600 64.100 1.000 64.200 ;
        RECT 3.800 64.100 4.200 64.200 ;
        RECT 37.400 64.100 37.800 64.200 ;
        RECT 43.000 64.100 43.400 64.200 ;
        RECT 0.600 63.800 43.400 64.100 ;
        RECT 62.200 64.100 62.600 64.200 ;
        RECT 67.000 64.100 67.300 64.800 ;
        RECT 71.000 64.100 71.400 64.200 ;
        RECT 62.200 63.800 71.400 64.100 ;
        RECT 108.600 64.100 109.000 64.200 ;
        RECT 110.200 64.100 110.600 64.200 ;
        RECT 108.600 63.800 110.600 64.100 ;
        RECT 121.400 64.100 121.800 64.200 ;
        RECT 122.200 64.100 122.600 64.200 ;
        RECT 121.400 63.800 122.600 64.100 ;
        RECT 144.600 64.100 145.000 64.200 ;
        RECT 151.800 64.100 152.200 64.200 ;
        RECT 144.600 63.800 152.200 64.100 ;
        RECT 163.800 64.100 164.100 64.800 ;
        RECT 186.200 64.200 186.500 64.800 ;
        RECT 167.800 64.100 168.200 64.200 ;
        RECT 163.800 63.800 168.200 64.100 ;
        RECT 186.200 63.800 186.600 64.200 ;
        RECT 193.400 64.100 193.800 64.200 ;
        RECT 194.200 64.100 194.600 64.200 ;
        RECT 193.400 63.800 194.600 64.100 ;
        RECT 201.400 64.100 201.800 64.200 ;
        RECT 212.600 64.100 213.000 64.200 ;
        RECT 201.400 63.800 213.700 64.100 ;
        RECT 29.400 63.100 29.800 63.200 ;
        RECT 39.800 63.100 40.200 63.200 ;
        RECT 29.400 62.800 40.200 63.100 ;
        RECT 47.000 62.800 47.400 63.200 ;
        RECT 58.200 63.100 58.600 63.200 ;
        RECT 76.600 63.100 77.000 63.200 ;
        RECT 58.200 62.800 77.000 63.100 ;
        RECT 91.000 63.100 91.400 63.200 ;
        RECT 109.400 63.100 109.800 63.200 ;
        RECT 91.000 62.800 109.800 63.100 ;
        RECT 122.200 63.100 122.600 63.200 ;
        RECT 126.200 63.100 126.600 63.200 ;
        RECT 122.200 62.800 126.600 63.100 ;
        RECT 144.600 63.100 145.000 63.200 ;
        RECT 163.000 63.100 163.400 63.200 ;
        RECT 144.600 62.800 163.400 63.100 ;
        RECT 177.400 63.100 177.800 63.200 ;
        RECT 199.800 63.100 200.200 63.200 ;
        RECT 177.400 62.800 200.200 63.100 ;
        RECT 210.200 63.100 210.600 63.200 ;
        RECT 211.000 63.100 211.400 63.200 ;
        RECT 229.400 63.100 229.800 63.200 ;
        RECT 210.200 62.800 229.800 63.100 ;
        RECT 47.000 62.100 47.300 62.800 ;
        RECT 162.200 62.100 162.600 62.200 ;
        RECT 47.000 61.800 162.600 62.100 ;
        RECT 211.000 62.100 211.400 62.200 ;
        RECT 214.200 62.100 214.600 62.200 ;
        RECT 211.000 61.800 214.600 62.100 ;
        RECT 70.200 61.100 70.600 61.200 ;
        RECT 111.000 61.100 111.400 61.200 ;
        RECT 138.200 61.100 138.600 61.200 ;
        RECT 70.200 60.800 110.500 61.100 ;
        RECT 111.000 60.800 138.600 61.100 ;
        RECT 143.000 61.100 143.400 61.200 ;
        RECT 191.000 61.100 191.400 61.200 ;
        RECT 143.000 60.800 191.400 61.100 ;
        RECT 16.600 60.100 17.000 60.200 ;
        RECT 17.400 60.100 17.800 60.200 ;
        RECT 16.600 59.800 17.800 60.100 ;
        RECT 44.600 60.100 45.000 60.200 ;
        RECT 59.000 60.100 59.400 60.200 ;
        RECT 61.400 60.100 61.800 60.200 ;
        RECT 72.600 60.100 73.000 60.200 ;
        RECT 44.600 59.800 73.000 60.100 ;
        RECT 79.000 60.100 79.400 60.200 ;
        RECT 80.600 60.100 81.000 60.200 ;
        RECT 79.000 59.800 81.000 60.100 ;
        RECT 84.600 60.100 85.000 60.200 ;
        RECT 94.200 60.100 94.600 60.200 ;
        RECT 84.600 59.800 94.600 60.100 ;
        RECT 110.200 60.100 110.500 60.800 ;
        RECT 116.600 60.100 117.000 60.200 ;
        RECT 110.200 59.800 117.000 60.100 ;
        RECT 155.000 60.100 155.400 60.200 ;
        RECT 160.600 60.100 161.000 60.200 ;
        RECT 155.000 59.800 161.000 60.100 ;
        RECT 189.400 60.100 189.800 60.200 ;
        RECT 193.400 60.100 193.800 60.200 ;
        RECT 206.200 60.100 206.600 60.200 ;
        RECT 189.400 59.800 206.600 60.100 ;
        RECT 43.000 59.100 43.400 59.200 ;
        RECT 71.800 59.100 72.200 59.200 ;
        RECT 43.000 58.800 72.200 59.100 ;
        RECT 79.000 59.100 79.400 59.200 ;
        RECT 115.800 59.100 116.200 59.200 ;
        RECT 132.600 59.100 133.000 59.200 ;
        RECT 147.000 59.100 147.400 59.200 ;
        RECT 79.000 58.800 116.200 59.100 ;
        RECT 131.800 58.800 147.400 59.100 ;
        RECT 161.400 59.100 161.800 59.200 ;
        RECT 166.200 59.100 166.600 59.200 ;
        RECT 161.400 58.800 166.600 59.100 ;
        RECT 178.200 59.100 178.600 59.200 ;
        RECT 215.000 59.100 215.400 59.200 ;
        RECT 178.200 58.800 215.400 59.100 ;
        RECT 16.600 57.800 17.000 58.200 ;
        RECT 19.000 57.800 19.400 58.200 ;
        RECT 34.200 58.100 34.600 58.200 ;
        RECT 55.000 58.100 55.400 58.200 ;
        RECT 34.200 57.800 55.400 58.100 ;
        RECT 56.600 57.800 57.000 58.200 ;
        RECT 72.600 58.100 73.000 58.200 ;
        RECT 95.800 58.100 96.200 58.200 ;
        RECT 72.600 57.800 96.200 58.100 ;
        RECT 96.600 58.100 97.000 58.200 ;
        RECT 102.200 58.100 102.600 58.200 ;
        RECT 96.600 57.800 102.600 58.100 ;
        RECT 115.800 58.100 116.200 58.200 ;
        RECT 120.600 58.100 121.000 58.200 ;
        RECT 115.800 57.800 121.000 58.100 ;
        RECT 121.400 57.800 121.800 58.200 ;
        RECT 142.200 58.100 142.600 58.200 ;
        RECT 161.400 58.100 161.800 58.200 ;
        RECT 179.800 58.100 180.200 58.200 ;
        RECT 142.200 57.800 180.200 58.100 ;
        RECT 183.800 58.100 184.200 58.200 ;
        RECT 188.600 58.100 189.000 58.200 ;
        RECT 183.800 57.800 189.000 58.100 ;
        RECT 7.000 57.100 7.400 57.200 ;
        RECT 16.600 57.100 16.900 57.800 ;
        RECT 7.000 56.800 16.900 57.100 ;
        RECT 19.000 57.200 19.300 57.800 ;
        RECT 19.000 57.100 19.400 57.200 ;
        RECT 29.400 57.100 29.800 57.200 ;
        RECT 19.000 56.800 29.800 57.100 ;
        RECT 30.200 57.100 30.600 57.200 ;
        RECT 31.000 57.100 31.400 57.200 ;
        RECT 35.000 57.100 35.400 57.200 ;
        RECT 30.200 56.800 35.400 57.100 ;
        RECT 42.200 57.100 42.600 57.200 ;
        RECT 43.000 57.100 43.400 57.200 ;
        RECT 42.200 56.800 43.400 57.100 ;
        RECT 45.400 57.100 45.800 57.200 ;
        RECT 50.200 57.100 50.600 57.200 ;
        RECT 45.400 56.800 50.600 57.100 ;
        RECT 53.400 57.100 53.800 57.200 ;
        RECT 56.600 57.100 56.900 57.800 ;
        RECT 53.400 56.800 56.900 57.100 ;
        RECT 65.400 57.100 65.800 57.200 ;
        RECT 75.000 57.100 75.400 57.200 ;
        RECT 65.400 56.800 75.400 57.100 ;
        RECT 103.000 57.100 103.400 57.200 ;
        RECT 104.600 57.100 105.000 57.200 ;
        RECT 103.000 56.800 105.000 57.100 ;
        RECT 107.800 57.100 108.200 57.200 ;
        RECT 109.400 57.100 109.800 57.200 ;
        RECT 107.800 56.800 109.800 57.100 ;
        RECT 117.400 57.100 117.800 57.200 ;
        RECT 119.000 57.100 119.400 57.200 ;
        RECT 117.400 56.800 119.400 57.100 ;
        RECT 120.600 57.100 121.000 57.200 ;
        RECT 121.400 57.100 121.700 57.800 ;
        RECT 120.600 56.800 121.700 57.100 ;
        RECT 123.000 57.100 123.400 57.200 ;
        RECT 123.800 57.100 124.200 57.200 ;
        RECT 123.000 56.800 124.200 57.100 ;
        RECT 128.600 57.100 129.000 57.200 ;
        RECT 129.400 57.100 129.800 57.200 ;
        RECT 128.600 56.800 129.800 57.100 ;
        RECT 131.800 57.100 132.200 57.200 ;
        RECT 132.600 57.100 133.000 57.200 ;
        RECT 131.800 56.800 133.000 57.100 ;
        RECT 135.800 57.100 136.200 57.200 ;
        RECT 151.800 57.100 152.200 57.200 ;
        RECT 166.200 57.100 166.600 57.200 ;
        RECT 174.200 57.100 174.600 57.200 ;
        RECT 135.800 56.800 152.200 57.100 ;
        RECT 165.400 56.800 174.600 57.100 ;
        RECT 195.800 57.100 196.200 57.200 ;
        RECT 203.000 57.100 203.400 57.200 ;
        RECT 195.800 56.800 203.400 57.100 ;
        RECT 12.600 56.100 13.000 56.200 ;
        RECT 20.600 56.100 21.000 56.200 ;
        RECT 12.600 55.800 21.000 56.100 ;
        RECT 45.400 56.100 45.800 56.200 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 59.800 56.100 60.200 56.200 ;
        RECT 45.400 55.800 60.200 56.100 ;
        RECT 77.400 55.800 77.800 56.200 ;
        RECT 103.800 56.100 104.200 56.200 ;
        RECT 105.400 56.100 105.800 56.200 ;
        RECT 103.800 55.800 105.800 56.100 ;
        RECT 107.000 56.100 107.400 56.200 ;
        RECT 111.800 56.100 112.200 56.200 ;
        RECT 115.800 56.100 116.200 56.200 ;
        RECT 107.000 55.800 116.200 56.100 ;
        RECT 120.600 56.100 121.000 56.200 ;
        RECT 124.600 56.100 125.000 56.200 ;
        RECT 135.000 56.100 135.400 56.200 ;
        RECT 120.600 55.800 135.400 56.100 ;
        RECT 143.800 56.100 144.200 56.200 ;
        RECT 183.800 56.100 184.200 56.200 ;
        RECT 143.800 55.800 184.200 56.100 ;
        RECT 184.600 55.800 185.000 56.200 ;
        RECT 190.200 56.100 190.600 56.200 ;
        RECT 206.200 56.100 206.600 56.200 ;
        RECT 190.200 55.800 206.600 56.100 ;
        RECT 207.000 56.100 207.400 56.200 ;
        RECT 213.400 56.100 213.800 56.200 ;
        RECT 227.000 56.100 227.400 56.200 ;
        RECT 207.000 55.800 227.400 56.100 ;
        RECT 8.600 55.100 9.000 55.200 ;
        RECT 15.000 55.100 15.400 55.200 ;
        RECT 8.600 54.800 15.400 55.100 ;
        RECT 15.800 55.100 16.200 55.200 ;
        RECT 19.000 55.100 19.400 55.200 ;
        RECT 15.800 54.800 19.400 55.100 ;
        RECT 27.000 55.100 27.400 55.200 ;
        RECT 36.600 55.100 37.000 55.200 ;
        RECT 27.000 54.800 37.000 55.100 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 40.600 54.800 46.600 55.100 ;
        RECT 51.800 55.100 52.200 55.200 ;
        RECT 55.800 55.100 56.200 55.200 ;
        RECT 51.800 54.800 56.200 55.100 ;
        RECT 61.400 54.800 61.800 55.200 ;
        RECT 77.400 55.100 77.700 55.800 ;
        RECT 111.800 55.100 112.200 55.200 ;
        RECT 141.400 55.100 141.800 55.200 ;
        RECT 77.400 54.800 141.800 55.100 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 148.600 54.800 149.000 55.200 ;
        RECT 163.000 55.100 163.400 55.200 ;
        RECT 164.600 55.100 165.000 55.200 ;
        RECT 163.000 54.800 165.000 55.100 ;
        RECT 172.600 54.800 173.000 55.200 ;
        RECT 173.400 55.100 173.800 55.200 ;
        RECT 182.200 55.100 182.600 55.200 ;
        RECT 184.600 55.100 184.900 55.800 ;
        RECT 173.400 54.800 184.900 55.100 ;
        RECT 191.000 55.100 191.400 55.200 ;
        RECT 194.200 55.100 194.600 55.200 ;
        RECT 191.000 54.800 194.600 55.100 ;
        RECT 200.600 55.100 201.000 55.200 ;
        RECT 201.400 55.100 201.800 55.200 ;
        RECT 200.600 54.800 201.800 55.100 ;
        RECT 203.000 55.100 203.400 55.200 ;
        RECT 209.400 55.100 209.800 55.200 ;
        RECT 217.400 55.100 217.800 55.200 ;
        RECT 221.400 55.100 221.800 55.200 ;
        RECT 203.000 54.800 209.800 55.100 ;
        RECT 216.600 54.800 221.800 55.100 ;
        RECT 3.000 54.100 3.400 54.200 ;
        RECT 9.400 54.100 9.800 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 3.000 53.800 15.400 54.100 ;
        RECT 20.600 54.100 21.000 54.200 ;
        RECT 27.800 54.100 28.200 54.200 ;
        RECT 20.600 53.800 28.200 54.100 ;
        RECT 32.600 54.100 33.000 54.200 ;
        RECT 45.400 54.100 45.800 54.200 ;
        RECT 46.200 54.100 46.600 54.200 ;
        RECT 32.600 53.800 46.600 54.100 ;
        RECT 56.600 54.100 57.000 54.200 ;
        RECT 57.400 54.100 57.800 54.200 ;
        RECT 56.600 53.800 57.800 54.100 ;
        RECT 61.400 54.100 61.700 54.800 ;
        RECT 147.800 54.200 148.100 54.800 ;
        RECT 64.600 54.100 65.000 54.200 ;
        RECT 61.400 53.800 65.000 54.100 ;
        RECT 74.200 54.100 74.600 54.200 ;
        RECT 78.200 54.100 78.600 54.200 ;
        RECT 74.200 53.800 78.600 54.100 ;
        RECT 81.400 54.100 81.800 54.200 ;
        RECT 85.400 54.100 85.800 54.200 ;
        RECT 81.400 53.800 85.800 54.100 ;
        RECT 87.000 54.100 87.400 54.200 ;
        RECT 89.400 54.100 89.800 54.200 ;
        RECT 87.000 53.800 89.800 54.100 ;
        RECT 118.200 54.100 118.600 54.200 ;
        RECT 122.200 54.100 122.600 54.200 ;
        RECT 118.200 53.800 122.600 54.100 ;
        RECT 125.400 54.100 125.800 54.200 ;
        RECT 126.200 54.100 126.600 54.200 ;
        RECT 125.400 53.800 126.600 54.100 ;
        RECT 127.000 54.100 127.400 54.200 ;
        RECT 130.200 54.100 130.600 54.200 ;
        RECT 127.000 53.800 130.600 54.100 ;
        RECT 134.200 54.100 134.600 54.200 ;
        RECT 136.600 54.100 137.000 54.200 ;
        RECT 134.200 53.800 137.000 54.100 ;
        RECT 138.200 54.100 138.600 54.200 ;
        RECT 146.200 54.100 146.600 54.200 ;
        RECT 138.200 53.800 146.600 54.100 ;
        RECT 147.800 53.800 148.200 54.200 ;
        RECT 148.600 54.100 148.900 54.800 ;
        RECT 149.400 54.100 149.800 54.200 ;
        RECT 148.600 53.800 149.800 54.100 ;
        RECT 157.400 54.100 157.800 54.200 ;
        RECT 172.600 54.100 172.900 54.800 ;
        RECT 157.400 53.800 172.900 54.100 ;
        RECT 185.400 54.100 185.800 54.200 ;
        RECT 188.600 54.100 189.000 54.200 ;
        RECT 228.600 54.100 229.000 54.200 ;
        RECT 185.400 53.800 189.000 54.100 ;
        RECT 214.200 53.800 229.000 54.100 ;
        RECT 214.200 53.200 214.500 53.800 ;
        RECT 19.800 53.100 20.200 53.200 ;
        RECT 28.600 53.100 29.000 53.200 ;
        RECT 31.800 53.100 32.200 53.200 ;
        RECT 41.400 53.100 41.800 53.200 ;
        RECT 19.800 52.800 41.800 53.100 ;
        RECT 76.600 53.100 77.000 53.200 ;
        RECT 84.600 53.100 85.000 53.200 ;
        RECT 91.000 53.100 91.400 53.200 ;
        RECT 76.600 52.800 91.400 53.100 ;
        RECT 124.600 53.100 125.000 53.200 ;
        RECT 125.400 53.100 125.800 53.200 ;
        RECT 124.600 52.800 125.800 53.100 ;
        RECT 143.000 53.100 143.400 53.200 ;
        RECT 144.600 53.100 145.000 53.200 ;
        RECT 150.200 53.100 150.600 53.200 ;
        RECT 143.000 52.800 145.000 53.100 ;
        RECT 145.400 52.800 150.600 53.100 ;
        RECT 167.000 53.100 167.400 53.200 ;
        RECT 179.000 53.100 179.400 53.200 ;
        RECT 167.000 52.800 179.400 53.100 ;
        RECT 187.800 53.100 188.200 53.200 ;
        RECT 202.200 53.100 202.600 53.200 ;
        RECT 187.800 52.800 203.300 53.100 ;
        RECT 214.200 52.800 214.600 53.200 ;
        RECT 145.400 52.200 145.700 52.800 ;
        RECT 56.600 52.100 57.000 52.200 ;
        RECT 99.000 52.100 99.400 52.200 ;
        RECT 56.600 51.800 99.400 52.100 ;
        RECT 109.400 52.100 109.800 52.200 ;
        RECT 123.000 52.100 123.400 52.200 ;
        RECT 132.600 52.100 133.000 52.200 ;
        RECT 143.800 52.100 144.200 52.200 ;
        RECT 109.400 51.800 144.200 52.100 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 146.200 52.100 146.600 52.200 ;
        RECT 169.400 52.100 169.800 52.200 ;
        RECT 146.200 51.800 169.800 52.100 ;
        RECT 200.600 52.100 201.000 52.200 ;
        RECT 214.200 52.100 214.600 52.200 ;
        RECT 216.600 52.100 217.000 52.200 ;
        RECT 200.600 51.800 217.000 52.100 ;
        RECT 15.000 51.100 15.400 51.200 ;
        RECT 17.400 51.100 17.800 51.200 ;
        RECT 32.600 51.100 33.000 51.200 ;
        RECT 15.000 50.800 33.000 51.100 ;
        RECT 95.000 51.100 95.400 51.200 ;
        RECT 119.000 51.100 119.400 51.200 ;
        RECT 190.200 51.100 190.600 51.200 ;
        RECT 95.000 50.800 190.600 51.100 ;
        RECT 201.400 51.100 201.800 51.200 ;
        RECT 205.400 51.100 205.800 51.200 ;
        RECT 201.400 50.800 205.800 51.100 ;
        RECT 94.200 50.100 94.600 50.200 ;
        RECT 101.400 50.100 101.800 50.200 ;
        RECT 94.200 49.800 101.800 50.100 ;
        RECT 103.000 50.100 103.400 50.200 ;
        RECT 127.800 50.100 128.200 50.200 ;
        RECT 140.600 50.100 141.000 50.200 ;
        RECT 147.800 50.100 148.200 50.200 ;
        RECT 163.000 50.100 163.400 50.200 ;
        RECT 165.400 50.100 165.800 50.200 ;
        RECT 166.200 50.100 166.600 50.200 ;
        RECT 103.000 49.800 166.600 50.100 ;
        RECT 195.000 50.100 195.400 50.200 ;
        RECT 210.200 50.100 210.600 50.200 ;
        RECT 195.000 49.800 210.600 50.100 ;
        RECT 211.000 50.100 211.400 50.200 ;
        RECT 219.800 50.100 220.200 50.200 ;
        RECT 211.000 49.800 220.200 50.100 ;
        RECT 12.600 48.800 13.000 49.200 ;
        RECT 30.200 48.800 30.600 49.200 ;
        RECT 47.000 49.100 47.400 49.200 ;
        RECT 51.800 49.100 52.200 49.200 ;
        RECT 47.000 48.800 52.200 49.100 ;
        RECT 99.800 49.100 100.200 49.200 ;
        RECT 107.800 49.100 108.200 49.200 ;
        RECT 108.600 49.100 109.000 49.200 ;
        RECT 99.800 48.800 109.000 49.100 ;
        RECT 131.800 49.100 132.200 49.200 ;
        RECT 137.400 49.100 137.800 49.200 ;
        RECT 131.800 48.800 137.800 49.100 ;
        RECT 151.000 49.100 151.400 49.200 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 167.800 49.100 168.200 49.200 ;
        RECT 151.000 48.800 168.200 49.100 ;
        RECT 192.600 49.100 193.000 49.200 ;
        RECT 194.200 49.100 194.600 49.200 ;
        RECT 192.600 48.800 194.600 49.100 ;
        RECT 203.800 49.100 204.200 49.200 ;
        RECT 217.400 49.100 217.800 49.200 ;
        RECT 219.000 49.100 219.400 49.200 ;
        RECT 203.800 48.800 219.400 49.100 ;
        RECT 3.800 48.100 4.200 48.200 ;
        RECT 12.600 48.100 12.900 48.800 ;
        RECT 15.800 48.100 16.200 48.200 ;
        RECT 3.800 47.800 12.900 48.100 ;
        RECT 13.400 47.800 16.200 48.100 ;
        RECT 22.200 48.100 22.600 48.200 ;
        RECT 30.200 48.100 30.500 48.800 ;
        RECT 22.200 47.800 30.500 48.100 ;
        RECT 73.400 48.100 73.800 48.200 ;
        RECT 95.000 48.100 95.400 48.200 ;
        RECT 73.400 47.800 95.400 48.100 ;
        RECT 113.400 48.100 113.800 48.200 ;
        RECT 125.400 48.100 125.800 48.200 ;
        RECT 142.200 48.100 142.600 48.200 ;
        RECT 147.000 48.100 147.400 48.200 ;
        RECT 113.400 47.800 147.400 48.100 ;
        RECT 181.400 48.100 181.800 48.200 ;
        RECT 201.400 48.100 201.800 48.200 ;
        RECT 181.400 47.800 201.800 48.100 ;
        RECT 205.400 48.100 205.800 48.200 ;
        RECT 207.000 48.100 207.400 48.200 ;
        RECT 208.600 48.100 209.000 48.200 ;
        RECT 205.400 47.800 209.000 48.100 ;
        RECT 10.200 47.100 10.600 47.200 ;
        RECT 13.400 47.100 13.700 47.800 ;
        RECT 10.200 46.800 13.700 47.100 ;
        RECT 14.200 47.100 14.600 47.200 ;
        RECT 47.800 47.100 48.200 47.200 ;
        RECT 50.200 47.100 50.600 47.200 ;
        RECT 14.200 46.800 50.600 47.100 ;
        RECT 75.000 46.800 75.400 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 87.800 47.100 88.200 47.200 ;
        RECT 81.400 46.800 88.200 47.100 ;
        RECT 97.400 47.100 97.800 47.200 ;
        RECT 103.000 47.100 103.400 47.200 ;
        RECT 97.400 46.800 103.400 47.100 ;
        RECT 137.400 46.800 137.800 47.200 ;
        RECT 149.400 46.800 149.800 47.200 ;
        RECT 180.600 47.100 181.000 47.200 ;
        RECT 183.800 47.100 184.200 47.200 ;
        RECT 196.600 47.100 197.000 47.200 ;
        RECT 200.600 47.100 201.000 47.200 ;
        RECT 203.000 47.100 203.400 47.200 ;
        RECT 180.600 46.800 203.400 47.100 ;
        RECT 203.800 47.100 204.200 47.200 ;
        RECT 211.800 47.100 212.200 47.200 ;
        RECT 216.600 47.100 217.000 47.200 ;
        RECT 203.800 46.800 212.200 47.100 ;
        RECT 213.400 46.800 217.000 47.100 ;
        RECT 11.800 46.100 12.200 46.200 ;
        RECT 13.400 46.100 13.800 46.200 ;
        RECT 11.800 45.800 13.800 46.100 ;
        RECT 27.000 46.100 27.400 46.200 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 27.000 45.800 28.200 46.100 ;
        RECT 29.400 46.100 29.800 46.200 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 29.400 45.800 32.200 46.100 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 33.400 46.100 33.800 46.200 ;
        RECT 32.600 45.800 33.800 46.100 ;
        RECT 41.400 46.100 41.800 46.200 ;
        RECT 49.400 46.100 49.800 46.200 ;
        RECT 41.400 45.800 49.800 46.100 ;
        RECT 58.200 46.100 58.600 46.200 ;
        RECT 62.200 46.100 62.600 46.200 ;
        RECT 58.200 45.800 62.600 46.100 ;
        RECT 70.200 46.100 70.600 46.200 ;
        RECT 75.000 46.100 75.300 46.800 ;
        RECT 137.400 46.200 137.700 46.800 ;
        RECT 70.200 45.800 75.300 46.100 ;
        RECT 96.600 46.100 97.000 46.200 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 96.600 45.800 98.600 46.100 ;
        RECT 106.200 46.100 106.600 46.200 ;
        RECT 137.400 46.100 137.800 46.200 ;
        RECT 139.000 46.100 139.400 46.200 ;
        RECT 148.600 46.100 149.000 46.200 ;
        RECT 106.200 45.800 117.700 46.100 ;
        RECT 137.400 45.800 149.000 46.100 ;
        RECT 149.400 46.100 149.700 46.800 ;
        RECT 213.400 46.200 213.700 46.800 ;
        RECT 166.200 46.100 166.600 46.200 ;
        RECT 173.400 46.100 173.800 46.200 ;
        RECT 149.400 45.800 153.700 46.100 ;
        RECT 166.200 45.800 173.800 46.100 ;
        RECT 179.000 46.100 179.400 46.200 ;
        RECT 207.800 46.100 208.200 46.200 ;
        RECT 208.600 46.100 209.000 46.200 ;
        RECT 179.000 45.800 209.000 46.100 ;
        RECT 210.200 46.100 210.600 46.200 ;
        RECT 210.200 45.800 212.900 46.100 ;
        RECT 213.400 45.800 213.800 46.200 ;
        RECT 219.800 46.100 220.200 46.200 ;
        RECT 223.800 46.100 224.200 46.200 ;
        RECT 219.800 45.800 224.200 46.100 ;
        RECT 117.400 45.200 117.700 45.800 ;
        RECT 153.400 45.200 153.700 45.800 ;
        RECT 212.600 45.200 212.900 45.800 ;
        RECT 16.600 45.100 17.000 45.200 ;
        RECT 35.000 45.100 35.400 45.200 ;
        RECT 16.600 44.800 35.400 45.100 ;
        RECT 44.600 45.100 45.000 45.200 ;
        RECT 55.800 45.100 56.200 45.200 ;
        RECT 44.600 44.800 56.200 45.100 ;
        RECT 64.600 45.100 65.000 45.200 ;
        RECT 77.400 45.100 77.800 45.200 ;
        RECT 64.600 44.800 77.800 45.100 ;
        RECT 79.000 45.100 79.400 45.200 ;
        RECT 80.600 45.100 81.000 45.200 ;
        RECT 79.000 44.800 81.000 45.100 ;
        RECT 109.400 45.100 109.800 45.200 ;
        RECT 112.600 45.100 113.000 45.200 ;
        RECT 109.400 44.800 113.000 45.100 ;
        RECT 117.400 44.800 117.800 45.200 ;
        RECT 132.600 45.100 133.000 45.200 ;
        RECT 144.600 45.100 145.000 45.200 ;
        RECT 132.600 44.800 145.000 45.100 ;
        RECT 153.400 44.800 153.800 45.200 ;
        RECT 163.800 45.100 164.200 45.200 ;
        RECT 167.000 45.100 167.400 45.200 ;
        RECT 203.000 45.100 203.400 45.200 ;
        RECT 163.800 44.800 203.400 45.100 ;
        RECT 212.600 44.800 213.000 45.200 ;
        RECT 14.200 44.100 14.600 44.200 ;
        RECT 52.600 44.100 53.000 44.200 ;
        RECT 14.200 43.800 53.000 44.100 ;
        RECT 71.000 44.100 71.400 44.200 ;
        RECT 82.200 44.100 82.600 44.200 ;
        RECT 90.200 44.100 90.600 44.200 ;
        RECT 71.000 43.800 90.600 44.100 ;
        RECT 99.000 44.100 99.400 44.200 ;
        RECT 110.200 44.100 110.600 44.200 ;
        RECT 99.000 43.800 110.600 44.100 ;
        RECT 120.600 44.100 121.000 44.200 ;
        RECT 125.400 44.100 125.800 44.200 ;
        RECT 135.800 44.100 136.200 44.200 ;
        RECT 120.600 43.800 136.200 44.100 ;
        RECT 153.400 43.800 153.800 44.200 ;
        RECT 184.600 44.100 185.000 44.200 ;
        RECT 185.400 44.100 185.800 44.200 ;
        RECT 184.600 43.800 185.800 44.100 ;
        RECT 207.000 44.100 207.400 44.200 ;
        RECT 219.800 44.100 220.200 44.200 ;
        RECT 207.000 43.800 220.200 44.100 ;
        RECT 153.400 43.200 153.700 43.800 ;
        RECT 16.600 43.100 17.000 43.200 ;
        RECT 53.400 43.100 53.800 43.200 ;
        RECT 103.800 43.100 104.200 43.200 ;
        RECT 112.600 43.100 113.000 43.200 ;
        RECT 16.600 42.800 113.000 43.100 ;
        RECT 113.400 43.100 113.800 43.200 ;
        RECT 121.400 43.100 121.800 43.200 ;
        RECT 113.400 42.800 121.800 43.100 ;
        RECT 150.200 43.100 150.600 43.200 ;
        RECT 151.800 43.100 152.200 43.200 ;
        RECT 150.200 42.800 152.200 43.100 ;
        RECT 153.400 42.800 153.800 43.200 ;
        RECT 6.200 42.100 6.600 42.200 ;
        RECT 21.400 42.100 21.800 42.200 ;
        RECT 6.200 41.800 21.800 42.100 ;
        RECT 29.400 42.100 29.800 42.200 ;
        RECT 59.000 42.100 59.400 42.200 ;
        RECT 29.400 41.800 59.400 42.100 ;
        RECT 59.800 42.100 60.200 42.200 ;
        RECT 62.200 42.100 62.600 42.200 ;
        RECT 59.800 41.800 62.600 42.100 ;
        RECT 80.600 42.100 81.000 42.200 ;
        RECT 98.200 42.100 98.600 42.200 ;
        RECT 80.600 41.800 98.600 42.100 ;
        RECT 110.200 42.100 110.600 42.200 ;
        RECT 148.600 42.100 149.000 42.200 ;
        RECT 110.200 41.800 149.000 42.100 ;
        RECT 150.200 42.100 150.600 42.200 ;
        RECT 157.400 42.100 157.800 42.200 ;
        RECT 150.200 41.800 157.800 42.100 ;
        RECT 69.400 41.100 69.800 41.200 ;
        RECT 87.000 41.100 87.400 41.200 ;
        RECT 69.400 40.800 87.400 41.100 ;
        RECT 148.600 41.100 148.900 41.800 ;
        RECT 195.800 41.100 196.200 41.200 ;
        RECT 215.800 41.100 216.200 41.200 ;
        RECT 148.600 40.800 216.200 41.100 ;
        RECT 76.600 40.100 77.000 40.200 ;
        RECT 83.800 40.100 84.200 40.200 ;
        RECT 76.600 39.800 84.200 40.100 ;
        RECT 85.400 40.100 85.800 40.200 ;
        RECT 115.000 40.100 115.400 40.200 ;
        RECT 85.400 39.800 115.400 40.100 ;
        RECT 155.000 40.100 155.400 40.200 ;
        RECT 168.600 40.100 169.000 40.200 ;
        RECT 155.000 39.800 169.000 40.100 ;
        RECT 40.600 39.100 41.000 39.200 ;
        RECT 83.000 39.100 83.400 39.200 ;
        RECT 40.600 38.800 83.400 39.100 ;
        RECT 98.200 39.100 98.600 39.200 ;
        RECT 104.600 39.100 105.000 39.200 ;
        RECT 111.000 39.100 111.400 39.200 ;
        RECT 98.200 38.800 111.400 39.100 ;
        RECT 116.600 39.100 117.000 39.200 ;
        RECT 152.600 39.100 153.000 39.200 ;
        RECT 116.600 38.800 136.900 39.100 ;
        RECT 152.600 38.800 184.100 39.100 ;
        RECT 47.000 38.100 47.400 38.200 ;
        RECT 59.800 38.100 60.200 38.200 ;
        RECT 64.600 38.100 65.000 38.200 ;
        RECT 47.000 37.800 65.000 38.100 ;
        RECT 103.000 37.800 103.400 38.200 ;
        RECT 110.200 38.100 110.600 38.200 ;
        RECT 136.600 38.100 136.900 38.800 ;
        RECT 183.800 38.200 184.100 38.800 ;
        RECT 160.600 38.100 161.000 38.200 ;
        RECT 110.200 37.800 135.300 38.100 ;
        RECT 136.600 37.800 161.000 38.100 ;
        RECT 163.800 37.800 164.200 38.200 ;
        RECT 164.600 37.800 165.000 38.200 ;
        RECT 183.800 37.800 184.200 38.200 ;
        RECT 42.200 37.100 42.600 37.200 ;
        RECT 44.600 37.100 45.000 37.200 ;
        RECT 42.200 36.800 45.000 37.100 ;
        RECT 61.400 36.800 61.800 37.200 ;
        RECT 72.600 37.100 73.000 37.200 ;
        RECT 73.400 37.100 73.800 37.200 ;
        RECT 72.600 36.800 73.800 37.100 ;
        RECT 95.800 37.100 96.200 37.200 ;
        RECT 103.000 37.100 103.300 37.800 ;
        RECT 135.000 37.200 135.300 37.800 ;
        RECT 163.800 37.200 164.100 37.800 ;
        RECT 164.600 37.200 164.900 37.800 ;
        RECT 95.800 36.800 103.300 37.100 ;
        RECT 103.800 36.800 104.200 37.200 ;
        RECT 110.200 37.100 110.600 37.200 ;
        RECT 113.400 37.100 113.800 37.200 ;
        RECT 110.200 36.800 113.800 37.100 ;
        RECT 124.600 37.100 125.000 37.200 ;
        RECT 130.200 37.100 130.600 37.200 ;
        RECT 124.600 36.800 130.600 37.100 ;
        RECT 135.000 37.100 135.400 37.200 ;
        RECT 141.400 37.100 141.800 37.200 ;
        RECT 135.000 36.800 141.800 37.100 ;
        RECT 143.000 37.100 143.400 37.200 ;
        RECT 154.200 37.100 154.600 37.200 ;
        RECT 143.000 36.800 154.600 37.100 ;
        RECT 161.400 36.800 161.800 37.200 ;
        RECT 163.800 36.800 164.200 37.200 ;
        RECT 164.600 36.800 165.000 37.200 ;
        RECT 167.000 37.100 167.400 37.200 ;
        RECT 167.800 37.100 168.200 37.200 ;
        RECT 167.000 36.800 168.200 37.100 ;
        RECT 173.400 37.100 173.800 37.200 ;
        RECT 180.600 37.100 181.000 37.200 ;
        RECT 173.400 36.800 181.000 37.100 ;
        RECT 199.000 37.100 199.400 37.200 ;
        RECT 201.400 37.100 201.800 37.200 ;
        RECT 199.000 36.800 201.800 37.100 ;
        RECT 203.000 36.800 203.400 37.200 ;
        RECT 61.400 36.200 61.700 36.800 ;
        RECT 103.800 36.200 104.100 36.800 ;
        RECT 161.400 36.200 161.700 36.800 ;
        RECT 203.000 36.200 203.300 36.800 ;
        RECT 1.400 36.100 1.800 36.200 ;
        RECT 2.200 36.100 2.600 36.200 ;
        RECT 1.400 35.800 2.600 36.100 ;
        RECT 18.200 36.100 18.600 36.200 ;
        RECT 51.000 36.100 51.400 36.200 ;
        RECT 18.200 35.800 51.400 36.100 ;
        RECT 61.400 35.800 61.800 36.200 ;
        RECT 62.200 36.100 62.600 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 90.200 36.100 90.600 36.200 ;
        RECT 62.200 35.800 90.600 36.100 ;
        RECT 101.400 36.100 101.800 36.200 ;
        RECT 103.800 36.100 104.200 36.200 ;
        RECT 101.400 35.800 104.200 36.100 ;
        RECT 104.600 36.100 105.000 36.200 ;
        RECT 107.000 36.100 107.400 36.200 ;
        RECT 116.600 36.100 117.000 36.200 ;
        RECT 104.600 35.800 117.000 36.100 ;
        RECT 117.400 36.100 117.800 36.200 ;
        RECT 118.200 36.100 118.600 36.200 ;
        RECT 125.400 36.100 125.800 36.200 ;
        RECT 130.200 36.100 130.600 36.200 ;
        RECT 139.800 36.100 140.200 36.200 ;
        RECT 147.800 36.100 148.200 36.200 ;
        RECT 117.400 35.800 130.600 36.100 ;
        RECT 139.000 35.800 148.200 36.100 ;
        RECT 159.800 36.100 160.200 36.200 ;
        RECT 161.400 36.100 161.800 36.200 ;
        RECT 174.200 36.100 174.600 36.200 ;
        RECT 177.400 36.100 177.800 36.200 ;
        RECT 159.800 35.800 177.800 36.100 ;
        RECT 191.000 35.800 191.400 36.200 ;
        RECT 198.200 35.800 198.600 36.200 ;
        RECT 200.600 36.100 201.000 36.200 ;
        RECT 203.000 36.100 203.400 36.200 ;
        RECT 200.600 35.800 203.400 36.100 ;
        RECT 215.800 36.100 216.200 36.200 ;
        RECT 217.400 36.100 217.800 36.200 ;
        RECT 226.200 36.100 226.600 36.200 ;
        RECT 215.800 35.800 226.600 36.100 ;
        RECT 51.000 35.200 51.300 35.800 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 6.200 35.100 6.600 35.200 ;
        RECT 7.800 35.100 8.200 35.200 ;
        RECT 6.200 34.800 8.200 35.100 ;
        RECT 13.400 35.100 13.800 35.200 ;
        RECT 28.600 35.100 29.000 35.200 ;
        RECT 32.600 35.100 33.000 35.200 ;
        RECT 13.400 34.800 33.000 35.100 ;
        RECT 47.000 35.100 47.400 35.200 ;
        RECT 49.400 35.100 49.800 35.200 ;
        RECT 50.200 35.100 50.600 35.200 ;
        RECT 47.000 34.800 50.600 35.100 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 52.600 35.100 53.000 35.200 ;
        RECT 56.600 35.100 57.000 35.200 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 52.600 34.800 59.400 35.100 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 63.800 35.100 64.200 35.200 ;
        RECT 79.000 35.100 79.400 35.200 ;
        RECT 80.600 35.100 81.000 35.200 ;
        RECT 60.600 34.800 81.000 35.100 ;
        RECT 82.200 35.100 82.600 35.200 ;
        RECT 86.200 35.100 86.600 35.200 ;
        RECT 82.200 34.800 86.600 35.100 ;
        RECT 89.400 35.100 89.800 35.200 ;
        RECT 99.000 35.100 99.400 35.200 ;
        RECT 89.400 34.800 99.400 35.100 ;
        RECT 103.000 34.800 103.400 35.200 ;
        RECT 108.600 35.100 109.000 35.200 ;
        RECT 111.000 35.100 111.400 35.200 ;
        RECT 108.600 34.800 111.400 35.100 ;
        RECT 113.400 35.100 113.800 35.200 ;
        RECT 115.000 35.100 115.400 35.200 ;
        RECT 113.400 34.800 115.400 35.100 ;
        RECT 128.600 35.100 129.000 35.200 ;
        RECT 136.600 35.100 137.000 35.200 ;
        RECT 139.800 35.100 140.200 35.200 ;
        RECT 166.200 35.100 166.600 35.200 ;
        RECT 128.600 34.800 131.300 35.100 ;
        RECT 136.600 34.800 166.600 35.100 ;
        RECT 171.000 35.100 171.400 35.200 ;
        RECT 178.200 35.100 178.600 35.200 ;
        RECT 171.000 34.800 178.600 35.100 ;
        RECT 191.000 35.100 191.300 35.800 ;
        RECT 198.200 35.100 198.500 35.800 ;
        RECT 191.000 34.800 198.500 35.100 ;
        RECT 199.800 34.800 200.200 35.200 ;
        RECT 215.000 35.100 215.400 35.200 ;
        RECT 216.600 35.100 217.000 35.200 ;
        RECT 215.000 34.800 217.000 35.100 ;
        RECT 218.200 35.100 218.600 35.200 ;
        RECT 218.200 34.800 226.500 35.100 ;
        RECT 3.800 34.100 4.100 34.800 ;
        RECT 103.000 34.200 103.300 34.800 ;
        RECT 131.000 34.200 131.300 34.800 ;
        RECT 14.200 34.100 14.600 34.200 ;
        RECT 3.800 33.800 14.600 34.100 ;
        RECT 23.800 34.100 24.200 34.200 ;
        RECT 26.200 34.100 26.600 34.200 ;
        RECT 23.800 33.800 26.600 34.100 ;
        RECT 29.400 34.100 29.800 34.200 ;
        RECT 30.200 34.100 30.600 34.200 ;
        RECT 29.400 33.800 30.600 34.100 ;
        RECT 37.400 34.100 37.800 34.200 ;
        RECT 47.000 34.100 47.400 34.200 ;
        RECT 37.400 33.800 47.400 34.100 ;
        RECT 51.800 34.100 52.200 34.200 ;
        RECT 56.600 34.100 57.000 34.200 ;
        RECT 51.800 33.800 57.000 34.100 ;
        RECT 58.200 34.100 58.600 34.200 ;
        RECT 71.000 34.100 71.400 34.200 ;
        RECT 87.000 34.100 87.400 34.200 ;
        RECT 58.200 33.800 87.400 34.100 ;
        RECT 103.000 33.800 103.400 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 104.600 33.800 116.200 34.100 ;
        RECT 120.600 34.100 121.000 34.200 ;
        RECT 125.400 34.100 125.800 34.200 ;
        RECT 120.600 33.800 125.800 34.100 ;
        RECT 131.000 33.800 131.400 34.200 ;
        RECT 134.200 34.100 134.600 34.200 ;
        RECT 145.400 34.100 145.800 34.200 ;
        RECT 134.200 33.800 145.800 34.100 ;
        RECT 151.000 34.100 151.400 34.200 ;
        RECT 152.600 34.100 153.000 34.200 ;
        RECT 151.000 33.800 153.000 34.100 ;
        RECT 161.400 34.100 161.800 34.200 ;
        RECT 171.000 34.100 171.400 34.200 ;
        RECT 161.400 33.800 171.400 34.100 ;
        RECT 190.200 34.100 190.600 34.200 ;
        RECT 199.800 34.100 200.100 34.800 ;
        RECT 215.000 34.100 215.300 34.800 ;
        RECT 190.200 33.800 215.300 34.100 ;
        RECT 226.200 34.200 226.500 34.800 ;
        RECT 226.200 33.800 226.600 34.200 ;
        RECT 19.000 33.100 19.400 33.200 ;
        RECT 27.000 33.100 27.400 33.200 ;
        RECT 19.000 32.800 27.400 33.100 ;
        RECT 50.200 33.100 50.600 33.200 ;
        RECT 61.400 33.100 61.800 33.200 ;
        RECT 50.200 32.800 61.800 33.100 ;
        RECT 63.000 33.100 63.400 33.200 ;
        RECT 71.800 33.100 72.200 33.200 ;
        RECT 63.000 32.800 72.200 33.100 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 75.000 32.800 76.200 33.100 ;
        RECT 76.600 33.100 77.000 33.200 ;
        RECT 100.600 33.100 101.000 33.200 ;
        RECT 76.600 32.800 101.000 33.100 ;
        RECT 133.400 33.100 133.800 33.200 ;
        RECT 146.200 33.100 146.600 33.200 ;
        RECT 133.400 32.800 146.600 33.100 ;
        RECT 159.000 33.100 159.400 33.200 ;
        RECT 163.000 33.100 163.400 33.200 ;
        RECT 159.000 32.800 163.400 33.100 ;
        RECT 171.800 33.100 172.200 33.200 ;
        RECT 178.200 33.100 178.600 33.200 ;
        RECT 196.600 33.100 197.000 33.200 ;
        RECT 171.800 32.800 197.000 33.100 ;
        RECT 202.200 32.800 202.600 33.200 ;
        RECT 219.800 33.100 220.200 33.200 ;
        RECT 220.600 33.100 221.000 33.200 ;
        RECT 219.800 32.800 221.000 33.100 ;
        RECT 225.400 33.100 225.800 33.200 ;
        RECT 230.200 33.100 230.600 33.200 ;
        RECT 225.400 32.800 230.600 33.100 ;
        RECT 15.000 32.100 15.400 32.200 ;
        RECT 29.400 32.100 29.800 32.200 ;
        RECT 15.000 31.800 29.800 32.100 ;
        RECT 80.600 32.100 81.000 32.200 ;
        RECT 91.000 32.100 91.400 32.200 ;
        RECT 80.600 31.800 91.400 32.100 ;
        RECT 97.400 32.100 97.800 32.200 ;
        RECT 107.000 32.100 107.400 32.200 ;
        RECT 97.400 31.800 107.400 32.100 ;
        RECT 111.000 32.100 111.400 32.200 ;
        RECT 115.800 32.100 116.200 32.200 ;
        RECT 111.000 31.800 116.200 32.100 ;
        RECT 163.000 32.100 163.300 32.800 ;
        RECT 167.800 32.100 168.200 32.200 ;
        RECT 163.000 31.800 168.200 32.100 ;
        RECT 169.400 32.100 169.800 32.200 ;
        RECT 173.400 32.100 173.800 32.200 ;
        RECT 177.400 32.100 177.800 32.200 ;
        RECT 169.400 31.800 177.800 32.100 ;
        RECT 183.000 32.100 183.400 32.200 ;
        RECT 186.200 32.100 186.600 32.200 ;
        RECT 199.800 32.100 200.200 32.200 ;
        RECT 183.000 31.800 200.200 32.100 ;
        RECT 202.200 32.100 202.500 32.800 ;
        RECT 227.000 32.100 227.400 32.200 ;
        RECT 202.200 31.800 227.400 32.100 ;
        RECT 7.000 31.100 7.400 31.200 ;
        RECT 17.400 31.100 17.800 31.200 ;
        RECT 7.000 30.800 17.800 31.100 ;
        RECT 28.600 31.100 29.000 31.200 ;
        RECT 76.600 31.100 77.000 31.200 ;
        RECT 28.600 30.800 77.000 31.100 ;
        RECT 91.000 31.100 91.400 31.200 ;
        RECT 97.400 31.100 97.800 31.200 ;
        RECT 143.000 31.100 143.400 31.200 ;
        RECT 91.000 30.800 143.400 31.100 ;
        RECT 148.600 31.100 149.000 31.200 ;
        RECT 163.000 31.100 163.400 31.200 ;
        RECT 165.400 31.100 165.800 31.200 ;
        RECT 148.600 30.800 165.800 31.100 ;
        RECT 168.600 31.100 169.000 31.200 ;
        RECT 172.600 31.100 173.000 31.200 ;
        RECT 168.600 30.800 173.000 31.100 ;
        RECT 175.800 31.100 176.200 31.200 ;
        RECT 181.400 31.100 181.800 31.200 ;
        RECT 175.800 30.800 181.800 31.100 ;
        RECT 193.400 31.100 193.800 31.200 ;
        RECT 202.200 31.100 202.600 31.200 ;
        RECT 193.400 30.800 202.600 31.100 ;
        RECT 204.600 31.100 205.000 31.200 ;
        RECT 221.400 31.100 221.800 31.200 ;
        RECT 204.600 30.800 221.800 31.100 ;
        RECT 61.400 30.100 61.800 30.200 ;
        RECT 83.800 30.100 84.200 30.200 ;
        RECT 61.400 29.800 84.200 30.100 ;
        RECT 99.800 30.100 100.200 30.200 ;
        RECT 102.200 30.100 102.600 30.200 ;
        RECT 99.800 29.800 102.600 30.100 ;
        RECT 114.200 30.100 114.600 30.200 ;
        RECT 117.400 30.100 117.800 30.200 ;
        RECT 127.000 30.100 127.400 30.200 ;
        RECT 142.200 30.100 142.600 30.200 ;
        RECT 114.200 29.800 116.900 30.100 ;
        RECT 117.400 29.800 142.600 30.100 ;
        RECT 155.800 30.100 156.200 30.200 ;
        RECT 157.400 30.100 157.800 30.200 ;
        RECT 160.600 30.100 161.000 30.200 ;
        RECT 155.800 29.800 161.000 30.100 ;
        RECT 161.400 29.800 161.800 30.200 ;
        RECT 196.600 30.100 197.000 30.200 ;
        RECT 203.800 30.100 204.200 30.200 ;
        RECT 211.000 30.100 211.400 30.200 ;
        RECT 196.600 29.800 211.400 30.100 ;
        RECT 10.200 29.100 10.600 29.200 ;
        RECT 12.600 29.100 13.000 29.200 ;
        RECT 10.200 28.800 13.000 29.100 ;
        RECT 31.800 29.100 32.200 29.200 ;
        RECT 39.800 29.100 40.200 29.200 ;
        RECT 51.800 29.100 52.200 29.200 ;
        RECT 31.800 28.800 52.200 29.100 ;
        RECT 70.200 29.100 70.600 29.200 ;
        RECT 79.000 29.100 79.400 29.200 ;
        RECT 70.200 28.800 79.400 29.100 ;
        RECT 101.400 29.100 101.800 29.200 ;
        RECT 102.200 29.100 102.600 29.200 ;
        RECT 101.400 28.800 102.600 29.100 ;
        RECT 106.200 29.100 106.600 29.200 ;
        RECT 114.200 29.100 114.600 29.200 ;
        RECT 106.200 28.800 114.600 29.100 ;
        RECT 116.600 29.100 116.900 29.800 ;
        RECT 161.400 29.200 161.700 29.800 ;
        RECT 121.400 29.100 121.800 29.200 ;
        RECT 116.600 28.800 121.800 29.100 ;
        RECT 129.400 29.100 129.800 29.200 ;
        RECT 143.800 29.100 144.200 29.200 ;
        RECT 148.600 29.100 149.000 29.200 ;
        RECT 129.400 28.800 149.000 29.100 ;
        RECT 161.400 28.800 161.800 29.200 ;
        RECT 185.400 29.100 185.800 29.200 ;
        RECT 185.400 28.800 209.700 29.100 ;
        RECT 209.400 28.200 209.700 28.800 ;
        RECT 11.800 27.800 12.200 28.200 ;
        RECT 21.400 27.800 21.800 28.200 ;
        RECT 23.800 28.100 24.200 28.200 ;
        RECT 31.000 28.100 31.400 28.200 ;
        RECT 23.800 27.800 31.400 28.100 ;
        RECT 95.800 27.800 96.200 28.200 ;
        RECT 139.800 28.100 140.200 28.200 ;
        RECT 143.000 28.100 143.400 28.200 ;
        RECT 162.200 28.100 162.600 28.200 ;
        RECT 139.800 27.800 162.600 28.100 ;
        RECT 163.000 28.100 163.400 28.200 ;
        RECT 187.800 28.100 188.200 28.200 ;
        RECT 163.000 27.800 188.200 28.100 ;
        RECT 209.400 27.800 209.800 28.200 ;
        RECT 3.800 27.100 4.200 27.200 ;
        RECT 4.600 27.100 5.000 27.200 ;
        RECT 3.800 26.800 5.000 27.100 ;
        RECT 11.800 27.100 12.100 27.800 ;
        RECT 21.400 27.100 21.700 27.800 ;
        RECT 30.200 27.100 30.600 27.200 ;
        RECT 33.400 27.100 33.800 27.200 ;
        RECT 42.200 27.100 42.600 27.200 ;
        RECT 11.800 26.800 42.600 27.100 ;
        RECT 45.400 27.100 45.800 27.200 ;
        RECT 51.000 27.100 51.400 27.200 ;
        RECT 45.400 26.800 51.400 27.100 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 81.400 27.100 81.800 27.200 ;
        RECT 75.800 26.800 81.800 27.100 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 95.800 27.100 96.100 27.800 ;
        RECT 94.200 26.800 96.100 27.100 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 151.000 27.100 151.400 27.200 ;
        RECT 125.400 26.800 151.400 27.100 ;
        RECT 152.600 27.100 153.000 27.200 ;
        RECT 161.400 27.100 161.800 27.200 ;
        RECT 152.600 26.800 161.800 27.100 ;
        RECT 166.200 27.100 166.600 27.200 ;
        RECT 167.000 27.100 167.400 27.200 ;
        RECT 196.600 27.100 197.000 27.200 ;
        RECT 166.200 26.800 197.000 27.100 ;
        RECT 200.600 26.800 201.000 27.200 ;
        RECT 206.200 27.100 206.600 27.200 ;
        RECT 215.000 27.100 215.400 27.200 ;
        RECT 206.200 26.800 215.400 27.100 ;
        RECT 215.800 27.100 216.200 27.200 ;
        RECT 224.600 27.100 225.000 27.200 ;
        RECT 215.800 26.800 225.000 27.100 ;
        RECT 228.600 27.100 229.000 27.200 ;
        RECT 229.400 27.100 229.800 27.200 ;
        RECT 228.600 26.800 229.800 27.100 ;
        RECT 3.000 26.100 3.400 26.200 ;
        RECT 23.000 26.100 23.400 26.200 ;
        RECT 26.200 26.100 26.600 26.200 ;
        RECT 3.000 25.800 26.600 26.100 ;
        RECT 48.600 25.800 49.000 26.200 ;
        RECT 50.200 26.100 50.600 26.200 ;
        RECT 53.400 26.100 53.800 26.200 ;
        RECT 50.200 25.800 53.800 26.100 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 90.200 26.100 90.600 26.200 ;
        RECT 72.600 25.800 90.600 26.100 ;
        RECT 104.600 26.100 104.900 26.800 ;
        RECT 108.600 26.100 108.900 26.800 ;
        RECT 200.600 26.200 200.900 26.800 ;
        RECT 104.600 25.800 108.900 26.100 ;
        RECT 145.400 26.100 145.800 26.200 ;
        RECT 147.000 26.100 147.400 26.200 ;
        RECT 197.400 26.100 197.800 26.200 ;
        RECT 198.200 26.100 198.600 26.200 ;
        RECT 145.400 25.800 198.600 26.100 ;
        RECT 200.600 25.800 201.000 26.200 ;
        RECT 203.800 26.100 204.200 26.200 ;
        RECT 204.600 26.100 205.000 26.200 ;
        RECT 207.000 26.100 207.400 26.200 ;
        RECT 203.800 25.800 207.400 26.100 ;
        RECT 219.000 25.800 219.400 26.200 ;
        RECT 220.600 26.100 221.000 26.200 ;
        RECT 225.400 26.100 225.800 26.200 ;
        RECT 220.600 25.800 225.800 26.100 ;
        RECT 48.600 25.200 48.900 25.800 ;
        RECT 219.000 25.200 219.300 25.800 ;
        RECT 9.400 25.100 9.800 25.200 ;
        RECT 2.200 24.800 9.800 25.100 ;
        RECT 27.000 25.100 27.400 25.200 ;
        RECT 28.600 25.100 29.000 25.200 ;
        RECT 27.000 24.800 29.000 25.100 ;
        RECT 48.600 24.800 49.000 25.200 ;
        RECT 51.800 25.100 52.200 25.200 ;
        RECT 57.400 25.100 57.800 25.200 ;
        RECT 51.800 24.800 57.800 25.100 ;
        RECT 81.400 25.100 81.800 25.200 ;
        RECT 84.600 25.100 85.000 25.200 ;
        RECT 110.200 25.100 110.600 25.200 ;
        RECT 81.400 24.800 110.600 25.100 ;
        RECT 111.800 25.100 112.200 25.200 ;
        RECT 134.200 25.100 134.600 25.200 ;
        RECT 155.000 25.100 155.400 25.200 ;
        RECT 111.800 24.800 134.600 25.100 ;
        RECT 147.800 24.800 155.400 25.100 ;
        RECT 160.600 25.100 161.000 25.200 ;
        RECT 161.400 25.100 161.800 25.200 ;
        RECT 160.600 24.800 161.800 25.100 ;
        RECT 164.600 25.100 165.000 25.200 ;
        RECT 191.000 25.100 191.400 25.200 ;
        RECT 164.600 24.800 191.400 25.100 ;
        RECT 219.000 24.800 219.400 25.200 ;
        RECT 2.200 24.200 2.500 24.800 ;
        RECT 147.800 24.200 148.100 24.800 ;
        RECT 2.200 23.800 2.600 24.200 ;
        RECT 55.800 24.100 56.200 24.200 ;
        RECT 58.200 24.100 58.600 24.200 ;
        RECT 67.000 24.100 67.400 24.200 ;
        RECT 72.600 24.100 73.000 24.200 ;
        RECT 55.800 23.800 73.000 24.100 ;
        RECT 78.200 24.100 78.600 24.200 ;
        RECT 83.000 24.100 83.400 24.200 ;
        RECT 78.200 23.800 83.400 24.100 ;
        RECT 90.200 24.100 90.600 24.200 ;
        RECT 121.400 24.100 121.800 24.200 ;
        RECT 145.400 24.100 145.800 24.200 ;
        RECT 90.200 23.800 145.800 24.100 ;
        RECT 147.800 23.800 148.200 24.200 ;
        RECT 148.600 24.100 149.000 24.200 ;
        RECT 159.000 24.100 159.400 24.200 ;
        RECT 148.600 23.800 159.400 24.100 ;
        RECT 167.800 24.100 168.200 24.200 ;
        RECT 179.000 24.100 179.400 24.200 ;
        RECT 167.800 23.800 179.400 24.100 ;
        RECT 184.600 24.100 185.000 24.200 ;
        RECT 203.800 24.100 204.200 24.200 ;
        RECT 184.600 23.800 204.200 24.100 ;
        RECT 68.600 23.100 69.000 23.200 ;
        RECT 131.000 23.100 131.400 23.200 ;
        RECT 68.600 22.800 131.400 23.100 ;
        RECT 140.600 22.800 141.000 23.200 ;
        RECT 142.200 23.100 142.600 23.200 ;
        RECT 147.800 23.100 148.200 23.200 ;
        RECT 193.400 23.100 193.800 23.200 ;
        RECT 142.200 22.800 193.800 23.100 ;
        RECT 47.000 22.100 47.400 22.200 ;
        RECT 60.600 22.100 61.000 22.200 ;
        RECT 47.000 21.800 61.000 22.100 ;
        RECT 81.400 22.100 81.800 22.200 ;
        RECT 99.800 22.100 100.200 22.200 ;
        RECT 81.400 21.800 100.200 22.100 ;
        RECT 118.200 22.100 118.600 22.200 ;
        RECT 119.800 22.100 120.200 22.200 ;
        RECT 118.200 21.800 120.200 22.100 ;
        RECT 123.800 22.100 124.200 22.200 ;
        RECT 134.200 22.100 134.600 22.200 ;
        RECT 123.800 21.800 134.600 22.100 ;
        RECT 137.400 22.100 137.800 22.200 ;
        RECT 140.600 22.100 140.900 22.800 ;
        RECT 149.400 22.100 149.800 22.200 ;
        RECT 153.400 22.100 153.800 22.200 ;
        RECT 160.600 22.100 161.000 22.200 ;
        RECT 171.000 22.100 171.400 22.200 ;
        RECT 137.400 21.800 171.400 22.100 ;
        RECT 224.600 22.100 225.000 22.200 ;
        RECT 228.600 22.100 229.000 22.200 ;
        RECT 224.600 21.800 229.000 22.100 ;
        RECT 79.800 21.100 80.200 21.200 ;
        RECT 97.400 21.100 97.800 21.200 ;
        RECT 79.800 20.800 97.800 21.100 ;
        RECT 99.800 21.100 100.200 21.200 ;
        RECT 117.400 21.100 117.800 21.200 ;
        RECT 99.800 20.800 117.800 21.100 ;
        RECT 109.400 19.800 109.800 20.200 ;
        RECT 141.400 20.100 141.800 20.200 ;
        RECT 201.400 20.100 201.800 20.200 ;
        RECT 141.400 19.800 201.800 20.100 ;
        RECT 10.200 19.100 10.600 19.200 ;
        RECT 23.000 19.100 23.400 19.200 ;
        RECT 10.200 18.800 23.400 19.100 ;
        RECT 23.800 19.100 24.200 19.200 ;
        RECT 36.600 19.100 37.000 19.200 ;
        RECT 43.800 19.100 44.200 19.200 ;
        RECT 23.800 18.800 44.200 19.100 ;
        RECT 54.200 19.100 54.600 19.200 ;
        RECT 55.000 19.100 55.400 19.200 ;
        RECT 54.200 18.800 55.400 19.100 ;
        RECT 79.000 19.100 79.400 19.200 ;
        RECT 102.200 19.100 102.600 19.200 ;
        RECT 79.000 18.800 102.600 19.100 ;
        RECT 109.400 19.100 109.700 19.800 ;
        RECT 115.000 19.100 115.400 19.200 ;
        RECT 126.200 19.100 126.600 19.200 ;
        RECT 148.600 19.100 149.000 19.200 ;
        RECT 109.400 18.800 126.600 19.100 ;
        RECT 127.800 18.800 149.000 19.100 ;
        RECT 186.200 19.100 186.600 19.200 ;
        RECT 187.000 19.100 187.400 19.200 ;
        RECT 186.200 18.800 187.400 19.100 ;
        RECT 127.800 18.200 128.100 18.800 ;
        RECT 29.400 18.100 29.800 18.200 ;
        RECT 63.800 18.100 64.200 18.200 ;
        RECT 77.400 18.100 77.800 18.200 ;
        RECT 82.200 18.100 82.600 18.200 ;
        RECT 90.200 18.100 90.600 18.200 ;
        RECT 29.400 17.800 90.600 18.100 ;
        RECT 108.600 18.100 109.000 18.200 ;
        RECT 126.200 18.100 126.600 18.200 ;
        RECT 108.600 17.800 126.600 18.100 ;
        RECT 127.800 17.800 128.200 18.200 ;
        RECT 11.000 17.100 11.400 17.200 ;
        RECT 49.400 17.100 49.800 17.200 ;
        RECT 11.000 16.800 49.800 17.100 ;
        RECT 83.000 17.100 83.400 17.200 ;
        RECT 85.400 17.100 85.800 17.200 ;
        RECT 103.800 17.100 104.200 17.200 ;
        RECT 83.000 16.800 104.200 17.100 ;
        RECT 111.000 16.800 111.400 17.200 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 161.400 17.100 161.800 17.200 ;
        RECT 168.600 17.100 169.000 17.200 ;
        RECT 161.400 16.800 169.000 17.100 ;
        RECT 172.600 17.100 173.000 17.200 ;
        RECT 177.400 17.100 177.800 17.200 ;
        RECT 172.600 16.800 177.800 17.100 ;
        RECT 11.800 16.100 12.200 16.200 ;
        RECT 14.200 16.100 14.600 16.200 ;
        RECT 11.800 15.800 14.600 16.100 ;
        RECT 21.400 16.100 21.800 16.200 ;
        RECT 29.400 16.100 29.800 16.200 ;
        RECT 21.400 15.800 29.800 16.100 ;
        RECT 35.000 16.100 35.400 16.200 ;
        RECT 39.800 16.100 40.200 16.200 ;
        RECT 35.000 15.800 40.200 16.100 ;
        RECT 43.000 15.800 43.400 16.200 ;
        RECT 64.600 16.100 65.000 16.200 ;
        RECT 67.000 16.100 67.400 16.200 ;
        RECT 64.600 15.800 67.400 16.100 ;
        RECT 67.800 16.100 68.200 16.200 ;
        RECT 71.800 16.100 72.200 16.200 ;
        RECT 67.800 15.800 72.200 16.100 ;
        RECT 92.600 15.800 93.000 16.200 ;
        RECT 103.800 16.100 104.200 16.200 ;
        RECT 111.000 16.100 111.300 16.800 ;
        RECT 126.200 16.200 126.500 16.800 ;
        RECT 103.800 15.800 111.300 16.100 ;
        RECT 115.000 16.100 115.400 16.200 ;
        RECT 115.800 16.100 116.200 16.200 ;
        RECT 115.000 15.800 116.200 16.100 ;
        RECT 116.600 16.100 117.000 16.200 ;
        RECT 120.600 16.100 121.000 16.200 ;
        RECT 116.600 15.800 121.000 16.100 ;
        RECT 121.400 16.100 121.800 16.200 ;
        RECT 123.000 16.100 123.400 16.200 ;
        RECT 121.400 15.800 123.400 16.100 ;
        RECT 126.200 15.800 126.600 16.200 ;
        RECT 135.800 16.100 136.200 16.200 ;
        RECT 141.400 16.100 141.800 16.200 ;
        RECT 135.800 15.800 141.800 16.100 ;
        RECT 142.200 16.100 142.600 16.200 ;
        RECT 170.200 16.100 170.600 16.200 ;
        RECT 172.600 16.100 173.000 16.200 ;
        RECT 142.200 15.800 173.000 16.100 ;
        RECT 187.000 16.100 187.400 16.200 ;
        RECT 189.400 16.100 189.800 16.200 ;
        RECT 187.000 15.800 189.800 16.100 ;
        RECT 225.400 16.100 225.800 16.200 ;
        RECT 226.200 16.100 226.600 16.200 ;
        RECT 228.600 16.100 229.000 16.200 ;
        RECT 225.400 15.800 229.000 16.100 ;
        RECT 43.000 15.200 43.300 15.800 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 35.000 15.100 35.400 15.200 ;
        RECT 29.400 14.800 35.400 15.100 ;
        RECT 43.000 14.800 43.400 15.200 ;
        RECT 58.200 15.100 58.600 15.200 ;
        RECT 59.800 15.100 60.200 15.200 ;
        RECT 83.000 15.100 83.400 15.200 ;
        RECT 58.200 14.800 83.400 15.100 ;
        RECT 85.400 15.100 85.800 15.200 ;
        RECT 92.600 15.100 92.900 15.800 ;
        RECT 85.400 14.800 92.900 15.100 ;
        RECT 110.200 15.100 110.600 15.200 ;
        RECT 113.400 15.100 113.800 15.200 ;
        RECT 138.200 15.100 138.600 15.200 ;
        RECT 141.400 15.100 141.800 15.200 ;
        RECT 110.200 14.800 141.800 15.100 ;
        RECT 162.200 15.100 162.600 15.200 ;
        RECT 211.800 15.100 212.200 15.200 ;
        RECT 215.000 15.100 215.400 15.200 ;
        RECT 162.200 14.800 215.400 15.100 ;
        RECT 12.600 14.100 12.900 14.800 ;
        RECT 15.800 14.100 16.200 14.200 ;
        RECT 12.600 13.800 16.200 14.100 ;
        RECT 46.200 14.100 46.600 14.200 ;
        RECT 55.800 14.100 56.200 14.200 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 77.400 14.100 77.800 14.200 ;
        RECT 46.200 13.800 59.400 14.100 ;
        RECT 68.600 13.800 77.800 14.100 ;
        RECT 79.000 14.100 79.400 14.200 ;
        RECT 79.800 14.100 80.200 14.200 ;
        RECT 79.000 13.800 80.200 14.100 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 94.200 14.100 94.600 14.200 ;
        RECT 81.400 13.800 94.600 14.100 ;
        RECT 105.400 14.100 105.800 14.200 ;
        RECT 116.600 14.100 117.000 14.200 ;
        RECT 105.400 13.800 117.000 14.100 ;
        RECT 119.000 14.100 119.400 14.200 ;
        RECT 128.600 14.100 129.000 14.200 ;
        RECT 119.000 13.800 129.000 14.100 ;
        RECT 135.000 14.100 135.400 14.200 ;
        RECT 136.600 14.100 137.000 14.200 ;
        RECT 135.000 13.800 137.000 14.100 ;
        RECT 157.400 14.100 157.800 14.200 ;
        RECT 207.800 14.100 208.200 14.200 ;
        RECT 210.200 14.100 210.600 14.200 ;
        RECT 217.400 14.100 217.800 14.200 ;
        RECT 157.400 13.800 217.800 14.100 ;
        RECT 68.600 13.200 68.900 13.800 ;
        RECT 10.200 13.100 10.600 13.200 ;
        RECT 21.400 13.100 21.800 13.200 ;
        RECT 10.200 12.800 21.800 13.100 ;
        RECT 68.600 12.800 69.000 13.200 ;
        RECT 88.600 13.100 89.000 13.200 ;
        RECT 98.200 13.100 98.600 13.200 ;
        RECT 88.600 12.800 98.600 13.100 ;
        RECT 147.800 13.100 148.200 13.200 ;
        RECT 188.600 13.100 189.000 13.200 ;
        RECT 147.800 12.800 189.000 13.100 ;
        RECT 34.200 12.100 34.600 12.200 ;
        RECT 43.000 12.100 43.400 12.200 ;
        RECT 34.200 11.800 43.400 12.100 ;
        RECT 94.200 12.100 94.600 12.200 ;
        RECT 158.200 12.100 158.600 12.200 ;
        RECT 94.200 11.800 158.600 12.100 ;
        RECT 171.000 12.100 171.400 12.200 ;
        RECT 174.200 12.100 174.600 12.200 ;
        RECT 183.000 12.100 183.400 12.200 ;
        RECT 185.400 12.100 185.800 12.200 ;
        RECT 171.000 11.800 174.600 12.100 ;
        RECT 182.200 11.800 185.800 12.100 ;
        RECT 189.400 12.100 189.800 12.200 ;
        RECT 193.400 12.100 193.800 12.200 ;
        RECT 189.400 11.800 193.800 12.100 ;
        RECT 209.400 12.100 209.800 12.200 ;
        RECT 213.400 12.100 213.800 12.200 ;
        RECT 209.400 11.800 213.800 12.100 ;
        RECT 4.600 11.100 5.000 11.200 ;
        RECT 36.600 11.100 37.000 11.200 ;
        RECT 4.600 10.800 37.000 11.100 ;
        RECT 47.800 11.100 48.200 11.200 ;
        RECT 68.600 11.100 69.000 11.200 ;
        RECT 47.800 10.800 69.000 11.100 ;
        RECT 125.400 11.100 125.800 11.200 ;
        RECT 128.600 11.100 129.000 11.200 ;
        RECT 132.600 11.100 133.000 11.200 ;
        RECT 125.400 10.800 133.000 11.100 ;
        RECT 149.400 11.100 149.800 11.200 ;
        RECT 182.200 11.100 182.600 11.200 ;
        RECT 183.800 11.100 184.200 11.200 ;
        RECT 149.400 10.800 184.200 11.100 ;
        RECT 206.200 11.100 206.600 11.200 ;
        RECT 209.400 11.100 209.800 11.200 ;
        RECT 206.200 10.800 209.800 11.100 ;
        RECT 36.600 10.100 36.900 10.800 ;
        RECT 48.600 10.100 49.000 10.200 ;
        RECT 36.600 9.800 49.000 10.100 ;
        RECT 49.400 10.100 49.800 10.200 ;
        RECT 61.400 10.100 61.800 10.200 ;
        RECT 49.400 9.800 61.800 10.100 ;
        RECT 77.400 10.100 77.800 10.200 ;
        RECT 80.600 10.100 81.000 10.200 ;
        RECT 77.400 9.800 81.000 10.100 ;
        RECT 103.000 10.100 103.400 10.200 ;
        RECT 110.200 10.100 110.600 10.200 ;
        RECT 127.800 10.100 128.200 10.200 ;
        RECT 103.000 9.800 128.200 10.100 ;
        RECT 132.600 10.100 133.000 10.200 ;
        RECT 135.000 10.100 135.400 10.200 ;
        RECT 132.600 9.800 135.400 10.100 ;
        RECT 147.000 10.100 147.400 10.200 ;
        RECT 164.600 10.100 165.000 10.200 ;
        RECT 147.000 9.800 165.000 10.100 ;
        RECT 176.600 10.100 177.000 10.200 ;
        RECT 183.000 10.100 183.400 10.200 ;
        RECT 176.600 9.800 183.400 10.100 ;
        RECT 202.200 10.100 202.600 10.200 ;
        RECT 216.600 10.100 217.000 10.200 ;
        RECT 221.400 10.100 221.800 10.200 ;
        RECT 202.200 9.800 221.800 10.100 ;
        RECT 1.400 9.100 1.800 9.200 ;
        RECT 3.000 9.100 3.400 9.200 ;
        RECT 1.400 8.800 3.400 9.100 ;
        RECT 12.600 9.100 13.000 9.200 ;
        RECT 23.800 9.100 24.200 9.200 ;
        RECT 12.600 8.800 24.200 9.100 ;
        RECT 35.800 9.100 36.200 9.200 ;
        RECT 52.600 9.100 53.000 9.200 ;
        RECT 35.800 8.800 53.000 9.100 ;
        RECT 55.800 9.100 56.200 9.200 ;
        RECT 59.000 9.100 59.400 9.200 ;
        RECT 55.800 8.800 59.400 9.100 ;
        RECT 68.600 9.100 69.000 9.200 ;
        RECT 79.000 9.100 79.400 9.200 ;
        RECT 68.600 8.800 79.400 9.100 ;
        RECT 85.400 9.100 85.800 9.200 ;
        RECT 91.800 9.100 92.200 9.200 ;
        RECT 94.200 9.100 94.600 9.200 ;
        RECT 85.400 8.800 94.600 9.100 ;
        RECT 95.800 9.100 96.200 9.200 ;
        RECT 104.600 9.100 105.000 9.200 ;
        RECT 95.800 8.800 105.000 9.100 ;
        RECT 120.600 9.100 121.000 9.200 ;
        RECT 131.800 9.100 132.200 9.200 ;
        RECT 143.000 9.100 143.400 9.200 ;
        RECT 120.600 8.800 143.400 9.100 ;
        RECT 183.800 9.100 184.200 9.200 ;
        RECT 200.600 9.100 201.000 9.200 ;
        RECT 207.800 9.100 208.200 9.200 ;
        RECT 183.800 8.800 185.700 9.100 ;
        RECT 200.600 8.800 208.200 9.100 ;
        RECT 185.400 8.200 185.700 8.800 ;
        RECT 15.000 7.800 15.400 8.200 ;
        RECT 43.800 7.800 44.200 8.200 ;
        RECT 69.400 7.800 69.800 8.200 ;
        RECT 72.600 8.100 73.000 8.200 ;
        RECT 79.000 8.100 79.400 8.200 ;
        RECT 72.600 7.800 79.400 8.100 ;
        RECT 100.600 8.100 101.000 8.200 ;
        RECT 106.200 8.100 106.600 8.200 ;
        RECT 114.200 8.100 114.600 8.200 ;
        RECT 123.800 8.100 124.200 8.200 ;
        RECT 137.400 8.100 137.800 8.200 ;
        RECT 100.600 7.800 137.800 8.100 ;
        RECT 143.800 8.100 144.200 8.200 ;
        RECT 153.400 8.100 153.800 8.200 ;
        RECT 143.800 7.800 153.800 8.100 ;
        RECT 185.400 7.800 185.800 8.200 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 6.200 7.100 6.600 7.200 ;
        RECT 4.600 6.800 6.600 7.100 ;
        RECT 15.000 7.100 15.300 7.800 ;
        RECT 19.000 7.100 19.400 7.200 ;
        RECT 35.000 7.100 35.400 7.200 ;
        RECT 37.400 7.100 37.800 7.200 ;
        RECT 15.000 6.800 19.400 7.100 ;
        RECT 29.400 6.800 31.300 7.100 ;
        RECT 35.000 6.800 37.800 7.100 ;
        RECT 39.000 7.100 39.400 7.200 ;
        RECT 43.800 7.100 44.100 7.800 ;
        RECT 39.000 6.800 44.100 7.100 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 45.400 6.800 46.600 7.100 ;
        RECT 64.600 7.100 65.000 7.200 ;
        RECT 69.400 7.100 69.700 7.800 ;
        RECT 64.600 6.800 69.700 7.100 ;
        RECT 78.200 7.100 78.600 7.200 ;
        RECT 87.000 7.100 87.400 7.200 ;
        RECT 78.200 6.800 87.400 7.100 ;
        RECT 214.200 7.100 214.600 7.200 ;
        RECT 227.000 7.100 227.400 7.200 ;
        RECT 214.200 6.800 227.400 7.100 ;
        RECT 29.400 6.200 29.700 6.800 ;
        RECT 31.000 6.200 31.300 6.800 ;
        RECT 0.600 6.100 1.000 6.200 ;
        RECT 4.600 6.100 5.000 6.200 ;
        RECT 0.600 5.800 5.000 6.100 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 37.400 6.100 37.800 6.200 ;
        RECT 41.400 6.100 41.800 6.200 ;
        RECT 85.400 6.100 85.800 6.200 ;
        RECT 37.400 5.800 85.800 6.100 ;
        RECT 93.400 6.100 93.800 6.200 ;
        RECT 115.000 6.100 115.400 6.200 ;
        RECT 129.400 6.100 129.800 6.200 ;
        RECT 93.400 5.800 99.300 6.100 ;
        RECT 115.000 5.800 129.800 6.100 ;
        RECT 131.000 6.100 131.400 6.200 ;
        RECT 155.000 6.100 155.400 6.200 ;
        RECT 156.600 6.100 157.000 6.200 ;
        RECT 131.000 5.800 157.000 6.100 ;
        RECT 161.400 6.100 161.800 6.200 ;
        RECT 169.400 6.100 169.800 6.200 ;
        RECT 161.400 5.800 169.800 6.100 ;
        RECT 198.200 6.100 198.600 6.200 ;
        RECT 204.600 6.100 205.000 6.200 ;
        RECT 217.400 6.100 217.800 6.200 ;
        RECT 223.000 6.100 223.400 6.200 ;
        RECT 225.400 6.100 225.800 6.200 ;
        RECT 198.200 5.800 225.800 6.100 ;
        RECT 99.000 5.200 99.300 5.800 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 11.000 5.100 11.400 5.200 ;
        RECT 14.200 5.100 14.600 5.200 ;
        RECT 4.600 4.800 14.600 5.100 ;
        RECT 46.200 5.100 46.600 5.200 ;
        RECT 47.800 5.100 48.200 5.200 ;
        RECT 46.200 4.800 48.200 5.100 ;
        RECT 62.200 5.100 62.600 5.200 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 83.000 5.100 83.400 5.200 ;
        RECT 62.200 4.800 78.500 5.100 ;
        RECT 79.000 4.800 83.400 5.100 ;
        RECT 99.000 4.800 99.400 5.200 ;
        RECT 139.000 5.100 139.400 5.200 ;
        RECT 140.600 5.100 141.000 5.200 ;
        RECT 139.000 4.800 141.000 5.100 ;
        RECT 150.200 5.100 150.600 5.200 ;
        RECT 155.800 5.100 156.200 5.200 ;
        RECT 150.200 4.800 156.200 5.100 ;
        RECT 158.200 5.100 158.600 5.200 ;
        RECT 161.400 5.100 161.800 5.200 ;
        RECT 202.200 5.100 202.600 5.200 ;
        RECT 158.200 4.800 161.800 5.100 ;
        RECT 189.400 4.800 202.600 5.100 ;
        RECT 203.000 5.100 203.400 5.200 ;
        RECT 203.000 4.800 219.300 5.100 ;
        RECT 78.200 4.200 78.500 4.800 ;
        RECT 189.400 4.200 189.700 4.800 ;
        RECT 219.000 4.200 219.300 4.800 ;
        RECT 78.200 3.800 78.600 4.200 ;
        RECT 189.400 3.800 189.800 4.200 ;
        RECT 219.000 3.800 219.400 4.200 ;
      LAYER via3 ;
        RECT 31.000 205.800 31.400 206.200 ;
        RECT 222.200 206.800 222.600 207.200 ;
        RECT 57.400 204.800 57.800 205.200 ;
        RECT 91.000 204.800 91.400 205.200 ;
        RECT 217.400 204.800 217.800 205.200 ;
        RECT 228.600 204.800 229.000 205.200 ;
        RECT 211.000 201.800 211.400 202.200 ;
        RECT 201.400 199.800 201.800 200.200 ;
        RECT 64.600 196.800 65.000 197.200 ;
        RECT 160.600 196.800 161.000 197.200 ;
        RECT 30.200 195.800 30.600 196.200 ;
        RECT 50.200 195.800 50.600 196.200 ;
        RECT 163.800 195.800 164.200 196.200 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 76.600 194.800 77.000 195.200 ;
        RECT 90.200 194.800 90.600 195.200 ;
        RECT 141.400 193.800 141.800 194.200 ;
        RECT 19.000 191.800 19.400 192.200 ;
        RECT 29.400 191.800 29.800 192.200 ;
        RECT 175.000 187.800 175.400 188.200 ;
        RECT 179.000 187.800 179.400 188.200 ;
        RECT 160.600 186.800 161.000 187.200 ;
        RECT 11.800 185.800 12.200 186.200 ;
        RECT 95.000 185.800 95.400 186.200 ;
        RECT 147.000 185.800 147.400 186.200 ;
        RECT 105.400 184.800 105.800 185.200 ;
        RECT 87.800 183.800 88.200 184.200 ;
        RECT 95.800 183.800 96.200 184.200 ;
        RECT 52.600 182.800 53.000 183.200 ;
        RECT 151.800 182.800 152.200 183.200 ;
        RECT 63.800 181.800 64.200 182.200 ;
        RECT 153.400 181.800 153.800 182.200 ;
        RECT 34.200 179.800 34.600 180.200 ;
        RECT 67.000 177.800 67.400 178.200 ;
        RECT 85.400 177.800 85.800 178.200 ;
        RECT 111.000 177.800 111.400 178.200 ;
        RECT 34.200 175.800 34.600 176.200 ;
        RECT 106.200 174.800 106.600 175.200 ;
        RECT 51.800 173.800 52.200 174.200 ;
        RECT 71.000 173.800 71.400 174.200 ;
        RECT 98.200 173.800 98.600 174.200 ;
        RECT 141.400 173.800 141.800 174.200 ;
        RECT 159.000 173.800 159.400 174.200 ;
        RECT 24.600 172.800 25.000 173.200 ;
        RECT 86.200 172.800 86.600 173.200 ;
        RECT 103.000 172.800 103.400 173.200 ;
        RECT 94.200 171.800 94.600 172.200 ;
        RECT 115.800 170.800 116.200 171.200 ;
        RECT 167.800 170.800 168.200 171.200 ;
        RECT 122.200 169.800 122.600 170.200 ;
        RECT 27.800 165.800 28.200 166.200 ;
        RECT 35.800 165.800 36.200 166.200 ;
        RECT 67.000 165.800 67.400 166.200 ;
        RECT 71.800 164.800 72.200 165.200 ;
        RECT 100.600 164.800 101.000 165.200 ;
        RECT 157.400 164.800 157.800 165.200 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 59.000 163.800 59.400 164.200 ;
        RECT 106.200 162.800 106.600 163.200 ;
        RECT 99.000 161.800 99.400 162.200 ;
        RECT 102.200 161.800 102.600 162.200 ;
        RECT 202.200 161.800 202.600 162.200 ;
        RECT 100.600 158.800 101.000 159.200 ;
        RECT 123.800 157.800 124.200 158.200 ;
        RECT 183.800 157.800 184.200 158.200 ;
        RECT 55.800 155.800 56.200 156.200 ;
        RECT 154.200 155.800 154.600 156.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 67.000 154.800 67.400 155.200 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 125.400 154.800 125.800 155.200 ;
        RECT 145.400 154.800 145.800 155.200 ;
        RECT 213.400 154.800 213.800 155.200 ;
        RECT 56.600 153.800 57.000 154.200 ;
        RECT 207.800 153.800 208.200 154.200 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 175.800 152.800 176.200 153.200 ;
        RECT 180.600 152.800 181.000 153.200 ;
        RECT 11.800 151.800 12.200 152.200 ;
        RECT 114.200 151.800 114.600 152.200 ;
        RECT 215.000 151.800 215.400 152.200 ;
        RECT 45.400 150.800 45.800 151.200 ;
        RECT 74.200 150.800 74.600 151.200 ;
        RECT 123.000 150.800 123.400 151.200 ;
        RECT 87.000 149.800 87.400 150.200 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 115.800 148.800 116.200 149.200 ;
        RECT 147.000 148.800 147.400 149.200 ;
        RECT 47.800 146.800 48.200 147.200 ;
        RECT 196.600 146.800 197.000 147.200 ;
        RECT 21.400 145.800 21.800 146.200 ;
        RECT 112.600 145.800 113.000 146.200 ;
        RECT 124.600 145.800 125.000 146.200 ;
        RECT 137.400 145.800 137.800 146.200 ;
        RECT 149.400 145.800 149.800 146.200 ;
        RECT 75.000 144.800 75.400 145.200 ;
        RECT 135.000 144.800 135.400 145.200 ;
        RECT 150.200 144.800 150.600 145.200 ;
        RECT 70.200 143.800 70.600 144.200 ;
        RECT 79.000 143.800 79.400 144.200 ;
        RECT 102.200 143.800 102.600 144.200 ;
        RECT 121.400 143.800 121.800 144.200 ;
        RECT 147.800 143.800 148.200 144.200 ;
        RECT 220.600 143.800 221.000 144.200 ;
        RECT 224.600 143.800 225.000 144.200 ;
        RECT 103.000 142.800 103.400 143.200 ;
        RECT 169.400 142.800 169.800 143.200 ;
        RECT 179.800 142.800 180.200 143.200 ;
        RECT 76.600 141.800 77.000 142.200 ;
        RECT 155.800 140.800 156.200 141.200 ;
        RECT 51.800 139.800 52.200 140.200 ;
        RECT 103.000 138.800 103.400 139.200 ;
        RECT 161.400 138.800 161.800 139.200 ;
        RECT 111.800 137.800 112.200 138.200 ;
        RECT 105.400 136.800 105.800 137.200 ;
        RECT 154.200 136.800 154.600 137.200 ;
        RECT 117.400 135.800 117.800 136.200 ;
        RECT 141.400 135.800 141.800 136.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 79.800 134.800 80.200 135.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 151.000 134.800 151.400 135.200 ;
        RECT 141.400 133.800 141.800 134.200 ;
        RECT 177.400 133.800 177.800 134.200 ;
        RECT 183.800 133.800 184.200 134.200 ;
        RECT 207.000 133.800 207.400 134.200 ;
        RECT 218.200 133.800 218.600 134.200 ;
        RECT 110.200 132.800 110.600 133.200 ;
        RECT 195.800 132.800 196.200 133.200 ;
        RECT 19.000 131.800 19.400 132.200 ;
        RECT 118.200 131.800 118.600 132.200 ;
        RECT 137.400 130.800 137.800 131.200 ;
        RECT 190.200 130.800 190.600 131.200 ;
        RECT 196.600 130.800 197.000 131.200 ;
        RECT 15.000 129.800 15.400 130.200 ;
        RECT 207.800 129.800 208.200 130.200 ;
        RECT 48.600 127.800 49.000 128.200 ;
        RECT 53.400 126.800 53.800 127.200 ;
        RECT 64.600 126.800 65.000 127.200 ;
        RECT 114.200 126.800 114.600 127.200 ;
        RECT 218.200 126.800 218.600 127.200 ;
        RECT 13.400 125.800 13.800 126.200 ;
        RECT 60.600 125.800 61.000 126.200 ;
        RECT 180.600 125.800 181.000 126.200 ;
        RECT 103.000 124.800 103.400 125.200 ;
        RECT 111.000 124.800 111.400 125.200 ;
        RECT 116.600 124.800 117.000 125.200 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 146.200 124.800 146.600 125.200 ;
        RECT 169.400 124.800 169.800 125.200 ;
        RECT 107.000 123.800 107.400 124.200 ;
        RECT 166.200 123.800 166.600 124.200 ;
        RECT 164.600 122.800 165.000 123.200 ;
        RECT 135.800 121.800 136.200 122.200 ;
        RECT 202.200 121.800 202.600 122.200 ;
        RECT 105.400 120.800 105.800 121.200 ;
        RECT 189.400 119.800 189.800 120.200 ;
        RECT 99.000 117.800 99.400 118.200 ;
        RECT 154.200 117.800 154.600 118.200 ;
        RECT 109.400 116.800 109.800 117.200 ;
        RECT 112.600 116.800 113.000 117.200 ;
        RECT 160.600 115.800 161.000 116.200 ;
        RECT 175.000 115.800 175.400 116.200 ;
        RECT 211.000 115.800 211.400 116.200 ;
        RECT 27.800 114.800 28.200 115.200 ;
        RECT 65.400 114.800 65.800 115.200 ;
        RECT 69.400 114.800 69.800 115.200 ;
        RECT 103.800 114.800 104.200 115.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 166.200 114.800 166.600 115.200 ;
        RECT 30.200 113.800 30.600 114.200 ;
        RECT 26.200 112.800 26.600 113.200 ;
        RECT 150.200 113.800 150.600 114.200 ;
        RECT 64.600 112.800 65.000 113.200 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 176.600 112.800 177.000 113.200 ;
        RECT 114.200 111.800 114.600 112.200 ;
        RECT 179.000 110.800 179.400 111.200 ;
        RECT 119.000 109.800 119.400 110.200 ;
        RECT 135.000 109.800 135.400 110.200 ;
        RECT 222.200 109.800 222.600 110.200 ;
        RECT 128.600 108.800 129.000 109.200 ;
        RECT 207.800 108.800 208.200 109.200 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 158.200 106.800 158.600 107.200 ;
        RECT 159.800 106.800 160.200 107.200 ;
        RECT 36.600 105.800 37.000 106.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 19.800 104.800 20.200 105.200 ;
        RECT 23.000 104.800 23.400 105.200 ;
        RECT 135.800 104.800 136.200 105.200 ;
        RECT 146.200 104.800 146.600 105.200 ;
        RECT 211.000 104.800 211.400 105.200 ;
        RECT 159.800 103.800 160.200 104.200 ;
        RECT 43.800 102.800 44.200 103.200 ;
        RECT 144.600 102.800 145.000 103.200 ;
        RECT 163.000 102.800 163.400 103.200 ;
        RECT 21.400 101.800 21.800 102.200 ;
        RECT 99.800 101.800 100.200 102.200 ;
        RECT 121.400 101.800 121.800 102.200 ;
        RECT 160.600 101.800 161.000 102.200 ;
        RECT 17.400 100.800 17.800 101.200 ;
        RECT 63.800 100.800 64.200 101.200 ;
        RECT 95.000 100.800 95.400 101.200 ;
        RECT 120.600 100.800 121.000 101.200 ;
        RECT 151.000 100.800 151.400 101.200 ;
        RECT 207.000 100.800 207.400 101.200 ;
        RECT 226.200 100.800 226.600 101.200 ;
        RECT 94.200 98.800 94.600 99.200 ;
        RECT 127.000 98.800 127.400 99.200 ;
        RECT 148.600 98.800 149.000 99.200 ;
        RECT 185.400 98.800 185.800 99.200 ;
        RECT 107.800 97.800 108.200 98.200 ;
        RECT 148.600 97.800 149.000 98.200 ;
        RECT 93.400 96.800 93.800 97.200 ;
        RECT 14.200 95.800 14.600 96.200 ;
        RECT 63.000 95.800 63.400 96.200 ;
        RECT 144.600 95.800 145.000 96.200 ;
        RECT 202.200 95.800 202.600 96.200 ;
        RECT 124.600 94.800 125.000 95.200 ;
        RECT 138.200 94.800 138.600 95.200 ;
        RECT 152.600 94.800 153.000 95.200 ;
        RECT 185.400 94.800 185.800 95.200 ;
        RECT 187.800 94.800 188.200 95.200 ;
        RECT 197.400 94.800 197.800 95.200 ;
        RECT 54.200 93.800 54.600 94.200 ;
        RECT 154.200 93.800 154.600 94.200 ;
        RECT 15.000 92.800 15.400 93.200 ;
        RECT 62.200 92.800 62.600 93.200 ;
        RECT 204.600 92.800 205.000 93.200 ;
        RECT 136.600 91.800 137.000 92.200 ;
        RECT 75.800 90.800 76.200 91.200 ;
        RECT 100.600 90.800 101.000 91.200 ;
        RECT 155.000 90.800 155.400 91.200 ;
        RECT 184.600 89.800 185.000 90.200 ;
        RECT 190.200 89.800 190.600 90.200 ;
        RECT 227.800 89.800 228.200 90.200 ;
        RECT 43.800 88.800 44.200 89.200 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 118.200 88.800 118.600 89.200 ;
        RECT 183.000 88.800 183.400 89.200 ;
        RECT 51.800 87.800 52.200 88.200 ;
        RECT 78.200 87.800 78.600 88.200 ;
        RECT 94.200 87.800 94.600 88.200 ;
        RECT 116.600 87.800 117.000 88.200 ;
        RECT 154.200 87.800 154.600 88.200 ;
        RECT 65.400 86.800 65.800 87.200 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 174.200 86.800 174.600 87.200 ;
        RECT 73.400 85.800 73.800 86.200 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 110.200 85.800 110.600 86.200 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 41.400 84.800 41.800 85.200 ;
        RECT 98.200 84.800 98.600 85.200 ;
        RECT 152.600 84.800 153.000 85.200 ;
        RECT 195.800 84.800 196.200 85.200 ;
        RECT 223.000 84.800 223.400 85.200 ;
        RECT 180.600 83.800 181.000 84.200 ;
        RECT 50.200 78.800 50.600 79.200 ;
        RECT 107.000 77.800 107.400 78.200 ;
        RECT 137.400 76.800 137.800 77.200 ;
        RECT 187.800 76.800 188.200 77.200 ;
        RECT 51.000 75.800 51.400 76.200 ;
        RECT 85.400 75.800 85.800 76.200 ;
        RECT 121.400 75.800 121.800 76.200 ;
        RECT 201.400 75.800 201.800 76.200 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.800 74.800 44.200 75.200 ;
        RECT 126.200 74.800 126.600 75.200 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 173.400 74.800 173.800 75.200 ;
        RECT 203.000 74.800 203.400 75.200 ;
        RECT 49.400 73.800 49.800 74.200 ;
        RECT 63.800 73.800 64.200 74.200 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 119.800 73.800 120.200 74.200 ;
        RECT 199.000 73.800 199.400 74.200 ;
        RECT 65.400 72.800 65.800 73.200 ;
        RECT 177.400 72.800 177.800 73.200 ;
        RECT 183.800 72.800 184.200 73.200 ;
        RECT 219.000 72.800 219.400 73.200 ;
        RECT 16.600 71.800 17.000 72.200 ;
        RECT 102.200 71.800 102.600 72.200 ;
        RECT 203.000 71.800 203.400 72.200 ;
        RECT 35.000 70.800 35.400 71.200 ;
        RECT 106.200 70.800 106.600 71.200 ;
        RECT 105.400 68.800 105.800 69.200 ;
        RECT 148.600 68.800 149.000 69.200 ;
        RECT 157.400 68.800 157.800 69.200 ;
        RECT 171.000 68.800 171.400 69.200 ;
        RECT 115.800 66.800 116.200 67.200 ;
        RECT 154.200 66.800 154.600 67.200 ;
        RECT 174.200 66.800 174.600 67.200 ;
        RECT 113.400 65.800 113.800 66.200 ;
        RECT 142.200 65.800 142.600 66.200 ;
        RECT 145.400 65.800 145.800 66.200 ;
        RECT 189.400 65.800 189.800 66.200 ;
        RECT 43.000 64.800 43.400 65.200 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 103.000 64.800 103.400 65.200 ;
        RECT 104.600 64.800 105.000 65.200 ;
        RECT 117.400 64.800 117.800 65.200 ;
        RECT 172.600 64.800 173.000 65.200 ;
        RECT 210.200 64.800 210.600 65.200 ;
        RECT 151.800 63.800 152.200 64.200 ;
        RECT 194.200 63.800 194.600 64.200 ;
        RECT 211.000 62.800 211.400 63.200 ;
        RECT 17.400 59.800 17.800 60.200 ;
        RECT 61.400 59.800 61.800 60.200 ;
        RECT 31.000 56.800 31.400 57.200 ;
        RECT 75.000 56.800 75.400 57.200 ;
        RECT 119.000 56.800 119.400 57.200 ;
        RECT 115.800 55.800 116.200 56.200 ;
        RECT 183.800 55.800 184.200 56.200 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 141.400 54.800 141.800 55.200 ;
        RECT 201.400 54.800 201.800 55.200 ;
        RECT 45.400 53.800 45.800 54.200 ;
        RECT 57.400 53.800 57.800 54.200 ;
        RECT 122.200 53.800 122.600 54.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 228.600 53.800 229.000 54.200 ;
        RECT 91.000 52.800 91.400 53.200 ;
        RECT 150.200 52.800 150.600 53.200 ;
        RECT 99.000 51.800 99.400 52.200 ;
        RECT 17.400 50.800 17.800 51.200 ;
        RECT 190.200 50.800 190.600 51.200 ;
        RECT 219.000 48.800 219.400 49.200 ;
        RECT 142.200 47.800 142.600 48.200 ;
        RECT 201.400 47.800 201.800 48.200 ;
        RECT 200.600 46.800 201.000 47.200 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 207.800 45.800 208.200 46.200 ;
        RECT 203.000 44.800 203.400 45.200 ;
        RECT 185.400 43.800 185.800 44.200 ;
        RECT 112.600 42.800 113.000 43.200 ;
        RECT 59.000 41.800 59.400 42.200 ;
        RECT 98.200 41.800 98.600 42.200 ;
        RECT 87.000 40.800 87.400 41.200 ;
        RECT 195.800 40.800 196.200 41.200 ;
        RECT 111.000 38.800 111.400 39.200 ;
        RECT 73.400 36.800 73.800 37.200 ;
        RECT 90.200 35.800 90.600 36.200 ;
        RECT 130.200 35.800 130.600 36.200 ;
        RECT 203.000 35.800 203.400 36.200 ;
        RECT 226.200 35.800 226.600 36.200 ;
        RECT 32.600 34.800 33.000 35.200 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 75.800 32.800 76.200 33.200 ;
        RECT 220.600 32.800 221.000 33.200 ;
        RECT 76.600 30.800 77.000 31.200 ;
        RECT 102.200 29.800 102.600 30.200 ;
        RECT 142.200 29.800 142.600 30.200 ;
        RECT 102.200 28.800 102.600 29.200 ;
        RECT 151.000 26.800 151.400 27.200 ;
        RECT 167.000 26.800 167.400 27.200 ;
        RECT 23.000 25.800 23.400 26.200 ;
        RECT 204.600 25.800 205.000 26.200 ;
        RECT 225.400 25.800 225.800 26.200 ;
        RECT 161.400 24.800 161.800 25.200 ;
        RECT 72.600 23.800 73.000 24.200 ;
        RECT 193.400 22.800 193.800 23.200 ;
        RECT 36.600 18.800 37.000 19.200 ;
        RECT 187.000 18.800 187.400 19.200 ;
        RECT 126.200 17.800 126.600 18.200 ;
        RECT 49.400 16.800 49.800 17.200 ;
        RECT 141.400 15.800 141.800 16.200 ;
        RECT 226.200 15.800 226.600 16.200 ;
        RECT 94.200 13.800 94.600 14.200 ;
        RECT 217.400 13.800 217.800 14.200 ;
        RECT 68.600 10.800 69.000 11.200 ;
        RECT 48.600 9.800 49.000 10.200 ;
        RECT 23.800 8.800 24.200 9.200 ;
        RECT 79.000 7.800 79.400 8.200 ;
        RECT 37.400 6.800 37.800 7.200 ;
        RECT 46.200 6.800 46.600 7.200 ;
        RECT 85.400 5.800 85.800 6.200 ;
      LAYER metal4 ;
        RECT 222.200 206.800 222.600 207.200 ;
        RECT 223.000 206.800 223.400 207.200 ;
        RECT 27.800 206.100 28.200 206.200 ;
        RECT 28.600 206.100 29.000 206.200 ;
        RECT 27.800 205.800 29.000 206.100 ;
        RECT 29.400 205.800 29.800 206.200 ;
        RECT 31.000 206.100 31.400 206.200 ;
        RECT 30.200 205.800 31.400 206.100 ;
        RECT 32.600 206.100 33.000 206.200 ;
        RECT 33.400 206.100 33.800 206.200 ;
        RECT 32.600 205.800 33.800 206.100 ;
        RECT 213.400 205.800 213.800 206.200 ;
        RECT 29.400 192.200 29.700 205.800 ;
        RECT 30.200 205.200 30.500 205.800 ;
        RECT 30.200 204.800 30.600 205.200 ;
        RECT 57.400 205.100 57.800 205.200 ;
        RECT 58.200 205.100 58.600 205.200 ;
        RECT 57.400 204.800 58.600 205.100 ;
        RECT 75.800 204.800 76.200 205.200 ;
        RECT 91.000 205.100 91.400 205.200 ;
        RECT 90.200 204.800 91.400 205.100 ;
        RECT 201.400 205.100 201.800 205.200 ;
        RECT 201.400 204.800 202.500 205.100 ;
        RECT 30.200 196.200 30.500 204.800 ;
        RECT 75.800 204.200 76.100 204.800 ;
        RECT 75.800 203.800 76.200 204.200 ;
        RECT 64.600 197.100 65.000 197.200 ;
        RECT 63.800 196.800 65.000 197.100 ;
        RECT 30.200 195.800 30.600 196.200 ;
        RECT 50.200 195.800 50.600 196.200 ;
        RECT 50.200 193.200 50.500 195.800 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 57.400 194.800 57.800 195.200 ;
        RECT 59.000 194.800 59.400 195.200 ;
        RECT 50.200 192.800 50.600 193.200 ;
        RECT 18.200 192.100 18.600 192.200 ;
        RECT 19.000 192.100 19.400 192.200 ;
        RECT 18.200 191.800 19.400 192.100 ;
        RECT 29.400 191.800 29.800 192.200 ;
        RECT 11.800 185.800 12.200 186.200 ;
        RECT 11.800 177.200 12.100 185.800 ;
        RECT 34.200 179.800 34.600 180.200 ;
        RECT 11.800 176.800 12.200 177.200 ;
        RECT 11.000 164.800 11.400 165.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 10.200 145.200 10.500 154.800 ;
        RECT 10.200 144.800 10.600 145.200 ;
        RECT 10.200 72.200 10.500 144.800 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 11.000 17.200 11.300 164.800 ;
        RECT 11.800 152.200 12.100 176.800 ;
        RECT 34.200 176.200 34.500 179.800 ;
        RECT 34.200 175.800 34.600 176.200 ;
        RECT 51.800 174.200 52.100 194.800 ;
        RECT 52.600 182.800 53.000 183.200 ;
        RECT 55.800 183.100 56.200 183.200 ;
        RECT 55.800 182.800 56.900 183.100 ;
        RECT 35.800 173.800 36.200 174.200 ;
        RECT 51.800 173.800 52.200 174.200 ;
        RECT 24.600 172.800 25.000 173.200 ;
        RECT 27.800 172.800 28.200 173.200 ;
        RECT 11.800 151.800 12.200 152.200 ;
        RECT 11.800 125.200 12.100 151.800 ;
        RECT 21.400 145.800 21.800 146.200 ;
        RECT 17.400 142.800 17.800 143.200 ;
        RECT 15.000 129.800 15.400 130.200 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 14.200 126.100 14.600 126.200 ;
        RECT 13.400 125.800 14.600 126.100 ;
        RECT 11.800 124.800 12.200 125.200 ;
        RECT 14.200 118.800 14.600 119.200 ;
        RECT 11.800 102.800 12.200 103.200 ;
        RECT 11.800 91.200 12.100 102.800 ;
        RECT 14.200 96.200 14.500 118.800 ;
        RECT 15.000 113.200 15.300 129.800 ;
        RECT 15.000 112.800 15.400 113.200 ;
        RECT 14.200 95.800 14.600 96.200 ;
        RECT 14.200 95.200 14.500 95.800 ;
        RECT 14.200 94.800 14.600 95.200 ;
        RECT 11.800 90.800 12.200 91.200 ;
        RECT 14.200 77.200 14.500 94.800 ;
        RECT 15.000 93.200 15.300 112.800 ;
        RECT 17.400 101.200 17.700 142.800 ;
        RECT 19.000 131.800 19.400 132.200 ;
        RECT 17.400 100.800 17.800 101.200 ;
        RECT 15.000 92.800 15.400 93.200 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 14.200 76.800 14.600 77.200 ;
        RECT 16.600 71.800 17.000 72.200 ;
        RECT 16.600 43.200 16.900 71.800 ;
        RECT 17.400 60.200 17.700 85.800 ;
        RECT 17.400 59.800 17.800 60.200 ;
        RECT 17.400 51.200 17.700 59.800 ;
        RECT 19.000 58.200 19.300 131.800 ;
        RECT 19.800 106.800 20.200 107.200 ;
        RECT 19.800 105.200 20.100 106.800 ;
        RECT 19.800 104.800 20.200 105.200 ;
        RECT 21.400 102.200 21.700 145.800 ;
        RECT 24.600 135.200 24.900 172.800 ;
        RECT 27.800 166.200 28.100 172.800 ;
        RECT 35.800 166.200 36.100 173.800 ;
        RECT 51.800 167.100 52.200 167.200 ;
        RECT 52.600 167.100 52.900 182.800 ;
        RECT 51.800 166.800 52.900 167.100 ;
        RECT 27.800 165.800 28.200 166.200 ;
        RECT 35.800 165.800 36.200 166.200 ;
        RECT 30.200 147.100 30.600 147.200 ;
        RECT 31.000 147.100 31.400 147.200 ;
        RECT 30.200 146.800 31.400 147.100 ;
        RECT 27.800 142.800 28.200 143.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 24.600 134.800 25.000 135.200 ;
        RECT 23.000 105.200 23.300 134.800 ;
        RECT 27.800 115.200 28.100 142.800 ;
        RECT 27.800 114.800 28.200 115.200 ;
        RECT 30.200 114.200 30.500 146.800 ;
        RECT 35.800 134.200 36.100 165.800 ;
        RECT 53.400 163.800 53.800 164.200 ;
        RECT 43.800 152.800 44.200 153.200 ;
        RECT 35.800 133.800 36.200 134.200 ;
        RECT 30.200 113.800 30.600 114.200 ;
        RECT 35.000 113.800 35.400 114.200 ;
        RECT 26.200 112.800 26.600 113.200 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 25.400 107.100 25.800 107.200 ;
        RECT 24.600 106.800 25.800 107.100 ;
        RECT 23.000 104.800 23.400 105.200 ;
        RECT 21.400 101.800 21.800 102.200 ;
        RECT 19.000 57.800 19.400 58.200 ;
        RECT 17.400 50.800 17.800 51.200 ;
        RECT 16.600 42.800 17.000 43.200 ;
        RECT 23.000 26.200 23.300 104.800 ;
        RECT 26.200 87.200 26.500 112.800 ;
        RECT 30.200 91.200 30.500 113.800 ;
        RECT 31.000 95.800 31.400 96.200 ;
        RECT 30.200 90.800 30.600 91.200 ;
        RECT 26.200 86.800 26.600 87.200 ;
        RECT 29.400 74.100 29.800 74.200 ;
        RECT 30.200 74.100 30.500 90.800 ;
        RECT 29.400 73.800 30.500 74.100 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 28.600 46.100 29.000 46.200 ;
        RECT 27.800 45.800 29.000 46.100 ;
        RECT 30.200 34.200 30.500 73.800 ;
        RECT 31.000 57.200 31.300 95.800 ;
        RECT 35.000 71.200 35.300 113.800 ;
        RECT 35.000 70.800 35.400 71.200 ;
        RECT 35.800 68.200 36.100 133.800 ;
        RECT 43.000 110.800 43.400 111.200 ;
        RECT 36.600 105.800 37.000 106.200 ;
        RECT 35.800 67.800 36.200 68.200 ;
        RECT 31.000 56.800 31.400 57.200 ;
        RECT 32.600 46.100 33.000 46.200 ;
        RECT 33.400 46.100 33.800 46.200 ;
        RECT 32.600 45.800 33.800 46.100 ;
        RECT 32.600 35.100 33.000 35.200 ;
        RECT 33.400 35.100 33.800 35.200 ;
        RECT 32.600 34.800 33.800 35.100 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 23.000 25.800 23.400 26.200 ;
        RECT 36.600 19.200 36.900 105.800 ;
        RECT 42.200 89.800 42.600 90.200 ;
        RECT 41.400 84.800 41.800 85.200 ;
        RECT 41.400 72.200 41.700 84.800 ;
        RECT 42.200 75.200 42.500 89.800 ;
        RECT 43.000 76.200 43.300 110.800 ;
        RECT 43.800 103.200 44.100 152.800 ;
        RECT 45.400 150.800 45.800 151.200 ;
        RECT 45.400 146.200 45.700 150.800 ;
        RECT 47.800 146.800 48.200 147.200 ;
        RECT 45.400 145.800 45.800 146.200 ;
        RECT 45.400 145.200 45.700 145.800 ;
        RECT 45.400 144.800 45.800 145.200 ;
        RECT 47.800 128.100 48.100 146.800 ;
        RECT 51.800 139.800 52.200 140.200 ;
        RECT 48.600 128.100 49.000 128.200 ;
        RECT 47.800 127.800 49.000 128.100 ;
        RECT 47.800 115.200 48.100 127.800 ;
        RECT 50.200 116.800 50.600 117.200 ;
        RECT 47.800 114.800 48.200 115.200 ;
        RECT 43.800 102.800 44.200 103.200 ;
        RECT 48.600 93.800 49.000 94.200 ;
        RECT 43.800 88.800 44.200 89.200 ;
        RECT 43.000 75.800 43.400 76.200 ;
        RECT 43.800 75.200 44.100 88.800 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.800 74.800 44.200 75.200 ;
        RECT 48.600 74.100 48.900 93.800 ;
        RECT 50.200 79.200 50.500 116.800 ;
        RECT 51.000 97.100 51.400 97.200 ;
        RECT 51.800 97.100 52.100 139.800 ;
        RECT 53.400 127.200 53.700 163.800 ;
        RECT 55.800 155.800 56.200 156.200 ;
        RECT 55.800 128.200 56.100 155.800 ;
        RECT 56.600 154.200 56.900 182.800 ;
        RECT 56.600 153.800 57.000 154.200 ;
        RECT 57.400 145.200 57.700 194.800 ;
        RECT 59.000 192.200 59.300 194.800 ;
        RECT 59.000 191.800 59.400 192.200 ;
        RECT 59.000 164.200 59.300 191.800 ;
        RECT 63.800 186.200 64.100 196.800 ;
        RECT 90.200 195.200 90.500 204.800 ;
        RECT 127.800 202.800 128.200 203.200 ;
        RECT 111.000 197.800 111.400 198.200 ;
        RECT 76.600 194.800 77.000 195.200 ;
        RECT 90.200 194.800 90.600 195.200 ;
        RECT 71.000 194.100 71.400 194.200 ;
        RECT 71.000 193.800 72.100 194.100 ;
        RECT 63.800 185.800 64.200 186.200 ;
        RECT 59.800 183.800 60.200 184.200 ;
        RECT 59.800 175.200 60.100 183.800 ;
        RECT 63.800 181.800 64.200 182.200 ;
        RECT 59.800 174.800 60.200 175.200 ;
        RECT 59.000 163.800 59.400 164.200 ;
        RECT 57.400 144.800 57.800 145.200 ;
        RECT 55.800 127.800 56.200 128.200 ;
        RECT 53.400 126.800 53.800 127.200 ;
        RECT 54.200 126.800 54.600 127.200 ;
        RECT 51.000 96.800 52.100 97.100 ;
        RECT 54.200 94.200 54.500 126.800 ;
        RECT 59.800 126.100 60.100 174.800 ;
        RECT 62.200 136.800 62.600 137.200 ;
        RECT 62.200 136.200 62.500 136.800 ;
        RECT 62.200 135.800 62.600 136.200 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 60.600 126.100 61.000 126.200 ;
        RECT 59.800 125.800 61.000 126.100 ;
        RECT 63.000 96.200 63.300 135.800 ;
        RECT 63.800 127.100 64.100 181.800 ;
        RECT 67.000 178.100 67.400 178.200 ;
        RECT 66.200 177.800 67.400 178.100 ;
        RECT 66.200 174.200 66.500 177.800 ;
        RECT 66.200 173.800 66.600 174.200 ;
        RECT 71.000 173.800 71.400 174.200 ;
        RECT 67.000 166.100 67.400 166.200 ;
        RECT 67.800 166.100 68.200 166.200 ;
        RECT 67.000 165.800 68.200 166.100 ;
        RECT 67.000 155.800 67.400 156.200 ;
        RECT 67.000 155.200 67.300 155.800 ;
        RECT 67.000 154.800 67.400 155.200 ;
        RECT 64.600 127.100 65.000 127.200 ;
        RECT 63.800 126.800 65.000 127.100 ;
        RECT 67.000 126.200 67.300 154.800 ;
        RECT 70.200 146.800 70.600 147.200 ;
        RECT 70.200 144.200 70.500 146.800 ;
        RECT 71.000 144.200 71.300 173.800 ;
        RECT 71.800 165.200 72.100 193.800 ;
        RECT 71.800 164.800 72.200 165.200 ;
        RECT 74.200 151.100 74.600 151.200 ;
        RECT 73.400 150.800 74.600 151.100 ;
        RECT 70.200 143.800 70.600 144.200 ;
        RECT 71.000 143.800 71.400 144.200 ;
        RECT 67.000 125.800 67.400 126.200 ;
        RECT 67.000 123.200 67.300 125.800 ;
        RECT 67.000 122.800 67.400 123.200 ;
        RECT 65.400 114.800 65.800 115.200 ;
        RECT 69.400 115.100 69.800 115.200 ;
        RECT 70.200 115.100 70.600 115.200 ;
        RECT 69.400 114.800 70.600 115.100 ;
        RECT 64.600 113.100 65.000 113.200 ;
        RECT 63.800 112.800 65.000 113.100 ;
        RECT 63.800 101.200 64.100 112.800 ;
        RECT 63.800 100.800 64.200 101.200 ;
        RECT 63.000 95.800 63.400 96.200 ;
        RECT 54.200 93.800 54.600 94.200 ;
        RECT 62.200 93.100 62.600 93.200 ;
        RECT 63.000 93.100 63.400 93.200 ;
        RECT 62.200 92.800 63.400 93.100 ;
        RECT 51.800 88.100 52.200 88.200 ;
        RECT 52.600 88.100 53.000 88.200 ;
        RECT 51.800 87.800 53.000 88.100 ;
        RECT 56.600 87.800 57.000 88.200 ;
        RECT 50.200 78.800 50.600 79.200 ;
        RECT 51.000 75.800 51.400 76.200 ;
        RECT 49.400 74.100 49.800 74.200 ;
        RECT 48.600 73.800 49.800 74.100 ;
        RECT 41.400 71.800 41.800 72.200 ;
        RECT 45.400 69.800 45.800 70.200 ;
        RECT 43.000 65.100 43.400 65.200 ;
        RECT 42.200 64.800 43.400 65.100 ;
        RECT 42.200 57.200 42.500 64.800 ;
        RECT 42.200 56.800 42.600 57.200 ;
        RECT 45.400 54.200 45.700 69.800 ;
        RECT 45.400 53.800 45.800 54.200 ;
        RECT 49.400 35.800 49.800 36.200 ;
        RECT 49.400 35.200 49.700 35.800 ;
        RECT 51.000 35.200 51.300 75.800 ;
        RECT 56.600 54.100 56.900 87.800 ;
        RECT 65.400 87.200 65.700 114.800 ;
        RECT 73.400 111.200 73.700 150.800 ;
        RECT 75.000 144.800 75.400 145.200 ;
        RECT 73.400 110.800 73.800 111.200 ;
        RECT 65.400 86.800 65.800 87.200 ;
        RECT 73.400 85.800 73.800 86.200 ;
        RECT 72.600 77.800 73.000 78.200 ;
        RECT 63.800 74.100 64.200 74.200 ;
        RECT 64.600 74.100 65.000 74.200 ;
        RECT 63.800 73.800 65.000 74.100 ;
        RECT 65.400 73.800 65.800 74.200 ;
        RECT 65.400 73.200 65.700 73.800 ;
        RECT 65.400 72.800 65.800 73.200 ;
        RECT 59.000 67.800 59.400 68.200 ;
        RECT 57.400 54.100 57.800 54.200 ;
        RECT 56.600 53.800 57.800 54.100 ;
        RECT 59.000 42.200 59.300 67.800 ;
        RECT 68.600 64.800 69.000 65.200 ;
        RECT 61.400 59.800 61.800 60.200 ;
        RECT 59.000 41.800 59.400 42.200 ;
        RECT 61.400 37.200 61.700 59.800 ;
        RECT 61.400 36.800 61.800 37.200 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 48.600 24.800 49.000 25.200 ;
        RECT 23.800 18.800 24.200 19.200 ;
        RECT 36.600 18.800 37.000 19.200 ;
        RECT 11.000 16.800 11.400 17.200 ;
        RECT 23.800 9.200 24.100 18.800 ;
        RECT 43.000 15.100 43.400 15.200 ;
        RECT 43.800 15.100 44.200 15.200 ;
        RECT 43.000 14.800 44.200 15.100 ;
        RECT 48.600 10.200 48.900 24.800 ;
        RECT 49.400 17.200 49.700 34.800 ;
        RECT 56.600 34.100 57.000 34.200 ;
        RECT 57.400 34.100 57.800 34.200 ;
        RECT 56.600 33.800 57.800 34.100 ;
        RECT 68.600 23.200 68.900 64.800 ;
        RECT 72.600 24.200 72.900 77.800 ;
        RECT 73.400 37.200 73.700 85.800 ;
        RECT 75.000 57.200 75.300 144.800 ;
        RECT 76.600 142.200 76.900 194.800 ;
        RECT 102.200 192.800 102.600 193.200 ;
        RECT 87.800 185.800 88.200 186.200 ;
        RECT 95.000 186.100 95.400 186.200 ;
        RECT 94.200 185.800 95.400 186.100 ;
        RECT 87.800 184.200 88.100 185.800 ;
        RECT 87.800 183.800 88.200 184.200 ;
        RECT 85.400 177.800 85.800 178.200 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 79.000 147.100 79.400 147.200 ;
        RECT 79.800 147.100 80.200 147.200 ;
        RECT 79.000 146.800 80.200 147.100 ;
        RECT 79.000 143.800 79.400 144.200 ;
        RECT 76.600 141.800 77.000 142.200 ;
        RECT 76.600 138.800 77.000 139.200 ;
        RECT 75.800 90.800 76.200 91.200 ;
        RECT 75.800 89.200 76.100 90.800 ;
        RECT 75.800 88.800 76.200 89.200 ;
        RECT 75.800 67.800 76.200 68.200 ;
        RECT 75.800 67.200 76.100 67.800 ;
        RECT 75.800 66.800 76.200 67.200 ;
        RECT 76.600 65.200 76.900 138.800 ;
        RECT 79.000 114.200 79.300 143.800 ;
        RECT 79.800 135.100 80.200 135.200 ;
        RECT 80.600 135.100 81.000 135.200 ;
        RECT 79.800 134.800 81.000 135.100 ;
        RECT 84.600 115.200 84.900 154.800 ;
        RECT 85.400 145.200 85.700 177.800 ;
        RECT 86.200 172.800 86.600 173.200 ;
        RECT 85.400 144.800 85.800 145.200 ;
        RECT 86.200 116.200 86.500 172.800 ;
        RECT 94.200 172.200 94.500 185.800 ;
        RECT 95.000 184.100 95.400 184.200 ;
        RECT 95.800 184.100 96.200 184.200 ;
        RECT 95.000 183.800 96.200 184.100 ;
        RECT 98.200 179.800 98.600 180.200 ;
        RECT 98.200 174.200 98.500 179.800 ;
        RECT 98.200 173.800 98.600 174.200 ;
        RECT 94.200 171.800 94.600 172.200 ;
        RECT 98.200 166.200 98.500 173.800 ;
        RECT 98.200 165.800 98.600 166.200 ;
        RECT 100.600 165.100 101.000 165.200 ;
        RECT 101.400 165.100 101.800 165.200 ;
        RECT 100.600 164.800 101.800 165.100 ;
        RECT 99.000 163.800 99.400 164.200 ;
        RECT 99.000 162.200 99.300 163.800 ;
        RECT 102.200 162.200 102.500 192.800 ;
        RECT 106.200 189.800 106.600 190.200 ;
        RECT 105.400 184.800 105.800 185.200 ;
        RECT 103.000 172.800 103.400 173.200 ;
        RECT 99.000 161.800 99.400 162.200 ;
        RECT 102.200 161.800 102.600 162.200 ;
        RECT 100.600 158.800 101.000 159.200 ;
        RECT 91.000 150.800 91.400 151.200 ;
        RECT 87.000 149.800 87.400 150.200 ;
        RECT 87.000 148.200 87.300 149.800 ;
        RECT 87.000 147.800 87.400 148.200 ;
        RECT 86.200 115.800 86.600 116.200 ;
        RECT 84.600 114.800 85.000 115.200 ;
        RECT 78.200 113.800 78.600 114.200 ;
        RECT 79.000 113.800 79.400 114.200 ;
        RECT 78.200 113.200 78.500 113.800 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 78.200 112.800 78.600 113.200 ;
        RECT 77.400 95.200 77.700 112.800 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 78.200 88.200 78.500 112.800 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 83.000 89.200 83.300 94.800 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 89.400 88.800 89.800 89.200 ;
        RECT 78.200 87.800 78.600 88.200 ;
        RECT 89.400 87.200 89.700 88.800 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 90.200 85.800 90.600 86.200 ;
        RECT 85.400 75.800 85.800 76.200 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 76.600 64.800 77.000 65.200 ;
        RECT 75.000 56.800 75.400 57.200 ;
        RECT 73.400 37.100 73.800 37.200 ;
        RECT 74.200 37.100 74.600 37.200 ;
        RECT 73.400 36.800 74.600 37.100 ;
        RECT 75.000 33.200 75.300 56.800 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 75.000 32.800 76.200 33.100 ;
        RECT 76.600 32.800 77.000 33.200 ;
        RECT 76.600 31.200 76.900 32.800 ;
        RECT 76.600 30.800 77.000 31.200 ;
        RECT 72.600 23.800 73.000 24.200 ;
        RECT 68.600 22.800 69.000 23.200 ;
        RECT 49.400 16.800 49.800 17.200 ;
        RECT 68.600 11.200 68.900 22.800 ;
        RECT 79.000 19.200 79.300 73.800 ;
        RECT 79.000 18.800 79.400 19.200 ;
        RECT 79.000 14.200 79.300 18.800 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 68.600 10.800 69.000 11.200 ;
        RECT 48.600 9.800 49.000 10.200 ;
        RECT 85.400 9.200 85.700 75.800 ;
        RECT 87.000 53.800 87.400 54.200 ;
        RECT 87.000 41.200 87.300 53.800 ;
        RECT 87.000 40.800 87.400 41.200 ;
        RECT 90.200 36.200 90.500 85.800 ;
        RECT 91.000 53.200 91.300 150.800 ;
        RECT 95.800 149.800 96.200 150.200 ;
        RECT 91.800 135.100 92.200 135.200 ;
        RECT 92.600 135.100 93.000 135.200 ;
        RECT 91.800 134.800 93.000 135.100 ;
        RECT 92.600 125.800 93.000 126.200 ;
        RECT 92.600 97.100 92.900 125.800 ;
        RECT 94.200 105.800 94.600 106.200 ;
        RECT 94.200 99.200 94.500 105.800 ;
        RECT 95.000 100.800 95.400 101.200 ;
        RECT 95.000 99.200 95.300 100.800 ;
        RECT 94.200 98.800 94.600 99.200 ;
        RECT 95.000 98.800 95.400 99.200 ;
        RECT 93.400 97.100 93.800 97.200 ;
        RECT 92.600 96.800 93.800 97.100 ;
        RECT 95.000 96.800 95.400 97.200 ;
        RECT 94.200 87.800 94.600 88.200 ;
        RECT 91.000 52.800 91.400 53.200 ;
        RECT 90.200 35.800 90.600 36.200 ;
        RECT 90.200 24.200 90.500 35.800 ;
        RECT 91.000 34.800 91.400 35.200 ;
        RECT 91.000 31.200 91.300 34.800 ;
        RECT 91.000 30.800 91.400 31.200 ;
        RECT 94.200 27.200 94.500 87.800 ;
        RECT 95.000 85.200 95.300 96.800 ;
        RECT 95.000 84.800 95.400 85.200 ;
        RECT 95.800 70.200 96.100 149.800 ;
        RECT 99.000 117.800 99.400 118.200 ;
        RECT 98.200 95.100 98.600 95.200 ;
        RECT 99.000 95.100 99.300 117.800 ;
        RECT 99.800 103.800 100.200 104.200 ;
        RECT 99.800 102.200 100.100 103.800 ;
        RECT 99.800 101.800 100.200 102.200 ;
        RECT 100.600 101.200 100.900 158.800 ;
        RECT 102.200 144.800 102.600 145.200 ;
        RECT 102.200 144.200 102.500 144.800 ;
        RECT 102.200 143.800 102.600 144.200 ;
        RECT 103.000 143.200 103.300 172.800 ;
        RECT 104.600 171.800 105.000 172.200 ;
        RECT 104.600 153.200 104.900 171.800 ;
        RECT 105.400 166.200 105.700 184.800 ;
        RECT 106.200 175.200 106.500 189.800 ;
        RECT 111.000 178.200 111.300 197.800 ;
        RECT 122.200 194.800 122.600 195.200 ;
        RECT 115.800 193.800 116.200 194.200 ;
        RECT 111.000 177.800 111.400 178.200 ;
        RECT 106.200 174.800 106.600 175.200 ;
        RECT 115.800 171.200 116.100 193.800 ;
        RECT 115.800 170.800 116.200 171.200 ;
        RECT 122.200 170.200 122.500 194.800 ;
        RECT 123.000 174.800 123.400 175.200 ;
        RECT 122.200 169.800 122.600 170.200 ;
        RECT 105.400 165.800 105.800 166.200 ;
        RECT 121.400 165.800 121.800 166.200 ;
        RECT 106.200 162.800 106.600 163.200 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 105.400 146.800 105.800 147.200 ;
        RECT 103.000 142.800 103.400 143.200 ;
        RECT 103.000 138.800 103.400 139.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 101.400 126.200 101.700 134.800 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 103.000 125.200 103.300 138.800 ;
        RECT 105.400 137.200 105.700 146.800 ;
        RECT 105.400 136.800 105.800 137.200 ;
        RECT 103.000 125.100 103.400 125.200 ;
        RECT 103.800 125.100 104.200 125.200 ;
        RECT 103.000 124.800 104.200 125.100 ;
        RECT 105.400 121.200 105.700 136.800 ;
        RECT 105.400 120.800 105.800 121.200 ;
        RECT 101.400 116.800 101.800 117.200 ;
        RECT 101.400 105.200 101.700 116.800 ;
        RECT 105.400 115.200 105.700 120.800 ;
        RECT 102.200 114.800 102.600 115.200 ;
        RECT 103.000 115.100 103.400 115.200 ;
        RECT 103.800 115.100 104.200 115.200 ;
        RECT 103.000 114.800 104.200 115.100 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 105.400 114.800 105.800 115.200 ;
        RECT 102.200 113.200 102.500 114.800 ;
        RECT 102.200 112.800 102.600 113.200 ;
        RECT 101.400 104.800 101.800 105.200 ;
        RECT 101.400 103.200 101.700 104.800 ;
        RECT 101.400 102.800 101.800 103.200 ;
        RECT 100.600 100.800 101.000 101.200 ;
        RECT 98.200 94.800 99.300 95.100 ;
        RECT 100.600 90.800 101.000 91.200 ;
        RECT 98.200 87.800 98.600 88.200 ;
        RECT 98.200 85.200 98.500 87.800 ;
        RECT 98.200 84.800 98.600 85.200 ;
        RECT 99.000 74.800 99.400 75.200 ;
        RECT 95.800 69.800 96.200 70.200 ;
        RECT 95.800 67.200 96.100 69.800 ;
        RECT 95.800 66.800 96.200 67.200 ;
        RECT 99.000 52.200 99.300 74.800 ;
        RECT 99.800 68.800 100.200 69.200 ;
        RECT 99.800 68.200 100.100 68.800 ;
        RECT 99.800 67.800 100.200 68.200 ;
        RECT 100.600 67.200 100.900 90.800 ;
        RECT 102.200 72.200 102.500 112.800 ;
        RECT 103.800 109.800 104.200 110.200 ;
        RECT 103.000 80.800 103.400 81.200 ;
        RECT 102.200 71.800 102.600 72.200 ;
        RECT 102.200 70.800 102.600 71.200 ;
        RECT 102.200 68.200 102.500 70.800 ;
        RECT 102.200 67.800 102.600 68.200 ;
        RECT 100.600 66.800 101.000 67.200 ;
        RECT 99.000 51.800 99.400 52.200 ;
        RECT 98.200 42.100 98.600 42.200 ;
        RECT 99.000 42.100 99.400 42.200 ;
        RECT 98.200 41.800 99.400 42.100 ;
        RECT 102.200 30.200 102.500 67.800 ;
        RECT 103.000 65.200 103.300 80.800 ;
        RECT 103.000 64.800 103.400 65.200 ;
        RECT 103.000 49.800 103.400 50.200 ;
        RECT 103.000 35.200 103.300 49.800 ;
        RECT 103.800 37.200 104.100 109.800 ;
        RECT 104.600 96.200 104.900 114.800 ;
        RECT 105.400 97.800 105.800 98.200 ;
        RECT 104.600 95.800 105.000 96.200 ;
        RECT 104.600 86.200 104.900 95.800 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 105.400 69.200 105.700 97.800 ;
        RECT 106.200 96.200 106.500 162.800 ;
        RECT 114.200 158.800 114.600 159.200 ;
        RECT 114.200 152.200 114.500 158.800 ;
        RECT 118.200 153.800 118.600 154.200 ;
        RECT 114.200 151.800 114.600 152.200 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 115.800 148.800 116.200 149.200 ;
        RECT 112.600 145.800 113.000 146.200 ;
        RECT 111.800 137.800 112.200 138.200 ;
        RECT 110.200 134.800 110.600 135.200 ;
        RECT 110.200 133.200 110.500 134.800 ;
        RECT 110.200 132.800 110.600 133.200 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 111.000 125.200 111.300 125.800 ;
        RECT 111.000 124.800 111.400 125.200 ;
        RECT 107.000 123.800 107.400 124.200 ;
        RECT 107.800 123.800 108.200 124.200 ;
        RECT 106.200 95.800 106.600 96.200 ;
        RECT 107.000 78.200 107.300 123.800 ;
        RECT 107.800 98.200 108.100 123.800 ;
        RECT 108.600 119.800 109.000 120.200 ;
        RECT 108.600 98.200 108.900 119.800 ;
        RECT 111.000 117.800 111.400 118.200 ;
        RECT 109.400 117.100 109.800 117.200 ;
        RECT 110.200 117.100 110.600 117.200 ;
        RECT 109.400 116.800 110.600 117.100 ;
        RECT 107.800 97.800 108.200 98.200 ;
        RECT 108.600 97.800 109.000 98.200 ;
        RECT 111.000 86.200 111.300 117.800 ;
        RECT 111.800 117.100 112.100 137.800 ;
        RECT 112.600 123.100 112.900 145.800 ;
        RECT 113.400 124.200 113.700 148.800 ;
        RECT 114.200 127.800 114.600 128.200 ;
        RECT 114.200 127.200 114.500 127.800 ;
        RECT 114.200 126.800 114.600 127.200 ;
        RECT 113.400 123.800 113.800 124.200 ;
        RECT 112.600 122.800 113.700 123.100 ;
        RECT 112.600 117.100 113.000 117.200 ;
        RECT 111.800 116.800 113.000 117.100 ;
        RECT 113.400 94.200 113.700 122.800 ;
        RECT 114.200 111.800 114.600 112.200 ;
        RECT 114.200 109.200 114.500 111.800 ;
        RECT 114.200 108.800 114.600 109.200 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 110.200 85.800 110.600 86.200 ;
        RECT 111.000 85.800 111.400 86.200 ;
        RECT 107.000 77.800 107.400 78.200 ;
        RECT 109.400 73.800 109.800 74.200 ;
        RECT 106.200 72.800 106.600 73.200 ;
        RECT 106.200 71.200 106.500 72.800 ;
        RECT 106.200 70.800 106.600 71.200 ;
        RECT 105.400 68.800 105.800 69.200 ;
        RECT 104.600 64.800 105.000 65.200 ;
        RECT 103.800 36.800 104.200 37.200 ;
        RECT 104.600 36.200 104.900 64.800 ;
        RECT 109.400 52.200 109.700 73.800 ;
        RECT 109.400 51.800 109.800 52.200 ;
        RECT 110.200 42.200 110.500 85.800 ;
        RECT 110.200 41.800 110.600 42.200 ;
        RECT 110.200 37.200 110.500 41.800 ;
        RECT 111.000 39.200 111.300 85.800 ;
        RECT 111.800 73.800 112.200 74.200 ;
        RECT 111.800 55.200 112.100 73.800 ;
        RECT 112.600 68.800 113.000 69.200 ;
        RECT 112.600 68.200 112.900 68.800 ;
        RECT 112.600 67.800 113.000 68.200 ;
        RECT 113.400 66.200 113.700 93.800 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 115.000 75.100 115.400 75.200 ;
        RECT 114.200 74.800 115.400 75.100 ;
        RECT 115.800 67.200 116.100 148.800 ;
        RECT 117.400 136.100 117.800 136.200 ;
        RECT 116.600 135.800 117.800 136.100 ;
        RECT 116.600 125.200 116.900 135.800 ;
        RECT 118.200 132.200 118.500 153.800 ;
        RECT 119.000 145.800 119.400 146.200 ;
        RECT 118.200 131.800 118.600 132.200 ;
        RECT 116.600 124.800 117.000 125.200 ;
        RECT 117.400 114.800 117.800 115.200 ;
        RECT 116.600 113.800 117.000 114.200 ;
        RECT 116.600 113.200 116.900 113.800 ;
        RECT 116.600 112.800 117.000 113.200 ;
        RECT 116.600 88.200 116.900 112.800 ;
        RECT 117.400 89.100 117.700 114.800 ;
        RECT 119.000 110.200 119.300 145.800 ;
        RECT 121.400 144.200 121.700 165.800 ;
        RECT 121.400 143.800 121.800 144.200 ;
        RECT 119.800 126.100 120.200 126.200 ;
        RECT 120.600 126.100 121.000 126.200 ;
        RECT 119.800 125.800 121.000 126.100 ;
        RECT 119.800 120.800 120.200 121.200 ;
        RECT 119.800 115.200 120.100 120.800 ;
        RECT 119.800 114.800 120.200 115.200 ;
        RECT 119.000 109.800 119.400 110.200 ;
        RECT 121.400 107.200 121.700 143.800 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 121.400 106.200 121.700 106.800 ;
        RECT 121.400 105.800 121.800 106.200 ;
        RECT 121.400 101.800 121.800 102.200 ;
        RECT 120.600 100.800 121.000 101.200 ;
        RECT 118.200 89.100 118.600 89.200 ;
        RECT 117.400 88.800 118.600 89.100 ;
        RECT 116.600 87.800 117.000 88.200 ;
        RECT 116.600 71.200 116.900 87.800 ;
        RECT 116.600 70.800 117.000 71.200 ;
        RECT 115.800 66.800 116.200 67.200 ;
        RECT 113.400 65.800 113.800 66.200 ;
        RECT 117.400 65.200 117.700 88.800 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 119.000 73.800 120.200 74.100 ;
        RECT 117.400 64.800 117.800 65.200 ;
        RECT 120.600 57.200 120.900 100.800 ;
        RECT 121.400 76.200 121.700 101.800 ;
        RECT 121.400 75.800 121.800 76.200 ;
        RECT 122.200 74.200 122.500 169.800 ;
        RECT 123.000 151.200 123.300 174.800 ;
        RECT 125.400 165.100 125.800 165.200 ;
        RECT 126.200 165.100 126.600 165.200 ;
        RECT 125.400 164.800 126.600 165.100 ;
        RECT 123.800 161.800 124.200 162.200 ;
        RECT 123.800 158.200 124.100 161.800 ;
        RECT 123.800 157.800 124.200 158.200 ;
        RECT 123.000 150.800 123.400 151.200 ;
        RECT 123.800 146.100 124.100 157.800 ;
        RECT 127.800 155.200 128.100 202.800 ;
        RECT 156.600 200.100 157.000 200.200 ;
        RECT 156.600 199.800 157.700 200.100 ;
        RECT 141.400 193.800 141.800 194.200 ;
        RECT 141.400 174.200 141.700 193.800 ;
        RECT 147.000 185.800 147.400 186.200 ;
        RECT 129.400 174.100 129.800 174.200 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 129.400 173.800 130.600 174.100 ;
        RECT 141.400 173.800 141.800 174.200 ;
        RECT 136.600 165.100 137.000 165.200 ;
        RECT 136.600 164.800 137.700 165.100 ;
        RECT 125.400 154.800 125.800 155.200 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 124.600 146.100 125.000 146.200 ;
        RECT 123.800 145.800 125.000 146.100 ;
        RECT 124.600 142.200 124.900 145.800 ;
        RECT 124.600 141.800 125.000 142.200 ;
        RECT 125.400 116.200 125.700 154.800 ;
        RECT 127.800 148.100 128.200 148.200 ;
        RECT 128.600 148.100 129.000 148.200 ;
        RECT 127.800 147.800 129.000 148.100 ;
        RECT 130.200 147.800 130.600 148.200 ;
        RECT 130.200 146.200 130.500 147.800 ;
        RECT 137.400 146.200 137.700 164.800 ;
        RECT 143.800 156.800 144.200 157.200 ;
        RECT 129.400 145.800 129.800 146.200 ;
        RECT 130.200 145.800 130.600 146.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 137.400 145.800 137.800 146.200 ;
        RECT 142.200 146.100 142.600 146.200 ;
        RECT 143.000 146.100 143.400 146.200 ;
        RECT 142.200 145.800 143.400 146.100 ;
        RECT 127.000 136.800 127.400 137.200 ;
        RECT 125.400 115.800 125.800 116.200 ;
        RECT 127.000 99.200 127.300 136.800 ;
        RECT 127.800 115.800 128.200 116.200 ;
        RECT 127.800 115.200 128.100 115.800 ;
        RECT 127.800 114.800 128.200 115.200 ;
        RECT 129.400 113.200 129.700 145.800 ;
        RECT 135.000 145.200 135.300 145.800 ;
        RECT 135.000 144.800 135.400 145.200 ;
        RECT 135.800 143.800 136.200 144.200 ;
        RECT 135.000 135.800 135.400 136.200 ;
        RECT 135.000 125.200 135.300 135.800 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 135.800 122.200 136.100 143.800 ;
        RECT 140.600 136.100 141.000 136.200 ;
        RECT 141.400 136.100 141.800 136.200 ;
        RECT 140.600 135.800 141.800 136.100 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 139.000 135.100 139.400 135.200 ;
        RECT 138.200 134.800 139.400 135.100 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 143.800 134.200 144.100 156.800 ;
        RECT 147.000 155.200 147.300 185.800 ;
        RECT 155.000 183.800 155.400 184.200 ;
        RECT 151.800 182.800 152.200 183.200 ;
        RECT 145.400 154.800 145.800 155.200 ;
        RECT 147.000 155.100 147.400 155.200 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 147.000 154.800 148.200 155.100 ;
        RECT 145.400 137.200 145.700 154.800 ;
        RECT 147.000 149.200 147.300 154.800 ;
        RECT 147.000 148.800 147.400 149.200 ;
        RECT 147.800 148.800 148.200 149.200 ;
        RECT 146.200 145.800 146.600 146.200 ;
        RECT 145.400 136.800 145.800 137.200 ;
        RECT 145.400 135.800 145.800 136.200 ;
        RECT 145.400 135.200 145.700 135.800 ;
        RECT 145.400 134.800 145.800 135.200 ;
        RECT 146.200 134.200 146.500 145.800 ;
        RECT 147.800 144.200 148.100 148.800 ;
        RECT 149.400 146.100 149.800 146.200 ;
        RECT 150.200 146.100 150.600 146.200 ;
        RECT 149.400 145.800 150.600 146.100 ;
        RECT 149.400 145.100 149.800 145.200 ;
        RECT 150.200 145.100 150.600 145.200 ;
        RECT 149.400 144.800 150.600 145.100 ;
        RECT 147.800 143.800 148.200 144.200 ;
        RECT 151.000 134.800 151.400 135.200 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 137.400 133.800 137.800 134.200 ;
        RECT 141.400 133.800 141.800 134.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 146.200 133.800 146.600 134.200 ;
        RECT 137.400 131.200 137.700 133.800 ;
        RECT 137.400 130.800 137.800 131.200 ;
        RECT 138.200 124.800 138.600 125.200 ;
        RECT 135.800 121.800 136.200 122.200 ;
        RECT 129.400 112.800 129.800 113.200 ;
        RECT 128.600 108.800 129.000 109.200 ;
        RECT 127.000 98.800 127.400 99.200 ;
        RECT 124.600 94.800 125.000 95.200 ;
        RECT 122.200 73.800 122.600 74.200 ;
        RECT 121.400 64.100 121.800 64.200 ;
        RECT 121.400 63.800 122.500 64.100 ;
        RECT 119.000 57.100 119.400 57.200 ;
        RECT 119.800 57.100 120.200 57.200 ;
        RECT 119.000 56.800 120.200 57.100 ;
        RECT 120.600 56.800 121.000 57.200 ;
        RECT 115.800 55.800 116.200 56.200 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 112.600 42.800 113.000 43.200 ;
        RECT 111.000 38.800 111.400 39.200 ;
        RECT 110.200 36.800 110.600 37.200 ;
        RECT 104.600 35.800 105.000 36.200 ;
        RECT 103.000 34.800 103.400 35.200 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 103.800 33.800 105.000 34.100 ;
        RECT 102.200 29.800 102.600 30.200 ;
        RECT 101.400 29.100 101.800 29.200 ;
        RECT 102.200 29.100 102.600 29.200 ;
        RECT 101.400 28.800 102.600 29.100 ;
        RECT 112.600 28.200 112.900 42.800 ;
        RECT 112.600 27.800 113.000 28.200 ;
        RECT 94.200 26.800 94.600 27.200 ;
        RECT 90.200 23.800 90.600 24.200 ;
        RECT 94.200 14.200 94.500 26.800 ;
        RECT 115.000 16.100 115.400 16.200 ;
        RECT 115.800 16.100 116.100 55.800 ;
        RECT 122.200 54.200 122.500 63.800 ;
        RECT 123.000 57.100 123.400 57.200 ;
        RECT 123.800 57.100 124.200 57.200 ;
        RECT 123.000 56.800 124.200 57.100 ;
        RECT 122.200 53.800 122.600 54.200 ;
        RECT 124.600 53.200 124.900 94.800 ;
        RECT 125.400 93.100 125.800 93.200 ;
        RECT 126.200 93.100 126.600 93.200 ;
        RECT 125.400 92.800 126.600 93.100 ;
        RECT 126.200 74.800 126.600 75.200 ;
        RECT 125.400 54.100 125.800 54.200 ;
        RECT 126.200 54.100 126.500 74.800 ;
        RECT 128.600 57.200 128.900 108.800 ;
        RECT 129.400 93.200 129.700 112.800 ;
        RECT 135.000 109.800 135.400 110.200 ;
        RECT 129.400 92.800 129.800 93.200 ;
        RECT 135.000 88.200 135.300 109.800 ;
        RECT 135.800 105.100 136.200 105.200 ;
        RECT 136.600 105.100 137.000 105.200 ;
        RECT 135.800 104.800 137.000 105.100 ;
        RECT 138.200 95.200 138.500 124.800 ;
        RECT 141.400 114.200 141.700 133.800 ;
        RECT 144.600 132.800 145.000 133.200 ;
        RECT 143.000 127.100 143.400 127.200 ;
        RECT 143.800 127.100 144.200 127.200 ;
        RECT 143.000 126.800 144.200 127.100 ;
        RECT 142.200 120.800 142.600 121.200 ;
        RECT 141.400 113.800 141.800 114.200 ;
        RECT 142.200 113.200 142.500 120.800 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 142.200 98.200 142.500 112.800 ;
        RECT 144.600 103.200 144.900 132.800 ;
        RECT 146.200 125.200 146.500 133.800 ;
        RECT 146.200 124.800 146.600 125.200 ;
        RECT 150.200 113.800 150.600 114.200 ;
        RECT 148.600 112.800 149.000 113.200 ;
        RECT 146.200 104.800 146.600 105.200 ;
        RECT 146.200 104.200 146.500 104.800 ;
        RECT 146.200 103.800 146.600 104.200 ;
        RECT 144.600 102.800 145.000 103.200 ;
        RECT 148.600 99.200 148.900 112.800 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 148.600 98.800 149.000 99.200 ;
        RECT 142.200 97.800 142.600 98.200 ;
        RECT 148.600 97.800 149.000 98.200 ;
        RECT 147.800 96.800 148.200 97.200 ;
        RECT 144.600 95.800 145.000 96.200 ;
        RECT 138.200 94.800 138.600 95.200 ;
        RECT 136.600 92.100 137.000 92.200 ;
        RECT 135.800 91.800 137.000 92.100 ;
        RECT 135.000 87.800 135.400 88.200 ;
        RECT 130.200 69.800 130.600 70.200 ;
        RECT 128.600 56.800 129.000 57.200 ;
        RECT 125.400 53.800 126.500 54.100 ;
        RECT 124.600 52.800 125.000 53.200 ;
        RECT 117.400 36.800 117.800 37.200 ;
        RECT 117.400 36.200 117.700 36.800 ;
        RECT 117.400 35.800 117.800 36.200 ;
        RECT 117.400 32.800 117.800 33.200 ;
        RECT 117.400 30.200 117.700 32.800 ;
        RECT 117.400 29.800 117.800 30.200 ;
        RECT 126.200 18.200 126.500 53.800 ;
        RECT 130.200 36.200 130.500 69.800 ;
        RECT 135.800 65.200 136.100 91.800 ;
        RECT 137.400 76.800 137.800 77.200 ;
        RECT 135.800 64.800 136.200 65.200 ;
        RECT 137.400 47.200 137.700 76.800 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 142.200 65.800 142.600 66.200 ;
        RECT 141.400 54.800 141.800 55.200 ;
        RECT 137.400 46.800 137.800 47.200 ;
        RECT 130.200 35.800 130.600 36.200 ;
        RECT 141.400 20.200 141.700 54.800 ;
        RECT 142.200 48.200 142.500 65.800 ;
        RECT 143.000 61.200 143.300 74.800 ;
        RECT 144.600 63.200 144.900 95.800 ;
        RECT 145.400 67.800 145.800 68.200 ;
        RECT 145.400 66.200 145.700 67.800 ;
        RECT 145.400 65.800 145.800 66.200 ;
        RECT 144.600 62.800 145.000 63.200 ;
        RECT 143.000 60.800 143.400 61.200 ;
        RECT 142.200 47.800 142.600 48.200 ;
        RECT 143.000 42.200 143.300 60.800 ;
        RECT 147.800 55.200 148.100 96.800 ;
        RECT 148.600 77.200 148.900 97.800 ;
        RECT 148.600 76.800 149.000 77.200 ;
        RECT 148.600 69.800 149.000 70.200 ;
        RECT 148.600 69.200 148.900 69.800 ;
        RECT 148.600 68.800 149.000 69.200 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 146.200 52.200 146.500 53.800 ;
        RECT 146.200 51.800 146.600 52.200 ;
        RECT 143.000 41.800 143.400 42.200 ;
        RECT 142.200 29.800 142.600 30.200 ;
        RECT 142.200 23.200 142.500 29.800 ;
        RECT 142.200 22.800 142.600 23.200 ;
        RECT 141.400 19.800 141.800 20.200 ;
        RECT 126.200 17.800 126.600 18.200 ;
        RECT 126.200 17.200 126.500 17.800 ;
        RECT 126.200 16.800 126.600 17.200 ;
        RECT 115.000 15.800 116.100 16.100 ;
        RECT 141.400 16.200 141.700 19.800 ;
        RECT 141.400 15.800 141.800 16.200 ;
        RECT 115.000 15.200 115.300 15.800 ;
        RECT 115.000 14.800 115.400 15.200 ;
        RECT 94.200 13.800 94.600 14.200 ;
        RECT 147.800 13.200 148.100 54.800 ;
        RECT 149.400 54.200 149.700 106.800 ;
        RECT 150.200 56.100 150.500 113.800 ;
        RECT 151.000 101.200 151.300 134.800 ;
        RECT 151.800 116.200 152.100 182.800 ;
        RECT 155.000 182.200 155.300 183.800 ;
        RECT 153.400 181.800 153.800 182.200 ;
        RECT 155.000 181.800 155.400 182.200 ;
        RECT 152.600 173.800 153.000 174.200 ;
        RECT 152.600 169.200 152.900 173.800 ;
        RECT 152.600 168.800 153.000 169.200 ;
        RECT 152.600 147.200 152.900 168.800 ;
        RECT 153.400 162.200 153.700 181.800 ;
        RECT 155.800 166.800 156.200 167.200 ;
        RECT 155.800 166.200 156.100 166.800 ;
        RECT 155.800 165.800 156.200 166.200 ;
        RECT 153.400 161.800 153.800 162.200 ;
        RECT 154.200 155.800 154.600 156.200 ;
        RECT 152.600 146.800 153.000 147.200 ;
        RECT 153.400 141.800 153.800 142.200 ;
        RECT 152.600 140.100 153.000 140.200 ;
        RECT 153.400 140.100 153.700 141.800 ;
        RECT 152.600 139.800 153.700 140.100 ;
        RECT 154.200 138.200 154.500 155.800 ;
        RECT 155.000 152.800 155.400 153.200 ;
        RECT 154.200 137.800 154.600 138.200 ;
        RECT 154.200 136.800 154.600 137.200 ;
        RECT 154.200 118.200 154.500 136.800 ;
        RECT 154.200 117.800 154.600 118.200 ;
        RECT 151.800 115.800 152.200 116.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 151.000 100.800 151.400 101.200 ;
        RECT 151.800 64.200 152.100 114.800 ;
        RECT 152.600 95.800 153.000 96.200 ;
        RECT 152.600 95.200 152.900 95.800 ;
        RECT 152.600 94.800 153.000 95.200 ;
        RECT 154.200 94.800 154.600 95.200 ;
        RECT 154.200 94.200 154.500 94.800 ;
        RECT 154.200 93.800 154.600 94.200 ;
        RECT 155.000 91.200 155.300 152.800 ;
        RECT 155.800 141.200 156.100 165.800 ;
        RECT 157.400 165.200 157.700 199.800 ;
        RECT 201.400 199.800 201.800 200.200 ;
        RECT 160.600 196.800 161.000 197.200 ;
        RECT 160.600 187.200 160.900 196.800 ;
        RECT 163.800 195.800 164.200 196.200 ;
        RECT 159.000 186.800 159.400 187.200 ;
        RECT 160.600 186.800 161.000 187.200 ;
        RECT 159.000 174.200 159.300 186.800 ;
        RECT 160.600 179.100 161.000 179.200 ;
        RECT 160.600 178.800 161.700 179.100 ;
        RECT 159.000 173.800 159.400 174.200 ;
        RECT 157.400 164.800 157.800 165.200 ;
        RECT 155.800 140.800 156.200 141.200 ;
        RECT 161.400 139.200 161.700 178.800 ;
        RECT 163.800 145.200 164.100 195.800 ;
        RECT 185.400 192.800 185.800 193.200 ;
        RECT 175.000 188.100 175.400 188.200 ;
        RECT 175.800 188.100 176.200 188.200 ;
        RECT 175.000 187.800 176.200 188.100 ;
        RECT 178.200 188.100 178.600 188.200 ;
        RECT 179.000 188.100 179.400 188.200 ;
        RECT 178.200 187.800 179.400 188.100 ;
        RECT 185.400 186.200 185.700 192.800 ;
        RECT 185.400 185.800 185.800 186.200 ;
        RECT 179.800 175.800 180.200 176.200 ;
        RECT 167.800 170.800 168.200 171.200 ;
        RECT 168.600 170.800 169.000 171.200 ;
        RECT 163.800 144.800 164.200 145.200 ;
        RECT 167.800 142.200 168.100 170.800 ;
        RECT 167.800 141.800 168.200 142.200 ;
        RECT 161.400 138.800 161.800 139.200 ;
        RECT 156.600 135.800 157.000 136.200 ;
        RECT 156.600 132.200 156.900 135.800 ;
        RECT 157.400 133.100 157.800 133.200 ;
        RECT 157.400 132.800 158.500 133.100 ;
        RECT 156.600 131.800 157.000 132.200 ;
        RECT 155.800 116.800 156.200 117.200 ;
        RECT 155.800 116.200 156.100 116.800 ;
        RECT 155.800 115.800 156.200 116.200 ;
        RECT 156.600 106.200 156.900 131.800 ;
        RECT 158.200 107.200 158.500 132.800 ;
        RECT 160.600 115.800 161.000 116.200 ;
        RECT 158.200 106.800 158.600 107.200 ;
        RECT 159.800 106.800 160.200 107.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 157.400 106.100 157.800 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 157.400 105.800 158.600 106.100 ;
        RECT 156.600 105.100 157.000 105.200 ;
        RECT 157.400 105.100 157.800 105.200 ;
        RECT 156.600 104.800 157.800 105.100 ;
        RECT 159.800 104.200 160.100 106.800 ;
        RECT 159.800 103.800 160.200 104.200 ;
        RECT 160.600 102.200 160.900 115.800 ;
        RECT 160.600 101.800 161.000 102.200 ;
        RECT 157.400 93.800 157.800 94.200 ;
        RECT 155.000 90.800 155.400 91.200 ;
        RECT 154.200 89.800 154.600 90.200 ;
        RECT 152.600 89.100 153.000 89.200 ;
        RECT 153.400 89.100 153.800 89.200 ;
        RECT 152.600 88.800 153.800 89.100 ;
        RECT 154.200 88.200 154.500 89.800 ;
        RECT 154.200 87.800 154.600 88.200 ;
        RECT 156.600 87.800 157.000 88.200 ;
        RECT 156.600 87.200 156.900 87.800 ;
        RECT 152.600 86.800 153.000 87.200 ;
        RECT 156.600 86.800 157.000 87.200 ;
        RECT 152.600 85.200 152.900 86.800 ;
        RECT 152.600 84.800 153.000 85.200 ;
        RECT 153.400 83.800 153.800 84.200 ;
        RECT 151.800 63.800 152.200 64.200 ;
        RECT 150.200 55.800 151.300 56.100 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 148.600 31.200 148.900 45.800 ;
        RECT 148.600 30.800 149.000 31.200 ;
        RECT 147.800 12.800 148.200 13.200 ;
        RECT 149.400 11.200 149.700 53.800 ;
        RECT 150.200 52.800 150.600 53.200 ;
        RECT 150.200 42.200 150.500 52.800 ;
        RECT 150.200 41.800 150.600 42.200 ;
        RECT 151.000 34.200 151.300 55.800 ;
        RECT 153.400 44.200 153.700 83.800 ;
        RECT 157.400 69.200 157.700 93.800 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 157.400 68.800 157.800 69.200 ;
        RECT 158.200 69.100 158.600 69.200 ;
        RECT 159.000 69.100 159.400 69.200 ;
        RECT 158.200 68.800 159.400 69.100 ;
        RECT 154.200 67.800 154.600 68.200 ;
        RECT 154.200 67.200 154.500 67.800 ;
        RECT 154.200 66.800 154.600 67.200 ;
        RECT 155.000 67.100 155.400 67.200 ;
        RECT 155.800 67.100 156.200 67.200 ;
        RECT 155.000 66.800 156.200 67.100 ;
        RECT 153.400 43.800 153.800 44.200 ;
        RECT 161.400 37.200 161.700 138.800 ;
        RECT 168.600 125.100 168.900 170.800 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 178.200 165.100 178.600 165.200 ;
        RECT 179.000 165.100 179.400 165.200 ;
        RECT 178.200 164.800 179.400 165.100 ;
        RECT 169.400 143.200 169.700 164.800 ;
        RECT 179.800 156.200 180.100 175.800 ;
        RECT 183.800 157.800 184.200 158.200 ;
        RECT 179.800 155.800 180.200 156.200 ;
        RECT 180.600 154.100 181.000 154.200 ;
        RECT 181.400 154.100 181.800 154.200 ;
        RECT 180.600 153.800 181.800 154.100 ;
        RECT 175.800 152.800 176.200 153.200 ;
        RECT 180.600 152.800 181.000 153.200 ;
        RECT 169.400 142.800 169.800 143.200 ;
        RECT 169.400 125.100 169.800 125.200 ;
        RECT 168.600 124.800 169.800 125.100 ;
        RECT 170.200 125.100 170.600 125.200 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 170.200 124.800 171.400 125.100 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 166.200 124.100 166.600 124.200 ;
        RECT 165.400 123.800 166.600 124.100 ;
        RECT 164.600 122.800 165.000 123.200 ;
        RECT 163.800 114.800 164.200 115.200 ;
        RECT 163.000 102.800 163.400 103.200 ;
        RECT 161.400 36.800 161.800 37.200 ;
        RECT 161.400 36.200 161.700 36.800 ;
        RECT 161.400 35.800 161.800 36.200 ;
        RECT 151.000 33.800 151.400 34.200 ;
        RECT 151.000 29.200 151.300 33.800 ;
        RECT 151.000 28.800 151.400 29.200 ;
        RECT 161.400 28.800 161.800 29.200 ;
        RECT 151.000 27.100 151.400 27.200 ;
        RECT 151.800 27.100 152.200 27.200 ;
        RECT 151.000 26.800 152.200 27.100 ;
        RECT 161.400 25.200 161.700 28.800 ;
        RECT 163.000 28.200 163.300 102.800 ;
        RECT 163.800 85.200 164.100 114.800 ;
        RECT 163.800 84.800 164.200 85.200 ;
        RECT 164.600 38.200 164.900 122.800 ;
        RECT 175.800 116.200 176.100 152.800 ;
        RECT 179.800 151.800 180.200 152.200 ;
        RECT 179.800 143.200 180.100 151.800 ;
        RECT 180.600 146.200 180.900 152.800 ;
        RECT 180.600 145.800 181.000 146.200 ;
        RECT 179.800 142.800 180.200 143.200 ;
        RECT 178.200 134.800 178.600 135.200 ;
        RECT 176.600 134.100 177.000 134.200 ;
        RECT 177.400 134.100 177.800 134.200 ;
        RECT 176.600 133.800 177.800 134.100 ;
        RECT 175.000 115.800 175.400 116.200 ;
        RECT 175.800 115.800 176.200 116.200 ;
        RECT 175.000 115.200 175.300 115.800 ;
        RECT 166.200 114.800 166.600 115.200 ;
        RECT 175.000 114.800 175.400 115.200 ;
        RECT 166.200 107.200 166.500 114.800 ;
        RECT 176.600 112.800 177.000 113.200 ;
        RECT 166.200 106.800 166.600 107.200 ;
        RECT 171.800 102.800 172.200 103.200 ;
        RECT 171.800 95.200 172.100 102.800 ;
        RECT 171.800 94.800 172.200 95.200 ;
        RECT 176.600 89.200 176.900 112.800 ;
        RECT 176.600 88.800 177.000 89.200 ;
        RECT 174.200 86.800 174.600 87.200 ;
        RECT 171.800 74.800 172.200 75.200 ;
        RECT 173.400 74.800 173.800 75.200 ;
        RECT 171.800 69.200 172.100 74.800 ;
        RECT 167.800 69.100 168.200 69.200 ;
        RECT 167.800 68.800 168.900 69.100 ;
        RECT 168.600 68.200 168.900 68.800 ;
        RECT 171.000 68.800 171.400 69.200 ;
        RECT 171.800 68.800 172.200 69.200 ;
        RECT 168.600 67.800 169.000 68.200 ;
        RECT 171.000 67.200 171.300 68.800 ;
        RECT 171.000 66.800 171.400 67.200 ;
        RECT 172.600 64.800 173.000 65.200 ;
        RECT 163.800 37.800 164.200 38.200 ;
        RECT 164.600 37.800 165.000 38.200 ;
        RECT 163.800 37.200 164.100 37.800 ;
        RECT 163.800 36.800 164.200 37.200 ;
        RECT 167.000 37.100 167.400 37.200 ;
        RECT 167.800 37.100 168.200 37.200 ;
        RECT 167.000 36.800 168.200 37.100 ;
        RECT 163.000 27.800 163.400 28.200 ;
        RECT 166.200 27.100 166.600 27.200 ;
        RECT 167.000 27.100 167.400 27.200 ;
        RECT 166.200 26.800 167.400 27.100 ;
        RECT 161.400 24.800 161.800 25.200 ;
        RECT 172.600 17.200 172.900 64.800 ;
        RECT 173.400 55.200 173.700 74.800 ;
        RECT 174.200 67.200 174.500 86.800 ;
        RECT 178.200 86.200 178.500 134.800 ;
        RECT 179.000 110.800 179.400 111.200 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 177.400 72.800 177.800 73.200 ;
        RECT 174.200 66.800 174.600 67.200 ;
        RECT 175.800 67.100 176.200 67.200 ;
        RECT 176.600 67.100 177.000 67.200 ;
        RECT 175.800 66.800 177.000 67.100 ;
        RECT 177.400 63.200 177.700 72.800 ;
        RECT 177.400 62.800 177.800 63.200 ;
        RECT 178.200 59.200 178.500 85.800 ;
        RECT 179.000 77.200 179.300 110.800 ;
        RECT 179.800 107.200 180.100 142.800 ;
        RECT 180.600 126.200 180.900 145.800 ;
        RECT 183.800 134.200 184.100 157.800 ;
        RECT 183.800 133.800 184.200 134.200 ;
        RECT 180.600 125.800 181.000 126.200 ;
        RECT 180.600 111.200 180.900 125.800 ;
        RECT 182.200 116.100 182.600 116.200 ;
        RECT 183.000 116.100 183.400 116.200 ;
        RECT 182.200 115.800 183.400 116.100 ;
        RECT 180.600 110.800 181.000 111.200 ;
        RECT 179.800 106.800 180.200 107.200 ;
        RECT 180.600 106.800 181.000 107.200 ;
        RECT 179.800 80.200 180.100 106.800 ;
        RECT 180.600 84.200 180.900 106.800 ;
        RECT 182.200 85.200 182.500 115.800 ;
        RECT 183.800 115.100 184.200 115.200 ;
        RECT 184.600 115.100 185.000 115.200 ;
        RECT 183.800 114.800 185.000 115.100 ;
        RECT 183.000 104.800 183.400 105.200 ;
        RECT 183.000 89.200 183.300 104.800 ;
        RECT 185.400 99.200 185.700 185.800 ;
        RECT 201.400 175.200 201.700 199.800 ;
        RECT 201.400 174.800 201.800 175.200 ;
        RECT 187.800 169.800 188.200 170.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 187.000 165.200 187.300 165.800 ;
        RECT 187.000 164.800 187.400 165.200 ;
        RECT 186.200 135.800 186.600 136.200 ;
        RECT 186.200 134.200 186.500 135.800 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 187.800 126.100 188.100 169.800 ;
        RECT 202.200 162.200 202.500 204.800 ;
        RECT 211.000 201.800 211.400 202.200 ;
        RECT 209.400 176.800 209.800 177.200 ;
        RECT 203.000 175.800 203.400 176.200 ;
        RECT 202.200 161.800 202.600 162.200 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 199.000 154.800 199.400 155.200 ;
        RECT 196.600 147.200 196.900 154.800 ;
        RECT 199.000 154.200 199.300 154.800 ;
        RECT 199.000 153.800 199.400 154.200 ;
        RECT 198.200 149.800 198.600 150.200 ;
        RECT 196.600 146.800 197.000 147.200 ;
        RECT 195.800 132.800 196.200 133.200 ;
        RECT 190.200 130.800 190.600 131.200 ;
        RECT 190.200 129.200 190.500 130.800 ;
        RECT 190.200 128.800 190.600 129.200 ;
        RECT 188.600 126.100 189.000 126.200 ;
        RECT 187.800 125.800 189.000 126.100 ;
        RECT 191.000 125.800 191.400 126.200 ;
        RECT 188.600 106.200 188.900 125.800 ;
        RECT 191.000 125.200 191.300 125.800 ;
        RECT 191.000 124.800 191.400 125.200 ;
        RECT 189.400 119.800 189.800 120.200 ;
        RECT 188.600 105.800 189.000 106.200 ;
        RECT 186.200 103.800 186.600 104.200 ;
        RECT 185.400 98.800 185.800 99.200 ;
        RECT 185.400 94.800 185.800 95.200 ;
        RECT 184.600 90.100 185.000 90.200 ;
        RECT 183.800 89.800 185.000 90.100 ;
        RECT 183.000 88.800 183.400 89.200 ;
        RECT 182.200 84.800 182.600 85.200 ;
        RECT 180.600 83.800 181.000 84.200 ;
        RECT 179.800 79.800 180.200 80.200 ;
        RECT 179.000 76.800 179.400 77.200 ;
        RECT 183.800 73.200 184.100 89.800 ;
        RECT 183.800 72.800 184.200 73.200 ;
        RECT 183.800 67.200 184.100 72.800 ;
        RECT 185.400 72.200 185.700 94.800 ;
        RECT 186.200 85.200 186.500 103.800 ;
        RECT 187.000 95.100 187.400 95.200 ;
        RECT 187.800 95.100 188.200 95.200 ;
        RECT 187.000 94.800 188.200 95.100 ;
        RECT 186.200 84.800 186.600 85.200 ;
        RECT 186.200 74.800 186.600 75.200 ;
        RECT 185.400 71.800 185.800 72.200 ;
        RECT 183.800 66.800 184.200 67.200 ;
        RECT 178.200 58.800 178.600 59.200 ;
        RECT 183.800 56.200 184.100 66.800 ;
        RECT 186.200 65.200 186.500 74.800 ;
        RECT 186.200 64.800 186.600 65.200 ;
        RECT 183.800 55.800 184.200 56.200 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 185.400 44.100 185.800 44.200 ;
        RECT 184.600 43.800 185.800 44.100 ;
        RECT 184.600 24.200 184.900 43.800 ;
        RECT 184.600 23.800 185.000 24.200 ;
        RECT 187.000 19.200 187.300 94.800 ;
        RECT 187.800 76.800 188.200 77.200 ;
        RECT 187.800 75.200 188.100 76.800 ;
        RECT 187.800 74.800 188.200 75.200 ;
        RECT 189.400 66.200 189.700 119.800 ;
        RECT 190.200 89.800 190.600 90.200 ;
        RECT 190.200 77.200 190.500 89.800 ;
        RECT 195.800 85.200 196.100 132.800 ;
        RECT 196.600 131.200 196.900 146.800 ;
        RECT 198.200 136.200 198.500 149.800 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 198.200 135.800 198.600 136.200 ;
        RECT 197.400 131.200 197.700 135.800 ;
        RECT 196.600 130.800 197.000 131.200 ;
        RECT 197.400 130.800 197.800 131.200 ;
        RECT 197.400 95.100 197.800 95.200 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 197.400 94.800 198.600 95.100 ;
        RECT 195.800 84.800 196.200 85.200 ;
        RECT 190.200 76.800 190.600 77.200 ;
        RECT 189.400 65.800 189.800 66.200 ;
        RECT 194.200 64.100 194.600 64.200 ;
        RECT 193.400 63.800 194.600 64.100 ;
        RECT 190.200 50.800 190.600 51.200 ;
        RECT 190.200 34.200 190.500 50.800 ;
        RECT 190.200 33.800 190.600 34.200 ;
        RECT 193.400 31.200 193.700 63.800 ;
        RECT 195.800 41.200 196.100 84.800 ;
        RECT 199.000 74.200 199.300 153.800 ;
        RECT 202.200 121.800 202.600 122.200 ;
        RECT 202.200 96.200 202.500 121.800 ;
        RECT 202.200 95.800 202.600 96.200 ;
        RECT 199.800 93.800 200.200 94.200 ;
        RECT 199.800 93.200 200.100 93.800 ;
        RECT 199.800 92.800 200.200 93.200 ;
        RECT 201.400 75.800 201.800 76.200 ;
        RECT 199.000 73.800 199.400 74.200 ;
        RECT 201.400 55.200 201.700 75.800 ;
        RECT 203.000 75.200 203.300 175.800 ;
        RECT 207.000 157.800 207.400 158.200 ;
        RECT 207.000 148.200 207.300 157.800 ;
        RECT 207.800 153.800 208.200 154.200 ;
        RECT 207.000 147.800 207.400 148.200 ;
        RECT 207.000 135.100 207.400 135.200 ;
        RECT 207.800 135.100 208.100 153.800 ;
        RECT 207.000 134.800 208.100 135.100 ;
        RECT 207.000 133.800 207.400 134.200 ;
        RECT 204.600 113.800 205.000 114.200 ;
        RECT 204.600 93.200 204.900 113.800 ;
        RECT 207.000 107.200 207.300 133.800 ;
        RECT 207.800 129.800 208.200 130.200 ;
        RECT 207.800 109.200 208.100 129.800 ;
        RECT 207.800 108.800 208.200 109.200 ;
        RECT 207.000 106.800 207.400 107.200 ;
        RECT 207.000 100.800 207.400 101.200 ;
        RECT 205.400 95.100 205.800 95.200 ;
        RECT 206.200 95.100 206.600 95.200 ;
        RECT 205.400 94.800 206.600 95.100 ;
        RECT 204.600 92.800 205.000 93.200 ;
        RECT 204.600 75.200 204.900 92.800 ;
        RECT 203.000 74.800 203.400 75.200 ;
        RECT 204.600 74.800 205.000 75.200 ;
        RECT 203.000 71.800 203.400 72.200 ;
        RECT 201.400 54.800 201.800 55.200 ;
        RECT 201.400 48.200 201.700 54.800 ;
        RECT 201.400 47.800 201.800 48.200 ;
        RECT 200.600 46.800 201.000 47.200 ;
        RECT 195.800 40.800 196.200 41.200 ;
        RECT 193.400 30.800 193.800 31.200 ;
        RECT 193.400 23.200 193.700 30.800 ;
        RECT 200.600 26.200 200.900 46.800 ;
        RECT 203.000 45.200 203.300 71.800 ;
        RECT 207.000 56.200 207.300 100.800 ;
        RECT 207.800 86.200 208.100 108.800 ;
        RECT 207.800 85.800 208.200 86.200 ;
        RECT 207.000 55.800 207.400 56.200 ;
        RECT 207.800 46.200 208.100 85.800 ;
        RECT 209.400 65.100 209.700 176.800 ;
        RECT 210.200 155.800 210.600 156.200 ;
        RECT 210.200 127.200 210.500 155.800 ;
        RECT 211.000 146.200 211.300 201.800 ;
        RECT 213.400 155.200 213.700 205.800 ;
        RECT 217.400 204.800 217.800 205.200 ;
        RECT 217.400 176.200 217.700 204.800 ;
        RECT 219.000 191.800 219.400 192.200 ;
        RECT 215.000 175.800 215.400 176.200 ;
        RECT 217.400 175.800 217.800 176.200 ;
        RECT 213.400 154.800 213.800 155.200 ;
        RECT 214.200 154.800 214.600 155.200 ;
        RECT 214.200 154.200 214.500 154.800 ;
        RECT 214.200 153.800 214.600 154.200 ;
        RECT 215.000 152.200 215.300 175.800 ;
        RECT 215.000 151.800 215.400 152.200 ;
        RECT 216.600 149.800 217.000 150.200 ;
        RECT 211.000 145.800 211.400 146.200 ;
        RECT 211.000 137.800 211.400 138.200 ;
        RECT 210.200 126.800 210.600 127.200 ;
        RECT 211.000 116.200 211.300 137.800 ;
        RECT 211.000 115.800 211.400 116.200 ;
        RECT 211.000 105.200 211.300 115.800 ;
        RECT 216.600 115.200 216.900 149.800 ;
        RECT 216.600 114.800 217.000 115.200 ;
        RECT 211.000 104.800 211.400 105.200 ;
        RECT 210.200 65.100 210.600 65.200 ;
        RECT 209.400 64.800 210.600 65.100 ;
        RECT 211.000 63.200 211.300 104.800 ;
        RECT 211.000 62.800 211.400 63.200 ;
        RECT 207.800 45.800 208.200 46.200 ;
        RECT 203.000 44.800 203.400 45.200 ;
        RECT 203.000 36.200 203.300 44.800 ;
        RECT 203.000 35.800 203.400 36.200 ;
        RECT 204.600 27.800 205.000 28.200 ;
        RECT 204.600 26.200 204.900 27.800 ;
        RECT 200.600 25.800 201.000 26.200 ;
        RECT 204.600 25.800 205.000 26.200 ;
        RECT 193.400 22.800 193.800 23.200 ;
        RECT 187.000 18.800 187.400 19.200 ;
        RECT 172.600 16.800 173.000 17.200 ;
        RECT 149.400 10.800 149.800 11.200 ;
        RECT 200.600 9.200 200.900 25.800 ;
        RECT 217.400 14.200 217.700 175.800 ;
        RECT 218.200 133.800 218.600 134.200 ;
        RECT 218.200 127.200 218.500 133.800 ;
        RECT 218.200 126.800 218.600 127.200 ;
        RECT 219.000 114.200 219.300 191.800 ;
        RECT 220.600 155.100 221.000 155.200 ;
        RECT 221.400 155.100 221.800 155.200 ;
        RECT 220.600 154.800 221.800 155.100 ;
        RECT 220.600 143.800 221.000 144.200 ;
        RECT 219.000 113.800 219.400 114.200 ;
        RECT 219.000 84.800 219.400 85.200 ;
        RECT 219.000 73.200 219.300 84.800 ;
        RECT 219.000 72.800 219.400 73.200 ;
        RECT 219.000 48.800 219.400 49.200 ;
        RECT 219.000 25.200 219.300 48.800 ;
        RECT 220.600 33.200 220.900 143.800 ;
        RECT 222.200 110.200 222.500 206.800 ;
        RECT 222.200 109.800 222.600 110.200 ;
        RECT 223.000 85.200 223.300 206.800 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 224.600 144.200 224.900 205.800 ;
        RECT 228.600 204.800 229.000 205.200 ;
        RECT 225.400 202.100 225.800 202.200 ;
        RECT 225.400 201.800 226.500 202.100 ;
        RECT 224.600 143.800 225.000 144.200 ;
        RECT 225.400 123.800 225.800 124.200 ;
        RECT 223.000 84.800 223.400 85.200 ;
        RECT 224.600 65.800 225.000 66.200 ;
        RECT 220.600 32.800 221.000 33.200 ;
        RECT 219.000 24.800 219.400 25.200 ;
        RECT 224.600 22.200 224.900 65.800 ;
        RECT 225.400 26.200 225.700 123.800 ;
        RECT 226.200 101.200 226.500 201.800 ;
        RECT 227.800 110.800 228.200 111.200 ;
        RECT 226.200 100.800 226.600 101.200 ;
        RECT 227.800 90.200 228.100 110.800 ;
        RECT 228.600 108.200 228.900 204.800 ;
        RECT 228.600 107.800 229.000 108.200 ;
        RECT 227.800 89.800 228.200 90.200 ;
        RECT 228.600 53.800 229.000 54.200 ;
        RECT 226.200 35.800 226.600 36.200 ;
        RECT 225.400 25.800 225.800 26.200 ;
        RECT 224.600 21.800 225.000 22.200 ;
        RECT 226.200 16.200 226.500 35.800 ;
        RECT 228.600 27.200 228.900 53.800 ;
        RECT 228.600 26.800 229.000 27.200 ;
        RECT 226.200 15.800 226.600 16.200 ;
        RECT 217.400 13.800 217.800 14.200 ;
        RECT 23.800 8.800 24.200 9.200 ;
        RECT 85.400 8.800 85.800 9.200 ;
        RECT 200.600 8.800 201.000 9.200 ;
        RECT 79.000 7.800 79.400 8.200 ;
        RECT 37.400 7.100 37.800 7.200 ;
        RECT 38.200 7.100 38.600 7.200 ;
        RECT 37.400 6.800 38.600 7.100 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 45.400 6.800 46.600 7.100 ;
        RECT 79.000 5.200 79.300 7.800 ;
        RECT 85.400 6.200 85.700 8.800 ;
        RECT 85.400 5.800 85.800 6.200 ;
        RECT 79.000 4.800 79.400 5.200 ;
      LAYER via4 ;
        RECT 28.600 205.800 29.000 206.200 ;
        RECT 58.200 204.800 58.600 205.200 ;
        RECT 14.200 125.800 14.600 126.200 ;
        RECT 31.000 146.800 31.400 147.200 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 33.400 45.800 33.800 46.200 ;
        RECT 33.400 34.800 33.800 35.200 ;
        RECT 67.800 165.800 68.200 166.200 ;
        RECT 70.200 114.800 70.600 115.200 ;
        RECT 63.000 92.800 63.400 93.200 ;
        RECT 52.600 87.800 53.000 88.200 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 57.400 33.800 57.800 34.200 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 101.400 164.800 101.800 165.200 ;
        RECT 74.200 36.800 74.600 37.200 ;
        RECT 103.800 124.800 104.200 125.200 ;
        RECT 99.000 41.800 99.400 42.200 ;
        RECT 110.200 116.800 110.600 117.200 ;
        RECT 115.000 74.800 115.400 75.200 ;
        RECT 120.600 125.800 121.000 126.200 ;
        RECT 126.200 164.800 126.600 165.200 ;
        RECT 130.200 173.800 130.600 174.200 ;
        RECT 128.600 147.800 129.000 148.200 ;
        RECT 139.000 134.800 139.400 135.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 150.200 145.800 150.600 146.200 ;
        RECT 119.800 56.800 120.200 57.200 ;
        RECT 123.800 56.800 124.200 57.200 ;
        RECT 126.200 92.800 126.600 93.200 ;
        RECT 136.600 104.800 137.000 105.200 ;
        RECT 143.800 126.800 144.200 127.200 ;
        RECT 175.800 187.800 176.200 188.200 ;
        RECT 158.200 105.800 158.600 106.200 ;
        RECT 153.400 88.800 153.800 89.200 ;
        RECT 159.000 68.800 159.400 69.200 ;
        RECT 179.000 164.800 179.400 165.200 ;
        RECT 181.400 153.800 181.800 154.200 ;
        RECT 171.000 124.800 171.400 125.200 ;
        RECT 151.800 26.800 152.200 27.200 ;
        RECT 167.800 36.800 168.200 37.200 ;
        RECT 176.600 66.800 177.000 67.200 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 221.400 154.800 221.800 155.200 ;
        RECT 38.200 6.800 38.600 7.200 ;
      LAYER metal5 ;
        RECT 28.600 206.100 29.000 206.200 ;
        RECT 32.600 206.100 33.000 206.200 ;
        RECT 28.600 205.800 33.000 206.100 ;
        RECT 30.200 205.100 30.600 205.200 ;
        RECT 58.200 205.100 58.600 205.200 ;
        RECT 75.800 205.100 76.200 205.200 ;
        RECT 30.200 204.800 76.200 205.100 ;
        RECT 18.200 192.100 18.600 192.200 ;
        RECT 59.000 192.100 59.400 192.200 ;
        RECT 18.200 191.800 59.400 192.100 ;
        RECT 175.800 188.100 176.200 188.200 ;
        RECT 178.200 188.100 178.600 188.200 ;
        RECT 175.800 187.800 178.600 188.100 ;
        RECT 59.800 184.100 60.200 184.200 ;
        RECT 95.000 184.100 95.400 184.200 ;
        RECT 155.000 184.100 155.400 184.200 ;
        RECT 59.800 183.800 155.400 184.100 ;
        RECT 71.000 174.100 71.400 174.200 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 152.600 174.100 153.000 174.200 ;
        RECT 71.000 173.800 153.000 174.100 ;
        RECT 67.800 166.100 68.200 166.200 ;
        RECT 155.800 166.100 156.200 166.200 ;
        RECT 67.800 165.800 156.200 166.100 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 101.400 165.100 101.800 165.200 ;
        RECT 126.200 165.100 126.600 165.200 ;
        RECT 101.400 164.800 126.600 165.100 ;
        RECT 179.000 165.100 179.400 165.200 ;
        RECT 187.000 165.100 187.300 165.800 ;
        RECT 179.000 164.800 187.300 165.100 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 199.000 155.100 199.400 155.200 ;
        RECT 147.800 154.800 199.400 155.100 ;
        RECT 214.200 155.100 214.600 155.200 ;
        RECT 221.400 155.100 221.800 155.200 ;
        RECT 214.200 154.800 221.800 155.100 ;
        RECT 118.200 154.100 118.600 154.200 ;
        RECT 181.400 154.100 181.800 154.200 ;
        RECT 118.200 153.800 181.800 154.100 ;
        RECT 87.000 148.100 87.400 148.200 ;
        RECT 128.600 148.100 129.000 148.200 ;
        RECT 87.000 147.800 129.000 148.100 ;
        RECT 31.000 147.100 31.400 147.200 ;
        RECT 79.000 147.100 79.400 147.200 ;
        RECT 31.000 146.800 79.400 147.100 ;
        RECT 45.400 146.100 45.800 146.200 ;
        RECT 130.200 146.100 130.600 146.200 ;
        RECT 45.400 145.800 130.600 146.100 ;
        RECT 135.000 146.100 135.400 146.200 ;
        RECT 142.200 146.100 142.600 146.200 ;
        RECT 135.000 145.800 142.600 146.100 ;
        RECT 150.200 146.100 150.600 146.200 ;
        RECT 180.600 146.100 181.000 146.200 ;
        RECT 150.200 145.800 181.000 146.100 ;
        RECT 102.200 145.100 102.600 145.200 ;
        RECT 149.400 145.100 149.800 145.200 ;
        RECT 102.200 144.800 149.800 145.100 ;
        RECT 124.600 142.100 125.000 142.200 ;
        RECT 153.400 142.100 153.800 142.200 ;
        RECT 124.600 141.800 153.800 142.100 ;
        RECT 62.200 136.100 62.600 136.200 ;
        RECT 140.600 136.100 141.000 136.200 ;
        RECT 62.200 135.800 141.000 136.100 ;
        RECT 80.600 135.100 81.000 135.200 ;
        RECT 91.800 135.100 92.200 135.200 ;
        RECT 80.600 134.800 92.200 135.100 ;
        RECT 110.200 135.100 110.600 135.200 ;
        RECT 139.000 135.100 139.400 135.200 ;
        RECT 145.400 135.100 145.800 135.200 ;
        RECT 110.200 134.800 136.900 135.100 ;
        RECT 139.000 134.800 145.800 135.100 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 176.600 134.100 177.000 134.200 ;
        RECT 186.200 134.100 186.600 134.200 ;
        RECT 176.600 133.800 186.600 134.100 ;
        RECT 114.200 127.800 114.600 128.200 ;
        RECT 114.200 127.100 114.500 127.800 ;
        RECT 143.800 127.100 144.200 127.200 ;
        RECT 114.200 126.800 144.200 127.100 ;
        RECT 14.200 126.100 14.600 126.200 ;
        RECT 67.000 126.100 67.400 126.200 ;
        RECT 14.200 125.800 67.400 126.100 ;
        RECT 111.000 126.100 111.400 126.200 ;
        RECT 120.600 126.100 121.000 126.200 ;
        RECT 111.000 125.800 121.000 126.100 ;
        RECT 103.800 125.100 104.200 125.200 ;
        RECT 116.600 125.100 117.000 125.200 ;
        RECT 103.800 124.800 117.000 125.100 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 191.000 125.100 191.400 125.200 ;
        RECT 171.000 124.800 191.400 125.100 ;
        RECT 113.400 124.100 113.800 124.200 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 113.400 123.800 165.800 124.100 ;
        RECT 110.200 117.100 110.600 117.200 ;
        RECT 155.800 117.100 156.200 117.200 ;
        RECT 110.200 116.800 156.200 117.100 ;
        RECT 86.200 116.100 86.600 116.200 ;
        RECT 127.800 116.100 128.200 116.200 ;
        RECT 86.200 115.800 128.200 116.100 ;
        RECT 160.600 116.100 161.000 116.200 ;
        RECT 182.200 116.100 182.600 116.200 ;
        RECT 160.600 115.800 182.600 116.100 ;
        RECT 47.800 115.100 48.200 115.200 ;
        RECT 70.200 115.100 70.600 115.200 ;
        RECT 84.600 115.100 85.000 115.200 ;
        RECT 103.000 115.100 103.400 115.200 ;
        RECT 119.800 115.100 120.200 115.200 ;
        RECT 47.800 114.800 120.200 115.100 ;
        RECT 175.000 115.100 175.400 115.200 ;
        RECT 183.800 115.100 184.200 115.200 ;
        RECT 175.000 114.800 184.200 115.100 ;
        RECT 116.600 114.100 117.000 114.200 ;
        RECT 78.200 113.800 117.000 114.100 ;
        RECT 78.200 113.200 78.500 113.800 ;
        RECT 78.200 112.800 78.600 113.200 ;
        RECT 102.200 113.100 102.600 113.200 ;
        RECT 129.400 113.100 129.800 113.200 ;
        RECT 102.200 112.800 129.800 113.100 ;
        RECT 19.800 107.100 20.200 107.200 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 19.800 106.800 25.000 107.100 ;
        RECT 121.400 106.100 121.800 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 121.400 105.800 158.600 106.100 ;
        RECT 136.600 105.100 137.000 105.200 ;
        RECT 156.600 105.100 157.000 105.200 ;
        RECT 136.600 104.800 157.000 105.100 ;
        RECT 99.800 104.100 100.200 104.200 ;
        RECT 146.200 104.100 146.600 104.200 ;
        RECT 99.800 103.800 146.600 104.100 ;
        RECT 101.400 103.100 101.800 103.200 ;
        RECT 171.800 103.100 172.200 103.200 ;
        RECT 101.400 102.800 172.200 103.100 ;
        RECT 105.400 98.100 105.800 98.200 ;
        RECT 108.600 98.100 109.000 98.200 ;
        RECT 105.400 97.800 109.000 98.100 ;
        RECT 152.600 95.800 153.000 96.200 ;
        RECT 77.400 95.100 77.800 95.200 ;
        RECT 152.600 95.100 152.900 95.800 ;
        RECT 77.400 94.800 152.900 95.100 ;
        RECT 154.200 95.100 154.600 95.200 ;
        RECT 187.000 95.100 187.400 95.200 ;
        RECT 154.200 94.800 187.400 95.100 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 205.400 95.100 205.800 95.200 ;
        RECT 198.200 94.800 205.800 95.100 ;
        RECT 157.400 94.100 157.800 94.200 ;
        RECT 157.400 93.800 200.100 94.100 ;
        RECT 199.800 93.200 200.100 93.800 ;
        RECT 63.000 93.100 63.400 93.200 ;
        RECT 126.200 93.100 126.600 93.200 ;
        RECT 63.000 92.800 126.600 93.100 ;
        RECT 199.800 92.800 200.200 93.200 ;
        RECT 75.800 89.100 76.200 89.200 ;
        RECT 153.400 89.100 153.800 89.200 ;
        RECT 75.800 88.800 153.800 89.100 ;
        RECT 52.600 88.100 53.000 88.200 ;
        RECT 156.600 88.100 157.000 88.200 ;
        RECT 52.600 87.800 157.000 88.100 ;
        RECT 152.600 87.100 153.000 87.200 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 152.600 86.800 159.400 87.100 ;
        RECT 115.000 75.100 115.400 75.200 ;
        RECT 171.800 75.100 172.200 75.200 ;
        RECT 115.000 74.800 172.200 75.100 ;
        RECT 64.600 74.100 65.000 74.200 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 64.600 73.800 119.400 74.100 ;
        RECT 65.400 73.100 65.800 73.200 ;
        RECT 106.200 73.100 106.600 73.200 ;
        RECT 65.400 72.800 106.600 73.100 ;
        RECT 102.200 71.100 102.600 71.200 ;
        RECT 116.600 71.100 117.000 71.200 ;
        RECT 102.200 70.800 117.000 71.100 ;
        RECT 148.600 69.800 149.000 70.200 ;
        RECT 99.800 68.800 100.200 69.200 ;
        RECT 112.600 68.800 113.000 69.200 ;
        RECT 148.600 69.100 148.900 69.800 ;
        RECT 159.000 69.100 159.400 69.200 ;
        RECT 148.600 68.800 159.400 69.100 ;
        RECT 99.800 68.100 100.100 68.800 ;
        RECT 112.600 68.100 112.900 68.800 ;
        RECT 99.800 67.800 112.900 68.100 ;
        RECT 154.200 68.100 154.600 68.200 ;
        RECT 168.600 68.100 169.000 68.200 ;
        RECT 154.200 67.800 169.000 68.100 ;
        RECT 75.800 67.100 76.200 67.200 ;
        RECT 155.000 67.100 155.400 67.200 ;
        RECT 75.800 66.800 155.400 67.100 ;
        RECT 171.000 67.100 171.400 67.200 ;
        RECT 176.600 67.100 177.000 67.200 ;
        RECT 171.000 66.800 177.000 67.100 ;
        RECT 119.800 57.100 120.200 57.200 ;
        RECT 123.800 57.100 124.200 57.200 ;
        RECT 119.800 56.800 124.200 57.100 ;
        RECT 28.600 46.100 29.000 46.200 ;
        RECT 33.400 46.100 33.800 46.200 ;
        RECT 28.600 45.800 33.800 46.100 ;
        RECT 99.000 42.100 99.400 42.200 ;
        RECT 143.000 42.100 143.400 42.200 ;
        RECT 99.000 41.800 143.400 42.100 ;
        RECT 74.200 37.100 74.600 37.200 ;
        RECT 117.400 37.100 117.800 37.200 ;
        RECT 74.200 36.800 117.800 37.100 ;
        RECT 163.800 37.100 164.200 37.200 ;
        RECT 167.800 37.100 168.200 37.200 ;
        RECT 163.800 36.800 168.200 37.100 ;
        RECT 49.400 36.100 49.800 36.200 ;
        RECT 161.400 36.100 161.800 36.200 ;
        RECT 49.400 35.800 161.800 36.100 ;
        RECT 33.400 35.100 33.800 35.200 ;
        RECT 91.000 35.100 91.400 35.200 ;
        RECT 33.400 34.800 91.400 35.100 ;
        RECT 57.400 34.100 57.800 34.200 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 57.400 33.800 104.200 34.100 ;
        RECT 75.000 33.100 75.400 33.200 ;
        RECT 117.400 33.100 117.800 33.200 ;
        RECT 75.000 32.800 117.800 33.100 ;
        RECT 101.400 29.100 101.800 29.200 ;
        RECT 151.000 29.100 151.400 29.200 ;
        RECT 101.400 28.800 151.400 29.100 ;
        RECT 112.600 28.100 113.000 28.200 ;
        RECT 204.600 28.100 205.000 28.200 ;
        RECT 112.600 27.800 205.000 28.100 ;
        RECT 151.800 27.100 152.200 27.200 ;
        RECT 166.200 27.100 166.600 27.200 ;
        RECT 151.800 26.800 166.600 27.100 ;
        RECT 43.800 15.100 44.200 15.200 ;
        RECT 115.000 15.100 115.400 15.200 ;
        RECT 43.800 14.800 115.400 15.100 ;
        RECT 38.200 7.100 38.600 7.200 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 38.200 6.800 45.800 7.100 ;
  END
END ram32_sdram_3split
END LIBRARY

