* NGSPICE file created from ram32_sdram_2split.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt ram32_sdram_2split vdd gnd en rw clk ras cas datain[0] datain[1] datain[2]
+ datain[3] datain[4] datain[5] datain[6] datain[7] address[0] address[1] address[2]
+ address[3] address[4] dataout[0] dataout[1] dataout[2] dataout[3] dataout[4] dataout[5]
+ dataout[6] dataout[7]
XFILL_23_3_0 gnd vdd FILL
XMUX2X1_17 INVX1_17/Y BUFX4_57/Y MUX2X1_17/S gnd MUX2X1_17/Y vdd MUX2X1
XFILL_14_3_0 gnd vdd FILL
XMUX2X1_28 INVX1_28/Y BUFX4_27/Y MUX2X1_27/S gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_39 INVX1_39/Y BUFX4_22/Y MUX2X1_39/S gnd MUX2X1_39/Y vdd MUX2X1
XNAND2X1_43 MUX2X1_178/A NAND3X1_4/Y gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_10 MUX2X1_76/A OAI21X1_9/B gnd OAI21X1_9/C vdd NAND2X1
XNAND2X1_32 NAND2X1_32/A OAI21X1_25/B gnd NAND2X1_32/Y vdd NAND2X1
XAOI22X1_30 MUX2X1_233/Y AND2X2_3/A AND2X2_2/B AOI22X1_30/D gnd AOI22X1_30/Y vdd AOI22X1
XNAND2X1_54 AND2X2_2/B NOR2X1_1/Y gnd NAND2X1_56/B vdd NAND2X1
XNAND2X1_87 MUX2X1_153/B NAND2X1_88/B gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_98 NAND2X1_98/A NAND3X1_7/Y gnd NAND2X1_98/Y vdd NAND2X1
XNAND2X1_76 MUX2X1_169/A NAND3X1_6/Y gnd OAI21X1_69/C vdd NAND2X1
XNAND2X1_65 MUX2X1_88/A NAND2X1_64/B gnd OAI21X1_58/C vdd NAND2X1
XNAND2X1_21 MUX2X1_99/B NAND3X1_3/Y gnd NAND2X1_21/Y vdd NAND2X1
XFILL_20_1_0 gnd vdd FILL
XOAI21X1_19 BUFX4_10/Y NAND3X1_3/Y NAND2X1_22/Y gnd OAI21X1_19/Y vdd OAI21X1
XFILL_19_2_0 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XDFFPOSX1_147 MUX2X1_232/A CLKBUF1_43/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 INVX1_19/A CLKBUF1_5/A MUX2X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_169 INVX1_30/A CLKBUF1_19/Y MUX2X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 MUX2X1_139/A CLKBUF1_25/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 NAND2X1_59/A CLKBUF1_21/Y OAI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 MUX2X1_202/A CLKBUF1_46/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_125 MUX2X1_90/A CLKBUF1_4/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XMUX2X1_245 MUX2X1_245/A MUX2X1_245/B BUFX4_18/Y gnd AOI22X1_32/A vdd MUX2X1
XMUX2X1_234 NOR2X1_19/A MUX2X1_234/B BUFX4_38/Y gnd MUX2X1_236/B vdd MUX2X1
XMUX2X1_256 INVX1_66/Y BUFX4_44/Y MUX2X1_249/S gnd MUX2X1_256/Y vdd MUX2X1
XMUX2X1_223 NAND2X1_98/A MUX2X1_223/B BUFX4_31/Y gnd MUX2X1_223/Y vdd MUX2X1
XMUX2X1_201 MUX2X1_201/A NAND2X1_89/A BUFX4_38/Y gnd MUX2X1_201/Y vdd MUX2X1
XMUX2X1_212 MUX2X1_212/A MUX2X1_210/Y BUFX4_15/Y gnd AOI22X1_26/D vdd MUX2X1
XBUFX4_41 INVX8_10/Y gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 BUFX4_34/A gnd BUFX4_30/Y vdd BUFX4
XBUFX4_52 INVX8_4/Y gnd BUFX4_52/Y vdd BUFX4
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XINVX8_11 INVX8_11/A gnd INVX8_11/Y vdd INVX8
XFILL_0_0_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XMUX2X1_29 INVX1_29/Y MUX2X1_5/B MUX2X1_27/S gnd MUX2X1_29/Y vdd MUX2X1
XMUX2X1_18 INVX1_18/Y MUX2X1_2/B MUX2X1_17/S gnd MUX2X1_18/Y vdd MUX2X1
XNAND2X1_88 NAND2X1_88/A NAND2X1_88/B gnd OAI21X1_78/C vdd NAND2X1
XNAND2X1_22 MUX2X1_123/B NAND3X1_3/Y gnd NAND2X1_22/Y vdd NAND2X1
XNAND2X1_66 MUX2X1_112/A NAND2X1_64/B gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_77 MUX2X1_193/A NAND3X1_6/Y gnd NAND2X1_77/Y vdd NAND2X1
XAOI22X1_1 AOI22X1_1/A INVX8_11/Y INVX8_1/Y AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_55 MUX2X1_66/B NAND2X1_56/B gnd OAI21X1_49/C vdd NAND2X1
XFILL_14_3_1 gnd vdd FILL
XNAND2X1_99 MUX2X1_247/A NAND3X1_7/Y gnd NAND2X1_99/Y vdd NAND2X1
XNAND2X1_33 MUX2X1_139/A OAI21X1_25/B gnd OAI21X1_28/C vdd NAND2X1
XNAND2X1_44 MUX2X1_202/A NAND3X1_4/Y gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_11 MUX2X1_100/A OAI21X1_9/B gnd OAI21X1_10/C vdd NAND2X1
XAOI22X1_31 AOI22X1_31/A INVX1_49/A INVX8_2/Y MUX2X1_242/Y gnd AOI22X1_31/Y vdd AOI22X1
XAOI22X1_20 AOI22X1_20/A AND2X2_4/B AND2X2_1/B MUX2X1_176/Y gnd AOI22X1_20/Y vdd AOI22X1
XFILL_20_1_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XDFFPOSX1_137 MUX2X1_186/B CLKBUF1_17/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_115 MUX2X1_226/A CLKBUF1_44/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 NOR2X1_14/A CLKBUF1_5/A AOI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 MUX2X1_73/A CLKBUF1_37/Y OAI21X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 MUX2X1_163/A CLKBUF1_21/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_159 INVX1_20/A CLKBUF1_2/A MUX2X1_20/Y gnd vdd DFFPOSX1
XMUX2X1_235 MUX2X1_235/A MUX2X1_235/B BUFX4_39/Y gnd MUX2X1_235/Y vdd MUX2X1
XMUX2X1_246 NOR2X1_9/A NAND2X1_8/A BUFX4_35/Y gnd MUX2X1_248/B vdd MUX2X1
XMUX2X1_213 INVX1_47/A INVX1_39/A BUFX4_35/Y gnd MUX2X1_213/Y vdd MUX2X1
XMUX2X1_224 MUX2X1_223/Y MUX2X1_222/Y BUFX4_11/Y gnd MUX2X1_224/Y vdd MUX2X1
XMUX2X1_202 MUX2X1_202/A MUX2X1_202/B BUFX4_39/Y gnd MUX2X1_202/Y vdd MUX2X1
XBUFX4_42 INVX8_10/Y gnd BUFX4_42/Y vdd BUFX4
XBUFX4_31 BUFX4_34/A gnd BUFX4_31/Y vdd BUFX4
XBUFX4_20 INVX8_9/Y gnd MUX2X1_7/B vdd BUFX4
XBUFX4_53 INVX8_4/Y gnd MUX2X1_2/B vdd BUFX4
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_12 MUX2X1_124/A OAI21X1_9/B gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_56 MUX2X1_90/B NAND2X1_56/B gnd OAI21X1_50/C vdd NAND2X1
XNAND2X1_45 MUX2X1_226/A NAND3X1_4/Y gnd NAND2X1_45/Y vdd NAND2X1
XAOI22X1_2 MUX2X1_65/Y AND2X2_3/A AND2X2_2/B AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XMUX2X1_19 INVX1_19/Y BUFX4_6/Y MUX2X1_17/S gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_67 MUX2X1_136/A NAND2X1_64/B gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_23 NAND2X1_23/A NAND3X1_3/Y gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_78 MUX2X1_217/A NAND3X1_6/Y gnd NAND2X1_78/Y vdd NAND2X1
XNAND2X1_89 NAND2X1_89/A NAND2X1_88/B gnd OAI21X1_79/C vdd NAND2X1
XNAND2X1_34 MUX2X1_163/A OAI21X1_25/B gnd NAND2X1_34/Y vdd NAND2X1
XAOI22X1_21 AOI22X1_21/A INVX8_11/Y INVX8_1/Y AOI22X1_21/D gnd AOI22X1_21/Y vdd AOI22X1
XAOI22X1_32 AOI22X1_32/A AND2X2_4/B AND2X2_1/B MUX2X1_248/Y gnd AOI22X1_32/Y vdd AOI22X1
XAOI22X1_10 AOI22X1_10/A AND2X2_3/A AND2X2_2/B AOI22X1_10/D gnd AOI22X1_10/Y vdd AOI22X1
XDFFPOSX1_116 MUX2X1_67/B CLKBUF1_40/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 MUX2X1_187/A CLKBUF1_18/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NOR2X1_15/A CLKBUF1_5/A AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 MUX2X1_210/B CLKBUF1_16/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 MUX2X1_97/A CLKBUF1_35/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XMUX2X1_225 MUX2X1_225/A NAND2X1_90/A BUFX4_32/Y gnd MUX2X1_227/B vdd MUX2X1
XMUX2X1_236 MUX2X1_235/Y MUX2X1_236/B BUFX4_15/Y gnd AOI22X1_30/D vdd MUX2X1
XMUX2X1_247 MUX2X1_247/A MUX2X1_247/B BUFX4_36/Y gnd MUX2X1_247/Y vdd MUX2X1
XMUX2X1_214 INVX1_56/A NOR2X1_38/A BUFX4_36/Y gnd MUX2X1_215/A vdd MUX2X1
XMUX2X1_203 MUX2X1_202/Y MUX2X1_201/Y BUFX4_12/Y gnd AOI22X1_25/A vdd MUX2X1
XBUFX4_43 INVX8_10/Y gnd BUFX4_43/Y vdd BUFX4
XBUFX4_10 INVX8_5/Y gnd BUFX4_10/Y vdd BUFX4
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XBUFX4_32 BUFX4_34/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_21 INVX8_9/Y gnd BUFX4_21/Y vdd BUFX4
XBUFX4_54 INVX8_4/Y gnd BUFX4_54/Y vdd BUFX4
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_1_3_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_160 BUFX4_40/Y NAND3X1_11/Y OAI21X1_160/C gnd DFFPOSX1_32/D vdd OAI21X1
XAOI22X1_3 AOI22X1_3/A INVX1_49/A INVX8_2/Y MUX2X1_74/Y gnd AOI22X1_3/Y vdd AOI22X1
XNAND2X1_46 MUX2X1_67/B NAND3X1_5/Y gnd NAND2X1_46/Y vdd NAND2X1
XNAND2X1_79 MUX2X1_241/A NAND3X1_6/Y gnd NAND2X1_79/Y vdd NAND2X1
XNAND2X1_57 MUX2X1_114/B NAND2X1_56/B gnd NAND2X1_57/Y vdd NAND2X1
XAOI22X1_22 MUX2X1_185/Y AND2X2_3/A AND2X2_2/B AOI22X1_22/D gnd AOI22X1_22/Y vdd AOI22X1
XNAND2X1_35 MUX2X1_187/A OAI21X1_25/B gnd NAND2X1_35/Y vdd NAND2X1
XAOI22X1_11 MUX2X1_119/Y INVX1_49/A INVX8_2/Y AOI22X1_11/D gnd AOI22X1_11/Y vdd AOI22X1
XNAND2X1_13 MUX2X1_148/A OAI21X1_9/B gnd NAND2X1_13/Y vdd NAND2X1
XNAND2X1_68 MUX2X1_160/A NAND2X1_64/B gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_24 MUX2X1_171/B NAND3X1_3/Y gnd OAI21X1_21/C vdd NAND2X1
XFILL_23_1_0 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_139 MUX2X1_234/B CLKBUF1_12/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 NOR2X1_16/A CLKBUF1_4/A AOI21X1_13/Y gnd vdd DFFPOSX1
XMUX2X1_204 NOR2X1_28/A INVX1_7/A BUFX4_29/Y gnd MUX2X1_204/Y vdd MUX2X1
XDFFPOSX1_117 MUX2X1_91/B CLKBUF1_36/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 NAND2X1_36/A CLKBUF1_15/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XMUX2X1_237 INVX1_48/A INVX1_40/A BUFX4_29/Y gnd MUX2X1_239/B vdd MUX2X1
XMUX2X1_226 MUX2X1_226/A MUX2X1_226/B BUFX4_33/Y gnd MUX2X1_226/Y vdd MUX2X1
XMUX2X1_248 MUX2X1_247/Y MUX2X1_248/B BUFX4_11/Y gnd MUX2X1_248/Y vdd MUX2X1
XINVX8_2 OR2X2_2/Y gnd INVX8_2/Y vdd INVX8
XMUX2X1_215 MUX2X1_215/A MUX2X1_213/Y BUFX4_16/Y gnd AOI22X1_27/A vdd MUX2X1
XFILL_3_0_0 gnd vdd FILL
XBUFX4_55 INVX8_3/Y gnd BUFX4_55/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_44 INVX8_10/Y gnd BUFX4_44/Y vdd BUFX4
XBUFX4_11 BUFX4_12/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_33 BUFX4_34/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_22 INVX8_9/Y gnd BUFX4_22/Y vdd BUFX4
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_1_3_1 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_161 BUFX4_55/Y NAND3X1_12/Y OAI21X1_161/C gnd OAI21X1_161/Y vdd OAI21X1
XAOI22X1_4 AOI22X1_4/A AND2X2_4/B AND2X2_1/B AOI22X1_4/D gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_150 OAI21X1_148/A BUFX4_23/Y OAI21X1_150/C gnd DFFPOSX1_15/D vdd OAI21X1
XAOI22X1_23 AOI22X1_23/A INVX1_49/A INVX8_2/Y MUX2X1_194/Y gnd AOI22X1_23/Y vdd AOI22X1
XNAND2X1_25 NAND2X1_25/A NAND3X1_3/Y gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_69 MUX2X1_184/A NAND2X1_64/B gnd NAND2X1_69/Y vdd NAND2X1
XAOI22X1_12 AOI22X1_12/A AND2X2_4/B AND2X2_1/B MUX2X1_128/Y gnd AOI22X1_12/Y vdd AOI22X1
XNAND2X1_58 NAND2X1_58/A NAND2X1_56/B gnd OAI21X1_52/C vdd NAND2X1
XNAND2X1_47 MUX2X1_91/B NAND3X1_5/Y gnd OAI21X1_42/C vdd NAND2X1
XNAND2X1_14 NAND2X1_14/A OAI21X1_9/B gnd NAND2X1_14/Y vdd NAND2X1
XNAND2X1_36 NAND2X1_36/A OAI21X1_25/B gnd NAND2X1_36/Y vdd NAND2X1
XFILL_23_1_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XDFFPOSX1_129 NOR2X1_17/A CLKBUF1_49/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 MUX2X1_235/A CLKBUF1_11/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_118 MUX2X1_115/B CLKBUF1_32/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XCLKBUF1_1 CLKBUF1_1/A gnd CLKBUF1_1/Y vdd CLKBUF1
XINVX8_3 datain[0] gnd INVX8_3/Y vdd INVX8
XMUX2X1_238 INVX1_57/A NOR2X1_39/A BUFX4_30/Y gnd MUX2X1_239/A vdd MUX2X1
XMUX2X1_227 MUX2X1_226/Y MUX2X1_227/B BUFX4_12/Y gnd AOI22X1_29/A vdd MUX2X1
XMUX2X1_249 INVX1_58/Y MUX2X1_9/B MUX2X1_249/S gnd DFFPOSX1_1/D vdd MUX2X1
XMUX2X1_216 NOR2X1_56/A MUX2X1_216/B INVX2_3/A gnd MUX2X1_216/Y vdd MUX2X1
XFILL_3_0_1 gnd vdd FILL
XMUX2X1_205 INVX1_23/A MUX2X1_205/B BUFX4_30/Y gnd MUX2X1_205/Y vdd MUX2X1
XBUFX4_56 INVX8_3/Y gnd BUFX4_56/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_12 BUFX4_12/A gnd BUFX4_12/Y vdd BUFX4
XBUFX4_34 BUFX4_34/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_23 INVX8_9/Y gnd BUFX4_23/Y vdd BUFX4
XBUFX4_45 INVX8_7/Y gnd BUFX4_45/Y vdd BUFX4
XOAI21X1_151 INVX2_5/A INVX8_11/A MUX2X1_225/A gnd OAI21X1_151/Y vdd OAI21X1
XNAND2X1_15 MUX2X1_196/A OAI21X1_9/B gnd NAND2X1_15/Y vdd NAND2X1
XAOI22X1_24 AOI22X1_24/A AND2X2_4/B AND2X2_1/B AOI22X1_24/D gnd AOI22X1_24/Y vdd AOI22X1
XNAND2X1_37 MUX2X1_235/A OAI21X1_25/B gnd NAND2X1_37/Y vdd NAND2X1
XNAND2X1_48 MUX2X1_115/B NAND3X1_5/Y gnd NAND2X1_48/Y vdd NAND2X1
XAOI22X1_13 MUX2X1_131/Y INVX8_11/Y INVX8_1/Y MUX2X1_134/Y gnd AOI22X1_13/Y vdd AOI22X1
XNAND2X1_59 NAND2X1_59/A NAND2X1_56/B gnd OAI21X1_53/C vdd NAND2X1
XOAI21X1_140 OAI21X1_148/A BUFX4_50/Y OAI21X1_140/C gnd DFFPOSX1_10/D vdd OAI21X1
XAOI22X1_5 AOI22X1_5/A INVX8_11/Y INVX8_1/Y MUX2X1_86/Y gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_26 MUX2X1_219/B NAND3X1_3/Y gnd NAND2X1_26/Y vdd NAND2X1
XOAI21X1_162 BUFX4_51/Y NAND3X1_12/Y NAND2X1_168/Y gnd DFFPOSX1_34/D vdd OAI21X1
XFILL_19_1 gnd vdd FILL
XMUX2X1_1 INVX1_1/Y BUFX4_57/Y MUX2X1_6/S gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_108 MUX2X1_58/A CLKBUF1_6/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_119 MUX2X1_139/B CLKBUF1_25/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XCLKBUF1_2 CLKBUF1_2/A gnd CLKBUF1_2/Y vdd CLKBUF1
XMUX2X1_239 MUX2X1_239/A MUX2X1_239/B BUFX4_16/Y gnd AOI22X1_31/A vdd MUX2X1
XMUX2X1_228 NOR2X1_29/A INVX1_8/A BUFX4_34/Y gnd MUX2X1_228/Y vdd MUX2X1
XMUX2X1_217 MUX2X1_217/A MUX2X1_217/B BUFX4_38/Y gnd MUX2X1_218/A vdd MUX2X1
XMUX2X1_206 MUX2X1_205/Y MUX2X1_204/Y INVX2_6/A gnd MUX2X1_206/Y vdd MUX2X1
XBUFX4_57 INVX8_3/Y gnd BUFX4_57/Y vdd BUFX4
XBUFX4_13 BUFX4_12/A gnd INVX2_6/A vdd BUFX4
XBUFX4_24 INVX8_6/Y gnd BUFX4_24/Y vdd BUFX4
XBUFX4_35 BUFX4_34/A gnd BUFX4_35/Y vdd BUFX4
XINVX8_4 datain[1] gnd INVX8_4/Y vdd INVX8
XBUFX4_46 INVX8_7/Y gnd BUFX4_46/Y vdd BUFX4
XDFFPOSX1_90 INVX1_10/A CLKBUF1_14/Y MUX2X1_10/Y gnd vdd DFFPOSX1
XFILL_21_2_0 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XNAND3X1_1 INVX2_2/A INVX2_7/Y AND2X2_1/B gnd NAND2X1_1/B vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XNAND2X1_27 MUX2X1_243/B NAND3X1_3/Y gnd NAND2X1_27/Y vdd NAND2X1
XOAI21X1_152 OAI21X1_148/A BUFX4_43/Y OAI21X1_151/Y gnd OAI21X1_152/Y vdd OAI21X1
XNAND2X1_38 MUX2X1_58/A NAND3X1_4/Y gnd OAI21X1_33/C vdd NAND2X1
XOAI21X1_141 INVX2_5/A INVX8_11/A MUX2X1_105/A gnd OAI21X1_141/Y vdd OAI21X1
XFILL_17_1_0 gnd vdd FILL
XNAND2X1_49 MUX2X1_139/B NAND3X1_5/Y gnd NAND2X1_49/Y vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XOAI21X1_163 BUFX4_8/Y NAND3X1_12/Y NAND2X1_169/Y gnd DFFPOSX1_35/D vdd OAI21X1
XOAI21X1_130 NAND2X1_132/Y NAND2X1_133/Y INVX4_1/Y gnd AOI21X1_39/B vdd OAI21X1
XAOI22X1_6 MUX2X1_89/Y AND2X2_3/A AND2X2_2/B MUX2X1_92/Y gnd AOI22X1_6/Y vdd AOI22X1
XNAND2X1_16 MUX2X1_220/A OAI21X1_9/B gnd OAI21X1_15/C vdd NAND2X1
XAOI22X1_14 MUX2X1_137/Y AND2X2_3/A AND2X2_2/B AOI22X1_14/D gnd AOI22X1_14/Y vdd AOI22X1
XAOI22X1_25 AOI22X1_25/A INVX8_11/Y INVX8_1/Y MUX2X1_206/Y gnd AOI22X1_25/Y vdd AOI22X1
XFILL_19_2 gnd vdd FILL
XCLKBUF1_3 CLKBUF1_3/A gnd CLKBUF1_3/Y vdd CLKBUF1
XDFFPOSX1_109 MUX2X1_82/A CLKBUF1_4/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XMUX2X1_2 INVX1_2/Y MUX2X1_2/B MUX2X1_6/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_6_0_0 gnd vdd FILL
XMUX2X1_229 INVX1_24/A MUX2X1_229/B BUFX4_35/Y gnd MUX2X1_229/Y vdd MUX2X1
XMUX2X1_218 MUX2X1_218/A MUX2X1_216/Y BUFX4_17/Y gnd AOI22X1_27/D vdd MUX2X1
XMUX2X1_207 INVX1_65/A INVX1_15/A BUFX4_31/Y gnd MUX2X1_207/Y vdd MUX2X1
XDFFPOSX1_80 MUX2X1_243/B CLKBUF1_3/A OAI21X1_24/Y gnd vdd DFFPOSX1
XBUFX4_58 INVX8_3/Y gnd BUFX4_58/Y vdd BUFX4
XDFFPOSX1_91 INVX1_11/A CLKBUF1_10/Y MUX2X1_11/Y gnd vdd DFFPOSX1
XINVX8_5 datain[2] gnd INVX8_5/Y vdd INVX8
XBUFX4_14 BUFX4_12/A gnd BUFX4_14/Y vdd BUFX4
XBUFX4_36 BUFX4_34/A gnd BUFX4_36/Y vdd BUFX4
XBUFX4_25 INVX8_6/Y gnd BUFX4_25/Y vdd BUFX4
XBUFX4_47 INVX8_7/Y gnd BUFX4_47/Y vdd BUFX4
XFILL_21_2_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XNAND3X1_2 INVX2_2/A INVX2_1/Y AND2X2_4/B gnd OAI21X1_9/B vdd NAND3X1
XNAND2X1_17 NAND2X1_17/A OAI21X1_9/B gnd NAND2X1_17/Y vdd NAND2X1
XOAI21X1_153 BUFX4_55/Y NAND3X1_11/Y OAI21X1_153/C gnd DFFPOSX1_25/D vdd OAI21X1
XOAI21X1_120 BUFX4_41/Y OAI21X1_118/B OAI21X1_120/C gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_142 OAI21X1_148/A BUFX4_7/Y OAI21X1_141/Y gnd OAI21X1_142/Y vdd OAI21X1
XOAI21X1_164 BUFX4_28/Y NAND3X1_12/Y NAND2X1_170/Y gnd DFFPOSX1_36/D vdd OAI21X1
XOAI21X1_131 OAI21X1_131/A NAND2X1_136/Y INVX4_1/Y gnd AOI21X1_40/B vdd OAI21X1
XNAND2X1_28 INVX2_7/Y AND2X2_3/Y gnd MUX2X1_9/S vdd NAND2X1
XNAND2X1_170 MUX2X1_151/B NAND3X1_12/Y gnd NAND2X1_170/Y vdd NAND2X1
XFILL_9_2_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_39 MUX2X1_82/A NAND3X1_4/Y gnd NAND2X1_39/Y vdd NAND2X1
XAOI22X1_7 MUX2X1_95/Y INVX1_49/A INVX8_2/Y AOI22X1_7/D gnd AOI22X1_7/Y vdd AOI22X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 AOI22X1_15/A INVX1_49/A INVX8_2/Y MUX2X1_146/Y gnd AOI22X1_15/Y vdd AOI22X1
XAOI22X1_26 MUX2X1_209/Y AND2X2_3/A AND2X2_2/B AOI22X1_26/D gnd AOI22X1_26/Y vdd AOI22X1
XFILL_19_3 gnd vdd FILL
XMUX2X1_3 INVX1_3/Y BUFX4_6/Y MUX2X1_6/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 CLKBUF1_4/A gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XFILL_24_1 gnd vdd FILL
XMUX2X1_219 NOR2X1_67/A MUX2X1_219/B BUFX4_39/Y gnd MUX2X1_221/B vdd MUX2X1
XMUX2X1_208 NAND2X1_70/A INVX1_31/A BUFX4_32/Y gnd MUX2X1_208/Y vdd MUX2X1
XDFFPOSX1_81 NOR2X1_2/A CLKBUF1_50/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_70 INVX1_6/A CLKBUF1_31/Y MUX2X1_6/Y gnd vdd DFFPOSX1
XBUFX4_59 INVX8_3/Y gnd MUX2X1_9/B vdd BUFX4
XBUFX4_15 BUFX4_12/A gnd BUFX4_15/Y vdd BUFX4
XBUFX4_26 INVX8_6/Y gnd BUFX4_26/Y vdd BUFX4
XINVX8_6 datain[3] gnd INVX8_6/Y vdd INVX8
XBUFX4_37 BUFX4_34/A gnd INVX2_3/A vdd BUFX4
XDFFPOSX1_92 INVX1_12/A CLKBUF1_8/Y MUX2X1_12/Y gnd vdd DFFPOSX1
XBUFX4_48 INVX8_7/Y gnd BUFX4_48/Y vdd BUFX4
XDFFPOSX1_260 MUX2X1_217/B CLKBUF1_39/Y OAI21X1_127/Y gnd vdd DFFPOSX1
XOAI21X1_110 BUFX4_3/Y NAND3X1_8/Y NAND2X1_108/Y gnd OAI21X1_110/Y vdd OAI21X1
XOAI21X1_121 BUFX4_56/Y NAND3X1_9/Y NAND2X1_120/Y gnd OAI21X1_121/Y vdd OAI21X1
XOAI21X1_132 NAND2X1_138/Y NAND2X1_139/Y INVX4_1/Y gnd AOI21X1_41/B vdd OAI21X1
XNAND3X1_3 INVX2_2/A INVX2_7/Y AND2X2_4/B gnd NAND3X1_3/Y vdd NAND3X1
XOAI21X1_143 INVX2_5/A INVX8_11/A MUX2X1_129/A gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_165 BUFX4_47/Y NAND3X1_12/Y OAI21X1_165/C gnd OAI21X1_165/Y vdd OAI21X1
XOAI21X1_154 BUFX4_52/Y NAND3X1_11/Y OAI21X1_154/C gnd DFFPOSX1_26/D vdd OAI21X1
XAOI22X1_8 AOI22X1_8/A AND2X2_4/B AND2X2_1/B AOI22X1_8/D gnd AOI22X1_8/Y vdd AOI22X1
XNAND2X1_29 AND2X2_2/B NOR2X1_11/Y gnd OAI21X1_25/B vdd NAND2X1
XAOI22X1_16 AOI22X1_16/A AND2X2_4/B AND2X2_1/B MUX2X1_152/Y gnd AOI22X1_16/Y vdd AOI22X1
XNAND2X1_18 INVX2_4/A NOR2X1_48/Y gnd INVX8_1/A vdd NAND2X1
XAOI22X1_27 AOI22X1_27/A INVX1_49/A INVX8_2/Y AOI22X1_27/D gnd AOI22X1_27/Y vdd AOI22X1
XNAND2X1_171 MUX2X1_175/B NAND3X1_12/Y gnd OAI21X1_165/C vdd NAND2X1
XNAND2X1_160 MUX2X1_100/B NAND3X1_11/Y gnd OAI21X1_154/C vdd NAND2X1
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_60 BUFX4_23/Y AND2X2_4/Y NOR2X1_67/Y gnd AOI21X1_60/Y vdd AOI21X1
XMUX2X1_4 INVX1_4/Y BUFX4_27/Y MUX2X1_6/S gnd MUX2X1_4/Y vdd MUX2X1
XFILL_24_2 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XCLKBUF1_5 CLKBUF1_5/A gnd CLKBUF1_5/Y vdd CLKBUF1
XMUX2X1_209 MUX2X1_208/Y MUX2X1_207/Y BUFX4_14/Y gnd MUX2X1_209/Y vdd MUX2X1
XDFFPOSX1_60 MUX2X1_148/A CLKBUF1_6/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XINVX8_7 datain[4] gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_82 NOR2X1_3/A CLKBUF1_47/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 INVX1_7/A CLKBUF1_26/Y MUX2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 INVX1_13/A CLKBUF1_2/Y MUX2X1_13/Y gnd vdd DFFPOSX1
XFILL_15_2_0 gnd vdd FILL
XBUFX4_16 BUFX4_12/A gnd BUFX4_16/Y vdd BUFX4
XBUFX4_38 BUFX4_34/A gnd BUFX4_38/Y vdd BUFX4
XBUFX4_27 INVX8_6/Y gnd BUFX4_27/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XBUFX4_49 INVX8_7/Y gnd MUX2X1_5/B vdd BUFX4
XBUFX4_1 INVX8_8/Y gnd BUFX4_1/Y vdd BUFX4
XFILL_21_0_0 gnd vdd FILL
XDFFPOSX1_261 MUX2X1_241/B CLKBUF1_33/Y OAI21X1_128/Y gnd vdd DFFPOSX1
XINVX4_1 rw gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XDFFPOSX1_250 MUX2X1_154/B CLKBUF1_16/Y OAI21X1_117/Y gnd vdd DFFPOSX1
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_155 BUFX4_10/Y NAND3X1_11/Y NAND2X1_161/Y gnd OAI21X1_155/Y vdd OAI21X1
XOAI21X1_166 BUFX4_3/Y NAND3X1_12/Y NAND2X1_172/Y gnd DFFPOSX1_38/D vdd OAI21X1
XNAND3X1_4 INVX2_1/Y INVX2_2/A INVX8_11/Y gnd NAND3X1_4/Y vdd NAND3X1
XAOI22X1_9 AOI22X1_9/A INVX8_11/Y INVX8_1/Y AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_100 BUFX4_28/Y NAND3X1_7/Y NAND2X1_95/Y gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_111 BUFX4_19/Y NAND3X1_8/Y OAI21X1_111/C gnd OAI21X1_111/Y vdd OAI21X1
XOAI21X1_144 OAI21X1_148/A BUFX4_25/Y OAI21X1_143/Y gnd DFFPOSX1_12/D vdd OAI21X1
XOAI21X1_133 NAND2X1_141/Y NAND2X1_142/Y INVX4_1/Y gnd AOI21X1_42/B vdd OAI21X1
XOAI21X1_122 BUFX4_52/Y NAND3X1_9/Y NAND2X1_121/Y gnd OAI21X1_122/Y vdd OAI21X1
XNAND2X1_161 MUX2X1_124/B NAND3X1_11/Y gnd NAND2X1_161/Y vdd NAND2X1
XNAND2X1_172 MUX2X1_199/B NAND3X1_12/Y gnd NAND2X1_172/Y vdd NAND2X1
XNAND2X1_150 AOI22X1_29/Y AOI22X1_30/Y gnd NAND2X1_150/Y vdd NAND2X1
XNAND2X1_19 INVX8_1/Y NOR2X1_1/Y gnd MUX2X1_6/S vdd NAND2X1
XAOI22X1_17 AOI22X1_17/A INVX8_11/Y INVX8_1/Y MUX2X1_158/Y gnd AOI22X1_17/Y vdd AOI22X1
XAOI22X1_28 AOI22X1_28/A AND2X2_4/B AND2X2_1/B MUX2X1_224/Y gnd AOI22X1_28/Y vdd AOI22X1
XAOI21X1_61 BUFX4_40/Y AND2X2_4/Y NOR2X1_68/Y gnd AOI21X1_61/Y vdd AOI21X1
XOAI21X1_1 BUFX4_55/Y NAND2X1_1/B OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_10_3_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XAOI21X1_50 BUFX4_48/Y NOR2X1_50/B NOR2X1_54/Y gnd AOI21X1_50/Y vdd AOI21X1
XMUX2X1_5 INVX1_5/Y MUX2X1_5/B MUX2X1_6/S gnd MUX2X1_5/Y vdd MUX2X1
XFILL_24_3 gnd vdd FILL
XCLKBUF1_6 CLKBUF1_5/A gnd CLKBUF1_6/Y vdd CLKBUF1
XINVX8_8 datain[5] gnd INVX8_8/Y vdd INVX8
XDFFPOSX1_94 INVX1_14/A CLKBUF1_67/Y MUX2X1_14/Y gnd vdd DFFPOSX1
XFILL_15_2_1 gnd vdd FILL
XDFFPOSX1_72 INVX1_8/A CLKBUF1_22/Y MUX2X1_8/Y gnd vdd DFFPOSX1
XBUFX4_17 BUFX4_12/A gnd BUFX4_17/Y vdd BUFX4
XDFFPOSX1_83 NOR2X1_4/A CLKBUF1_41/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XBUFX4_28 INVX8_6/Y gnd BUFX4_28/Y vdd BUFX4
XBUFX4_39 BUFX4_34/A gnd BUFX4_39/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XDFFPOSX1_50 NAND2X1_2/A CLKBUF1_47/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 NAND2X1_14/A CLKBUF1_1/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_251 MUX2X1_178/B CLKBUF1_10/Y OAI21X1_118/Y gnd vdd DFFPOSX1
XFILL_21_0_1 gnd vdd FILL
XBUFX4_2 INVX8_8/Y gnd BUFX4_2/Y vdd BUFX4
XDFFPOSX1_262 BUFX2_1/A CLKBUF1_32/Y AOI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_240 MUX2X1_120/B CLKBUF1_41/A OAI21X1_107/Y gnd vdd DFFPOSX1
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XOAI21X1_112 BUFX4_42/Y NAND3X1_8/Y NAND2X1_110/Y gnd OAI21X1_112/Y vdd OAI21X1
XNAND3X1_5 INVX2_2/A NAND3X1_5/B AND2X2_2/B gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_101 MUX2X1_5/B NAND3X1_7/Y NAND2X1_96/Y gnd OAI21X1_101/Y vdd OAI21X1
XNAND2X1_151 AOI22X1_31/Y AOI22X1_32/Y gnd OAI21X1_136/B vdd NAND2X1
XOAI21X1_134 NAND2X1_144/Y NAND2X1_145/Y INVX4_1/Y gnd AOI21X1_43/B vdd OAI21X1
XAOI22X1_29 AOI22X1_29/A INVX8_11/Y INVX8_1/Y MUX2X1_230/Y gnd AOI22X1_29/Y vdd AOI22X1
XOAI21X1_123 BUFX4_9/Y NAND3X1_9/Y NAND2X1_122/Y gnd OAI21X1_123/Y vdd OAI21X1
XNAND2X1_162 MUX2X1_148/B NAND3X1_11/Y gnd OAI21X1_156/C vdd NAND2X1
XOAI21X1_156 BUFX4_24/Y NAND3X1_11/Y OAI21X1_156/C gnd OAI21X1_156/Y vdd OAI21X1
XNAND2X1_140 rw BUFX2_5/A gnd AOI21X1_42/A vdd NAND2X1
XOAI21X1_145 INVX2_5/A INVX8_11/A MUX2X1_153/A gnd OAI21X1_145/Y vdd OAI21X1
XAOI22X1_18 MUX2X1_161/Y AND2X2_3/A AND2X2_2/B AOI22X1_18/D gnd AOI22X1_18/Y vdd AOI22X1
XOAI21X1_167 BUFX4_21/Y NAND3X1_12/Y NAND2X1_173/Y gnd OAI21X1_167/Y vdd OAI21X1
XNAND2X1_173 MUX2X1_223/B NAND3X1_12/Y gnd NAND2X1_173/Y vdd NAND2X1
XMUX2X1_190 INVX1_55/A NOR2X1_37/A BUFX4_31/Y gnd MUX2X1_191/A vdd MUX2X1
XAOI21X1_51 BUFX4_1/Y NOR2X1_50/B NOR2X1_55/Y gnd AOI21X1_51/Y vdd AOI21X1
XAOI21X1_40 AOI21X1_40/A AOI21X1_40/B NOR2X1_46/B gnd AOI21X1_40/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 BUFX4_51/Y NAND2X1_1/B OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XCLKBUF1_7 CLKBUF1_7/A gnd CLKBUF1_7/Y vdd CLKBUF1
XMUX2X1_6 INVX1_6/Y BUFX4_5/Y MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XDFFPOSX1_73 MUX2X1_75/B CLKBUF1_17/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_62 MUX2X1_196/A CLKBUF1_67/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XBUFX4_18 BUFX4_12/A gnd BUFX4_18/Y vdd BUFX4
XDFFPOSX1_51 NAND2X1_3/A CLKBUF1_41/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 MUX2X1_247/B CLKBUF1_23/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_84 NOR2X1_5/A CLKBUF1_39/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XBUFX4_29 BUFX4_34/A gnd BUFX4_29/Y vdd BUFX4
XINVX8_9 datain[6] gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_95 INVX1_15/A CLKBUF1_27/A MUX2X1_15/Y gnd vdd DFFPOSX1
XFILL_22_1 gnd vdd FILL
XBUFX4_3 INVX8_8/Y gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_230 INVX1_50/A CLKBUF1_30/Y MUX2X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_241 MUX2X1_144/B CLKBUF1_51/Y OAI21X1_108/Y gnd vdd DFFPOSX1
XDFFPOSX1_263 BUFX2_2/A CLKBUF1_26/Y AOI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_252 MUX2X1_202/B CLKBUF1_5/Y OAI21X1_119/Y gnd vdd DFFPOSX1
XNAND3X1_6 INVX2_2/A INVX2_1/Y INVX8_2/Y gnd NAND3X1_6/Y vdd NAND3X1
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 BUFX4_3/Y NAND3X1_7/Y NAND2X1_97/Y gnd OAI21X1_102/Y vdd OAI21X1
XOAI21X1_113 BUFX4_58/Y OAI21X1_118/B NAND2X1_112/Y gnd OAI21X1_113/Y vdd OAI21X1
XNAND2X1_130 AOI22X1_3/Y AOI22X1_4/Y gnd OAI21X1_129/B vdd NAND2X1
XFILL_13_3_0 gnd vdd FILL
XOAI21X1_124 BUFX4_26/Y NAND3X1_9/Y OAI21X1_124/C gnd OAI21X1_124/Y vdd OAI21X1
XNAND2X1_174 MUX2X1_247/B NAND3X1_12/Y gnd OAI21X1_168/C vdd NAND2X1
XOAI21X1_168 BUFX4_44/Y NAND3X1_12/Y OAI21X1_168/C gnd DFFPOSX1_40/D vdd OAI21X1
XNAND2X1_152 INVX1_67/A INVX1_59/Y gnd NOR2X1_47/B vdd NAND2X1
XOAI21X1_146 OAI21X1_148/A BUFX4_45/Y OAI21X1_145/Y gnd OAI21X1_146/Y vdd OAI21X1
XOAI21X1_135 NAND2X1_147/Y NAND2X1_148/Y INVX4_1/Y gnd AOI21X1_44/B vdd OAI21X1
XNAND2X1_141 AOI22X1_17/Y AOI22X1_18/Y gnd NAND2X1_141/Y vdd NAND2X1
XNAND2X1_163 MUX2X1_172/B NAND3X1_11/Y gnd NAND2X1_163/Y vdd NAND2X1
XOAI21X1_157 BUFX4_46/Y NAND3X1_11/Y NAND2X1_163/Y gnd DFFPOSX1_29/D vdd OAI21X1
XMUX2X1_180 NOR2X1_27/A INVX1_6/A BUFX4_35/Y gnd MUX2X1_180/Y vdd MUX2X1
XMUX2X1_191 MUX2X1_191/A MUX2X1_191/B BUFX4_16/Y gnd AOI22X1_23/A vdd MUX2X1
XAOI22X1_19 MUX2X1_167/Y INVX1_49/A INVX8_2/Y MUX2X1_170/Y gnd AOI22X1_19/Y vdd AOI22X1
XAOI21X1_30 BUFX4_1/Y NOR2X1_39/B NOR2X1_37/Y gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_41 AOI21X1_41/A AOI21X1_41/B NOR2X1_46/B gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_52 BUFX4_19/Y NOR2X1_50/B NOR2X1_56/Y gnd AOI21X1_52/Y vdd AOI21X1
XOAI21X1_3 BUFX4_9/Y NAND2X1_1/B OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XFILL_10_1_0 gnd vdd FILL
XCLKBUF1_8 CLKBUF1_8/A gnd CLKBUF1_8/Y vdd CLKBUF1
XMUX2X1_7 INVX1_7/Y MUX2X1_7/B MUX2X1_6/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_2_2_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XDFFPOSX1_41 MUX2X1_75/A CLKBUF1_17/Y AOI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 MUX2X1_196/B CLKBUF1_67/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_96 INVX1_16/A CLKBUF1_67/Y MUX2X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 NAND2X1_4/A CLKBUF1_37/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XBUFX4_19 INVX8_9/Y gnd BUFX4_19/Y vdd BUFX4
XDFFPOSX1_85 NOR2X1_6/A CLKBUF1_35/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 MUX2X1_99/B CLKBUF1_13/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 MUX2X1_220/A CLKBUF1_2/A OAI21X1_15/Y gnd vdd DFFPOSX1
XFILL_15_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XBUFX4_4 INVX8_8/Y gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_253 MUX2X1_226/B CLKBUF1_3/Y OAI21X1_120/Y gnd vdd DFFPOSX1
XDFFPOSX1_264 BUFX2_3/A CLKBUF1_21/Y AOI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_220 INVX1_47/A CLKBUF1_8/Y MUX2X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_231 INVX1_51/A CLKBUF1_28/Y MUX2X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_242 MUX2X1_168/B CLKBUF1_45/Y OAI21X1_109/Y gnd vdd DFFPOSX1
XNAND3X1_7 INVX2_2/A INVX2_1/Y AND2X2_1/B gnd NAND3X1_7/Y vdd NAND3X1
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_147 INVX2_5/A INVX8_11/A MUX2X1_177/A gnd OAI21X1_147/Y vdd OAI21X1
XOAI21X1_158 BUFX4_2/Y NAND3X1_11/Y NAND2X1_164/Y gnd DFFPOSX1_30/D vdd OAI21X1
XNAND2X1_164 MUX2X1_196/B NAND3X1_11/Y gnd NAND2X1_164/Y vdd NAND2X1
XBUFX2_1 BUFX2_1/A gnd dataout[0] vdd BUFX2
XOAI21X1_136 NAND2X1_150/Y OAI21X1_136/B INVX4_1/Y gnd AOI21X1_45/B vdd OAI21X1
XNAND2X1_120 MUX2X1_73/B NAND3X1_9/Y gnd NAND2X1_120/Y vdd NAND2X1
XNAND2X1_175 INVX2_3/Y INVX2_6/Y gnd INVX2_7/A vdd NAND2X1
XNAND2X1_153 NOR2X1_45/Y AND2X2_3/Y gnd MUX2X1_249/S vdd NAND2X1
XNAND2X1_131 rw BUFX2_2/A gnd AOI21X1_39/A vdd NAND2X1
XNAND2X1_142 AOI22X1_19/Y AOI22X1_20/Y gnd NAND2X1_142/Y vdd NAND2X1
XOAI21X1_103 BUFX4_22/Y NAND3X1_7/Y NAND2X1_98/Y gnd OAI21X1_103/Y vdd OAI21X1
XOAI21X1_114 BUFX4_50/Y OAI21X1_118/B NAND2X1_113/Y gnd OAI21X1_114/Y vdd OAI21X1
XOAI21X1_125 BUFX4_47/Y NAND3X1_9/Y OAI21X1_125/C gnd OAI21X1_125/Y vdd OAI21X1
XAOI21X1_1 BUFX4_55/Y NOR2X1_2/B NOR2X1_2/Y gnd AOI21X1_1/Y vdd AOI21X1
XMUX2X1_192 NOR2X1_55/A MUX2X1_192/B BUFX4_32/Y gnd MUX2X1_194/B vdd MUX2X1
XMUX2X1_181 INVX1_22/A MUX2X1_181/B BUFX4_36/Y gnd MUX2X1_182/A vdd MUX2X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XMUX2X1_170 MUX2X1_169/Y MUX2X1_168/Y BUFX4_17/Y gnd MUX2X1_170/Y vdd MUX2X1
XAOI21X1_53 BUFX4_42/Y NOR2X1_50/B NOR2X1_57/Y gnd AOI21X1_53/Y vdd AOI21X1
XOAI21X1_4 BUFX4_28/Y NAND2X1_1/B OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_31 BUFX4_19/Y NOR2X1_39/B NOR2X1_38/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_42 AOI21X1_42/A AOI21X1_42/B NOR2X1_46/B gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_20 BUFX4_27/Y NOR2X1_22/B NOR2X1_25/Y gnd AOI21X1_20/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XCLKBUF1_9 CLKBUF1_9/A gnd CLKBUF1_9/Y vdd CLKBUF1
XMUX2X1_8 INVX1_8/Y BUFX4_41/Y MUX2X1_6/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XFILL_18_2_1 gnd vdd FILL
XDFFPOSX1_64 NAND2X1_17/A CLKBUF1_67/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 MUX2X1_123/B CLKBUF1_12/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 NOR2X1_7/A CLKBUF1_29/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX2_4/A CLKBUF1_49/Y AOI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 NOR2X1_53/A CLKBUF1_39/Y AOI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 MUX2X1_220/B CLKBUF1_2/A OAI21X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_53 NAND2X1_5/A CLKBUF1_35/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 NOR2X1_62/A CLKBUF1_13/Y AOI21X1_55/Y gnd vdd DFFPOSX1
XFILL_15_2 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX4_5 INVX8_8/Y gnd BUFX4_5/Y vdd BUFX4
XDFFPOSX1_243 MUX2X1_192/B CLKBUF1_43/Y OAI21X1_110/Y gnd vdd DFFPOSX1
XDFFPOSX1_221 INVX1_48/A CLKBUF1_3/Y MUX2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_254 MUX2X1_73/B CLKBUF1_67/Y OAI21X1_121/Y gnd vdd DFFPOSX1
XDFFPOSX1_265 BUFX2_4/A CLKBUF1_18/Y AOI21X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_232 INVX1_52/A CLKBUF1_23/Y MUX2X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_210 INVX1_37/A CLKBUF1_48/Y MUX2X1_37/Y gnd vdd DFFPOSX1
XOAI21X1_148 OAI21X1_148/A BUFX4_5/Y OAI21X1_147/Y gnd OAI21X1_148/Y vdd OAI21X1
XOAI21X1_137 INVX2_5/A INVX8_11/A MUX2X1_57/A gnd OAI21X1_138/C vdd OAI21X1
XNAND2X1_110 MUX2X1_240/B NAND3X1_8/Y gnd NAND2X1_110/Y vdd NAND2X1
XNAND2X1_143 rw BUFX2_6/A gnd AOI21X1_43/A vdd NAND2X1
XOAI21X1_126 BUFX4_1/Y NAND3X1_9/Y NAND2X1_125/Y gnd OAI21X1_126/Y vdd OAI21X1
XOAI21X1_115 BUFX4_6/Y OAI21X1_118/B OAI21X1_115/C gnd OAI21X1_115/Y vdd OAI21X1
XNAND3X1_8 INVX2_2/A INVX2_7/Y INVX8_2/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_104 BUFX4_44/Y NAND3X1_7/Y NAND2X1_99/Y gnd OAI21X1_104/Y vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd dataout[1] vdd BUFX2
XOAI21X1_159 BUFX4_22/Y NAND3X1_11/Y OAI21X1_159/C gnd OAI21X1_159/Y vdd OAI21X1
XNAND2X1_121 MUX2X1_97/B NAND3X1_9/Y gnd NAND2X1_121/Y vdd NAND2X1
XNAND2X1_132 AOI22X1_5/Y AOI22X1_6/Y gnd NAND2X1_132/Y vdd NAND2X1
XMUX2X1_182 MUX2X1_182/A MUX2X1_180/Y INVX2_6/A gnd AOI22X1_21/D vdd MUX2X1
XMUX2X1_193 MUX2X1_193/A MUX2X1_193/B BUFX4_33/Y gnd MUX2X1_193/Y vdd MUX2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XNAND2X1_154 INVX2_4/Y NOR2X1_48/Y gnd INVX8_11/A vdd NAND2X1
XNAND2X1_165 MUX2X1_220/B NAND3X1_11/Y gnd OAI21X1_159/C vdd NAND2X1
XAOI21X1_2 BUFX4_54/Y NOR2X1_2/B NOR2X1_3/Y gnd AOI21X1_2/Y vdd AOI21X1
XMUX2X1_160 MUX2X1_160/A INVX1_29/A BUFX4_33/Y gnd MUX2X1_160/Y vdd MUX2X1
XMUX2X1_171 NOR2X1_65/A MUX2X1_171/B BUFX4_29/Y gnd MUX2X1_173/B vdd MUX2X1
XAOI21X1_54 BUFX4_57/Y AND2X2_4/Y NOR2X1_61/Y gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_32 BUFX4_40/Y NOR2X1_39/B NOR2X1_39/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_43 AOI21X1_43/A AOI21X1_43/B NOR2X1_46/B gnd AOI21X1_43/Y vdd AOI21X1
XOAI21X1_5 BUFX4_47/Y NAND2X1_1/B OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_21 BUFX4_46/Y NOR2X1_22/B NOR2X1_26/Y gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_10 MUX2X1_2/B AND2X2_2/Y NOR2X1_13/Y gnd AOI21X1_10/Y vdd AOI21X1
XFILL_3_2 gnd vdd FILL
XMUX2X1_9 INVX1_9/Y MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XDFFPOSX1_32 MUX2X1_244/B CLKBUF1_67/Y DFFPOSX1_32/D gnd vdd DFFPOSX1
XDFFPOSX1_43 NOR2X1_63/A CLKBUF1_9/Y AOI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_65 INVX1_1/A CLKBUF1_52/Y MUX2X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 NAND2X1_6/A CLKBUF1_30/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_67/A CLKBUF1_46/Y AOI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 NAND2X1_23/A CLKBUF1_5/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 MUX2X1_81/A CLKBUF1_15/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XDFFPOSX1_87 NOR2X1_8/A CLKBUF1_27/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 NOR2X1_54/A CLKBUF1_35/Y AOI21X1_50/Y gnd vdd DFFPOSX1
XFILL_20_1 gnd vdd FILL
XDFFPOSX1_211 INVX1_38/A CLKBUF1_43/Y MUX2X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_233 INVX1_53/A CLKBUF1_20/Y MUX2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_222 NOR2X1_32/A CLKBUF1_65/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XBUFX4_6 INVX8_5/Y gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_266 BUFX2_5/A CLKBUF1_15/Y AOI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_244 MUX2X1_216/B CLKBUF1_39/Y OAI21X1_111/Y gnd vdd DFFPOSX1
XDFFPOSX1_200 NAND2X1_94/A CLKBUF1_24/Y OAI21X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_255 MUX2X1_97/B CLKBUF1_2/A OAI21X1_122/Y gnd vdd DFFPOSX1
XFILL_0_3_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XOAI21X1_138 OAI21X1_148/A BUFX4_57/Y OAI21X1_138/C gnd DFFPOSX1_9/D vdd OAI21X1
XOAI21X1_105 BUFX4_56/Y NAND3X1_8/Y OAI21X1_105/C gnd OAI21X1_105/Y vdd OAI21X1
XNAND3X1_9 INVX2_2/A NAND3X1_5/B INVX8_2/Y gnd NAND3X1_9/Y vdd NAND3X1
XBUFX2_3 BUFX2_3/A gnd dataout[2] vdd BUFX2
XOAI21X1_116 BUFX4_24/Y OAI21X1_118/B OAI21X1_116/C gnd OAI21X1_116/Y vdd OAI21X1
XOAI21X1_127 BUFX4_19/Y NAND3X1_9/Y NAND2X1_126/Y gnd OAI21X1_127/Y vdd OAI21X1
XOAI21X1_149 INVX2_5/A INVX8_11/A MUX2X1_201/A gnd OAI21X1_150/C vdd OAI21X1
XNAND2X1_166 MUX2X1_244/B NAND3X1_11/Y gnd OAI21X1_160/C vdd NAND2X1
XNAND2X1_144 AOI22X1_21/Y AOI22X1_22/Y gnd NAND2X1_144/Y vdd NAND2X1
XMUX2X1_183 INVX1_64/A INVX1_14/A INVX2_3/A gnd MUX2X1_183/Y vdd MUX2X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XNAND2X1_155 NOR2X1_45/Y INVX2_2/A gnd INVX2_5/A vdd NAND2X1
XNAND2X1_111 NAND3X1_5/B NOR2X1_20/Y gnd OAI21X1_118/B vdd NAND2X1
XNAND2X1_100 INVX1_49/A NOR2X1_1/Y gnd MUX2X1_39/S vdd NAND2X1
XAOI21X1_3 BUFX4_9/Y NOR2X1_2/B NOR2X1_4/Y gnd AOI21X1_3/Y vdd AOI21X1
XNAND2X1_122 MUX2X1_121/B NAND3X1_9/Y gnd NAND2X1_122/Y vdd NAND2X1
XMUX2X1_150 NOR2X1_5/A NAND2X1_4/A INVX2_3/A gnd MUX2X1_150/Y vdd MUX2X1
XNAND2X1_133 AOI22X1_7/Y AOI22X1_8/Y gnd NAND2X1_133/Y vdd NAND2X1
XMUX2X1_161 MUX2X1_160/Y MUX2X1_159/Y BUFX4_14/Y gnd MUX2X1_161/Y vdd MUX2X1
XMUX2X1_172 NAND2X1_14/A MUX2X1_172/B BUFX4_30/Y gnd MUX2X1_172/Y vdd MUX2X1
XMUX2X1_194 MUX2X1_193/Y MUX2X1_194/B BUFX4_17/Y gnd MUX2X1_194/Y vdd MUX2X1
XNOR2X1_1 INVX2_7/A INVX2_2/Y gnd NOR2X1_1/Y vdd NOR2X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_22 BUFX4_5/Y NOR2X1_22/B NOR2X1_27/Y gnd AOI21X1_22/Y vdd AOI21X1
XOAI21X1_6 BUFX4_3/Y NAND2X1_1/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_11 BUFX4_7/Y AND2X2_2/Y NOR2X1_14/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_33 ras INVX2_4/Y NOR2X1_40/Y gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_44 AOI21X1_44/A AOI21X1_44/B NOR2X1_46/B gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_55 MUX2X1_2/B AND2X2_4/Y NOR2X1_62/Y gnd AOI21X1_55/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XFILL_3_3 gnd vdd FILL
XDFFPOSX1_11 MUX2X1_105/A CLKBUF1_10/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 MUX2X1_79/B CLKBUF1_50/Y OAI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 NOR2X1_55/A CLKBUF1_29/Y AOI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 NOR2X1_9/A CLKBUF1_22/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX1_59/A CLKBUF1_42/Y AOI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 NOR2X1_64/A CLKBUF1_8/Y AOI21X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 NAND2X1_7/A CLKBUF1_27/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_77 MUX2X1_171/B CLKBUF1_1/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_2/A CLKBUF1_45/Y MUX2X1_2/Y gnd vdd DFFPOSX1
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_245 MUX2X1_240/B CLKBUF1_33/Y OAI21X1_112/Y gnd vdd DFFPOSX1
XBUFX4_7 INVX8_5/Y gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_201 NAND2X1_95/A CLKBUF1_19/Y OAI21X1_100/Y gnd vdd DFFPOSX1
XDFFPOSX1_256 MUX2X1_121/B CLKBUF1_41/A OAI21X1_123/Y gnd vdd DFFPOSX1
XDFFPOSX1_267 BUFX2_6/A CLKBUF1_10/Y AOI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_212 INVX1_39/A CLKBUF1_38/Y MUX2X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_223 NOR2X1_33/A CLKBUF1_25/A AOI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_234 INVX1_54/A CLKBUF1_14/Y MUX2X1_53/Y gnd vdd DFFPOSX1
XFILL_16_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XOAI21X1_128 BUFX4_42/Y NAND3X1_9/Y NAND2X1_127/Y gnd OAI21X1_128/Y vdd OAI21X1
XOAI21X1_106 BUFX4_51/Y NAND3X1_8/Y NAND2X1_104/Y gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_117 BUFX4_46/Y OAI21X1_118/B OAI21X1_117/C gnd OAI21X1_117/Y vdd OAI21X1
XNAND2X1_167 MUX2X1_79/B NAND3X1_12/Y gnd OAI21X1_161/C vdd NAND2X1
XNAND2X1_112 MUX2X1_58/B OAI21X1_118/B gnd NAND2X1_112/Y vdd NAND2X1
XNAND2X1_145 AOI22X1_23/Y AOI22X1_24/Y gnd NAND2X1_145/Y vdd NAND2X1
XNAND2X1_134 rw BUFX2_3/A gnd AOI21X1_40/A vdd NAND2X1
XBUFX2_4 BUFX2_4/A gnd dataout[3] vdd BUFX2
XNAND2X1_123 MUX2X1_145/B NAND3X1_9/Y gnd OAI21X1_124/C vdd NAND2X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XAOI21X1_4 BUFX4_28/Y NOR2X1_2/B NOR2X1_5/Y gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_139 INVX2_5/A INVX8_11/A MUX2X1_81/A gnd OAI21X1_140/C vdd OAI21X1
XNAND2X1_156 INVX8_11/Y INVX2_5/Y gnd OAI21X1_148/A vdd NAND2X1
XNAND2X1_101 INVX1_49/A INVX2_5/Y gnd MUX2X1_46/S vdd NAND2X1
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XMUX2X1_195 NOR2X1_66/A NAND2X1_25/A BUFX4_34/Y gnd MUX2X1_195/Y vdd MUX2X1
XMUX2X1_184 MUX2X1_184/A INVX1_30/A BUFX4_38/Y gnd MUX2X1_184/Y vdd MUX2X1
XMUX2X1_151 NAND2X1_95/A MUX2X1_151/B BUFX4_38/Y gnd MUX2X1_152/A vdd MUX2X1
XMUX2X1_140 MUX2X1_139/Y MUX2X1_140/B BUFX4_15/Y gnd AOI22X1_14/D vdd MUX2X1
XMUX2X1_162 NOR2X1_16/A NAND2X1_59/A BUFX4_34/Y gnd MUX2X1_164/B vdd MUX2X1
XMUX2X1_173 MUX2X1_172/Y MUX2X1_173/B BUFX4_18/Y gnd AOI22X1_20/A vdd MUX2X1
XAOI21X1_56 BUFX4_10/Y AND2X2_4/Y NOR2X1_63/Y gnd AOI21X1_56/Y vdd AOI21X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B NOR2X1_46/B gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_12 BUFX4_25/Y AND2X2_2/Y NOR2X1_15/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_34 ras INVX1_67/Y NOR2X1_41/Y gnd AOI21X1_34/Y vdd AOI21X1
XOAI21X1_7 BUFX4_22/Y NAND2X1_1/B OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_23 MUX2X1_7/B NOR2X1_22/B NOR2X1_28/Y gnd AOI21X1_23/Y vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_89 INVX1_9/A CLKBUF1_17/Y MUX2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 NAND2X1_25/A CLKBUF1_67/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 NAND2X1_8/A CLKBUF1_23/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_3/A CLKBUF1_42/Y MUX2X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 MUX2X1_129/A CLKBUF1_5/Y DFFPOSX1_12/D gnd vdd DFFPOSX1
XDFFPOSX1_23 NOR2X1_56/A CLKBUF1_28/Y AOI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 MUX2X1_103/B CLKBUF1_47/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_45 NOR2X1_65/A CLKBUF1_1/Y AOI21X1_58/Y gnd vdd DFFPOSX1
XFILL_18_0_1 gnd vdd FILL
XDFFPOSX1_213 INVX1_40/A CLKBUF1_33/Y MUX2X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_235 INVX1_55/A CLKBUF1_9/Y MUX2X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_246 MUX2X1_58/B CLKBUF1_31/Y OAI21X1_113/Y gnd vdd DFFPOSX1
XDFFPOSX1_257 MUX2X1_145/B CLKBUF1_51/Y OAI21X1_124/Y gnd vdd DFFPOSX1
XBUFX4_8 INVX8_5/Y gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_268 BUFX2_7/A CLKBUF1_6/Y AOI21X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_224 NOR2X1_34/A CLKBUF1_41/A AOI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_202 NAND2X1_96/A CLKBUF1_13/Y OAI21X1_101/Y gnd vdd DFFPOSX1
XOAI21X1_118 BUFX4_5/Y OAI21X1_118/B NAND2X1_117/Y gnd OAI21X1_118/Y vdd OAI21X1
XOAI21X1_129 OAI21X1_129/A OAI21X1_129/B INVX4_1/Y gnd AOI21X1_38/B vdd OAI21X1
XNAND2X1_102 INVX1_49/A NOR2X1_11/Y gnd MUX2X1_56/S vdd NAND2X1
XNAND2X1_135 AOI22X1_9/Y AOI22X1_10/Y gnd OAI21X1_131/A vdd NAND2X1
XOAI21X1_107 BUFX4_9/Y NAND3X1_8/Y OAI21X1_107/C gnd OAI21X1_107/Y vdd OAI21X1
XNAND2X1_157 INVX1_67/A INVX1_59/A gnd OR2X2_2/A vdd NAND2X1
XNAND2X1_146 rw BUFX2_7/A gnd AOI21X1_44/A vdd NAND2X1
XBUFX2_5 BUFX2_5/A gnd dataout[4] vdd BUFX2
XNAND2X1_168 MUX2X1_103/B NAND3X1_12/Y gnd NAND2X1_168/Y vdd NAND2X1
XNAND2X1_113 MUX2X1_82/B OAI21X1_118/B gnd NAND2X1_113/Y vdd NAND2X1
XNAND2X1_124 MUX2X1_169/B NAND3X1_9/Y gnd OAI21X1_125/C vdd NAND2X1
XMUX2X1_196 MUX2X1_196/A MUX2X1_196/B BUFX4_35/Y gnd MUX2X1_197/A vdd MUX2X1
XMUX2X1_185 MUX2X1_184/Y MUX2X1_183/Y BUFX4_14/Y gnd MUX2X1_185/Y vdd MUX2X1
XMUX2X1_141 INVX1_44/A INVX1_36/A BUFX4_31/Y gnd MUX2X1_143/B vdd MUX2X1
XMUX2X1_130 NAND2X1_41/A MUX2X1_130/B BUFX4_35/Y gnd MUX2X1_131/A vdd MUX2X1
XMUX2X1_152 MUX2X1_152/A MUX2X1_150/Y BUFX4_11/Y gnd MUX2X1_152/Y vdd MUX2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XAOI21X1_5 BUFX4_47/Y NOR2X1_2/B NOR2X1_6/Y gnd AOI21X1_5/Y vdd AOI21X1
XMUX2X1_174 NOR2X1_6/A NAND2X1_5/A BUFX4_31/Y gnd MUX2X1_174/Y vdd MUX2X1
XMUX2X1_163 MUX2X1_163/A MUX2X1_163/B BUFX4_35/Y gnd MUX2X1_164/A vdd MUX2X1
XAOI21X1_46 BUFX4_55/Y NOR2X1_50/B NOR2X1_50/Y gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_24 BUFX4_41/Y NOR2X1_22/B NOR2X1_29/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_35 ras INVX1_59/Y NOR2X1_42/Y gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_57 BUFX4_24/Y AND2X2_4/Y NOR2X1_64/Y gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_13 BUFX4_45/Y AND2X2_2/Y NOR2X1_16/Y gnd AOI21X1_13/Y vdd AOI21X1
XNOR2X1_3 NOR2X1_3/A NOR2X1_2/B gnd NOR2X1_3/Y vdd NOR2X1
XOAI21X1_8 BUFX4_44/Y NAND2X1_1/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XDFFPOSX1_57 MUX2X1_76/A CLKBUF1_20/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 NOR2X1_57/A CLKBUF1_22/Y AOI21X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_46 NOR2X1_66/A CLKBUF1_67/Y AOI21X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 MUX2X1_153/A CLKBUF1_4/Y OAI21X1_146/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 MUX2X1_127/B CLKBUF1_41/Y DFFPOSX1_35/D gnd vdd DFFPOSX1
XDFFPOSX1_68 INVX1_4/A CLKBUF1_38/Y MUX2X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_79 MUX2X1_219/B CLKBUF1_8/A OAI21X1_23/Y gnd vdd DFFPOSX1
XFILL_20_2_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XDFFPOSX1_225 NOR2X1_35/A CLKBUF1_50/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_203 MUX2X1_199/A CLKBUF1_9/Y OAI21X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_214 INVX1_41/A CLKBUF1_29/Y MUX2X1_41/Y gnd vdd DFFPOSX1
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_269 BUFX2_8/A CLKBUF1_3/Y AOI21X1_45/Y gnd vdd DFFPOSX1
XBUFX4_9 INVX8_5/Y gnd BUFX4_9/Y vdd BUFX4
XDFFPOSX1_236 INVX1_56/A CLKBUF1_8/Y MUX2X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_258 MUX2X1_169/B CLKBUF1_47/Y OAI21X1_125/Y gnd vdd DFFPOSX1
XDFFPOSX1_247 MUX2X1_82/B CLKBUF1_26/Y OAI21X1_114/Y gnd vdd DFFPOSX1
XNAND2X1_1 MUX2X1_78/B NAND2X1_1/B gnd OAI21X1_1/C vdd NAND2X1
XNAND2X1_103 MUX2X1_72/B NAND3X1_8/Y gnd OAI21X1_105/C vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd dataout[5] vdd BUFX2
XNAND2X1_125 MUX2X1_193/B NAND3X1_9/Y gnd NAND2X1_125/Y vdd NAND2X1
XOAI21X1_108 BUFX4_26/Y NAND3X1_8/Y OAI21X1_108/C gnd OAI21X1_108/Y vdd OAI21X1
XNAND2X1_114 MUX2X1_106/B OAI21X1_118/B gnd OAI21X1_115/C vdd NAND2X1
XNAND2X1_136 AOI22X1_11/Y AOI22X1_12/Y gnd NAND2X1_136/Y vdd NAND2X1
XNAND2X1_158 INVX1_59/A INVX1_67/Y gnd NOR2X1_60/B vdd NAND2X1
XNAND2X1_169 MUX2X1_127/B NAND3X1_12/Y gnd NAND2X1_169/Y vdd NAND2X1
XNAND2X1_147 AOI22X1_25/Y AOI22X1_26/Y gnd NAND2X1_147/Y vdd NAND2X1
XOAI21X1_119 BUFX4_21/Y OAI21X1_118/B OAI21X1_119/C gnd OAI21X1_119/Y vdd OAI21X1
XMUX2X1_142 INVX1_53/A NOR2X1_35/A BUFX4_32/Y gnd MUX2X1_143/A vdd MUX2X1
XAOI21X1_6 BUFX4_3/Y NOR2X1_2/B NOR2X1_7/Y gnd AOI21X1_6/Y vdd AOI21X1
XMUX2X1_186 NOR2X1_17/A MUX2X1_186/B BUFX4_39/Y gnd MUX2X1_188/B vdd MUX2X1
XDFFPOSX1_1 INVX1_58/A CLKBUF1_49/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XMUX2X1_197 MUX2X1_197/A MUX2X1_195/Y BUFX4_18/Y gnd AOI22X1_24/A vdd MUX2X1
XFILL_16_1_0 gnd vdd FILL
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XMUX2X1_120 NOR2X1_52/A MUX2X1_120/B BUFX4_39/Y gnd MUX2X1_120/Y vdd MUX2X1
XMUX2X1_131 MUX2X1_131/A MUX2X1_131/B BUFX4_12/Y gnd MUX2X1_131/Y vdd MUX2X1
XFILL_8_2_0 gnd vdd FILL
XMUX2X1_153 MUX2X1_153/A MUX2X1_153/B BUFX4_39/Y gnd MUX2X1_155/B vdd MUX2X1
XMUX2X1_164 MUX2X1_164/A MUX2X1_164/B BUFX4_15/Y gnd AOI22X1_18/D vdd MUX2X1
XFILL_0_1_0 gnd vdd FILL
XMUX2X1_175 NAND2X1_96/A MUX2X1_175/B BUFX4_32/Y gnd MUX2X1_175/Y vdd MUX2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XNOR2X1_4 NOR2X1_4/A NOR2X1_2/B gnd NOR2X1_4/Y vdd NOR2X1
XOAI21X1_9 BUFX4_55/Y OAI21X1_9/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_25 BUFX4_56/Y NOR2X1_39/B NOR2X1_32/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_14 BUFX4_4/Y AND2X2_2/Y NOR2X1_17/Y gnd AOI21X1_14/Y vdd AOI21X1
XAOI21X1_36 cas INVX2_3/Y NOR2X1_43/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_58 BUFX4_45/Y AND2X2_4/Y NOR2X1_65/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_47 BUFX4_51/Y NOR2X1_50/B NOR2X1_51/Y gnd AOI21X1_47/Y vdd AOI21X1
XFILL_1_3 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_25 MUX2X1_76/B CLKBUF1_20/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_14 MUX2X1_177/A CLKBUF1_56/Y OAI21X1_148/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 MUX2X1_151/B CLKBUF1_37/Y DFFPOSX1_36/D gnd vdd DFFPOSX1
XDFFPOSX1_47 NOR2X1_67/A CLKBUF1_5/A AOI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 INVX1_5/A CLKBUF1_34/Y MUX2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 MUX2X1_100/A CLKBUF1_13/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XFILL_20_2_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XDFFPOSX1_237 INVX1_57/A CLKBUF1_3/Y MUX2X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_259 MUX2X1_193/B CLKBUF1_41/Y OAI21X1_126/Y gnd vdd DFFPOSX1
XDFFPOSX1_248 MUX2X1_106/B CLKBUF1_21/Y OAI21X1_115/Y gnd vdd DFFPOSX1
XDFFPOSX1_226 NOR2X1_36/A CLKBUF1_48/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_204 NAND2X1_98/A CLKBUF1_5/Y OAI21X1_103/Y gnd vdd DFFPOSX1
XDFFPOSX1_215 INVX1_42/A CLKBUF1_28/Y MUX2X1_42/Y gnd vdd DFFPOSX1
XNAND2X1_159 MUX2X1_76/B NAND3X1_11/Y gnd OAI21X1_153/C vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd dataout[6] vdd BUFX2
XNAND2X1_137 rw BUFX2_4/A gnd AOI21X1_41/A vdd NAND2X1
XNAND2X1_115 MUX2X1_130/B OAI21X1_118/B gnd OAI21X1_116/C vdd NAND2X1
XFILL_11_1 gnd vdd FILL
XNAND2X1_126 MUX2X1_217/B NAND3X1_9/Y gnd NAND2X1_126/Y vdd NAND2X1
XNAND2X1_148 AOI22X1_27/Y AOI22X1_28/Y gnd NAND2X1_148/Y vdd NAND2X1
XNAND2X1_104 MUX2X1_96/B NAND3X1_8/Y gnd NAND2X1_104/Y vdd NAND2X1
XOAI21X1_109 BUFX4_48/Y NAND3X1_8/Y OAI21X1_109/C gnd OAI21X1_109/Y vdd OAI21X1
XMUX2X1_198 NOR2X1_7/A NAND2X1_6/A BUFX4_36/Y gnd MUX2X1_198/Y vdd MUX2X1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XMUX2X1_187 MUX2X1_187/A NAND2X1_51/A BUFX4_29/Y gnd MUX2X1_187/Y vdd MUX2X1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XMUX2X1_143 MUX2X1_143/A MUX2X1_143/B BUFX4_16/Y gnd AOI22X1_15/A vdd MUX2X1
XMUX2X1_110 MUX2X1_110/A MUX2X1_108/Y INVX2_6/A gnd AOI22X1_9/D vdd MUX2X1
XMUX2X1_121 NAND2X1_74/A MUX2X1_121/B BUFX4_29/Y gnd MUX2X1_122/A vdd MUX2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XFILL_8_2_1 gnd vdd FILL
XMUX2X1_132 NOR2X1_25/A INVX1_4/A BUFX4_36/Y gnd MUX2X1_134/B vdd MUX2X1
XAOI21X1_7 BUFX4_22/Y NOR2X1_2/B NOR2X1_8/Y gnd AOI21X1_7/Y vdd AOI21X1
XFILL_0_1_1 gnd vdd FILL
XNAND2X1_2 NAND2X1_2/A NAND2X1_1/B gnd OAI21X1_2/C vdd NAND2X1
XMUX2X1_176 MUX2X1_175/Y MUX2X1_174/Y BUFX4_11/Y gnd MUX2X1_176/Y vdd MUX2X1
XMUX2X1_165 INVX1_45/A INVX1_37/A BUFX4_36/Y gnd MUX2X1_165/Y vdd MUX2X1
XMUX2X1_154 MUX2X1_154/A MUX2X1_154/B BUFX4_29/Y gnd MUX2X1_154/Y vdd MUX2X1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_2/B gnd NOR2X1_5/Y vdd NOR2X1
XDFFPOSX1_2 INVX1_60/A CLKBUF1_48/Y MUX2X1_250/Y gnd vdd DFFPOSX1
XAOI21X1_59 BUFX4_2/Y AND2X2_4/Y NOR2X1_66/Y gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_37 cas INVX2_6/Y NOR2X1_44/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_48 BUFX4_9/Y NOR2X1_50/B NOR2X1_52/Y gnd AOI21X1_48/Y vdd AOI21X1
XAOI21X1_26 BUFX4_51/Y NOR2X1_39/B NOR2X1_33/Y gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_15 MUX2X1_7/B AND2X2_2/Y NOR2X1_18/Y gnd AOI21X1_15/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_59 MUX2X1_124/A CLKBUF1_12/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 NOR2X1_68/A CLKBUF1_3/A AOI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 MUX2X1_201/A CLKBUF1_5/A DFFPOSX1_15/D gnd vdd DFFPOSX1
XDFFPOSX1_37 MUX2X1_175/B CLKBUF1_34/Y OAI21X1_165/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 MUX2X1_100/B CLKBUF1_13/Y DFFPOSX1_26/D gnd vdd DFFPOSX1
XDFFPOSX1_227 NOR2X1_37/A CLKBUF1_43/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_238 MUX2X1_72/B CLKBUF1_65/Y OAI21X1_105/Y gnd vdd DFFPOSX1
XDFFPOSX1_249 MUX2X1_130/B CLKBUF1_19/Y OAI21X1_116/Y gnd vdd DFFPOSX1
XDFFPOSX1_216 INVX1_43/A CLKBUF1_23/Y MUX2X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_205 MUX2X1_247/A CLKBUF1_2/Y OAI21X1_104/Y gnd vdd DFFPOSX1
XBUFX2_8 BUFX2_8/A gnd dataout[7] vdd BUFX2
XMUX2X1_177 MUX2X1_177/A NAND2X1_88/A BUFX4_33/Y gnd MUX2X1_179/B vdd MUX2X1
XMUX2X1_199 MUX2X1_199/A MUX2X1_199/B INVX2_3/A gnd MUX2X1_200/A vdd MUX2X1
XNAND2X1_149 rw BUFX2_8/A gnd AOI21X1_45/A vdd NAND2X1
XMUX2X1_111 INVX1_61/A INVX1_11/A BUFX4_33/Y gnd MUX2X1_111/Y vdd MUX2X1
XMUX2X1_188 MUX2X1_187/Y MUX2X1_188/B BUFX4_15/Y gnd AOI22X1_22/D vdd MUX2X1
XNAND2X1_127 MUX2X1_241/B NAND3X1_9/Y gnd NAND2X1_127/Y vdd NAND2X1
XAOI21X1_8 BUFX4_44/Y NOR2X1_2/B NOR2X1_9/Y gnd AOI21X1_8/Y vdd AOI21X1
XNAND2X1_3 NAND2X1_3/A NAND2X1_1/B gnd OAI21X1_3/C vdd NAND2X1
XMUX2X1_144 NOR2X1_53/A MUX2X1_144/B BUFX4_33/Y gnd MUX2X1_146/B vdd MUX2X1
XMUX2X1_122 MUX2X1_122/A MUX2X1_120/Y BUFX4_17/Y gnd AOI22X1_11/D vdd MUX2X1
XNAND2X1_105 MUX2X1_120/B NAND3X1_8/Y gnd OAI21X1_107/C vdd NAND2X1
XNAND2X1_138 AOI22X1_13/Y AOI22X1_14/Y gnd NAND2X1_138/Y vdd NAND2X1
XMUX2X1_155 MUX2X1_154/Y MUX2X1_155/B BUFX4_12/Y gnd AOI22X1_17/A vdd MUX2X1
XNAND2X1_116 MUX2X1_154/B OAI21X1_118/B gnd OAI21X1_117/C vdd NAND2X1
XMUX2X1_100 MUX2X1_100/A MUX2X1_100/B INVX2_3/A gnd MUX2X1_100/Y vdd MUX2X1
XMUX2X1_133 INVX1_20/A MUX2X1_133/B INVX2_3/A gnd MUX2X1_133/Y vdd MUX2X1
XMUX2X1_166 INVX1_54/A NOR2X1_36/A INVX2_3/A gnd MUX2X1_166/Y vdd MUX2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XDFFPOSX1_3 INVX1_61/A CLKBUF1_42/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_2/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B NOR2X1_46/B gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_16 BUFX4_41/Y AND2X2_2/Y NOR2X1_19/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_49 BUFX4_26/Y NOR2X1_50/B NOR2X1_53/Y gnd AOI21X1_49/Y vdd AOI21X1
XAOI21X1_27 BUFX4_8/Y NOR2X1_39/B NOR2X1_34/Y gnd AOI21X1_27/Y vdd AOI21X1
XOAI21X1_90 OR2X2_1/Y BUFX4_46/Y OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XDFFPOSX1_27 MUX2X1_124/B CLKBUF1_9/Y OAI21X1_155/Y gnd vdd DFFPOSX1
XDFFPOSX1_16 MUX2X1_225/A CLKBUF1_3/A OAI21X1_152/Y gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XDFFPOSX1_38 MUX2X1_199/B CLKBUF1_29/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 MUX2X1_78/B CLKBUF1_49/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XDFFPOSX1_206 INVX1_33/A CLKBUF1_67/Y MUX2X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_217 INVX1_44/A CLKBUF1_19/Y MUX2X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_228 NOR2X1_38/A CLKBUF1_38/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_239 MUX2X1_96/B CLKBUF1_14/A OAI21X1_106/Y gnd vdd DFFPOSX1
XFILL_20_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_60 INVX2_4/Y NOR2X1_60/B gnd AND2X2_1/B vdd NOR2X1
XFILL_11_0_0 gnd vdd FILL
XNAND2X1_117 MUX2X1_178/B OAI21X1_118/B gnd NAND2X1_117/Y vdd NAND2X1
XNAND2X1_128 rw BUFX2_1/A gnd AOI21X1_38/A vdd NAND2X1
XAOI21X1_9 BUFX4_58/Y AND2X2_2/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XNAND2X1_139 AOI22X1_15/Y AOI22X1_16/Y gnd NAND2X1_139/Y vdd NAND2X1
XNAND2X1_4 NAND2X1_4/A NAND2X1_1/B gnd OAI21X1_4/C vdd NAND2X1
XNAND2X1_106 MUX2X1_144/B NAND3X1_8/Y gnd OAI21X1_108/C vdd NAND2X1
XMUX2X1_178 MUX2X1_178/A MUX2X1_178/B BUFX4_34/Y gnd MUX2X1_179/A vdd MUX2X1
XMUX2X1_123 NOR2X1_63/A MUX2X1_123/B BUFX4_30/Y gnd MUX2X1_125/B vdd MUX2X1
XMUX2X1_189 INVX1_46/A INVX1_38/A BUFX4_30/Y gnd MUX2X1_191/B vdd MUX2X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_2/B gnd NOR2X1_7/Y vdd NOR2X1
XMUX2X1_112 MUX2X1_112/A INVX1_27/A BUFX4_34/Y gnd MUX2X1_113/A vdd MUX2X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XMUX2X1_145 MUX2X1_145/A MUX2X1_145/B BUFX4_34/Y gnd MUX2X1_145/Y vdd MUX2X1
XDFFPOSX1_4 INVX1_62/A CLKBUF1_38/Y MUX2X1_252/Y gnd vdd DFFPOSX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XMUX2X1_134 MUX2X1_133/Y MUX2X1_134/B INVX2_6/A gnd MUX2X1_134/Y vdd MUX2X1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XMUX2X1_156 NOR2X1_26/A INVX1_5/A BUFX4_30/Y gnd MUX2X1_156/Y vdd MUX2X1
XMUX2X1_167 MUX2X1_166/Y MUX2X1_165/Y BUFX4_16/Y gnd MUX2X1_167/Y vdd MUX2X1
XMUX2X1_101 MUX2X1_100/Y MUX2X1_99/Y BUFX4_18/Y gnd AOI22X1_8/A vdd MUX2X1
XAOI21X1_17 BUFX4_57/Y NOR2X1_22/B NOR2X1_22/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 BUFX4_28/Y NOR2X1_39/B NOR2X1_35/Y gnd AOI21X1_28/Y vdd AOI21X1
XAOI21X1_39 AOI21X1_39/A AOI21X1_39/B NOR2X1_46/B gnd AOI21X1_39/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_80 BUFX4_43/Y NAND2X1_88/B OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 OR2X2_1/A INVX8_1/A MUX2X1_181/B gnd OAI21X1_92/C vdd OAI21X1
XFILL_23_2_1 gnd vdd FILL
XDFFPOSX1_17 NOR2X1_50/A CLKBUF1_50/Y AOI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 MUX2X1_148/B CLKBUF1_5/Y OAI21X1_156/Y gnd vdd DFFPOSX1
XDFFPOSX1_39 MUX2X1_223/B CLKBUF1_27/Y OAI21X1_167/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XDFFPOSX1_229 NOR2X1_39/A CLKBUF1_33/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_218 INVX1_45/A CLKBUF1_14/Y MUX2X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_207 INVX1_34/A CLKBUF1_25/A MUX2X1_34/Y gnd vdd DFFPOSX1
XFILL_20_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_61 MUX2X1_75/A AND2X2_4/Y gnd NOR2X1_61/Y vdd NOR2X1
XNOR2X1_50 NOR2X1_50/A NOR2X1_50/B gnd NOR2X1_50/Y vdd NOR2X1
XFILL_19_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND2X1_129 AOI22X1_1/Y AOI22X1_2/Y gnd OAI21X1_129/A vdd NAND2X1
XNAND2X1_118 MUX2X1_202/B OAI21X1_118/B gnd OAI21X1_119/C vdd NAND2X1
XNAND2X1_5 NAND2X1_5/A NAND2X1_1/B gnd OAI21X1_5/C vdd NAND2X1
XMUX2X1_90 MUX2X1_90/A MUX2X1_90/B BUFX4_30/Y gnd MUX2X1_90/Y vdd MUX2X1
XNAND2X1_107 MUX2X1_168/B NAND3X1_8/Y gnd OAI21X1_109/C vdd NAND2X1
XMUX2X1_124 MUX2X1_124/A MUX2X1_124/B BUFX4_31/Y gnd MUX2X1_125/A vdd MUX2X1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XMUX2X1_179 MUX2X1_179/A MUX2X1_179/B BUFX4_12/Y gnd AOI22X1_21/A vdd MUX2X1
XMUX2X1_113 MUX2X1_113/A MUX2X1_111/Y BUFX4_14/Y gnd AOI22X1_10/A vdd MUX2X1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XMUX2X1_146 MUX2X1_145/Y MUX2X1_146/B BUFX4_17/Y gnd MUX2X1_146/Y vdd MUX2X1
XMUX2X1_135 INVX1_62/A INVX1_12/A BUFX4_38/Y gnd MUX2X1_135/Y vdd MUX2X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XDFFPOSX1_5 INVX1_63/A CLKBUF1_34/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XMUX2X1_102 NOR2X1_3/A NAND2X1_2/A BUFX4_38/Y gnd MUX2X1_102/Y vdd MUX2X1
XMUX2X1_157 INVX1_21/A OAI21X1_89/C BUFX4_31/Y gnd MUX2X1_157/Y vdd MUX2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XMUX2X1_168 NOR2X1_54/A MUX2X1_168/B BUFX4_38/Y gnd MUX2X1_168/Y vdd MUX2X1
XAOI21X1_29 BUFX4_48/Y NOR2X1_39/B NOR2X1_36/Y gnd AOI21X1_29/Y vdd AOI21X1
XNOR2X1_8 NOR2X1_8/A NOR2X1_2/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 MUX2X1_2/B NOR2X1_22/B NOR2X1_23/Y gnd AOI21X1_18/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_70 BUFX4_1/Y NAND3X1_6/Y NAND2X1_77/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 OR2X2_1/Y BUFX4_4/Y OAI21X1_92/C gnd OAI21X1_92/Y vdd OAI21X1
XOAI21X1_81 OR2X2_1/A INVX8_1/A MUX2X1_61/B gnd OAI21X1_82/C vdd OAI21X1
XDFFPOSX1_29 MUX2X1_172/B CLKBUF1_2/Y DFFPOSX1_29/D gnd vdd DFFPOSX1
XDFFPOSX1_18 NOR2X1_51/A CLKBUF1_48/Y AOI21X1_47/Y gnd vdd DFFPOSX1
XCLKBUF1_60 clk gnd CLKBUF1_41/A vdd CLKBUF1
XDFFPOSX1_219 INVX1_46/A CLKBUF1_9/Y MUX2X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_208 INVX1_35/A CLKBUF1_14/A MUX2X1_35/Y gnd vdd DFFPOSX1
XNAND2X1_108 MUX2X1_192/B NAND3X1_8/Y gnd NAND2X1_108/Y vdd NAND2X1
XNAND2X1_119 MUX2X1_226/B OAI21X1_118/B gnd OAI21X1_120/C vdd NAND2X1
XNAND2X1_6 NAND2X1_6/A NAND2X1_1/B gnd OAI21X1_6/C vdd NAND2X1
XNOR2X1_40 ras address[2] gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_62 NOR2X1_62/A AND2X2_4/Y gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_51 NOR2X1_51/A NOR2X1_50/B gnd NOR2X1_51/Y vdd NOR2X1
XMUX2X1_125 MUX2X1_125/A MUX2X1_125/B BUFX4_18/Y gnd AOI22X1_12/A vdd MUX2X1
XFILL_21_3_0 gnd vdd FILL
XMUX2X1_80 MUX2X1_80/A MUX2X1_80/B BUFX4_11/Y gnd AOI22X1_4/D vdd MUX2X1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XMUX2X1_114 NOR2X1_14/A MUX2X1_114/B BUFX4_35/Y gnd MUX2X1_116/B vdd MUX2X1
XDFFPOSX1_6 INVX1_64/A CLKBUF1_30/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XMUX2X1_147 NOR2X1_64/A NAND2X1_23/A BUFX4_35/Y gnd MUX2X1_147/Y vdd MUX2X1
XMUX2X1_136 MUX2X1_136/A INVX1_28/A BUFX4_39/Y gnd MUX2X1_136/Y vdd MUX2X1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XMUX2X1_103 MUX2X1_103/A MUX2X1_103/B BUFX4_39/Y gnd MUX2X1_103/Y vdd MUX2X1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XMUX2X1_91 MUX2X1_91/A MUX2X1_91/B BUFX4_31/Y gnd MUX2X1_91/Y vdd MUX2X1
XMUX2X1_169 MUX2X1_169/A MUX2X1_169/B BUFX4_39/Y gnd MUX2X1_169/Y vdd MUX2X1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XMUX2X1_158 MUX2X1_157/Y MUX2X1_156/Y INVX2_6/A gnd MUX2X1_158/Y vdd MUX2X1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_2/B gnd NOR2X1_9/Y vdd NOR2X1
XFILL_12_3_0 gnd vdd FILL
XAOI21X1_19 BUFX4_6/Y NOR2X1_22/B NOR2X1_24/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_82 OR2X2_1/Y MUX2X1_9/B OAI21X1_82/C gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_60 BUFX4_24/Y NAND2X1_64/B NAND2X1_67/Y gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_71 BUFX4_19/Y NAND3X1_6/Y NAND2X1_78/Y gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_93 OR2X2_1/A INVX8_1/A MUX2X1_205/B gnd OAI21X1_93/Y vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XDFFPOSX1_19 NOR2X1_52/A CLKBUF1_41/Y AOI21X1_48/Y gnd vdd DFFPOSX1
XCLKBUF1_50 CLKBUF1_9/A gnd CLKBUF1_50/Y vdd CLKBUF1
XCLKBUF1_61 clk gnd CLKBUF1_27/A vdd CLKBUF1
XFILL_23_0_0 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XDFFPOSX1_209 INVX1_36/A CLKBUF1_51/Y MUX2X1_36/Y gnd vdd DFFPOSX1
XNOR2X1_63 NOR2X1_63/A AND2X2_4/Y gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 NOR2X1_52/A NOR2X1_50/B gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_30 INVX2_4/A OR2X2_2/A gnd INVX1_49/A vdd NOR2X1
XNOR2X1_41 ras address[3] gnd NOR2X1_41/Y vdd NOR2X1
XNAND2X1_109 MUX2X1_216/B NAND3X1_8/Y gnd OAI21X1_111/C vdd NAND2X1
XNAND2X1_7 NAND2X1_7/A NAND2X1_1/B gnd OAI21X1_7/C vdd NAND2X1
XFILL_21_3_1 gnd vdd FILL
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XMUX2X1_70 INVX1_50/A NOR2X1_32/A BUFX4_39/Y gnd MUX2X1_70/Y vdd MUX2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XMUX2X1_115 NAND2X1_32/A MUX2X1_115/B BUFX4_36/Y gnd MUX2X1_116/A vdd MUX2X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XMUX2X1_126 NOR2X1_4/A NAND2X1_3/A BUFX4_32/Y gnd MUX2X1_128/B vdd MUX2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XMUX2X1_148 MUX2X1_148/A MUX2X1_148/B BUFX4_36/Y gnd MUX2X1_148/Y vdd MUX2X1
XMUX2X1_137 MUX2X1_136/Y MUX2X1_135/Y BUFX4_14/Y gnd MUX2X1_137/Y vdd MUX2X1
XMUX2X1_81 MUX2X1_81/A MUX2X1_81/B BUFX4_35/Y gnd MUX2X1_83/B vdd MUX2X1
XMUX2X1_104 MUX2X1_103/Y MUX2X1_102/Y BUFX4_11/Y gnd AOI22X1_8/D vdd MUX2X1
XMUX2X1_159 INVX1_63/A INVX1_13/A BUFX4_32/Y gnd MUX2X1_159/Y vdd MUX2X1
XMUX2X1_92 MUX2X1_91/Y MUX2X1_90/Y BUFX4_15/Y gnd MUX2X1_92/Y vdd MUX2X1
XFILL_12_3_1 gnd vdd FILL
XDFFPOSX1_7 INVX1_65/A CLKBUF1_27/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XOAI21X1_72 BUFX4_42/Y NAND3X1_6/Y NAND2X1_79/Y gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_94 OR2X2_1/Y MUX2X1_7/B OAI21X1_93/Y gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_50 BUFX4_50/Y NAND2X1_56/B OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 BUFX4_47/Y NAND2X1_64/B OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_83 OR2X2_1/A INVX8_1/A MUX2X1_85/B gnd OAI21X1_84/C vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XFILL_9_3_1 gnd vdd FILL
XCLKBUF1_40 CLKBUF1_56/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XCLKBUF1_51 CLKBUF1_67/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XCLKBUF1_62 clk gnd CLKBUF1_14/A vdd CLKBUF1
XFILL_23_0_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_20 INVX8_11/A INVX2_2/Y gnd NOR2X1_20/Y vdd NOR2X1
XNOR2X1_53 NOR2X1_53/A NOR2X1_50/B gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_42 ras address[4] gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A AND2X2_4/Y gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_31 INVX1_49/Y OR2X2_1/A gnd NOR2X1_39/B vdd NOR2X1
XMUX2X1_60 MUX2X1_60/A INVX1_1/A BUFX4_32/Y gnd MUX2X1_62/B vdd MUX2X1
XMUX2X1_71 MUX2X1_70/Y MUX2X1_71/B BUFX4_16/Y gnd AOI22X1_3/A vdd MUX2X1
XMUX2X1_105 MUX2X1_105/A NAND2X1_85/A BUFX4_29/Y gnd MUX2X1_107/B vdd MUX2X1
XMUX2X1_116 MUX2X1_116/A MUX2X1_116/B BUFX4_15/Y gnd AOI22X1_10/D vdd MUX2X1
XNAND2X1_8 NAND2X1_8/A NAND2X1_1/B gnd OAI21X1_8/C vdd NAND2X1
XMUX2X1_149 MUX2X1_148/Y MUX2X1_147/Y BUFX4_18/Y gnd AOI22X1_16/A vdd MUX2X1
XMUX2X1_138 NOR2X1_15/A NAND2X1_58/A BUFX4_29/Y gnd MUX2X1_140/B vdd MUX2X1
XMUX2X1_127 NAND2X1_94/A MUX2X1_127/B BUFX4_33/Y gnd MUX2X1_127/Y vdd MUX2X1
XMUX2X1_82 MUX2X1_82/A MUX2X1_82/B BUFX4_36/Y gnd MUX2X1_82/Y vdd MUX2X1
XMUX2X1_93 INVX1_42/A INVX1_34/A BUFX4_32/Y gnd MUX2X1_93/Y vdd MUX2X1
XDFFPOSX1_8 INVX1_66/A CLKBUF1_22/Y MUX2X1_256/Y gnd vdd DFFPOSX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XOAI21X1_73 BUFX4_57/Y NAND2X1_88/B NAND2X1_83/Y gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_40 BUFX4_43/Y NAND3X1_4/Y NAND2X1_45/Y gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_51 BUFX4_7/Y NAND2X1_56/B NAND2X1_57/Y gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_95 OR2X2_1/A INVX8_1/A MUX2X1_229/B gnd OAI21X1_96/C vdd OAI21X1
XOAI21X1_62 BUFX4_2/Y NAND2X1_64/B NAND2X1_69/Y gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_84 OR2X2_1/Y MUX2X1_2/B OAI21X1_84/C gnd OAI21X1_84/Y vdd OAI21X1
XDFFPOSX1_190 NOR2X1_24/A CLKBUF1_5/A AOI21X1_19/Y gnd vdd DFFPOSX1
XCLKBUF1_63 clk gnd CLKBUF1_9/A vdd CLKBUF1
XCLKBUF1_52 CLKBUF1_56/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XCLKBUF1_30 CLKBUF1_65/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XCLKBUF1_41 CLKBUF1_41/A gnd CLKBUF1_41/Y vdd CLKBUF1
XFILL_18_1 gnd vdd FILL
XNOR2X1_32 NOR2X1_32/A NOR2X1_39/B gnd NOR2X1_32/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNOR2X1_43 cas address[0] gnd NOR2X1_43/Y vdd NOR2X1
XNAND3X1_10 ras en cas gnd NOR2X1_46/B vdd NAND3X1
XNOR2X1_21 INVX8_1/A INVX2_5/A gnd NOR2X1_22/B vdd NOR2X1
XNOR2X1_10 INVX2_4/Y NOR2X1_47/B gnd AND2X2_2/B vdd NOR2X1
XNOR2X1_54 NOR2X1_54/A NOR2X1_50/B gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_65 NOR2X1_65/A AND2X2_4/Y gnd NOR2X1_65/Y vdd NOR2X1
XMUX2X1_72 NOR2X1_50/A MUX2X1_72/B BUFX4_29/Y gnd MUX2X1_74/B vdd MUX2X1
XMUX2X1_61 INVX1_17/A MUX2X1_61/B BUFX4_33/Y gnd MUX2X1_61/Y vdd MUX2X1
XNAND2X1_9 BUFX4_29/Y BUFX4_11/Y gnd INVX2_1/A vdd NAND2X1
XMUX2X1_83 MUX2X1_82/Y MUX2X1_83/B BUFX4_12/Y gnd AOI22X1_5/A vdd MUX2X1
XMUX2X1_94 INVX1_51/A NOR2X1_33/A BUFX4_33/Y gnd MUX2X1_94/Y vdd MUX2X1
XMUX2X1_50 INVX1_51/Y BUFX4_54/Y MUX2X1_56/S gnd MUX2X1_50/Y vdd MUX2X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XDFFPOSX1_9 MUX2X1_57/A CLKBUF1_17/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XMUX2X1_128 MUX2X1_127/Y MUX2X1_128/B BUFX4_11/Y gnd MUX2X1_128/Y vdd MUX2X1
XMUX2X1_106 MUX2X1_106/A MUX2X1_106/B BUFX4_30/Y gnd MUX2X1_107/A vdd MUX2X1
XMUX2X1_117 INVX1_43/A INVX1_35/A INVX2_3/A gnd MUX2X1_117/Y vdd MUX2X1
XMUX2X1_139 MUX2X1_139/A MUX2X1_139/B BUFX4_30/Y gnd MUX2X1_139/Y vdd MUX2X1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XFILL_21_1_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_41 BUFX4_58/Y NAND3X1_5/Y NAND2X1_46/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_30 BUFX4_4/Y OAI21X1_25/B NAND2X1_35/Y gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_96 OR2X2_1/Y BUFX4_41/Y OAI21X1_96/C gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_85 OR2X2_1/A INVX8_1/A MUX2X1_109/B gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_52 BUFX4_25/Y NAND2X1_56/B OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_63 BUFX4_21/Y NAND2X1_64/B OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_74 BUFX4_50/Y NAND2X1_88/B OAI21X1_74/C gnd OAI21X1_74/Y vdd OAI21X1
XDFFPOSX1_180 MUX2X1_61/B CLKBUF1_37/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_191 NOR2X1_25/A CLKBUF1_8/A AOI21X1_20/Y gnd vdd DFFPOSX1
XFILL_6_1 gnd vdd FILL
XCLKBUF1_20 CLKBUF1_9/A gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_64 clk gnd CLKBUF1_3/A vdd CLKBUF1
XCLKBUF1_31 CLKBUF1_5/A gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_42 CLKBUF1_5/A gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_53 clk gnd CLKBUF1_4/A vdd CLKBUF1
XFILL_1_0_0 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XFILL_18_2 gnd vdd FILL
XNOR2X1_22 MUX2X1_60/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_55 NOR2X1_55/A NOR2X1_50/B gnd NOR2X1_55/Y vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_66 NOR2X1_66/A AND2X2_4/Y gnd NOR2X1_66/Y vdd NOR2X1
XNAND3X1_11 INVX2_2/A NAND3X1_5/B AND2X2_4/B gnd NAND3X1_11/Y vdd NAND3X1
XNOR2X1_11 INVX2_1/A INVX2_2/Y gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_44 cas address[1] gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_39/B gnd NOR2X1_33/Y vdd NOR2X1
XMUX2X1_40 INVX1_40/Y BUFX4_40/Y MUX2X1_39/S gnd MUX2X1_40/Y vdd MUX2X1
XMUX2X1_62 MUX2X1_61/Y MUX2X1_62/B INVX2_6/A gnd AOI22X1_1/D vdd MUX2X1
XMUX2X1_73 MUX2X1_73/A MUX2X1_73/B BUFX4_30/Y gnd MUX2X1_73/Y vdd MUX2X1
XMUX2X1_51 INVX1_52/Y BUFX4_8/Y MUX2X1_56/S gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_84 MUX2X1_84/A INVX1_2/A INVX2_3/A gnd MUX2X1_84/Y vdd MUX2X1
XMUX2X1_95 MUX2X1_94/Y MUX2X1_93/Y BUFX4_16/Y gnd MUX2X1_95/Y vdd MUX2X1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XMUX2X1_107 MUX2X1_107/A MUX2X1_107/B BUFX4_12/Y gnd AOI22X1_9/A vdd MUX2X1
XMUX2X1_118 INVX1_52/A NOR2X1_34/A BUFX4_38/Y gnd MUX2X1_118/Y vdd MUX2X1
XMUX2X1_129 MUX2X1_129/A NAND2X1_86/A BUFX4_34/Y gnd MUX2X1_131/B vdd MUX2X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XFILL_21_1_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XOAI21X1_75 BUFX4_10/Y NAND2X1_88/B OAI21X1_75/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_97 BUFX4_55/Y NAND3X1_7/Y OAI21X1_97/C gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_64 BUFX4_40/Y NAND2X1_64/B NAND2X1_71/Y gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_86 OR2X2_1/Y BUFX4_6/Y OAI21X1_85/Y gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_20 BUFX4_25/Y NAND3X1_3/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_53 BUFX4_45/Y NAND2X1_56/B OAI21X1_53/C gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_42 BUFX4_50/Y NAND3X1_5/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_31 BUFX4_23/Y OAI21X1_25/B NAND2X1_36/Y gnd OAI21X1_31/Y vdd OAI21X1
XDFFPOSX1_170 INVX1_31/A CLKBUF1_16/Y MUX2X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_192 NOR2X1_26/A CLKBUF1_27/A AOI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_181 MUX2X1_85/B CLKBUF1_36/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XFILL_6_2 gnd vdd FILL
XCLKBUF1_54 clk gnd CLKBUF1_7/A vdd CLKBUF1
XCLKBUF1_43 CLKBUF1_9/A gnd CLKBUF1_43/Y vdd CLKBUF1
XCLKBUF1_65 clk gnd CLKBUF1_65/Y vdd CLKBUF1
XCLKBUF1_10 CLKBUF1_56/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XCLKBUF1_32 CLKBUF1_5/A gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_21 CLKBUF1_4/A gnd CLKBUF1_21/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XFILL_18_3 gnd vdd FILL
XNOR2X1_12 MUX2X1_66/A AND2X2_2/Y gnd AOI21X1_9/C vdd NOR2X1
XNAND3X1_12 INVX2_2/A NAND3X1_5/B AND2X2_1/B gnd NAND3X1_12/Y vdd NAND3X1
XMUX2X1_52 INVX1_53/Y BUFX4_28/Y MUX2X1_56/S gnd MUX2X1_52/Y vdd MUX2X1
XMUX2X1_41 INVX1_41/Y BUFX4_56/Y MUX2X1_46/S gnd MUX2X1_41/Y vdd MUX2X1
XMUX2X1_63 INVX1_58/A INVX1_9/A BUFX4_34/Y gnd MUX2X1_65/B vdd MUX2X1
XMUX2X1_30 INVX1_30/Y BUFX4_2/Y MUX2X1_27/S gnd MUX2X1_30/Y vdd MUX2X1
XNOR2X1_45 BUFX4_12/Y INVX2_3/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_39/B gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_56 NOR2X1_56/A NOR2X1_50/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A AND2X2_4/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_23 MUX2X1_84/A NOR2X1_22/B gnd NOR2X1_23/Y vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XMUX2X1_74 MUX2X1_73/Y MUX2X1_74/B BUFX4_17/Y gnd MUX2X1_74/Y vdd MUX2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XMUX2X1_108 NOR2X1_24/A INVX1_3/A BUFX4_31/Y gnd MUX2X1_108/Y vdd MUX2X1
XMUX2X1_119 MUX2X1_118/Y MUX2X1_117/Y BUFX4_16/Y gnd MUX2X1_119/Y vdd MUX2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XMUX2X1_85 INVX1_18/A MUX2X1_85/B BUFX4_38/Y gnd MUX2X1_85/Y vdd MUX2X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XMUX2X1_96 NOR2X1_51/A MUX2X1_96/B BUFX4_34/Y gnd MUX2X1_96/Y vdd MUX2X1
XOAI21X1_54 BUFX4_4/Y NAND2X1_56/B NAND2X1_60/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_32 BUFX4_41/Y OAI21X1_25/B NAND2X1_37/Y gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_65 BUFX4_56/Y NAND3X1_6/Y OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_43 BUFX4_6/Y NAND3X1_5/Y NAND2X1_48/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_76 BUFX4_25/Y NAND2X1_88/B NAND2X1_86/Y gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_98 BUFX4_54/Y NAND3X1_7/Y NAND2X1_93/Y gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_10 BUFX4_52/Y OAI21X1_9/B OAI21X1_10/C gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_87 OR2X2_1/A INVX8_1/A MUX2X1_133/B gnd OAI21X1_88/C vdd OAI21X1
XOAI21X1_21 BUFX4_46/Y NAND3X1_3/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XDFFPOSX1_193 NOR2X1_27/A CLKBUF1_52/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_171 INVX1_32/A CLKBUF1_11/Y MUX2X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_182 MUX2X1_109/B CLKBUF1_32/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_160 INVX1_21/A CLKBUF1_27/A MUX2X1_21/Y gnd vdd DFFPOSX1
XCLKBUF1_33 CLKBUF1_67/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_44 CLKBUF1_67/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XCLKBUF1_11 CLKBUF1_67/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XCLKBUF1_22 CLKBUF1_67/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_66 clk gnd CLKBUF1_2/A vdd CLKBUF1
XCLKBUF1_55 clk gnd CLKBUF1_1/A vdd CLKBUF1
XFILL_10_2_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_18_3_0 gnd vdd FILL
XNOR2X1_68 NOR2X1_68/A AND2X2_4/Y gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_35 NOR2X1_35/A NOR2X1_39/B gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_57 NOR2X1_57/A NOR2X1_50/B gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_46 INVX4_1/Y NOR2X1_46/B gnd INVX2_2/A vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A NOR2X1_22/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_13 MUX2X1_90/A AND2X2_2/Y gnd NOR2X1_13/Y vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XMUX2X1_75 MUX2X1_75/A MUX2X1_75/B BUFX4_31/Y gnd MUX2X1_77/B vdd MUX2X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XMUX2X1_64 MUX2X1_64/A INVX1_25/A BUFX4_35/Y gnd MUX2X1_65/A vdd MUX2X1
XMUX2X1_109 INVX1_19/A MUX2X1_109/B BUFX4_32/Y gnd MUX2X1_110/A vdd MUX2X1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XMUX2X1_31 INVX1_31/Y BUFX4_21/Y MUX2X1_27/S gnd MUX2X1_31/Y vdd MUX2X1
XMUX2X1_42 INVX1_42/Y BUFX4_54/Y MUX2X1_46/S gnd MUX2X1_42/Y vdd MUX2X1
XMUX2X1_20 INVX1_20/Y BUFX4_27/Y MUX2X1_17/S gnd MUX2X1_20/Y vdd MUX2X1
XMUX2X1_53 INVX1_54/Y BUFX4_48/Y MUX2X1_56/S gnd MUX2X1_53/Y vdd MUX2X1
XMUX2X1_86 MUX2X1_85/Y MUX2X1_84/Y INVX2_6/A gnd MUX2X1_86/Y vdd MUX2X1
XMUX2X1_97 MUX2X1_97/A MUX2X1_97/B BUFX4_35/Y gnd MUX2X1_98/A vdd MUX2X1
XNAND2X1_90 NAND2X1_90/A NAND2X1_88/B gnd OAI21X1_80/C vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_11 BUFX4_10/Y OAI21X1_9/B NAND2X1_12/Y gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_33 BUFX4_58/Y NAND3X1_4/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_22 BUFX4_2/Y NAND3X1_3/Y NAND2X1_25/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_44 BUFX4_25/Y NAND3X1_5/Y NAND2X1_49/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_99 BUFX4_8/Y NAND3X1_7/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_77 BUFX4_45/Y NAND2X1_88/B NAND2X1_87/Y gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_55 MUX2X1_7/B NAND2X1_56/B OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_66 BUFX4_54/Y NAND3X1_6/Y NAND2X1_73/Y gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_88 OR2X2_1/Y BUFX4_27/Y OAI21X1_88/C gnd OAI21X1_88/Y vdd OAI21X1
XDFFPOSX1_172 MUX2X1_57/B CLKBUF1_7/Y OAI21X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_161 INVX1_22/A CLKBUF1_49/Y MUX2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_150 NAND2X1_74/A CLKBUF1_30/Y OAI21X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_194 NOR2X1_28/A CLKBUF1_45/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XFILL_4_0_0 gnd vdd FILL
XDFFPOSX1_183 MUX2X1_133/B CLKBUF1_25/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XCLKBUF1_56 clk gnd CLKBUF1_56/Y vdd CLKBUF1
XCLKBUF1_12 CLKBUF1_7/A gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_23 CLKBUF1_67/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_45 CLKBUF1_2/A gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_34 CLKBUF1_35/A gnd CLKBUF1_34/Y vdd CLKBUF1
XCLKBUF1_67 clk gnd CLKBUF1_67/Y vdd CLKBUF1
XFILL_4_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_14 NOR2X1_14/A AND2X2_2/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_58 BUFX4_38/Y INVX2_6/Y gnd NAND3X1_5/B vdd NOR2X1
XNOR2X1_47 INVX2_4/A NOR2X1_47/B gnd AND2X2_3/A vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_22/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_36 NOR2X1_36/A NOR2X1_39/B gnd NOR2X1_36/Y vdd NOR2X1
XMUX2X1_76 MUX2X1_76/A MUX2X1_76/B BUFX4_32/Y gnd MUX2X1_77/A vdd MUX2X1
XMUX2X1_54 INVX1_55/Y BUFX4_1/Y MUX2X1_56/S gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_32 INVX1_32/Y BUFX4_42/Y MUX2X1_27/S gnd MUX2X1_32/Y vdd MUX2X1
XMUX2X1_65 MUX2X1_65/A MUX2X1_65/B BUFX4_14/Y gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_43 INVX1_43/Y BUFX4_8/Y MUX2X1_46/S gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_87 INVX1_60/A INVX1_10/A BUFX4_39/Y gnd MUX2X1_87/Y vdd MUX2X1
XMUX2X1_21 INVX1_21/Y MUX2X1_5/B MUX2X1_17/S gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_98 MUX2X1_98/A MUX2X1_96/Y BUFX4_17/Y gnd AOI22X1_7/D vdd MUX2X1
XMUX2X1_10 INVX1_10/Y BUFX4_52/Y MUX2X1_9/S gnd MUX2X1_10/Y vdd MUX2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XNAND2X1_80 INVX8_1/Y NOR2X1_11/Y gnd MUX2X1_17/S vdd NAND2X1
XNAND2X1_91 NAND3X1_5/B INVX2_2/A gnd OR2X2_1/A vdd NAND2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_12 BUFX4_25/Y OAI21X1_9/B NAND2X1_13/Y gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_23 BUFX4_23/Y NAND3X1_3/Y NAND2X1_26/Y gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_34 BUFX4_50/Y NAND3X1_4/Y NAND2X1_39/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 BUFX4_45/Y NAND3X1_5/Y NAND2X1_50/Y gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_78 BUFX4_5/Y NAND2X1_88/B OAI21X1_78/C gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_56 BUFX4_43/Y NAND2X1_56/B OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_67 BUFX4_9/Y NAND3X1_6/Y OAI21X1_67/C gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_89 OR2X2_1/A INVX8_1/A OAI21X1_89/C gnd OAI21X1_90/C vdd OAI21X1
XDFFPOSX1_140 MUX2X1_64/A CLKBUF1_7/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_195 NOR2X1_29/A CLKBUF1_44/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_151 MUX2X1_145/A CLKBUF1_25/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 INVX1_23/A CLKBUF1_45/Y MUX2X1_23/Y gnd vdd DFFPOSX1
XFILL_4_0_1 gnd vdd FILL
XDFFPOSX1_184 OAI21X1_89/C CLKBUF1_24/Y OAI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_173 MUX2X1_81/B CLKBUF1_4/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XCLKBUF1_68 clk gnd CLKBUF1_5/A vdd CLKBUF1
XCLKBUF1_35 CLKBUF1_35/A gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_24 CLKBUF1_35/A gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_57 clk gnd CLKBUF1_25/A vdd CLKBUF1
XCLKBUF1_46 CLKBUF1_1/A gnd CLKBUF1_46/Y vdd CLKBUF1
XCLKBUF1_13 CLKBUF1_2/A gnd CLKBUF1_13/Y vdd CLKBUF1
XNOR2X1_37 NOR2X1_37/A NOR2X1_39/B gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_59 INVX2_4/A NOR2X1_60/B gnd AND2X2_4/B vdd NOR2X1
XNOR2X1_48 INVX1_67/A INVX1_59/A gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_15 NOR2X1_15/A AND2X2_2/Y gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A NOR2X1_22/B gnd NOR2X1_26/Y vdd NOR2X1
XMUX2X1_77 MUX2X1_77/A MUX2X1_77/B BUFX4_18/Y gnd AOI22X1_4/A vdd MUX2X1
XMUX2X1_33 INVX1_33/Y BUFX4_56/Y MUX2X1_39/S gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_22 INVX1_22/Y BUFX4_4/Y MUX2X1_17/S gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_11 INVX1_11/Y BUFX4_7/Y MUX2X1_9/S gnd MUX2X1_11/Y vdd MUX2X1
XMUX2X1_66 MUX2X1_66/A MUX2X1_66/B BUFX4_36/Y gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_44 INVX1_44/Y BUFX4_26/Y MUX2X1_46/S gnd MUX2X1_44/Y vdd MUX2X1
XMUX2X1_55 INVX1_56/Y BUFX4_19/Y MUX2X1_56/S gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_88 MUX2X1_88/A INVX1_26/A BUFX4_29/Y gnd MUX2X1_88/Y vdd MUX2X1
XMUX2X1_99 NOR2X1_62/A MUX2X1_99/B BUFX4_36/Y gnd MUX2X1_99/Y vdd MUX2X1
XNAND2X1_92 MUX2X1_79/A NAND3X1_7/Y gnd OAI21X1_97/C vdd NAND2X1
XNAND2X1_81 NAND3X1_5/B AND2X2_3/Y gnd MUX2X1_27/S vdd NAND2X1
XNAND2X1_70 NAND2X1_70/A NAND2X1_64/B gnd OAI21X1_63/C vdd NAND2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XFILL_21_1 gnd vdd FILL
XOAI21X1_24 BUFX4_43/Y NAND3X1_3/Y NAND2X1_27/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_57 MUX2X1_9/B NAND2X1_64/B OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_46 BUFX4_4/Y NAND3X1_5/Y OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_35 BUFX4_6/Y NAND3X1_4/Y NAND2X1_40/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_68 BUFX4_26/Y NAND3X1_6/Y NAND2X1_75/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_13 BUFX4_46/Y OAI21X1_9/B NAND2X1_14/Y gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_79 BUFX4_23/Y NAND2X1_88/B OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XDFFPOSX1_174 NAND2X1_85/A CLKBUF1_7/A OAI21X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_163 INVX1_24/A CLKBUF1_44/Y MUX2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_185 MUX2X1_181/B CLKBUF1_18/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_196 BUFX4_34/A CLKBUF1_40/Y AOI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 MUX2X1_169/A CLKBUF1_24/Y OAI21X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_130 NOR2X1_18/A CLKBUF1_46/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_141 MUX2X1_88/A CLKBUF1_2/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XMUX2X1_250 INVX1_60/Y BUFX4_51/Y MUX2X1_249/S gnd MUX2X1_250/Y vdd MUX2X1
XFILL_22_2_0 gnd vdd FILL
XCLKBUF1_58 clk gnd CLKBUF1_8/A vdd CLKBUF1
XCLKBUF1_36 CLKBUF1_1/A gnd CLKBUF1_36/Y vdd CLKBUF1
XCLKBUF1_47 CLKBUF1_25/A gnd CLKBUF1_47/Y vdd CLKBUF1
XCLKBUF1_25 CLKBUF1_25/A gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_14 CLKBUF1_14/A gnd CLKBUF1_14/Y vdd CLKBUF1
XFILL_13_2_0 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XNOR2X1_27 NOR2X1_27/A NOR2X1_22/B gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_49 OR2X2_2/Y INVX2_5/A gnd NOR2X1_50/B vdd NOR2X1
XNOR2X1_38 NOR2X1_38/A NOR2X1_39/B gnd NOR2X1_38/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_16 NOR2X1_16/A AND2X2_2/Y gnd NOR2X1_16/Y vdd NOR2X1
XMUX2X1_56 INVX1_57/Y BUFX4_40/Y MUX2X1_56/S gnd MUX2X1_56/Y vdd MUX2X1
XMUX2X1_78 NOR2X1_2/A MUX2X1_78/B BUFX4_33/Y gnd MUX2X1_80/B vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_67 MUX2X1_67/A MUX2X1_67/B INVX2_3/A gnd MUX2X1_68/A vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XMUX2X1_12 INVX1_12/Y BUFX4_24/Y MUX2X1_9/S gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_45 INVX1_45/Y BUFX4_48/Y MUX2X1_46/S gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_89 MUX2X1_88/Y MUX2X1_87/Y BUFX4_14/Y gnd MUX2X1_89/Y vdd MUX2X1
XMUX2X1_23 INVX1_23/Y MUX2X1_7/B MUX2X1_17/S gnd MUX2X1_23/Y vdd MUX2X1
XMUX2X1_34 INVX1_34/Y BUFX4_51/Y MUX2X1_39/S gnd MUX2X1_34/Y vdd MUX2X1
XNAND2X1_60 MUX2X1_186/B NAND2X1_56/B gnd NAND2X1_60/Y vdd NAND2X1
XNAND2X1_71 MUX2X1_232/A NAND2X1_64/B gnd NAND2X1_71/Y vdd NAND2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_82 INVX2_7/Y NOR2X1_20/Y gnd NAND2X1_88/B vdd NAND2X1
XNAND2X1_93 MUX2X1_103/A NAND3X1_7/Y gnd NAND2X1_93/Y vdd NAND2X1
XFILL_21_2 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_14 BUFX4_2/Y OAI21X1_9/B NAND2X1_15/Y gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_25 BUFX4_58/Y OAI21X1_25/B NAND2X1_30/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_36 BUFX4_24/Y NAND3X1_4/Y OAI21X1_36/C gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_69 BUFX4_47/Y NAND3X1_6/Y OAI21X1_69/C gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_58 BUFX4_52/Y NAND2X1_64/B OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_47 BUFX4_23/Y NAND3X1_5/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XDFFPOSX1_142 MUX2X1_112/A CLKBUF1_5/A OAI21X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 MUX2X1_193/A CLKBUF1_20/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_164 INVX1_25/A CLKBUF1_37/Y MUX2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 NOR2X1_19/A CLKBUF1_42/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_197 BUFX4_12/A CLKBUF1_33/Y AOI21X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_175 NAND2X1_86/A CLKBUF1_5/A OAI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 MUX2X1_163/B CLKBUF1_21/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_186 MUX2X1_205/B CLKBUF1_16/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XMUX2X1_240 NOR2X1_57/A MUX2X1_240/B BUFX4_31/Y gnd MUX2X1_240/Y vdd MUX2X1
XMUX2X1_251 INVX1_61/Y BUFX4_10/Y MUX2X1_249/S gnd DFFPOSX1_3/D vdd MUX2X1
XFILL_22_2_1 gnd vdd FILL
XCLKBUF1_37 CLKBUF1_2/A gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_26 CLKBUF1_5/A gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_15 CLKBUF1_8/A gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_59 clk gnd CLKBUF1_35/A vdd CLKBUF1
XCLKBUF1_48 CLKBUF1_14/A gnd CLKBUF1_48/Y vdd CLKBUF1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XAND2X2_1 INVX2_5/Y AND2X2_1/B gnd NOR2X1_2/B vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_17 NOR2X1_17/A AND2X2_2/Y gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 NOR2X1_28/A NOR2X1_22/B gnd NOR2X1_28/Y vdd NOR2X1
XMUX2X1_79 MUX2X1_79/A MUX2X1_79/B BUFX4_34/Y gnd MUX2X1_80/A vdd MUX2X1
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B gnd NOR2X1_39/Y vdd NOR2X1
XMUX2X1_46 INVX1_46/Y BUFX4_3/Y MUX2X1_46/S gnd MUX2X1_46/Y vdd MUX2X1
XMUX2X1_57 MUX2X1_57/A MUX2X1_57/B BUFX4_30/Y gnd MUX2X1_57/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_24 INVX1_24/Y BUFX4_41/Y MUX2X1_17/S gnd MUX2X1_24/Y vdd MUX2X1
XMUX2X1_68 MUX2X1_68/A MUX2X1_66/Y BUFX4_15/Y gnd AOI22X1_2/D vdd MUX2X1
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_35 INVX1_35/Y BUFX4_8/Y MUX2X1_39/S gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_13 INVX1_13/Y MUX2X1_5/B MUX2X1_9/S gnd MUX2X1_13/Y vdd MUX2X1
XFILL_2_1_1 gnd vdd FILL
XNAND2X1_83 MUX2X1_57/B NAND2X1_88/B gnd NAND2X1_83/Y vdd NAND2X1
XNAND2X1_72 MUX2X1_73/A NAND3X1_6/Y gnd OAI21X1_65/C vdd NAND2X1
XNAND2X1_94 NAND2X1_94/A NAND3X1_7/Y gnd OAI21X1_99/C vdd NAND2X1
XNAND2X1_61 MUX2X1_210/B NAND2X1_56/B gnd OAI21X1_55/C vdd NAND2X1
XNAND2X1_50 MUX2X1_163/B NAND3X1_5/Y gnd NAND2X1_50/Y vdd NAND2X1
XFILL_21_3 gnd vdd FILL
XFILL_14_2 gnd vdd FILL
XOAI21X1_48 BUFX4_43/Y NAND3X1_5/Y OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_59 BUFX4_7/Y NAND2X1_64/B OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_26 BUFX4_50/Y OAI21X1_25/B NAND2X1_31/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_15 BUFX4_22/Y OAI21X1_9/B OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_37 BUFX4_46/Y NAND3X1_4/Y OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XDFFPOSX1_198 MUX2X1_79/A CLKBUF1_29/Y OAI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_187 MUX2X1_229/B CLKBUF1_11/Y OAI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_132 MUX2X1_66/B CLKBUF1_40/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 NAND2X1_51/A CLKBUF1_18/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_110 MUX2X1_106/A CLKBUF1_5/A OAI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_143 MUX2X1_136/A CLKBUF1_2/A OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_154 MUX2X1_217/A CLKBUF1_14/Y OAI21X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_176 MUX2X1_153/B CLKBUF1_4/A OAI21X1_77/Y gnd vdd DFFPOSX1
XDFFPOSX1_165 INVX1_26/A CLKBUF1_34/Y MUX2X1_26/Y gnd vdd DFFPOSX1
XMUX2X1_241 MUX2X1_241/A MUX2X1_241/B BUFX4_32/Y gnd MUX2X1_242/A vdd MUX2X1
XMUX2X1_230 MUX2X1_229/Y MUX2X1_228/Y INVX2_6/A gnd MUX2X1_230/Y vdd MUX2X1
XMUX2X1_252 INVX1_62/Y BUFX4_24/Y MUX2X1_249/S gnd MUX2X1_252/Y vdd MUX2X1
XCLKBUF1_49 CLKBUF1_2/A gnd CLKBUF1_49/Y vdd CLKBUF1
XCLKBUF1_38 CLKBUF1_2/A gnd CLKBUF1_38/Y vdd CLKBUF1
XCLKBUF1_27 CLKBUF1_27/A gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_16 CLKBUF1_1/A gnd CLKBUF1_16/Y vdd CLKBUF1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XAND2X2_2 INVX2_5/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_29 NOR2X1_29/A NOR2X1_22/B gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_18 NOR2X1_18/A AND2X2_2/Y gnd NOR2X1_18/Y vdd NOR2X1
XNAND2X1_62 MUX2X1_234/B NAND2X1_56/B gnd OAI21X1_56/C vdd NAND2X1
XMUX2X1_58 MUX2X1_58/A MUX2X1_58/B BUFX4_31/Y gnd MUX2X1_59/A vdd MUX2X1
XMUX2X1_14 INVX1_14/Y BUFX4_2/Y MUX2X1_9/S gnd MUX2X1_14/Y vdd MUX2X1
XMUX2X1_69 INVX1_41/A INVX1_33/A BUFX4_38/Y gnd MUX2X1_71/B vdd MUX2X1
XMUX2X1_25 INVX1_25/Y MUX2X1_9/B MUX2X1_27/S gnd MUX2X1_25/Y vdd MUX2X1
XNAND2X1_51 NAND2X1_51/A NAND3X1_5/Y gnd OAI21X1_46/C vdd NAND2X1
XMUX2X1_36 INVX1_36/Y BUFX4_26/Y MUX2X1_39/S gnd MUX2X1_36/Y vdd MUX2X1
XNAND2X1_40 MUX2X1_106/A NAND3X1_4/Y gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_95 NAND2X1_95/A NAND3X1_7/Y gnd NAND2X1_95/Y vdd NAND2X1
XMUX2X1_47 INVX1_47/Y BUFX4_19/Y MUX2X1_46/S gnd MUX2X1_47/Y vdd MUX2X1
XNAND2X1_73 MUX2X1_97/A NAND3X1_6/Y gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_84 MUX2X1_81/B NAND2X1_88/B gnd OAI21X1_74/C vdd NAND2X1
XFILL_20_3_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XOAI21X1_16 BUFX4_40/Y OAI21X1_9/B NAND2X1_17/Y gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_38 BUFX4_5/Y NAND3X1_4/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_27 BUFX4_7/Y OAI21X1_25/B NAND2X1_32/Y gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_49 BUFX4_58/Y NAND2X1_56/B OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XDFFPOSX1_155 MUX2X1_241/A CLKBUF1_11/Y OAI21X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 MUX2X1_67/A CLKBUF1_40/Y OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 NAND2X1_41/A CLKBUF1_2/A OAI21X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_144 MUX2X1_160/A CLKBUF1_2/A OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 MUX2X1_90/B CLKBUF1_36/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 MUX2X1_211/B CLKBUF1_15/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_188 MUX2X1_60/A CLKBUF1_7/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_177 NAND2X1_88/A CLKBUF1_52/Y OAI21X1_78/Y gnd vdd DFFPOSX1
XDFFPOSX1_166 INVX1_27/A CLKBUF1_31/Y MUX2X1_27/Y gnd vdd DFFPOSX1
XMUX2X1_242 MUX2X1_242/A MUX2X1_240/Y BUFX4_17/Y gnd MUX2X1_242/Y vdd MUX2X1
XMUX2X1_231 INVX1_66/A INVX1_16/A BUFX4_36/Y gnd MUX2X1_231/Y vdd MUX2X1
XFILL_8_3_0 gnd vdd FILL
XMUX2X1_220 MUX2X1_220/A MUX2X1_220/B BUFX4_29/Y gnd MUX2X1_220/Y vdd MUX2X1
XFILL_0_2_0 gnd vdd FILL
XMUX2X1_253 INVX1_63/Y MUX2X1_5/B MUX2X1_249/S gnd DFFPOSX1_5/D vdd MUX2X1
XDFFPOSX1_199 MUX2X1_103/A CLKBUF1_28/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XCLKBUF1_17 CLKBUF1_7/A gnd CLKBUF1_17/Y vdd CLKBUF1
XFILL_16_2_0 gnd vdd FILL
XCLKBUF1_39 CLKBUF1_2/A gnd CLKBUF1_39/Y vdd CLKBUF1
XCLKBUF1_28 CLKBUF1_35/A gnd CLKBUF1_28/Y vdd CLKBUF1
XOR2X2_1 OR2X2_1/A INVX8_1/A gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_22_0_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 AND2X2_3/A INVX2_2/A gnd AND2X2_3/Y vdd AND2X2
XNOR2X1_19 NOR2X1_19/A AND2X2_2/Y gnd NOR2X1_19/Y vdd NOR2X1
XMUX2X1_48 INVX1_48/Y BUFX4_42/Y MUX2X1_46/S gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_59 MUX2X1_59/A MUX2X1_57/Y BUFX4_12/Y gnd AOI22X1_1/A vdd MUX2X1
XMUX2X1_15 INVX1_15/Y BUFX4_21/Y MUX2X1_9/S gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_26 INVX1_26/Y BUFX4_54/Y MUX2X1_27/S gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_37 INVX1_37/Y BUFX4_48/Y MUX2X1_39/S gnd MUX2X1_37/Y vdd MUX2X1
XNAND2X1_85 NAND2X1_85/A NAND2X1_88/B gnd OAI21X1_75/C vdd NAND2X1
XFILL_20_3_1 gnd vdd FILL
XNAND2X1_30 MUX2X1_67/A OAI21X1_25/B gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_74 NAND2X1_74/A NAND3X1_6/Y gnd OAI21X1_67/C vdd NAND2X1
XNAND2X1_63 INVX2_1/Y AND2X2_3/Y gnd NAND2X1_64/B vdd NAND2X1
XNAND2X1_41 NAND2X1_41/A NAND3X1_4/Y gnd OAI21X1_36/C vdd NAND2X1
XNAND2X1_96 NAND2X1_96/A NAND3X1_7/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_52 MUX2X1_211/B NAND3X1_5/Y gnd OAI21X1_47/C vdd NAND2X1
XFILL_11_3_1 gnd vdd FILL
XOAI21X1_17 MUX2X1_9/B NAND3X1_3/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 BUFX4_27/Y OAI21X1_25/B OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_39 MUX2X1_7/B NAND3X1_4/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XDFFPOSX1_123 MUX2X1_235/B CLKBUF1_12/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 INVX1_17/A CLKBUF1_7/Y MUX2X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 MUX2X1_114/B CLKBUF1_31/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 MUX2X1_184/A CLKBUF1_51/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_167 INVX1_28/A CLKBUF1_25/Y MUX2X1_28/Y gnd vdd DFFPOSX1
XFILL_0_2_1 gnd vdd FILL
XDFFPOSX1_101 MUX2X1_91/A CLKBUF1_36/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_189 MUX2X1_84/A CLKBUF1_1/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_178 NAND2X1_89/A CLKBUF1_46/Y OAI21X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 MUX2X1_154/A CLKBUF1_2/A OAI21X1_37/Y gnd vdd DFFPOSX1
XMUX2X1_243 NOR2X1_68/A MUX2X1_243/B BUFX4_33/Y gnd MUX2X1_245/B vdd MUX2X1
XMUX2X1_232 MUX2X1_232/A INVX1_32/A INVX2_3/A gnd MUX2X1_233/A vdd MUX2X1
XFILL_16_2_1 gnd vdd FILL
XMUX2X1_254 INVX1_64/Y BUFX4_1/Y MUX2X1_249/S gnd DFFPOSX1_6/D vdd MUX2X1
XFILL_8_3_1 gnd vdd FILL
XMUX2X1_221 MUX2X1_220/Y MUX2X1_221/B BUFX4_18/Y gnd AOI22X1_28/A vdd MUX2X1
XMUX2X1_210 NOR2X1_18/A MUX2X1_210/B BUFX4_33/Y gnd MUX2X1_210/Y vdd MUX2X1
XCLKBUF1_29 CLKBUF1_65/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XCLKBUF1_18 CLKBUF1_5/A gnd CLKBUF1_18/Y vdd CLKBUF1
XOR2X2_2 OR2X2_2/A INVX2_4/Y gnd OR2X2_2/Y vdd OR2X2
XBUFX4_50 INVX8_4/Y gnd BUFX4_50/Y vdd BUFX4
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XAND2X2_4 INVX2_5/Y AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XMUX2X1_38 INVX1_38/Y BUFX4_1/Y MUX2X1_39/S gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_27 INVX1_27/Y BUFX4_7/Y MUX2X1_27/S gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_49 INVX1_50/Y BUFX4_56/Y MUX2X1_56/S gnd MUX2X1_49/Y vdd MUX2X1
XMUX2X1_16 INVX1_16/Y BUFX4_44/Y MUX2X1_9/S gnd MUX2X1_16/Y vdd MUX2X1
XNAND2X1_20 MUX2X1_75/B NAND3X1_3/Y gnd OAI21X1_17/C vdd NAND2X1
XNAND2X1_64 MUX2X1_64/A NAND2X1_64/B gnd OAI21X1_57/C vdd NAND2X1
XNAND2X1_97 MUX2X1_199/A NAND3X1_7/Y gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_53 MUX2X1_235/B NAND3X1_5/Y gnd OAI21X1_48/C vdd NAND2X1
XNAND2X1_86 NAND2X1_86/A NAND2X1_88/B gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_75 MUX2X1_145/A NAND3X1_6/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_31 MUX2X1_91/A OAI21X1_25/B gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_42 MUX2X1_154/A NAND3X1_4/Y gnd OAI21X1_37/C vdd NAND2X1
XOAI21X1_18 BUFX4_52/Y NAND3X1_3/Y NAND2X1_21/Y gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 BUFX4_45/Y OAI21X1_25/B NAND2X1_34/Y gnd OAI21X1_29/Y vdd OAI21X1
XDFFPOSX1_113 MUX2X1_178/A CLKBUF1_52/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_179 NAND2X1_90/A CLKBUF1_44/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_102 NAND2X1_32/A CLKBUF1_32/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 MUX2X1_66/A CLKBUF1_6/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_135 NAND2X1_58/A CLKBUF1_26/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 INVX1_18/A CLKBUF1_1/Y MUX2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_146 NAND2X1_70/A CLKBUF1_45/Y OAI21X1_63/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 INVX1_29/A CLKBUF1_24/Y MUX2X1_29/Y gnd vdd DFFPOSX1
XMUX2X1_244 NAND2X1_17/A MUX2X1_244/B BUFX4_34/Y gnd MUX2X1_245/A vdd MUX2X1
XMUX2X1_200 MUX2X1_200/A MUX2X1_198/Y BUFX4_11/Y gnd AOI22X1_24/D vdd MUX2X1
XMUX2X1_233 MUX2X1_233/A MUX2X1_231/Y BUFX4_14/Y gnd MUX2X1_233/Y vdd MUX2X1
XMUX2X1_255 INVX1_65/Y BUFX4_21/Y MUX2X1_249/S gnd DFFPOSX1_7/D vdd MUX2X1
XMUX2X1_222 NOR2X1_8/A NAND2X1_7/A BUFX4_30/Y gnd MUX2X1_222/Y vdd MUX2X1
XMUX2X1_211 NAND2X1_36/A MUX2X1_211/B BUFX4_34/Y gnd MUX2X1_212/A vdd MUX2X1
XBUFX4_40 INVX8_10/Y gnd BUFX4_40/Y vdd BUFX4
XCLKBUF1_19 CLKBUF1_2/A gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_51 INVX8_4/Y gnd BUFX4_51/Y vdd BUFX4
XINVX8_10 datain[7] gnd INVX8_10/Y vdd INVX8
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends

