VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram32_sram
  CLASS BLOCK ;
  FOREIGN ram32_sram ;
  ORIGIN 2.600 3.000 ;
  SIZE 258.000 BY 246.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 240.200 252.600 240.800 ;
        RECT 0.600 235.900 1.000 240.200 ;
        RECT 4.600 236.500 5.000 240.200 ;
        RECT 6.200 235.900 6.600 240.200 ;
        RECT 8.300 237.900 8.700 240.200 ;
        RECT 9.400 237.900 9.800 240.200 ;
        RECT 11.000 237.900 11.400 240.200 ;
        RECT 12.600 235.900 13.000 240.200 ;
        RECT 15.400 237.900 15.800 240.200 ;
        RECT 17.000 237.900 17.400 240.200 ;
        RECT 19.800 236.000 20.200 240.200 ;
        RECT 21.400 235.900 21.800 240.200 ;
        RECT 23.000 236.500 23.400 240.200 ;
        RECT 24.600 235.900 25.000 240.200 ;
        RECT 26.200 235.900 26.600 240.200 ;
        RECT 27.800 235.900 28.200 240.200 ;
        RECT 28.600 235.900 29.000 240.200 ;
        RECT 30.700 237.900 31.100 240.200 ;
        RECT 31.800 237.900 32.200 240.200 ;
        RECT 33.400 237.900 33.800 240.200 ;
        RECT 35.000 236.000 35.400 240.200 ;
        RECT 37.800 237.900 38.200 240.200 ;
        RECT 39.400 237.900 39.800 240.200 ;
        RECT 42.200 235.900 42.600 240.200 ;
        RECT 46.200 235.900 46.600 240.200 ;
        RECT 49.000 237.900 49.400 240.200 ;
        RECT 50.600 237.900 51.000 240.200 ;
        RECT 53.400 236.000 53.800 240.200 ;
        RECT 55.000 237.900 55.400 240.200 ;
        RECT 56.600 237.900 57.000 240.200 ;
        RECT 57.700 237.900 58.100 240.200 ;
        RECT 59.800 235.900 60.200 240.200 ;
        RECT 61.400 236.000 61.800 240.200 ;
        RECT 64.200 237.900 64.600 240.200 ;
        RECT 65.800 237.900 66.200 240.200 ;
        RECT 68.600 235.900 69.000 240.200 ;
        RECT 70.200 237.900 70.600 240.200 ;
        RECT 71.800 237.900 72.200 240.200 ;
        RECT 72.900 237.900 73.300 240.200 ;
        RECT 75.000 235.900 75.400 240.200 ;
        RECT 76.600 235.900 77.000 240.200 ;
        RECT 79.400 237.900 79.800 240.200 ;
        RECT 81.000 237.900 81.400 240.200 ;
        RECT 83.800 236.000 84.200 240.200 ;
        RECT 86.200 236.500 86.600 240.200 ;
        RECT 87.800 235.900 88.200 240.200 ;
        RECT 89.400 236.500 89.800 240.200 ;
        RECT 91.000 235.900 91.400 240.200 ;
        RECT 92.600 235.900 93.000 240.200 ;
        RECT 94.200 235.900 94.600 240.200 ;
        RECT 95.800 235.900 96.200 240.200 ;
        RECT 97.400 235.900 97.800 240.200 ;
        RECT 100.600 236.000 101.000 240.200 ;
        RECT 103.400 237.900 103.800 240.200 ;
        RECT 105.000 237.900 105.400 240.200 ;
        RECT 107.800 235.900 108.200 240.200 ;
        RECT 109.400 235.900 109.800 240.200 ;
        RECT 111.500 237.900 111.900 240.200 ;
        RECT 112.600 235.900 113.000 240.200 ;
        RECT 114.200 235.900 114.600 240.200 ;
        RECT 115.800 235.900 116.200 240.200 ;
        RECT 117.400 236.000 117.800 240.200 ;
        RECT 120.200 237.900 120.600 240.200 ;
        RECT 121.800 237.900 122.200 240.200 ;
        RECT 124.600 235.900 125.000 240.200 ;
        RECT 126.200 237.900 126.600 240.200 ;
        RECT 127.800 237.900 128.200 240.200 ;
        RECT 128.900 237.900 129.300 240.200 ;
        RECT 131.000 235.900 131.400 240.200 ;
        RECT 131.800 235.900 132.200 240.200 ;
        RECT 133.900 237.900 134.300 240.200 ;
        RECT 135.000 237.900 135.400 240.200 ;
        RECT 136.600 237.900 137.000 240.200 ;
        RECT 138.200 236.000 138.600 240.200 ;
        RECT 141.000 237.900 141.400 240.200 ;
        RECT 142.600 237.900 143.000 240.200 ;
        RECT 145.400 235.900 145.800 240.200 ;
        RECT 147.800 236.500 148.200 240.200 ;
        RECT 153.400 235.900 153.800 240.200 ;
        RECT 155.000 236.500 155.400 240.200 ;
        RECT 156.600 235.900 157.000 240.200 ;
        RECT 158.700 237.900 159.100 240.200 ;
        RECT 159.800 237.900 160.200 240.200 ;
        RECT 161.400 237.900 161.800 240.200 ;
        RECT 163.000 235.900 163.400 240.200 ;
        RECT 165.800 237.900 166.200 240.200 ;
        RECT 167.400 237.900 167.800 240.200 ;
        RECT 170.200 236.000 170.600 240.200 ;
        RECT 172.600 235.900 173.000 240.200 ;
        RECT 175.400 237.900 175.800 240.200 ;
        RECT 177.000 237.900 177.400 240.200 ;
        RECT 179.800 236.000 180.200 240.200 ;
        RECT 182.200 236.000 182.600 240.200 ;
        RECT 185.000 237.900 185.400 240.200 ;
        RECT 186.600 237.900 187.000 240.200 ;
        RECT 189.400 235.900 189.800 240.200 ;
        RECT 191.000 235.900 191.400 240.200 ;
        RECT 193.100 237.900 193.500 240.200 ;
        RECT 195.000 236.000 195.400 240.200 ;
        RECT 197.800 237.900 198.200 240.200 ;
        RECT 199.400 237.900 199.800 240.200 ;
        RECT 202.200 235.900 202.600 240.200 ;
        RECT 205.400 237.900 205.800 240.200 ;
        RECT 207.000 237.900 207.400 240.200 ;
        RECT 208.100 237.900 208.500 240.200 ;
        RECT 210.200 235.900 210.600 240.200 ;
        RECT 211.800 236.000 212.200 240.200 ;
        RECT 214.600 237.900 215.000 240.200 ;
        RECT 216.200 237.900 216.600 240.200 ;
        RECT 219.000 235.900 219.400 240.200 ;
        RECT 220.600 237.900 221.000 240.200 ;
        RECT 222.200 237.900 222.600 240.200 ;
        RECT 223.800 236.000 224.200 240.200 ;
        RECT 226.600 237.900 227.000 240.200 ;
        RECT 228.200 237.900 228.600 240.200 ;
        RECT 231.000 235.900 231.400 240.200 ;
        RECT 233.400 236.000 233.800 240.200 ;
        RECT 236.200 237.900 236.600 240.200 ;
        RECT 237.800 237.900 238.200 240.200 ;
        RECT 240.600 235.900 241.000 240.200 ;
        RECT 242.200 235.900 242.600 240.200 ;
        RECT 243.800 235.900 244.200 240.200 ;
        RECT 245.400 235.900 245.800 240.200 ;
        RECT 246.200 235.900 246.600 240.200 ;
        RECT 248.300 237.900 248.700 240.200 ;
        RECT 249.400 237.900 249.800 240.200 ;
        RECT 251.000 237.900 251.400 240.200 ;
        RECT 1.400 220.800 1.800 225.100 ;
        RECT 4.200 220.800 4.600 223.100 ;
        RECT 5.800 220.800 6.200 223.100 ;
        RECT 8.600 220.800 9.000 225.000 ;
        RECT 10.200 220.800 10.600 225.100 ;
        RECT 11.800 220.800 12.200 225.100 ;
        RECT 13.400 220.800 13.800 225.100 ;
        RECT 15.000 220.800 15.400 225.100 ;
        RECT 16.600 220.800 17.000 225.100 ;
        RECT 17.400 220.800 17.800 225.100 ;
        RECT 19.500 220.800 19.900 223.100 ;
        RECT 20.600 220.800 21.000 223.100 ;
        RECT 22.200 220.800 22.600 223.100 ;
        RECT 23.800 220.800 24.200 225.000 ;
        RECT 26.600 220.800 27.000 223.100 ;
        RECT 28.200 220.800 28.600 223.100 ;
        RECT 31.000 220.800 31.400 225.100 ;
        RECT 33.400 220.800 33.800 224.900 ;
        RECT 36.000 220.800 36.400 225.100 ;
        RECT 37.400 220.800 37.800 225.100 ;
        RECT 39.500 220.800 39.900 223.100 ;
        RECT 40.600 220.800 41.000 223.100 ;
        RECT 42.200 220.800 42.600 223.100 ;
        RECT 43.800 220.800 44.200 225.000 ;
        RECT 46.600 220.800 47.000 223.100 ;
        RECT 48.200 220.800 48.600 223.100 ;
        RECT 51.000 220.800 51.400 225.100 ;
        RECT 55.000 220.800 55.400 224.900 ;
        RECT 57.600 220.800 58.000 225.100 ;
        RECT 59.800 220.800 60.200 224.900 ;
        RECT 62.400 220.800 62.800 225.100 ;
        RECT 64.600 220.800 65.000 224.900 ;
        RECT 67.200 220.800 67.600 225.100 ;
        RECT 68.600 220.800 69.000 225.100 ;
        RECT 70.200 220.800 70.600 225.100 ;
        RECT 71.800 220.800 72.200 225.100 ;
        RECT 73.400 220.800 73.800 225.100 ;
        RECT 75.000 220.800 75.400 225.100 ;
        RECT 76.600 220.800 77.000 225.100 ;
        RECT 79.400 220.800 79.800 223.100 ;
        RECT 81.000 220.800 81.400 223.100 ;
        RECT 83.800 220.800 84.200 225.000 ;
        RECT 85.400 220.800 85.800 223.100 ;
        RECT 87.000 220.800 87.400 223.100 ;
        RECT 88.100 220.800 88.500 223.100 ;
        RECT 90.200 220.800 90.600 225.100 ;
        RECT 91.600 220.800 92.000 225.100 ;
        RECT 94.200 220.800 94.600 224.900 ;
        RECT 98.200 220.800 98.600 225.100 ;
        RECT 101.000 220.800 101.400 223.100 ;
        RECT 102.600 220.800 103.000 223.100 ;
        RECT 105.400 220.800 105.800 225.000 ;
        RECT 107.000 220.800 107.400 225.100 ;
        RECT 109.100 220.800 109.500 223.100 ;
        RECT 110.200 220.800 110.600 223.100 ;
        RECT 111.800 220.800 112.200 223.100 ;
        RECT 112.900 220.800 113.300 223.100 ;
        RECT 115.000 220.800 115.400 225.100 ;
        RECT 115.800 220.800 116.200 225.100 ;
        RECT 119.800 220.800 120.200 224.500 ;
        RECT 121.400 220.800 121.800 223.100 ;
        RECT 123.000 220.800 123.400 223.100 ;
        RECT 124.400 220.800 124.800 225.100 ;
        RECT 127.000 220.800 127.400 224.900 ;
        RECT 129.400 220.800 129.800 225.100 ;
        RECT 132.200 220.800 132.600 223.100 ;
        RECT 133.800 220.800 134.200 223.100 ;
        RECT 136.600 220.800 137.000 225.000 ;
        RECT 138.200 220.800 138.600 225.100 ;
        RECT 140.300 220.800 140.700 223.100 ;
        RECT 141.400 220.800 141.800 223.100 ;
        RECT 143.000 220.800 143.400 223.100 ;
        RECT 144.400 220.800 144.800 225.100 ;
        RECT 147.000 220.800 147.400 224.900 ;
        RECT 151.000 220.800 151.400 225.100 ;
        RECT 153.800 220.800 154.200 223.100 ;
        RECT 155.400 220.800 155.800 223.100 ;
        RECT 158.200 220.800 158.600 225.000 ;
        RECT 160.600 220.800 161.000 224.500 ;
        RECT 164.600 220.800 165.000 225.100 ;
        RECT 165.400 220.800 165.800 225.100 ;
        RECT 167.000 220.800 167.400 225.100 ;
        RECT 168.600 220.800 169.000 225.100 ;
        RECT 170.200 220.800 170.600 225.100 ;
        RECT 171.800 220.800 172.200 225.100 ;
        RECT 173.400 220.800 173.800 225.000 ;
        RECT 176.200 220.800 176.600 223.100 ;
        RECT 177.800 220.800 178.200 223.100 ;
        RECT 180.600 220.800 181.000 225.100 ;
        RECT 183.000 220.800 183.400 224.900 ;
        RECT 185.600 220.800 186.000 225.100 ;
        RECT 187.600 220.800 188.000 225.100 ;
        RECT 190.200 220.800 190.600 224.900 ;
        RECT 192.600 220.800 193.000 224.900 ;
        RECT 195.200 220.800 195.600 225.100 ;
        RECT 196.600 220.800 197.000 225.100 ;
        RECT 198.700 220.800 199.100 223.100 ;
        RECT 199.800 220.800 200.200 223.100 ;
        RECT 201.400 220.800 201.800 223.100 ;
        RECT 203.800 220.800 204.200 223.100 ;
        RECT 205.400 220.800 205.800 223.100 ;
        RECT 207.000 220.800 207.400 225.000 ;
        RECT 209.800 220.800 210.200 223.100 ;
        RECT 211.400 220.800 211.800 223.100 ;
        RECT 214.200 220.800 214.600 225.100 ;
        RECT 216.600 220.800 217.000 224.900 ;
        RECT 219.200 220.800 219.600 225.100 ;
        RECT 221.200 220.800 221.600 225.100 ;
        RECT 223.800 220.800 224.200 224.900 ;
        RECT 225.400 220.800 225.800 225.100 ;
        RECT 227.500 220.800 227.900 223.100 ;
        RECT 228.600 220.800 229.000 223.100 ;
        RECT 230.200 220.800 230.600 223.100 ;
        RECT 231.800 220.800 232.200 225.100 ;
        RECT 234.600 220.800 235.000 223.100 ;
        RECT 236.200 220.800 236.600 223.100 ;
        RECT 239.000 220.800 239.400 225.000 ;
        RECT 241.400 220.800 241.800 225.100 ;
        RECT 244.200 220.800 244.600 223.100 ;
        RECT 245.800 220.800 246.200 223.100 ;
        RECT 248.600 220.800 249.000 225.000 ;
        RECT 0.200 220.200 252.600 220.800 ;
        RECT 1.400 215.900 1.800 220.200 ;
        RECT 4.200 217.900 4.600 220.200 ;
        RECT 5.800 217.900 6.200 220.200 ;
        RECT 8.600 216.000 9.000 220.200 ;
        RECT 10.200 215.900 10.600 220.200 ;
        RECT 12.300 217.900 12.700 220.200 ;
        RECT 13.400 217.900 13.800 220.200 ;
        RECT 15.000 217.900 15.400 220.200 ;
        RECT 16.600 216.000 17.000 220.200 ;
        RECT 19.400 217.900 19.800 220.200 ;
        RECT 21.000 217.900 21.400 220.200 ;
        RECT 23.800 215.900 24.200 220.200 ;
        RECT 26.000 215.900 26.400 220.200 ;
        RECT 28.600 216.100 29.000 220.200 ;
        RECT 31.800 215.900 32.200 220.200 ;
        RECT 34.200 216.500 34.600 220.200 ;
        RECT 36.600 215.900 37.000 220.200 ;
        RECT 39.400 217.900 39.800 220.200 ;
        RECT 41.000 217.900 41.400 220.200 ;
        RECT 43.800 216.000 44.200 220.200 ;
        RECT 46.200 216.500 46.600 220.200 ;
        RECT 50.200 215.900 50.600 220.200 ;
        RECT 53.000 217.900 53.400 220.200 ;
        RECT 54.600 217.900 55.000 220.200 ;
        RECT 57.400 216.000 57.800 220.200 ;
        RECT 59.800 215.900 60.200 220.200 ;
        RECT 62.600 217.900 63.000 220.200 ;
        RECT 64.200 217.900 64.600 220.200 ;
        RECT 67.000 216.000 67.400 220.200 ;
        RECT 68.900 217.900 69.300 220.200 ;
        RECT 71.000 215.900 71.400 220.200 ;
        RECT 72.600 216.500 73.000 220.200 ;
        RECT 75.800 216.500 76.200 220.200 ;
        RECT 77.400 215.900 77.800 220.200 ;
        RECT 78.200 215.900 78.600 220.200 ;
        RECT 79.800 216.500 80.200 220.200 ;
        RECT 82.200 216.000 82.600 220.200 ;
        RECT 85.000 217.900 85.400 220.200 ;
        RECT 86.600 217.900 87.000 220.200 ;
        RECT 89.400 215.900 89.800 220.200 ;
        RECT 91.000 215.900 91.400 220.200 ;
        RECT 93.100 217.900 93.500 220.200 ;
        RECT 94.200 217.900 94.600 220.200 ;
        RECT 95.800 217.900 96.200 220.200 ;
        RECT 97.200 215.900 97.600 220.200 ;
        RECT 99.800 216.100 100.200 220.200 ;
        RECT 103.300 217.900 103.700 220.200 ;
        RECT 105.400 215.900 105.800 220.200 ;
        RECT 106.200 217.900 106.600 220.200 ;
        RECT 107.800 217.900 108.200 220.200 ;
        RECT 109.400 215.900 109.800 220.200 ;
        RECT 112.200 217.900 112.600 220.200 ;
        RECT 113.800 217.900 114.200 220.200 ;
        RECT 116.600 216.000 117.000 220.200 ;
        RECT 118.200 217.900 118.600 220.200 ;
        RECT 119.800 217.900 120.200 220.200 ;
        RECT 121.400 215.900 121.800 220.200 ;
        RECT 124.200 217.900 124.600 220.200 ;
        RECT 125.800 217.900 126.200 220.200 ;
        RECT 128.600 216.000 129.000 220.200 ;
        RECT 130.200 215.900 130.600 220.200 ;
        RECT 132.300 217.900 132.700 220.200 ;
        RECT 133.400 217.900 133.800 220.200 ;
        RECT 135.000 217.900 135.400 220.200 ;
        RECT 136.600 216.000 137.000 220.200 ;
        RECT 139.400 217.900 139.800 220.200 ;
        RECT 141.000 217.900 141.400 220.200 ;
        RECT 143.800 215.900 144.200 220.200 ;
        RECT 146.200 215.900 146.600 220.200 ;
        RECT 149.000 217.900 149.400 220.200 ;
        RECT 150.600 217.900 151.000 220.200 ;
        RECT 153.400 216.000 153.800 220.200 ;
        RECT 156.600 215.900 157.000 220.200 ;
        RECT 158.700 217.900 159.100 220.200 ;
        RECT 159.800 217.900 160.200 220.200 ;
        RECT 161.400 217.900 161.800 220.200 ;
        RECT 162.200 215.900 162.600 220.200 ;
        RECT 164.300 217.900 164.700 220.200 ;
        RECT 165.400 217.900 165.800 220.200 ;
        RECT 167.000 217.900 167.400 220.200 ;
        RECT 168.600 216.000 169.000 220.200 ;
        RECT 171.400 217.900 171.800 220.200 ;
        RECT 173.000 217.900 173.400 220.200 ;
        RECT 175.800 215.900 176.200 220.200 ;
        RECT 177.400 215.900 177.800 220.200 ;
        RECT 179.000 216.500 179.400 220.200 ;
        RECT 180.600 217.900 181.000 220.200 ;
        RECT 182.200 217.900 182.600 220.200 ;
        RECT 183.800 215.900 184.200 220.200 ;
        RECT 186.600 217.900 187.000 220.200 ;
        RECT 188.200 217.900 188.600 220.200 ;
        RECT 191.000 216.000 191.400 220.200 ;
        RECT 192.600 215.900 193.000 220.200 ;
        RECT 194.200 215.900 194.600 220.200 ;
        RECT 195.800 215.900 196.200 220.200 ;
        RECT 197.400 215.900 197.800 220.200 ;
        RECT 199.000 215.900 199.400 220.200 ;
        RECT 200.600 216.500 201.000 220.200 ;
        RECT 202.200 215.900 202.600 220.200 ;
        RECT 204.600 215.900 205.000 220.200 ;
        RECT 206.700 217.900 207.100 220.200 ;
        RECT 207.800 217.900 208.200 220.200 ;
        RECT 209.400 217.900 209.800 220.200 ;
        RECT 210.200 215.900 210.600 220.200 ;
        RECT 211.800 215.900 212.200 220.200 ;
        RECT 213.400 215.900 213.800 220.200 ;
        RECT 215.000 215.900 215.400 220.200 ;
        RECT 216.600 215.900 217.000 220.200 ;
        RECT 217.400 217.900 217.800 220.200 ;
        RECT 219.000 217.900 219.400 220.200 ;
        RECT 220.100 217.900 220.500 220.200 ;
        RECT 222.200 215.900 222.600 220.200 ;
        RECT 223.800 216.000 224.200 220.200 ;
        RECT 226.600 217.900 227.000 220.200 ;
        RECT 228.200 217.900 228.600 220.200 ;
        RECT 231.000 215.900 231.400 220.200 ;
        RECT 232.900 217.900 233.300 220.200 ;
        RECT 235.000 215.900 235.400 220.200 ;
        RECT 235.800 217.900 236.200 220.200 ;
        RECT 237.400 217.900 237.800 220.200 ;
        RECT 238.500 217.900 238.900 220.200 ;
        RECT 240.600 215.900 241.000 220.200 ;
        RECT 242.200 215.900 242.600 220.200 ;
        RECT 245.000 217.900 245.400 220.200 ;
        RECT 246.600 217.900 247.000 220.200 ;
        RECT 249.400 216.000 249.800 220.200 ;
        RECT 1.400 200.800 1.800 205.100 ;
        RECT 4.200 200.800 4.600 203.100 ;
        RECT 5.800 200.800 6.200 203.100 ;
        RECT 8.600 200.800 9.000 205.000 ;
        RECT 10.200 200.800 10.600 205.100 ;
        RECT 12.300 200.800 12.700 203.100 ;
        RECT 13.400 200.800 13.800 203.100 ;
        RECT 15.000 200.800 15.400 203.100 ;
        RECT 15.800 200.800 16.200 205.100 ;
        RECT 17.900 200.800 18.300 203.100 ;
        RECT 19.000 200.800 19.400 203.100 ;
        RECT 20.600 200.800 21.000 203.100 ;
        RECT 22.200 200.800 22.600 204.900 ;
        RECT 24.800 200.800 25.200 205.100 ;
        RECT 27.000 200.800 27.400 205.100 ;
        RECT 29.800 200.800 30.200 203.100 ;
        RECT 31.400 200.800 31.800 203.100 ;
        RECT 34.200 200.800 34.600 205.000 ;
        RECT 35.800 200.800 36.200 203.100 ;
        RECT 37.400 200.800 37.800 203.100 ;
        RECT 38.500 200.800 38.900 203.100 ;
        RECT 40.600 200.800 41.000 205.100 ;
        RECT 42.200 200.800 42.600 205.000 ;
        RECT 45.000 200.800 45.400 203.100 ;
        RECT 46.600 200.800 47.000 203.100 ;
        RECT 49.400 200.800 49.800 205.100 ;
        RECT 52.600 200.800 53.000 203.100 ;
        RECT 54.200 200.800 54.600 203.100 ;
        RECT 55.800 200.800 56.200 204.500 ;
        RECT 58.800 200.800 59.200 205.100 ;
        RECT 61.400 200.800 61.800 204.900 ;
        RECT 63.000 200.800 63.400 203.100 ;
        RECT 64.600 200.800 65.000 203.100 ;
        RECT 66.200 200.800 66.600 205.100 ;
        RECT 69.000 200.800 69.400 203.100 ;
        RECT 70.600 200.800 71.000 203.100 ;
        RECT 73.400 200.800 73.800 205.000 ;
        RECT 75.000 200.800 75.400 205.100 ;
        RECT 77.400 200.800 77.800 203.100 ;
        RECT 79.000 200.800 79.400 203.100 ;
        RECT 80.600 200.800 81.000 205.000 ;
        RECT 83.400 200.800 83.800 203.100 ;
        RECT 85.000 200.800 85.400 203.100 ;
        RECT 87.800 200.800 88.200 205.100 ;
        RECT 90.200 200.800 90.600 204.900 ;
        RECT 92.800 200.800 93.200 205.100 ;
        RECT 94.800 200.800 95.200 205.100 ;
        RECT 97.400 200.800 97.800 204.900 ;
        RECT 100.600 200.800 101.000 203.100 ;
        RECT 102.200 200.800 102.600 203.100 ;
        RECT 103.800 200.800 104.200 205.100 ;
        RECT 106.600 200.800 107.000 203.100 ;
        RECT 108.200 200.800 108.600 203.100 ;
        RECT 111.000 200.800 111.400 205.000 ;
        RECT 113.400 200.800 113.800 204.900 ;
        RECT 116.000 200.800 116.400 205.100 ;
        RECT 118.200 200.800 118.600 204.500 ;
        RECT 119.800 200.800 120.200 205.100 ;
        RECT 121.400 200.800 121.800 204.500 ;
        RECT 124.600 200.800 125.000 204.900 ;
        RECT 127.200 200.800 127.600 205.100 ;
        RECT 129.400 200.800 129.800 205.100 ;
        RECT 132.200 200.800 132.600 203.100 ;
        RECT 133.800 200.800 134.200 203.100 ;
        RECT 136.600 200.800 137.000 205.000 ;
        RECT 138.200 200.800 138.600 205.100 ;
        RECT 142.200 200.800 142.600 204.500 ;
        RECT 145.400 200.800 145.800 205.100 ;
        RECT 147.800 200.800 148.200 204.500 ;
        RECT 151.800 200.800 152.200 205.000 ;
        RECT 154.600 200.800 155.000 203.100 ;
        RECT 156.200 200.800 156.600 203.100 ;
        RECT 159.000 200.800 159.400 205.100 ;
        RECT 161.400 200.800 161.800 204.900 ;
        RECT 164.000 200.800 164.400 205.100 ;
        RECT 165.400 200.800 165.800 205.100 ;
        RECT 167.500 200.800 167.900 203.100 ;
        RECT 168.600 200.800 169.000 203.100 ;
        RECT 170.200 200.800 170.600 203.100 ;
        RECT 171.800 200.800 172.200 205.000 ;
        RECT 174.600 200.800 175.000 203.100 ;
        RECT 176.200 200.800 176.600 203.100 ;
        RECT 179.000 200.800 179.400 205.100 ;
        RECT 182.200 200.800 182.600 204.500 ;
        RECT 184.400 200.800 184.800 205.100 ;
        RECT 187.000 200.800 187.400 204.900 ;
        RECT 189.200 200.800 189.600 205.100 ;
        RECT 191.800 200.800 192.200 204.900 ;
        RECT 195.000 200.800 195.400 205.100 ;
        RECT 197.400 200.800 197.800 204.500 ;
        RECT 199.000 200.800 199.400 205.100 ;
        RECT 201.100 200.800 201.500 203.100 ;
        RECT 204.600 200.800 205.000 205.100 ;
        RECT 207.400 200.800 207.800 203.100 ;
        RECT 209.000 200.800 209.400 203.100 ;
        RECT 211.800 200.800 212.200 205.000 ;
        RECT 213.400 200.800 213.800 205.100 ;
        RECT 215.000 200.800 215.400 205.100 ;
        RECT 216.600 200.800 217.000 205.100 ;
        RECT 218.200 200.800 218.600 205.100 ;
        RECT 219.800 200.800 220.200 205.100 ;
        RECT 221.200 200.800 221.600 205.100 ;
        RECT 223.800 200.800 224.200 204.900 ;
        RECT 226.200 200.800 226.600 204.900 ;
        RECT 228.800 200.800 229.200 205.100 ;
        RECT 230.200 200.800 230.600 203.100 ;
        RECT 231.800 200.800 232.200 203.100 ;
        RECT 233.400 200.800 233.800 205.100 ;
        RECT 236.200 200.800 236.600 203.100 ;
        RECT 237.800 200.800 238.200 203.100 ;
        RECT 240.600 200.800 241.000 205.000 ;
        RECT 242.200 200.800 242.600 203.100 ;
        RECT 243.800 200.800 244.200 203.100 ;
        RECT 244.600 200.800 245.000 205.100 ;
        RECT 247.800 200.800 248.200 204.500 ;
        RECT 0.200 200.200 252.600 200.800 ;
        RECT 1.400 195.900 1.800 200.200 ;
        RECT 4.200 197.900 4.600 200.200 ;
        RECT 5.800 197.900 6.200 200.200 ;
        RECT 8.600 196.000 9.000 200.200 ;
        RECT 11.000 196.000 11.400 200.200 ;
        RECT 13.800 197.900 14.200 200.200 ;
        RECT 15.400 197.900 15.800 200.200 ;
        RECT 18.200 195.900 18.600 200.200 ;
        RECT 19.800 195.900 20.200 200.200 ;
        RECT 21.400 195.900 21.800 200.200 ;
        RECT 23.000 195.900 23.400 200.200 ;
        RECT 24.600 195.900 25.000 200.200 ;
        RECT 26.200 195.900 26.600 200.200 ;
        RECT 27.000 197.900 27.400 200.200 ;
        RECT 28.600 197.900 29.000 200.200 ;
        RECT 29.700 197.900 30.100 200.200 ;
        RECT 31.800 195.900 32.200 200.200 ;
        RECT 33.400 196.000 33.800 200.200 ;
        RECT 36.200 197.900 36.600 200.200 ;
        RECT 37.800 197.900 38.200 200.200 ;
        RECT 40.600 195.900 41.000 200.200 ;
        RECT 42.200 195.900 42.600 200.200 ;
        RECT 43.800 196.500 44.200 200.200 ;
        RECT 46.200 196.100 46.600 200.200 ;
        RECT 48.800 195.900 49.200 200.200 ;
        RECT 52.600 196.100 53.000 200.200 ;
        RECT 55.200 195.900 55.600 200.200 ;
        RECT 56.600 197.900 57.000 200.200 ;
        RECT 58.200 197.900 58.600 200.200 ;
        RECT 59.300 197.900 59.700 200.200 ;
        RECT 61.400 195.900 61.800 200.200 ;
        RECT 62.200 195.900 62.600 200.200 ;
        RECT 64.300 197.900 64.700 200.200 ;
        RECT 66.200 196.500 66.600 200.200 ;
        RECT 69.400 197.900 69.800 200.200 ;
        RECT 71.000 197.900 71.400 200.200 ;
        RECT 71.800 195.900 72.200 200.200 ;
        RECT 73.400 196.500 73.800 200.200 ;
        RECT 75.800 196.500 76.200 200.200 ;
        RECT 77.400 195.900 77.800 200.200 ;
        RECT 78.500 197.900 78.900 200.200 ;
        RECT 80.600 195.900 81.000 200.200 ;
        RECT 82.200 195.900 82.600 200.200 ;
        RECT 85.000 197.900 85.400 200.200 ;
        RECT 86.600 197.900 87.000 200.200 ;
        RECT 89.400 196.000 89.800 200.200 ;
        RECT 91.600 195.900 92.000 200.200 ;
        RECT 94.200 196.100 94.600 200.200 ;
        RECT 95.800 195.900 96.200 200.200 ;
        RECT 97.900 197.900 98.300 200.200 ;
        RECT 100.600 197.900 101.000 200.200 ;
        RECT 102.200 197.900 102.600 200.200 ;
        RECT 103.800 195.900 104.200 200.200 ;
        RECT 106.600 197.900 107.000 200.200 ;
        RECT 108.200 197.900 108.600 200.200 ;
        RECT 111.000 196.000 111.400 200.200 ;
        RECT 113.200 195.900 113.600 200.200 ;
        RECT 115.800 196.100 116.200 200.200 ;
        RECT 118.200 195.900 118.600 200.200 ;
        RECT 121.000 197.900 121.400 200.200 ;
        RECT 122.600 197.900 123.000 200.200 ;
        RECT 125.400 196.000 125.800 200.200 ;
        RECT 127.600 195.900 128.000 200.200 ;
        RECT 130.200 196.100 130.600 200.200 ;
        RECT 132.400 195.900 132.800 200.200 ;
        RECT 135.000 196.100 135.400 200.200 ;
        RECT 137.400 196.500 137.800 200.200 ;
        RECT 141.200 195.900 141.600 200.200 ;
        RECT 143.800 196.100 144.200 200.200 ;
        RECT 145.400 195.900 145.800 200.200 ;
        RECT 147.500 197.900 147.900 200.200 ;
        RECT 151.000 196.000 151.400 200.200 ;
        RECT 153.800 197.900 154.200 200.200 ;
        RECT 155.400 197.900 155.800 200.200 ;
        RECT 158.200 195.900 158.600 200.200 ;
        RECT 160.600 195.900 161.000 200.200 ;
        RECT 163.400 197.900 163.800 200.200 ;
        RECT 165.000 197.900 165.400 200.200 ;
        RECT 167.800 196.000 168.200 200.200 ;
        RECT 169.400 197.900 169.800 200.200 ;
        RECT 171.000 197.900 171.400 200.200 ;
        RECT 172.100 197.900 172.500 200.200 ;
        RECT 174.200 195.900 174.600 200.200 ;
        RECT 175.000 195.900 175.400 200.200 ;
        RECT 176.600 195.900 177.000 200.200 ;
        RECT 178.200 195.900 178.600 200.200 ;
        RECT 179.800 195.900 180.200 200.200 ;
        RECT 181.400 195.900 181.800 200.200 ;
        RECT 182.500 197.900 182.900 200.200 ;
        RECT 184.600 195.900 185.000 200.200 ;
        RECT 185.400 197.900 185.800 200.200 ;
        RECT 187.000 197.900 187.400 200.200 ;
        RECT 190.200 196.500 190.600 200.200 ;
        RECT 192.600 196.100 193.000 200.200 ;
        RECT 195.200 195.900 195.600 200.200 ;
        RECT 197.200 195.900 197.600 200.200 ;
        RECT 199.800 196.100 200.200 200.200 ;
        RECT 203.800 195.900 204.200 200.200 ;
        RECT 206.600 197.900 207.000 200.200 ;
        RECT 208.200 197.900 208.600 200.200 ;
        RECT 211.000 196.000 211.400 200.200 ;
        RECT 212.600 195.900 213.000 200.200 ;
        RECT 214.700 197.900 215.100 200.200 ;
        RECT 215.800 195.900 216.200 200.200 ;
        RECT 217.900 197.900 218.300 200.200 ;
        RECT 219.000 197.900 219.400 200.200 ;
        RECT 220.600 197.900 221.000 200.200 ;
        RECT 222.200 195.900 222.600 200.200 ;
        RECT 225.000 197.900 225.400 200.200 ;
        RECT 226.600 197.900 227.000 200.200 ;
        RECT 229.400 196.000 229.800 200.200 ;
        RECT 231.000 195.900 231.400 200.200 ;
        RECT 233.100 197.900 233.500 200.200 ;
        RECT 235.000 195.900 235.400 200.200 ;
        RECT 237.800 197.900 238.200 200.200 ;
        RECT 239.400 197.900 239.800 200.200 ;
        RECT 242.200 196.000 242.600 200.200 ;
        RECT 244.100 197.900 244.500 200.200 ;
        RECT 246.200 195.900 246.600 200.200 ;
        RECT 247.800 196.500 248.200 200.200 ;
        RECT 249.400 195.900 249.800 200.200 ;
        RECT 0.600 180.800 1.000 183.100 ;
        RECT 2.200 180.800 2.600 183.100 ;
        RECT 3.300 180.800 3.700 183.100 ;
        RECT 5.400 180.800 5.800 185.100 ;
        RECT 6.200 180.800 6.600 185.100 ;
        RECT 8.300 180.800 8.700 183.100 ;
        RECT 9.400 180.800 9.800 183.100 ;
        RECT 11.000 180.800 11.400 183.100 ;
        RECT 12.400 180.800 12.800 185.100 ;
        RECT 15.000 180.800 15.400 184.900 ;
        RECT 16.600 180.800 17.000 185.100 ;
        RECT 18.200 180.800 18.600 185.100 ;
        RECT 19.800 180.800 20.200 185.100 ;
        RECT 21.400 180.800 21.800 185.100 ;
        RECT 23.000 180.800 23.400 185.100 ;
        RECT 24.400 180.800 24.800 185.100 ;
        RECT 27.000 180.800 27.400 184.900 ;
        RECT 29.200 180.800 29.600 185.100 ;
        RECT 31.800 180.800 32.200 184.900 ;
        RECT 33.400 180.800 33.800 185.100 ;
        RECT 35.000 180.800 35.400 185.100 ;
        RECT 36.600 180.800 37.000 185.100 ;
        RECT 38.200 180.800 38.600 185.100 ;
        RECT 39.800 180.800 40.200 185.100 ;
        RECT 40.600 180.800 41.000 185.100 ;
        RECT 44.600 180.800 45.000 184.500 ;
        RECT 48.600 180.800 49.000 185.100 ;
        RECT 51.400 180.800 51.800 183.100 ;
        RECT 53.000 180.800 53.400 183.100 ;
        RECT 55.800 180.800 56.200 185.000 ;
        RECT 58.200 180.800 58.600 184.900 ;
        RECT 60.800 180.800 61.200 185.100 ;
        RECT 62.800 180.800 63.200 185.100 ;
        RECT 65.400 180.800 65.800 184.900 ;
        RECT 67.800 180.800 68.200 184.900 ;
        RECT 70.400 180.800 70.800 185.100 ;
        RECT 74.200 180.800 74.600 184.500 ;
        RECT 76.600 180.800 77.000 185.000 ;
        RECT 79.400 180.800 79.800 183.100 ;
        RECT 81.000 180.800 81.400 183.100 ;
        RECT 83.800 180.800 84.200 185.100 ;
        RECT 85.400 180.800 85.800 183.100 ;
        RECT 87.000 180.800 87.400 183.100 ;
        RECT 88.100 180.800 88.500 183.100 ;
        RECT 90.200 180.800 90.600 185.100 ;
        RECT 91.000 180.800 91.400 183.100 ;
        RECT 92.600 180.800 93.000 183.100 ;
        RECT 93.700 180.800 94.100 183.100 ;
        RECT 95.800 180.800 96.200 185.100 ;
        RECT 97.200 180.800 97.600 185.100 ;
        RECT 99.800 180.800 100.200 184.900 ;
        RECT 103.800 180.800 104.200 185.000 ;
        RECT 106.600 180.800 107.000 183.100 ;
        RECT 108.200 180.800 108.600 183.100 ;
        RECT 111.000 180.800 111.400 185.100 ;
        RECT 112.600 180.800 113.000 183.100 ;
        RECT 114.200 180.800 114.600 183.100 ;
        RECT 115.300 180.800 115.700 183.100 ;
        RECT 117.400 180.800 117.800 185.100 ;
        RECT 118.200 180.800 118.600 185.100 ;
        RECT 120.300 180.800 120.700 183.100 ;
        RECT 122.200 180.800 122.600 185.100 ;
        RECT 125.000 180.800 125.400 183.100 ;
        RECT 126.600 180.800 127.000 183.100 ;
        RECT 129.400 180.800 129.800 185.000 ;
        RECT 131.000 180.800 131.400 185.100 ;
        RECT 133.100 180.800 133.500 183.100 ;
        RECT 134.200 180.800 134.600 185.100 ;
        RECT 135.800 180.800 136.200 185.100 ;
        RECT 137.400 180.800 137.800 185.100 ;
        RECT 139.000 180.800 139.400 185.100 ;
        RECT 140.600 180.800 141.000 185.100 ;
        RECT 141.400 180.800 141.800 185.100 ;
        RECT 145.400 180.800 145.800 184.500 ;
        RECT 147.000 180.800 147.400 183.100 ;
        RECT 148.600 180.800 149.000 183.100 ;
        RECT 151.800 180.800 152.200 184.500 ;
        RECT 155.800 180.800 156.200 184.500 ;
        RECT 157.400 180.800 157.800 185.100 ;
        RECT 158.200 180.800 158.600 183.100 ;
        RECT 159.800 180.800 160.200 183.100 ;
        RECT 160.600 180.800 161.000 183.100 ;
        RECT 162.200 180.800 162.600 183.100 ;
        RECT 163.000 180.800 163.400 185.100 ;
        RECT 165.100 180.800 165.500 183.100 ;
        RECT 167.000 180.800 167.400 185.100 ;
        RECT 169.800 180.800 170.200 183.100 ;
        RECT 171.400 180.800 171.800 183.100 ;
        RECT 174.200 180.800 174.600 185.000 ;
        RECT 176.600 180.800 177.000 184.900 ;
        RECT 179.200 180.800 179.600 185.100 ;
        RECT 180.600 180.800 181.000 185.100 ;
        RECT 182.700 180.800 183.100 183.100 ;
        RECT 183.800 180.800 184.200 183.100 ;
        RECT 185.400 180.800 185.800 183.100 ;
        RECT 188.600 180.800 189.000 184.500 ;
        RECT 191.000 180.800 191.400 185.100 ;
        RECT 193.800 180.800 194.200 183.100 ;
        RECT 195.400 180.800 195.800 183.100 ;
        RECT 198.200 180.800 198.600 185.000 ;
        RECT 199.800 180.800 200.200 183.100 ;
        RECT 201.400 180.800 201.800 183.100 ;
        RECT 204.600 180.800 205.000 185.100 ;
        RECT 207.400 180.800 207.800 183.100 ;
        RECT 209.000 180.800 209.400 183.100 ;
        RECT 211.800 180.800 212.200 185.000 ;
        RECT 213.400 180.800 213.800 183.100 ;
        RECT 215.000 180.800 215.400 183.100 ;
        RECT 216.600 180.800 217.000 184.900 ;
        RECT 219.200 180.800 219.600 185.100 ;
        RECT 221.200 180.800 221.600 185.100 ;
        RECT 223.800 180.800 224.200 184.900 ;
        RECT 225.400 180.800 225.800 185.100 ;
        RECT 227.500 180.800 227.900 183.100 ;
        RECT 228.600 180.800 229.000 183.100 ;
        RECT 230.200 180.800 230.600 183.100 ;
        RECT 231.800 180.800 232.200 185.000 ;
        RECT 234.600 180.800 235.000 183.100 ;
        RECT 236.200 180.800 236.600 183.100 ;
        RECT 239.000 180.800 239.400 185.100 ;
        RECT 240.600 180.800 241.000 185.100 ;
        RECT 242.200 180.800 242.600 185.100 ;
        RECT 243.800 180.800 244.200 185.100 ;
        RECT 245.400 180.800 245.800 185.100 ;
        RECT 247.000 180.800 247.400 185.100 ;
        RECT 247.800 180.800 248.200 185.100 ;
        RECT 249.400 180.800 249.800 184.500 ;
        RECT 0.200 180.200 252.600 180.800 ;
        RECT 1.400 175.900 1.800 180.200 ;
        RECT 4.200 177.900 4.600 180.200 ;
        RECT 5.800 177.900 6.200 180.200 ;
        RECT 8.600 176.000 9.000 180.200 ;
        RECT 10.500 177.900 10.900 180.200 ;
        RECT 12.600 175.900 13.000 180.200 ;
        RECT 13.400 177.900 13.800 180.200 ;
        RECT 15.000 177.900 15.400 180.200 ;
        RECT 15.800 177.900 16.200 180.200 ;
        RECT 17.400 177.900 17.800 180.200 ;
        RECT 18.200 175.900 18.600 180.200 ;
        RECT 20.300 177.900 20.700 180.200 ;
        RECT 21.400 177.900 21.800 180.200 ;
        RECT 23.000 177.900 23.400 180.200 ;
        RECT 24.600 176.000 25.000 180.200 ;
        RECT 27.400 177.900 27.800 180.200 ;
        RECT 29.000 177.900 29.400 180.200 ;
        RECT 31.800 175.900 32.200 180.200 ;
        RECT 34.200 175.900 34.600 180.200 ;
        RECT 37.000 177.900 37.400 180.200 ;
        RECT 38.600 177.900 39.000 180.200 ;
        RECT 41.400 176.000 41.800 180.200 ;
        RECT 43.300 177.900 43.700 180.200 ;
        RECT 45.400 175.900 45.800 180.200 ;
        RECT 48.600 176.100 49.000 180.200 ;
        RECT 51.200 175.900 51.600 180.200 ;
        RECT 52.600 177.900 53.000 180.200 ;
        RECT 54.200 177.900 54.600 180.200 ;
        RECT 55.800 176.500 56.200 180.200 ;
        RECT 59.000 177.900 59.400 180.200 ;
        RECT 60.600 177.900 61.000 180.200 ;
        RECT 61.700 177.900 62.100 180.200 ;
        RECT 63.800 175.900 64.200 180.200 ;
        RECT 65.400 175.900 65.800 180.200 ;
        RECT 68.200 177.900 68.600 180.200 ;
        RECT 69.800 177.900 70.200 180.200 ;
        RECT 72.600 176.000 73.000 180.200 ;
        RECT 74.800 175.900 75.200 180.200 ;
        RECT 77.400 176.100 77.800 180.200 ;
        RECT 79.800 176.000 80.200 180.200 ;
        RECT 82.600 177.900 83.000 180.200 ;
        RECT 84.200 177.900 84.600 180.200 ;
        RECT 87.000 175.900 87.400 180.200 ;
        RECT 89.200 175.900 89.600 180.200 ;
        RECT 91.800 176.100 92.200 180.200 ;
        RECT 94.000 175.900 94.400 180.200 ;
        RECT 96.600 176.100 97.000 180.200 ;
        RECT 100.400 175.900 100.800 180.200 ;
        RECT 103.000 176.100 103.400 180.200 ;
        RECT 105.400 175.900 105.800 180.200 ;
        RECT 108.200 177.900 108.600 180.200 ;
        RECT 109.800 177.900 110.200 180.200 ;
        RECT 112.600 176.000 113.000 180.200 ;
        RECT 114.200 177.900 114.600 180.200 ;
        RECT 115.800 177.900 116.200 180.200 ;
        RECT 116.900 177.900 117.300 180.200 ;
        RECT 119.000 175.900 119.400 180.200 ;
        RECT 119.800 177.900 120.200 180.200 ;
        RECT 121.400 177.900 121.800 180.200 ;
        RECT 122.200 175.900 122.600 180.200 ;
        RECT 123.800 176.500 124.200 180.200 ;
        RECT 126.000 175.900 126.400 180.200 ;
        RECT 128.600 176.100 129.000 180.200 ;
        RECT 131.000 176.500 131.400 180.200 ;
        RECT 134.800 175.900 135.200 180.200 ;
        RECT 137.400 176.100 137.800 180.200 ;
        RECT 139.600 175.900 140.000 180.200 ;
        RECT 142.200 176.100 142.600 180.200 ;
        RECT 144.400 175.900 144.800 180.200 ;
        RECT 147.000 176.100 147.400 180.200 ;
        RECT 148.600 177.900 149.000 180.200 ;
        RECT 150.200 177.900 150.600 180.200 ;
        RECT 152.900 177.900 153.300 180.200 ;
        RECT 155.000 175.900 155.400 180.200 ;
        RECT 156.600 175.900 157.000 180.200 ;
        RECT 159.400 177.900 159.800 180.200 ;
        RECT 161.000 177.900 161.400 180.200 ;
        RECT 163.800 176.000 164.200 180.200 ;
        RECT 166.000 175.900 166.400 180.200 ;
        RECT 168.600 176.100 169.000 180.200 ;
        RECT 170.200 177.900 170.600 180.200 ;
        RECT 171.800 177.900 172.200 180.200 ;
        RECT 172.900 177.900 173.300 180.200 ;
        RECT 175.000 175.900 175.400 180.200 ;
        RECT 176.600 175.900 177.000 180.200 ;
        RECT 179.400 177.900 179.800 180.200 ;
        RECT 181.000 177.900 181.400 180.200 ;
        RECT 183.800 176.000 184.200 180.200 ;
        RECT 186.200 176.500 186.600 180.200 ;
        RECT 187.800 175.900 188.200 180.200 ;
        RECT 189.400 176.000 189.800 180.200 ;
        RECT 192.200 177.900 192.600 180.200 ;
        RECT 193.800 177.900 194.200 180.200 ;
        RECT 196.600 175.900 197.000 180.200 ;
        RECT 199.000 176.100 199.400 180.200 ;
        RECT 201.600 175.900 202.000 180.200 ;
        RECT 207.000 176.500 207.400 180.200 ;
        RECT 208.600 175.900 209.000 180.200 ;
        RECT 210.700 177.900 211.100 180.200 ;
        RECT 212.600 175.900 213.000 180.200 ;
        RECT 215.400 177.900 215.800 180.200 ;
        RECT 217.000 177.900 217.400 180.200 ;
        RECT 219.800 176.000 220.200 180.200 ;
        RECT 222.000 175.900 222.400 180.200 ;
        RECT 224.600 176.100 225.000 180.200 ;
        RECT 227.000 176.100 227.400 180.200 ;
        RECT 229.600 175.900 230.000 180.200 ;
        RECT 231.600 175.900 232.000 180.200 ;
        RECT 234.200 176.100 234.600 180.200 ;
        RECT 235.800 177.900 236.200 180.200 ;
        RECT 237.400 177.900 237.800 180.200 ;
        RECT 239.000 175.900 239.400 180.200 ;
        RECT 241.800 177.900 242.200 180.200 ;
        RECT 243.400 177.900 243.800 180.200 ;
        RECT 246.200 176.000 246.600 180.200 ;
        RECT 247.800 175.900 248.200 180.200 ;
        RECT 249.900 177.900 250.300 180.200 ;
        RECT 0.600 160.800 1.000 165.100 ;
        RECT 2.200 160.800 2.600 165.100 ;
        RECT 3.800 160.800 4.200 165.100 ;
        RECT 5.400 160.800 5.800 165.100 ;
        RECT 7.000 160.800 7.400 165.100 ;
        RECT 8.600 160.800 9.000 165.000 ;
        RECT 11.400 160.800 11.800 163.100 ;
        RECT 13.000 160.800 13.400 163.100 ;
        RECT 15.800 160.800 16.200 165.100 ;
        RECT 17.700 160.800 18.100 163.100 ;
        RECT 19.800 160.800 20.200 165.100 ;
        RECT 21.400 160.800 21.800 165.000 ;
        RECT 24.200 160.800 24.600 163.100 ;
        RECT 25.800 160.800 26.200 163.100 ;
        RECT 28.600 160.800 29.000 165.100 ;
        RECT 30.200 160.800 30.600 163.100 ;
        RECT 31.800 160.800 32.200 163.100 ;
        RECT 32.900 160.800 33.300 163.100 ;
        RECT 35.000 160.800 35.400 165.100 ;
        RECT 36.400 160.800 36.800 165.100 ;
        RECT 39.000 160.800 39.400 164.900 ;
        RECT 40.600 160.800 41.000 163.100 ;
        RECT 42.200 160.800 42.600 163.100 ;
        RECT 43.600 160.800 44.000 165.100 ;
        RECT 46.200 160.800 46.600 164.900 ;
        RECT 51.800 160.800 52.200 164.500 ;
        RECT 54.200 160.800 54.600 165.000 ;
        RECT 57.000 160.800 57.400 163.100 ;
        RECT 58.600 160.800 59.000 163.100 ;
        RECT 61.400 160.800 61.800 165.100 ;
        RECT 63.000 160.800 63.400 165.100 ;
        RECT 65.100 160.800 65.500 163.100 ;
        RECT 66.200 160.800 66.600 163.100 ;
        RECT 67.800 160.800 68.200 163.100 ;
        RECT 69.400 160.800 69.800 164.900 ;
        RECT 72.000 160.800 72.400 165.100 ;
        RECT 74.000 160.800 74.400 165.100 ;
        RECT 76.600 160.800 77.000 164.900 ;
        RECT 78.200 160.800 78.600 165.100 ;
        RECT 80.300 160.800 80.700 163.100 ;
        RECT 81.400 160.800 81.800 163.100 ;
        RECT 83.000 160.800 83.400 163.100 ;
        RECT 86.200 160.800 86.600 164.500 ;
        RECT 88.600 160.800 89.000 165.100 ;
        RECT 91.400 160.800 91.800 163.100 ;
        RECT 93.000 160.800 93.400 163.100 ;
        RECT 95.800 160.800 96.200 165.000 ;
        RECT 97.400 160.800 97.800 163.100 ;
        RECT 99.000 160.800 99.400 163.100 ;
        RECT 101.700 160.800 102.100 163.100 ;
        RECT 103.800 160.800 104.200 165.100 ;
        RECT 105.400 160.800 105.800 165.000 ;
        RECT 108.200 160.800 108.600 163.100 ;
        RECT 109.800 160.800 110.200 163.100 ;
        RECT 112.600 160.800 113.000 165.100 ;
        RECT 114.200 160.800 114.600 165.100 ;
        RECT 116.300 160.800 116.700 163.100 ;
        RECT 117.400 160.800 117.800 163.100 ;
        RECT 119.000 160.800 119.400 163.100 ;
        RECT 120.400 160.800 120.800 165.100 ;
        RECT 123.000 160.800 123.400 164.900 ;
        RECT 124.600 160.800 125.000 163.100 ;
        RECT 126.200 160.800 126.600 163.100 ;
        RECT 127.300 160.800 127.700 163.100 ;
        RECT 129.400 160.800 129.800 165.100 ;
        RECT 130.200 160.800 130.600 163.100 ;
        RECT 131.800 160.800 132.200 163.100 ;
        RECT 133.400 160.800 133.800 165.100 ;
        RECT 136.200 160.800 136.600 163.100 ;
        RECT 137.800 160.800 138.200 163.100 ;
        RECT 140.600 160.800 141.000 165.000 ;
        RECT 142.200 160.800 142.600 165.100 ;
        RECT 144.300 160.800 144.700 163.100 ;
        RECT 146.200 160.800 146.600 165.100 ;
        RECT 149.000 160.800 149.400 163.100 ;
        RECT 150.600 160.800 151.000 163.100 ;
        RECT 153.400 160.800 153.800 165.000 ;
        RECT 157.400 160.800 157.800 164.900 ;
        RECT 160.000 160.800 160.400 165.100 ;
        RECT 163.800 160.800 164.200 164.500 ;
        RECT 165.400 160.800 165.800 165.100 ;
        RECT 167.500 160.800 167.900 163.100 ;
        RECT 168.600 160.800 169.000 163.100 ;
        RECT 170.200 160.800 170.600 163.100 ;
        RECT 171.800 160.800 172.200 164.900 ;
        RECT 174.400 160.800 174.800 165.100 ;
        RECT 176.600 160.800 177.000 164.900 ;
        RECT 179.200 160.800 179.600 165.100 ;
        RECT 180.600 160.800 181.000 163.100 ;
        RECT 182.200 160.800 182.600 163.100 ;
        RECT 183.800 160.800 184.200 165.100 ;
        RECT 186.600 160.800 187.000 163.100 ;
        RECT 188.200 160.800 188.600 163.100 ;
        RECT 191.000 160.800 191.400 165.000 ;
        RECT 192.600 160.800 193.000 165.100 ;
        RECT 194.700 160.800 195.100 163.100 ;
        RECT 195.800 160.800 196.200 163.100 ;
        RECT 197.400 160.800 197.800 163.100 ;
        RECT 199.000 160.800 199.400 164.900 ;
        RECT 201.600 160.800 202.000 165.100 ;
        RECT 205.400 160.800 205.800 164.900 ;
        RECT 208.000 160.800 208.400 165.100 ;
        RECT 209.400 160.800 209.800 163.100 ;
        RECT 211.000 160.800 211.400 163.100 ;
        RECT 211.800 160.800 212.200 163.100 ;
        RECT 213.400 160.800 213.800 163.100 ;
        RECT 214.500 160.800 214.900 163.100 ;
        RECT 216.600 160.800 217.000 165.100 ;
        RECT 218.200 160.800 218.600 165.100 ;
        RECT 221.000 160.800 221.400 163.100 ;
        RECT 222.600 160.800 223.000 163.100 ;
        RECT 225.400 160.800 225.800 165.000 ;
        RECT 227.000 160.800 227.400 165.100 ;
        RECT 228.600 160.800 229.000 165.100 ;
        RECT 230.200 160.800 230.600 165.100 ;
        RECT 231.800 160.800 232.200 165.100 ;
        RECT 233.400 160.800 233.800 165.100 ;
        RECT 235.000 160.800 235.400 165.100 ;
        RECT 237.800 160.800 238.200 163.100 ;
        RECT 239.400 160.800 239.800 163.100 ;
        RECT 242.200 160.800 242.600 165.000 ;
        RECT 243.800 160.800 244.200 165.100 ;
        RECT 245.400 160.800 245.800 164.500 ;
        RECT 247.300 160.800 247.700 163.100 ;
        RECT 249.400 160.800 249.800 165.100 ;
        RECT 0.200 160.200 252.600 160.800 ;
        RECT 1.400 156.000 1.800 160.200 ;
        RECT 4.200 157.900 4.600 160.200 ;
        RECT 5.800 157.900 6.200 160.200 ;
        RECT 8.600 155.900 9.000 160.200 ;
        RECT 10.200 157.900 10.600 160.200 ;
        RECT 11.800 157.900 12.200 160.200 ;
        RECT 12.900 157.900 13.300 160.200 ;
        RECT 15.000 155.900 15.400 160.200 ;
        RECT 16.400 155.900 16.800 160.200 ;
        RECT 19.000 156.100 19.400 160.200 ;
        RECT 20.600 155.900 21.000 160.200 ;
        RECT 22.700 157.900 23.100 160.200 ;
        RECT 23.800 157.900 24.200 160.200 ;
        RECT 25.400 157.900 25.800 160.200 ;
        RECT 27.000 155.900 27.400 160.200 ;
        RECT 29.800 157.900 30.200 160.200 ;
        RECT 31.400 157.900 31.800 160.200 ;
        RECT 34.200 156.000 34.600 160.200 ;
        RECT 37.400 155.900 37.800 160.200 ;
        RECT 39.800 155.900 40.200 160.200 ;
        RECT 41.400 155.900 41.800 160.200 ;
        RECT 42.800 155.900 43.200 160.200 ;
        RECT 45.400 156.100 45.800 160.200 ;
        RECT 48.600 155.900 49.000 160.200 ;
        RECT 52.600 155.900 53.000 160.200 ;
        RECT 54.200 155.900 54.600 160.200 ;
        RECT 57.000 157.900 57.400 160.200 ;
        RECT 58.600 157.900 59.000 160.200 ;
        RECT 61.400 156.000 61.800 160.200 ;
        RECT 63.000 157.900 63.400 160.200 ;
        RECT 64.600 157.900 65.000 160.200 ;
        RECT 65.700 157.900 66.100 160.200 ;
        RECT 67.800 155.900 68.200 160.200 ;
        RECT 68.600 155.900 69.000 160.200 ;
        RECT 70.200 155.900 70.600 160.200 ;
        RECT 71.800 155.900 72.200 160.200 ;
        RECT 73.400 155.900 73.800 160.200 ;
        RECT 75.000 155.900 75.400 160.200 ;
        RECT 75.800 155.900 76.200 160.200 ;
        RECT 77.900 157.900 78.300 160.200 ;
        RECT 79.000 157.900 79.400 160.200 ;
        RECT 80.600 157.900 81.000 160.200 ;
        RECT 82.200 155.900 82.600 160.200 ;
        RECT 85.000 157.900 85.400 160.200 ;
        RECT 86.600 157.900 87.000 160.200 ;
        RECT 89.400 156.000 89.800 160.200 ;
        RECT 91.800 156.500 92.200 160.200 ;
        RECT 94.200 156.500 94.600 160.200 ;
        RECT 98.200 155.900 98.600 160.200 ;
        RECT 101.400 156.500 101.800 160.200 ;
        RECT 105.400 155.900 105.800 160.200 ;
        RECT 107.000 156.500 107.400 160.200 ;
        RECT 111.000 155.900 111.400 160.200 ;
        RECT 111.800 155.900 112.200 160.200 ;
        RECT 113.400 155.900 113.800 160.200 ;
        RECT 115.000 156.000 115.400 160.200 ;
        RECT 117.800 157.900 118.200 160.200 ;
        RECT 119.400 157.900 119.800 160.200 ;
        RECT 122.200 155.900 122.600 160.200 ;
        RECT 123.800 157.900 124.200 160.200 ;
        RECT 125.400 157.900 125.800 160.200 ;
        RECT 126.500 157.900 126.900 160.200 ;
        RECT 128.600 155.900 129.000 160.200 ;
        RECT 130.200 156.100 130.600 160.200 ;
        RECT 132.800 155.900 133.200 160.200 ;
        RECT 135.000 156.000 135.400 160.200 ;
        RECT 137.800 157.900 138.200 160.200 ;
        RECT 139.400 157.900 139.800 160.200 ;
        RECT 142.200 155.900 142.600 160.200 ;
        RECT 143.800 157.900 144.200 160.200 ;
        RECT 145.400 157.900 145.800 160.200 ;
        RECT 146.200 157.900 146.600 160.200 ;
        RECT 147.800 157.900 148.200 160.200 ;
        RECT 150.800 155.900 151.200 160.200 ;
        RECT 153.400 156.100 153.800 160.200 ;
        RECT 155.000 155.900 155.400 160.200 ;
        RECT 157.100 157.900 157.500 160.200 ;
        RECT 158.200 157.900 158.600 160.200 ;
        RECT 159.800 157.900 160.200 160.200 ;
        RECT 161.400 155.900 161.800 160.200 ;
        RECT 164.200 157.900 164.600 160.200 ;
        RECT 165.800 157.900 166.200 160.200 ;
        RECT 168.600 156.000 169.000 160.200 ;
        RECT 170.200 157.900 170.600 160.200 ;
        RECT 171.800 157.900 172.200 160.200 ;
        RECT 172.600 155.900 173.000 160.200 ;
        RECT 174.700 157.900 175.100 160.200 ;
        RECT 175.800 157.900 176.200 160.200 ;
        RECT 177.400 157.900 177.800 160.200 ;
        RECT 179.000 156.100 179.400 160.200 ;
        RECT 181.600 155.900 182.000 160.200 ;
        RECT 183.800 155.900 184.200 160.200 ;
        RECT 186.600 157.900 187.000 160.200 ;
        RECT 188.200 157.900 188.600 160.200 ;
        RECT 191.000 156.000 191.400 160.200 ;
        RECT 192.600 157.900 193.000 160.200 ;
        RECT 194.200 157.900 194.600 160.200 ;
        RECT 195.300 157.900 195.700 160.200 ;
        RECT 197.400 155.900 197.800 160.200 ;
        RECT 198.200 155.900 198.600 160.200 ;
        RECT 200.300 157.900 200.700 160.200 ;
        RECT 203.000 157.900 203.400 160.200 ;
        RECT 204.600 157.900 205.000 160.200 ;
        RECT 206.200 155.900 206.600 160.200 ;
        RECT 209.000 157.900 209.400 160.200 ;
        RECT 210.600 157.900 211.000 160.200 ;
        RECT 213.400 156.000 213.800 160.200 ;
        RECT 215.800 155.900 216.200 160.200 ;
        RECT 218.600 157.900 219.000 160.200 ;
        RECT 220.200 157.900 220.600 160.200 ;
        RECT 223.000 156.000 223.400 160.200 ;
        RECT 224.600 155.900 225.000 160.200 ;
        RECT 226.200 155.900 226.600 160.200 ;
        RECT 227.800 155.900 228.200 160.200 ;
        RECT 229.400 155.900 229.800 160.200 ;
        RECT 231.000 155.900 231.400 160.200 ;
        RECT 231.800 155.900 232.200 160.200 ;
        RECT 233.900 157.900 234.300 160.200 ;
        RECT 235.000 157.900 235.400 160.200 ;
        RECT 236.600 157.900 237.000 160.200 ;
        RECT 238.200 155.900 238.600 160.200 ;
        RECT 241.000 157.900 241.400 160.200 ;
        RECT 242.600 157.900 243.000 160.200 ;
        RECT 245.400 156.000 245.800 160.200 ;
        RECT 247.000 155.900 247.400 160.200 ;
        RECT 249.400 157.900 249.800 160.200 ;
        RECT 251.000 157.900 251.400 160.200 ;
        RECT 1.400 140.800 1.800 145.000 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.100 ;
        RECT 10.200 140.800 10.600 143.100 ;
        RECT 11.800 140.800 12.200 143.100 ;
        RECT 12.900 140.800 13.300 143.100 ;
        RECT 15.000 140.800 15.400 145.100 ;
        RECT 16.600 140.800 17.000 145.000 ;
        RECT 19.400 140.800 19.800 143.100 ;
        RECT 21.000 140.800 21.400 143.100 ;
        RECT 23.800 140.800 24.200 145.100 ;
        RECT 25.400 140.800 25.800 145.100 ;
        RECT 27.500 140.800 27.900 143.100 ;
        RECT 28.600 140.800 29.000 143.100 ;
        RECT 30.200 140.800 30.600 143.100 ;
        RECT 31.000 140.800 31.400 143.100 ;
        RECT 32.600 140.800 33.000 143.100 ;
        RECT 34.200 140.800 34.600 143.100 ;
        RECT 35.000 140.800 35.400 143.100 ;
        RECT 36.600 140.800 37.000 143.100 ;
        RECT 38.200 140.800 38.600 143.100 ;
        RECT 39.600 140.800 40.000 145.100 ;
        RECT 42.200 140.800 42.600 144.900 ;
        RECT 43.800 140.800 44.200 143.100 ;
        RECT 45.400 140.800 45.800 143.100 ;
        RECT 46.200 140.800 46.600 143.100 ;
        RECT 47.800 140.800 48.200 143.100 ;
        RECT 50.200 140.800 50.600 145.100 ;
        RECT 54.200 140.800 54.600 145.100 ;
        RECT 55.000 140.800 55.400 145.100 ;
        RECT 58.700 140.800 59.100 145.100 ;
        RECT 60.600 140.800 61.000 145.100 ;
        RECT 62.200 140.800 62.600 145.100 ;
        RECT 63.800 140.800 64.200 145.100 ;
        RECT 65.400 140.800 65.800 145.000 ;
        RECT 68.200 140.800 68.600 143.100 ;
        RECT 69.800 140.800 70.200 143.100 ;
        RECT 72.600 140.800 73.000 145.100 ;
        RECT 75.800 140.800 76.200 144.500 ;
        RECT 77.400 140.800 77.800 143.100 ;
        RECT 79.000 140.800 79.400 143.100 ;
        RECT 80.600 140.800 81.000 145.100 ;
        RECT 83.400 140.800 83.800 143.100 ;
        RECT 85.000 140.800 85.400 143.100 ;
        RECT 87.800 140.800 88.200 145.000 ;
        RECT 89.400 140.800 89.800 145.100 ;
        RECT 91.000 140.800 91.400 145.100 ;
        RECT 92.600 140.800 93.000 145.100 ;
        RECT 94.200 140.800 94.600 145.100 ;
        RECT 95.800 140.800 96.200 145.100 ;
        RECT 99.000 140.800 99.400 145.000 ;
        RECT 101.800 140.800 102.200 143.100 ;
        RECT 103.400 140.800 103.800 143.100 ;
        RECT 106.200 140.800 106.600 145.100 ;
        RECT 108.600 140.800 109.000 145.000 ;
        RECT 111.400 140.800 111.800 143.100 ;
        RECT 113.000 140.800 113.400 143.100 ;
        RECT 115.800 140.800 116.200 145.100 ;
        RECT 118.200 140.800 118.600 144.900 ;
        RECT 120.800 140.800 121.200 145.100 ;
        RECT 123.000 140.800 123.400 145.000 ;
        RECT 125.800 140.800 126.200 143.100 ;
        RECT 127.400 140.800 127.800 143.100 ;
        RECT 130.200 140.800 130.600 145.100 ;
        RECT 132.400 140.800 132.800 145.100 ;
        RECT 135.000 140.800 135.400 144.900 ;
        RECT 137.400 140.800 137.800 145.100 ;
        RECT 140.200 140.800 140.600 143.100 ;
        RECT 141.800 140.800 142.200 143.100 ;
        RECT 144.600 140.800 145.000 145.000 ;
        RECT 146.200 140.800 146.600 145.100 ;
        RECT 148.300 140.800 148.700 143.100 ;
        RECT 149.400 140.800 149.800 143.100 ;
        RECT 151.000 140.800 151.400 143.100 ;
        RECT 153.700 140.800 154.100 143.100 ;
        RECT 155.800 140.800 156.200 145.100 ;
        RECT 156.600 140.800 157.000 145.100 ;
        RECT 158.700 140.800 159.100 143.100 ;
        RECT 159.800 140.800 160.200 143.100 ;
        RECT 161.400 140.800 161.800 143.100 ;
        RECT 163.000 140.800 163.400 145.000 ;
        RECT 165.800 140.800 166.200 143.100 ;
        RECT 167.400 140.800 167.800 143.100 ;
        RECT 170.200 140.800 170.600 145.100 ;
        RECT 172.100 140.800 172.500 143.100 ;
        RECT 174.200 140.800 174.600 145.100 ;
        RECT 175.800 140.800 176.200 145.100 ;
        RECT 178.600 140.800 179.000 143.100 ;
        RECT 180.200 140.800 180.600 143.100 ;
        RECT 183.000 140.800 183.400 145.000 ;
        RECT 184.600 140.800 185.000 145.100 ;
        RECT 186.200 140.800 186.600 145.100 ;
        RECT 187.800 140.800 188.200 145.100 ;
        RECT 189.400 140.800 189.800 145.100 ;
        RECT 191.000 140.800 191.400 145.100 ;
        RECT 192.600 140.800 193.000 144.900 ;
        RECT 195.200 140.800 195.600 145.100 ;
        RECT 196.600 140.800 197.000 145.100 ;
        RECT 198.700 140.800 199.100 143.100 ;
        RECT 199.800 140.800 200.200 143.100 ;
        RECT 201.400 140.800 201.800 143.100 ;
        RECT 204.600 140.800 205.000 144.900 ;
        RECT 207.200 140.800 207.600 145.100 ;
        RECT 209.400 140.800 209.800 145.100 ;
        RECT 212.200 140.800 212.600 143.100 ;
        RECT 213.800 140.800 214.200 143.100 ;
        RECT 216.600 140.800 217.000 145.000 ;
        RECT 218.800 140.800 219.200 145.100 ;
        RECT 221.400 140.800 221.800 144.900 ;
        RECT 223.000 140.800 223.400 143.100 ;
        RECT 224.600 140.800 225.000 143.100 ;
        RECT 225.700 140.800 226.100 143.100 ;
        RECT 227.800 140.800 228.200 145.100 ;
        RECT 229.400 140.800 229.800 145.100 ;
        RECT 232.200 140.800 232.600 143.100 ;
        RECT 233.800 140.800 234.200 143.100 ;
        RECT 236.600 140.800 237.000 145.000 ;
        RECT 238.200 140.800 238.600 145.100 ;
        RECT 240.300 140.800 240.700 143.100 ;
        RECT 242.200 140.800 242.600 145.000 ;
        RECT 245.000 140.800 245.400 143.100 ;
        RECT 246.600 140.800 247.000 143.100 ;
        RECT 249.400 140.800 249.800 145.100 ;
        RECT 0.200 140.200 252.600 140.800 ;
        RECT 0.600 135.900 1.000 140.200 ;
        RECT 2.200 135.900 2.600 140.200 ;
        RECT 3.800 135.900 4.200 140.200 ;
        RECT 5.400 136.000 5.800 140.200 ;
        RECT 8.200 137.900 8.600 140.200 ;
        RECT 9.800 137.900 10.200 140.200 ;
        RECT 12.600 135.900 13.000 140.200 ;
        RECT 14.200 135.900 14.600 140.200 ;
        RECT 16.300 137.900 16.700 140.200 ;
        RECT 17.400 137.900 17.800 140.200 ;
        RECT 19.000 137.900 19.400 140.200 ;
        RECT 19.800 137.900 20.200 140.200 ;
        RECT 21.400 137.900 21.800 140.200 ;
        RECT 23.000 136.100 23.400 140.200 ;
        RECT 25.600 135.900 26.000 140.200 ;
        RECT 27.800 136.500 28.200 140.200 ;
        RECT 29.400 135.900 29.800 140.200 ;
        RECT 30.200 135.900 30.600 140.200 ;
        RECT 31.800 135.900 32.200 140.200 ;
        RECT 33.400 135.900 33.800 140.200 ;
        RECT 35.000 135.900 35.400 140.200 ;
        RECT 36.600 135.900 37.000 140.200 ;
        RECT 38.000 135.900 38.400 140.200 ;
        RECT 40.600 136.100 41.000 140.200 ;
        RECT 43.000 136.500 43.400 140.200 ;
        RECT 48.600 136.100 49.000 140.200 ;
        RECT 51.200 135.900 51.600 140.200 ;
        RECT 53.400 135.900 53.800 140.200 ;
        RECT 56.200 137.900 56.600 140.200 ;
        RECT 57.800 137.900 58.200 140.200 ;
        RECT 60.600 136.000 61.000 140.200 ;
        RECT 63.000 136.500 63.400 140.200 ;
        RECT 66.200 137.900 66.600 140.200 ;
        RECT 67.800 137.900 68.200 140.200 ;
        RECT 68.600 135.900 69.000 140.200 ;
        RECT 70.700 137.900 71.100 140.200 ;
        RECT 72.600 136.500 73.000 140.200 ;
        RECT 74.200 135.900 74.600 140.200 ;
        RECT 75.800 136.100 76.200 140.200 ;
        RECT 78.400 135.900 78.800 140.200 ;
        RECT 79.800 137.900 80.200 140.200 ;
        RECT 81.400 137.900 81.800 140.200 ;
        RECT 82.500 137.900 82.900 140.200 ;
        RECT 84.600 135.900 85.000 140.200 ;
        RECT 85.400 135.900 85.800 140.200 ;
        RECT 87.500 137.900 87.900 140.200 ;
        RECT 88.600 137.900 89.000 140.200 ;
        RECT 90.200 137.900 90.600 140.200 ;
        RECT 91.800 136.000 92.200 140.200 ;
        RECT 94.600 137.900 95.000 140.200 ;
        RECT 96.200 137.900 96.600 140.200 ;
        RECT 99.000 135.900 99.400 140.200 ;
        RECT 103.000 136.000 103.400 140.200 ;
        RECT 105.800 137.900 106.200 140.200 ;
        RECT 107.400 137.900 107.800 140.200 ;
        RECT 110.200 135.900 110.600 140.200 ;
        RECT 111.800 137.900 112.200 140.200 ;
        RECT 113.400 137.900 113.800 140.200 ;
        RECT 114.500 137.900 114.900 140.200 ;
        RECT 116.600 135.900 117.000 140.200 ;
        RECT 118.000 135.900 118.400 140.200 ;
        RECT 120.600 136.100 121.000 140.200 ;
        RECT 122.200 137.900 122.600 140.200 ;
        RECT 123.800 137.900 124.200 140.200 ;
        RECT 124.900 137.900 125.300 140.200 ;
        RECT 127.000 135.900 127.400 140.200 ;
        RECT 128.600 135.900 129.000 140.200 ;
        RECT 131.400 137.900 131.800 140.200 ;
        RECT 133.000 137.900 133.400 140.200 ;
        RECT 135.800 136.000 136.200 140.200 ;
        RECT 138.200 136.000 138.600 140.200 ;
        RECT 141.000 137.900 141.400 140.200 ;
        RECT 142.600 137.900 143.000 140.200 ;
        RECT 145.400 135.900 145.800 140.200 ;
        RECT 147.000 137.900 147.400 140.200 ;
        RECT 148.600 137.900 149.000 140.200 ;
        RECT 151.600 135.900 152.000 140.200 ;
        RECT 154.200 136.100 154.600 140.200 ;
        RECT 156.600 136.000 157.000 140.200 ;
        RECT 159.400 137.900 159.800 140.200 ;
        RECT 161.000 137.900 161.400 140.200 ;
        RECT 163.800 135.900 164.200 140.200 ;
        RECT 166.200 136.100 166.600 140.200 ;
        RECT 168.800 135.900 169.200 140.200 ;
        RECT 170.200 137.900 170.600 140.200 ;
        RECT 171.800 137.900 172.200 140.200 ;
        RECT 172.900 137.900 173.300 140.200 ;
        RECT 175.000 135.900 175.400 140.200 ;
        RECT 176.600 136.100 177.000 140.200 ;
        RECT 179.200 135.900 179.600 140.200 ;
        RECT 183.000 136.500 183.400 140.200 ;
        RECT 184.600 137.900 185.000 140.200 ;
        RECT 186.200 137.900 186.600 140.200 ;
        RECT 187.800 136.500 188.200 140.200 ;
        RECT 189.400 135.900 189.800 140.200 ;
        RECT 190.800 135.900 191.200 140.200 ;
        RECT 193.400 136.100 193.800 140.200 ;
        RECT 195.000 135.900 195.400 140.200 ;
        RECT 197.100 137.900 197.500 140.200 ;
        RECT 198.200 137.900 198.600 140.200 ;
        RECT 199.800 137.900 200.200 140.200 ;
        RECT 203.000 135.900 203.400 140.200 ;
        RECT 205.800 137.900 206.200 140.200 ;
        RECT 207.400 137.900 207.800 140.200 ;
        RECT 210.200 136.000 210.600 140.200 ;
        RECT 211.800 137.900 212.200 140.200 ;
        RECT 213.400 137.900 213.800 140.200 ;
        RECT 214.500 137.900 214.900 140.200 ;
        RECT 216.600 135.900 217.000 140.200 ;
        RECT 218.200 135.900 218.600 140.200 ;
        RECT 221.000 137.900 221.400 140.200 ;
        RECT 222.600 137.900 223.000 140.200 ;
        RECT 225.400 136.000 225.800 140.200 ;
        RECT 227.800 135.900 228.200 140.200 ;
        RECT 230.600 137.900 231.000 140.200 ;
        RECT 232.200 137.900 232.600 140.200 ;
        RECT 235.000 136.000 235.400 140.200 ;
        RECT 236.900 137.900 237.300 140.200 ;
        RECT 239.000 135.900 239.400 140.200 ;
        RECT 239.800 135.900 240.200 140.200 ;
        RECT 241.400 136.500 241.800 140.200 ;
        RECT 243.000 135.900 243.400 140.200 ;
        RECT 244.600 135.900 245.000 140.200 ;
        RECT 246.200 135.900 246.600 140.200 ;
        RECT 247.800 135.900 248.200 140.200 ;
        RECT 249.400 135.900 249.800 140.200 ;
        RECT 1.400 120.800 1.800 125.000 ;
        RECT 4.200 120.800 4.600 123.100 ;
        RECT 5.800 120.800 6.200 123.100 ;
        RECT 8.600 120.800 9.000 125.100 ;
        RECT 10.200 120.800 10.600 123.100 ;
        RECT 11.800 120.800 12.200 123.100 ;
        RECT 12.900 120.800 13.300 123.100 ;
        RECT 15.000 120.800 15.400 125.100 ;
        RECT 15.800 120.800 16.200 125.100 ;
        RECT 17.900 120.800 18.300 123.100 ;
        RECT 19.800 120.800 20.200 125.000 ;
        RECT 22.600 120.800 23.000 123.100 ;
        RECT 24.200 120.800 24.600 123.100 ;
        RECT 27.000 120.800 27.400 125.100 ;
        RECT 29.200 120.800 29.600 125.100 ;
        RECT 31.800 120.800 32.200 124.900 ;
        RECT 34.200 120.800 34.600 124.900 ;
        RECT 36.800 120.800 37.200 125.100 ;
        RECT 39.000 120.800 39.400 124.900 ;
        RECT 41.600 120.800 42.000 125.100 ;
        RECT 44.600 120.800 45.000 125.100 ;
        RECT 47.000 120.800 47.400 124.500 ;
        RECT 51.000 120.800 51.400 125.100 ;
        RECT 53.800 120.800 54.200 123.100 ;
        RECT 55.400 120.800 55.800 123.100 ;
        RECT 58.200 120.800 58.600 125.000 ;
        RECT 59.800 120.800 60.200 123.100 ;
        RECT 61.400 120.800 61.800 123.100 ;
        RECT 62.500 120.800 62.900 123.100 ;
        RECT 64.600 120.800 65.000 125.100 ;
        RECT 66.200 120.800 66.600 124.500 ;
        RECT 67.800 120.800 68.200 125.100 ;
        RECT 68.600 120.800 69.000 125.100 ;
        RECT 70.200 120.800 70.600 125.100 ;
        RECT 71.800 120.800 72.200 125.100 ;
        RECT 73.400 120.800 73.800 125.100 ;
        RECT 75.000 120.800 75.400 125.100 ;
        RECT 76.400 120.800 76.800 125.100 ;
        RECT 79.000 120.800 79.400 124.900 ;
        RECT 81.400 120.800 81.800 124.500 ;
        RECT 84.600 120.800 85.000 123.100 ;
        RECT 86.200 120.800 86.600 123.100 ;
        RECT 87.800 120.800 88.200 124.500 ;
        RECT 89.400 120.800 89.800 125.100 ;
        RECT 90.800 120.800 91.200 125.100 ;
        RECT 93.400 120.800 93.800 124.900 ;
        RECT 95.800 120.800 96.200 124.900 ;
        RECT 98.400 120.800 98.800 125.100 ;
        RECT 103.800 120.800 104.200 124.500 ;
        RECT 106.000 120.800 106.400 125.100 ;
        RECT 108.600 120.800 109.000 124.900 ;
        RECT 110.800 120.800 111.200 125.100 ;
        RECT 113.400 120.800 113.800 124.900 ;
        RECT 115.000 120.800 115.400 125.100 ;
        RECT 117.100 120.800 117.500 123.100 ;
        RECT 118.200 120.800 118.600 123.100 ;
        RECT 119.800 120.800 120.200 123.100 ;
        RECT 121.400 120.800 121.800 125.000 ;
        RECT 124.200 120.800 124.600 123.100 ;
        RECT 125.800 120.800 126.200 123.100 ;
        RECT 128.600 120.800 129.000 125.100 ;
        RECT 131.000 120.800 131.400 125.100 ;
        RECT 133.800 120.800 134.200 123.100 ;
        RECT 135.400 120.800 135.800 123.100 ;
        RECT 138.200 120.800 138.600 125.000 ;
        RECT 139.800 120.800 140.200 123.100 ;
        RECT 141.400 120.800 141.800 123.100 ;
        RECT 142.500 120.800 142.900 123.100 ;
        RECT 144.600 120.800 145.000 125.100 ;
        RECT 145.400 120.800 145.800 125.100 ;
        RECT 147.500 120.800 147.900 123.100 ;
        RECT 151.000 120.800 151.400 125.100 ;
        RECT 153.800 120.800 154.200 123.100 ;
        RECT 155.400 120.800 155.800 123.100 ;
        RECT 158.200 120.800 158.600 125.000 ;
        RECT 159.800 120.800 160.200 123.100 ;
        RECT 161.400 120.800 161.800 123.100 ;
        RECT 162.500 120.800 162.900 123.100 ;
        RECT 164.600 120.800 165.000 125.100 ;
        RECT 166.200 120.800 166.600 124.900 ;
        RECT 168.800 120.800 169.200 125.100 ;
        RECT 170.200 120.800 170.600 125.100 ;
        RECT 172.300 120.800 172.700 123.100 ;
        RECT 173.400 120.800 173.800 123.100 ;
        RECT 175.000 120.800 175.400 123.100 ;
        RECT 176.600 120.800 177.000 125.000 ;
        RECT 179.400 120.800 179.800 123.100 ;
        RECT 181.000 120.800 181.400 123.100 ;
        RECT 183.800 120.800 184.200 125.100 ;
        RECT 186.200 120.800 186.600 124.900 ;
        RECT 188.800 120.800 189.200 125.100 ;
        RECT 192.600 120.800 193.000 124.500 ;
        RECT 194.800 120.800 195.200 125.100 ;
        RECT 197.400 120.800 197.800 124.900 ;
        RECT 201.400 120.800 201.800 125.100 ;
        RECT 204.200 120.800 204.600 123.100 ;
        RECT 205.800 120.800 206.200 123.100 ;
        RECT 208.600 120.800 209.000 125.000 ;
        RECT 210.200 120.800 210.600 123.100 ;
        RECT 211.800 120.800 212.200 123.100 ;
        RECT 212.900 120.800 213.300 123.100 ;
        RECT 215.000 120.800 215.400 125.100 ;
        RECT 216.600 120.800 217.000 124.900 ;
        RECT 219.200 120.800 219.600 125.100 ;
        RECT 220.600 120.800 221.000 123.100 ;
        RECT 222.200 120.800 222.600 123.100 ;
        RECT 223.300 120.800 223.700 123.100 ;
        RECT 225.400 120.800 225.800 125.100 ;
        RECT 227.000 120.800 227.400 125.100 ;
        RECT 229.800 120.800 230.200 123.100 ;
        RECT 231.400 120.800 231.800 123.100 ;
        RECT 234.200 120.800 234.600 125.000 ;
        RECT 235.800 120.800 236.200 123.100 ;
        RECT 237.400 120.800 237.800 123.100 ;
        RECT 239.000 120.800 239.400 124.500 ;
        RECT 242.200 120.800 242.600 125.100 ;
        RECT 245.000 120.800 245.400 123.100 ;
        RECT 246.600 120.800 247.000 123.100 ;
        RECT 249.400 120.800 249.800 125.000 ;
        RECT 0.200 120.200 252.600 120.800 ;
        RECT 0.600 115.900 1.000 120.200 ;
        RECT 2.200 115.900 2.600 120.200 ;
        RECT 3.800 115.900 4.200 120.200 ;
        RECT 5.400 115.900 5.800 120.200 ;
        RECT 7.000 115.900 7.400 120.200 ;
        RECT 7.800 117.900 8.200 120.200 ;
        RECT 9.400 117.900 9.800 120.200 ;
        RECT 10.500 117.900 10.900 120.200 ;
        RECT 12.600 115.900 13.000 120.200 ;
        RECT 14.200 116.000 14.600 120.200 ;
        RECT 17.000 117.900 17.400 120.200 ;
        RECT 18.600 117.900 19.000 120.200 ;
        RECT 21.400 115.900 21.800 120.200 ;
        RECT 23.800 116.100 24.200 120.200 ;
        RECT 26.400 115.900 26.800 120.200 ;
        RECT 27.800 117.900 28.200 120.200 ;
        RECT 29.400 117.900 29.800 120.200 ;
        RECT 30.200 115.900 30.600 120.200 ;
        RECT 32.300 117.900 32.700 120.200 ;
        RECT 34.200 116.000 34.600 120.200 ;
        RECT 37.000 117.900 37.400 120.200 ;
        RECT 38.600 117.900 39.000 120.200 ;
        RECT 41.400 115.900 41.800 120.200 ;
        RECT 43.300 117.900 43.700 120.200 ;
        RECT 45.400 115.900 45.800 120.200 ;
        RECT 48.600 115.900 49.000 120.200 ;
        RECT 51.400 117.900 51.800 120.200 ;
        RECT 53.000 117.900 53.400 120.200 ;
        RECT 55.800 116.000 56.200 120.200 ;
        RECT 57.400 115.900 57.800 120.200 ;
        RECT 59.500 117.900 59.900 120.200 ;
        RECT 60.600 117.900 61.000 120.200 ;
        RECT 62.200 117.900 62.600 120.200 ;
        RECT 63.600 115.900 64.000 120.200 ;
        RECT 66.200 116.100 66.600 120.200 ;
        RECT 68.600 116.100 69.000 120.200 ;
        RECT 71.200 115.900 71.600 120.200 ;
        RECT 72.600 117.900 73.000 120.200 ;
        RECT 74.200 117.900 74.600 120.200 ;
        RECT 75.600 115.900 76.000 120.200 ;
        RECT 78.200 116.100 78.600 120.200 ;
        RECT 79.800 115.900 80.200 120.200 ;
        RECT 81.900 117.900 82.300 120.200 ;
        RECT 83.000 117.900 83.400 120.200 ;
        RECT 84.600 117.900 85.000 120.200 ;
        RECT 86.200 116.000 86.600 120.200 ;
        RECT 89.000 117.900 89.400 120.200 ;
        RECT 90.600 117.900 91.000 120.200 ;
        RECT 93.400 115.900 93.800 120.200 ;
        RECT 95.000 117.900 95.400 120.200 ;
        RECT 96.600 117.900 97.000 120.200 ;
        RECT 97.400 117.900 97.800 120.200 ;
        RECT 99.000 117.900 99.400 120.200 ;
        RECT 101.700 117.900 102.100 120.200 ;
        RECT 103.800 115.900 104.200 120.200 ;
        RECT 104.600 117.900 105.000 120.200 ;
        RECT 106.200 117.900 106.600 120.200 ;
        RECT 107.300 117.900 107.700 120.200 ;
        RECT 109.400 115.900 109.800 120.200 ;
        RECT 111.000 115.900 111.400 120.200 ;
        RECT 113.800 117.900 114.200 120.200 ;
        RECT 115.400 117.900 115.800 120.200 ;
        RECT 118.200 116.000 118.600 120.200 ;
        RECT 120.600 115.900 121.000 120.200 ;
        RECT 123.400 117.900 123.800 120.200 ;
        RECT 125.000 117.900 125.400 120.200 ;
        RECT 127.800 116.000 128.200 120.200 ;
        RECT 129.400 115.900 129.800 120.200 ;
        RECT 131.000 115.900 131.400 120.200 ;
        RECT 132.600 115.900 133.000 120.200 ;
        RECT 134.200 115.900 134.600 120.200 ;
        RECT 135.800 115.900 136.200 120.200 ;
        RECT 137.400 116.100 137.800 120.200 ;
        RECT 140.000 115.900 140.400 120.200 ;
        RECT 141.400 117.900 141.800 120.200 ;
        RECT 143.000 117.900 143.400 120.200 ;
        RECT 144.100 117.900 144.500 120.200 ;
        RECT 146.200 115.900 146.600 120.200 ;
        RECT 149.400 115.900 149.800 120.200 ;
        RECT 152.200 117.900 152.600 120.200 ;
        RECT 153.800 117.900 154.200 120.200 ;
        RECT 156.600 116.000 157.000 120.200 ;
        RECT 158.500 117.900 158.900 120.200 ;
        RECT 160.600 115.900 161.000 120.200 ;
        RECT 162.200 116.000 162.600 120.200 ;
        RECT 165.000 117.900 165.400 120.200 ;
        RECT 166.600 117.900 167.000 120.200 ;
        RECT 169.400 115.900 169.800 120.200 ;
        RECT 171.000 115.900 171.400 120.200 ;
        RECT 173.100 117.900 173.500 120.200 ;
        RECT 174.200 117.900 174.600 120.200 ;
        RECT 175.800 117.900 176.200 120.200 ;
        RECT 177.400 116.100 177.800 120.200 ;
        RECT 180.000 115.900 180.400 120.200 ;
        RECT 181.400 115.900 181.800 120.200 ;
        RECT 183.000 116.500 183.400 120.200 ;
        RECT 184.600 117.900 185.000 120.200 ;
        RECT 186.200 117.900 186.600 120.200 ;
        RECT 187.000 117.900 187.400 120.200 ;
        RECT 188.600 117.900 189.000 120.200 ;
        RECT 189.700 117.900 190.100 120.200 ;
        RECT 191.800 115.900 192.200 120.200 ;
        RECT 192.600 115.900 193.000 120.200 ;
        RECT 194.700 117.900 195.100 120.200 ;
        RECT 195.800 117.900 196.200 120.200 ;
        RECT 197.400 117.900 197.800 120.200 ;
        RECT 200.600 115.900 201.000 120.200 ;
        RECT 203.400 117.900 203.800 120.200 ;
        RECT 205.000 117.900 205.400 120.200 ;
        RECT 207.800 116.000 208.200 120.200 ;
        RECT 210.200 116.000 210.600 120.200 ;
        RECT 213.000 117.900 213.400 120.200 ;
        RECT 214.600 117.900 215.000 120.200 ;
        RECT 217.400 115.900 217.800 120.200 ;
        RECT 219.000 115.900 219.400 120.200 ;
        RECT 221.100 117.900 221.500 120.200 ;
        RECT 222.200 115.900 222.600 120.200 ;
        RECT 223.800 116.500 224.200 120.200 ;
        RECT 226.200 116.100 226.600 120.200 ;
        RECT 228.800 115.900 229.200 120.200 ;
        RECT 231.000 116.100 231.400 120.200 ;
        RECT 233.600 115.900 234.000 120.200 ;
        RECT 235.800 116.500 236.200 120.200 ;
        RECT 237.400 115.900 237.800 120.200 ;
        RECT 238.200 117.900 238.600 120.200 ;
        RECT 239.800 117.900 240.200 120.200 ;
        RECT 241.400 116.000 241.800 120.200 ;
        RECT 244.200 117.900 244.600 120.200 ;
        RECT 245.800 117.900 246.200 120.200 ;
        RECT 248.600 115.900 249.000 120.200 ;
        RECT 1.400 100.800 1.800 105.000 ;
        RECT 4.200 100.800 4.600 103.100 ;
        RECT 5.800 100.800 6.200 103.100 ;
        RECT 8.600 100.800 9.000 105.100 ;
        RECT 10.200 100.800 10.600 105.100 ;
        RECT 11.800 100.800 12.200 104.500 ;
        RECT 14.200 100.800 14.600 105.100 ;
        RECT 17.000 100.800 17.400 103.100 ;
        RECT 18.600 100.800 19.000 103.100 ;
        RECT 21.400 100.800 21.800 105.000 ;
        RECT 23.000 100.800 23.400 103.100 ;
        RECT 24.600 100.800 25.000 103.100 ;
        RECT 25.700 100.800 26.100 103.100 ;
        RECT 27.800 100.800 28.200 105.100 ;
        RECT 29.400 100.800 29.800 105.100 ;
        RECT 32.200 100.800 32.600 103.100 ;
        RECT 33.800 100.800 34.200 103.100 ;
        RECT 36.600 100.800 37.000 105.000 ;
        RECT 38.200 100.800 38.600 105.100 ;
        RECT 39.800 100.800 40.200 105.100 ;
        RECT 41.400 100.800 41.800 105.100 ;
        RECT 43.000 100.800 43.400 105.100 ;
        RECT 44.600 100.800 45.000 105.100 ;
        RECT 45.400 100.800 45.800 103.100 ;
        RECT 47.000 100.800 47.400 103.100 ;
        RECT 50.200 100.800 50.600 104.900 ;
        RECT 52.800 100.800 53.200 105.100 ;
        RECT 55.000 100.800 55.400 105.100 ;
        RECT 57.800 100.800 58.200 103.100 ;
        RECT 59.400 100.800 59.800 103.100 ;
        RECT 62.200 100.800 62.600 105.000 ;
        RECT 63.800 100.800 64.200 103.100 ;
        RECT 65.400 100.800 65.800 103.100 ;
        RECT 66.500 100.800 66.900 103.100 ;
        RECT 68.600 100.800 69.000 105.100 ;
        RECT 69.400 100.800 69.800 105.100 ;
        RECT 71.500 100.800 71.900 103.100 ;
        RECT 72.600 100.800 73.000 103.100 ;
        RECT 74.200 100.800 74.600 103.100 ;
        RECT 75.800 100.800 76.200 105.100 ;
        RECT 78.600 100.800 79.000 103.100 ;
        RECT 80.200 100.800 80.600 103.100 ;
        RECT 83.000 100.800 83.400 105.000 ;
        RECT 85.400 100.800 85.800 105.000 ;
        RECT 88.200 100.800 88.600 103.100 ;
        RECT 89.800 100.800 90.200 103.100 ;
        RECT 92.600 100.800 93.000 105.100 ;
        RECT 94.200 100.800 94.600 105.100 ;
        RECT 96.300 100.800 96.700 103.100 ;
        RECT 97.400 100.800 97.800 103.100 ;
        RECT 99.000 100.800 99.400 103.100 ;
        RECT 101.400 100.800 101.800 103.100 ;
        RECT 103.000 100.800 103.400 103.100 ;
        RECT 103.800 100.800 104.200 103.100 ;
        RECT 105.400 100.800 105.800 103.100 ;
        RECT 106.200 100.800 106.600 103.100 ;
        RECT 107.800 100.800 108.200 103.100 ;
        RECT 108.600 100.800 109.000 103.100 ;
        RECT 110.200 100.800 110.600 103.100 ;
        RECT 111.000 100.800 111.400 103.100 ;
        RECT 112.600 100.800 113.000 103.100 ;
        RECT 113.400 100.800 113.800 105.100 ;
        RECT 115.000 100.800 115.400 105.100 ;
        RECT 116.600 100.800 117.000 105.100 ;
        RECT 118.200 100.800 118.600 105.100 ;
        RECT 119.800 100.800 120.200 105.100 ;
        RECT 120.600 100.800 121.000 103.100 ;
        RECT 122.200 100.800 122.600 103.100 ;
        RECT 123.000 100.800 123.400 103.100 ;
        RECT 124.600 100.800 125.000 103.100 ;
        RECT 125.700 100.800 126.100 103.100 ;
        RECT 127.800 100.800 128.200 105.100 ;
        RECT 128.600 100.800 129.000 103.100 ;
        RECT 130.200 100.800 130.600 103.100 ;
        RECT 131.000 100.800 131.400 103.100 ;
        RECT 132.600 100.800 133.000 103.100 ;
        RECT 133.400 100.800 133.800 103.100 ;
        RECT 135.000 100.800 135.400 103.100 ;
        RECT 136.600 100.800 137.000 105.100 ;
        RECT 139.400 100.800 139.800 103.100 ;
        RECT 141.000 100.800 141.400 103.100 ;
        RECT 143.800 100.800 144.200 105.000 ;
        RECT 145.400 100.800 145.800 105.100 ;
        RECT 147.000 100.800 147.400 105.100 ;
        RECT 148.600 100.800 149.000 105.100 ;
        RECT 150.200 100.800 150.600 105.100 ;
        RECT 151.800 100.800 152.200 105.100 ;
        RECT 154.200 100.800 154.600 103.100 ;
        RECT 155.800 100.800 156.200 103.100 ;
        RECT 157.400 100.800 157.800 104.900 ;
        RECT 160.000 100.800 160.400 105.100 ;
        RECT 163.800 100.800 164.200 104.500 ;
        RECT 165.400 100.800 165.800 103.100 ;
        RECT 167.000 100.800 167.400 103.100 ;
        RECT 167.800 100.800 168.200 105.100 ;
        RECT 169.900 100.800 170.300 103.100 ;
        RECT 172.600 100.800 173.000 104.500 ;
        RECT 174.200 100.800 174.600 103.100 ;
        RECT 175.800 100.800 176.200 103.100 ;
        RECT 177.400 100.800 177.800 105.100 ;
        RECT 180.200 100.800 180.600 103.100 ;
        RECT 181.800 100.800 182.200 103.100 ;
        RECT 184.600 100.800 185.000 105.000 ;
        RECT 186.500 100.800 186.900 103.100 ;
        RECT 188.600 100.800 189.000 105.100 ;
        RECT 190.200 100.800 190.600 105.100 ;
        RECT 193.000 100.800 193.400 103.100 ;
        RECT 194.600 100.800 195.000 103.100 ;
        RECT 197.400 100.800 197.800 105.000 ;
        RECT 201.400 100.800 201.800 104.500 ;
        RECT 205.200 100.800 205.600 105.100 ;
        RECT 207.800 100.800 208.200 104.900 ;
        RECT 209.400 100.800 209.800 105.100 ;
        RECT 211.500 100.800 211.900 103.100 ;
        RECT 213.400 100.800 213.800 105.000 ;
        RECT 216.200 100.800 216.600 103.100 ;
        RECT 217.800 100.800 218.200 103.100 ;
        RECT 220.600 100.800 221.000 105.100 ;
        RECT 222.200 100.800 222.600 103.100 ;
        RECT 223.800 100.800 224.200 103.100 ;
        RECT 225.400 100.800 225.800 104.900 ;
        RECT 228.000 100.800 228.400 105.100 ;
        RECT 230.200 100.800 230.600 104.500 ;
        RECT 231.800 100.800 232.200 105.100 ;
        RECT 233.400 100.800 233.800 105.100 ;
        RECT 235.000 100.800 235.400 105.100 ;
        RECT 236.600 100.800 237.000 105.100 ;
        RECT 238.200 100.800 238.600 105.100 ;
        RECT 239.000 100.800 239.400 103.100 ;
        RECT 240.600 100.800 241.000 103.100 ;
        RECT 241.700 100.800 242.100 103.100 ;
        RECT 243.800 100.800 244.200 105.100 ;
        RECT 244.600 100.800 245.000 105.100 ;
        RECT 246.200 100.800 246.600 105.100 ;
        RECT 247.800 100.800 248.200 105.100 ;
        RECT 249.400 100.800 249.800 105.100 ;
        RECT 251.000 100.800 251.400 105.100 ;
        RECT 0.200 100.200 252.600 100.800 ;
        RECT 0.900 97.900 1.300 100.200 ;
        RECT 3.000 95.900 3.400 100.200 ;
        RECT 4.600 96.000 5.000 100.200 ;
        RECT 7.400 97.900 7.800 100.200 ;
        RECT 9.000 97.900 9.400 100.200 ;
        RECT 11.800 95.900 12.200 100.200 ;
        RECT 14.000 95.900 14.400 100.200 ;
        RECT 16.600 96.100 17.000 100.200 ;
        RECT 18.200 97.900 18.600 100.200 ;
        RECT 19.800 97.900 20.200 100.200 ;
        RECT 20.900 97.900 21.300 100.200 ;
        RECT 23.000 95.900 23.400 100.200 ;
        RECT 23.800 97.900 24.200 100.200 ;
        RECT 25.400 97.900 25.800 100.200 ;
        RECT 26.500 97.900 26.900 100.200 ;
        RECT 28.600 95.900 29.000 100.200 ;
        RECT 29.400 95.900 29.800 100.200 ;
        RECT 31.500 97.900 31.900 100.200 ;
        RECT 33.400 96.000 33.800 100.200 ;
        RECT 36.200 97.900 36.600 100.200 ;
        RECT 37.800 97.900 38.200 100.200 ;
        RECT 40.600 95.900 41.000 100.200 ;
        RECT 42.500 97.900 42.900 100.200 ;
        RECT 44.600 95.900 45.000 100.200 ;
        RECT 46.200 96.100 46.600 100.200 ;
        RECT 48.800 95.900 49.200 100.200 ;
        RECT 52.600 96.000 53.000 100.200 ;
        RECT 55.400 97.900 55.800 100.200 ;
        RECT 57.000 97.900 57.400 100.200 ;
        RECT 59.800 95.900 60.200 100.200 ;
        RECT 62.200 96.100 62.600 100.200 ;
        RECT 64.800 95.900 65.200 100.200 ;
        RECT 66.200 97.900 66.600 100.200 ;
        RECT 67.800 97.900 68.200 100.200 ;
        RECT 68.900 97.900 69.300 100.200 ;
        RECT 71.000 95.900 71.400 100.200 ;
        RECT 71.800 95.900 72.200 100.200 ;
        RECT 73.900 97.900 74.300 100.200 ;
        RECT 75.800 96.000 76.200 100.200 ;
        RECT 78.600 97.900 79.000 100.200 ;
        RECT 80.200 97.900 80.600 100.200 ;
        RECT 83.000 95.900 83.400 100.200 ;
        RECT 85.400 96.000 85.800 100.200 ;
        RECT 88.200 97.900 88.600 100.200 ;
        RECT 89.800 97.900 90.200 100.200 ;
        RECT 92.600 95.900 93.000 100.200 ;
        RECT 94.200 97.900 94.600 100.200 ;
        RECT 95.800 97.900 96.200 100.200 ;
        RECT 96.600 97.900 97.000 100.200 ;
        RECT 98.200 97.900 98.600 100.200 ;
        RECT 100.900 97.900 101.300 100.200 ;
        RECT 103.000 95.900 103.400 100.200 ;
        RECT 104.600 96.000 105.000 100.200 ;
        RECT 107.400 97.900 107.800 100.200 ;
        RECT 109.000 97.900 109.400 100.200 ;
        RECT 111.800 95.900 112.200 100.200 ;
        RECT 113.400 97.900 113.800 100.200 ;
        RECT 115.000 97.900 115.400 100.200 ;
        RECT 115.800 97.900 116.200 100.200 ;
        RECT 117.400 97.900 117.800 100.200 ;
        RECT 118.800 95.900 119.200 100.200 ;
        RECT 121.400 96.100 121.800 100.200 ;
        RECT 123.800 96.100 124.200 100.200 ;
        RECT 125.400 97.900 125.800 100.200 ;
        RECT 126.200 95.900 126.600 100.200 ;
        RECT 127.800 95.900 128.200 100.200 ;
        RECT 129.400 95.900 129.800 100.200 ;
        RECT 131.000 95.900 131.400 100.200 ;
        RECT 132.600 95.900 133.000 100.200 ;
        RECT 133.400 97.900 133.800 100.200 ;
        RECT 135.000 97.900 135.400 100.200 ;
        RECT 135.800 95.900 136.200 100.200 ;
        RECT 137.400 96.500 137.800 100.200 ;
        RECT 139.000 95.900 139.400 100.200 ;
        RECT 140.600 96.500 141.000 100.200 ;
        RECT 142.200 95.900 142.600 100.200 ;
        RECT 143.800 96.500 144.200 100.200 ;
        RECT 146.200 96.500 146.600 100.200 ;
        RECT 147.800 95.900 148.200 100.200 ;
        RECT 148.600 95.900 149.000 100.200 ;
        RECT 150.200 96.500 150.600 100.200 ;
        RECT 154.000 95.900 154.400 100.200 ;
        RECT 156.600 96.100 157.000 100.200 ;
        RECT 159.800 95.900 160.200 100.200 ;
        RECT 161.400 95.900 161.800 100.200 ;
        RECT 164.200 97.900 164.600 100.200 ;
        RECT 165.800 97.900 166.200 100.200 ;
        RECT 168.600 96.000 169.000 100.200 ;
        RECT 171.000 96.000 171.400 100.200 ;
        RECT 173.800 97.900 174.200 100.200 ;
        RECT 175.400 97.900 175.800 100.200 ;
        RECT 178.200 95.900 178.600 100.200 ;
        RECT 180.600 95.900 181.000 100.200 ;
        RECT 183.400 97.900 183.800 100.200 ;
        RECT 185.000 97.900 185.400 100.200 ;
        RECT 187.800 96.000 188.200 100.200 ;
        RECT 189.400 97.900 189.800 100.200 ;
        RECT 191.000 97.900 191.400 100.200 ;
        RECT 192.100 97.900 192.500 100.200 ;
        RECT 194.200 95.900 194.600 100.200 ;
        RECT 195.800 95.900 196.200 100.200 ;
        RECT 198.600 97.900 199.000 100.200 ;
        RECT 200.200 97.900 200.600 100.200 ;
        RECT 203.000 96.000 203.400 100.200 ;
        RECT 206.500 97.900 206.900 100.200 ;
        RECT 208.600 95.900 209.000 100.200 ;
        RECT 210.200 96.100 210.600 100.200 ;
        RECT 212.800 95.900 213.200 100.200 ;
        RECT 214.200 97.900 214.600 100.200 ;
        RECT 215.800 97.900 216.200 100.200 ;
        RECT 217.400 95.900 217.800 100.200 ;
        RECT 220.200 97.900 220.600 100.200 ;
        RECT 221.800 97.900 222.200 100.200 ;
        RECT 224.600 96.000 225.000 100.200 ;
        RECT 226.500 97.900 226.900 100.200 ;
        RECT 228.600 95.900 229.000 100.200 ;
        RECT 229.400 95.900 229.800 100.200 ;
        RECT 231.500 97.900 231.900 100.200 ;
        RECT 232.600 97.900 233.000 100.200 ;
        RECT 234.200 97.900 234.600 100.200 ;
        RECT 235.800 96.000 236.200 100.200 ;
        RECT 238.600 97.900 239.000 100.200 ;
        RECT 240.200 97.900 240.600 100.200 ;
        RECT 243.000 95.900 243.400 100.200 ;
        RECT 244.600 97.900 245.000 100.200 ;
        RECT 246.200 97.900 246.600 100.200 ;
        RECT 247.800 96.100 248.200 100.200 ;
        RECT 250.400 95.900 250.800 100.200 ;
        RECT 0.600 80.800 1.000 85.100 ;
        RECT 2.200 80.800 2.600 85.100 ;
        RECT 3.800 80.800 4.200 85.100 ;
        RECT 5.400 80.800 5.800 85.100 ;
        RECT 7.000 80.800 7.400 85.100 ;
        RECT 7.800 80.800 8.200 83.100 ;
        RECT 9.400 80.800 9.800 83.100 ;
        RECT 11.000 80.800 11.400 85.000 ;
        RECT 13.800 80.800 14.200 83.100 ;
        RECT 15.400 80.800 15.800 83.100 ;
        RECT 18.200 80.800 18.600 85.100 ;
        RECT 20.600 80.800 21.000 85.100 ;
        RECT 23.400 80.800 23.800 83.100 ;
        RECT 25.000 80.800 25.400 83.100 ;
        RECT 27.800 80.800 28.200 85.000 ;
        RECT 30.000 80.800 30.400 85.100 ;
        RECT 32.600 80.800 33.000 84.900 ;
        RECT 34.200 80.800 34.600 83.100 ;
        RECT 35.800 80.800 36.200 83.100 ;
        RECT 37.400 80.800 37.800 84.900 ;
        RECT 40.000 80.800 40.400 85.100 ;
        RECT 41.400 80.800 41.800 83.100 ;
        RECT 43.000 80.800 43.400 83.100 ;
        RECT 46.200 80.800 46.600 85.100 ;
        RECT 49.000 80.800 49.400 83.100 ;
        RECT 50.600 80.800 51.000 83.100 ;
        RECT 53.400 80.800 53.800 85.000 ;
        RECT 55.000 80.800 55.400 85.100 ;
        RECT 57.100 80.800 57.500 83.100 ;
        RECT 58.200 80.800 58.600 83.100 ;
        RECT 59.800 80.800 60.200 83.100 ;
        RECT 61.200 80.800 61.600 85.100 ;
        RECT 63.800 80.800 64.200 84.900 ;
        RECT 66.200 80.800 66.600 85.100 ;
        RECT 69.000 80.800 69.400 83.100 ;
        RECT 70.600 80.800 71.000 83.100 ;
        RECT 73.400 80.800 73.800 85.000 ;
        RECT 75.000 80.800 75.400 85.100 ;
        RECT 76.600 80.800 77.000 85.100 ;
        RECT 78.200 80.800 78.600 85.100 ;
        RECT 79.800 80.800 80.200 85.100 ;
        RECT 81.400 80.800 81.800 85.100 ;
        RECT 82.200 80.800 82.600 83.100 ;
        RECT 83.800 80.800 84.200 83.100 ;
        RECT 84.600 80.800 85.000 83.100 ;
        RECT 86.200 80.800 86.600 83.100 ;
        RECT 87.000 80.800 87.400 83.100 ;
        RECT 88.600 80.800 89.000 83.100 ;
        RECT 89.400 80.800 89.800 83.100 ;
        RECT 91.000 80.800 91.400 83.100 ;
        RECT 91.800 80.800 92.200 83.100 ;
        RECT 93.400 80.800 93.800 83.100 ;
        RECT 94.200 80.800 94.600 83.100 ;
        RECT 95.800 80.800 96.200 83.100 ;
        RECT 96.600 80.800 97.000 83.100 ;
        RECT 98.200 80.800 98.600 83.100 ;
        RECT 100.600 80.800 101.000 83.100 ;
        RECT 102.200 80.800 102.600 83.100 ;
        RECT 103.000 80.800 103.400 83.100 ;
        RECT 104.600 80.800 105.000 83.100 ;
        RECT 106.200 80.800 106.600 85.000 ;
        RECT 109.000 80.800 109.400 83.100 ;
        RECT 110.600 80.800 111.000 83.100 ;
        RECT 113.400 80.800 113.800 85.100 ;
        RECT 115.000 80.800 115.400 85.100 ;
        RECT 117.100 80.800 117.500 83.100 ;
        RECT 118.200 80.800 118.600 83.100 ;
        RECT 119.800 80.800 120.200 83.100 ;
        RECT 121.400 80.800 121.800 84.900 ;
        RECT 124.000 80.800 124.400 85.100 ;
        RECT 125.400 80.800 125.800 85.100 ;
        RECT 127.500 80.800 127.900 83.100 ;
        RECT 128.600 80.800 129.000 83.100 ;
        RECT 130.200 80.800 130.600 83.100 ;
        RECT 131.800 80.800 132.200 85.100 ;
        RECT 134.600 80.800 135.000 83.100 ;
        RECT 136.200 80.800 136.600 83.100 ;
        RECT 139.000 80.800 139.400 85.000 ;
        RECT 141.400 80.800 141.800 85.100 ;
        RECT 144.200 80.800 144.600 83.100 ;
        RECT 145.800 80.800 146.200 83.100 ;
        RECT 148.600 80.800 149.000 85.000 ;
        RECT 151.800 80.800 152.200 83.100 ;
        RECT 153.400 80.800 153.800 83.100 ;
        RECT 154.500 80.800 154.900 83.100 ;
        RECT 156.600 80.800 157.000 85.100 ;
        RECT 158.200 80.800 158.600 84.500 ;
        RECT 161.200 80.800 161.600 85.100 ;
        RECT 163.800 80.800 164.200 84.900 ;
        RECT 165.400 80.800 165.800 85.100 ;
        RECT 169.400 80.800 169.800 84.500 ;
        RECT 171.800 80.800 172.200 85.100 ;
        RECT 174.600 80.800 175.000 83.100 ;
        RECT 176.200 80.800 176.600 83.100 ;
        RECT 179.000 80.800 179.400 85.000 ;
        RECT 181.200 80.800 181.600 85.100 ;
        RECT 183.800 80.800 184.200 84.900 ;
        RECT 186.200 80.800 186.600 84.900 ;
        RECT 188.800 80.800 189.200 85.100 ;
        RECT 191.000 80.800 191.400 84.900 ;
        RECT 193.600 80.800 194.000 85.100 ;
        RECT 195.000 80.800 195.400 83.100 ;
        RECT 196.600 80.800 197.000 83.100 ;
        RECT 197.400 80.800 197.800 83.100 ;
        RECT 199.000 80.800 199.400 83.100 ;
        RECT 200.100 80.800 200.500 83.100 ;
        RECT 202.200 80.800 202.600 85.100 ;
        RECT 205.400 80.800 205.800 85.100 ;
        RECT 208.200 80.800 208.600 83.100 ;
        RECT 209.800 80.800 210.200 83.100 ;
        RECT 212.600 80.800 213.000 85.000 ;
        RECT 214.800 80.800 215.200 85.100 ;
        RECT 217.400 80.800 217.800 84.900 ;
        RECT 219.000 80.800 219.400 83.100 ;
        RECT 220.600 80.800 221.000 83.100 ;
        RECT 222.200 80.800 222.600 84.900 ;
        RECT 224.800 80.800 225.200 85.100 ;
        RECT 226.200 80.800 226.600 83.100 ;
        RECT 227.800 80.800 228.200 83.100 ;
        RECT 228.900 80.800 229.300 83.100 ;
        RECT 231.000 80.800 231.400 85.100 ;
        RECT 232.600 80.800 233.000 85.000 ;
        RECT 235.400 80.800 235.800 83.100 ;
        RECT 237.000 80.800 237.400 83.100 ;
        RECT 239.800 80.800 240.200 85.100 ;
        RECT 241.400 80.800 241.800 85.100 ;
        RECT 243.500 80.800 243.900 83.100 ;
        RECT 244.600 80.800 245.000 85.100 ;
        RECT 246.200 80.800 246.600 85.100 ;
        RECT 247.800 80.800 248.200 85.100 ;
        RECT 249.400 80.800 249.800 85.100 ;
        RECT 251.000 80.800 251.400 85.100 ;
        RECT 0.200 80.200 252.600 80.800 ;
        RECT 1.400 76.000 1.800 80.200 ;
        RECT 4.200 77.900 4.600 80.200 ;
        RECT 5.800 77.900 6.200 80.200 ;
        RECT 8.600 75.900 9.000 80.200 ;
        RECT 11.000 76.500 11.400 80.200 ;
        RECT 13.400 76.500 13.800 80.200 ;
        RECT 17.400 75.900 17.800 80.200 ;
        RECT 18.200 75.900 18.600 80.200 ;
        RECT 20.300 77.900 20.700 80.200 ;
        RECT 21.400 77.900 21.800 80.200 ;
        RECT 23.000 77.900 23.400 80.200 ;
        RECT 24.600 76.500 25.000 80.200 ;
        RECT 28.600 75.900 29.000 80.200 ;
        RECT 29.400 75.900 29.800 80.200 ;
        RECT 31.500 77.900 31.900 80.200 ;
        RECT 32.600 77.900 33.000 80.200 ;
        RECT 34.200 77.900 34.600 80.200 ;
        RECT 35.800 76.000 36.200 80.200 ;
        RECT 38.600 77.900 39.000 80.200 ;
        RECT 40.200 77.900 40.600 80.200 ;
        RECT 43.000 75.900 43.400 80.200 ;
        RECT 45.400 76.100 45.800 80.200 ;
        RECT 48.000 75.900 48.400 80.200 ;
        RECT 51.000 75.900 51.400 80.200 ;
        RECT 55.000 76.500 55.400 80.200 ;
        RECT 57.400 75.900 57.800 80.200 ;
        RECT 60.200 77.900 60.600 80.200 ;
        RECT 61.800 77.900 62.200 80.200 ;
        RECT 64.600 76.000 65.000 80.200 ;
        RECT 66.200 75.900 66.600 80.200 ;
        RECT 67.800 76.500 68.200 80.200 ;
        RECT 70.200 76.500 70.600 80.200 ;
        RECT 71.800 75.900 72.200 80.200 ;
        RECT 72.600 75.900 73.000 80.200 ;
        RECT 74.700 77.900 75.100 80.200 ;
        RECT 75.800 77.900 76.200 80.200 ;
        RECT 77.400 77.900 77.800 80.200 ;
        RECT 79.000 76.000 79.400 80.200 ;
        RECT 81.800 77.900 82.200 80.200 ;
        RECT 83.400 77.900 83.800 80.200 ;
        RECT 86.200 75.900 86.600 80.200 ;
        RECT 88.600 76.500 89.000 80.200 ;
        RECT 91.800 77.900 92.200 80.200 ;
        RECT 93.400 77.900 93.800 80.200 ;
        RECT 94.200 77.900 94.600 80.200 ;
        RECT 95.800 77.900 96.200 80.200 ;
        RECT 96.600 77.900 97.000 80.200 ;
        RECT 98.200 77.900 98.600 80.200 ;
        RECT 100.900 77.900 101.300 80.200 ;
        RECT 103.000 75.900 103.400 80.200 ;
        RECT 103.800 77.900 104.200 80.200 ;
        RECT 105.400 76.100 105.800 80.200 ;
        RECT 107.000 77.900 107.400 80.200 ;
        RECT 108.600 77.900 109.000 80.200 ;
        RECT 111.000 75.900 111.400 80.200 ;
        RECT 113.400 75.900 113.800 80.200 ;
        RECT 114.800 75.900 115.200 80.200 ;
        RECT 117.400 76.100 117.800 80.200 ;
        RECT 119.000 77.900 119.400 80.200 ;
        RECT 120.600 77.900 121.000 80.200 ;
        RECT 123.000 75.900 123.400 80.200 ;
        RECT 124.400 75.900 124.800 80.200 ;
        RECT 127.000 76.100 127.400 80.200 ;
        RECT 131.000 76.500 131.400 80.200 ;
        RECT 133.400 76.100 133.800 80.200 ;
        RECT 136.000 75.900 136.400 80.200 ;
        RECT 137.400 77.900 137.800 80.200 ;
        RECT 139.000 76.100 139.400 80.200 ;
        RECT 140.600 77.900 141.000 80.200 ;
        RECT 142.200 77.900 142.600 80.200 ;
        RECT 143.800 76.500 144.200 80.200 ;
        RECT 145.400 75.900 145.800 80.200 ;
        RECT 148.600 75.900 149.000 80.200 ;
        RECT 151.400 77.900 151.800 80.200 ;
        RECT 153.000 77.900 153.400 80.200 ;
        RECT 155.800 76.000 156.200 80.200 ;
        RECT 157.400 77.900 157.800 80.200 ;
        RECT 159.000 77.900 159.400 80.200 ;
        RECT 160.600 76.500 161.000 80.200 ;
        RECT 163.000 75.900 163.400 80.200 ;
        RECT 164.600 76.500 165.000 80.200 ;
        RECT 166.200 75.900 166.600 80.200 ;
        RECT 168.300 77.900 168.700 80.200 ;
        RECT 169.400 77.900 169.800 80.200 ;
        RECT 171.000 77.900 171.400 80.200 ;
        RECT 172.600 76.000 173.000 80.200 ;
        RECT 175.400 77.900 175.800 80.200 ;
        RECT 177.000 77.900 177.400 80.200 ;
        RECT 179.800 75.900 180.200 80.200 ;
        RECT 181.700 77.900 182.100 80.200 ;
        RECT 183.800 75.900 184.200 80.200 ;
        RECT 185.400 76.100 185.800 80.200 ;
        RECT 188.000 75.900 188.400 80.200 ;
        RECT 190.200 76.100 190.600 80.200 ;
        RECT 192.800 75.900 193.200 80.200 ;
        RECT 194.200 75.900 194.600 80.200 ;
        RECT 196.300 77.900 196.700 80.200 ;
        RECT 197.400 77.900 197.800 80.200 ;
        RECT 199.000 77.900 199.400 80.200 ;
        RECT 199.800 77.900 200.200 80.200 ;
        RECT 201.400 77.900 201.800 80.200 ;
        RECT 206.200 76.500 206.600 80.200 ;
        RECT 208.600 76.100 209.000 80.200 ;
        RECT 211.200 75.900 211.600 80.200 ;
        RECT 212.600 77.900 213.000 80.200 ;
        RECT 214.200 77.900 214.600 80.200 ;
        RECT 215.000 77.900 215.400 80.200 ;
        RECT 216.600 77.900 217.000 80.200 ;
        RECT 217.400 75.900 217.800 80.200 ;
        RECT 219.500 77.900 219.900 80.200 ;
        RECT 221.200 75.900 221.600 80.200 ;
        RECT 223.800 76.100 224.200 80.200 ;
        RECT 226.200 75.900 226.600 80.200 ;
        RECT 229.000 77.900 229.400 80.200 ;
        RECT 230.600 77.900 231.000 80.200 ;
        RECT 233.400 76.000 233.800 80.200 ;
        RECT 235.000 75.900 235.400 80.200 ;
        RECT 236.600 75.900 237.000 80.200 ;
        RECT 238.200 75.900 238.600 80.200 ;
        RECT 239.800 75.900 240.200 80.200 ;
        RECT 241.400 75.900 241.800 80.200 ;
        RECT 242.200 75.900 242.600 80.200 ;
        RECT 246.200 76.500 246.600 80.200 ;
        RECT 248.100 77.900 248.500 80.200 ;
        RECT 250.200 75.900 250.600 80.200 ;
        RECT 0.600 60.800 1.000 63.100 ;
        RECT 2.200 60.800 2.600 63.100 ;
        RECT 3.300 60.800 3.700 63.100 ;
        RECT 5.400 60.800 5.800 65.100 ;
        RECT 6.800 60.800 7.200 65.100 ;
        RECT 9.400 60.800 9.800 64.900 ;
        RECT 11.800 60.800 12.200 65.000 ;
        RECT 14.600 60.800 15.000 63.100 ;
        RECT 16.200 60.800 16.600 63.100 ;
        RECT 19.000 60.800 19.400 65.100 ;
        RECT 21.400 60.800 21.800 65.000 ;
        RECT 24.200 60.800 24.600 63.100 ;
        RECT 25.800 60.800 26.200 63.100 ;
        RECT 28.600 60.800 29.000 65.100 ;
        RECT 31.000 60.800 31.400 64.900 ;
        RECT 33.600 60.800 34.000 65.100 ;
        RECT 35.800 60.800 36.200 64.900 ;
        RECT 38.400 60.800 38.800 65.100 ;
        RECT 40.400 60.800 40.800 65.100 ;
        RECT 43.000 60.800 43.400 64.900 ;
        RECT 45.200 60.800 45.600 65.100 ;
        RECT 47.800 60.800 48.200 64.900 ;
        RECT 53.400 60.800 53.800 64.500 ;
        RECT 55.800 60.800 56.200 64.500 ;
        RECT 59.000 60.800 59.400 63.100 ;
        RECT 60.600 60.800 61.000 63.100 ;
        RECT 61.400 60.800 61.800 65.100 ;
        RECT 63.500 60.800 63.900 63.100 ;
        RECT 67.000 60.800 67.400 64.500 ;
        RECT 68.600 60.800 69.000 63.100 ;
        RECT 70.200 60.800 70.600 63.100 ;
        RECT 71.600 60.800 72.000 65.100 ;
        RECT 74.200 60.800 74.600 64.900 ;
        RECT 76.600 60.800 77.000 64.500 ;
        RECT 80.100 60.800 80.500 63.100 ;
        RECT 82.200 60.800 82.600 65.100 ;
        RECT 83.000 60.800 83.400 63.100 ;
        RECT 84.600 60.800 85.000 63.100 ;
        RECT 85.400 60.800 85.800 63.100 ;
        RECT 87.000 60.800 87.400 64.900 ;
        RECT 89.400 60.800 89.800 64.500 ;
        RECT 92.600 60.800 93.000 63.100 ;
        RECT 94.200 60.800 94.600 63.100 ;
        RECT 97.400 60.800 97.800 65.100 ;
        RECT 100.200 60.800 100.600 63.100 ;
        RECT 101.800 60.800 102.200 63.100 ;
        RECT 104.600 60.800 105.000 65.000 ;
        RECT 106.200 60.800 106.600 63.100 ;
        RECT 107.800 60.800 108.200 63.100 ;
        RECT 109.400 60.800 109.800 63.100 ;
        RECT 110.200 60.800 110.600 63.100 ;
        RECT 111.800 60.800 112.200 63.100 ;
        RECT 112.600 60.800 113.000 63.100 ;
        RECT 114.200 60.800 114.600 63.100 ;
        RECT 117.400 60.800 117.800 64.500 ;
        RECT 119.800 60.800 120.200 65.100 ;
        RECT 122.600 60.800 123.000 63.100 ;
        RECT 124.200 60.800 124.600 63.100 ;
        RECT 127.000 60.800 127.400 65.000 ;
        RECT 128.600 60.800 129.000 63.100 ;
        RECT 130.200 60.800 130.600 63.100 ;
        RECT 131.300 60.800 131.700 63.100 ;
        RECT 133.400 60.800 133.800 65.100 ;
        RECT 135.000 60.800 135.400 64.500 ;
        RECT 139.000 60.800 139.400 65.100 ;
        RECT 140.600 60.800 141.000 65.000 ;
        RECT 143.400 60.800 143.800 63.100 ;
        RECT 145.000 60.800 145.400 63.100 ;
        RECT 147.800 60.800 148.200 65.100 ;
        RECT 151.800 60.800 152.200 65.000 ;
        RECT 154.600 60.800 155.000 63.100 ;
        RECT 156.200 60.800 156.600 63.100 ;
        RECT 159.000 60.800 159.400 65.100 ;
        RECT 160.600 60.800 161.000 63.100 ;
        RECT 162.200 60.800 162.600 63.100 ;
        RECT 163.300 60.800 163.700 63.100 ;
        RECT 165.400 60.800 165.800 65.100 ;
        RECT 168.600 60.800 169.000 64.500 ;
        RECT 171.000 60.800 171.400 64.900 ;
        RECT 173.600 60.800 174.000 65.100 ;
        RECT 175.800 60.800 176.200 65.000 ;
        RECT 178.600 60.800 179.000 63.100 ;
        RECT 180.200 60.800 180.600 63.100 ;
        RECT 183.000 60.800 183.400 65.100 ;
        RECT 184.600 60.800 185.000 63.100 ;
        RECT 186.200 60.800 186.600 63.100 ;
        RECT 187.600 60.800 188.000 65.100 ;
        RECT 190.200 60.800 190.600 64.900 ;
        RECT 194.200 60.800 194.600 64.500 ;
        RECT 196.400 60.800 196.800 65.100 ;
        RECT 199.000 60.800 199.400 64.900 ;
        RECT 204.600 60.800 205.000 64.500 ;
        RECT 206.200 60.800 206.600 65.100 ;
        RECT 207.800 60.800 208.200 64.500 ;
        RECT 210.200 60.800 210.600 64.500 ;
        RECT 211.800 60.800 212.200 65.100 ;
        RECT 212.600 60.800 213.000 65.100 ;
        RECT 214.700 60.800 215.100 63.100 ;
        RECT 216.600 60.800 217.000 65.100 ;
        RECT 219.400 60.800 219.800 63.100 ;
        RECT 221.000 60.800 221.400 63.100 ;
        RECT 223.800 60.800 224.200 65.000 ;
        RECT 226.000 60.800 226.400 65.100 ;
        RECT 228.600 60.800 229.000 64.900 ;
        RECT 230.200 60.800 230.600 63.100 ;
        RECT 231.800 60.800 232.200 63.100 ;
        RECT 233.400 60.800 233.800 65.100 ;
        RECT 236.200 60.800 236.600 63.100 ;
        RECT 237.800 60.800 238.200 63.100 ;
        RECT 240.600 60.800 241.000 65.000 ;
        RECT 243.000 60.800 243.400 65.000 ;
        RECT 245.800 60.800 246.200 63.100 ;
        RECT 247.400 60.800 247.800 63.100 ;
        RECT 250.200 60.800 250.600 65.100 ;
        RECT 0.200 60.200 252.600 60.800 ;
        RECT 0.600 57.900 1.000 60.200 ;
        RECT 2.200 57.900 2.600 60.200 ;
        RECT 3.300 57.900 3.700 60.200 ;
        RECT 5.400 55.900 5.800 60.200 ;
        RECT 7.000 56.000 7.400 60.200 ;
        RECT 9.800 57.900 10.200 60.200 ;
        RECT 11.400 57.900 11.800 60.200 ;
        RECT 14.200 55.900 14.600 60.200 ;
        RECT 16.600 56.000 17.000 60.200 ;
        RECT 19.400 57.900 19.800 60.200 ;
        RECT 21.000 57.900 21.400 60.200 ;
        RECT 23.800 55.900 24.200 60.200 ;
        RECT 25.400 57.900 25.800 60.200 ;
        RECT 27.000 57.900 27.400 60.200 ;
        RECT 28.100 57.900 28.500 60.200 ;
        RECT 30.200 55.900 30.600 60.200 ;
        RECT 31.800 55.900 32.200 60.200 ;
        RECT 34.600 57.900 35.000 60.200 ;
        RECT 36.200 57.900 36.600 60.200 ;
        RECT 39.000 56.000 39.400 60.200 ;
        RECT 41.200 55.900 41.600 60.200 ;
        RECT 43.800 56.100 44.200 60.200 ;
        RECT 46.200 56.100 46.600 60.200 ;
        RECT 48.800 55.900 49.200 60.200 ;
        RECT 52.600 56.100 53.000 60.200 ;
        RECT 55.200 55.900 55.600 60.200 ;
        RECT 57.400 56.500 57.800 60.200 ;
        RECT 61.400 56.500 61.800 60.200 ;
        RECT 63.000 55.900 63.400 60.200 ;
        RECT 65.100 57.900 65.500 60.200 ;
        RECT 66.200 57.900 66.600 60.200 ;
        RECT 67.800 57.900 68.200 60.200 ;
        RECT 69.400 56.000 69.800 60.200 ;
        RECT 72.200 57.900 72.600 60.200 ;
        RECT 73.800 57.900 74.200 60.200 ;
        RECT 76.600 55.900 77.000 60.200 ;
        RECT 78.800 55.900 79.200 60.200 ;
        RECT 81.400 56.100 81.800 60.200 ;
        RECT 83.600 55.900 84.000 60.200 ;
        RECT 86.200 56.100 86.600 60.200 ;
        RECT 88.600 56.100 89.000 60.200 ;
        RECT 91.200 55.900 91.600 60.200 ;
        RECT 93.400 56.100 93.800 60.200 ;
        RECT 96.000 55.900 96.400 60.200 ;
        RECT 99.800 55.900 100.200 60.200 ;
        RECT 102.600 57.900 103.000 60.200 ;
        RECT 104.200 57.900 104.600 60.200 ;
        RECT 107.000 56.000 107.400 60.200 ;
        RECT 108.600 57.900 109.000 60.200 ;
        RECT 110.200 57.900 110.600 60.200 ;
        RECT 111.300 57.900 111.700 60.200 ;
        RECT 113.400 55.900 113.800 60.200 ;
        RECT 114.200 55.900 114.600 60.200 ;
        RECT 116.600 57.900 117.000 60.200 ;
        RECT 118.200 57.900 118.600 60.200 ;
        RECT 119.800 57.900 120.200 60.200 ;
        RECT 121.400 56.100 121.800 60.200 ;
        RECT 124.000 55.900 124.400 60.200 ;
        RECT 125.400 57.900 125.800 60.200 ;
        RECT 127.000 57.900 127.400 60.200 ;
        RECT 128.100 57.900 128.500 60.200 ;
        RECT 130.200 55.900 130.600 60.200 ;
        RECT 131.800 56.000 132.200 60.200 ;
        RECT 134.600 57.900 135.000 60.200 ;
        RECT 136.200 57.900 136.600 60.200 ;
        RECT 139.000 55.900 139.400 60.200 ;
        RECT 141.400 56.500 141.800 60.200 ;
        RECT 145.400 55.900 145.800 60.200 ;
        RECT 146.800 55.900 147.200 60.200 ;
        RECT 149.400 56.100 149.800 60.200 ;
        RECT 152.600 55.900 153.000 60.200 ;
        RECT 154.700 57.900 155.100 60.200 ;
        RECT 155.800 57.900 156.200 60.200 ;
        RECT 157.400 57.900 157.800 60.200 ;
        RECT 159.000 56.000 159.400 60.200 ;
        RECT 161.800 57.900 162.200 60.200 ;
        RECT 163.400 57.900 163.800 60.200 ;
        RECT 166.200 55.900 166.600 60.200 ;
        RECT 168.600 55.900 169.000 60.200 ;
        RECT 171.400 57.900 171.800 60.200 ;
        RECT 173.000 57.900 173.400 60.200 ;
        RECT 175.800 56.000 176.200 60.200 ;
        RECT 178.200 56.000 178.600 60.200 ;
        RECT 181.000 57.900 181.400 60.200 ;
        RECT 182.600 57.900 183.000 60.200 ;
        RECT 185.400 55.900 185.800 60.200 ;
        RECT 188.600 56.500 189.000 60.200 ;
        RECT 191.800 55.900 192.200 60.200 ;
        RECT 193.200 55.900 193.600 60.200 ;
        RECT 195.800 56.100 196.200 60.200 ;
        RECT 197.400 55.900 197.800 60.200 ;
        RECT 201.400 56.500 201.800 60.200 ;
        RECT 205.400 56.500 205.800 60.200 ;
        RECT 207.000 55.900 207.400 60.200 ;
        RECT 207.800 55.900 208.200 60.200 ;
        RECT 209.400 55.900 209.800 60.200 ;
        RECT 211.000 55.900 211.400 60.200 ;
        RECT 212.600 55.900 213.000 60.200 ;
        RECT 214.200 55.900 214.600 60.200 ;
        RECT 215.800 55.900 216.200 60.200 ;
        RECT 218.600 57.900 219.000 60.200 ;
        RECT 220.200 57.900 220.600 60.200 ;
        RECT 223.000 56.000 223.400 60.200 ;
        RECT 226.200 56.500 226.600 60.200 ;
        RECT 228.600 55.900 229.000 60.200 ;
        RECT 231.400 57.900 231.800 60.200 ;
        RECT 233.000 57.900 233.400 60.200 ;
        RECT 235.800 56.000 236.200 60.200 ;
        RECT 237.700 57.900 238.100 60.200 ;
        RECT 239.800 55.900 240.200 60.200 ;
        RECT 241.400 55.900 241.800 60.200 ;
        RECT 244.200 57.900 244.600 60.200 ;
        RECT 245.800 57.900 246.200 60.200 ;
        RECT 248.600 56.000 249.000 60.200 ;
        RECT 1.400 40.800 1.800 44.500 ;
        RECT 3.000 40.800 3.400 45.100 ;
        RECT 4.600 40.800 5.000 45.100 ;
        RECT 6.200 40.800 6.600 45.100 ;
        RECT 7.800 40.800 8.200 45.100 ;
        RECT 9.400 40.800 9.800 45.100 ;
        RECT 10.200 40.800 10.600 43.100 ;
        RECT 11.800 40.800 12.200 43.100 ;
        RECT 12.900 40.800 13.300 43.100 ;
        RECT 15.000 40.800 15.400 45.100 ;
        RECT 16.600 40.800 17.000 45.000 ;
        RECT 19.400 40.800 19.800 43.100 ;
        RECT 21.000 40.800 21.400 43.100 ;
        RECT 23.800 40.800 24.200 45.100 ;
        RECT 26.000 40.800 26.400 45.100 ;
        RECT 28.600 40.800 29.000 44.900 ;
        RECT 30.200 40.800 30.600 43.100 ;
        RECT 31.800 40.800 32.200 43.100 ;
        RECT 32.900 40.800 33.300 43.100 ;
        RECT 35.000 40.800 35.400 45.100 ;
        RECT 36.600 40.800 37.000 45.100 ;
        RECT 39.400 40.800 39.800 43.100 ;
        RECT 41.000 40.800 41.400 43.100 ;
        RECT 43.800 40.800 44.200 45.000 ;
        RECT 45.400 40.800 45.800 43.100 ;
        RECT 47.000 40.800 47.400 43.100 ;
        RECT 49.400 40.800 49.800 43.100 ;
        RECT 51.000 40.800 51.400 43.100 ;
        RECT 52.600 40.800 53.000 45.100 ;
        RECT 55.400 40.800 55.800 43.100 ;
        RECT 57.000 40.800 57.400 43.100 ;
        RECT 59.800 40.800 60.200 45.000 ;
        RECT 62.200 40.800 62.600 45.000 ;
        RECT 65.000 40.800 65.400 43.100 ;
        RECT 66.600 40.800 67.000 43.100 ;
        RECT 69.400 40.800 69.800 45.100 ;
        RECT 71.000 40.800 71.400 45.100 ;
        RECT 73.100 40.800 73.500 43.100 ;
        RECT 74.200 40.800 74.600 43.100 ;
        RECT 75.800 40.800 76.200 43.100 ;
        RECT 77.400 40.800 77.800 45.000 ;
        RECT 80.200 40.800 80.600 43.100 ;
        RECT 81.800 40.800 82.200 43.100 ;
        RECT 84.600 40.800 85.000 45.100 ;
        RECT 86.200 40.800 86.600 43.100 ;
        RECT 87.800 40.800 88.200 43.100 ;
        RECT 88.900 40.800 89.300 43.100 ;
        RECT 91.000 40.800 91.400 45.100 ;
        RECT 92.600 40.800 93.000 45.100 ;
        RECT 95.400 40.800 95.800 43.100 ;
        RECT 97.000 40.800 97.400 43.100 ;
        RECT 99.800 40.800 100.200 45.000 ;
        RECT 103.000 40.800 103.400 43.100 ;
        RECT 104.600 40.800 105.000 43.100 ;
        RECT 105.700 40.800 106.100 43.100 ;
        RECT 107.800 40.800 108.200 45.100 ;
        RECT 108.600 40.800 109.000 45.100 ;
        RECT 110.200 40.800 110.600 44.500 ;
        RECT 111.800 40.800 112.200 45.100 ;
        RECT 113.400 40.800 113.800 45.100 ;
        RECT 115.000 40.800 115.400 45.100 ;
        RECT 116.600 40.800 117.000 45.100 ;
        RECT 118.200 40.800 118.600 45.100 ;
        RECT 119.000 40.800 119.400 45.100 ;
        RECT 121.100 40.800 121.500 43.100 ;
        RECT 122.200 40.800 122.600 43.100 ;
        RECT 123.800 40.800 124.200 43.100 ;
        RECT 125.400 40.800 125.800 45.100 ;
        RECT 128.200 40.800 128.600 43.100 ;
        RECT 129.800 40.800 130.200 43.100 ;
        RECT 132.600 40.800 133.000 45.000 ;
        RECT 135.000 40.800 135.400 44.500 ;
        RECT 136.600 40.800 137.000 45.100 ;
        RECT 137.400 40.800 137.800 43.100 ;
        RECT 139.000 40.800 139.400 43.100 ;
        RECT 140.600 40.800 141.000 45.000 ;
        RECT 143.400 40.800 143.800 43.100 ;
        RECT 145.000 40.800 145.400 43.100 ;
        RECT 147.800 40.800 148.200 45.100 ;
        RECT 151.600 40.800 152.000 45.100 ;
        RECT 154.200 40.800 154.600 44.900 ;
        RECT 155.800 40.800 156.200 43.100 ;
        RECT 157.400 40.800 157.800 43.100 ;
        RECT 158.500 40.800 158.900 43.100 ;
        RECT 160.600 40.800 161.000 45.100 ;
        RECT 161.400 40.800 161.800 45.100 ;
        RECT 163.000 40.800 163.400 44.500 ;
        RECT 164.600 40.800 165.000 45.100 ;
        RECT 166.200 40.800 166.600 44.500 ;
        RECT 167.800 40.800 168.200 45.100 ;
        RECT 169.400 40.800 169.800 44.500 ;
        RECT 171.800 40.800 172.200 44.500 ;
        RECT 173.400 40.800 173.800 45.100 ;
        RECT 175.000 40.800 175.400 44.500 ;
        RECT 176.600 40.800 177.000 45.100 ;
        RECT 177.400 40.800 177.800 45.100 ;
        RECT 179.000 40.800 179.400 44.500 ;
        RECT 180.600 40.800 181.000 45.100 ;
        RECT 182.200 40.800 182.600 45.100 ;
        RECT 183.800 40.800 184.200 45.100 ;
        RECT 185.400 40.800 185.800 45.100 ;
        RECT 187.000 40.800 187.400 45.100 ;
        RECT 188.600 40.800 189.000 44.900 ;
        RECT 191.200 40.800 191.600 45.100 ;
        RECT 193.400 40.800 193.800 45.100 ;
        RECT 196.200 40.800 196.600 43.100 ;
        RECT 197.800 40.800 198.200 43.100 ;
        RECT 200.600 40.800 201.000 45.000 ;
        RECT 204.400 40.800 204.800 45.100 ;
        RECT 207.000 40.800 207.400 44.900 ;
        RECT 209.400 40.800 209.800 45.100 ;
        RECT 212.200 40.800 212.600 43.100 ;
        RECT 213.800 40.800 214.200 43.100 ;
        RECT 216.600 40.800 217.000 45.000 ;
        RECT 218.200 40.800 218.600 43.100 ;
        RECT 219.800 40.800 220.200 43.100 ;
        RECT 220.900 40.800 221.300 43.100 ;
        RECT 223.000 40.800 223.400 45.100 ;
        RECT 223.800 40.800 224.200 45.100 ;
        RECT 227.000 40.800 227.400 44.900 ;
        RECT 229.600 40.800 230.000 45.100 ;
        RECT 231.600 40.800 232.000 45.100 ;
        RECT 234.200 40.800 234.600 44.900 ;
        RECT 235.800 40.800 236.200 45.100 ;
        RECT 237.900 40.800 238.300 43.100 ;
        RECT 239.000 40.800 239.400 43.100 ;
        RECT 240.600 40.800 241.000 43.100 ;
        RECT 242.200 40.800 242.600 45.000 ;
        RECT 245.000 40.800 245.400 43.100 ;
        RECT 246.600 40.800 247.000 43.100 ;
        RECT 249.400 40.800 249.800 45.100 ;
        RECT 0.200 40.200 252.600 40.800 ;
        RECT 1.400 36.000 1.800 40.200 ;
        RECT 4.200 37.900 4.600 40.200 ;
        RECT 5.800 37.900 6.200 40.200 ;
        RECT 8.600 35.900 9.000 40.200 ;
        RECT 10.800 35.900 11.200 40.200 ;
        RECT 13.400 36.100 13.800 40.200 ;
        RECT 15.000 35.900 15.400 40.200 ;
        RECT 17.100 37.900 17.500 40.200 ;
        RECT 18.200 37.900 18.600 40.200 ;
        RECT 19.800 37.900 20.200 40.200 ;
        RECT 21.400 36.000 21.800 40.200 ;
        RECT 24.200 37.900 24.600 40.200 ;
        RECT 25.800 37.900 26.200 40.200 ;
        RECT 28.600 35.900 29.000 40.200 ;
        RECT 31.000 36.100 31.400 40.200 ;
        RECT 33.600 35.900 34.000 40.200 ;
        RECT 35.600 35.900 36.000 40.200 ;
        RECT 38.200 36.100 38.600 40.200 ;
        RECT 39.800 37.900 40.200 40.200 ;
        RECT 41.400 37.900 41.800 40.200 ;
        RECT 42.500 37.900 42.900 40.200 ;
        RECT 44.600 35.900 45.000 40.200 ;
        RECT 45.400 35.900 45.800 40.200 ;
        RECT 47.000 36.500 47.400 40.200 ;
        RECT 50.200 37.900 50.600 40.200 ;
        RECT 51.800 37.900 52.200 40.200 ;
        RECT 52.900 37.900 53.300 40.200 ;
        RECT 55.000 35.900 55.400 40.200 ;
        RECT 56.600 36.100 57.000 40.200 ;
        RECT 59.200 35.900 59.600 40.200 ;
        RECT 61.200 35.900 61.600 40.200 ;
        RECT 63.800 36.100 64.200 40.200 ;
        RECT 66.000 35.900 66.400 40.200 ;
        RECT 68.600 36.100 69.000 40.200 ;
        RECT 70.200 35.900 70.600 40.200 ;
        RECT 71.800 36.500 72.200 40.200 ;
        RECT 74.200 36.000 74.600 40.200 ;
        RECT 77.000 37.900 77.400 40.200 ;
        RECT 78.600 37.900 79.000 40.200 ;
        RECT 81.400 35.900 81.800 40.200 ;
        RECT 83.000 37.900 83.400 40.200 ;
        RECT 84.600 37.900 85.000 40.200 ;
        RECT 86.200 36.500 86.600 40.200 ;
        RECT 88.600 35.900 89.000 40.200 ;
        RECT 91.600 35.900 92.000 40.200 ;
        RECT 94.200 36.100 94.600 40.200 ;
        RECT 95.800 35.900 96.200 40.200 ;
        RECT 97.400 36.500 97.800 40.200 ;
        RECT 101.200 35.900 101.600 40.200 ;
        RECT 103.800 36.100 104.200 40.200 ;
        RECT 105.400 35.900 105.800 40.200 ;
        RECT 107.500 37.900 107.900 40.200 ;
        RECT 108.600 37.900 109.000 40.200 ;
        RECT 110.200 37.900 110.600 40.200 ;
        RECT 111.800 36.000 112.200 40.200 ;
        RECT 114.600 37.900 115.000 40.200 ;
        RECT 116.200 37.900 116.600 40.200 ;
        RECT 119.000 35.900 119.400 40.200 ;
        RECT 121.400 36.100 121.800 40.200 ;
        RECT 124.000 35.900 124.400 40.200 ;
        RECT 126.000 35.900 126.400 40.200 ;
        RECT 128.600 36.100 129.000 40.200 ;
        RECT 131.000 35.900 131.400 40.200 ;
        RECT 133.800 37.900 134.200 40.200 ;
        RECT 135.400 37.900 135.800 40.200 ;
        RECT 138.200 36.000 138.600 40.200 ;
        RECT 139.800 37.900 140.200 40.200 ;
        RECT 141.400 37.900 141.800 40.200 ;
        RECT 142.200 35.900 142.600 40.200 ;
        RECT 143.800 35.900 144.200 40.200 ;
        RECT 145.200 35.900 145.600 40.200 ;
        RECT 147.800 36.100 148.200 40.200 ;
        RECT 151.800 35.900 152.200 40.200 ;
        RECT 154.600 37.900 155.000 40.200 ;
        RECT 156.200 37.900 156.600 40.200 ;
        RECT 159.000 36.000 159.400 40.200 ;
        RECT 160.600 35.900 161.000 40.200 ;
        RECT 162.200 36.500 162.600 40.200 ;
        RECT 164.600 36.500 165.000 40.200 ;
        RECT 166.200 35.900 166.600 40.200 ;
        RECT 167.000 37.900 167.400 40.200 ;
        RECT 168.600 37.900 169.000 40.200 ;
        RECT 170.200 36.100 170.600 40.200 ;
        RECT 172.800 35.900 173.200 40.200 ;
        RECT 175.000 36.500 175.400 40.200 ;
        RECT 176.600 35.900 177.000 40.200 ;
        RECT 178.200 36.100 178.600 40.200 ;
        RECT 180.800 35.900 181.200 40.200 ;
        RECT 182.200 37.900 182.600 40.200 ;
        RECT 183.800 37.900 184.200 40.200 ;
        RECT 184.900 37.900 185.300 40.200 ;
        RECT 187.000 35.900 187.400 40.200 ;
        RECT 188.600 35.900 189.000 40.200 ;
        RECT 191.400 37.900 191.800 40.200 ;
        RECT 193.000 37.900 193.400 40.200 ;
        RECT 195.800 36.000 196.200 40.200 ;
        RECT 198.200 36.100 198.600 40.200 ;
        RECT 200.800 35.900 201.200 40.200 ;
        RECT 204.600 35.900 205.000 40.200 ;
        RECT 207.400 37.900 207.800 40.200 ;
        RECT 209.000 37.900 209.400 40.200 ;
        RECT 211.800 36.000 212.200 40.200 ;
        RECT 213.400 37.900 213.800 40.200 ;
        RECT 215.000 37.900 215.400 40.200 ;
        RECT 216.600 36.100 217.000 40.200 ;
        RECT 219.200 35.900 219.600 40.200 ;
        RECT 220.600 35.900 221.000 40.200 ;
        RECT 222.700 37.900 223.100 40.200 ;
        RECT 223.800 37.900 224.200 40.200 ;
        RECT 225.400 37.900 225.800 40.200 ;
        RECT 226.800 35.900 227.200 40.200 ;
        RECT 229.400 36.100 229.800 40.200 ;
        RECT 231.000 35.900 231.400 40.200 ;
        RECT 235.000 36.500 235.400 40.200 ;
        RECT 236.600 35.900 237.000 40.200 ;
        RECT 238.700 37.900 239.100 40.200 ;
        RECT 239.800 37.900 240.200 40.200 ;
        RECT 241.400 37.900 241.800 40.200 ;
        RECT 243.000 36.000 243.400 40.200 ;
        RECT 245.800 37.900 246.200 40.200 ;
        RECT 247.400 37.900 247.800 40.200 ;
        RECT 250.200 35.900 250.600 40.200 ;
        RECT 0.600 20.800 1.000 23.100 ;
        RECT 2.200 20.800 2.600 23.100 ;
        RECT 3.300 20.800 3.700 23.100 ;
        RECT 5.400 20.800 5.800 25.100 ;
        RECT 6.200 20.800 6.600 23.100 ;
        RECT 7.800 20.800 8.200 23.100 ;
        RECT 8.900 20.800 9.300 23.100 ;
        RECT 11.000 20.800 11.400 25.100 ;
        RECT 12.600 20.800 13.000 25.000 ;
        RECT 15.400 20.800 15.800 23.100 ;
        RECT 17.000 20.800 17.400 23.100 ;
        RECT 19.800 20.800 20.200 25.100 ;
        RECT 22.200 20.800 22.600 25.000 ;
        RECT 25.000 20.800 25.400 23.100 ;
        RECT 26.600 20.800 27.000 23.100 ;
        RECT 29.400 20.800 29.800 25.100 ;
        RECT 31.800 20.800 32.200 25.100 ;
        RECT 34.600 20.800 35.000 23.100 ;
        RECT 36.200 20.800 36.600 23.100 ;
        RECT 39.000 20.800 39.400 25.000 ;
        RECT 41.400 20.800 41.800 25.100 ;
        RECT 44.200 20.800 44.600 23.100 ;
        RECT 45.800 20.800 46.200 23.100 ;
        RECT 48.600 20.800 49.000 25.000 ;
        RECT 52.600 20.800 53.000 24.900 ;
        RECT 55.200 20.800 55.600 25.100 ;
        RECT 56.600 20.800 57.000 25.100 ;
        RECT 58.700 20.800 59.100 23.100 ;
        RECT 59.800 20.800 60.200 23.100 ;
        RECT 61.400 20.800 61.800 23.100 ;
        RECT 63.000 20.800 63.400 25.000 ;
        RECT 65.800 20.800 66.200 23.100 ;
        RECT 67.400 20.800 67.800 23.100 ;
        RECT 70.200 20.800 70.600 25.100 ;
        RECT 72.400 20.800 72.800 25.100 ;
        RECT 75.000 20.800 75.400 24.900 ;
        RECT 76.600 20.800 77.000 23.100 ;
        RECT 78.200 20.800 78.600 23.100 ;
        RECT 79.300 20.800 79.700 23.100 ;
        RECT 81.400 20.800 81.800 25.100 ;
        RECT 82.200 20.800 82.600 25.100 ;
        RECT 84.300 20.800 84.700 23.100 ;
        RECT 86.200 20.800 86.600 25.100 ;
        RECT 89.000 20.800 89.400 23.100 ;
        RECT 90.600 20.800 91.000 23.100 ;
        RECT 93.400 20.800 93.800 25.000 ;
        RECT 97.400 20.800 97.800 25.100 ;
        RECT 100.200 20.800 100.600 23.100 ;
        RECT 101.800 20.800 102.200 23.100 ;
        RECT 104.600 20.800 105.000 25.000 ;
        RECT 106.200 20.800 106.600 23.100 ;
        RECT 107.800 20.800 108.200 23.100 ;
        RECT 108.900 20.800 109.300 23.100 ;
        RECT 111.000 20.800 111.400 25.100 ;
        RECT 111.800 20.800 112.200 25.100 ;
        RECT 113.900 20.800 114.300 23.100 ;
        RECT 115.000 20.800 115.400 23.100 ;
        RECT 116.600 20.800 117.000 23.100 ;
        RECT 118.200 20.800 118.600 25.000 ;
        RECT 121.000 20.800 121.400 23.100 ;
        RECT 122.600 20.800 123.000 23.100 ;
        RECT 125.400 20.800 125.800 25.100 ;
        RECT 127.000 20.800 127.400 25.100 ;
        RECT 129.100 20.800 129.500 23.100 ;
        RECT 130.200 20.800 130.600 23.100 ;
        RECT 131.800 20.800 132.200 23.100 ;
        RECT 133.400 20.800 133.800 25.000 ;
        RECT 136.200 20.800 136.600 23.100 ;
        RECT 137.800 20.800 138.200 23.100 ;
        RECT 140.600 20.800 141.000 25.100 ;
        RECT 142.500 20.800 142.900 23.100 ;
        RECT 144.600 20.800 145.000 25.100 ;
        RECT 146.200 20.800 146.600 24.900 ;
        RECT 148.800 20.800 149.200 25.100 ;
        RECT 152.600 20.800 153.000 24.900 ;
        RECT 155.200 20.800 155.600 25.100 ;
        RECT 157.400 20.800 157.800 24.500 ;
        RECT 159.000 20.800 159.400 25.100 ;
        RECT 159.800 20.800 160.200 23.100 ;
        RECT 161.400 20.800 161.800 23.100 ;
        RECT 162.500 20.800 162.900 23.100 ;
        RECT 164.600 20.800 165.000 25.100 ;
        RECT 166.200 20.800 166.600 24.500 ;
        RECT 167.800 20.800 168.200 25.100 ;
        RECT 168.900 20.800 169.300 23.100 ;
        RECT 171.000 20.800 171.400 25.100 ;
        RECT 172.600 20.800 173.000 25.100 ;
        RECT 175.400 20.800 175.800 23.100 ;
        RECT 177.000 20.800 177.400 23.100 ;
        RECT 179.800 20.800 180.200 25.000 ;
        RECT 181.400 20.800 181.800 23.100 ;
        RECT 183.000 20.800 183.400 23.100 ;
        RECT 184.100 20.800 184.500 23.100 ;
        RECT 186.200 20.800 186.600 25.100 ;
        RECT 187.800 20.800 188.200 25.100 ;
        RECT 190.600 20.800 191.000 23.100 ;
        RECT 192.200 20.800 192.600 23.100 ;
        RECT 195.000 20.800 195.400 25.000 ;
        RECT 197.400 20.800 197.800 24.900 ;
        RECT 200.000 20.800 200.400 25.100 ;
        RECT 203.800 20.800 204.200 24.500 ;
        RECT 205.400 20.800 205.800 25.100 ;
        RECT 206.200 20.800 206.600 23.100 ;
        RECT 207.800 20.800 208.200 23.100 ;
        RECT 208.900 20.800 209.300 23.100 ;
        RECT 211.000 20.800 211.400 25.100 ;
        RECT 211.800 20.800 212.200 25.100 ;
        RECT 213.900 20.800 214.300 23.100 ;
        RECT 215.000 20.800 215.400 25.100 ;
        RECT 216.600 20.800 217.000 24.500 ;
        RECT 219.000 20.800 219.400 25.100 ;
        RECT 221.800 20.800 222.200 23.100 ;
        RECT 223.400 20.800 223.800 23.100 ;
        RECT 226.200 20.800 226.600 25.000 ;
        RECT 227.800 20.800 228.200 23.100 ;
        RECT 229.400 20.800 229.800 23.100 ;
        RECT 231.000 20.800 231.400 25.100 ;
        RECT 233.800 20.800 234.200 23.100 ;
        RECT 235.400 20.800 235.800 23.100 ;
        RECT 238.200 20.800 238.600 25.000 ;
        RECT 240.600 20.800 241.000 25.100 ;
        RECT 243.400 20.800 243.800 23.100 ;
        RECT 245.000 20.800 245.400 23.100 ;
        RECT 247.800 20.800 248.200 25.000 ;
        RECT 249.400 20.800 249.800 25.100 ;
        RECT 251.500 20.800 251.900 23.100 ;
        RECT 0.200 20.200 252.600 20.800 ;
        RECT 1.400 15.900 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 16.000 9.000 20.200 ;
        RECT 10.200 17.900 10.600 20.200 ;
        RECT 11.800 17.900 12.200 20.200 ;
        RECT 12.900 17.900 13.300 20.200 ;
        RECT 15.000 15.900 15.400 20.200 ;
        RECT 15.800 17.900 16.200 20.200 ;
        RECT 17.400 17.900 17.800 20.200 ;
        RECT 19.000 16.500 19.400 20.200 ;
        RECT 23.000 15.900 23.400 20.200 ;
        RECT 24.600 16.000 25.000 20.200 ;
        RECT 27.400 17.900 27.800 20.200 ;
        RECT 29.000 17.900 29.400 20.200 ;
        RECT 31.800 15.900 32.200 20.200 ;
        RECT 33.400 15.900 33.800 20.200 ;
        RECT 35.000 15.900 35.400 20.200 ;
        RECT 36.600 15.900 37.000 20.200 ;
        RECT 38.200 15.900 38.600 20.200 ;
        RECT 39.800 15.900 40.200 20.200 ;
        RECT 40.600 15.900 41.000 20.200 ;
        RECT 42.200 15.900 42.600 20.200 ;
        RECT 43.800 15.900 44.200 20.200 ;
        RECT 45.200 15.900 45.600 20.200 ;
        RECT 47.800 16.100 48.200 20.200 ;
        RECT 51.800 16.500 52.200 20.200 ;
        RECT 53.400 15.900 53.800 20.200 ;
        RECT 55.000 15.900 55.400 20.200 ;
        RECT 56.600 15.900 57.000 20.200 ;
        RECT 58.200 15.900 58.600 20.200 ;
        RECT 59.800 15.900 60.200 20.200 ;
        RECT 60.600 17.900 61.000 20.200 ;
        RECT 62.200 17.900 62.600 20.200 ;
        RECT 63.300 17.900 63.700 20.200 ;
        RECT 65.400 15.900 65.800 20.200 ;
        RECT 66.800 15.900 67.200 20.200 ;
        RECT 69.400 16.100 69.800 20.200 ;
        RECT 71.800 16.000 72.200 20.200 ;
        RECT 74.600 17.900 75.000 20.200 ;
        RECT 76.200 17.900 76.600 20.200 ;
        RECT 79.000 15.900 79.400 20.200 ;
        RECT 80.600 17.900 81.000 20.200 ;
        RECT 82.200 17.900 82.600 20.200 ;
        RECT 83.300 17.900 83.700 20.200 ;
        RECT 85.400 15.900 85.800 20.200 ;
        RECT 86.200 15.900 86.600 20.200 ;
        RECT 87.800 15.900 88.200 20.200 ;
        RECT 89.400 15.900 89.800 20.200 ;
        RECT 90.200 15.900 90.600 20.200 ;
        RECT 91.800 15.900 92.200 20.200 ;
        RECT 93.400 15.900 93.800 20.200 ;
        RECT 95.000 15.900 95.400 20.200 ;
        RECT 96.600 15.900 97.000 20.200 ;
        RECT 99.600 15.900 100.000 20.200 ;
        RECT 102.200 16.100 102.600 20.200 ;
        RECT 104.400 15.900 104.800 20.200 ;
        RECT 107.000 16.100 107.400 20.200 ;
        RECT 108.600 17.900 109.000 20.200 ;
        RECT 110.200 17.900 110.600 20.200 ;
        RECT 111.300 17.900 111.700 20.200 ;
        RECT 113.400 15.900 113.800 20.200 ;
        RECT 115.000 15.900 115.400 20.200 ;
        RECT 117.800 17.900 118.200 20.200 ;
        RECT 119.400 17.900 119.800 20.200 ;
        RECT 122.200 16.000 122.600 20.200 ;
        RECT 124.600 16.100 125.000 20.200 ;
        RECT 127.200 15.900 127.600 20.200 ;
        RECT 129.400 15.900 129.800 20.200 ;
        RECT 132.200 17.900 132.600 20.200 ;
        RECT 133.800 17.900 134.200 20.200 ;
        RECT 136.600 16.000 137.000 20.200 ;
        RECT 138.200 17.900 138.600 20.200 ;
        RECT 139.800 17.900 140.200 20.200 ;
        RECT 140.900 17.900 141.300 20.200 ;
        RECT 143.000 15.900 143.400 20.200 ;
        RECT 143.800 17.900 144.200 20.200 ;
        RECT 145.400 17.900 145.800 20.200 ;
        RECT 146.200 17.900 146.600 20.200 ;
        RECT 147.800 17.900 148.200 20.200 ;
        RECT 150.800 15.900 151.200 20.200 ;
        RECT 153.400 16.100 153.800 20.200 ;
        RECT 155.000 17.900 155.400 20.200 ;
        RECT 156.600 17.900 157.000 20.200 ;
        RECT 157.700 17.900 158.100 20.200 ;
        RECT 159.800 15.900 160.200 20.200 ;
        RECT 161.400 16.000 161.800 20.200 ;
        RECT 164.200 17.900 164.600 20.200 ;
        RECT 165.800 17.900 166.200 20.200 ;
        RECT 168.600 15.900 169.000 20.200 ;
        RECT 170.200 17.900 170.600 20.200 ;
        RECT 171.800 17.900 172.200 20.200 ;
        RECT 172.900 17.900 173.300 20.200 ;
        RECT 175.000 15.900 175.400 20.200 ;
        RECT 176.600 15.900 177.000 20.200 ;
        RECT 179.400 17.900 179.800 20.200 ;
        RECT 181.000 17.900 181.400 20.200 ;
        RECT 183.800 16.000 184.200 20.200 ;
        RECT 185.400 15.900 185.800 20.200 ;
        RECT 187.500 17.900 187.900 20.200 ;
        RECT 188.600 17.900 189.000 20.200 ;
        RECT 190.200 17.900 190.600 20.200 ;
        RECT 191.800 16.000 192.200 20.200 ;
        RECT 194.600 17.900 195.000 20.200 ;
        RECT 196.200 17.900 196.600 20.200 ;
        RECT 199.000 15.900 199.400 20.200 ;
        RECT 202.800 15.900 203.200 20.200 ;
        RECT 205.400 16.100 205.800 20.200 ;
        RECT 207.000 15.900 207.400 20.200 ;
        RECT 208.600 16.500 209.000 20.200 ;
        RECT 211.000 16.100 211.400 20.200 ;
        RECT 213.600 15.900 214.000 20.200 ;
        RECT 215.000 15.900 215.400 20.200 ;
        RECT 217.100 17.900 217.500 20.200 ;
        RECT 218.200 17.900 218.600 20.200 ;
        RECT 219.800 17.900 220.200 20.200 ;
        RECT 220.600 15.900 221.000 20.200 ;
        RECT 222.700 17.900 223.100 20.200 ;
        RECT 223.800 17.900 224.200 20.200 ;
        RECT 225.400 17.900 225.800 20.200 ;
        RECT 227.000 15.900 227.400 20.200 ;
        RECT 229.800 17.900 230.200 20.200 ;
        RECT 231.400 17.900 231.800 20.200 ;
        RECT 234.200 16.000 234.600 20.200 ;
        RECT 235.800 15.900 236.200 20.200 ;
        RECT 237.400 15.900 237.800 20.200 ;
        RECT 239.000 15.900 239.400 20.200 ;
        RECT 240.600 15.900 241.000 20.200 ;
        RECT 242.200 15.900 242.600 20.200 ;
        RECT 243.000 15.900 243.400 20.200 ;
        RECT 244.600 15.900 245.000 20.200 ;
        RECT 246.200 15.900 246.600 20.200 ;
        RECT 247.800 15.900 248.200 20.200 ;
        RECT 249.400 15.900 249.800 20.200 ;
        RECT 250.200 17.900 250.600 20.200 ;
        RECT 251.800 17.900 252.200 20.200 ;
        RECT 0.600 0.800 1.000 5.100 ;
        RECT 2.200 0.800 2.600 5.100 ;
        RECT 3.800 0.800 4.200 5.100 ;
        RECT 5.400 0.800 5.800 5.100 ;
        RECT 7.000 0.800 7.400 5.100 ;
        RECT 7.800 0.800 8.200 5.100 ;
        RECT 9.400 0.800 9.800 5.100 ;
        RECT 11.000 0.800 11.400 5.100 ;
        RECT 12.600 0.800 13.000 5.100 ;
        RECT 14.200 0.800 14.600 5.100 ;
        RECT 15.000 0.800 15.400 5.100 ;
        RECT 17.100 0.800 17.500 3.100 ;
        RECT 19.000 0.800 19.400 5.000 ;
        RECT 21.800 0.800 22.200 3.100 ;
        RECT 23.400 0.800 23.800 3.100 ;
        RECT 26.200 0.800 26.600 5.100 ;
        RECT 29.400 0.800 29.800 5.100 ;
        RECT 31.800 0.800 32.200 4.500 ;
        RECT 34.200 0.800 34.600 5.000 ;
        RECT 37.000 0.800 37.400 3.100 ;
        RECT 38.600 0.800 39.000 3.100 ;
        RECT 41.400 0.800 41.800 5.100 ;
        RECT 43.000 0.800 43.400 5.100 ;
        RECT 45.100 0.800 45.500 3.100 ;
        RECT 46.200 0.800 46.600 3.100 ;
        RECT 47.800 0.800 48.200 3.100 ;
        RECT 51.000 0.800 51.400 5.100 ;
        RECT 53.800 0.800 54.200 3.100 ;
        RECT 55.400 0.800 55.800 3.100 ;
        RECT 58.200 0.800 58.600 5.000 ;
        RECT 60.600 0.800 61.000 5.100 ;
        RECT 63.400 0.800 63.800 3.100 ;
        RECT 65.000 0.800 65.400 3.100 ;
        RECT 67.800 0.800 68.200 5.000 ;
        RECT 70.200 0.800 70.600 4.500 ;
        RECT 71.800 0.800 72.200 5.100 ;
        RECT 73.400 0.800 73.800 5.000 ;
        RECT 76.200 0.800 76.600 3.100 ;
        RECT 77.800 0.800 78.200 3.100 ;
        RECT 80.600 0.800 81.000 5.100 ;
        RECT 82.200 0.800 82.600 3.100 ;
        RECT 83.800 0.800 84.200 3.100 ;
        RECT 84.900 0.800 85.300 3.100 ;
        RECT 87.000 0.800 87.400 5.100 ;
        RECT 88.600 0.800 89.000 4.500 ;
        RECT 90.200 0.800 90.600 5.100 ;
        RECT 91.800 0.800 92.200 5.100 ;
        RECT 94.600 0.800 95.000 3.100 ;
        RECT 96.200 0.800 96.600 3.100 ;
        RECT 99.000 0.800 99.400 5.000 ;
        RECT 102.200 0.800 102.600 3.100 ;
        RECT 103.800 0.800 104.200 3.100 ;
        RECT 104.900 0.800 105.300 3.100 ;
        RECT 107.000 0.800 107.400 5.100 ;
        RECT 107.800 0.800 108.200 5.100 ;
        RECT 109.400 0.800 109.800 5.100 ;
        RECT 111.000 0.800 111.400 5.100 ;
        RECT 112.600 0.800 113.000 5.100 ;
        RECT 114.200 0.800 114.600 5.100 ;
        RECT 115.800 0.800 116.200 5.000 ;
        RECT 118.600 0.800 119.000 3.100 ;
        RECT 120.200 0.800 120.600 3.100 ;
        RECT 123.000 0.800 123.400 5.100 ;
        RECT 124.600 0.800 125.000 3.100 ;
        RECT 126.200 0.800 126.600 3.100 ;
        RECT 127.300 0.800 127.700 3.100 ;
        RECT 129.400 0.800 129.800 5.100 ;
        RECT 131.000 0.800 131.400 5.000 ;
        RECT 133.800 0.800 134.200 3.100 ;
        RECT 135.400 0.800 135.800 3.100 ;
        RECT 138.200 0.800 138.600 5.100 ;
        RECT 140.100 0.800 140.500 3.100 ;
        RECT 142.200 0.800 142.600 5.100 ;
        RECT 143.000 0.800 143.400 5.100 ;
        RECT 145.100 0.800 145.500 3.100 ;
        RECT 148.600 0.800 149.000 5.100 ;
        RECT 151.400 0.800 151.800 3.100 ;
        RECT 153.000 0.800 153.400 3.100 ;
        RECT 155.800 0.800 156.200 5.000 ;
        RECT 157.400 0.800 157.800 5.100 ;
        RECT 159.000 0.800 159.400 5.100 ;
        RECT 160.600 0.800 161.000 5.100 ;
        RECT 162.200 0.800 162.600 5.100 ;
        RECT 163.800 0.800 164.200 5.100 ;
        RECT 164.600 0.800 165.000 5.100 ;
        RECT 166.700 0.800 167.100 3.100 ;
        RECT 167.800 0.800 168.200 3.100 ;
        RECT 169.400 0.800 169.800 3.100 ;
        RECT 171.000 0.800 171.400 5.100 ;
        RECT 173.800 0.800 174.200 3.100 ;
        RECT 175.400 0.800 175.800 3.100 ;
        RECT 178.200 0.800 178.600 5.000 ;
        RECT 179.800 0.800 180.200 3.100 ;
        RECT 181.400 0.800 181.800 3.100 ;
        RECT 182.500 0.800 182.900 3.100 ;
        RECT 184.600 0.800 185.000 5.100 ;
        RECT 186.200 0.800 186.600 5.000 ;
        RECT 189.000 0.800 189.400 3.100 ;
        RECT 190.600 0.800 191.000 3.100 ;
        RECT 193.400 0.800 193.800 5.100 ;
        RECT 195.000 0.800 195.400 5.100 ;
        RECT 197.100 0.800 197.500 3.100 ;
        RECT 198.200 0.800 198.600 3.100 ;
        RECT 199.800 0.800 200.200 3.100 ;
        RECT 203.000 0.800 203.400 5.000 ;
        RECT 205.800 0.800 206.200 3.100 ;
        RECT 207.400 0.800 207.800 3.100 ;
        RECT 210.200 0.800 210.600 5.100 ;
        RECT 212.600 0.800 213.000 5.000 ;
        RECT 215.400 0.800 215.800 3.100 ;
        RECT 217.000 0.800 217.400 3.100 ;
        RECT 219.800 0.800 220.200 5.100 ;
        RECT 221.400 0.800 221.800 5.100 ;
        RECT 223.500 0.800 223.900 3.100 ;
        RECT 224.600 0.800 225.000 3.100 ;
        RECT 226.200 0.800 226.600 3.100 ;
        RECT 227.800 0.800 228.200 5.100 ;
        RECT 230.600 0.800 231.000 3.100 ;
        RECT 232.200 0.800 232.600 3.100 ;
        RECT 235.000 0.800 235.400 5.000 ;
        RECT 236.600 0.800 237.000 5.100 ;
        RECT 238.200 0.800 238.600 5.100 ;
        RECT 239.800 0.800 240.200 5.100 ;
        RECT 241.400 0.800 241.800 5.100 ;
        RECT 243.000 0.800 243.400 5.100 ;
        RECT 243.800 0.800 244.200 5.100 ;
        RECT 245.400 0.800 245.800 5.100 ;
        RECT 247.000 0.800 247.400 5.100 ;
        RECT 247.800 0.800 248.200 5.100 ;
        RECT 249.400 0.800 249.800 5.100 ;
        RECT 251.000 0.800 251.400 5.100 ;
        RECT 0.200 0.200 252.600 0.800 ;
      LAYER via1 ;
        RECT 48.200 240.300 48.600 240.700 ;
        RECT 48.900 240.300 49.300 240.700 ;
        RECT 149.800 240.300 150.200 240.700 ;
        RECT 150.500 240.300 150.900 240.700 ;
        RECT 48.200 220.300 48.600 220.700 ;
        RECT 48.900 220.300 49.300 220.700 ;
        RECT 149.800 220.300 150.200 220.700 ;
        RECT 150.500 220.300 150.900 220.700 ;
        RECT 48.200 200.300 48.600 200.700 ;
        RECT 48.900 200.300 49.300 200.700 ;
        RECT 149.800 200.300 150.200 200.700 ;
        RECT 150.500 200.300 150.900 200.700 ;
        RECT 48.200 180.300 48.600 180.700 ;
        RECT 48.900 180.300 49.300 180.700 ;
        RECT 149.800 180.300 150.200 180.700 ;
        RECT 150.500 180.300 150.900 180.700 ;
        RECT 48.200 160.300 48.600 160.700 ;
        RECT 48.900 160.300 49.300 160.700 ;
        RECT 149.800 160.300 150.200 160.700 ;
        RECT 150.500 160.300 150.900 160.700 ;
        RECT 48.200 140.300 48.600 140.700 ;
        RECT 48.900 140.300 49.300 140.700 ;
        RECT 149.800 140.300 150.200 140.700 ;
        RECT 150.500 140.300 150.900 140.700 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 149.800 120.300 150.200 120.700 ;
        RECT 150.500 120.300 150.900 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 149.800 100.300 150.200 100.700 ;
        RECT 150.500 100.300 150.900 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 149.800 80.300 150.200 80.700 ;
        RECT 150.500 80.300 150.900 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 149.800 60.300 150.200 60.700 ;
        RECT 150.500 60.300 150.900 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 149.800 40.300 150.200 40.700 ;
        RECT 150.500 40.300 150.900 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 149.800 20.300 150.200 20.700 ;
        RECT 150.500 20.300 150.900 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
        RECT 149.800 0.300 150.200 0.700 ;
        RECT 150.500 0.300 150.900 0.700 ;
      LAYER metal2 ;
        RECT 48.000 240.300 49.600 240.700 ;
        RECT 149.600 240.300 151.200 240.700 ;
        RECT 48.000 220.300 49.600 220.700 ;
        RECT 149.600 220.300 151.200 220.700 ;
        RECT 48.000 200.300 49.600 200.700 ;
        RECT 149.600 200.300 151.200 200.700 ;
        RECT 48.000 180.300 49.600 180.700 ;
        RECT 149.600 180.300 151.200 180.700 ;
        RECT 48.000 160.300 49.600 160.700 ;
        RECT 149.600 160.300 151.200 160.700 ;
        RECT 48.000 140.300 49.600 140.700 ;
        RECT 149.600 140.300 151.200 140.700 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 149.600 120.300 151.200 120.700 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 149.600 100.300 151.200 100.700 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 149.600 80.300 151.200 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 149.600 60.300 151.200 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 149.600 40.300 151.200 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 149.600 20.300 151.200 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
        RECT 149.600 0.300 151.200 0.700 ;
      LAYER via2 ;
        RECT 48.200 240.300 48.600 240.700 ;
        RECT 48.900 240.300 49.300 240.700 ;
        RECT 149.800 240.300 150.200 240.700 ;
        RECT 150.500 240.300 150.900 240.700 ;
        RECT 48.200 220.300 48.600 220.700 ;
        RECT 48.900 220.300 49.300 220.700 ;
        RECT 149.800 220.300 150.200 220.700 ;
        RECT 150.500 220.300 150.900 220.700 ;
        RECT 48.200 200.300 48.600 200.700 ;
        RECT 48.900 200.300 49.300 200.700 ;
        RECT 149.800 200.300 150.200 200.700 ;
        RECT 150.500 200.300 150.900 200.700 ;
        RECT 48.200 180.300 48.600 180.700 ;
        RECT 48.900 180.300 49.300 180.700 ;
        RECT 149.800 180.300 150.200 180.700 ;
        RECT 150.500 180.300 150.900 180.700 ;
        RECT 48.200 160.300 48.600 160.700 ;
        RECT 48.900 160.300 49.300 160.700 ;
        RECT 149.800 160.300 150.200 160.700 ;
        RECT 150.500 160.300 150.900 160.700 ;
        RECT 48.200 140.300 48.600 140.700 ;
        RECT 48.900 140.300 49.300 140.700 ;
        RECT 149.800 140.300 150.200 140.700 ;
        RECT 150.500 140.300 150.900 140.700 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 149.800 120.300 150.200 120.700 ;
        RECT 150.500 120.300 150.900 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 149.800 100.300 150.200 100.700 ;
        RECT 150.500 100.300 150.900 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 149.800 80.300 150.200 80.700 ;
        RECT 150.500 80.300 150.900 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 149.800 60.300 150.200 60.700 ;
        RECT 150.500 60.300 150.900 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 149.800 40.300 150.200 40.700 ;
        RECT 150.500 40.300 150.900 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 149.800 20.300 150.200 20.700 ;
        RECT 150.500 20.300 150.900 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
        RECT 149.800 0.300 150.200 0.700 ;
        RECT 150.500 0.300 150.900 0.700 ;
      LAYER metal3 ;
        RECT 48.000 240.300 49.600 240.700 ;
        RECT 149.600 240.300 151.200 240.700 ;
        RECT 48.000 220.300 49.600 220.700 ;
        RECT 149.600 220.300 151.200 220.700 ;
        RECT 48.000 200.300 49.600 200.700 ;
        RECT 149.600 200.300 151.200 200.700 ;
        RECT 48.000 180.300 49.600 180.700 ;
        RECT 149.600 180.300 151.200 180.700 ;
        RECT 48.000 160.300 49.600 160.700 ;
        RECT 149.600 160.300 151.200 160.700 ;
        RECT 48.000 140.300 49.600 140.700 ;
        RECT 149.600 140.300 151.200 140.700 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 149.600 120.300 151.200 120.700 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 149.600 100.300 151.200 100.700 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 149.600 80.300 151.200 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 149.600 60.300 151.200 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 149.600 40.300 151.200 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 149.600 20.300 151.200 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
        RECT 149.600 0.300 151.200 0.700 ;
      LAYER via3 ;
        RECT 48.200 240.300 48.600 240.700 ;
        RECT 49.000 240.300 49.400 240.700 ;
        RECT 149.800 240.300 150.200 240.700 ;
        RECT 150.600 240.300 151.000 240.700 ;
        RECT 48.200 220.300 48.600 220.700 ;
        RECT 49.000 220.300 49.400 220.700 ;
        RECT 149.800 220.300 150.200 220.700 ;
        RECT 150.600 220.300 151.000 220.700 ;
        RECT 48.200 200.300 48.600 200.700 ;
        RECT 49.000 200.300 49.400 200.700 ;
        RECT 149.800 200.300 150.200 200.700 ;
        RECT 150.600 200.300 151.000 200.700 ;
        RECT 48.200 180.300 48.600 180.700 ;
        RECT 49.000 180.300 49.400 180.700 ;
        RECT 149.800 180.300 150.200 180.700 ;
        RECT 150.600 180.300 151.000 180.700 ;
        RECT 48.200 160.300 48.600 160.700 ;
        RECT 49.000 160.300 49.400 160.700 ;
        RECT 149.800 160.300 150.200 160.700 ;
        RECT 150.600 160.300 151.000 160.700 ;
        RECT 48.200 140.300 48.600 140.700 ;
        RECT 49.000 140.300 49.400 140.700 ;
        RECT 149.800 140.300 150.200 140.700 ;
        RECT 150.600 140.300 151.000 140.700 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 49.000 120.300 49.400 120.700 ;
        RECT 149.800 120.300 150.200 120.700 ;
        RECT 150.600 120.300 151.000 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 49.000 100.300 49.400 100.700 ;
        RECT 149.800 100.300 150.200 100.700 ;
        RECT 150.600 100.300 151.000 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 49.000 80.300 49.400 80.700 ;
        RECT 149.800 80.300 150.200 80.700 ;
        RECT 150.600 80.300 151.000 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 49.000 60.300 49.400 60.700 ;
        RECT 149.800 60.300 150.200 60.700 ;
        RECT 150.600 60.300 151.000 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 49.000 40.300 49.400 40.700 ;
        RECT 149.800 40.300 150.200 40.700 ;
        RECT 150.600 40.300 151.000 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 49.000 20.300 49.400 20.700 ;
        RECT 149.800 20.300 150.200 20.700 ;
        RECT 150.600 20.300 151.000 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 49.000 0.300 49.400 0.700 ;
        RECT 149.800 0.300 150.200 0.700 ;
        RECT 150.600 0.300 151.000 0.700 ;
      LAYER metal4 ;
        RECT 48.000 240.300 49.600 240.700 ;
        RECT 149.600 240.300 151.200 240.700 ;
        RECT 48.000 220.300 49.600 220.700 ;
        RECT 149.600 220.300 151.200 220.700 ;
        RECT 48.000 200.300 49.600 200.700 ;
        RECT 149.600 200.300 151.200 200.700 ;
        RECT 48.000 180.300 49.600 180.700 ;
        RECT 149.600 180.300 151.200 180.700 ;
        RECT 48.000 160.300 49.600 160.700 ;
        RECT 149.600 160.300 151.200 160.700 ;
        RECT 48.000 140.300 49.600 140.700 ;
        RECT 149.600 140.300 151.200 140.700 ;
        RECT 48.000 120.300 49.600 120.700 ;
        RECT 149.600 120.300 151.200 120.700 ;
        RECT 48.000 100.300 49.600 100.700 ;
        RECT 149.600 100.300 151.200 100.700 ;
        RECT 48.000 80.300 49.600 80.700 ;
        RECT 149.600 80.300 151.200 80.700 ;
        RECT 48.000 60.300 49.600 60.700 ;
        RECT 149.600 60.300 151.200 60.700 ;
        RECT 48.000 40.300 49.600 40.700 ;
        RECT 149.600 40.300 151.200 40.700 ;
        RECT 48.000 20.300 49.600 20.700 ;
        RECT 149.600 20.300 151.200 20.700 ;
        RECT 48.000 0.300 49.600 0.700 ;
        RECT 149.600 0.300 151.200 0.700 ;
      LAYER via4 ;
        RECT 48.200 240.300 48.600 240.700 ;
        RECT 48.900 240.300 49.300 240.700 ;
        RECT 149.800 240.300 150.200 240.700 ;
        RECT 150.500 240.300 150.900 240.700 ;
        RECT 48.200 220.300 48.600 220.700 ;
        RECT 48.900 220.300 49.300 220.700 ;
        RECT 149.800 220.300 150.200 220.700 ;
        RECT 150.500 220.300 150.900 220.700 ;
        RECT 48.200 200.300 48.600 200.700 ;
        RECT 48.900 200.300 49.300 200.700 ;
        RECT 149.800 200.300 150.200 200.700 ;
        RECT 150.500 200.300 150.900 200.700 ;
        RECT 48.200 180.300 48.600 180.700 ;
        RECT 48.900 180.300 49.300 180.700 ;
        RECT 149.800 180.300 150.200 180.700 ;
        RECT 150.500 180.300 150.900 180.700 ;
        RECT 48.200 160.300 48.600 160.700 ;
        RECT 48.900 160.300 49.300 160.700 ;
        RECT 149.800 160.300 150.200 160.700 ;
        RECT 150.500 160.300 150.900 160.700 ;
        RECT 48.200 140.300 48.600 140.700 ;
        RECT 48.900 140.300 49.300 140.700 ;
        RECT 149.800 140.300 150.200 140.700 ;
        RECT 150.500 140.300 150.900 140.700 ;
        RECT 48.200 120.300 48.600 120.700 ;
        RECT 48.900 120.300 49.300 120.700 ;
        RECT 149.800 120.300 150.200 120.700 ;
        RECT 150.500 120.300 150.900 120.700 ;
        RECT 48.200 100.300 48.600 100.700 ;
        RECT 48.900 100.300 49.300 100.700 ;
        RECT 149.800 100.300 150.200 100.700 ;
        RECT 150.500 100.300 150.900 100.700 ;
        RECT 48.200 80.300 48.600 80.700 ;
        RECT 48.900 80.300 49.300 80.700 ;
        RECT 149.800 80.300 150.200 80.700 ;
        RECT 150.500 80.300 150.900 80.700 ;
        RECT 48.200 60.300 48.600 60.700 ;
        RECT 48.900 60.300 49.300 60.700 ;
        RECT 149.800 60.300 150.200 60.700 ;
        RECT 150.500 60.300 150.900 60.700 ;
        RECT 48.200 40.300 48.600 40.700 ;
        RECT 48.900 40.300 49.300 40.700 ;
        RECT 149.800 40.300 150.200 40.700 ;
        RECT 150.500 40.300 150.900 40.700 ;
        RECT 48.200 20.300 48.600 20.700 ;
        RECT 48.900 20.300 49.300 20.700 ;
        RECT 149.800 20.300 150.200 20.700 ;
        RECT 150.500 20.300 150.900 20.700 ;
        RECT 48.200 0.300 48.600 0.700 ;
        RECT 48.900 0.300 49.300 0.700 ;
        RECT 149.800 0.300 150.200 0.700 ;
        RECT 150.500 0.300 150.900 0.700 ;
      LAYER metal5 ;
        RECT 48.000 240.200 49.600 240.700 ;
        RECT 149.600 240.200 151.200 240.700 ;
        RECT 48.000 220.200 49.600 220.700 ;
        RECT 149.600 220.200 151.200 220.700 ;
        RECT 48.000 200.200 49.600 200.700 ;
        RECT 149.600 200.200 151.200 200.700 ;
        RECT 48.000 180.200 49.600 180.700 ;
        RECT 149.600 180.200 151.200 180.700 ;
        RECT 48.000 160.200 49.600 160.700 ;
        RECT 149.600 160.200 151.200 160.700 ;
        RECT 48.000 140.200 49.600 140.700 ;
        RECT 149.600 140.200 151.200 140.700 ;
        RECT 48.000 120.200 49.600 120.700 ;
        RECT 149.600 120.200 151.200 120.700 ;
        RECT 48.000 100.200 49.600 100.700 ;
        RECT 149.600 100.200 151.200 100.700 ;
        RECT 48.000 80.200 49.600 80.700 ;
        RECT 149.600 80.200 151.200 80.700 ;
        RECT 48.000 60.200 49.600 60.700 ;
        RECT 149.600 60.200 151.200 60.700 ;
        RECT 48.000 40.200 49.600 40.700 ;
        RECT 149.600 40.200 151.200 40.700 ;
        RECT 48.000 20.200 49.600 20.700 ;
        RECT 149.600 20.200 151.200 20.700 ;
        RECT 48.000 0.200 49.600 0.700 ;
        RECT 149.600 0.200 151.200 0.700 ;
      LAYER via5 ;
        RECT 49.000 240.200 49.500 240.700 ;
        RECT 150.600 240.200 151.100 240.700 ;
        RECT 49.000 220.200 49.500 220.700 ;
        RECT 150.600 220.200 151.100 220.700 ;
        RECT 49.000 200.200 49.500 200.700 ;
        RECT 150.600 200.200 151.100 200.700 ;
        RECT 49.000 180.200 49.500 180.700 ;
        RECT 150.600 180.200 151.100 180.700 ;
        RECT 49.000 160.200 49.500 160.700 ;
        RECT 150.600 160.200 151.100 160.700 ;
        RECT 49.000 140.200 49.500 140.700 ;
        RECT 150.600 140.200 151.100 140.700 ;
        RECT 49.000 120.200 49.500 120.700 ;
        RECT 150.600 120.200 151.100 120.700 ;
        RECT 49.000 100.200 49.500 100.700 ;
        RECT 150.600 100.200 151.100 100.700 ;
        RECT 49.000 80.200 49.500 80.700 ;
        RECT 150.600 80.200 151.100 80.700 ;
        RECT 49.000 60.200 49.500 60.700 ;
        RECT 150.600 60.200 151.100 60.700 ;
        RECT 49.000 40.200 49.500 40.700 ;
        RECT 150.600 40.200 151.100 40.700 ;
        RECT 49.000 20.200 49.500 20.700 ;
        RECT 150.600 20.200 151.100 20.700 ;
        RECT 49.000 0.200 49.500 0.700 ;
        RECT 150.600 0.200 151.100 0.700 ;
      LAYER metal6 ;
        RECT 48.000 -3.000 49.600 243.000 ;
        RECT 149.600 -3.000 151.200 243.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 230.800 1.000 232.100 ;
        RECT 2.200 230.800 2.600 232.100 ;
        RECT 3.000 230.800 3.400 232.100 ;
        RECT 5.100 230.800 5.500 233.100 ;
        RECT 7.000 230.800 7.400 232.700 ;
        RECT 11.000 230.800 11.400 233.100 ;
        RECT 12.600 230.800 13.000 233.000 ;
        RECT 15.400 230.800 15.800 232.100 ;
        RECT 17.000 230.800 17.500 232.100 ;
        RECT 19.800 230.800 20.200 233.100 ;
        RECT 21.400 230.800 21.800 233.100 ;
        RECT 23.000 230.800 23.400 233.100 ;
        RECT 24.600 230.800 25.000 233.100 ;
        RECT 26.200 230.800 26.600 233.100 ;
        RECT 27.800 230.800 28.200 233.100 ;
        RECT 29.400 230.800 29.800 232.700 ;
        RECT 33.400 230.800 33.800 233.100 ;
        RECT 35.000 230.800 35.400 233.100 ;
        RECT 37.700 230.800 38.200 232.100 ;
        RECT 39.400 230.800 39.800 232.100 ;
        RECT 42.200 230.800 42.600 233.000 ;
        RECT 46.200 230.800 46.600 233.000 ;
        RECT 49.000 230.800 49.400 232.100 ;
        RECT 50.600 230.800 51.100 232.100 ;
        RECT 53.400 230.800 53.800 233.100 ;
        RECT 55.000 230.800 55.400 233.100 ;
        RECT 59.000 230.800 59.400 232.700 ;
        RECT 61.400 230.800 61.800 233.100 ;
        RECT 64.100 230.800 64.600 232.100 ;
        RECT 65.800 230.800 66.200 232.100 ;
        RECT 68.600 230.800 69.000 233.000 ;
        RECT 70.200 230.800 70.600 233.100 ;
        RECT 74.200 230.800 74.600 232.700 ;
        RECT 76.600 230.800 77.000 233.000 ;
        RECT 79.400 230.800 79.800 232.100 ;
        RECT 81.000 230.800 81.500 232.100 ;
        RECT 83.800 230.800 84.200 233.100 ;
        RECT 86.200 230.800 86.600 233.100 ;
        RECT 87.800 230.800 88.200 233.100 ;
        RECT 89.400 230.800 89.800 233.100 ;
        RECT 91.000 230.800 91.400 233.100 ;
        RECT 92.600 230.800 93.000 233.100 ;
        RECT 94.200 230.800 94.600 233.100 ;
        RECT 95.800 230.800 96.200 233.100 ;
        RECT 97.400 230.800 97.800 233.100 ;
        RECT 100.600 230.800 101.000 233.100 ;
        RECT 103.300 230.800 103.800 232.100 ;
        RECT 105.000 230.800 105.400 232.100 ;
        RECT 107.800 230.800 108.200 233.000 ;
        RECT 110.200 230.800 110.600 232.700 ;
        RECT 112.600 230.800 113.000 233.100 ;
        RECT 114.200 230.800 114.600 233.100 ;
        RECT 115.800 230.800 116.200 233.100 ;
        RECT 117.400 230.800 117.800 233.100 ;
        RECT 120.100 230.800 120.600 232.100 ;
        RECT 121.800 230.800 122.200 232.100 ;
        RECT 124.600 230.800 125.000 233.000 ;
        RECT 126.200 230.800 126.600 233.100 ;
        RECT 130.200 230.800 130.600 232.700 ;
        RECT 132.600 230.800 133.000 232.700 ;
        RECT 136.600 230.800 137.000 233.100 ;
        RECT 138.200 230.800 138.600 233.100 ;
        RECT 140.900 230.800 141.400 232.100 ;
        RECT 142.600 230.800 143.000 232.100 ;
        RECT 145.400 230.800 145.800 233.000 ;
        RECT 147.300 230.800 147.700 233.100 ;
        RECT 149.400 230.800 149.800 232.100 ;
        RECT 151.800 230.800 152.200 232.100 ;
        RECT 153.400 230.800 153.800 232.100 ;
        RECT 155.000 230.800 155.400 233.100 ;
        RECT 157.400 230.800 157.800 232.700 ;
        RECT 161.400 230.800 161.800 233.100 ;
        RECT 163.000 230.800 163.400 233.000 ;
        RECT 165.800 230.800 166.200 232.100 ;
        RECT 167.400 230.800 167.900 232.100 ;
        RECT 170.200 230.800 170.600 233.100 ;
        RECT 172.600 230.800 173.000 233.000 ;
        RECT 175.400 230.800 175.800 232.100 ;
        RECT 177.000 230.800 177.500 232.100 ;
        RECT 179.800 230.800 180.200 233.100 ;
        RECT 182.200 230.800 182.600 233.100 ;
        RECT 184.900 230.800 185.400 232.100 ;
        RECT 186.600 230.800 187.000 232.100 ;
        RECT 189.400 230.800 189.800 233.000 ;
        RECT 191.800 230.800 192.200 232.700 ;
        RECT 195.000 230.800 195.400 233.100 ;
        RECT 197.700 230.800 198.200 232.100 ;
        RECT 199.400 230.800 199.800 232.100 ;
        RECT 202.200 230.800 202.600 233.000 ;
        RECT 205.400 230.800 205.800 233.100 ;
        RECT 209.400 230.800 209.800 232.700 ;
        RECT 211.800 230.800 212.200 233.100 ;
        RECT 214.500 230.800 215.000 232.100 ;
        RECT 216.200 230.800 216.600 232.100 ;
        RECT 219.000 230.800 219.400 233.000 ;
        RECT 222.200 230.800 222.600 233.100 ;
        RECT 223.800 230.800 224.200 233.100 ;
        RECT 226.500 230.800 227.000 232.100 ;
        RECT 228.200 230.800 228.600 232.100 ;
        RECT 231.000 230.800 231.400 233.000 ;
        RECT 233.400 230.800 233.800 233.100 ;
        RECT 236.100 230.800 236.600 232.100 ;
        RECT 237.800 230.800 238.200 232.100 ;
        RECT 240.600 230.800 241.000 233.000 ;
        RECT 242.200 230.800 242.600 233.100 ;
        RECT 243.800 230.800 244.200 233.100 ;
        RECT 245.400 230.800 245.800 233.100 ;
        RECT 247.000 230.800 247.400 232.700 ;
        RECT 251.000 230.800 251.400 233.100 ;
        RECT 0.200 230.200 252.600 230.800 ;
        RECT 1.400 228.000 1.800 230.200 ;
        RECT 4.200 228.900 4.600 230.200 ;
        RECT 5.800 228.900 6.300 230.200 ;
        RECT 8.600 227.900 9.000 230.200 ;
        RECT 10.200 227.900 10.600 230.200 ;
        RECT 11.800 227.900 12.200 230.200 ;
        RECT 13.400 227.900 13.800 230.200 ;
        RECT 15.000 227.900 15.400 230.200 ;
        RECT 16.600 227.900 17.000 230.200 ;
        RECT 18.200 228.300 18.600 230.200 ;
        RECT 22.200 227.900 22.600 230.200 ;
        RECT 23.800 227.900 24.200 230.200 ;
        RECT 26.500 228.900 27.000 230.200 ;
        RECT 28.200 228.900 28.600 230.200 ;
        RECT 31.000 228.000 31.400 230.200 ;
        RECT 33.400 227.700 33.800 230.200 ;
        RECT 36.000 227.500 36.400 230.200 ;
        RECT 38.200 228.300 38.600 230.200 ;
        RECT 42.200 227.900 42.600 230.200 ;
        RECT 43.800 227.900 44.200 230.200 ;
        RECT 46.500 228.900 47.000 230.200 ;
        RECT 48.200 228.900 48.600 230.200 ;
        RECT 51.000 228.000 51.400 230.200 ;
        RECT 55.000 227.700 55.400 230.200 ;
        RECT 57.600 227.500 58.000 230.200 ;
        RECT 59.800 227.700 60.200 230.200 ;
        RECT 62.400 227.500 62.800 230.200 ;
        RECT 64.600 227.700 65.000 230.200 ;
        RECT 67.200 227.500 67.600 230.200 ;
        RECT 68.600 227.900 69.000 230.200 ;
        RECT 70.200 227.900 70.600 230.200 ;
        RECT 71.800 227.900 72.200 230.200 ;
        RECT 73.400 227.900 73.800 230.200 ;
        RECT 75.000 227.900 75.400 230.200 ;
        RECT 76.600 228.000 77.000 230.200 ;
        RECT 79.400 228.900 79.800 230.200 ;
        RECT 81.000 228.900 81.500 230.200 ;
        RECT 83.800 227.900 84.200 230.200 ;
        RECT 85.400 227.900 85.800 230.200 ;
        RECT 89.400 228.300 89.800 230.200 ;
        RECT 91.600 227.500 92.000 230.200 ;
        RECT 94.200 227.700 94.600 230.200 ;
        RECT 98.200 228.000 98.600 230.200 ;
        RECT 101.000 228.900 101.400 230.200 ;
        RECT 102.600 228.900 103.100 230.200 ;
        RECT 105.400 227.900 105.800 230.200 ;
        RECT 107.800 228.300 108.200 230.200 ;
        RECT 110.200 227.900 110.600 230.200 ;
        RECT 114.200 228.300 114.600 230.200 ;
        RECT 115.800 228.900 116.200 230.200 ;
        RECT 117.400 228.900 117.800 230.200 ;
        RECT 118.200 228.900 118.600 230.200 ;
        RECT 120.300 227.900 120.700 230.200 ;
        RECT 123.000 227.900 123.400 230.200 ;
        RECT 124.400 227.500 124.800 230.200 ;
        RECT 127.000 227.700 127.400 230.200 ;
        RECT 129.400 228.000 129.800 230.200 ;
        RECT 132.200 228.900 132.600 230.200 ;
        RECT 133.800 228.900 134.300 230.200 ;
        RECT 136.600 227.900 137.000 230.200 ;
        RECT 139.000 228.300 139.400 230.200 ;
        RECT 141.400 227.900 141.800 230.200 ;
        RECT 144.400 227.500 144.800 230.200 ;
        RECT 147.000 227.700 147.400 230.200 ;
        RECT 151.000 228.000 151.400 230.200 ;
        RECT 153.800 228.900 154.200 230.200 ;
        RECT 155.400 228.900 155.900 230.200 ;
        RECT 158.200 227.900 158.600 230.200 ;
        RECT 160.100 227.900 160.500 230.200 ;
        RECT 162.200 228.900 162.600 230.200 ;
        RECT 163.000 228.900 163.400 230.200 ;
        RECT 164.600 228.900 165.000 230.200 ;
        RECT 165.400 227.900 165.800 230.200 ;
        RECT 167.000 227.900 167.400 230.200 ;
        RECT 168.600 227.900 169.000 230.200 ;
        RECT 170.200 227.900 170.600 230.200 ;
        RECT 171.800 227.900 172.200 230.200 ;
        RECT 173.400 227.900 173.800 230.200 ;
        RECT 176.100 228.900 176.600 230.200 ;
        RECT 177.800 228.900 178.200 230.200 ;
        RECT 180.600 228.000 181.000 230.200 ;
        RECT 183.000 227.700 183.400 230.200 ;
        RECT 185.600 227.500 186.000 230.200 ;
        RECT 187.600 227.500 188.000 230.200 ;
        RECT 190.200 227.700 190.600 230.200 ;
        RECT 192.600 227.700 193.000 230.200 ;
        RECT 195.200 227.500 195.600 230.200 ;
        RECT 197.400 228.300 197.800 230.200 ;
        RECT 201.400 227.900 201.800 230.200 ;
        RECT 203.800 227.900 204.200 230.200 ;
        RECT 207.000 227.900 207.400 230.200 ;
        RECT 209.700 228.900 210.200 230.200 ;
        RECT 211.400 228.900 211.800 230.200 ;
        RECT 214.200 228.000 214.600 230.200 ;
        RECT 216.600 227.700 217.000 230.200 ;
        RECT 219.200 227.500 219.600 230.200 ;
        RECT 221.200 227.500 221.600 230.200 ;
        RECT 223.800 227.700 224.200 230.200 ;
        RECT 226.200 228.300 226.600 230.200 ;
        RECT 230.200 227.900 230.600 230.200 ;
        RECT 231.800 228.000 232.200 230.200 ;
        RECT 234.600 228.900 235.000 230.200 ;
        RECT 236.200 228.900 236.700 230.200 ;
        RECT 239.000 227.900 239.400 230.200 ;
        RECT 241.400 228.000 241.800 230.200 ;
        RECT 244.200 228.900 244.600 230.200 ;
        RECT 245.800 228.900 246.300 230.200 ;
        RECT 248.600 227.900 249.000 230.200 ;
        RECT 1.400 210.800 1.800 213.000 ;
        RECT 4.200 210.800 4.600 212.100 ;
        RECT 5.800 210.800 6.300 212.100 ;
        RECT 8.600 210.800 9.000 213.100 ;
        RECT 11.000 210.800 11.400 212.700 ;
        RECT 15.000 210.800 15.400 213.100 ;
        RECT 16.600 210.800 17.000 213.100 ;
        RECT 19.300 210.800 19.800 212.100 ;
        RECT 21.000 210.800 21.400 212.100 ;
        RECT 23.800 210.800 24.200 213.000 ;
        RECT 26.000 210.800 26.400 213.500 ;
        RECT 28.600 210.800 29.000 213.300 ;
        RECT 30.200 210.800 30.600 212.100 ;
        RECT 31.800 210.800 32.200 212.100 ;
        RECT 32.600 210.800 33.000 212.100 ;
        RECT 34.700 210.800 35.100 213.100 ;
        RECT 36.600 210.800 37.000 213.000 ;
        RECT 39.400 210.800 39.800 212.100 ;
        RECT 41.000 210.800 41.500 212.100 ;
        RECT 43.800 210.800 44.200 213.100 ;
        RECT 46.200 210.800 46.600 213.100 ;
        RECT 50.200 210.800 50.600 213.000 ;
        RECT 53.000 210.800 53.400 212.100 ;
        RECT 54.600 210.800 55.100 212.100 ;
        RECT 57.400 210.800 57.800 213.100 ;
        RECT 59.800 210.800 60.200 213.000 ;
        RECT 62.600 210.800 63.000 212.100 ;
        RECT 64.200 210.800 64.700 212.100 ;
        RECT 67.000 210.800 67.400 213.100 ;
        RECT 70.200 210.800 70.600 212.700 ;
        RECT 72.100 210.800 72.500 213.100 ;
        RECT 74.200 210.800 74.600 212.100 ;
        RECT 75.800 210.800 76.200 213.100 ;
        RECT 77.400 210.800 77.800 213.100 ;
        RECT 78.200 210.800 78.600 213.100 ;
        RECT 79.800 210.800 80.200 213.100 ;
        RECT 82.200 210.800 82.600 213.100 ;
        RECT 84.900 210.800 85.400 212.100 ;
        RECT 86.600 210.800 87.000 212.100 ;
        RECT 89.400 210.800 89.800 213.000 ;
        RECT 91.800 210.800 92.200 212.700 ;
        RECT 94.200 210.800 94.600 213.100 ;
        RECT 97.200 210.800 97.600 213.500 ;
        RECT 99.800 210.800 100.200 213.300 ;
        RECT 104.600 210.800 105.000 212.700 ;
        RECT 106.200 210.800 106.600 213.100 ;
        RECT 109.400 210.800 109.800 213.000 ;
        RECT 112.200 210.800 112.600 212.100 ;
        RECT 113.800 210.800 114.300 212.100 ;
        RECT 116.600 210.800 117.000 213.100 ;
        RECT 118.200 210.800 118.600 213.100 ;
        RECT 121.400 210.800 121.800 213.000 ;
        RECT 124.200 210.800 124.600 212.100 ;
        RECT 125.800 210.800 126.300 212.100 ;
        RECT 128.600 210.800 129.000 213.100 ;
        RECT 131.000 210.800 131.400 212.700 ;
        RECT 135.000 210.800 135.400 213.100 ;
        RECT 136.600 210.800 137.000 213.100 ;
        RECT 139.300 210.800 139.800 212.100 ;
        RECT 141.000 210.800 141.400 212.100 ;
        RECT 143.800 210.800 144.200 213.000 ;
        RECT 146.200 210.800 146.600 213.000 ;
        RECT 149.000 210.800 149.400 212.100 ;
        RECT 150.600 210.800 151.100 212.100 ;
        RECT 153.400 210.800 153.800 213.100 ;
        RECT 157.400 210.800 157.800 212.700 ;
        RECT 161.400 210.800 161.800 213.100 ;
        RECT 163.000 210.800 163.400 212.700 ;
        RECT 167.000 210.800 167.400 213.100 ;
        RECT 168.600 210.800 169.000 213.100 ;
        RECT 171.300 210.800 171.800 212.100 ;
        RECT 173.000 210.800 173.400 212.100 ;
        RECT 175.800 210.800 176.200 213.000 ;
        RECT 177.400 210.800 177.800 213.100 ;
        RECT 179.000 210.800 179.400 213.100 ;
        RECT 180.600 210.800 181.000 213.100 ;
        RECT 183.800 210.800 184.200 213.000 ;
        RECT 186.600 210.800 187.000 212.100 ;
        RECT 188.200 210.800 188.700 212.100 ;
        RECT 191.000 210.800 191.400 213.100 ;
        RECT 192.600 210.800 193.000 213.100 ;
        RECT 194.200 210.800 194.600 213.100 ;
        RECT 195.800 210.800 196.200 213.100 ;
        RECT 197.400 210.800 197.800 213.100 ;
        RECT 199.000 210.800 199.400 213.100 ;
        RECT 200.600 210.800 201.000 213.100 ;
        RECT 202.200 210.800 202.600 213.100 ;
        RECT 205.400 210.800 205.800 212.700 ;
        RECT 209.400 210.800 209.800 213.100 ;
        RECT 210.200 210.800 210.600 213.100 ;
        RECT 211.800 210.800 212.200 213.100 ;
        RECT 213.400 210.800 213.800 213.100 ;
        RECT 215.000 210.800 215.400 213.100 ;
        RECT 216.600 210.800 217.000 213.100 ;
        RECT 219.000 210.800 219.400 213.100 ;
        RECT 221.400 210.800 221.800 212.700 ;
        RECT 223.800 210.800 224.200 213.100 ;
        RECT 226.500 210.800 227.000 212.100 ;
        RECT 228.200 210.800 228.600 212.100 ;
        RECT 231.000 210.800 231.400 213.000 ;
        RECT 234.200 210.800 234.600 212.700 ;
        RECT 235.800 210.800 236.200 213.100 ;
        RECT 239.800 210.800 240.200 212.700 ;
        RECT 242.200 210.800 242.600 213.000 ;
        RECT 245.000 210.800 245.400 212.100 ;
        RECT 246.600 210.800 247.100 212.100 ;
        RECT 249.400 210.800 249.800 213.100 ;
        RECT 0.200 210.200 252.600 210.800 ;
        RECT 1.400 208.000 1.800 210.200 ;
        RECT 4.200 208.900 4.600 210.200 ;
        RECT 5.800 208.900 6.300 210.200 ;
        RECT 8.600 207.900 9.000 210.200 ;
        RECT 11.000 208.300 11.400 210.200 ;
        RECT 15.000 207.900 15.400 210.200 ;
        RECT 16.600 208.300 17.000 210.200 ;
        RECT 20.600 207.900 21.000 210.200 ;
        RECT 22.200 207.700 22.600 210.200 ;
        RECT 24.800 207.500 25.200 210.200 ;
        RECT 27.000 208.000 27.400 210.200 ;
        RECT 29.800 208.900 30.200 210.200 ;
        RECT 31.400 208.900 31.900 210.200 ;
        RECT 34.200 207.900 34.600 210.200 ;
        RECT 35.800 207.900 36.200 210.200 ;
        RECT 39.800 208.300 40.200 210.200 ;
        RECT 42.200 207.900 42.600 210.200 ;
        RECT 44.900 208.900 45.400 210.200 ;
        RECT 46.600 208.900 47.000 210.200 ;
        RECT 49.400 208.000 49.800 210.200 ;
        RECT 54.200 207.900 54.600 210.200 ;
        RECT 55.300 207.900 55.700 210.200 ;
        RECT 57.400 208.900 57.800 210.200 ;
        RECT 58.800 207.500 59.200 210.200 ;
        RECT 61.400 207.700 61.800 210.200 ;
        RECT 63.000 207.900 63.400 210.200 ;
        RECT 66.200 208.000 66.600 210.200 ;
        RECT 69.000 208.900 69.400 210.200 ;
        RECT 70.600 208.900 71.100 210.200 ;
        RECT 73.400 207.900 73.800 210.200 ;
        RECT 75.000 208.900 75.400 210.200 ;
        RECT 76.600 208.900 77.000 210.200 ;
        RECT 77.400 207.900 77.800 210.200 ;
        RECT 80.600 207.900 81.000 210.200 ;
        RECT 83.300 208.900 83.800 210.200 ;
        RECT 85.000 208.900 85.400 210.200 ;
        RECT 87.800 208.000 88.200 210.200 ;
        RECT 90.200 207.700 90.600 210.200 ;
        RECT 92.800 207.500 93.200 210.200 ;
        RECT 94.800 207.500 95.200 210.200 ;
        RECT 97.400 207.700 97.800 210.200 ;
        RECT 100.600 207.900 101.000 210.200 ;
        RECT 103.800 208.000 104.200 210.200 ;
        RECT 106.600 208.900 107.000 210.200 ;
        RECT 108.200 208.900 108.700 210.200 ;
        RECT 111.000 207.900 111.400 210.200 ;
        RECT 113.400 207.700 113.800 210.200 ;
        RECT 116.000 207.500 116.400 210.200 ;
        RECT 118.200 207.900 118.600 210.200 ;
        RECT 119.800 207.900 120.200 210.200 ;
        RECT 120.900 207.900 121.300 210.200 ;
        RECT 123.000 208.900 123.400 210.200 ;
        RECT 124.600 207.700 125.000 210.200 ;
        RECT 127.200 207.500 127.600 210.200 ;
        RECT 129.400 208.000 129.800 210.200 ;
        RECT 132.200 208.900 132.600 210.200 ;
        RECT 133.800 208.900 134.300 210.200 ;
        RECT 136.600 207.900 137.000 210.200 ;
        RECT 138.200 208.900 138.600 210.200 ;
        RECT 139.800 208.900 140.200 210.200 ;
        RECT 140.600 208.900 141.000 210.200 ;
        RECT 142.700 207.900 143.100 210.200 ;
        RECT 143.800 208.900 144.200 210.200 ;
        RECT 145.400 208.900 145.800 210.200 ;
        RECT 146.200 208.900 146.600 210.200 ;
        RECT 148.300 207.900 148.700 210.200 ;
        RECT 151.800 207.900 152.200 210.200 ;
        RECT 154.500 208.900 155.000 210.200 ;
        RECT 156.200 208.900 156.600 210.200 ;
        RECT 159.000 208.000 159.400 210.200 ;
        RECT 161.400 207.700 161.800 210.200 ;
        RECT 164.000 207.500 164.400 210.200 ;
        RECT 166.200 208.300 166.600 210.200 ;
        RECT 170.200 207.900 170.600 210.200 ;
        RECT 171.800 207.900 172.200 210.200 ;
        RECT 174.500 208.900 175.000 210.200 ;
        RECT 176.200 208.900 176.600 210.200 ;
        RECT 179.000 208.000 179.400 210.200 ;
        RECT 180.600 208.900 181.000 210.200 ;
        RECT 182.700 207.900 183.100 210.200 ;
        RECT 184.400 207.500 184.800 210.200 ;
        RECT 187.000 207.700 187.400 210.200 ;
        RECT 189.200 207.500 189.600 210.200 ;
        RECT 191.800 207.700 192.200 210.200 ;
        RECT 193.400 208.900 193.800 210.200 ;
        RECT 195.000 208.900 195.400 210.200 ;
        RECT 195.800 208.900 196.200 210.200 ;
        RECT 197.900 207.900 198.300 210.200 ;
        RECT 199.800 208.300 200.200 210.200 ;
        RECT 204.600 208.000 205.000 210.200 ;
        RECT 207.400 208.900 207.800 210.200 ;
        RECT 209.000 208.900 209.500 210.200 ;
        RECT 211.800 207.900 212.200 210.200 ;
        RECT 213.400 207.900 213.800 210.200 ;
        RECT 215.000 207.900 215.400 210.200 ;
        RECT 216.600 207.900 217.000 210.200 ;
        RECT 218.200 207.900 218.600 210.200 ;
        RECT 219.800 207.900 220.200 210.200 ;
        RECT 221.200 207.500 221.600 210.200 ;
        RECT 223.800 207.700 224.200 210.200 ;
        RECT 226.200 207.700 226.600 210.200 ;
        RECT 228.800 207.500 229.200 210.200 ;
        RECT 230.200 207.900 230.600 210.200 ;
        RECT 233.400 208.000 233.800 210.200 ;
        RECT 236.200 208.900 236.600 210.200 ;
        RECT 237.800 208.900 238.300 210.200 ;
        RECT 240.600 207.900 241.000 210.200 ;
        RECT 242.200 207.900 242.600 210.200 ;
        RECT 244.600 208.900 245.000 210.200 ;
        RECT 246.200 208.900 246.600 210.200 ;
        RECT 247.300 207.900 247.700 210.200 ;
        RECT 249.400 208.900 249.800 210.200 ;
        RECT 1.400 190.800 1.800 193.000 ;
        RECT 4.200 190.800 4.600 192.100 ;
        RECT 5.800 190.800 6.300 192.100 ;
        RECT 8.600 190.800 9.000 193.100 ;
        RECT 11.000 190.800 11.400 193.100 ;
        RECT 13.700 190.800 14.200 192.100 ;
        RECT 15.400 190.800 15.800 192.100 ;
        RECT 18.200 190.800 18.600 193.000 ;
        RECT 19.800 190.800 20.200 193.100 ;
        RECT 21.400 190.800 21.800 193.100 ;
        RECT 23.000 190.800 23.400 193.100 ;
        RECT 24.600 190.800 25.000 193.100 ;
        RECT 26.200 190.800 26.600 193.100 ;
        RECT 27.000 190.800 27.400 193.100 ;
        RECT 31.000 190.800 31.400 192.700 ;
        RECT 33.400 190.800 33.800 193.100 ;
        RECT 36.100 190.800 36.600 192.100 ;
        RECT 37.800 190.800 38.200 192.100 ;
        RECT 40.600 190.800 41.000 193.000 ;
        RECT 42.200 190.800 42.600 193.100 ;
        RECT 43.800 190.800 44.200 193.100 ;
        RECT 46.200 190.800 46.600 193.300 ;
        RECT 48.800 190.800 49.200 193.500 ;
        RECT 52.600 190.800 53.000 193.300 ;
        RECT 55.200 190.800 55.600 193.500 ;
        RECT 56.600 190.800 57.000 193.100 ;
        RECT 60.600 190.800 61.000 192.700 ;
        RECT 63.000 190.800 63.400 192.700 ;
        RECT 65.600 190.800 66.000 193.100 ;
        RECT 68.600 190.800 69.000 193.100 ;
        RECT 71.000 190.800 71.400 193.100 ;
        RECT 71.800 190.800 72.200 193.100 ;
        RECT 73.400 190.800 73.800 193.100 ;
        RECT 75.800 190.800 76.200 193.100 ;
        RECT 77.400 190.800 77.800 193.100 ;
        RECT 79.800 190.800 80.200 192.700 ;
        RECT 82.200 190.800 82.600 193.000 ;
        RECT 85.000 190.800 85.400 192.100 ;
        RECT 86.600 190.800 87.100 192.100 ;
        RECT 89.400 190.800 89.800 193.100 ;
        RECT 91.600 190.800 92.000 193.500 ;
        RECT 94.200 190.800 94.600 193.300 ;
        RECT 96.600 190.800 97.000 192.700 ;
        RECT 102.200 190.800 102.600 193.100 ;
        RECT 103.800 190.800 104.200 193.000 ;
        RECT 106.600 190.800 107.000 192.100 ;
        RECT 108.200 190.800 108.700 192.100 ;
        RECT 111.000 190.800 111.400 193.100 ;
        RECT 113.200 190.800 113.600 193.500 ;
        RECT 115.800 190.800 116.200 193.300 ;
        RECT 118.200 190.800 118.600 193.000 ;
        RECT 121.000 190.800 121.400 192.100 ;
        RECT 122.600 190.800 123.100 192.100 ;
        RECT 125.400 190.800 125.800 193.100 ;
        RECT 127.600 190.800 128.000 193.500 ;
        RECT 130.200 190.800 130.600 193.300 ;
        RECT 132.400 190.800 132.800 193.500 ;
        RECT 135.000 190.800 135.400 193.300 ;
        RECT 136.800 190.800 137.200 193.100 ;
        RECT 139.800 190.800 140.200 193.100 ;
        RECT 141.200 190.800 141.600 193.500 ;
        RECT 143.800 190.800 144.200 193.300 ;
        RECT 146.200 190.800 146.600 192.700 ;
        RECT 151.000 190.800 151.400 193.100 ;
        RECT 153.700 190.800 154.200 192.100 ;
        RECT 155.400 190.800 155.800 192.100 ;
        RECT 158.200 190.800 158.600 193.000 ;
        RECT 160.600 190.800 161.000 193.000 ;
        RECT 163.400 190.800 163.800 192.100 ;
        RECT 165.000 190.800 165.500 192.100 ;
        RECT 167.800 190.800 168.200 193.100 ;
        RECT 169.400 190.800 169.800 193.100 ;
        RECT 173.400 190.800 173.800 192.700 ;
        RECT 175.000 190.800 175.400 193.100 ;
        RECT 176.600 190.800 177.000 193.100 ;
        RECT 178.200 190.800 178.600 193.100 ;
        RECT 179.800 190.800 180.200 193.100 ;
        RECT 181.400 190.800 181.800 193.100 ;
        RECT 183.800 190.800 184.200 192.700 ;
        RECT 187.000 190.800 187.400 193.100 ;
        RECT 187.800 190.800 188.200 193.100 ;
        RECT 190.800 190.800 191.200 193.100 ;
        RECT 192.600 190.800 193.000 193.300 ;
        RECT 195.200 190.800 195.600 193.500 ;
        RECT 197.200 190.800 197.600 193.500 ;
        RECT 199.800 190.800 200.200 193.300 ;
        RECT 203.800 190.800 204.200 193.000 ;
        RECT 206.600 190.800 207.000 192.100 ;
        RECT 208.200 190.800 208.700 192.100 ;
        RECT 211.000 190.800 211.400 193.100 ;
        RECT 213.400 190.800 213.800 192.700 ;
        RECT 216.600 190.800 217.000 192.700 ;
        RECT 220.600 190.800 221.000 193.100 ;
        RECT 222.200 190.800 222.600 193.000 ;
        RECT 225.000 190.800 225.400 192.100 ;
        RECT 226.600 190.800 227.100 192.100 ;
        RECT 229.400 190.800 229.800 193.100 ;
        RECT 231.800 190.800 232.200 192.700 ;
        RECT 235.000 190.800 235.400 193.000 ;
        RECT 237.800 190.800 238.200 192.100 ;
        RECT 239.400 190.800 239.900 192.100 ;
        RECT 242.200 190.800 242.600 193.100 ;
        RECT 245.400 190.800 245.800 192.700 ;
        RECT 247.800 190.800 248.200 193.100 ;
        RECT 249.400 190.800 249.800 193.100 ;
        RECT 0.200 190.200 252.600 190.800 ;
        RECT 0.600 187.900 1.000 190.200 ;
        RECT 4.600 188.300 5.000 190.200 ;
        RECT 7.000 188.300 7.400 190.200 ;
        RECT 11.000 187.900 11.400 190.200 ;
        RECT 12.400 187.500 12.800 190.200 ;
        RECT 15.000 187.700 15.400 190.200 ;
        RECT 16.600 187.900 17.000 190.200 ;
        RECT 18.200 187.900 18.600 190.200 ;
        RECT 19.800 187.900 20.200 190.200 ;
        RECT 21.400 187.900 21.800 190.200 ;
        RECT 23.000 187.900 23.400 190.200 ;
        RECT 24.400 187.500 24.800 190.200 ;
        RECT 27.000 187.700 27.400 190.200 ;
        RECT 29.200 187.500 29.600 190.200 ;
        RECT 31.800 187.700 32.200 190.200 ;
        RECT 33.400 187.900 33.800 190.200 ;
        RECT 35.000 187.900 35.400 190.200 ;
        RECT 36.600 187.900 37.000 190.200 ;
        RECT 38.200 187.900 38.600 190.200 ;
        RECT 39.800 187.900 40.200 190.200 ;
        RECT 40.600 188.900 41.000 190.200 ;
        RECT 42.200 188.900 42.600 190.200 ;
        RECT 43.000 188.900 43.400 190.200 ;
        RECT 45.100 187.900 45.500 190.200 ;
        RECT 48.600 188.000 49.000 190.200 ;
        RECT 51.400 188.900 51.800 190.200 ;
        RECT 53.000 188.900 53.500 190.200 ;
        RECT 55.800 187.900 56.200 190.200 ;
        RECT 58.200 187.700 58.600 190.200 ;
        RECT 60.800 187.500 61.200 190.200 ;
        RECT 62.800 187.500 63.200 190.200 ;
        RECT 65.400 187.700 65.800 190.200 ;
        RECT 67.800 187.700 68.200 190.200 ;
        RECT 70.400 187.500 70.800 190.200 ;
        RECT 71.800 187.900 72.200 190.200 ;
        RECT 74.800 187.900 75.200 190.200 ;
        RECT 76.600 187.900 77.000 190.200 ;
        RECT 79.300 188.900 79.800 190.200 ;
        RECT 81.000 188.900 81.400 190.200 ;
        RECT 83.800 188.000 84.200 190.200 ;
        RECT 85.400 187.900 85.800 190.200 ;
        RECT 89.400 188.300 89.800 190.200 ;
        RECT 91.000 187.900 91.400 190.200 ;
        RECT 95.000 188.300 95.400 190.200 ;
        RECT 97.200 187.500 97.600 190.200 ;
        RECT 99.800 187.700 100.200 190.200 ;
        RECT 103.800 187.900 104.200 190.200 ;
        RECT 106.500 188.900 107.000 190.200 ;
        RECT 108.200 188.900 108.600 190.200 ;
        RECT 111.000 188.000 111.400 190.200 ;
        RECT 112.600 187.900 113.000 190.200 ;
        RECT 116.600 188.300 117.000 190.200 ;
        RECT 119.000 188.300 119.400 190.200 ;
        RECT 122.200 188.000 122.600 190.200 ;
        RECT 125.000 188.900 125.400 190.200 ;
        RECT 126.600 188.900 127.100 190.200 ;
        RECT 129.400 187.900 129.800 190.200 ;
        RECT 131.800 188.300 132.200 190.200 ;
        RECT 134.200 187.900 134.600 190.200 ;
        RECT 135.800 187.900 136.200 190.200 ;
        RECT 137.400 187.900 137.800 190.200 ;
        RECT 139.000 187.900 139.400 190.200 ;
        RECT 140.600 187.900 141.000 190.200 ;
        RECT 141.400 188.900 141.800 190.200 ;
        RECT 143.000 188.900 143.400 190.200 ;
        RECT 143.800 188.900 144.200 190.200 ;
        RECT 145.900 187.900 146.300 190.200 ;
        RECT 148.600 187.900 149.000 190.200 ;
        RECT 151.200 187.900 151.600 190.200 ;
        RECT 154.200 187.900 154.600 190.200 ;
        RECT 155.800 187.900 156.200 190.200 ;
        RECT 157.400 187.900 157.800 190.200 ;
        RECT 159.800 187.900 160.200 190.200 ;
        RECT 160.600 187.900 161.000 190.200 ;
        RECT 163.800 188.300 164.200 190.200 ;
        RECT 167.000 188.000 167.400 190.200 ;
        RECT 169.800 188.900 170.200 190.200 ;
        RECT 171.400 188.900 171.900 190.200 ;
        RECT 174.200 187.900 174.600 190.200 ;
        RECT 176.600 187.700 177.000 190.200 ;
        RECT 179.200 187.500 179.600 190.200 ;
        RECT 181.400 188.300 181.800 190.200 ;
        RECT 185.400 187.900 185.800 190.200 ;
        RECT 186.200 187.900 186.600 190.200 ;
        RECT 189.200 187.900 189.600 190.200 ;
        RECT 191.000 188.000 191.400 190.200 ;
        RECT 193.800 188.900 194.200 190.200 ;
        RECT 195.400 188.900 195.900 190.200 ;
        RECT 198.200 187.900 198.600 190.200 ;
        RECT 201.400 187.900 201.800 190.200 ;
        RECT 204.600 188.000 205.000 190.200 ;
        RECT 207.400 188.900 207.800 190.200 ;
        RECT 209.000 188.900 209.500 190.200 ;
        RECT 211.800 187.900 212.200 190.200 ;
        RECT 213.400 187.900 213.800 190.200 ;
        RECT 216.600 187.700 217.000 190.200 ;
        RECT 219.200 187.500 219.600 190.200 ;
        RECT 221.200 187.500 221.600 190.200 ;
        RECT 223.800 187.700 224.200 190.200 ;
        RECT 226.200 188.300 226.600 190.200 ;
        RECT 230.200 187.900 230.600 190.200 ;
        RECT 231.800 187.900 232.200 190.200 ;
        RECT 234.500 188.900 235.000 190.200 ;
        RECT 236.200 188.900 236.600 190.200 ;
        RECT 239.000 188.000 239.400 190.200 ;
        RECT 240.600 187.900 241.000 190.200 ;
        RECT 242.200 187.900 242.600 190.200 ;
        RECT 243.800 187.900 244.200 190.200 ;
        RECT 245.400 187.900 245.800 190.200 ;
        RECT 247.000 187.900 247.400 190.200 ;
        RECT 247.800 187.900 248.200 190.200 ;
        RECT 249.400 187.900 249.800 190.200 ;
        RECT 1.400 170.800 1.800 173.000 ;
        RECT 4.200 170.800 4.600 172.100 ;
        RECT 5.800 170.800 6.300 172.100 ;
        RECT 8.600 170.800 9.000 173.100 ;
        RECT 11.800 170.800 12.200 172.700 ;
        RECT 15.000 170.800 15.400 173.100 ;
        RECT 15.800 170.800 16.200 173.100 ;
        RECT 19.000 170.800 19.400 172.700 ;
        RECT 23.000 170.800 23.400 173.100 ;
        RECT 24.600 170.800 25.000 173.100 ;
        RECT 27.300 170.800 27.800 172.100 ;
        RECT 29.000 170.800 29.400 172.100 ;
        RECT 31.800 170.800 32.200 173.000 ;
        RECT 34.200 170.800 34.600 173.000 ;
        RECT 37.000 170.800 37.400 172.100 ;
        RECT 38.600 170.800 39.100 172.100 ;
        RECT 41.400 170.800 41.800 173.100 ;
        RECT 44.600 170.800 45.000 172.700 ;
        RECT 48.600 170.800 49.000 173.300 ;
        RECT 51.200 170.800 51.600 173.500 ;
        RECT 54.200 170.800 54.600 173.100 ;
        RECT 55.200 170.800 55.600 173.100 ;
        RECT 58.200 170.800 58.600 173.100 ;
        RECT 59.000 170.800 59.400 173.100 ;
        RECT 63.000 170.800 63.400 172.700 ;
        RECT 65.400 170.800 65.800 173.000 ;
        RECT 68.200 170.800 68.600 172.100 ;
        RECT 69.800 170.800 70.300 172.100 ;
        RECT 72.600 170.800 73.000 173.100 ;
        RECT 74.800 170.800 75.200 173.500 ;
        RECT 77.400 170.800 77.800 173.300 ;
        RECT 79.800 170.800 80.200 173.100 ;
        RECT 82.500 170.800 83.000 172.100 ;
        RECT 84.200 170.800 84.600 172.100 ;
        RECT 87.000 170.800 87.400 173.000 ;
        RECT 89.200 170.800 89.600 173.500 ;
        RECT 91.800 170.800 92.200 173.300 ;
        RECT 94.000 170.800 94.400 173.500 ;
        RECT 96.600 170.800 97.000 173.300 ;
        RECT 100.400 170.800 100.800 173.500 ;
        RECT 103.000 170.800 103.400 173.300 ;
        RECT 105.400 170.800 105.800 173.000 ;
        RECT 108.200 170.800 108.600 172.100 ;
        RECT 109.800 170.800 110.300 172.100 ;
        RECT 112.600 170.800 113.000 173.100 ;
        RECT 114.200 170.800 114.600 173.100 ;
        RECT 118.200 170.800 118.600 172.700 ;
        RECT 121.400 170.800 121.800 173.100 ;
        RECT 122.200 170.800 122.600 173.100 ;
        RECT 123.800 170.800 124.200 173.100 ;
        RECT 126.000 170.800 126.400 173.500 ;
        RECT 128.600 170.800 129.000 173.300 ;
        RECT 130.400 170.800 130.800 173.100 ;
        RECT 133.400 170.800 133.800 173.100 ;
        RECT 134.800 170.800 135.200 173.500 ;
        RECT 137.400 170.800 137.800 173.300 ;
        RECT 139.600 170.800 140.000 173.500 ;
        RECT 142.200 170.800 142.600 173.300 ;
        RECT 144.400 170.800 144.800 173.500 ;
        RECT 147.000 170.800 147.400 173.300 ;
        RECT 148.600 170.800 149.000 173.100 ;
        RECT 154.200 170.800 154.600 172.700 ;
        RECT 156.600 170.800 157.000 173.000 ;
        RECT 159.400 170.800 159.800 172.100 ;
        RECT 161.000 170.800 161.500 172.100 ;
        RECT 163.800 170.800 164.200 173.100 ;
        RECT 166.000 170.800 166.400 173.500 ;
        RECT 168.600 170.800 169.000 173.300 ;
        RECT 170.200 170.800 170.600 173.100 ;
        RECT 174.200 170.800 174.600 172.700 ;
        RECT 176.600 170.800 177.000 173.000 ;
        RECT 179.400 170.800 179.800 172.100 ;
        RECT 181.000 170.800 181.500 172.100 ;
        RECT 183.800 170.800 184.200 173.100 ;
        RECT 186.200 170.800 186.600 173.100 ;
        RECT 187.800 170.800 188.200 173.100 ;
        RECT 189.400 170.800 189.800 173.100 ;
        RECT 192.100 170.800 192.600 172.100 ;
        RECT 193.800 170.800 194.200 172.100 ;
        RECT 196.600 170.800 197.000 173.000 ;
        RECT 199.000 170.800 199.400 173.300 ;
        RECT 201.600 170.800 202.000 173.500 ;
        RECT 204.600 170.800 205.000 173.100 ;
        RECT 207.600 170.800 208.000 173.100 ;
        RECT 209.400 170.800 209.800 172.700 ;
        RECT 212.600 170.800 213.000 173.000 ;
        RECT 215.400 170.800 215.800 172.100 ;
        RECT 217.000 170.800 217.500 172.100 ;
        RECT 219.800 170.800 220.200 173.100 ;
        RECT 222.000 170.800 222.400 173.500 ;
        RECT 224.600 170.800 225.000 173.300 ;
        RECT 227.000 170.800 227.400 173.300 ;
        RECT 229.600 170.800 230.000 173.500 ;
        RECT 231.600 170.800 232.000 173.500 ;
        RECT 234.200 170.800 234.600 173.300 ;
        RECT 235.800 170.800 236.200 173.100 ;
        RECT 239.000 170.800 239.400 173.000 ;
        RECT 241.800 170.800 242.200 172.100 ;
        RECT 243.400 170.800 243.900 172.100 ;
        RECT 246.200 170.800 246.600 173.100 ;
        RECT 248.600 170.800 249.000 172.700 ;
        RECT 0.200 170.200 252.600 170.800 ;
        RECT 0.600 167.900 1.000 170.200 ;
        RECT 2.200 167.900 2.600 170.200 ;
        RECT 3.800 167.900 4.200 170.200 ;
        RECT 5.400 167.900 5.800 170.200 ;
        RECT 7.000 167.900 7.400 170.200 ;
        RECT 8.600 167.900 9.000 170.200 ;
        RECT 11.300 168.900 11.800 170.200 ;
        RECT 13.000 168.900 13.400 170.200 ;
        RECT 15.800 168.000 16.200 170.200 ;
        RECT 19.000 168.300 19.400 170.200 ;
        RECT 21.400 167.900 21.800 170.200 ;
        RECT 24.100 168.900 24.600 170.200 ;
        RECT 25.800 168.900 26.200 170.200 ;
        RECT 28.600 168.000 29.000 170.200 ;
        RECT 30.200 167.900 30.600 170.200 ;
        RECT 34.200 168.300 34.600 170.200 ;
        RECT 36.400 167.500 36.800 170.200 ;
        RECT 39.000 167.700 39.400 170.200 ;
        RECT 40.600 167.900 41.000 170.200 ;
        RECT 43.600 167.500 44.000 170.200 ;
        RECT 46.200 167.700 46.600 170.200 ;
        RECT 49.400 167.900 49.800 170.200 ;
        RECT 52.400 167.900 52.800 170.200 ;
        RECT 54.200 167.900 54.600 170.200 ;
        RECT 56.900 168.900 57.400 170.200 ;
        RECT 58.600 168.900 59.000 170.200 ;
        RECT 61.400 168.000 61.800 170.200 ;
        RECT 63.800 168.300 64.200 170.200 ;
        RECT 67.800 167.900 68.200 170.200 ;
        RECT 69.400 167.700 69.800 170.200 ;
        RECT 72.000 167.500 72.400 170.200 ;
        RECT 74.000 167.500 74.400 170.200 ;
        RECT 76.600 167.700 77.000 170.200 ;
        RECT 79.000 168.300 79.400 170.200 ;
        RECT 83.000 167.900 83.400 170.200 ;
        RECT 83.800 167.900 84.200 170.200 ;
        RECT 86.800 167.900 87.200 170.200 ;
        RECT 88.600 168.000 89.000 170.200 ;
        RECT 91.400 168.900 91.800 170.200 ;
        RECT 93.000 168.900 93.500 170.200 ;
        RECT 95.800 167.900 96.200 170.200 ;
        RECT 97.400 167.900 97.800 170.200 ;
        RECT 103.000 168.300 103.400 170.200 ;
        RECT 105.400 167.900 105.800 170.200 ;
        RECT 108.100 168.900 108.600 170.200 ;
        RECT 109.800 168.900 110.200 170.200 ;
        RECT 112.600 168.000 113.000 170.200 ;
        RECT 115.000 168.300 115.400 170.200 ;
        RECT 119.000 167.900 119.400 170.200 ;
        RECT 120.400 167.500 120.800 170.200 ;
        RECT 123.000 167.700 123.400 170.200 ;
        RECT 124.600 167.900 125.000 170.200 ;
        RECT 128.600 168.300 129.000 170.200 ;
        RECT 131.800 167.900 132.200 170.200 ;
        RECT 133.400 168.000 133.800 170.200 ;
        RECT 136.200 168.900 136.600 170.200 ;
        RECT 137.800 168.900 138.300 170.200 ;
        RECT 140.600 167.900 141.000 170.200 ;
        RECT 143.000 168.300 143.400 170.200 ;
        RECT 146.200 168.000 146.600 170.200 ;
        RECT 149.000 168.900 149.400 170.200 ;
        RECT 150.600 168.900 151.100 170.200 ;
        RECT 153.400 167.900 153.800 170.200 ;
        RECT 157.400 167.700 157.800 170.200 ;
        RECT 160.000 167.500 160.400 170.200 ;
        RECT 161.400 167.900 161.800 170.200 ;
        RECT 164.400 167.900 164.800 170.200 ;
        RECT 166.200 168.300 166.600 170.200 ;
        RECT 170.200 167.900 170.600 170.200 ;
        RECT 171.800 167.700 172.200 170.200 ;
        RECT 174.400 167.500 174.800 170.200 ;
        RECT 176.600 167.700 177.000 170.200 ;
        RECT 179.200 167.500 179.600 170.200 ;
        RECT 182.200 167.900 182.600 170.200 ;
        RECT 183.800 168.000 184.200 170.200 ;
        RECT 186.600 168.900 187.000 170.200 ;
        RECT 188.200 168.900 188.700 170.200 ;
        RECT 191.000 167.900 191.400 170.200 ;
        RECT 193.400 168.300 193.800 170.200 ;
        RECT 197.400 167.900 197.800 170.200 ;
        RECT 199.000 167.700 199.400 170.200 ;
        RECT 201.600 167.500 202.000 170.200 ;
        RECT 205.400 167.700 205.800 170.200 ;
        RECT 208.000 167.500 208.400 170.200 ;
        RECT 209.400 167.900 209.800 170.200 ;
        RECT 211.800 167.900 212.200 170.200 ;
        RECT 215.800 168.300 216.200 170.200 ;
        RECT 218.200 168.000 218.600 170.200 ;
        RECT 221.000 168.900 221.400 170.200 ;
        RECT 222.600 168.900 223.100 170.200 ;
        RECT 225.400 167.900 225.800 170.200 ;
        RECT 227.000 167.900 227.400 170.200 ;
        RECT 228.600 167.900 229.000 170.200 ;
        RECT 230.200 167.900 230.600 170.200 ;
        RECT 231.800 167.900 232.200 170.200 ;
        RECT 233.400 167.900 233.800 170.200 ;
        RECT 235.000 168.000 235.400 170.200 ;
        RECT 237.800 168.900 238.200 170.200 ;
        RECT 239.400 168.900 239.900 170.200 ;
        RECT 242.200 167.900 242.600 170.200 ;
        RECT 243.800 167.900 244.200 170.200 ;
        RECT 245.400 167.900 245.800 170.200 ;
        RECT 248.600 168.300 249.000 170.200 ;
        RECT 1.400 150.800 1.800 153.100 ;
        RECT 4.100 150.800 4.600 152.100 ;
        RECT 5.800 150.800 6.200 152.100 ;
        RECT 8.600 150.800 9.000 153.000 ;
        RECT 10.200 150.800 10.600 153.100 ;
        RECT 14.200 150.800 14.600 152.700 ;
        RECT 16.400 150.800 16.800 153.500 ;
        RECT 19.000 150.800 19.400 153.300 ;
        RECT 21.400 150.800 21.800 152.700 ;
        RECT 25.400 150.800 25.800 153.100 ;
        RECT 27.000 150.800 27.400 153.000 ;
        RECT 29.800 150.800 30.200 152.100 ;
        RECT 31.400 150.800 31.900 152.100 ;
        RECT 34.200 150.800 34.600 153.100 ;
        RECT 35.800 150.800 36.200 152.100 ;
        RECT 37.400 150.800 37.800 152.100 ;
        RECT 38.200 150.800 38.600 152.100 ;
        RECT 39.800 150.800 40.200 152.100 ;
        RECT 41.400 150.800 41.800 153.100 ;
        RECT 42.800 150.800 43.200 153.500 ;
        RECT 45.400 150.800 45.800 153.300 ;
        RECT 47.000 150.800 47.400 152.100 ;
        RECT 48.600 150.800 49.000 152.100 ;
        RECT 51.000 150.800 51.400 152.100 ;
        RECT 52.600 150.800 53.000 152.100 ;
        RECT 54.200 150.800 54.600 153.000 ;
        RECT 57.000 150.800 57.400 152.100 ;
        RECT 58.600 150.800 59.100 152.100 ;
        RECT 61.400 150.800 61.800 153.100 ;
        RECT 63.000 150.800 63.400 153.100 ;
        RECT 67.000 150.800 67.400 152.700 ;
        RECT 68.600 150.800 69.000 153.100 ;
        RECT 70.200 150.800 70.600 153.100 ;
        RECT 71.800 150.800 72.200 153.100 ;
        RECT 73.400 150.800 73.800 153.100 ;
        RECT 75.000 150.800 75.400 153.100 ;
        RECT 76.600 150.800 77.000 152.700 ;
        RECT 79.000 150.800 79.400 153.100 ;
        RECT 82.200 150.800 82.600 153.000 ;
        RECT 85.000 150.800 85.400 152.100 ;
        RECT 86.600 150.800 87.100 152.100 ;
        RECT 89.400 150.800 89.800 153.100 ;
        RECT 91.800 150.800 92.200 153.100 ;
        RECT 93.700 150.800 94.100 153.100 ;
        RECT 95.800 150.800 96.200 152.100 ;
        RECT 96.600 150.800 97.000 152.100 ;
        RECT 98.200 150.800 98.600 152.100 ;
        RECT 100.900 150.800 101.300 153.100 ;
        RECT 103.000 150.800 103.400 152.100 ;
        RECT 103.800 150.800 104.200 152.100 ;
        RECT 105.400 150.800 105.800 152.100 ;
        RECT 106.500 150.800 106.900 153.100 ;
        RECT 108.600 150.800 109.000 152.100 ;
        RECT 109.400 150.800 109.800 152.100 ;
        RECT 111.000 150.800 111.400 152.100 ;
        RECT 111.800 150.800 112.200 153.100 ;
        RECT 113.400 150.800 113.800 153.100 ;
        RECT 115.000 150.800 115.400 153.100 ;
        RECT 117.700 150.800 118.200 152.100 ;
        RECT 119.400 150.800 119.800 152.100 ;
        RECT 122.200 150.800 122.600 153.000 ;
        RECT 123.800 150.800 124.200 153.100 ;
        RECT 127.800 150.800 128.200 152.700 ;
        RECT 130.200 150.800 130.600 153.300 ;
        RECT 132.800 150.800 133.200 153.500 ;
        RECT 135.000 150.800 135.400 153.100 ;
        RECT 137.700 150.800 138.200 152.100 ;
        RECT 139.400 150.800 139.800 152.100 ;
        RECT 142.200 150.800 142.600 153.000 ;
        RECT 145.400 150.800 145.800 153.100 ;
        RECT 146.200 150.800 146.600 153.100 ;
        RECT 150.800 150.800 151.200 153.500 ;
        RECT 153.400 150.800 153.800 153.300 ;
        RECT 155.800 150.800 156.200 152.700 ;
        RECT 159.800 150.800 160.200 153.100 ;
        RECT 161.400 150.800 161.800 153.000 ;
        RECT 164.200 150.800 164.600 152.100 ;
        RECT 165.800 150.800 166.300 152.100 ;
        RECT 168.600 150.800 169.000 153.100 ;
        RECT 170.200 150.800 170.600 153.100 ;
        RECT 173.400 150.800 173.800 152.700 ;
        RECT 177.400 150.800 177.800 153.100 ;
        RECT 179.000 150.800 179.400 153.300 ;
        RECT 181.600 150.800 182.000 153.500 ;
        RECT 183.800 150.800 184.200 153.000 ;
        RECT 186.600 150.800 187.000 152.100 ;
        RECT 188.200 150.800 188.700 152.100 ;
        RECT 191.000 150.800 191.400 153.100 ;
        RECT 192.600 150.800 193.000 153.100 ;
        RECT 196.600 150.800 197.000 152.700 ;
        RECT 199.000 150.800 199.400 152.700 ;
        RECT 204.600 150.800 205.000 153.100 ;
        RECT 206.200 150.800 206.600 153.000 ;
        RECT 209.000 150.800 209.400 152.100 ;
        RECT 210.600 150.800 211.100 152.100 ;
        RECT 213.400 150.800 213.800 153.100 ;
        RECT 215.800 150.800 216.200 153.000 ;
        RECT 218.600 150.800 219.000 152.100 ;
        RECT 220.200 150.800 220.700 152.100 ;
        RECT 223.000 150.800 223.400 153.100 ;
        RECT 224.600 150.800 225.000 153.100 ;
        RECT 226.200 150.800 226.600 153.100 ;
        RECT 227.800 150.800 228.200 153.100 ;
        RECT 229.400 150.800 229.800 153.100 ;
        RECT 231.000 150.800 231.400 153.100 ;
        RECT 232.600 150.800 233.000 152.700 ;
        RECT 236.600 150.800 237.000 153.100 ;
        RECT 238.200 150.800 238.600 153.000 ;
        RECT 241.000 150.800 241.400 152.100 ;
        RECT 242.600 150.800 243.100 152.100 ;
        RECT 245.400 150.800 245.800 153.100 ;
        RECT 247.000 150.800 247.400 152.100 ;
        RECT 248.600 150.800 249.000 152.100 ;
        RECT 249.400 150.800 249.800 153.100 ;
        RECT 0.200 150.200 252.600 150.800 ;
        RECT 1.400 147.900 1.800 150.200 ;
        RECT 4.100 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.200 150.200 ;
        RECT 8.600 148.000 9.000 150.200 ;
        RECT 10.200 147.900 10.600 150.200 ;
        RECT 14.200 148.300 14.600 150.200 ;
        RECT 16.600 147.900 17.000 150.200 ;
        RECT 19.300 148.900 19.800 150.200 ;
        RECT 21.000 148.900 21.400 150.200 ;
        RECT 23.800 148.000 24.200 150.200 ;
        RECT 26.200 148.300 26.600 150.200 ;
        RECT 30.200 147.900 30.600 150.200 ;
        RECT 31.000 148.900 31.400 150.200 ;
        RECT 32.600 147.900 33.000 150.200 ;
        RECT 36.600 147.900 37.000 150.200 ;
        RECT 38.200 148.900 38.600 150.200 ;
        RECT 39.600 147.500 40.000 150.200 ;
        RECT 42.200 147.700 42.600 150.200 ;
        RECT 43.800 147.900 44.200 150.200 ;
        RECT 46.200 147.900 46.600 150.200 ;
        RECT 50.200 148.900 50.600 150.200 ;
        RECT 51.800 148.900 52.200 150.200 ;
        RECT 52.600 148.900 53.000 150.200 ;
        RECT 54.200 148.900 54.600 150.200 ;
        RECT 55.000 148.900 55.400 150.200 ;
        RECT 56.600 148.900 57.000 150.200 ;
        RECT 57.400 148.900 57.800 150.200 ;
        RECT 59.000 148.100 59.400 150.200 ;
        RECT 60.600 147.900 61.000 150.200 ;
        RECT 62.200 147.900 62.600 150.200 ;
        RECT 63.800 147.900 64.200 150.200 ;
        RECT 65.400 147.900 65.800 150.200 ;
        RECT 68.100 148.900 68.600 150.200 ;
        RECT 69.800 148.900 70.200 150.200 ;
        RECT 72.600 148.000 73.000 150.200 ;
        RECT 74.200 148.900 74.600 150.200 ;
        RECT 76.300 147.900 76.700 150.200 ;
        RECT 79.000 147.900 79.400 150.200 ;
        RECT 80.600 148.000 81.000 150.200 ;
        RECT 83.400 148.900 83.800 150.200 ;
        RECT 85.000 148.900 85.500 150.200 ;
        RECT 87.800 147.900 88.200 150.200 ;
        RECT 89.400 147.900 89.800 150.200 ;
        RECT 91.000 147.900 91.400 150.200 ;
        RECT 92.600 147.900 93.000 150.200 ;
        RECT 94.200 147.900 94.600 150.200 ;
        RECT 95.800 147.900 96.200 150.200 ;
        RECT 99.000 147.900 99.400 150.200 ;
        RECT 101.700 148.900 102.200 150.200 ;
        RECT 103.400 148.900 103.800 150.200 ;
        RECT 106.200 148.000 106.600 150.200 ;
        RECT 108.600 147.900 109.000 150.200 ;
        RECT 111.300 148.900 111.800 150.200 ;
        RECT 113.000 148.900 113.400 150.200 ;
        RECT 115.800 148.000 116.200 150.200 ;
        RECT 118.200 147.700 118.600 150.200 ;
        RECT 120.800 147.500 121.200 150.200 ;
        RECT 123.000 147.900 123.400 150.200 ;
        RECT 125.700 148.900 126.200 150.200 ;
        RECT 127.400 148.900 127.800 150.200 ;
        RECT 130.200 148.000 130.600 150.200 ;
        RECT 132.400 147.500 132.800 150.200 ;
        RECT 135.000 147.700 135.400 150.200 ;
        RECT 137.400 148.000 137.800 150.200 ;
        RECT 140.200 148.900 140.600 150.200 ;
        RECT 141.800 148.900 142.300 150.200 ;
        RECT 144.600 147.900 145.000 150.200 ;
        RECT 147.000 148.300 147.400 150.200 ;
        RECT 149.400 147.900 149.800 150.200 ;
        RECT 155.000 148.300 155.400 150.200 ;
        RECT 157.400 148.300 157.800 150.200 ;
        RECT 161.400 147.900 161.800 150.200 ;
        RECT 163.000 147.900 163.400 150.200 ;
        RECT 165.700 148.900 166.200 150.200 ;
        RECT 167.400 148.900 167.800 150.200 ;
        RECT 170.200 148.000 170.600 150.200 ;
        RECT 173.400 148.300 173.800 150.200 ;
        RECT 175.800 148.000 176.200 150.200 ;
        RECT 178.600 148.900 179.000 150.200 ;
        RECT 180.200 148.900 180.700 150.200 ;
        RECT 183.000 147.900 183.400 150.200 ;
        RECT 184.600 147.900 185.000 150.200 ;
        RECT 186.200 147.900 186.600 150.200 ;
        RECT 187.800 147.900 188.200 150.200 ;
        RECT 189.400 147.900 189.800 150.200 ;
        RECT 191.000 147.900 191.400 150.200 ;
        RECT 192.600 147.700 193.000 150.200 ;
        RECT 195.200 147.500 195.600 150.200 ;
        RECT 197.400 148.300 197.800 150.200 ;
        RECT 201.400 147.900 201.800 150.200 ;
        RECT 204.600 147.700 205.000 150.200 ;
        RECT 207.200 147.500 207.600 150.200 ;
        RECT 209.400 148.000 209.800 150.200 ;
        RECT 212.200 148.900 212.600 150.200 ;
        RECT 213.800 148.900 214.300 150.200 ;
        RECT 216.600 147.900 217.000 150.200 ;
        RECT 218.800 147.500 219.200 150.200 ;
        RECT 221.400 147.700 221.800 150.200 ;
        RECT 223.000 147.900 223.400 150.200 ;
        RECT 227.000 148.300 227.400 150.200 ;
        RECT 229.400 148.000 229.800 150.200 ;
        RECT 232.200 148.900 232.600 150.200 ;
        RECT 233.800 148.900 234.300 150.200 ;
        RECT 236.600 147.900 237.000 150.200 ;
        RECT 239.000 148.300 239.400 150.200 ;
        RECT 242.200 147.900 242.600 150.200 ;
        RECT 244.900 148.900 245.400 150.200 ;
        RECT 246.600 148.900 247.000 150.200 ;
        RECT 249.400 148.000 249.800 150.200 ;
        RECT 0.600 130.800 1.000 133.100 ;
        RECT 2.200 130.800 2.600 133.100 ;
        RECT 3.800 130.800 4.200 133.100 ;
        RECT 5.400 130.800 5.800 133.100 ;
        RECT 8.100 130.800 8.600 132.100 ;
        RECT 9.800 130.800 10.200 132.100 ;
        RECT 12.600 130.800 13.000 133.000 ;
        RECT 15.000 130.800 15.400 132.700 ;
        RECT 19.000 130.800 19.400 133.100 ;
        RECT 21.400 130.800 21.800 133.100 ;
        RECT 23.000 130.800 23.400 133.300 ;
        RECT 25.600 130.800 26.000 133.500 ;
        RECT 27.800 130.800 28.200 133.100 ;
        RECT 29.400 130.800 29.800 133.100 ;
        RECT 30.200 130.800 30.600 133.100 ;
        RECT 31.800 130.800 32.200 133.100 ;
        RECT 33.400 130.800 33.800 133.100 ;
        RECT 35.000 130.800 35.400 133.100 ;
        RECT 36.600 130.800 37.000 133.100 ;
        RECT 38.000 130.800 38.400 133.500 ;
        RECT 40.600 130.800 41.000 133.300 ;
        RECT 42.400 130.800 42.800 133.100 ;
        RECT 45.400 130.800 45.800 133.100 ;
        RECT 48.600 130.800 49.000 133.300 ;
        RECT 51.200 130.800 51.600 133.500 ;
        RECT 53.400 130.800 53.800 133.000 ;
        RECT 56.200 130.800 56.600 132.100 ;
        RECT 57.800 130.800 58.300 132.100 ;
        RECT 60.600 130.800 61.000 133.100 ;
        RECT 62.400 130.800 62.800 133.100 ;
        RECT 65.400 130.800 65.800 133.100 ;
        RECT 66.200 130.800 66.600 133.100 ;
        RECT 69.400 130.800 69.800 132.700 ;
        RECT 72.600 130.800 73.000 133.100 ;
        RECT 74.200 130.800 74.600 133.100 ;
        RECT 75.800 130.800 76.200 133.300 ;
        RECT 78.400 130.800 78.800 133.500 ;
        RECT 79.800 130.800 80.200 133.100 ;
        RECT 83.800 130.800 84.200 132.700 ;
        RECT 86.200 130.800 86.600 132.700 ;
        RECT 90.200 130.800 90.600 133.100 ;
        RECT 91.800 130.800 92.200 133.100 ;
        RECT 94.500 130.800 95.000 132.100 ;
        RECT 96.200 130.800 96.600 132.100 ;
        RECT 99.000 130.800 99.400 133.000 ;
        RECT 103.000 130.800 103.400 133.100 ;
        RECT 105.700 130.800 106.200 132.100 ;
        RECT 107.400 130.800 107.800 132.100 ;
        RECT 110.200 130.800 110.600 133.000 ;
        RECT 111.800 130.800 112.200 133.100 ;
        RECT 115.800 130.800 116.200 132.700 ;
        RECT 118.000 130.800 118.400 133.500 ;
        RECT 120.600 130.800 121.000 133.300 ;
        RECT 122.200 130.800 122.600 133.100 ;
        RECT 126.200 130.800 126.600 132.700 ;
        RECT 128.600 130.800 129.000 133.000 ;
        RECT 131.400 130.800 131.800 132.100 ;
        RECT 133.000 130.800 133.500 132.100 ;
        RECT 135.800 130.800 136.200 133.100 ;
        RECT 138.200 130.800 138.600 133.100 ;
        RECT 140.900 130.800 141.400 132.100 ;
        RECT 142.600 130.800 143.000 132.100 ;
        RECT 145.400 130.800 145.800 133.000 ;
        RECT 147.000 130.800 147.400 133.100 ;
        RECT 151.600 130.800 152.000 133.500 ;
        RECT 154.200 130.800 154.600 133.300 ;
        RECT 156.600 130.800 157.000 133.100 ;
        RECT 159.300 130.800 159.800 132.100 ;
        RECT 161.000 130.800 161.400 132.100 ;
        RECT 163.800 130.800 164.200 133.000 ;
        RECT 166.200 130.800 166.600 133.300 ;
        RECT 168.800 130.800 169.200 133.500 ;
        RECT 170.200 130.800 170.600 133.100 ;
        RECT 174.200 130.800 174.600 132.700 ;
        RECT 176.600 130.800 177.000 133.300 ;
        RECT 179.200 130.800 179.600 133.500 ;
        RECT 180.600 130.800 181.000 133.100 ;
        RECT 183.600 130.800 184.000 133.100 ;
        RECT 186.200 130.800 186.600 133.100 ;
        RECT 187.800 130.800 188.200 133.100 ;
        RECT 189.400 130.800 189.800 133.100 ;
        RECT 190.800 130.800 191.200 133.500 ;
        RECT 193.400 130.800 193.800 133.300 ;
        RECT 195.800 130.800 196.200 132.700 ;
        RECT 199.800 130.800 200.200 133.100 ;
        RECT 203.000 130.800 203.400 133.000 ;
        RECT 205.800 130.800 206.200 132.100 ;
        RECT 207.400 130.800 207.900 132.100 ;
        RECT 210.200 130.800 210.600 133.100 ;
        RECT 211.800 130.800 212.200 133.100 ;
        RECT 215.800 130.800 216.200 132.700 ;
        RECT 218.200 130.800 218.600 133.000 ;
        RECT 221.000 130.800 221.400 132.100 ;
        RECT 222.600 130.800 223.100 132.100 ;
        RECT 225.400 130.800 225.800 133.100 ;
        RECT 227.800 130.800 228.200 133.000 ;
        RECT 230.600 130.800 231.000 132.100 ;
        RECT 232.200 130.800 232.700 132.100 ;
        RECT 235.000 130.800 235.400 133.100 ;
        RECT 238.200 130.800 238.600 132.700 ;
        RECT 239.800 130.800 240.200 133.100 ;
        RECT 241.400 130.800 241.800 133.100 ;
        RECT 243.000 130.800 243.400 133.100 ;
        RECT 244.600 130.800 245.000 133.100 ;
        RECT 246.200 130.800 246.600 133.100 ;
        RECT 247.800 130.800 248.200 133.100 ;
        RECT 249.400 130.800 249.800 133.100 ;
        RECT 0.200 130.200 252.600 130.800 ;
        RECT 1.400 127.900 1.800 130.200 ;
        RECT 4.100 128.900 4.600 130.200 ;
        RECT 5.800 128.900 6.200 130.200 ;
        RECT 8.600 128.000 9.000 130.200 ;
        RECT 11.800 127.900 12.200 130.200 ;
        RECT 14.200 128.300 14.600 130.200 ;
        RECT 16.600 128.300 17.000 130.200 ;
        RECT 19.800 127.900 20.200 130.200 ;
        RECT 22.500 128.900 23.000 130.200 ;
        RECT 24.200 128.900 24.600 130.200 ;
        RECT 27.000 128.000 27.400 130.200 ;
        RECT 29.200 127.500 29.600 130.200 ;
        RECT 31.800 127.700 32.200 130.200 ;
        RECT 34.200 127.700 34.600 130.200 ;
        RECT 36.800 127.500 37.200 130.200 ;
        RECT 39.000 127.700 39.400 130.200 ;
        RECT 41.600 127.500 42.000 130.200 ;
        RECT 43.000 128.900 43.400 130.200 ;
        RECT 44.600 128.900 45.000 130.200 ;
        RECT 45.400 128.900 45.800 130.200 ;
        RECT 47.500 127.900 47.900 130.200 ;
        RECT 51.000 128.000 51.400 130.200 ;
        RECT 53.800 128.900 54.200 130.200 ;
        RECT 55.400 128.900 55.900 130.200 ;
        RECT 58.200 127.900 58.600 130.200 ;
        RECT 59.800 127.900 60.200 130.200 ;
        RECT 63.800 128.300 64.200 130.200 ;
        RECT 66.200 127.900 66.600 130.200 ;
        RECT 67.800 127.900 68.200 130.200 ;
        RECT 68.600 127.900 69.000 130.200 ;
        RECT 70.200 127.900 70.600 130.200 ;
        RECT 71.800 127.900 72.200 130.200 ;
        RECT 73.400 127.900 73.800 130.200 ;
        RECT 75.000 127.900 75.400 130.200 ;
        RECT 76.400 127.500 76.800 130.200 ;
        RECT 79.000 127.700 79.400 130.200 ;
        RECT 80.800 127.900 81.200 130.200 ;
        RECT 83.800 127.900 84.200 130.200 ;
        RECT 86.200 127.900 86.600 130.200 ;
        RECT 87.800 127.900 88.200 130.200 ;
        RECT 89.400 127.900 89.800 130.200 ;
        RECT 90.800 127.500 91.200 130.200 ;
        RECT 93.400 127.700 93.800 130.200 ;
        RECT 95.800 127.700 96.200 130.200 ;
        RECT 98.400 127.500 98.800 130.200 ;
        RECT 101.400 127.900 101.800 130.200 ;
        RECT 104.400 127.900 104.800 130.200 ;
        RECT 106.000 127.500 106.400 130.200 ;
        RECT 108.600 127.700 109.000 130.200 ;
        RECT 110.800 127.500 111.200 130.200 ;
        RECT 113.400 127.700 113.800 130.200 ;
        RECT 115.800 128.300 116.200 130.200 ;
        RECT 119.800 127.900 120.200 130.200 ;
        RECT 121.400 127.900 121.800 130.200 ;
        RECT 124.100 128.900 124.600 130.200 ;
        RECT 125.800 128.900 126.200 130.200 ;
        RECT 128.600 128.000 129.000 130.200 ;
        RECT 131.000 128.000 131.400 130.200 ;
        RECT 133.800 128.900 134.200 130.200 ;
        RECT 135.400 128.900 135.900 130.200 ;
        RECT 138.200 127.900 138.600 130.200 ;
        RECT 139.800 127.900 140.200 130.200 ;
        RECT 143.800 128.300 144.200 130.200 ;
        RECT 146.200 128.300 146.600 130.200 ;
        RECT 151.000 128.000 151.400 130.200 ;
        RECT 153.800 128.900 154.200 130.200 ;
        RECT 155.400 128.900 155.900 130.200 ;
        RECT 158.200 127.900 158.600 130.200 ;
        RECT 159.800 127.900 160.200 130.200 ;
        RECT 163.800 128.300 164.200 130.200 ;
        RECT 166.200 127.700 166.600 130.200 ;
        RECT 168.800 127.500 169.200 130.200 ;
        RECT 171.000 128.300 171.400 130.200 ;
        RECT 175.000 127.900 175.400 130.200 ;
        RECT 176.600 127.900 177.000 130.200 ;
        RECT 179.300 128.900 179.800 130.200 ;
        RECT 181.000 128.900 181.400 130.200 ;
        RECT 183.800 128.000 184.200 130.200 ;
        RECT 186.200 127.700 186.600 130.200 ;
        RECT 188.800 127.500 189.200 130.200 ;
        RECT 190.200 127.900 190.600 130.200 ;
        RECT 193.200 127.900 193.600 130.200 ;
        RECT 194.800 127.500 195.200 130.200 ;
        RECT 197.400 127.700 197.800 130.200 ;
        RECT 201.400 128.000 201.800 130.200 ;
        RECT 204.200 128.900 204.600 130.200 ;
        RECT 205.800 128.900 206.300 130.200 ;
        RECT 208.600 127.900 209.000 130.200 ;
        RECT 210.200 127.900 210.600 130.200 ;
        RECT 214.200 128.300 214.600 130.200 ;
        RECT 216.600 127.700 217.000 130.200 ;
        RECT 219.200 127.500 219.600 130.200 ;
        RECT 222.200 127.900 222.600 130.200 ;
        RECT 224.600 128.300 225.000 130.200 ;
        RECT 227.000 128.000 227.400 130.200 ;
        RECT 229.800 128.900 230.200 130.200 ;
        RECT 231.400 128.900 231.900 130.200 ;
        RECT 234.200 127.900 234.600 130.200 ;
        RECT 235.800 127.900 236.200 130.200 ;
        RECT 238.500 127.900 238.900 130.200 ;
        RECT 240.600 128.900 241.000 130.200 ;
        RECT 242.200 128.000 242.600 130.200 ;
        RECT 245.000 128.900 245.400 130.200 ;
        RECT 246.600 128.900 247.100 130.200 ;
        RECT 249.400 127.900 249.800 130.200 ;
        RECT 0.600 110.800 1.000 113.100 ;
        RECT 2.200 110.800 2.600 113.100 ;
        RECT 3.800 110.800 4.200 113.100 ;
        RECT 5.400 110.800 5.800 113.100 ;
        RECT 7.000 110.800 7.400 113.100 ;
        RECT 7.800 110.800 8.200 113.100 ;
        RECT 11.800 110.800 12.200 112.700 ;
        RECT 14.200 110.800 14.600 113.100 ;
        RECT 16.900 110.800 17.400 112.100 ;
        RECT 18.600 110.800 19.000 112.100 ;
        RECT 21.400 110.800 21.800 113.000 ;
        RECT 23.800 110.800 24.200 113.300 ;
        RECT 26.400 110.800 26.800 113.500 ;
        RECT 27.800 110.800 28.200 113.100 ;
        RECT 31.000 110.800 31.400 112.700 ;
        RECT 34.200 110.800 34.600 113.100 ;
        RECT 36.900 110.800 37.400 112.100 ;
        RECT 38.600 110.800 39.000 112.100 ;
        RECT 41.400 110.800 41.800 113.000 ;
        RECT 44.600 110.800 45.000 112.700 ;
        RECT 48.600 110.800 49.000 113.000 ;
        RECT 51.400 110.800 51.800 112.100 ;
        RECT 53.000 110.800 53.500 112.100 ;
        RECT 55.800 110.800 56.200 113.100 ;
        RECT 58.200 110.800 58.600 112.700 ;
        RECT 62.200 110.800 62.600 113.100 ;
        RECT 63.600 110.800 64.000 113.500 ;
        RECT 66.200 110.800 66.600 113.300 ;
        RECT 68.600 110.800 69.000 113.300 ;
        RECT 71.200 110.800 71.600 113.500 ;
        RECT 72.600 110.800 73.000 113.100 ;
        RECT 75.600 110.800 76.000 113.500 ;
        RECT 78.200 110.800 78.600 113.300 ;
        RECT 80.600 110.800 81.000 112.700 ;
        RECT 84.600 110.800 85.000 113.100 ;
        RECT 86.200 110.800 86.600 113.100 ;
        RECT 88.900 110.800 89.400 112.100 ;
        RECT 90.600 110.800 91.000 112.100 ;
        RECT 93.400 110.800 93.800 113.000 ;
        RECT 95.000 110.800 95.400 113.100 ;
        RECT 97.400 110.800 97.800 113.100 ;
        RECT 103.000 110.800 103.400 112.700 ;
        RECT 104.600 110.800 105.000 113.100 ;
        RECT 108.600 110.800 109.000 112.700 ;
        RECT 111.000 110.800 111.400 113.000 ;
        RECT 113.800 110.800 114.200 112.100 ;
        RECT 115.400 110.800 115.900 112.100 ;
        RECT 118.200 110.800 118.600 113.100 ;
        RECT 120.600 110.800 121.000 113.000 ;
        RECT 123.400 110.800 123.800 112.100 ;
        RECT 125.000 110.800 125.500 112.100 ;
        RECT 127.800 110.800 128.200 113.100 ;
        RECT 129.400 110.800 129.800 113.100 ;
        RECT 131.000 110.800 131.400 113.100 ;
        RECT 132.600 110.800 133.000 113.100 ;
        RECT 134.200 110.800 134.600 113.100 ;
        RECT 135.800 110.800 136.200 113.100 ;
        RECT 137.400 110.800 137.800 113.300 ;
        RECT 140.000 110.800 140.400 113.500 ;
        RECT 141.400 110.800 141.800 113.100 ;
        RECT 145.400 110.800 145.800 112.700 ;
        RECT 149.400 110.800 149.800 113.000 ;
        RECT 152.200 110.800 152.600 112.100 ;
        RECT 153.800 110.800 154.300 112.100 ;
        RECT 156.600 110.800 157.000 113.100 ;
        RECT 159.800 110.800 160.200 112.700 ;
        RECT 162.200 110.800 162.600 113.100 ;
        RECT 164.900 110.800 165.400 112.100 ;
        RECT 166.600 110.800 167.000 112.100 ;
        RECT 169.400 110.800 169.800 113.000 ;
        RECT 171.800 110.800 172.200 112.700 ;
        RECT 175.800 110.800 176.200 113.100 ;
        RECT 177.400 110.800 177.800 113.300 ;
        RECT 180.000 110.800 180.400 113.500 ;
        RECT 181.400 110.800 181.800 113.100 ;
        RECT 183.000 110.800 183.400 113.100 ;
        RECT 184.600 110.800 185.000 113.100 ;
        RECT 188.600 110.800 189.000 113.100 ;
        RECT 191.000 110.800 191.400 112.700 ;
        RECT 193.400 110.800 193.800 112.700 ;
        RECT 197.400 110.800 197.800 113.100 ;
        RECT 200.600 110.800 201.000 113.000 ;
        RECT 203.400 110.800 203.800 112.100 ;
        RECT 205.000 110.800 205.500 112.100 ;
        RECT 207.800 110.800 208.200 113.100 ;
        RECT 210.200 110.800 210.600 113.100 ;
        RECT 212.900 110.800 213.400 112.100 ;
        RECT 214.600 110.800 215.000 112.100 ;
        RECT 217.400 110.800 217.800 113.000 ;
        RECT 219.800 110.800 220.200 112.700 ;
        RECT 222.200 110.800 222.600 113.100 ;
        RECT 223.800 110.800 224.200 113.100 ;
        RECT 226.200 110.800 226.600 113.300 ;
        RECT 228.800 110.800 229.200 113.500 ;
        RECT 231.000 110.800 231.400 113.300 ;
        RECT 233.600 110.800 234.000 113.500 ;
        RECT 235.800 110.800 236.200 113.100 ;
        RECT 237.400 110.800 237.800 113.100 ;
        RECT 238.200 110.800 238.600 113.100 ;
        RECT 241.400 110.800 241.800 113.100 ;
        RECT 244.100 110.800 244.600 112.100 ;
        RECT 245.800 110.800 246.200 112.100 ;
        RECT 248.600 110.800 249.000 113.000 ;
        RECT 0.200 110.200 252.600 110.800 ;
        RECT 1.400 107.900 1.800 110.200 ;
        RECT 4.100 108.900 4.600 110.200 ;
        RECT 5.800 108.900 6.200 110.200 ;
        RECT 8.600 108.000 9.000 110.200 ;
        RECT 10.200 107.900 10.600 110.200 ;
        RECT 11.800 107.900 12.200 110.200 ;
        RECT 14.200 108.000 14.600 110.200 ;
        RECT 17.000 108.900 17.400 110.200 ;
        RECT 18.600 108.900 19.100 110.200 ;
        RECT 21.400 107.900 21.800 110.200 ;
        RECT 23.000 107.900 23.400 110.200 ;
        RECT 27.000 108.300 27.400 110.200 ;
        RECT 29.400 108.000 29.800 110.200 ;
        RECT 32.200 108.900 32.600 110.200 ;
        RECT 33.800 108.900 34.300 110.200 ;
        RECT 36.600 107.900 37.000 110.200 ;
        RECT 38.200 107.900 38.600 110.200 ;
        RECT 39.800 107.900 40.200 110.200 ;
        RECT 41.400 107.900 41.800 110.200 ;
        RECT 43.000 107.900 43.400 110.200 ;
        RECT 44.600 107.900 45.000 110.200 ;
        RECT 47.000 107.900 47.400 110.200 ;
        RECT 50.200 107.700 50.600 110.200 ;
        RECT 52.800 107.500 53.200 110.200 ;
        RECT 55.000 108.000 55.400 110.200 ;
        RECT 57.800 108.900 58.200 110.200 ;
        RECT 59.400 108.900 59.900 110.200 ;
        RECT 62.200 107.900 62.600 110.200 ;
        RECT 65.400 107.900 65.800 110.200 ;
        RECT 67.800 108.300 68.200 110.200 ;
        RECT 70.200 108.300 70.600 110.200 ;
        RECT 74.200 107.900 74.600 110.200 ;
        RECT 75.800 108.000 76.200 110.200 ;
        RECT 78.600 108.900 79.000 110.200 ;
        RECT 80.200 108.900 80.700 110.200 ;
        RECT 83.000 107.900 83.400 110.200 ;
        RECT 85.400 107.900 85.800 110.200 ;
        RECT 88.100 108.900 88.600 110.200 ;
        RECT 89.800 108.900 90.200 110.200 ;
        RECT 92.600 108.000 93.000 110.200 ;
        RECT 95.000 108.300 95.400 110.200 ;
        RECT 99.000 107.900 99.400 110.200 ;
        RECT 103.000 107.900 103.400 110.200 ;
        RECT 105.400 107.900 105.800 110.200 ;
        RECT 106.200 107.900 106.600 110.200 ;
        RECT 110.200 107.900 110.600 110.200 ;
        RECT 111.000 107.900 111.400 110.200 ;
        RECT 113.400 107.900 113.800 110.200 ;
        RECT 115.000 107.900 115.400 110.200 ;
        RECT 116.600 107.900 117.000 110.200 ;
        RECT 118.200 107.900 118.600 110.200 ;
        RECT 119.800 107.900 120.200 110.200 ;
        RECT 120.600 107.900 121.000 110.200 ;
        RECT 123.000 107.900 123.400 110.200 ;
        RECT 127.000 108.300 127.400 110.200 ;
        RECT 128.600 107.900 129.000 110.200 ;
        RECT 132.600 107.900 133.000 110.200 ;
        RECT 133.400 107.900 133.800 110.200 ;
        RECT 136.600 108.000 137.000 110.200 ;
        RECT 139.400 108.900 139.800 110.200 ;
        RECT 141.000 108.900 141.500 110.200 ;
        RECT 143.800 107.900 144.200 110.200 ;
        RECT 145.400 107.900 145.800 110.200 ;
        RECT 147.000 107.900 147.400 110.200 ;
        RECT 148.600 107.900 149.000 110.200 ;
        RECT 150.200 107.900 150.600 110.200 ;
        RECT 151.800 107.900 152.200 110.200 ;
        RECT 154.200 107.900 154.600 110.200 ;
        RECT 157.400 107.700 157.800 110.200 ;
        RECT 160.000 107.500 160.400 110.200 ;
        RECT 161.400 107.900 161.800 110.200 ;
        RECT 164.400 107.900 164.800 110.200 ;
        RECT 167.000 107.900 167.400 110.200 ;
        RECT 168.600 108.300 169.000 110.200 ;
        RECT 171.000 108.900 171.400 110.200 ;
        RECT 173.100 107.900 173.500 110.200 ;
        RECT 174.200 107.900 174.600 110.200 ;
        RECT 177.400 108.000 177.800 110.200 ;
        RECT 180.200 108.900 180.600 110.200 ;
        RECT 181.800 108.900 182.300 110.200 ;
        RECT 184.600 107.900 185.000 110.200 ;
        RECT 187.800 108.300 188.200 110.200 ;
        RECT 190.200 108.000 190.600 110.200 ;
        RECT 193.000 108.900 193.400 110.200 ;
        RECT 194.600 108.900 195.100 110.200 ;
        RECT 197.400 107.900 197.800 110.200 ;
        RECT 199.000 107.900 199.400 110.200 ;
        RECT 202.000 107.900 202.400 110.200 ;
        RECT 205.200 107.500 205.600 110.200 ;
        RECT 207.800 107.700 208.200 110.200 ;
        RECT 210.200 108.300 210.600 110.200 ;
        RECT 213.400 107.900 213.800 110.200 ;
        RECT 216.100 108.900 216.600 110.200 ;
        RECT 217.800 108.900 218.200 110.200 ;
        RECT 220.600 108.000 221.000 110.200 ;
        RECT 223.800 107.900 224.200 110.200 ;
        RECT 225.400 107.700 225.800 110.200 ;
        RECT 228.000 107.500 228.400 110.200 ;
        RECT 230.200 107.900 230.600 110.200 ;
        RECT 231.800 107.900 232.200 110.200 ;
        RECT 233.400 107.900 233.800 110.200 ;
        RECT 235.000 107.900 235.400 110.200 ;
        RECT 236.600 107.900 237.000 110.200 ;
        RECT 238.200 107.900 238.600 110.200 ;
        RECT 239.000 107.900 239.400 110.200 ;
        RECT 243.000 108.300 243.400 110.200 ;
        RECT 244.600 107.900 245.000 110.200 ;
        RECT 246.200 107.900 246.600 110.200 ;
        RECT 247.800 107.900 248.200 110.200 ;
        RECT 249.400 107.900 249.800 110.200 ;
        RECT 251.000 107.900 251.400 110.200 ;
        RECT 2.200 90.800 2.600 92.700 ;
        RECT 4.600 90.800 5.000 93.100 ;
        RECT 7.300 90.800 7.800 92.100 ;
        RECT 9.000 90.800 9.400 92.100 ;
        RECT 11.800 90.800 12.200 93.000 ;
        RECT 14.000 90.800 14.400 93.500 ;
        RECT 16.600 90.800 17.000 93.300 ;
        RECT 18.200 90.800 18.600 93.100 ;
        RECT 22.200 90.800 22.600 92.700 ;
        RECT 23.800 90.800 24.200 93.100 ;
        RECT 27.800 90.800 28.200 92.700 ;
        RECT 30.200 90.800 30.600 92.700 ;
        RECT 33.400 90.800 33.800 93.100 ;
        RECT 36.100 90.800 36.600 92.100 ;
        RECT 37.800 90.800 38.200 92.100 ;
        RECT 40.600 90.800 41.000 93.000 ;
        RECT 43.800 90.800 44.200 92.700 ;
        RECT 46.200 90.800 46.600 93.300 ;
        RECT 48.800 90.800 49.200 93.500 ;
        RECT 52.600 90.800 53.000 93.100 ;
        RECT 55.300 90.800 55.800 92.100 ;
        RECT 57.000 90.800 57.400 92.100 ;
        RECT 59.800 90.800 60.200 93.000 ;
        RECT 62.200 90.800 62.600 93.300 ;
        RECT 64.800 90.800 65.200 93.500 ;
        RECT 66.200 90.800 66.600 93.100 ;
        RECT 70.200 90.800 70.600 92.700 ;
        RECT 72.600 90.800 73.000 92.700 ;
        RECT 75.800 90.800 76.200 93.100 ;
        RECT 78.500 90.800 79.000 92.100 ;
        RECT 80.200 90.800 80.600 92.100 ;
        RECT 83.000 90.800 83.400 93.000 ;
        RECT 85.400 90.800 85.800 93.100 ;
        RECT 88.100 90.800 88.600 92.100 ;
        RECT 89.800 90.800 90.200 92.100 ;
        RECT 92.600 90.800 93.000 93.000 ;
        RECT 95.800 90.800 96.200 93.100 ;
        RECT 98.200 90.800 98.600 93.100 ;
        RECT 102.200 90.800 102.600 92.700 ;
        RECT 104.600 90.800 105.000 93.100 ;
        RECT 107.300 90.800 107.800 92.100 ;
        RECT 109.000 90.800 109.400 92.100 ;
        RECT 111.800 90.800 112.200 93.000 ;
        RECT 113.400 90.800 113.800 93.100 ;
        RECT 115.800 90.800 116.200 93.100 ;
        RECT 118.800 90.800 119.200 93.500 ;
        RECT 121.400 90.800 121.800 93.300 ;
        RECT 124.100 90.800 124.500 93.000 ;
        RECT 126.200 90.800 126.600 93.100 ;
        RECT 127.800 90.800 128.200 93.100 ;
        RECT 129.400 90.800 129.800 93.100 ;
        RECT 131.000 90.800 131.400 93.100 ;
        RECT 132.600 90.800 133.000 93.100 ;
        RECT 133.400 90.800 133.800 93.100 ;
        RECT 135.800 90.800 136.200 93.100 ;
        RECT 137.400 90.800 137.800 93.100 ;
        RECT 139.000 90.800 139.400 93.100 ;
        RECT 140.600 90.800 141.000 93.100 ;
        RECT 142.200 90.800 142.600 93.100 ;
        RECT 143.800 90.800 144.200 93.100 ;
        RECT 146.200 90.800 146.600 93.100 ;
        RECT 147.800 90.800 148.200 93.100 ;
        RECT 148.600 90.800 149.000 93.100 ;
        RECT 150.200 90.800 150.600 93.100 ;
        RECT 154.000 90.800 154.400 93.500 ;
        RECT 156.600 90.800 157.000 93.300 ;
        RECT 158.200 90.800 158.600 92.100 ;
        RECT 159.800 90.800 160.200 92.100 ;
        RECT 161.400 90.800 161.800 93.000 ;
        RECT 164.200 90.800 164.600 92.100 ;
        RECT 165.800 90.800 166.300 92.100 ;
        RECT 168.600 90.800 169.000 93.100 ;
        RECT 171.000 90.800 171.400 93.100 ;
        RECT 173.700 90.800 174.200 92.100 ;
        RECT 175.400 90.800 175.800 92.100 ;
        RECT 178.200 90.800 178.600 93.000 ;
        RECT 180.600 90.800 181.000 93.000 ;
        RECT 183.400 90.800 183.800 92.100 ;
        RECT 185.000 90.800 185.500 92.100 ;
        RECT 187.800 90.800 188.200 93.100 ;
        RECT 189.400 90.800 189.800 93.100 ;
        RECT 193.400 90.800 193.800 92.700 ;
        RECT 195.800 90.800 196.200 93.000 ;
        RECT 198.600 90.800 199.000 92.100 ;
        RECT 200.200 90.800 200.700 92.100 ;
        RECT 203.000 90.800 203.400 93.100 ;
        RECT 207.800 90.800 208.200 92.700 ;
        RECT 210.200 90.800 210.600 93.300 ;
        RECT 212.800 90.800 213.200 93.500 ;
        RECT 215.800 90.800 216.200 93.100 ;
        RECT 217.400 90.800 217.800 93.000 ;
        RECT 220.200 90.800 220.600 92.100 ;
        RECT 221.800 90.800 222.300 92.100 ;
        RECT 224.600 90.800 225.000 93.100 ;
        RECT 227.800 90.800 228.200 92.700 ;
        RECT 230.200 90.800 230.600 92.700 ;
        RECT 234.200 90.800 234.600 93.100 ;
        RECT 235.800 90.800 236.200 93.100 ;
        RECT 238.500 90.800 239.000 92.100 ;
        RECT 240.200 90.800 240.600 92.100 ;
        RECT 243.000 90.800 243.400 93.000 ;
        RECT 246.200 90.800 246.600 93.100 ;
        RECT 247.800 90.800 248.200 93.300 ;
        RECT 250.400 90.800 250.800 93.500 ;
        RECT 0.200 90.200 252.600 90.800 ;
        RECT 0.600 87.900 1.000 90.200 ;
        RECT 2.200 87.900 2.600 90.200 ;
        RECT 3.800 87.900 4.200 90.200 ;
        RECT 5.400 87.900 5.800 90.200 ;
        RECT 7.000 87.900 7.400 90.200 ;
        RECT 9.400 87.900 9.800 90.200 ;
        RECT 11.000 87.900 11.400 90.200 ;
        RECT 13.700 88.900 14.200 90.200 ;
        RECT 15.400 88.900 15.800 90.200 ;
        RECT 18.200 88.000 18.600 90.200 ;
        RECT 20.600 88.000 21.000 90.200 ;
        RECT 23.400 88.900 23.800 90.200 ;
        RECT 25.000 88.900 25.500 90.200 ;
        RECT 27.800 87.900 28.200 90.200 ;
        RECT 30.000 87.500 30.400 90.200 ;
        RECT 32.600 87.700 33.000 90.200 ;
        RECT 35.800 87.900 36.200 90.200 ;
        RECT 37.400 87.700 37.800 90.200 ;
        RECT 40.000 87.500 40.400 90.200 ;
        RECT 41.400 87.900 41.800 90.200 ;
        RECT 46.200 88.000 46.600 90.200 ;
        RECT 49.000 88.900 49.400 90.200 ;
        RECT 50.600 88.900 51.100 90.200 ;
        RECT 53.400 87.900 53.800 90.200 ;
        RECT 55.800 88.300 56.200 90.200 ;
        RECT 59.800 87.900 60.200 90.200 ;
        RECT 61.200 87.500 61.600 90.200 ;
        RECT 63.800 87.700 64.200 90.200 ;
        RECT 66.200 88.000 66.600 90.200 ;
        RECT 69.000 88.900 69.400 90.200 ;
        RECT 70.600 88.900 71.100 90.200 ;
        RECT 73.400 87.900 73.800 90.200 ;
        RECT 75.000 87.900 75.400 90.200 ;
        RECT 76.600 87.900 77.000 90.200 ;
        RECT 78.200 87.900 78.600 90.200 ;
        RECT 79.800 87.900 80.200 90.200 ;
        RECT 81.400 87.900 81.800 90.200 ;
        RECT 83.800 87.900 84.200 90.200 ;
        RECT 86.200 87.900 86.600 90.200 ;
        RECT 88.600 87.900 89.000 90.200 ;
        RECT 89.400 87.900 89.800 90.200 ;
        RECT 93.400 87.900 93.800 90.200 ;
        RECT 94.200 87.900 94.600 90.200 ;
        RECT 98.200 87.900 98.600 90.200 ;
        RECT 100.600 87.900 101.000 90.200 ;
        RECT 103.000 87.900 103.400 90.200 ;
        RECT 106.200 87.900 106.600 90.200 ;
        RECT 108.900 88.900 109.400 90.200 ;
        RECT 110.600 88.900 111.000 90.200 ;
        RECT 113.400 88.000 113.800 90.200 ;
        RECT 115.800 88.300 116.200 90.200 ;
        RECT 119.800 87.900 120.200 90.200 ;
        RECT 121.400 87.700 121.800 90.200 ;
        RECT 124.000 87.500 124.400 90.200 ;
        RECT 126.200 88.300 126.600 90.200 ;
        RECT 130.200 87.900 130.600 90.200 ;
        RECT 131.800 88.000 132.200 90.200 ;
        RECT 134.600 88.900 135.000 90.200 ;
        RECT 136.200 88.900 136.700 90.200 ;
        RECT 139.000 87.900 139.400 90.200 ;
        RECT 141.400 88.000 141.800 90.200 ;
        RECT 144.200 88.900 144.600 90.200 ;
        RECT 145.800 88.900 146.300 90.200 ;
        RECT 148.600 87.900 149.000 90.200 ;
        RECT 151.800 87.900 152.200 90.200 ;
        RECT 155.800 88.300 156.200 90.200 ;
        RECT 157.700 87.900 158.100 90.200 ;
        RECT 159.800 88.900 160.200 90.200 ;
        RECT 161.200 87.500 161.600 90.200 ;
        RECT 163.800 87.700 164.200 90.200 ;
        RECT 165.400 88.900 165.800 90.200 ;
        RECT 167.000 88.900 167.400 90.200 ;
        RECT 167.800 88.900 168.200 90.200 ;
        RECT 169.900 87.900 170.300 90.200 ;
        RECT 171.800 88.000 172.200 90.200 ;
        RECT 174.600 88.900 175.000 90.200 ;
        RECT 176.200 88.900 176.700 90.200 ;
        RECT 179.000 87.900 179.400 90.200 ;
        RECT 181.200 87.500 181.600 90.200 ;
        RECT 183.800 87.700 184.200 90.200 ;
        RECT 186.200 87.700 186.600 90.200 ;
        RECT 188.800 87.500 189.200 90.200 ;
        RECT 191.000 87.700 191.400 90.200 ;
        RECT 193.600 87.500 194.000 90.200 ;
        RECT 195.000 87.900 195.400 90.200 ;
        RECT 197.400 87.900 197.800 90.200 ;
        RECT 201.400 88.300 201.800 90.200 ;
        RECT 205.400 88.000 205.800 90.200 ;
        RECT 208.200 88.900 208.600 90.200 ;
        RECT 209.800 88.900 210.300 90.200 ;
        RECT 212.600 87.900 213.000 90.200 ;
        RECT 214.800 87.500 215.200 90.200 ;
        RECT 217.400 87.700 217.800 90.200 ;
        RECT 219.000 87.900 219.400 90.200 ;
        RECT 222.200 87.700 222.600 90.200 ;
        RECT 224.800 87.500 225.200 90.200 ;
        RECT 226.200 87.900 226.600 90.200 ;
        RECT 230.200 88.300 230.600 90.200 ;
        RECT 232.600 87.900 233.000 90.200 ;
        RECT 235.300 88.900 235.800 90.200 ;
        RECT 237.000 88.900 237.400 90.200 ;
        RECT 239.800 88.000 240.200 90.200 ;
        RECT 242.200 88.300 242.600 90.200 ;
        RECT 244.600 87.900 245.000 90.200 ;
        RECT 246.200 87.900 246.600 90.200 ;
        RECT 247.800 87.900 248.200 90.200 ;
        RECT 249.400 87.900 249.800 90.200 ;
        RECT 251.000 87.900 251.400 90.200 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 4.100 70.800 4.600 72.100 ;
        RECT 5.800 70.800 6.200 72.100 ;
        RECT 8.600 70.800 9.000 73.000 ;
        RECT 11.000 70.800 11.400 73.100 ;
        RECT 12.900 70.800 13.300 73.100 ;
        RECT 15.000 70.800 15.400 72.100 ;
        RECT 15.800 70.800 16.200 72.100 ;
        RECT 17.400 70.800 17.800 72.100 ;
        RECT 19.000 70.800 19.400 72.700 ;
        RECT 23.000 70.800 23.400 73.100 ;
        RECT 24.100 70.800 24.500 73.100 ;
        RECT 26.200 70.800 26.600 72.100 ;
        RECT 27.000 70.800 27.400 72.100 ;
        RECT 28.600 70.800 29.000 72.100 ;
        RECT 30.200 70.800 30.600 72.700 ;
        RECT 34.200 70.800 34.600 73.100 ;
        RECT 35.800 70.800 36.200 73.100 ;
        RECT 38.500 70.800 39.000 72.100 ;
        RECT 40.200 70.800 40.600 72.100 ;
        RECT 43.000 70.800 43.400 73.000 ;
        RECT 45.400 70.800 45.800 73.300 ;
        RECT 48.000 70.800 48.400 73.500 ;
        RECT 51.000 70.800 51.400 72.100 ;
        RECT 52.600 70.800 53.000 72.100 ;
        RECT 53.400 70.800 53.800 72.100 ;
        RECT 55.500 70.800 55.900 73.100 ;
        RECT 57.400 70.800 57.800 73.000 ;
        RECT 60.200 70.800 60.600 72.100 ;
        RECT 61.800 70.800 62.300 72.100 ;
        RECT 64.600 70.800 65.000 73.100 ;
        RECT 66.200 70.800 66.600 73.100 ;
        RECT 67.800 70.800 68.200 73.100 ;
        RECT 70.200 70.800 70.600 73.100 ;
        RECT 71.800 70.800 72.200 73.100 ;
        RECT 73.400 70.800 73.800 72.700 ;
        RECT 77.400 70.800 77.800 73.100 ;
        RECT 79.000 70.800 79.400 73.100 ;
        RECT 81.700 70.800 82.200 72.100 ;
        RECT 83.400 70.800 83.800 72.100 ;
        RECT 86.200 70.800 86.600 73.000 ;
        RECT 88.000 70.800 88.400 73.100 ;
        RECT 91.000 70.800 91.400 73.100 ;
        RECT 91.800 70.800 92.200 73.100 ;
        RECT 95.800 70.800 96.200 73.100 ;
        RECT 96.600 70.800 97.000 73.100 ;
        RECT 102.200 70.800 102.600 72.700 ;
        RECT 105.100 70.800 105.500 73.000 ;
        RECT 107.000 70.800 107.400 73.100 ;
        RECT 109.400 70.800 109.800 72.100 ;
        RECT 111.000 70.800 111.400 72.100 ;
        RECT 111.800 70.800 112.200 72.100 ;
        RECT 113.400 70.800 113.800 72.100 ;
        RECT 114.800 70.800 115.200 73.500 ;
        RECT 117.400 70.800 117.800 73.300 ;
        RECT 119.000 70.800 119.400 73.100 ;
        RECT 121.400 70.800 121.800 72.100 ;
        RECT 123.000 70.800 123.400 72.100 ;
        RECT 124.400 70.800 124.800 73.500 ;
        RECT 127.000 70.800 127.400 73.300 ;
        RECT 128.600 70.800 129.000 73.100 ;
        RECT 131.600 70.800 132.000 73.100 ;
        RECT 133.400 70.800 133.800 73.300 ;
        RECT 136.000 70.800 136.400 73.500 ;
        RECT 138.700 70.800 139.100 73.000 ;
        RECT 140.600 70.800 141.000 73.100 ;
        RECT 143.800 70.800 144.200 73.100 ;
        RECT 145.400 70.800 145.800 73.100 ;
        RECT 148.600 70.800 149.000 73.000 ;
        RECT 151.400 70.800 151.800 72.100 ;
        RECT 153.000 70.800 153.500 72.100 ;
        RECT 155.800 70.800 156.200 73.100 ;
        RECT 159.000 70.800 159.400 73.100 ;
        RECT 160.100 70.800 160.500 73.100 ;
        RECT 162.200 70.800 162.600 72.100 ;
        RECT 163.000 70.800 163.400 73.100 ;
        RECT 164.600 70.800 165.000 73.100 ;
        RECT 167.000 70.800 167.400 72.700 ;
        RECT 171.000 70.800 171.400 73.100 ;
        RECT 172.600 70.800 173.000 73.100 ;
        RECT 175.300 70.800 175.800 72.100 ;
        RECT 177.000 70.800 177.400 72.100 ;
        RECT 179.800 70.800 180.200 73.000 ;
        RECT 183.000 70.800 183.400 72.700 ;
        RECT 185.400 70.800 185.800 73.300 ;
        RECT 188.000 70.800 188.400 73.500 ;
        RECT 190.200 70.800 190.600 73.300 ;
        RECT 192.800 70.800 193.200 73.500 ;
        RECT 195.000 70.800 195.400 72.700 ;
        RECT 199.000 70.800 199.400 73.100 ;
        RECT 199.800 70.800 200.200 73.100 ;
        RECT 203.800 70.800 204.200 73.100 ;
        RECT 206.800 70.800 207.200 73.100 ;
        RECT 208.600 70.800 209.000 73.300 ;
        RECT 211.200 70.800 211.600 73.500 ;
        RECT 212.600 70.800 213.000 73.100 ;
        RECT 215.000 70.800 215.400 73.100 ;
        RECT 218.200 70.800 218.600 72.700 ;
        RECT 221.200 70.800 221.600 73.500 ;
        RECT 223.800 70.800 224.200 73.300 ;
        RECT 226.200 70.800 226.600 73.000 ;
        RECT 229.000 70.800 229.400 72.100 ;
        RECT 230.600 70.800 231.100 72.100 ;
        RECT 233.400 70.800 233.800 73.100 ;
        RECT 235.000 70.800 235.400 73.100 ;
        RECT 236.600 70.800 237.000 73.100 ;
        RECT 238.200 70.800 238.600 73.100 ;
        RECT 239.800 70.800 240.200 73.100 ;
        RECT 241.400 70.800 241.800 73.100 ;
        RECT 242.200 70.800 242.600 72.100 ;
        RECT 243.800 70.800 244.200 72.100 ;
        RECT 244.600 70.800 245.000 72.100 ;
        RECT 246.700 70.800 247.100 73.100 ;
        RECT 249.400 70.800 249.800 72.700 ;
        RECT 0.200 70.200 252.600 70.800 ;
        RECT 0.600 67.900 1.000 70.200 ;
        RECT 4.600 68.300 5.000 70.200 ;
        RECT 6.800 67.500 7.200 70.200 ;
        RECT 9.400 67.700 9.800 70.200 ;
        RECT 11.800 67.900 12.200 70.200 ;
        RECT 14.500 68.900 15.000 70.200 ;
        RECT 16.200 68.900 16.600 70.200 ;
        RECT 19.000 68.000 19.400 70.200 ;
        RECT 21.400 67.900 21.800 70.200 ;
        RECT 24.100 68.900 24.600 70.200 ;
        RECT 25.800 68.900 26.200 70.200 ;
        RECT 28.600 68.000 29.000 70.200 ;
        RECT 31.000 67.700 31.400 70.200 ;
        RECT 33.600 67.500 34.000 70.200 ;
        RECT 35.800 67.700 36.200 70.200 ;
        RECT 38.400 67.500 38.800 70.200 ;
        RECT 40.400 67.500 40.800 70.200 ;
        RECT 43.000 67.700 43.400 70.200 ;
        RECT 45.200 67.500 45.600 70.200 ;
        RECT 47.800 67.700 48.200 70.200 ;
        RECT 51.000 67.900 51.400 70.200 ;
        RECT 54.000 67.900 54.400 70.200 ;
        RECT 55.200 67.900 55.600 70.200 ;
        RECT 58.200 67.900 58.600 70.200 ;
        RECT 59.000 67.900 59.400 70.200 ;
        RECT 62.200 68.300 62.600 70.200 ;
        RECT 64.600 67.900 65.000 70.200 ;
        RECT 67.600 67.900 68.000 70.200 ;
        RECT 68.600 67.900 69.000 70.200 ;
        RECT 71.600 67.500 72.000 70.200 ;
        RECT 74.200 67.700 74.600 70.200 ;
        RECT 76.000 67.900 76.400 70.200 ;
        RECT 79.000 67.900 79.400 70.200 ;
        RECT 81.400 68.300 81.800 70.200 ;
        RECT 83.000 67.900 83.400 70.200 ;
        RECT 86.700 68.000 87.100 70.200 ;
        RECT 88.800 67.900 89.200 70.200 ;
        RECT 91.800 67.900 92.200 70.200 ;
        RECT 92.600 67.900 93.000 70.200 ;
        RECT 97.400 68.000 97.800 70.200 ;
        RECT 100.200 68.900 100.600 70.200 ;
        RECT 101.800 68.900 102.300 70.200 ;
        RECT 104.600 67.900 105.000 70.200 ;
        RECT 106.200 68.900 106.600 70.200 ;
        RECT 107.800 67.900 108.200 70.200 ;
        RECT 110.200 67.900 110.600 70.200 ;
        RECT 114.200 67.900 114.600 70.200 ;
        RECT 115.000 67.900 115.400 70.200 ;
        RECT 118.000 67.900 118.400 70.200 ;
        RECT 119.800 68.000 120.200 70.200 ;
        RECT 122.600 68.900 123.000 70.200 ;
        RECT 124.200 68.900 124.700 70.200 ;
        RECT 127.000 67.900 127.400 70.200 ;
        RECT 128.600 67.900 129.000 70.200 ;
        RECT 132.600 68.300 133.000 70.200 ;
        RECT 134.500 67.900 134.900 70.200 ;
        RECT 136.600 68.900 137.000 70.200 ;
        RECT 137.400 68.900 137.800 70.200 ;
        RECT 139.000 68.900 139.400 70.200 ;
        RECT 140.600 67.900 141.000 70.200 ;
        RECT 143.300 68.900 143.800 70.200 ;
        RECT 145.000 68.900 145.400 70.200 ;
        RECT 147.800 68.000 148.200 70.200 ;
        RECT 151.800 67.900 152.200 70.200 ;
        RECT 154.500 68.900 155.000 70.200 ;
        RECT 156.200 68.900 156.600 70.200 ;
        RECT 159.000 68.000 159.400 70.200 ;
        RECT 160.600 67.900 161.000 70.200 ;
        RECT 164.600 68.300 165.000 70.200 ;
        RECT 166.200 67.900 166.600 70.200 ;
        RECT 169.200 67.900 169.600 70.200 ;
        RECT 171.000 67.700 171.400 70.200 ;
        RECT 173.600 67.500 174.000 70.200 ;
        RECT 175.800 67.900 176.200 70.200 ;
        RECT 178.500 68.900 179.000 70.200 ;
        RECT 180.200 68.900 180.600 70.200 ;
        RECT 183.000 68.000 183.400 70.200 ;
        RECT 186.200 67.900 186.600 70.200 ;
        RECT 187.600 67.500 188.000 70.200 ;
        RECT 190.200 67.700 190.600 70.200 ;
        RECT 191.800 67.900 192.200 70.200 ;
        RECT 194.800 67.900 195.200 70.200 ;
        RECT 196.400 67.500 196.800 70.200 ;
        RECT 199.000 67.700 199.400 70.200 ;
        RECT 202.200 67.900 202.600 70.200 ;
        RECT 205.200 67.900 205.600 70.200 ;
        RECT 206.200 67.900 206.600 70.200 ;
        RECT 207.800 67.900 208.200 70.200 ;
        RECT 210.200 67.900 210.600 70.200 ;
        RECT 211.800 67.900 212.200 70.200 ;
        RECT 213.400 68.300 213.800 70.200 ;
        RECT 216.600 68.000 217.000 70.200 ;
        RECT 219.400 68.900 219.800 70.200 ;
        RECT 221.000 68.900 221.500 70.200 ;
        RECT 223.800 67.900 224.200 70.200 ;
        RECT 226.000 67.500 226.400 70.200 ;
        RECT 228.600 67.700 229.000 70.200 ;
        RECT 230.200 67.900 230.600 70.200 ;
        RECT 233.400 68.000 233.800 70.200 ;
        RECT 236.200 68.900 236.600 70.200 ;
        RECT 237.800 68.900 238.300 70.200 ;
        RECT 240.600 67.900 241.000 70.200 ;
        RECT 243.000 67.900 243.400 70.200 ;
        RECT 245.700 68.900 246.200 70.200 ;
        RECT 247.400 68.900 247.800 70.200 ;
        RECT 250.200 68.000 250.600 70.200 ;
        RECT 0.600 50.800 1.000 53.100 ;
        RECT 4.600 50.800 5.000 52.700 ;
        RECT 7.000 50.800 7.400 53.100 ;
        RECT 9.700 50.800 10.200 52.100 ;
        RECT 11.400 50.800 11.800 52.100 ;
        RECT 14.200 50.800 14.600 53.000 ;
        RECT 16.600 50.800 17.000 53.100 ;
        RECT 19.300 50.800 19.800 52.100 ;
        RECT 21.000 50.800 21.400 52.100 ;
        RECT 23.800 50.800 24.200 53.000 ;
        RECT 25.400 50.800 25.800 53.100 ;
        RECT 29.400 50.800 29.800 52.700 ;
        RECT 31.800 50.800 32.200 53.000 ;
        RECT 34.600 50.800 35.000 52.100 ;
        RECT 36.200 50.800 36.700 52.100 ;
        RECT 39.000 50.800 39.400 53.100 ;
        RECT 41.200 50.800 41.600 53.500 ;
        RECT 43.800 50.800 44.200 53.300 ;
        RECT 46.200 50.800 46.600 53.300 ;
        RECT 48.800 50.800 49.200 53.500 ;
        RECT 52.600 50.800 53.000 53.300 ;
        RECT 55.200 50.800 55.600 53.500 ;
        RECT 56.900 50.800 57.300 53.100 ;
        RECT 59.000 50.800 59.400 52.100 ;
        RECT 59.800 50.800 60.200 52.100 ;
        RECT 61.900 50.800 62.300 53.100 ;
        RECT 63.800 50.800 64.200 52.700 ;
        RECT 67.800 50.800 68.200 53.100 ;
        RECT 69.400 50.800 69.800 53.100 ;
        RECT 72.100 50.800 72.600 52.100 ;
        RECT 73.800 50.800 74.200 52.100 ;
        RECT 76.600 50.800 77.000 53.000 ;
        RECT 78.800 50.800 79.200 53.500 ;
        RECT 81.400 50.800 81.800 53.300 ;
        RECT 83.600 50.800 84.000 53.500 ;
        RECT 86.200 50.800 86.600 53.300 ;
        RECT 88.600 50.800 89.000 53.300 ;
        RECT 91.200 50.800 91.600 53.500 ;
        RECT 93.400 50.800 93.800 53.300 ;
        RECT 96.000 50.800 96.400 53.500 ;
        RECT 99.800 50.800 100.200 53.000 ;
        RECT 102.600 50.800 103.000 52.100 ;
        RECT 104.200 50.800 104.700 52.100 ;
        RECT 107.000 50.800 107.400 53.100 ;
        RECT 108.600 50.800 109.000 53.100 ;
        RECT 112.600 50.800 113.000 52.700 ;
        RECT 114.200 50.800 114.600 52.100 ;
        RECT 115.800 50.800 116.200 52.100 ;
        RECT 118.200 50.800 118.600 53.100 ;
        RECT 119.800 50.800 120.200 52.100 ;
        RECT 121.400 50.800 121.800 53.300 ;
        RECT 124.000 50.800 124.400 53.500 ;
        RECT 127.000 50.800 127.400 53.100 ;
        RECT 129.400 50.800 129.800 52.700 ;
        RECT 131.800 50.800 132.200 53.100 ;
        RECT 134.500 50.800 135.000 52.100 ;
        RECT 136.200 50.800 136.600 52.100 ;
        RECT 139.000 50.800 139.400 53.000 ;
        RECT 140.900 50.800 141.300 53.100 ;
        RECT 143.000 50.800 143.400 52.100 ;
        RECT 143.800 50.800 144.200 52.100 ;
        RECT 145.400 50.800 145.800 52.100 ;
        RECT 146.800 50.800 147.200 53.500 ;
        RECT 149.400 50.800 149.800 53.300 ;
        RECT 153.400 50.800 153.800 52.700 ;
        RECT 157.400 50.800 157.800 53.100 ;
        RECT 159.000 50.800 159.400 53.100 ;
        RECT 161.700 50.800 162.200 52.100 ;
        RECT 163.400 50.800 163.800 52.100 ;
        RECT 166.200 50.800 166.600 53.000 ;
        RECT 168.600 50.800 169.000 53.000 ;
        RECT 171.400 50.800 171.800 52.100 ;
        RECT 173.000 50.800 173.500 52.100 ;
        RECT 175.800 50.800 176.200 53.100 ;
        RECT 178.200 50.800 178.600 53.100 ;
        RECT 180.900 50.800 181.400 52.100 ;
        RECT 182.600 50.800 183.000 52.100 ;
        RECT 185.400 50.800 185.800 53.000 ;
        RECT 187.000 50.800 187.400 52.100 ;
        RECT 189.100 50.800 189.500 53.100 ;
        RECT 190.200 50.800 190.600 52.100 ;
        RECT 191.800 50.800 192.200 52.100 ;
        RECT 193.200 50.800 193.600 53.500 ;
        RECT 195.800 50.800 196.200 53.300 ;
        RECT 197.400 50.800 197.800 52.100 ;
        RECT 199.000 50.800 199.400 52.100 ;
        RECT 199.800 50.800 200.200 52.100 ;
        RECT 201.900 50.800 202.300 53.100 ;
        RECT 205.400 50.800 205.800 53.100 ;
        RECT 207.000 50.800 207.400 53.100 ;
        RECT 207.800 50.800 208.200 53.100 ;
        RECT 209.400 50.800 209.800 53.100 ;
        RECT 211.000 50.800 211.400 53.100 ;
        RECT 212.600 50.800 213.000 53.100 ;
        RECT 214.200 50.800 214.600 53.100 ;
        RECT 215.800 50.800 216.200 53.000 ;
        RECT 218.600 50.800 219.000 52.100 ;
        RECT 220.200 50.800 220.700 52.100 ;
        RECT 223.000 50.800 223.400 53.100 ;
        RECT 224.600 50.800 225.000 52.100 ;
        RECT 226.700 50.800 227.100 53.100 ;
        RECT 228.600 50.800 229.000 53.000 ;
        RECT 231.400 50.800 231.800 52.100 ;
        RECT 233.000 50.800 233.500 52.100 ;
        RECT 235.800 50.800 236.200 53.100 ;
        RECT 239.000 50.800 239.400 52.700 ;
        RECT 241.400 50.800 241.800 53.000 ;
        RECT 244.200 50.800 244.600 52.100 ;
        RECT 245.800 50.800 246.300 52.100 ;
        RECT 248.600 50.800 249.000 53.100 ;
        RECT 0.200 50.200 252.600 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 3.000 47.900 3.400 50.200 ;
        RECT 4.600 47.900 5.000 50.200 ;
        RECT 6.200 47.900 6.600 50.200 ;
        RECT 7.800 47.900 8.200 50.200 ;
        RECT 9.400 47.900 9.800 50.200 ;
        RECT 10.200 47.900 10.600 50.200 ;
        RECT 14.200 48.300 14.600 50.200 ;
        RECT 16.600 47.900 17.000 50.200 ;
        RECT 19.300 48.900 19.800 50.200 ;
        RECT 21.000 48.900 21.400 50.200 ;
        RECT 23.800 48.000 24.200 50.200 ;
        RECT 26.000 47.500 26.400 50.200 ;
        RECT 28.600 47.700 29.000 50.200 ;
        RECT 30.200 47.900 30.600 50.200 ;
        RECT 34.200 48.300 34.600 50.200 ;
        RECT 36.600 48.000 37.000 50.200 ;
        RECT 39.400 48.900 39.800 50.200 ;
        RECT 41.000 48.900 41.500 50.200 ;
        RECT 43.800 47.900 44.200 50.200 ;
        RECT 47.000 47.900 47.400 50.200 ;
        RECT 49.400 47.900 49.800 50.200 ;
        RECT 52.600 48.000 53.000 50.200 ;
        RECT 55.400 48.900 55.800 50.200 ;
        RECT 57.000 48.900 57.500 50.200 ;
        RECT 59.800 47.900 60.200 50.200 ;
        RECT 62.200 47.900 62.600 50.200 ;
        RECT 64.900 48.900 65.400 50.200 ;
        RECT 66.600 48.900 67.000 50.200 ;
        RECT 69.400 48.000 69.800 50.200 ;
        RECT 71.800 48.300 72.200 50.200 ;
        RECT 75.800 47.900 76.200 50.200 ;
        RECT 77.400 47.900 77.800 50.200 ;
        RECT 80.100 48.900 80.600 50.200 ;
        RECT 81.800 48.900 82.200 50.200 ;
        RECT 84.600 48.000 85.000 50.200 ;
        RECT 86.200 47.900 86.600 50.200 ;
        RECT 90.200 48.300 90.600 50.200 ;
        RECT 92.600 48.000 93.000 50.200 ;
        RECT 95.400 48.900 95.800 50.200 ;
        RECT 97.000 48.900 97.500 50.200 ;
        RECT 99.800 47.900 100.200 50.200 ;
        RECT 103.000 47.900 103.400 50.200 ;
        RECT 107.000 48.300 107.400 50.200 ;
        RECT 108.600 47.900 109.000 50.200 ;
        RECT 110.200 47.900 110.600 50.200 ;
        RECT 111.800 47.900 112.200 50.200 ;
        RECT 113.400 47.900 113.800 50.200 ;
        RECT 115.000 47.900 115.400 50.200 ;
        RECT 116.600 47.900 117.000 50.200 ;
        RECT 118.200 47.900 118.600 50.200 ;
        RECT 119.800 48.300 120.200 50.200 ;
        RECT 123.800 47.900 124.200 50.200 ;
        RECT 125.400 48.000 125.800 50.200 ;
        RECT 128.200 48.900 128.600 50.200 ;
        RECT 129.800 48.900 130.300 50.200 ;
        RECT 132.600 47.900 133.000 50.200 ;
        RECT 135.000 47.900 135.400 50.200 ;
        RECT 136.600 47.900 137.000 50.200 ;
        RECT 137.400 47.900 137.800 50.200 ;
        RECT 140.600 47.900 141.000 50.200 ;
        RECT 143.300 48.900 143.800 50.200 ;
        RECT 145.000 48.900 145.400 50.200 ;
        RECT 147.800 48.000 148.200 50.200 ;
        RECT 151.600 47.500 152.000 50.200 ;
        RECT 154.200 47.700 154.600 50.200 ;
        RECT 155.800 47.900 156.200 50.200 ;
        RECT 159.800 48.300 160.200 50.200 ;
        RECT 161.400 47.900 161.800 50.200 ;
        RECT 163.000 47.900 163.400 50.200 ;
        RECT 164.600 47.900 165.000 50.200 ;
        RECT 166.200 47.900 166.600 50.200 ;
        RECT 167.800 47.900 168.200 50.200 ;
        RECT 169.400 47.900 169.800 50.200 ;
        RECT 171.800 47.900 172.200 50.200 ;
        RECT 173.400 47.900 173.800 50.200 ;
        RECT 175.000 47.900 175.400 50.200 ;
        RECT 176.600 47.900 177.000 50.200 ;
        RECT 177.400 47.900 177.800 50.200 ;
        RECT 179.000 47.900 179.400 50.200 ;
        RECT 180.600 47.900 181.000 50.200 ;
        RECT 182.200 47.900 182.600 50.200 ;
        RECT 183.800 47.900 184.200 50.200 ;
        RECT 185.400 47.900 185.800 50.200 ;
        RECT 187.000 47.900 187.400 50.200 ;
        RECT 188.600 47.700 189.000 50.200 ;
        RECT 191.200 47.500 191.600 50.200 ;
        RECT 193.400 48.000 193.800 50.200 ;
        RECT 196.200 48.900 196.600 50.200 ;
        RECT 197.800 48.900 198.300 50.200 ;
        RECT 200.600 47.900 201.000 50.200 ;
        RECT 204.400 47.500 204.800 50.200 ;
        RECT 207.000 47.700 207.400 50.200 ;
        RECT 209.400 48.000 209.800 50.200 ;
        RECT 212.200 48.900 212.600 50.200 ;
        RECT 213.800 48.900 214.300 50.200 ;
        RECT 216.600 47.900 217.000 50.200 ;
        RECT 218.200 47.900 218.600 50.200 ;
        RECT 222.200 48.300 222.600 50.200 ;
        RECT 223.800 48.900 224.200 50.200 ;
        RECT 225.400 48.900 225.800 50.200 ;
        RECT 227.000 47.700 227.400 50.200 ;
        RECT 229.600 47.500 230.000 50.200 ;
        RECT 231.600 47.500 232.000 50.200 ;
        RECT 234.200 47.700 234.600 50.200 ;
        RECT 236.600 48.300 237.000 50.200 ;
        RECT 240.600 47.900 241.000 50.200 ;
        RECT 242.200 47.900 242.600 50.200 ;
        RECT 244.900 48.900 245.400 50.200 ;
        RECT 246.600 48.900 247.000 50.200 ;
        RECT 249.400 48.000 249.800 50.200 ;
        RECT 1.400 30.800 1.800 33.100 ;
        RECT 4.100 30.800 4.600 32.100 ;
        RECT 5.800 30.800 6.200 32.100 ;
        RECT 8.600 30.800 9.000 33.000 ;
        RECT 10.800 30.800 11.200 33.500 ;
        RECT 13.400 30.800 13.800 33.300 ;
        RECT 15.800 30.800 16.200 32.700 ;
        RECT 19.800 30.800 20.200 33.100 ;
        RECT 21.400 30.800 21.800 33.100 ;
        RECT 24.100 30.800 24.600 32.100 ;
        RECT 25.800 30.800 26.200 32.100 ;
        RECT 28.600 30.800 29.000 33.000 ;
        RECT 31.000 30.800 31.400 33.300 ;
        RECT 33.600 30.800 34.000 33.500 ;
        RECT 35.600 30.800 36.000 33.500 ;
        RECT 38.200 30.800 38.600 33.300 ;
        RECT 39.800 30.800 40.200 33.100 ;
        RECT 43.800 30.800 44.200 32.700 ;
        RECT 45.400 30.800 45.800 33.100 ;
        RECT 47.000 30.800 47.400 33.100 ;
        RECT 50.200 30.800 50.600 33.100 ;
        RECT 54.200 30.800 54.600 32.700 ;
        RECT 56.600 30.800 57.000 33.300 ;
        RECT 59.200 30.800 59.600 33.500 ;
        RECT 61.200 30.800 61.600 33.500 ;
        RECT 63.800 30.800 64.200 33.300 ;
        RECT 66.000 30.800 66.400 33.500 ;
        RECT 68.600 30.800 69.000 33.300 ;
        RECT 70.200 30.800 70.600 33.100 ;
        RECT 71.800 30.800 72.200 33.100 ;
        RECT 74.200 30.800 74.600 33.100 ;
        RECT 76.900 30.800 77.400 32.100 ;
        RECT 78.600 30.800 79.000 32.100 ;
        RECT 81.400 30.800 81.800 33.000 ;
        RECT 83.000 30.800 83.400 33.100 ;
        RECT 85.700 30.800 86.100 33.100 ;
        RECT 87.800 30.800 88.200 32.100 ;
        RECT 88.600 30.800 89.000 32.100 ;
        RECT 90.200 30.800 90.600 32.100 ;
        RECT 91.600 30.800 92.000 33.500 ;
        RECT 94.200 30.800 94.600 33.300 ;
        RECT 95.800 30.800 96.200 33.100 ;
        RECT 97.400 30.800 97.800 33.100 ;
        RECT 101.200 30.800 101.600 33.500 ;
        RECT 103.800 30.800 104.200 33.300 ;
        RECT 106.200 30.800 106.600 32.700 ;
        RECT 110.200 30.800 110.600 33.100 ;
        RECT 111.800 30.800 112.200 33.100 ;
        RECT 114.500 30.800 115.000 32.100 ;
        RECT 116.200 30.800 116.600 32.100 ;
        RECT 119.000 30.800 119.400 33.000 ;
        RECT 121.400 30.800 121.800 33.300 ;
        RECT 124.000 30.800 124.400 33.500 ;
        RECT 126.000 30.800 126.400 33.500 ;
        RECT 128.600 30.800 129.000 33.300 ;
        RECT 131.000 30.800 131.400 33.000 ;
        RECT 133.800 30.800 134.200 32.100 ;
        RECT 135.400 30.800 135.900 32.100 ;
        RECT 138.200 30.800 138.600 33.100 ;
        RECT 139.800 30.800 140.200 33.100 ;
        RECT 142.200 30.800 142.600 33.100 ;
        RECT 143.800 30.800 144.200 33.100 ;
        RECT 145.200 30.800 145.600 33.500 ;
        RECT 147.800 30.800 148.200 33.300 ;
        RECT 151.800 30.800 152.200 33.000 ;
        RECT 154.600 30.800 155.000 32.100 ;
        RECT 156.200 30.800 156.700 32.100 ;
        RECT 159.000 30.800 159.400 33.100 ;
        RECT 160.600 30.800 161.000 33.100 ;
        RECT 162.200 30.800 162.600 33.100 ;
        RECT 164.600 30.800 165.000 33.100 ;
        RECT 166.200 30.800 166.600 33.100 ;
        RECT 168.600 30.800 169.000 33.100 ;
        RECT 170.200 30.800 170.600 33.300 ;
        RECT 172.800 30.800 173.200 33.500 ;
        RECT 175.000 30.800 175.400 33.100 ;
        RECT 176.600 30.800 177.000 33.100 ;
        RECT 178.200 30.800 178.600 33.300 ;
        RECT 180.800 30.800 181.200 33.500 ;
        RECT 182.200 30.800 182.600 33.100 ;
        RECT 186.200 30.800 186.600 32.700 ;
        RECT 188.600 30.800 189.000 33.000 ;
        RECT 191.400 30.800 191.800 32.100 ;
        RECT 193.000 30.800 193.500 32.100 ;
        RECT 195.800 30.800 196.200 33.100 ;
        RECT 198.200 30.800 198.600 33.300 ;
        RECT 200.800 30.800 201.200 33.500 ;
        RECT 204.600 30.800 205.000 33.000 ;
        RECT 207.400 30.800 207.800 32.100 ;
        RECT 209.000 30.800 209.500 32.100 ;
        RECT 211.800 30.800 212.200 33.100 ;
        RECT 215.000 30.800 215.400 33.100 ;
        RECT 216.600 30.800 217.000 33.300 ;
        RECT 219.200 30.800 219.600 33.500 ;
        RECT 221.400 30.800 221.800 32.700 ;
        RECT 225.400 30.800 225.800 33.100 ;
        RECT 226.800 30.800 227.200 33.500 ;
        RECT 229.400 30.800 229.800 33.300 ;
        RECT 231.000 30.800 231.400 32.100 ;
        RECT 232.600 30.800 233.000 32.100 ;
        RECT 233.400 30.800 233.800 32.100 ;
        RECT 235.500 30.800 235.900 33.100 ;
        RECT 237.400 30.800 237.800 32.700 ;
        RECT 241.400 30.800 241.800 33.100 ;
        RECT 243.000 30.800 243.400 33.100 ;
        RECT 245.700 30.800 246.200 32.100 ;
        RECT 247.400 30.800 247.800 32.100 ;
        RECT 250.200 30.800 250.600 33.000 ;
        RECT 0.200 30.200 252.600 30.800 ;
        RECT 0.600 27.900 1.000 30.200 ;
        RECT 4.600 28.300 5.000 30.200 ;
        RECT 6.200 27.900 6.600 30.200 ;
        RECT 10.200 28.300 10.600 30.200 ;
        RECT 12.600 27.900 13.000 30.200 ;
        RECT 15.300 28.900 15.800 30.200 ;
        RECT 17.000 28.900 17.400 30.200 ;
        RECT 19.800 28.000 20.200 30.200 ;
        RECT 22.200 27.900 22.600 30.200 ;
        RECT 24.900 28.900 25.400 30.200 ;
        RECT 26.600 28.900 27.000 30.200 ;
        RECT 29.400 28.000 29.800 30.200 ;
        RECT 31.800 28.000 32.200 30.200 ;
        RECT 34.600 28.900 35.000 30.200 ;
        RECT 36.200 28.900 36.700 30.200 ;
        RECT 39.000 27.900 39.400 30.200 ;
        RECT 41.400 28.000 41.800 30.200 ;
        RECT 44.200 28.900 44.600 30.200 ;
        RECT 45.800 28.900 46.300 30.200 ;
        RECT 48.600 27.900 49.000 30.200 ;
        RECT 52.600 27.700 53.000 30.200 ;
        RECT 55.200 27.500 55.600 30.200 ;
        RECT 57.400 28.300 57.800 30.200 ;
        RECT 61.400 27.900 61.800 30.200 ;
        RECT 63.000 27.900 63.400 30.200 ;
        RECT 65.700 28.900 66.200 30.200 ;
        RECT 67.400 28.900 67.800 30.200 ;
        RECT 70.200 28.000 70.600 30.200 ;
        RECT 72.400 27.500 72.800 30.200 ;
        RECT 75.000 27.700 75.400 30.200 ;
        RECT 76.600 27.900 77.000 30.200 ;
        RECT 80.600 28.300 81.000 30.200 ;
        RECT 83.000 28.300 83.400 30.200 ;
        RECT 86.200 28.000 86.600 30.200 ;
        RECT 89.000 28.900 89.400 30.200 ;
        RECT 90.600 28.900 91.100 30.200 ;
        RECT 93.400 27.900 93.800 30.200 ;
        RECT 97.400 28.000 97.800 30.200 ;
        RECT 100.200 28.900 100.600 30.200 ;
        RECT 101.800 28.900 102.300 30.200 ;
        RECT 104.600 27.900 105.000 30.200 ;
        RECT 106.200 27.900 106.600 30.200 ;
        RECT 110.200 28.300 110.600 30.200 ;
        RECT 112.600 28.300 113.000 30.200 ;
        RECT 116.600 27.900 117.000 30.200 ;
        RECT 118.200 27.900 118.600 30.200 ;
        RECT 120.900 28.900 121.400 30.200 ;
        RECT 122.600 28.900 123.000 30.200 ;
        RECT 125.400 28.000 125.800 30.200 ;
        RECT 127.800 28.300 128.200 30.200 ;
        RECT 131.800 27.900 132.200 30.200 ;
        RECT 133.400 27.900 133.800 30.200 ;
        RECT 136.100 28.900 136.600 30.200 ;
        RECT 137.800 28.900 138.200 30.200 ;
        RECT 140.600 28.000 141.000 30.200 ;
        RECT 143.800 28.300 144.200 30.200 ;
        RECT 146.200 27.700 146.600 30.200 ;
        RECT 148.800 27.500 149.200 30.200 ;
        RECT 152.600 27.700 153.000 30.200 ;
        RECT 155.200 27.500 155.600 30.200 ;
        RECT 157.400 27.900 157.800 30.200 ;
        RECT 159.000 27.900 159.400 30.200 ;
        RECT 159.800 27.900 160.200 30.200 ;
        RECT 163.800 28.300 164.200 30.200 ;
        RECT 166.200 27.900 166.600 30.200 ;
        RECT 167.800 27.900 168.200 30.200 ;
        RECT 170.200 28.300 170.600 30.200 ;
        RECT 172.600 28.000 173.000 30.200 ;
        RECT 175.400 28.900 175.800 30.200 ;
        RECT 177.000 28.900 177.500 30.200 ;
        RECT 179.800 27.900 180.200 30.200 ;
        RECT 181.400 27.900 181.800 30.200 ;
        RECT 185.400 28.300 185.800 30.200 ;
        RECT 187.800 28.000 188.200 30.200 ;
        RECT 190.600 28.900 191.000 30.200 ;
        RECT 192.200 28.900 192.700 30.200 ;
        RECT 195.000 27.900 195.400 30.200 ;
        RECT 197.400 27.700 197.800 30.200 ;
        RECT 200.000 27.500 200.400 30.200 ;
        RECT 203.800 27.900 204.200 30.200 ;
        RECT 205.400 27.900 205.800 30.200 ;
        RECT 206.200 27.900 206.600 30.200 ;
        RECT 210.200 28.300 210.600 30.200 ;
        RECT 212.600 28.300 213.000 30.200 ;
        RECT 215.000 27.900 215.400 30.200 ;
        RECT 216.600 27.900 217.000 30.200 ;
        RECT 219.000 28.000 219.400 30.200 ;
        RECT 221.800 28.900 222.200 30.200 ;
        RECT 223.400 28.900 223.900 30.200 ;
        RECT 226.200 27.900 226.600 30.200 ;
        RECT 227.800 27.900 228.200 30.200 ;
        RECT 231.000 28.000 231.400 30.200 ;
        RECT 233.800 28.900 234.200 30.200 ;
        RECT 235.400 28.900 235.900 30.200 ;
        RECT 238.200 27.900 238.600 30.200 ;
        RECT 240.600 28.000 241.000 30.200 ;
        RECT 243.400 28.900 243.800 30.200 ;
        RECT 245.000 28.900 245.500 30.200 ;
        RECT 247.800 27.900 248.200 30.200 ;
        RECT 250.200 28.300 250.600 30.200 ;
        RECT 1.400 10.800 1.800 13.000 ;
        RECT 4.200 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.300 12.100 ;
        RECT 8.600 10.800 9.000 13.100 ;
        RECT 10.200 10.800 10.600 13.100 ;
        RECT 14.200 10.800 14.600 12.700 ;
        RECT 17.400 10.800 17.800 13.100 ;
        RECT 18.500 10.800 18.900 13.100 ;
        RECT 20.600 10.800 21.000 12.100 ;
        RECT 21.400 10.800 21.800 12.100 ;
        RECT 23.000 10.800 23.400 12.100 ;
        RECT 24.600 10.800 25.000 13.100 ;
        RECT 27.300 10.800 27.800 12.100 ;
        RECT 29.000 10.800 29.400 12.100 ;
        RECT 31.800 10.800 32.200 13.000 ;
        RECT 33.400 10.800 33.800 13.100 ;
        RECT 35.000 10.800 35.400 13.100 ;
        RECT 36.600 10.800 37.000 13.100 ;
        RECT 38.200 10.800 38.600 13.100 ;
        RECT 39.800 10.800 40.200 13.100 ;
        RECT 40.600 10.800 41.000 13.100 ;
        RECT 42.200 10.800 42.600 13.100 ;
        RECT 43.800 10.800 44.200 13.100 ;
        RECT 45.200 10.800 45.600 13.500 ;
        RECT 47.800 10.800 48.200 13.300 ;
        RECT 51.800 10.800 52.200 13.100 ;
        RECT 53.400 10.800 53.800 13.100 ;
        RECT 55.000 10.800 55.400 13.100 ;
        RECT 56.600 10.800 57.000 13.100 ;
        RECT 58.200 10.800 58.600 13.100 ;
        RECT 59.800 10.800 60.200 13.100 ;
        RECT 60.600 10.800 61.000 13.100 ;
        RECT 64.600 10.800 65.000 12.700 ;
        RECT 66.800 10.800 67.200 13.500 ;
        RECT 69.400 10.800 69.800 13.300 ;
        RECT 71.800 10.800 72.200 13.100 ;
        RECT 74.500 10.800 75.000 12.100 ;
        RECT 76.200 10.800 76.600 12.100 ;
        RECT 79.000 10.800 79.400 13.000 ;
        RECT 80.600 10.800 81.000 13.100 ;
        RECT 84.600 10.800 85.000 12.700 ;
        RECT 86.200 10.800 86.600 13.100 ;
        RECT 87.800 10.800 88.200 13.100 ;
        RECT 89.400 10.800 89.800 13.100 ;
        RECT 90.200 10.800 90.600 13.100 ;
        RECT 91.800 10.800 92.200 13.100 ;
        RECT 93.400 10.800 93.800 13.100 ;
        RECT 95.000 10.800 95.400 13.100 ;
        RECT 96.600 10.800 97.000 13.100 ;
        RECT 99.600 10.800 100.000 13.500 ;
        RECT 102.200 10.800 102.600 13.300 ;
        RECT 104.400 10.800 104.800 13.500 ;
        RECT 107.000 10.800 107.400 13.300 ;
        RECT 108.600 10.800 109.000 13.100 ;
        RECT 112.600 10.800 113.000 12.700 ;
        RECT 115.000 10.800 115.400 13.000 ;
        RECT 117.800 10.800 118.200 12.100 ;
        RECT 119.400 10.800 119.900 12.100 ;
        RECT 122.200 10.800 122.600 13.100 ;
        RECT 124.600 10.800 125.000 13.300 ;
        RECT 127.200 10.800 127.600 13.500 ;
        RECT 129.400 10.800 129.800 13.000 ;
        RECT 132.200 10.800 132.600 12.100 ;
        RECT 133.800 10.800 134.300 12.100 ;
        RECT 136.600 10.800 137.000 13.100 ;
        RECT 138.200 10.800 138.600 13.100 ;
        RECT 142.200 10.800 142.600 12.700 ;
        RECT 145.400 10.800 145.800 13.100 ;
        RECT 147.800 10.800 148.200 13.100 ;
        RECT 150.800 10.800 151.200 13.500 ;
        RECT 153.400 10.800 153.800 13.300 ;
        RECT 155.000 10.800 155.400 13.100 ;
        RECT 159.000 10.800 159.400 12.700 ;
        RECT 161.400 10.800 161.800 13.100 ;
        RECT 164.100 10.800 164.600 12.100 ;
        RECT 165.800 10.800 166.200 12.100 ;
        RECT 168.600 10.800 169.000 13.000 ;
        RECT 171.800 10.800 172.200 13.100 ;
        RECT 174.200 10.800 174.600 12.700 ;
        RECT 176.600 10.800 177.000 13.000 ;
        RECT 179.400 10.800 179.800 12.100 ;
        RECT 181.000 10.800 181.500 12.100 ;
        RECT 183.800 10.800 184.200 13.100 ;
        RECT 186.200 10.800 186.600 12.700 ;
        RECT 190.200 10.800 190.600 13.100 ;
        RECT 191.800 10.800 192.200 13.100 ;
        RECT 194.500 10.800 195.000 12.100 ;
        RECT 196.200 10.800 196.600 12.100 ;
        RECT 199.000 10.800 199.400 13.000 ;
        RECT 202.800 10.800 203.200 13.500 ;
        RECT 205.400 10.800 205.800 13.300 ;
        RECT 207.000 10.800 207.400 13.100 ;
        RECT 208.600 10.800 209.000 13.100 ;
        RECT 211.000 10.800 211.400 13.300 ;
        RECT 213.600 10.800 214.000 13.500 ;
        RECT 215.800 10.800 216.200 12.700 ;
        RECT 219.800 10.800 220.200 13.100 ;
        RECT 221.400 10.800 221.800 12.700 ;
        RECT 225.400 10.800 225.800 13.100 ;
        RECT 227.000 10.800 227.400 13.000 ;
        RECT 229.800 10.800 230.200 12.100 ;
        RECT 231.400 10.800 231.900 12.100 ;
        RECT 234.200 10.800 234.600 13.100 ;
        RECT 235.800 10.800 236.200 13.100 ;
        RECT 237.400 10.800 237.800 13.100 ;
        RECT 239.000 10.800 239.400 13.100 ;
        RECT 240.600 10.800 241.000 13.100 ;
        RECT 242.200 10.800 242.600 13.100 ;
        RECT 243.000 10.800 243.400 13.100 ;
        RECT 244.600 10.800 245.000 13.100 ;
        RECT 246.200 10.800 246.600 13.100 ;
        RECT 247.800 10.800 248.200 13.100 ;
        RECT 249.400 10.800 249.800 13.100 ;
        RECT 251.800 10.800 252.200 13.100 ;
        RECT 0.200 10.200 252.600 10.800 ;
        RECT 0.600 7.900 1.000 10.200 ;
        RECT 2.200 7.900 2.600 10.200 ;
        RECT 3.800 7.900 4.200 10.200 ;
        RECT 5.400 7.900 5.800 10.200 ;
        RECT 7.000 7.900 7.400 10.200 ;
        RECT 7.800 7.900 8.200 10.200 ;
        RECT 9.400 7.900 9.800 10.200 ;
        RECT 11.000 7.900 11.400 10.200 ;
        RECT 12.600 7.900 13.000 10.200 ;
        RECT 14.200 7.900 14.600 10.200 ;
        RECT 15.800 8.300 16.200 10.200 ;
        RECT 19.000 7.900 19.400 10.200 ;
        RECT 21.700 8.900 22.200 10.200 ;
        RECT 23.400 8.900 23.800 10.200 ;
        RECT 26.200 8.000 26.600 10.200 ;
        RECT 27.800 8.900 28.200 10.200 ;
        RECT 29.400 8.900 29.800 10.200 ;
        RECT 30.200 8.900 30.600 10.200 ;
        RECT 32.300 7.900 32.700 10.200 ;
        RECT 34.200 7.900 34.600 10.200 ;
        RECT 36.900 8.900 37.400 10.200 ;
        RECT 38.600 8.900 39.000 10.200 ;
        RECT 41.400 8.000 41.800 10.200 ;
        RECT 43.800 8.300 44.200 10.200 ;
        RECT 47.800 7.900 48.200 10.200 ;
        RECT 51.000 8.000 51.400 10.200 ;
        RECT 53.800 8.900 54.200 10.200 ;
        RECT 55.400 8.900 55.900 10.200 ;
        RECT 58.200 7.900 58.600 10.200 ;
        RECT 60.600 8.000 61.000 10.200 ;
        RECT 63.400 8.900 63.800 10.200 ;
        RECT 65.000 8.900 65.500 10.200 ;
        RECT 67.800 7.900 68.200 10.200 ;
        RECT 70.200 7.900 70.600 10.200 ;
        RECT 71.800 7.900 72.200 10.200 ;
        RECT 73.400 7.900 73.800 10.200 ;
        RECT 76.100 8.900 76.600 10.200 ;
        RECT 77.800 8.900 78.200 10.200 ;
        RECT 80.600 8.000 81.000 10.200 ;
        RECT 82.200 7.900 82.600 10.200 ;
        RECT 86.200 8.300 86.600 10.200 ;
        RECT 88.600 7.900 89.000 10.200 ;
        RECT 90.200 7.900 90.600 10.200 ;
        RECT 91.800 8.000 92.200 10.200 ;
        RECT 94.600 8.900 95.000 10.200 ;
        RECT 96.200 8.900 96.700 10.200 ;
        RECT 99.000 7.900 99.400 10.200 ;
        RECT 102.200 7.900 102.600 10.200 ;
        RECT 106.200 8.300 106.600 10.200 ;
        RECT 107.800 7.900 108.200 10.200 ;
        RECT 109.400 7.900 109.800 10.200 ;
        RECT 111.000 7.900 111.400 10.200 ;
        RECT 112.600 7.900 113.000 10.200 ;
        RECT 114.200 7.900 114.600 10.200 ;
        RECT 115.800 7.900 116.200 10.200 ;
        RECT 118.500 8.900 119.000 10.200 ;
        RECT 120.200 8.900 120.600 10.200 ;
        RECT 123.000 8.000 123.400 10.200 ;
        RECT 124.600 7.900 125.000 10.200 ;
        RECT 128.600 8.300 129.000 10.200 ;
        RECT 131.000 7.900 131.400 10.200 ;
        RECT 133.700 8.900 134.200 10.200 ;
        RECT 135.400 8.900 135.800 10.200 ;
        RECT 138.200 8.000 138.600 10.200 ;
        RECT 141.400 8.300 141.800 10.200 ;
        RECT 143.800 8.300 144.200 10.200 ;
        RECT 148.600 8.000 149.000 10.200 ;
        RECT 151.400 8.900 151.800 10.200 ;
        RECT 153.000 8.900 153.500 10.200 ;
        RECT 155.800 7.900 156.200 10.200 ;
        RECT 157.400 7.900 157.800 10.200 ;
        RECT 159.000 7.900 159.400 10.200 ;
        RECT 160.600 7.900 161.000 10.200 ;
        RECT 162.200 7.900 162.600 10.200 ;
        RECT 163.800 7.900 164.200 10.200 ;
        RECT 165.400 8.300 165.800 10.200 ;
        RECT 167.800 7.900 168.200 10.200 ;
        RECT 171.000 8.000 171.400 10.200 ;
        RECT 173.800 8.900 174.200 10.200 ;
        RECT 175.400 8.900 175.900 10.200 ;
        RECT 178.200 7.900 178.600 10.200 ;
        RECT 181.400 7.900 181.800 10.200 ;
        RECT 183.800 8.300 184.200 10.200 ;
        RECT 186.200 7.900 186.600 10.200 ;
        RECT 188.900 8.900 189.400 10.200 ;
        RECT 190.600 8.900 191.000 10.200 ;
        RECT 193.400 8.000 193.800 10.200 ;
        RECT 195.800 8.300 196.200 10.200 ;
        RECT 199.800 7.900 200.200 10.200 ;
        RECT 203.000 7.900 203.400 10.200 ;
        RECT 205.700 8.900 206.200 10.200 ;
        RECT 207.400 8.900 207.800 10.200 ;
        RECT 210.200 8.000 210.600 10.200 ;
        RECT 212.600 7.900 213.000 10.200 ;
        RECT 215.300 8.900 215.800 10.200 ;
        RECT 217.000 8.900 217.400 10.200 ;
        RECT 219.800 8.000 220.200 10.200 ;
        RECT 222.200 8.300 222.600 10.200 ;
        RECT 226.200 7.900 226.600 10.200 ;
        RECT 227.800 8.000 228.200 10.200 ;
        RECT 230.600 8.900 231.000 10.200 ;
        RECT 232.200 8.900 232.700 10.200 ;
        RECT 235.000 7.900 235.400 10.200 ;
        RECT 236.600 7.900 237.000 10.200 ;
        RECT 238.200 7.900 238.600 10.200 ;
        RECT 239.800 7.900 240.200 10.200 ;
        RECT 241.400 7.900 241.800 10.200 ;
        RECT 243.000 7.900 243.400 10.200 ;
        RECT 243.800 7.900 244.200 10.200 ;
        RECT 245.400 7.900 245.800 10.200 ;
        RECT 247.000 7.900 247.400 10.200 ;
        RECT 247.800 7.900 248.200 10.200 ;
        RECT 249.400 7.900 249.800 10.200 ;
        RECT 251.000 7.900 251.400 10.200 ;
      LAYER via1 ;
        RECT 98.600 230.300 99.000 230.700 ;
        RECT 99.300 230.300 99.700 230.700 ;
        RECT 201.800 230.300 202.200 230.700 ;
        RECT 202.500 230.300 202.900 230.700 ;
        RECT 98.600 210.300 99.000 210.700 ;
        RECT 99.300 210.300 99.700 210.700 ;
        RECT 201.800 210.300 202.200 210.700 ;
        RECT 202.500 210.300 202.900 210.700 ;
        RECT 98.600 190.300 99.000 190.700 ;
        RECT 99.300 190.300 99.700 190.700 ;
        RECT 201.800 190.300 202.200 190.700 ;
        RECT 202.500 190.300 202.900 190.700 ;
        RECT 98.600 170.300 99.000 170.700 ;
        RECT 99.300 170.300 99.700 170.700 ;
        RECT 201.800 170.300 202.200 170.700 ;
        RECT 202.500 170.300 202.900 170.700 ;
        RECT 98.600 150.300 99.000 150.700 ;
        RECT 99.300 150.300 99.700 150.700 ;
        RECT 201.800 150.300 202.200 150.700 ;
        RECT 202.500 150.300 202.900 150.700 ;
        RECT 98.600 130.300 99.000 130.700 ;
        RECT 99.300 130.300 99.700 130.700 ;
        RECT 201.800 130.300 202.200 130.700 ;
        RECT 202.500 130.300 202.900 130.700 ;
        RECT 98.600 110.300 99.000 110.700 ;
        RECT 99.300 110.300 99.700 110.700 ;
        RECT 201.800 110.300 202.200 110.700 ;
        RECT 202.500 110.300 202.900 110.700 ;
        RECT 98.600 90.300 99.000 90.700 ;
        RECT 99.300 90.300 99.700 90.700 ;
        RECT 201.800 90.300 202.200 90.700 ;
        RECT 202.500 90.300 202.900 90.700 ;
        RECT 98.600 70.300 99.000 70.700 ;
        RECT 99.300 70.300 99.700 70.700 ;
        RECT 201.800 70.300 202.200 70.700 ;
        RECT 202.500 70.300 202.900 70.700 ;
        RECT 98.600 50.300 99.000 50.700 ;
        RECT 99.300 50.300 99.700 50.700 ;
        RECT 201.800 50.300 202.200 50.700 ;
        RECT 202.500 50.300 202.900 50.700 ;
        RECT 98.600 30.300 99.000 30.700 ;
        RECT 99.300 30.300 99.700 30.700 ;
        RECT 201.800 30.300 202.200 30.700 ;
        RECT 202.500 30.300 202.900 30.700 ;
        RECT 98.600 10.300 99.000 10.700 ;
        RECT 99.300 10.300 99.700 10.700 ;
        RECT 201.800 10.300 202.200 10.700 ;
        RECT 202.500 10.300 202.900 10.700 ;
      LAYER metal2 ;
        RECT 98.400 230.300 100.000 230.700 ;
        RECT 201.600 230.300 203.200 230.700 ;
        RECT 98.400 210.300 100.000 210.700 ;
        RECT 201.600 210.300 203.200 210.700 ;
        RECT 98.400 190.300 100.000 190.700 ;
        RECT 201.600 190.300 203.200 190.700 ;
        RECT 98.400 170.300 100.000 170.700 ;
        RECT 201.600 170.300 203.200 170.700 ;
        RECT 98.400 150.300 100.000 150.700 ;
        RECT 201.600 150.300 203.200 150.700 ;
        RECT 98.400 130.300 100.000 130.700 ;
        RECT 201.600 130.300 203.200 130.700 ;
        RECT 98.400 110.300 100.000 110.700 ;
        RECT 201.600 110.300 203.200 110.700 ;
        RECT 98.400 90.300 100.000 90.700 ;
        RECT 201.600 90.300 203.200 90.700 ;
        RECT 98.400 70.300 100.000 70.700 ;
        RECT 201.600 70.300 203.200 70.700 ;
        RECT 98.400 50.300 100.000 50.700 ;
        RECT 201.600 50.300 203.200 50.700 ;
        RECT 98.400 30.300 100.000 30.700 ;
        RECT 201.600 30.300 203.200 30.700 ;
        RECT 98.400 10.300 100.000 10.700 ;
        RECT 201.600 10.300 203.200 10.700 ;
      LAYER via2 ;
        RECT 98.600 230.300 99.000 230.700 ;
        RECT 99.300 230.300 99.700 230.700 ;
        RECT 201.800 230.300 202.200 230.700 ;
        RECT 202.500 230.300 202.900 230.700 ;
        RECT 98.600 210.300 99.000 210.700 ;
        RECT 99.300 210.300 99.700 210.700 ;
        RECT 201.800 210.300 202.200 210.700 ;
        RECT 202.500 210.300 202.900 210.700 ;
        RECT 98.600 190.300 99.000 190.700 ;
        RECT 99.300 190.300 99.700 190.700 ;
        RECT 201.800 190.300 202.200 190.700 ;
        RECT 202.500 190.300 202.900 190.700 ;
        RECT 98.600 170.300 99.000 170.700 ;
        RECT 99.300 170.300 99.700 170.700 ;
        RECT 201.800 170.300 202.200 170.700 ;
        RECT 202.500 170.300 202.900 170.700 ;
        RECT 98.600 150.300 99.000 150.700 ;
        RECT 99.300 150.300 99.700 150.700 ;
        RECT 201.800 150.300 202.200 150.700 ;
        RECT 202.500 150.300 202.900 150.700 ;
        RECT 98.600 130.300 99.000 130.700 ;
        RECT 99.300 130.300 99.700 130.700 ;
        RECT 201.800 130.300 202.200 130.700 ;
        RECT 202.500 130.300 202.900 130.700 ;
        RECT 98.600 110.300 99.000 110.700 ;
        RECT 99.300 110.300 99.700 110.700 ;
        RECT 201.800 110.300 202.200 110.700 ;
        RECT 202.500 110.300 202.900 110.700 ;
        RECT 98.600 90.300 99.000 90.700 ;
        RECT 99.300 90.300 99.700 90.700 ;
        RECT 201.800 90.300 202.200 90.700 ;
        RECT 202.500 90.300 202.900 90.700 ;
        RECT 98.600 70.300 99.000 70.700 ;
        RECT 99.300 70.300 99.700 70.700 ;
        RECT 201.800 70.300 202.200 70.700 ;
        RECT 202.500 70.300 202.900 70.700 ;
        RECT 98.600 50.300 99.000 50.700 ;
        RECT 99.300 50.300 99.700 50.700 ;
        RECT 201.800 50.300 202.200 50.700 ;
        RECT 202.500 50.300 202.900 50.700 ;
        RECT 98.600 30.300 99.000 30.700 ;
        RECT 99.300 30.300 99.700 30.700 ;
        RECT 201.800 30.300 202.200 30.700 ;
        RECT 202.500 30.300 202.900 30.700 ;
        RECT 98.600 10.300 99.000 10.700 ;
        RECT 99.300 10.300 99.700 10.700 ;
        RECT 201.800 10.300 202.200 10.700 ;
        RECT 202.500 10.300 202.900 10.700 ;
      LAYER metal3 ;
        RECT 98.400 230.300 100.000 230.700 ;
        RECT 201.600 230.300 203.200 230.700 ;
        RECT 98.400 210.300 100.000 210.700 ;
        RECT 201.600 210.300 203.200 210.700 ;
        RECT 98.400 190.300 100.000 190.700 ;
        RECT 201.600 190.300 203.200 190.700 ;
        RECT 98.400 170.300 100.000 170.700 ;
        RECT 201.600 170.300 203.200 170.700 ;
        RECT 98.400 150.300 100.000 150.700 ;
        RECT 201.600 150.300 203.200 150.700 ;
        RECT 98.400 130.300 100.000 130.700 ;
        RECT 201.600 130.300 203.200 130.700 ;
        RECT 98.400 110.300 100.000 110.700 ;
        RECT 201.600 110.300 203.200 110.700 ;
        RECT 98.400 90.300 100.000 90.700 ;
        RECT 201.600 90.300 203.200 90.700 ;
        RECT 98.400 70.300 100.000 70.700 ;
        RECT 201.600 70.300 203.200 70.700 ;
        RECT 98.400 50.300 100.000 50.700 ;
        RECT 201.600 50.300 203.200 50.700 ;
        RECT 98.400 30.300 100.000 30.700 ;
        RECT 201.600 30.300 203.200 30.700 ;
        RECT 98.400 10.300 100.000 10.700 ;
        RECT 201.600 10.300 203.200 10.700 ;
      LAYER via3 ;
        RECT 98.600 230.300 99.000 230.700 ;
        RECT 99.400 230.300 99.800 230.700 ;
        RECT 201.800 230.300 202.200 230.700 ;
        RECT 202.600 230.300 203.000 230.700 ;
        RECT 98.600 210.300 99.000 210.700 ;
        RECT 99.400 210.300 99.800 210.700 ;
        RECT 201.800 210.300 202.200 210.700 ;
        RECT 202.600 210.300 203.000 210.700 ;
        RECT 98.600 190.300 99.000 190.700 ;
        RECT 99.400 190.300 99.800 190.700 ;
        RECT 201.800 190.300 202.200 190.700 ;
        RECT 202.600 190.300 203.000 190.700 ;
        RECT 98.600 170.300 99.000 170.700 ;
        RECT 99.400 170.300 99.800 170.700 ;
        RECT 201.800 170.300 202.200 170.700 ;
        RECT 202.600 170.300 203.000 170.700 ;
        RECT 98.600 150.300 99.000 150.700 ;
        RECT 99.400 150.300 99.800 150.700 ;
        RECT 201.800 150.300 202.200 150.700 ;
        RECT 202.600 150.300 203.000 150.700 ;
        RECT 98.600 130.300 99.000 130.700 ;
        RECT 99.400 130.300 99.800 130.700 ;
        RECT 201.800 130.300 202.200 130.700 ;
        RECT 202.600 130.300 203.000 130.700 ;
        RECT 98.600 110.300 99.000 110.700 ;
        RECT 99.400 110.300 99.800 110.700 ;
        RECT 201.800 110.300 202.200 110.700 ;
        RECT 202.600 110.300 203.000 110.700 ;
        RECT 98.600 90.300 99.000 90.700 ;
        RECT 99.400 90.300 99.800 90.700 ;
        RECT 201.800 90.300 202.200 90.700 ;
        RECT 202.600 90.300 203.000 90.700 ;
        RECT 98.600 70.300 99.000 70.700 ;
        RECT 99.400 70.300 99.800 70.700 ;
        RECT 201.800 70.300 202.200 70.700 ;
        RECT 202.600 70.300 203.000 70.700 ;
        RECT 98.600 50.300 99.000 50.700 ;
        RECT 99.400 50.300 99.800 50.700 ;
        RECT 201.800 50.300 202.200 50.700 ;
        RECT 202.600 50.300 203.000 50.700 ;
        RECT 98.600 30.300 99.000 30.700 ;
        RECT 99.400 30.300 99.800 30.700 ;
        RECT 201.800 30.300 202.200 30.700 ;
        RECT 202.600 30.300 203.000 30.700 ;
        RECT 98.600 10.300 99.000 10.700 ;
        RECT 99.400 10.300 99.800 10.700 ;
        RECT 201.800 10.300 202.200 10.700 ;
        RECT 202.600 10.300 203.000 10.700 ;
      LAYER metal4 ;
        RECT 98.400 230.300 100.000 230.700 ;
        RECT 201.600 230.300 203.200 230.700 ;
        RECT 98.400 210.300 100.000 210.700 ;
        RECT 201.600 210.300 203.200 210.700 ;
        RECT 98.400 190.300 100.000 190.700 ;
        RECT 201.600 190.300 203.200 190.700 ;
        RECT 98.400 170.300 100.000 170.700 ;
        RECT 201.600 170.300 203.200 170.700 ;
        RECT 98.400 150.300 100.000 150.700 ;
        RECT 201.600 150.300 203.200 150.700 ;
        RECT 98.400 130.300 100.000 130.700 ;
        RECT 201.600 130.300 203.200 130.700 ;
        RECT 98.400 110.300 100.000 110.700 ;
        RECT 201.600 110.300 203.200 110.700 ;
        RECT 98.400 90.300 100.000 90.700 ;
        RECT 201.600 90.300 203.200 90.700 ;
        RECT 98.400 70.300 100.000 70.700 ;
        RECT 201.600 70.300 203.200 70.700 ;
        RECT 98.400 50.300 100.000 50.700 ;
        RECT 201.600 50.300 203.200 50.700 ;
        RECT 98.400 30.300 100.000 30.700 ;
        RECT 201.600 30.300 203.200 30.700 ;
        RECT 98.400 10.300 100.000 10.700 ;
        RECT 201.600 10.300 203.200 10.700 ;
      LAYER via4 ;
        RECT 98.600 230.300 99.000 230.700 ;
        RECT 99.300 230.300 99.700 230.700 ;
        RECT 201.800 230.300 202.200 230.700 ;
        RECT 202.500 230.300 202.900 230.700 ;
        RECT 98.600 210.300 99.000 210.700 ;
        RECT 99.300 210.300 99.700 210.700 ;
        RECT 201.800 210.300 202.200 210.700 ;
        RECT 202.500 210.300 202.900 210.700 ;
        RECT 98.600 190.300 99.000 190.700 ;
        RECT 99.300 190.300 99.700 190.700 ;
        RECT 201.800 190.300 202.200 190.700 ;
        RECT 202.500 190.300 202.900 190.700 ;
        RECT 98.600 170.300 99.000 170.700 ;
        RECT 99.300 170.300 99.700 170.700 ;
        RECT 201.800 170.300 202.200 170.700 ;
        RECT 202.500 170.300 202.900 170.700 ;
        RECT 98.600 150.300 99.000 150.700 ;
        RECT 99.300 150.300 99.700 150.700 ;
        RECT 201.800 150.300 202.200 150.700 ;
        RECT 202.500 150.300 202.900 150.700 ;
        RECT 98.600 130.300 99.000 130.700 ;
        RECT 99.300 130.300 99.700 130.700 ;
        RECT 201.800 130.300 202.200 130.700 ;
        RECT 202.500 130.300 202.900 130.700 ;
        RECT 98.600 110.300 99.000 110.700 ;
        RECT 99.300 110.300 99.700 110.700 ;
        RECT 201.800 110.300 202.200 110.700 ;
        RECT 202.500 110.300 202.900 110.700 ;
        RECT 98.600 90.300 99.000 90.700 ;
        RECT 99.300 90.300 99.700 90.700 ;
        RECT 201.800 90.300 202.200 90.700 ;
        RECT 202.500 90.300 202.900 90.700 ;
        RECT 98.600 70.300 99.000 70.700 ;
        RECT 99.300 70.300 99.700 70.700 ;
        RECT 201.800 70.300 202.200 70.700 ;
        RECT 202.500 70.300 202.900 70.700 ;
        RECT 98.600 50.300 99.000 50.700 ;
        RECT 99.300 50.300 99.700 50.700 ;
        RECT 201.800 50.300 202.200 50.700 ;
        RECT 202.500 50.300 202.900 50.700 ;
        RECT 98.600 30.300 99.000 30.700 ;
        RECT 99.300 30.300 99.700 30.700 ;
        RECT 201.800 30.300 202.200 30.700 ;
        RECT 202.500 30.300 202.900 30.700 ;
        RECT 98.600 10.300 99.000 10.700 ;
        RECT 99.300 10.300 99.700 10.700 ;
        RECT 201.800 10.300 202.200 10.700 ;
        RECT 202.500 10.300 202.900 10.700 ;
      LAYER metal5 ;
        RECT 98.400 230.200 100.000 230.700 ;
        RECT 201.600 230.200 203.200 230.700 ;
        RECT 98.400 210.200 100.000 210.700 ;
        RECT 201.600 210.200 203.200 210.700 ;
        RECT 98.400 190.200 100.000 190.700 ;
        RECT 201.600 190.200 203.200 190.700 ;
        RECT 98.400 170.200 100.000 170.700 ;
        RECT 201.600 170.200 203.200 170.700 ;
        RECT 98.400 150.200 100.000 150.700 ;
        RECT 201.600 150.200 203.200 150.700 ;
        RECT 98.400 130.200 100.000 130.700 ;
        RECT 201.600 130.200 203.200 130.700 ;
        RECT 98.400 110.200 100.000 110.700 ;
        RECT 201.600 110.200 203.200 110.700 ;
        RECT 98.400 90.200 100.000 90.700 ;
        RECT 201.600 90.200 203.200 90.700 ;
        RECT 98.400 70.200 100.000 70.700 ;
        RECT 201.600 70.200 203.200 70.700 ;
        RECT 98.400 50.200 100.000 50.700 ;
        RECT 201.600 50.200 203.200 50.700 ;
        RECT 98.400 30.200 100.000 30.700 ;
        RECT 201.600 30.200 203.200 30.700 ;
        RECT 98.400 10.200 100.000 10.700 ;
        RECT 201.600 10.200 203.200 10.700 ;
      LAYER via5 ;
        RECT 99.400 230.200 99.900 230.700 ;
        RECT 202.600 230.200 203.100 230.700 ;
        RECT 99.400 210.200 99.900 210.700 ;
        RECT 202.600 210.200 203.100 210.700 ;
        RECT 99.400 190.200 99.900 190.700 ;
        RECT 202.600 190.200 203.100 190.700 ;
        RECT 99.400 170.200 99.900 170.700 ;
        RECT 202.600 170.200 203.100 170.700 ;
        RECT 99.400 150.200 99.900 150.700 ;
        RECT 202.600 150.200 203.100 150.700 ;
        RECT 99.400 130.200 99.900 130.700 ;
        RECT 202.600 130.200 203.100 130.700 ;
        RECT 99.400 110.200 99.900 110.700 ;
        RECT 202.600 110.200 203.100 110.700 ;
        RECT 99.400 90.200 99.900 90.700 ;
        RECT 202.600 90.200 203.100 90.700 ;
        RECT 99.400 70.200 99.900 70.700 ;
        RECT 202.600 70.200 203.100 70.700 ;
        RECT 99.400 50.200 99.900 50.700 ;
        RECT 202.600 50.200 203.100 50.700 ;
        RECT 99.400 30.200 99.900 30.700 ;
        RECT 202.600 30.200 203.100 30.700 ;
        RECT 99.400 10.200 99.900 10.700 ;
        RECT 202.600 10.200 203.100 10.700 ;
      LAYER metal6 ;
        RECT 98.400 -3.000 100.000 243.000 ;
        RECT 201.600 -3.000 203.200 243.000 ;
    END
  END gnd
  PIN enable
    PORT
      LAYER metal1 ;
        RECT 139.000 44.400 139.400 45.200 ;
        RECT 142.200 33.400 142.600 34.200 ;
      LAYER via1 ;
        RECT 139.000 44.800 139.400 45.200 ;
        RECT 142.200 33.800 142.600 34.200 ;
      LAYER metal2 ;
        RECT 139.000 44.800 139.400 45.200 ;
        RECT 142.200 44.800 142.600 45.200 ;
        RECT 139.000 44.200 139.300 44.800 ;
        RECT 139.000 43.800 139.400 44.200 ;
        RECT 142.200 34.200 142.500 44.800 ;
        RECT 142.200 33.800 142.600 34.200 ;
        RECT 142.200 33.100 142.500 33.800 ;
        RECT 143.000 33.100 143.400 33.200 ;
        RECT 142.200 32.800 143.400 33.100 ;
        RECT 142.200 0.800 142.600 1.200 ;
        RECT 142.200 -1.800 142.500 0.800 ;
        RECT 142.200 -2.200 142.600 -1.800 ;
      LAYER via2 ;
        RECT 143.000 32.800 143.400 33.200 ;
      LAYER metal3 ;
        RECT 142.200 45.100 142.600 45.200 ;
        RECT 139.000 44.800 142.600 45.100 ;
        RECT 139.000 44.200 139.300 44.800 ;
        RECT 139.000 43.800 139.400 44.200 ;
        RECT 142.200 33.100 142.600 33.200 ;
        RECT 143.000 33.100 143.400 33.200 ;
        RECT 142.200 32.800 143.400 33.100 ;
        RECT 142.200 1.800 142.600 2.200 ;
        RECT 142.200 1.200 142.500 1.800 ;
        RECT 142.200 0.800 142.600 1.200 ;
      LAYER metal4 ;
        RECT 142.200 32.800 142.600 33.200 ;
        RECT 142.200 2.200 142.500 32.800 ;
        RECT 142.200 1.800 142.600 2.200 ;
    END
  END enable
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 192.600 214.100 193.500 214.500 ;
        RECT 192.600 213.800 193.000 214.100 ;
        RECT 25.700 194.100 26.600 194.500 ;
        RECT 180.900 194.100 181.800 194.500 ;
        RECT 26.200 193.800 26.600 194.100 ;
        RECT 181.400 193.800 181.800 194.100 ;
        RECT 247.000 186.900 247.400 187.200 ;
        RECT 246.500 186.500 247.400 186.900 ;
        RECT 224.600 154.100 225.500 154.500 ;
        RECT 224.600 153.800 225.000 154.100 ;
        RECT 191.000 146.900 191.400 147.200 ;
        RECT 190.500 146.500 191.400 146.900 ;
        RECT 30.200 134.100 31.100 134.500 ;
        RECT 30.200 133.800 30.600 134.100 ;
        RECT 44.600 106.900 45.000 107.200 ;
        RECT 44.100 106.500 45.000 106.900 ;
        RECT 113.400 106.900 113.800 107.200 ;
        RECT 244.600 106.900 245.000 107.200 ;
        RECT 113.400 106.500 114.300 106.900 ;
        RECT 244.600 106.500 245.500 106.900 ;
        RECT 126.200 94.100 127.100 94.500 ;
        RECT 126.200 93.800 126.600 94.100 ;
        RECT 0.600 86.900 1.000 87.200 ;
        RECT 0.600 86.500 1.500 86.900 ;
        RECT 90.200 14.100 91.100 14.500 ;
        RECT 248.900 14.100 249.800 14.500 ;
        RECT 90.200 13.800 90.600 14.100 ;
        RECT 249.400 13.800 249.800 14.100 ;
        RECT 0.600 6.900 1.000 7.200 ;
        RECT 236.600 6.900 237.000 7.200 ;
        RECT 0.600 6.500 1.500 6.900 ;
        RECT 236.600 6.500 237.500 6.900 ;
      LAYER via1 ;
        RECT 247.000 186.800 247.400 187.200 ;
        RECT 191.000 146.800 191.400 147.200 ;
        RECT 44.600 106.800 45.000 107.200 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 244.600 106.800 245.000 107.200 ;
        RECT 0.600 86.800 1.000 87.200 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 236.600 6.800 237.000 7.200 ;
      LAYER metal2 ;
        RECT 192.600 213.800 193.000 214.200 ;
        RECT 192.600 213.200 192.900 213.800 ;
        RECT 192.600 212.800 193.000 213.200 ;
        RECT 26.200 193.800 26.600 194.200 ;
        RECT 181.400 194.100 181.800 194.200 ;
        RECT 182.200 194.100 182.600 194.200 ;
        RECT 181.400 193.800 182.600 194.100 ;
        RECT 191.000 193.800 191.400 194.200 ;
        RECT 26.200 181.200 26.500 193.800 ;
        RECT 26.200 180.800 26.600 181.200 ;
        RECT 191.000 154.200 191.300 193.800 ;
        RECT 246.200 187.100 246.600 187.200 ;
        RECT 247.000 187.100 247.400 187.200 ;
        RECT 246.200 186.800 247.400 187.100 ;
        RECT 191.000 153.800 191.400 154.200 ;
        RECT 224.600 154.100 225.000 154.200 ;
        RECT 225.400 154.100 225.800 154.200 ;
        RECT 224.600 153.800 225.800 154.100 ;
        RECT 191.000 147.200 191.300 153.800 ;
        RECT 191.000 146.800 191.400 147.200 ;
        RECT 30.200 133.800 30.600 134.200 ;
        RECT 30.200 128.200 30.500 133.800 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 44.600 107.800 45.000 108.200 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 126.200 107.800 126.600 108.200 ;
        RECT 244.600 107.800 245.000 108.200 ;
        RECT 44.600 107.200 44.900 107.800 ;
        RECT 113.400 107.200 113.700 107.800 ;
        RECT 44.600 106.800 45.000 107.200 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 126.200 94.200 126.500 107.800 ;
        RECT 244.600 107.200 244.900 107.800 ;
        RECT 244.600 106.800 245.000 107.200 ;
        RECT 126.200 93.800 126.600 94.200 ;
        RECT 0.600 87.100 1.000 87.200 ;
        RECT 1.400 87.100 1.800 87.200 ;
        RECT 0.600 86.800 1.800 87.100 ;
        RECT 90.200 17.800 90.600 18.200 ;
        RECT 90.200 14.200 90.500 17.800 ;
        RECT 90.200 13.800 90.600 14.200 ;
        RECT 236.600 13.800 237.000 14.200 ;
        RECT 248.600 14.100 249.000 14.200 ;
        RECT 249.400 14.100 249.800 14.200 ;
        RECT 248.600 13.800 249.800 14.100 ;
        RECT 0.600 7.800 1.000 8.200 ;
        RECT 0.600 7.200 0.900 7.800 ;
        RECT 236.600 7.200 236.900 13.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 236.600 6.800 237.000 7.200 ;
      LAYER via2 ;
        RECT 182.200 193.800 182.600 194.200 ;
        RECT 225.400 153.800 225.800 154.200 ;
        RECT 1.400 86.800 1.800 87.200 ;
      LAYER metal3 ;
        RECT 191.800 214.100 192.200 214.200 ;
        RECT 191.800 213.800 192.900 214.100 ;
        RECT 192.600 213.200 192.900 213.800 ;
        RECT 192.600 212.800 193.000 213.200 ;
        RECT 182.200 194.100 182.600 194.200 ;
        RECT 191.000 194.100 191.400 194.200 ;
        RECT 191.800 194.100 192.200 194.200 ;
        RECT 182.200 193.800 192.200 194.100 ;
        RECT 234.200 187.100 234.600 187.200 ;
        RECT 246.200 187.100 246.600 187.200 ;
        RECT 234.200 186.800 246.600 187.100 ;
        RECT 26.200 181.100 26.600 181.200 ;
        RECT 30.200 181.100 30.600 181.200 ;
        RECT 26.200 180.800 30.600 181.100 ;
        RECT 191.000 154.100 191.400 154.200 ;
        RECT 224.600 154.100 225.000 154.200 ;
        RECT 225.400 154.100 225.800 154.200 ;
        RECT 234.200 154.100 234.600 154.200 ;
        RECT 191.000 153.800 234.600 154.100 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 30.200 127.200 30.500 127.800 ;
        RECT 30.200 126.800 30.600 127.200 ;
        RECT 0.600 108.100 1.000 108.200 ;
        RECT 30.200 108.100 30.600 108.200 ;
        RECT 44.600 108.100 45.000 108.200 ;
        RECT 90.200 108.100 90.600 108.200 ;
        RECT 113.400 108.100 113.800 108.200 ;
        RECT 126.200 108.100 126.600 108.200 ;
        RECT 224.600 108.100 225.000 108.200 ;
        RECT 244.600 108.100 245.000 108.200 ;
        RECT 0.600 107.800 245.000 108.100 ;
        RECT -2.600 87.100 -2.200 87.200 ;
        RECT 0.600 87.100 1.000 87.200 ;
        RECT 1.400 87.100 1.800 87.200 ;
        RECT -2.600 86.800 1.800 87.100 ;
        RECT 90.200 18.800 90.600 19.200 ;
        RECT 90.200 18.200 90.500 18.800 ;
        RECT 90.200 17.800 90.600 18.200 ;
        RECT 236.600 14.100 237.000 14.200 ;
        RECT 244.600 14.100 245.000 14.200 ;
        RECT 248.600 14.100 249.000 14.200 ;
        RECT 236.600 13.800 249.000 14.100 ;
        RECT 0.600 7.800 1.000 8.200 ;
        RECT 0.600 7.200 0.900 7.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
      LAYER via3 ;
        RECT 191.800 193.800 192.200 194.200 ;
        RECT 30.200 180.800 30.600 181.200 ;
        RECT 224.600 153.800 225.000 154.200 ;
        RECT 234.200 153.800 234.600 154.200 ;
        RECT 30.200 107.800 30.600 108.200 ;
        RECT 90.200 107.800 90.600 108.200 ;
        RECT 224.600 107.800 225.000 108.200 ;
        RECT 244.600 107.800 245.000 108.200 ;
        RECT 0.600 86.800 1.000 87.200 ;
        RECT 244.600 13.800 245.000 14.200 ;
      LAYER metal4 ;
        RECT 191.800 213.800 192.200 214.200 ;
        RECT 191.800 194.200 192.100 213.800 ;
        RECT 191.800 193.800 192.200 194.200 ;
        RECT 234.200 186.800 234.600 187.200 ;
        RECT 30.200 180.800 30.600 181.200 ;
        RECT 30.200 127.200 30.500 180.800 ;
        RECT 234.200 154.200 234.500 186.800 ;
        RECT 224.600 153.800 225.000 154.200 ;
        RECT 234.200 153.800 234.600 154.200 ;
        RECT 30.200 126.800 30.600 127.200 ;
        RECT 30.200 108.200 30.500 126.800 ;
        RECT 224.600 108.200 224.900 153.800 ;
        RECT 0.600 107.800 1.000 108.200 ;
        RECT 30.200 107.800 30.600 108.200 ;
        RECT 90.200 107.800 90.600 108.200 ;
        RECT 224.600 107.800 225.000 108.200 ;
        RECT 244.600 107.800 245.000 108.200 ;
        RECT 0.600 87.200 0.900 107.800 ;
        RECT 0.600 86.800 1.000 87.200 ;
        RECT 0.600 7.200 0.900 86.800 ;
        RECT 90.200 19.200 90.500 107.800 ;
        RECT 90.200 18.800 90.600 19.200 ;
        RECT 244.600 14.200 244.900 107.800 ;
        RECT 244.600 13.800 245.000 14.200 ;
        RECT 0.600 6.800 1.000 7.200 ;
    END
  END clk
  PIN r_w
    PORT
      LAYER metal1 ;
        RECT 118.200 213.400 118.600 214.200 ;
        RECT 180.600 213.400 181.000 214.200 ;
        RECT 54.200 207.100 54.600 207.600 ;
        RECT 55.000 207.100 55.400 207.200 ;
        RECT 54.200 206.800 55.400 207.100 ;
        RECT 113.400 153.400 113.800 154.200 ;
        RECT 79.000 146.800 79.400 147.600 ;
        RECT 174.200 106.800 174.600 107.600 ;
        RECT 159.000 73.400 159.400 74.200 ;
        RECT 47.000 47.100 47.400 47.600 ;
        RECT 49.400 47.100 49.800 47.600 ;
        RECT 47.000 46.800 49.800 47.100 ;
        RECT 137.400 46.800 137.800 47.600 ;
      LAYER via1 ;
        RECT 118.200 213.800 118.600 214.200 ;
        RECT 180.600 213.800 181.000 214.200 ;
        RECT 55.000 206.800 55.400 207.200 ;
        RECT 113.400 153.800 113.800 154.200 ;
        RECT 159.000 73.800 159.400 74.200 ;
        RECT 49.400 46.800 49.800 47.200 ;
      LAYER metal2 ;
        RECT 180.600 242.800 181.000 243.200 ;
        RECT 180.600 240.200 180.900 242.800 ;
        RECT 180.600 239.800 181.000 240.200 ;
        RECT 118.200 213.800 118.600 214.200 ;
        RECT 180.600 213.800 181.000 214.200 ;
        RECT 118.200 213.200 118.500 213.800 ;
        RECT 180.600 213.200 180.900 213.800 ;
        RECT 118.200 212.800 118.600 213.200 ;
        RECT 180.600 212.800 181.000 213.200 ;
        RECT 55.000 206.800 55.400 207.200 ;
        RECT 55.000 196.200 55.300 206.800 ;
        RECT 118.200 197.200 118.500 212.800 ;
        RECT 118.200 196.800 118.600 197.200 ;
        RECT 55.000 195.800 55.400 196.200 ;
        RECT 113.400 153.800 113.800 154.200 ;
        RECT 113.400 153.200 113.700 153.800 ;
        RECT 79.000 152.800 79.400 153.200 ;
        RECT 113.400 152.800 113.800 153.200 ;
        RECT 79.000 150.200 79.300 152.800 ;
        RECT 79.000 149.800 79.400 150.200 ;
        RECT 79.000 147.200 79.300 149.800 ;
        RECT 79.000 146.800 79.400 147.200 ;
        RECT 174.200 110.800 174.600 111.200 ;
        RECT 174.200 107.200 174.500 110.800 ;
        RECT 174.200 106.800 174.600 107.200 ;
        RECT 174.200 79.200 174.500 106.800 ;
        RECT 159.000 78.800 159.400 79.200 ;
        RECT 174.200 78.800 174.600 79.200 ;
        RECT 159.000 74.200 159.300 78.800 ;
        RECT 159.000 73.800 159.400 74.200 ;
        RECT 159.000 58.200 159.300 73.800 ;
        RECT 159.000 57.800 159.400 58.200 ;
        RECT 49.400 49.800 49.800 50.200 ;
        RECT 49.400 47.200 49.700 49.800 ;
        RECT 49.400 46.800 49.800 47.200 ;
        RECT 137.400 47.100 137.800 47.200 ;
        RECT 138.200 47.100 138.600 47.200 ;
        RECT 137.400 46.800 138.600 47.100 ;
      LAYER via2 ;
        RECT 138.200 46.800 138.600 47.200 ;
      LAYER metal3 ;
        RECT 180.600 239.800 181.000 240.200 ;
        RECT 180.600 239.200 180.900 239.800 ;
        RECT 180.600 238.800 181.000 239.200 ;
        RECT 118.200 213.100 118.600 213.200 ;
        RECT 174.200 213.100 174.600 213.200 ;
        RECT 180.600 213.100 181.000 213.200 ;
        RECT 118.200 212.800 181.000 213.100 ;
        RECT 117.400 197.100 117.800 197.200 ;
        RECT 118.200 197.100 118.600 197.200 ;
        RECT 117.400 196.800 118.600 197.100 ;
        RECT 55.000 196.100 55.400 196.200 ;
        RECT 56.600 196.100 57.000 196.200 ;
        RECT 55.000 195.800 57.000 196.100 ;
        RECT 79.000 153.100 79.400 153.200 ;
        RECT 113.400 153.100 113.800 153.200 ;
        RECT 118.200 153.100 118.600 153.200 ;
        RECT 79.000 152.800 118.600 153.100 ;
        RECT 56.600 150.100 57.000 150.200 ;
        RECT 57.400 150.100 57.800 150.200 ;
        RECT 79.000 150.100 79.400 150.200 ;
        RECT 56.600 149.800 79.400 150.100 ;
        RECT 174.200 111.100 174.600 111.200 ;
        RECT 175.000 111.100 175.400 111.200 ;
        RECT 174.200 110.800 175.400 111.100 ;
        RECT 159.000 79.100 159.400 79.200 ;
        RECT 174.200 79.100 174.600 79.200 ;
        RECT 159.000 78.800 174.600 79.100 ;
        RECT 139.800 58.100 140.200 58.200 ;
        RECT 159.000 58.100 159.400 58.200 ;
        RECT 139.800 57.800 159.400 58.100 ;
        RECT 49.400 50.100 49.800 50.200 ;
        RECT 57.400 50.100 57.800 50.200 ;
        RECT 49.400 49.800 57.800 50.100 ;
        RECT 138.200 47.100 138.600 47.200 ;
        RECT 139.800 47.100 140.200 47.200 ;
        RECT 138.200 46.800 140.200 47.100 ;
      LAYER via3 ;
        RECT 174.200 212.800 174.600 213.200 ;
        RECT 180.600 212.800 181.000 213.200 ;
        RECT 56.600 195.800 57.000 196.200 ;
        RECT 118.200 152.800 118.600 153.200 ;
        RECT 57.400 149.800 57.800 150.200 ;
        RECT 175.000 110.800 175.400 111.200 ;
        RECT 57.400 49.800 57.800 50.200 ;
        RECT 139.800 46.800 140.200 47.200 ;
      LAYER metal4 ;
        RECT 180.600 238.800 181.000 239.200 ;
        RECT 180.600 213.200 180.900 238.800 ;
        RECT 174.200 212.800 174.600 213.200 ;
        RECT 180.600 212.800 181.000 213.200 ;
        RECT 117.400 197.100 117.800 197.200 ;
        RECT 117.400 196.800 118.500 197.100 ;
        RECT 56.600 195.800 57.000 196.200 ;
        RECT 56.600 150.200 56.900 195.800 ;
        RECT 118.200 153.200 118.500 196.800 ;
        RECT 118.200 152.800 118.600 153.200 ;
        RECT 56.600 149.800 57.000 150.200 ;
        RECT 57.400 149.800 57.800 150.200 ;
        RECT 57.400 50.200 57.700 149.800 ;
        RECT 174.200 111.100 174.500 212.800 ;
        RECT 175.000 111.100 175.400 111.200 ;
        RECT 174.200 110.800 175.400 111.100 ;
        RECT 139.800 57.800 140.200 58.200 ;
        RECT 57.400 49.800 57.800 50.200 ;
        RECT 139.800 47.200 140.100 57.800 ;
        RECT 139.800 46.800 140.200 47.200 ;
    END
  END r_w
  PIN datain[0]
    PORT
      LAYER metal1 ;
        RECT 24.600 233.400 25.000 234.200 ;
      LAYER via1 ;
        RECT 24.600 233.800 25.000 234.200 ;
      LAYER metal2 ;
        RECT 26.200 242.800 26.600 243.200 ;
        RECT 26.200 240.200 26.500 242.800 ;
        RECT 24.600 239.800 25.000 240.200 ;
        RECT 26.200 239.800 26.600 240.200 ;
        RECT 24.600 234.200 24.900 239.800 ;
        RECT 24.600 233.800 25.000 234.200 ;
      LAYER metal3 ;
        RECT 24.600 240.100 25.000 240.200 ;
        RECT 26.200 240.100 26.600 240.200 ;
        RECT 24.600 239.800 26.600 240.100 ;
    END
  END datain[0]
  PIN datain[1]
    PORT
      LAYER metal1 ;
        RECT 0.600 133.400 1.000 134.200 ;
      LAYER via1 ;
        RECT 0.600 133.800 1.000 134.200 ;
      LAYER metal2 ;
        RECT 0.600 134.800 1.000 135.200 ;
        RECT 0.600 134.200 0.900 134.800 ;
        RECT 0.600 133.800 1.000 134.200 ;
      LAYER metal3 ;
        RECT -2.600 135.100 -2.200 135.200 ;
        RECT 0.600 135.100 1.000 135.200 ;
        RECT -2.600 134.800 1.000 135.100 ;
    END
  END datain[1]
  PIN datain[2]
    PORT
      LAYER metal1 ;
        RECT 115.800 233.400 116.200 234.200 ;
      LAYER via1 ;
        RECT 115.800 233.800 116.200 234.200 ;
      LAYER metal2 ;
        RECT 114.200 242.800 114.600 243.200 ;
        RECT 114.200 240.200 114.500 242.800 ;
        RECT 114.200 239.800 114.600 240.200 ;
        RECT 115.800 239.800 116.200 240.200 ;
        RECT 115.800 234.200 116.100 239.800 ;
        RECT 115.800 233.800 116.200 234.200 ;
      LAYER metal3 ;
        RECT 114.200 240.100 114.600 240.200 ;
        RECT 115.800 240.100 116.200 240.200 ;
        RECT 114.200 239.800 116.200 240.100 ;
    END
  END datain[2]
  PIN datain[3]
    PORT
      LAYER metal1 ;
        RECT 251.800 7.800 252.200 8.200 ;
        RECT 251.000 7.100 251.400 7.600 ;
        RECT 251.800 7.100 252.100 7.800 ;
        RECT 251.000 6.800 252.100 7.100 ;
      LAYER metal2 ;
        RECT 251.800 7.800 252.200 8.200 ;
        RECT 251.800 7.200 252.100 7.800 ;
        RECT 251.800 6.800 252.200 7.200 ;
      LAYER metal3 ;
        RECT 251.800 7.100 252.200 7.200 ;
        RECT 255.000 7.100 255.400 7.200 ;
        RECT 251.800 6.800 255.400 7.100 ;
    END
  END datain[3]
  PIN datain[4]
    PORT
      LAYER metal1 ;
        RECT 43.800 13.400 44.200 14.200 ;
      LAYER via1 ;
        RECT 43.800 13.800 44.200 14.200 ;
      LAYER metal2 ;
        RECT 43.800 13.800 44.200 14.200 ;
        RECT 43.800 8.200 44.100 13.800 ;
        RECT 42.200 7.800 42.600 8.200 ;
        RECT 43.800 7.800 44.200 8.200 ;
        RECT 42.200 -1.800 42.500 7.800 ;
        RECT 42.200 -2.200 42.600 -1.800 ;
      LAYER metal3 ;
        RECT 42.200 8.100 42.600 8.200 ;
        RECT 43.800 8.100 44.200 8.200 ;
        RECT 42.200 7.800 44.200 8.100 ;
    END
  END datain[4]
  PIN datain[5]
    PORT
      LAYER metal1 ;
        RECT 247.000 7.100 247.400 7.600 ;
        RECT 247.800 7.100 248.200 7.200 ;
        RECT 247.000 6.800 248.200 7.100 ;
      LAYER via1 ;
        RECT 247.800 6.800 248.200 7.200 ;
      LAYER metal2 ;
        RECT 247.800 6.800 248.200 7.200 ;
        RECT 247.800 5.200 248.100 6.800 ;
        RECT 247.800 4.800 248.200 5.200 ;
      LAYER metal3 ;
        RECT 247.800 5.100 248.200 5.200 ;
        RECT 255.000 5.100 255.400 5.200 ;
        RECT 247.800 4.800 255.400 5.100 ;
    END
  END datain[5]
  PIN datain[6]
    PORT
      LAYER metal1 ;
        RECT 89.400 13.400 89.800 14.200 ;
      LAYER via1 ;
        RECT 89.400 13.800 89.800 14.200 ;
      LAYER metal2 ;
        RECT 89.400 13.800 89.800 14.200 ;
        RECT 89.400 10.100 89.700 13.800 ;
        RECT 88.600 9.800 89.700 10.100 ;
        RECT 87.800 -1.900 88.200 -1.800 ;
        RECT 88.600 -1.900 88.900 9.800 ;
        RECT 87.800 -2.200 88.900 -1.900 ;
    END
  END datain[6]
  PIN datain[7]
    PORT
      LAYER metal1 ;
        RECT 245.400 233.400 245.800 234.200 ;
      LAYER via1 ;
        RECT 245.400 233.800 245.800 234.200 ;
      LAYER metal2 ;
        RECT 245.400 235.800 245.800 236.200 ;
        RECT 245.400 234.200 245.700 235.800 ;
        RECT 245.400 233.800 245.800 234.200 ;
      LAYER metal3 ;
        RECT 245.400 236.100 245.800 236.200 ;
        RECT 245.400 235.800 255.300 236.100 ;
        RECT 255.000 235.200 255.300 235.800 ;
        RECT 255.000 234.800 255.400 235.200 ;
    END
  END datain[7]
  PIN address[0]
    PORT
      LAYER metal1 ;
        RECT 203.800 55.100 204.200 55.200 ;
        RECT 204.600 55.100 205.100 55.200 ;
        RECT 203.800 54.800 205.100 55.100 ;
        RECT 204.700 54.400 205.100 54.800 ;
        RECT 163.700 46.200 164.100 46.600 ;
        RECT 166.900 46.200 167.300 46.600 ;
        RECT 170.100 46.200 170.500 46.600 ;
        RECT 171.100 46.200 171.500 46.600 ;
        RECT 174.300 46.200 174.700 46.600 ;
        RECT 163.700 45.800 164.200 46.200 ;
        RECT 166.900 46.100 167.400 46.200 ;
        RECT 167.800 46.100 168.200 46.200 ;
        RECT 166.900 45.800 168.200 46.100 ;
        RECT 170.100 46.100 170.600 46.200 ;
        RECT 171.000 46.100 171.500 46.200 ;
        RECT 170.100 45.800 171.500 46.100 ;
        RECT 174.200 45.800 174.700 46.200 ;
        RECT 179.700 46.200 180.100 46.600 ;
        RECT 179.700 45.800 180.200 46.200 ;
        RECT 162.900 35.100 163.400 35.200 ;
        RECT 163.800 35.100 164.300 35.200 ;
        RECT 162.900 34.800 164.300 35.100 ;
        RECT 174.200 34.800 174.700 35.200 ;
        RECT 162.900 34.400 163.300 34.800 ;
        RECT 163.900 34.400 164.300 34.800 ;
        RECT 174.300 34.400 174.700 34.800 ;
        RECT 203.100 26.200 203.500 26.600 ;
        RECT 203.000 25.800 203.500 26.200 ;
      LAYER via1 ;
        RECT 163.800 45.800 164.200 46.200 ;
        RECT 167.800 45.800 168.200 46.200 ;
        RECT 170.200 45.800 170.600 46.200 ;
        RECT 179.800 45.800 180.200 46.200 ;
        RECT 163.800 34.800 164.200 35.200 ;
      LAYER metal2 ;
        RECT 203.800 54.800 204.200 55.200 ;
        RECT 203.800 48.200 204.100 54.800 ;
        RECT 179.800 47.800 180.200 48.200 ;
        RECT 203.800 47.800 204.200 48.200 ;
        RECT 179.800 46.200 180.100 47.800 ;
        RECT 163.800 46.100 164.200 46.200 ;
        RECT 164.600 46.100 165.000 46.200 ;
        RECT 163.800 45.800 165.000 46.100 ;
        RECT 167.800 46.100 168.200 46.200 ;
        RECT 168.600 46.100 169.000 46.200 ;
        RECT 167.800 45.800 169.000 46.100 ;
        RECT 170.200 45.800 170.600 46.200 ;
        RECT 174.200 45.800 174.600 46.200 ;
        RECT 179.000 46.100 179.400 46.200 ;
        RECT 179.800 46.100 180.200 46.200 ;
        RECT 179.000 45.800 180.200 46.100 ;
        RECT 163.800 35.200 164.100 45.800 ;
        RECT 170.200 45.200 170.500 45.800 ;
        RECT 170.200 44.800 170.600 45.200 ;
        RECT 174.200 35.200 174.500 45.800 ;
        RECT 163.800 34.800 164.200 35.200 ;
        RECT 174.200 34.800 174.600 35.200 ;
        RECT 203.000 26.100 203.400 26.200 ;
        RECT 203.800 26.100 204.100 47.800 ;
        RECT 203.000 25.800 204.100 26.100 ;
        RECT 203.800 11.200 204.100 25.800 ;
        RECT 203.800 10.800 204.200 11.200 ;
        RECT 203.800 0.800 204.200 1.200 ;
        RECT 203.800 -1.800 204.100 0.800 ;
        RECT 203.800 -2.200 204.200 -1.800 ;
      LAYER via2 ;
        RECT 164.600 45.800 165.000 46.200 ;
        RECT 168.600 45.800 169.000 46.200 ;
      LAYER metal3 ;
        RECT 179.800 48.100 180.200 48.200 ;
        RECT 203.800 48.100 204.200 48.200 ;
        RECT 179.800 47.800 204.200 48.100 ;
        RECT 164.600 46.100 165.000 46.200 ;
        RECT 168.600 46.100 169.000 46.200 ;
        RECT 174.200 46.100 174.600 46.200 ;
        RECT 179.000 46.100 179.400 46.200 ;
        RECT 164.600 45.800 179.400 46.100 ;
        RECT 170.200 45.200 170.500 45.800 ;
        RECT 170.200 44.800 170.600 45.200 ;
        RECT 203.800 10.800 204.200 11.200 ;
        RECT 203.800 10.200 204.100 10.800 ;
        RECT 203.800 9.800 204.200 10.200 ;
        RECT 203.800 1.800 204.200 2.200 ;
        RECT 203.800 1.200 204.100 1.800 ;
        RECT 203.800 0.800 204.200 1.200 ;
      LAYER metal4 ;
        RECT 203.800 9.800 204.200 10.200 ;
        RECT 203.800 2.200 204.100 9.800 ;
        RECT 203.800 1.800 204.200 2.200 ;
    END
  END address[0]
  PIN address[1]
    PORT
      LAYER metal1 ;
        RECT 138.100 94.800 138.600 95.200 ;
        RECT 141.300 94.800 141.800 95.200 ;
        RECT 144.500 95.100 145.000 95.200 ;
        RECT 145.400 95.100 145.900 95.200 ;
        RECT 144.500 94.800 145.900 95.100 ;
        RECT 138.100 94.400 138.500 94.800 ;
        RECT 141.300 94.400 141.700 94.800 ;
        RECT 144.500 94.400 144.900 94.800 ;
        RECT 145.500 94.400 145.900 94.800 ;
        RECT 150.900 94.800 151.400 95.200 ;
        RECT 150.900 94.400 151.300 94.800 ;
        RECT 143.000 74.800 143.500 75.200 ;
        RECT 143.100 74.400 143.500 74.800 ;
        RECT 165.300 74.800 165.800 75.200 ;
        RECT 165.300 74.400 165.700 74.800 ;
        RECT 165.500 26.200 165.900 26.600 ;
        RECT 165.400 25.800 165.900 26.200 ;
      LAYER via1 ;
        RECT 138.200 94.800 138.600 95.200 ;
        RECT 141.400 94.800 141.800 95.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 151.000 94.800 151.400 95.200 ;
        RECT 165.400 74.800 165.800 75.200 ;
      LAYER metal2 ;
        RECT 138.200 95.100 138.600 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 138.200 94.800 139.400 95.100 ;
        RECT 141.400 95.100 141.800 95.200 ;
        RECT 142.200 95.100 142.600 95.200 ;
        RECT 141.400 94.800 142.600 95.100 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 150.200 95.100 150.600 95.200 ;
        RECT 151.000 95.100 151.400 95.200 ;
        RECT 150.200 94.800 151.400 95.100 ;
        RECT 145.400 76.200 145.700 94.800 ;
        RECT 143.000 75.800 143.400 76.200 ;
        RECT 145.400 75.800 145.800 76.200 ;
        RECT 165.400 75.800 165.800 76.200 ;
        RECT 143.000 75.200 143.300 75.800 ;
        RECT 165.400 75.200 165.700 75.800 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 165.400 73.200 165.700 74.800 ;
        RECT 165.400 72.800 165.800 73.200 ;
        RECT 164.600 26.100 165.000 26.200 ;
        RECT 165.400 26.100 165.800 26.200 ;
        RECT 164.600 25.800 165.800 26.100 ;
        RECT 165.400 0.800 165.800 1.200 ;
        RECT 165.400 -1.800 165.700 0.800 ;
        RECT 165.400 -2.200 165.800 -1.800 ;
      LAYER via2 ;
        RECT 139.000 94.800 139.400 95.200 ;
        RECT 142.200 94.800 142.600 95.200 ;
      LAYER metal3 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 142.200 95.100 142.600 95.200 ;
        RECT 145.400 95.100 145.800 95.200 ;
        RECT 150.200 95.100 150.600 95.200 ;
        RECT 139.000 94.800 150.600 95.100 ;
        RECT 143.000 76.100 143.400 76.200 ;
        RECT 145.400 76.100 145.800 76.200 ;
        RECT 165.400 76.100 165.800 76.200 ;
        RECT 143.000 75.800 165.800 76.100 ;
        RECT 165.400 73.800 165.800 74.200 ;
        RECT 165.400 73.200 165.700 73.800 ;
        RECT 165.400 72.800 165.800 73.200 ;
        RECT 164.600 26.100 165.000 26.200 ;
        RECT 165.400 26.100 165.800 26.200 ;
        RECT 164.600 25.800 165.800 26.100 ;
        RECT 165.400 1.800 165.800 2.200 ;
        RECT 165.400 1.200 165.700 1.800 ;
        RECT 165.400 0.800 165.800 1.200 ;
      LAYER via3 ;
        RECT 165.400 25.800 165.800 26.200 ;
      LAYER metal4 ;
        RECT 165.400 73.800 165.800 74.200 ;
        RECT 165.400 26.200 165.700 73.800 ;
        RECT 165.400 25.800 165.800 26.200 ;
        RECT 165.400 2.200 165.700 25.800 ;
        RECT 165.400 1.800 165.800 2.200 ;
    END
  END address[1]
  PIN address[2]
    PORT
      LAYER metal1 ;
        RECT 41.400 153.400 41.800 154.200 ;
        RECT 37.400 152.400 37.800 153.200 ;
        RECT 52.600 152.400 53.000 153.200 ;
        RECT 50.200 147.800 50.600 148.600 ;
        RECT 55.000 147.800 55.400 148.600 ;
      LAYER via1 ;
        RECT 41.400 153.800 41.800 154.200 ;
        RECT 37.400 152.800 37.800 153.200 ;
        RECT 52.600 152.800 53.000 153.200 ;
      LAYER metal2 ;
        RECT 41.400 153.800 41.800 154.200 ;
        RECT 37.400 152.800 37.800 153.200 ;
        RECT 37.400 150.200 37.700 152.800 ;
        RECT 37.400 149.800 37.800 150.200 ;
        RECT 37.400 149.200 37.700 149.800 ;
        RECT 41.400 149.200 41.700 153.800 ;
        RECT 52.600 152.800 53.000 153.200 ;
        RECT 52.600 149.200 52.900 152.800 ;
        RECT 37.400 148.800 37.800 149.200 ;
        RECT 41.400 148.800 41.800 149.200 ;
        RECT 50.200 148.800 50.600 149.200 ;
        RECT 52.600 148.800 53.000 149.200 ;
        RECT 55.000 148.800 55.400 149.200 ;
        RECT 50.200 148.200 50.500 148.800 ;
        RECT 55.000 148.200 55.300 148.800 ;
        RECT 50.200 147.800 50.600 148.200 ;
        RECT 55.000 147.800 55.400 148.200 ;
      LAYER metal3 ;
        RECT -2.600 155.100 -2.200 155.200 ;
        RECT 0.600 155.100 1.000 155.200 ;
        RECT -2.600 154.800 1.000 155.100 ;
        RECT 0.600 150.100 1.000 150.200 ;
        RECT 37.400 150.100 37.800 150.200 ;
        RECT 0.600 149.800 37.800 150.100 ;
        RECT 37.400 149.100 37.800 149.200 ;
        RECT 41.400 149.100 41.800 149.200 ;
        RECT 50.200 149.100 50.600 149.200 ;
        RECT 52.600 149.100 53.000 149.200 ;
        RECT 55.000 149.100 55.400 149.200 ;
        RECT 37.400 148.800 55.400 149.100 ;
      LAYER via3 ;
        RECT 0.600 154.800 1.000 155.200 ;
      LAYER metal4 ;
        RECT 0.600 154.800 1.000 155.200 ;
        RECT 0.600 150.200 0.900 154.800 ;
        RECT 0.600 149.800 1.000 150.200 ;
    END
  END address[2]
  PIN address[3]
    PORT
      LAYER metal1 ;
        RECT 38.200 147.800 38.600 148.600 ;
        RECT 32.600 146.800 33.000 147.600 ;
        RECT 43.800 146.800 44.200 147.600 ;
      LAYER metal2 ;
        RECT 32.600 147.800 33.000 148.200 ;
        RECT 37.400 148.100 37.800 148.200 ;
        RECT 38.200 148.100 38.600 148.200 ;
        RECT 37.400 147.800 38.600 148.100 ;
        RECT 32.600 147.200 32.900 147.800 ;
        RECT 38.200 147.200 38.500 147.800 ;
        RECT 32.600 146.800 33.000 147.200 ;
        RECT 38.200 146.800 38.600 147.200 ;
        RECT 43.000 147.100 43.400 147.200 ;
        RECT 43.800 147.100 44.200 147.200 ;
        RECT 43.000 146.800 44.200 147.100 ;
      LAYER metal3 ;
        RECT 3.000 148.100 3.400 148.200 ;
        RECT 32.600 148.100 33.000 148.200 ;
        RECT 37.400 148.100 37.800 148.200 ;
        RECT 3.000 147.800 37.800 148.100 ;
        RECT 38.200 147.100 38.600 147.200 ;
        RECT 43.000 147.100 43.400 147.200 ;
        RECT 38.200 146.800 43.400 147.100 ;
        RECT 3.000 146.100 3.400 146.200 ;
        RECT -2.600 145.800 3.400 146.100 ;
        RECT -2.600 145.200 -2.300 145.800 ;
        RECT -2.600 144.800 -2.200 145.200 ;
      LAYER via3 ;
        RECT 3.000 145.800 3.400 146.200 ;
      LAYER metal4 ;
        RECT 3.000 147.800 3.400 148.200 ;
        RECT 3.000 146.200 3.300 147.800 ;
        RECT 3.000 145.800 3.400 146.200 ;
    END
  END address[3]
  PIN address[4]
    PORT
      LAYER metal1 ;
        RECT 31.000 147.800 31.400 148.600 ;
        RECT 46.200 146.800 46.600 147.600 ;
        RECT 45.400 144.400 45.800 145.200 ;
      LAYER via1 ;
        RECT 45.400 144.800 45.800 145.200 ;
      LAYER metal2 ;
        RECT 31.000 147.800 31.400 148.200 ;
        RECT 31.000 145.200 31.300 147.800 ;
        RECT 46.200 146.800 46.600 147.200 ;
        RECT 31.000 144.800 31.400 145.200 ;
        RECT 44.600 145.100 45.000 145.200 ;
        RECT 45.400 145.100 45.800 145.200 ;
        RECT 46.200 145.100 46.500 146.800 ;
        RECT 44.600 144.800 46.500 145.100 ;
      LAYER metal3 ;
        RECT -2.600 147.100 -2.200 147.200 ;
        RECT 0.600 147.100 1.000 147.200 ;
        RECT -2.600 146.800 1.000 147.100 ;
        RECT 0.600 145.100 1.000 145.200 ;
        RECT 31.000 145.100 31.400 145.200 ;
        RECT 44.600 145.100 45.000 145.200 ;
        RECT 0.600 144.800 45.000 145.100 ;
      LAYER via3 ;
        RECT 0.600 146.800 1.000 147.200 ;
      LAYER metal4 ;
        RECT 0.600 146.800 1.000 147.200 ;
        RECT 0.600 145.200 0.900 146.800 ;
        RECT 0.600 144.800 1.000 145.200 ;
    END
  END address[4]
  PIN dataout[0]
    PORT
      LAYER metal1 ;
        RECT 45.400 215.900 45.800 219.900 ;
        RECT 45.400 214.800 45.700 215.900 ;
        RECT 45.400 211.100 45.800 214.800 ;
      LAYER via1 ;
        RECT 45.400 218.800 45.800 219.200 ;
      LAYER metal2 ;
        RECT 46.200 242.800 46.600 243.200 ;
        RECT 46.200 224.100 46.500 242.800 ;
        RECT 45.400 223.800 46.500 224.100 ;
        RECT 45.400 219.200 45.700 223.800 ;
        RECT 45.400 218.800 45.800 219.200 ;
    END
  END dataout[0]
  PIN dataout[1]
    PORT
      LAYER metal1 ;
        RECT 92.600 155.900 93.000 159.900 ;
        RECT 92.700 154.800 93.000 155.900 ;
        RECT 92.600 151.100 93.000 154.800 ;
      LAYER via1 ;
        RECT 92.600 158.800 93.000 159.200 ;
      LAYER metal2 ;
        RECT 91.800 242.800 92.200 243.200 ;
        RECT 91.800 240.200 92.100 242.800 ;
        RECT 91.800 239.800 92.200 240.200 ;
        RECT 92.600 165.800 93.000 166.200 ;
        RECT 92.600 159.200 92.900 165.800 ;
        RECT 92.600 158.800 93.000 159.200 ;
      LAYER metal3 ;
        RECT 91.800 240.100 92.200 240.200 ;
        RECT 92.600 240.100 93.000 240.200 ;
        RECT 91.800 239.800 93.000 240.100 ;
        RECT 91.800 166.100 92.200 166.200 ;
        RECT 92.600 166.100 93.000 166.200 ;
        RECT 91.800 165.800 93.000 166.100 ;
      LAYER via3 ;
        RECT 92.600 239.800 93.000 240.200 ;
      LAYER metal4 ;
        RECT 92.600 240.100 93.000 240.200 ;
        RECT 91.800 239.800 93.000 240.100 ;
        RECT 91.800 166.200 92.100 239.800 ;
        RECT 91.800 165.800 92.200 166.200 ;
    END
  END dataout[1]
  PIN dataout[2]
    PORT
      LAYER metal1 ;
        RECT 88.600 235.900 89.000 239.900 ;
        RECT 88.600 234.800 88.900 235.900 ;
        RECT 88.600 231.100 89.000 234.800 ;
      LAYER via1 ;
        RECT 88.600 238.800 89.000 239.200 ;
      LAYER metal2 ;
        RECT 89.400 243.100 89.800 243.200 ;
        RECT 88.600 242.800 89.800 243.100 ;
        RECT 88.600 239.200 88.900 242.800 ;
        RECT 88.600 238.800 89.000 239.200 ;
    END
  END dataout[2]
  PIN dataout[3]
    PORT
      LAYER metal1 ;
        RECT 231.000 106.200 231.400 109.900 ;
        RECT 231.100 105.100 231.400 106.200 ;
        RECT 231.000 101.100 231.400 105.100 ;
      LAYER via1 ;
        RECT 231.000 103.800 231.400 104.200 ;
      LAYER metal2 ;
        RECT 231.000 104.800 231.400 105.200 ;
        RECT 231.000 104.200 231.300 104.800 ;
        RECT 231.000 103.800 231.400 104.200 ;
      LAYER metal3 ;
        RECT 231.000 105.100 231.400 105.200 ;
        RECT 255.000 105.100 255.400 105.200 ;
        RECT 231.000 104.800 255.400 105.100 ;
    END
  END dataout[3]
  PIN dataout[4]
    PORT
      LAYER metal1 ;
        RECT 0.600 46.200 1.000 49.900 ;
        RECT 0.600 45.100 0.900 46.200 ;
        RECT 0.600 41.100 1.000 45.100 ;
      LAYER via1 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal2 ;
        RECT 0.600 44.800 1.000 45.200 ;
        RECT 0.600 44.200 0.900 44.800 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal3 ;
        RECT -2.600 45.100 -2.200 45.200 ;
        RECT 0.600 45.100 1.000 45.200 ;
        RECT -2.600 44.800 1.000 45.100 ;
    END
  END dataout[4]
  PIN dataout[5]
    PORT
      LAYER metal1 ;
        RECT 10.200 75.900 10.600 79.900 ;
        RECT 10.200 74.800 10.500 75.900 ;
        RECT 10.200 71.100 10.600 74.800 ;
      LAYER via1 ;
        RECT 10.200 76.800 10.600 77.200 ;
      LAYER metal2 ;
        RECT 10.200 76.800 10.600 77.200 ;
        RECT 10.200 75.200 10.500 76.800 ;
        RECT 10.200 74.800 10.600 75.200 ;
      LAYER metal3 ;
        RECT -2.600 75.100 -2.200 75.200 ;
        RECT 10.200 75.100 10.600 75.200 ;
        RECT -2.600 74.800 10.600 75.100 ;
    END
  END dataout[5]
  PIN dataout[6]
    PORT
      LAYER metal1 ;
        RECT 52.600 15.900 53.000 19.900 ;
        RECT 52.700 14.800 53.000 15.900 ;
        RECT 52.600 11.100 53.000 14.800 ;
      LAYER via1 ;
        RECT 52.600 11.800 53.000 12.200 ;
      LAYER metal2 ;
        RECT 52.600 11.800 53.000 12.200 ;
        RECT 52.600 10.100 52.900 11.800 ;
        RECT 51.800 9.800 52.900 10.100 ;
        RECT 51.800 -1.800 52.100 9.800 ;
        RECT 51.800 -2.200 52.200 -1.800 ;
    END
  END dataout[6]
  PIN dataout[7]
    PORT
      LAYER metal1 ;
        RECT 154.200 235.900 154.600 239.900 ;
        RECT 154.200 234.800 154.500 235.900 ;
        RECT 154.200 231.100 154.600 234.800 ;
      LAYER via1 ;
        RECT 154.200 238.800 154.600 239.200 ;
      LAYER metal2 ;
        RECT 155.000 243.100 155.400 243.200 ;
        RECT 154.200 242.800 155.400 243.100 ;
        RECT 154.200 239.200 154.500 242.800 ;
        RECT 154.200 238.800 154.600 239.200 ;
    END
  END dataout[7]
  OBS
      LAYER metal1 ;
        RECT 1.900 236.300 2.300 239.900 ;
        RECT 1.400 235.900 2.300 236.300 ;
        RECT 3.000 235.900 3.400 239.900 ;
        RECT 3.800 236.200 4.200 239.900 ;
        RECT 5.400 236.200 5.800 239.900 ;
        RECT 3.800 235.900 5.800 236.200 ;
        RECT 7.500 236.200 7.900 239.900 ;
        RECT 8.200 236.800 8.600 237.200 ;
        RECT 8.300 236.200 8.600 236.800 ;
        RECT 7.500 235.900 8.000 236.200 ;
        RECT 8.300 235.900 9.000 236.200 ;
        RECT 1.500 234.200 1.800 235.900 ;
        RECT 2.200 234.800 2.600 235.600 ;
        RECT 3.100 235.200 3.400 235.900 ;
        RECT 5.000 235.200 5.400 235.400 ;
        RECT 3.000 234.900 4.200 235.200 ;
        RECT 5.000 235.100 5.800 235.200 ;
        RECT 5.000 234.900 6.500 235.100 ;
        RECT 3.000 234.800 3.400 234.900 ;
        RECT 1.400 233.800 1.800 234.200 ;
        RECT 0.600 232.400 1.000 233.200 ;
        RECT 1.500 233.100 1.800 233.800 ;
        RECT 3.000 233.100 3.400 233.200 ;
        RECT 3.900 233.100 4.200 234.900 ;
        RECT 5.400 234.800 6.500 234.900 ;
        RECT 4.600 233.800 5.000 234.600 ;
        RECT 6.200 234.200 6.500 234.800 ;
        RECT 7.000 234.400 7.400 235.200 ;
        RECT 7.700 234.200 8.000 235.900 ;
        RECT 8.600 235.800 9.000 235.900 ;
        RECT 9.400 235.800 9.800 236.600 ;
        RECT 8.600 235.100 8.900 235.800 ;
        RECT 10.200 235.100 10.600 239.900 ;
        RECT 11.000 237.100 11.400 237.200 ;
        RECT 11.800 237.100 12.200 239.900 ;
        RECT 13.900 237.900 14.500 239.900 ;
        RECT 16.200 237.900 16.600 239.900 ;
        RECT 18.400 238.200 18.800 239.900 ;
        RECT 18.400 237.900 19.400 238.200 ;
        RECT 14.200 237.500 14.600 237.900 ;
        RECT 16.300 237.600 16.600 237.900 ;
        RECT 15.900 237.300 17.700 237.600 ;
        RECT 19.000 237.500 19.400 237.900 ;
        RECT 15.900 237.200 16.300 237.300 ;
        RECT 17.300 237.200 17.700 237.300 ;
        RECT 11.000 236.800 12.200 237.100 ;
        RECT 8.600 234.800 10.600 235.100 ;
        RECT 6.200 234.100 6.600 234.200 ;
        RECT 7.700 234.100 9.000 234.200 ;
        RECT 9.400 234.100 9.800 234.200 ;
        RECT 6.200 233.800 7.000 234.100 ;
        RECT 7.700 233.800 9.800 234.100 ;
        RECT 6.600 233.600 7.000 233.800 ;
        RECT 6.300 233.100 8.100 233.300 ;
        RECT 8.600 233.100 8.900 233.800 ;
        RECT 10.200 233.100 10.600 234.800 ;
        RECT 11.800 235.600 12.200 236.800 ;
        RECT 13.800 236.600 14.500 237.000 ;
        RECT 14.200 236.100 14.500 236.600 ;
        RECT 15.300 236.500 16.400 236.800 ;
        RECT 15.300 236.400 15.700 236.500 ;
        RECT 14.200 235.800 15.400 236.100 ;
        RECT 11.800 235.300 13.900 235.600 ;
        RECT 11.000 233.400 11.400 234.200 ;
        RECT 11.800 233.600 12.200 235.300 ;
        RECT 13.500 235.200 13.900 235.300 ;
        RECT 12.700 234.900 13.100 235.000 ;
        RECT 12.700 234.600 14.600 234.900 ;
        RECT 14.200 234.500 14.600 234.600 ;
        RECT 15.100 234.200 15.400 235.800 ;
        RECT 16.100 235.900 16.400 236.500 ;
        RECT 16.700 236.500 17.100 236.600 ;
        RECT 19.000 236.500 19.400 236.600 ;
        RECT 16.700 236.200 19.400 236.500 ;
        RECT 16.100 235.700 18.500 235.900 ;
        RECT 20.600 235.700 21.000 239.900 ;
        RECT 22.200 236.400 22.600 239.900 ;
        RECT 16.100 235.600 21.000 235.700 ;
        RECT 18.100 235.500 21.000 235.600 ;
        RECT 18.200 235.400 21.000 235.500 ;
        RECT 22.100 235.900 22.600 236.400 ;
        RECT 23.800 236.200 24.200 239.900 ;
        RECT 22.900 235.900 24.200 236.200 ;
        RECT 17.400 235.100 17.800 235.200 ;
        RECT 17.400 234.800 19.900 235.100 ;
        RECT 19.500 234.700 19.900 234.800 ;
        RECT 18.700 234.200 19.100 234.300 ;
        RECT 22.100 234.200 22.400 235.900 ;
        RECT 22.900 234.900 23.200 235.900 ;
        RECT 25.400 235.600 25.800 239.900 ;
        RECT 27.000 235.600 27.400 239.900 ;
        RECT 29.900 236.200 30.300 239.900 ;
        RECT 30.600 236.800 31.000 237.200 ;
        RECT 30.700 236.200 31.000 236.800 ;
        RECT 29.900 235.900 30.400 236.200 ;
        RECT 30.700 235.900 31.400 236.200 ;
        RECT 25.400 235.200 27.400 235.600 ;
        RECT 22.700 234.500 23.200 234.900 ;
        RECT 15.100 234.100 20.600 234.200 ;
        RECT 21.400 234.100 21.800 234.200 ;
        RECT 15.100 233.900 21.800 234.100 ;
        RECT 15.300 233.800 15.700 233.900 ;
        RECT 1.400 232.800 3.400 233.100 ;
        RECT 1.500 232.100 1.800 232.800 ;
        RECT 3.100 232.400 3.500 232.800 ;
        RECT 1.400 231.100 1.800 232.100 ;
        RECT 3.800 231.100 4.200 233.100 ;
        RECT 6.200 233.000 8.200 233.100 ;
        RECT 6.200 231.100 6.600 233.000 ;
        RECT 7.800 231.100 8.200 233.000 ;
        RECT 8.600 231.100 9.000 233.100 ;
        RECT 9.700 232.800 10.600 233.100 ;
        RECT 11.800 233.300 13.700 233.600 ;
        RECT 9.700 231.100 10.100 232.800 ;
        RECT 11.800 231.100 12.200 233.300 ;
        RECT 13.300 233.200 13.700 233.300 ;
        RECT 18.200 232.800 18.500 233.900 ;
        RECT 19.800 233.800 21.800 233.900 ;
        RECT 22.100 233.800 22.600 234.200 ;
        RECT 17.300 232.700 17.700 232.800 ;
        RECT 14.200 232.100 14.600 232.500 ;
        RECT 16.300 232.400 17.700 232.700 ;
        RECT 18.200 232.400 18.600 232.800 ;
        RECT 16.300 232.100 16.600 232.400 ;
        RECT 19.000 232.100 19.400 232.500 ;
        RECT 13.900 231.800 14.600 232.100 ;
        RECT 13.900 231.100 14.500 231.800 ;
        RECT 16.200 231.100 16.600 232.100 ;
        RECT 18.400 231.800 19.400 232.100 ;
        RECT 18.400 231.100 18.800 231.800 ;
        RECT 20.600 231.100 21.000 233.500 ;
        RECT 22.100 233.100 22.400 233.800 ;
        RECT 22.900 233.700 23.200 234.500 ;
        RECT 23.700 235.100 24.200 235.200 ;
        RECT 25.400 235.100 25.800 235.200 ;
        RECT 23.700 234.800 25.800 235.100 ;
        RECT 23.700 234.400 24.100 234.800 ;
        RECT 27.000 233.800 27.400 235.200 ;
        RECT 29.400 234.400 29.800 235.200 ;
        RECT 30.100 234.200 30.400 235.900 ;
        RECT 31.000 235.800 31.400 235.900 ;
        RECT 31.800 235.800 32.200 236.600 ;
        RECT 31.000 235.100 31.300 235.800 ;
        RECT 32.600 235.100 33.000 239.900 ;
        RECT 34.200 235.700 34.600 239.900 ;
        RECT 36.400 238.200 36.800 239.900 ;
        RECT 35.800 237.900 36.800 238.200 ;
        RECT 38.600 237.900 39.000 239.900 ;
        RECT 40.700 237.900 41.300 239.900 ;
        RECT 35.800 237.500 36.200 237.900 ;
        RECT 38.600 237.600 38.900 237.900 ;
        RECT 37.500 237.300 39.300 237.600 ;
        RECT 40.600 237.500 41.000 237.900 ;
        RECT 37.500 237.200 37.900 237.300 ;
        RECT 38.900 237.200 39.300 237.300 ;
        RECT 35.800 236.500 36.200 236.600 ;
        RECT 38.100 236.500 38.500 236.600 ;
        RECT 35.800 236.200 38.500 236.500 ;
        RECT 38.800 236.500 39.900 236.800 ;
        RECT 38.800 235.900 39.100 236.500 ;
        RECT 39.500 236.400 39.900 236.500 ;
        RECT 40.700 236.600 41.400 237.000 ;
        RECT 40.700 236.100 41.000 236.600 ;
        RECT 36.700 235.700 39.100 235.900 ;
        RECT 34.200 235.600 39.100 235.700 ;
        RECT 39.800 235.800 41.000 236.100 ;
        RECT 34.200 235.500 37.100 235.600 ;
        RECT 34.200 235.400 37.000 235.500 ;
        RECT 37.400 235.100 37.800 235.200 ;
        RECT 31.000 234.800 33.000 235.100 ;
        RECT 28.600 234.100 29.000 234.200 ;
        RECT 30.100 234.100 31.400 234.200 ;
        RECT 31.800 234.100 32.200 234.200 ;
        RECT 28.600 233.800 29.400 234.100 ;
        RECT 30.100 233.800 32.200 234.100 ;
        RECT 22.900 233.400 24.200 233.700 ;
        RECT 22.100 232.800 22.600 233.100 ;
        RECT 22.200 231.100 22.600 232.800 ;
        RECT 23.800 231.100 24.200 233.400 ;
        RECT 25.400 233.400 27.400 233.800 ;
        RECT 29.000 233.600 29.400 233.800 ;
        RECT 25.400 231.100 25.800 233.400 ;
        RECT 27.000 231.100 27.400 233.400 ;
        RECT 28.700 233.100 30.500 233.300 ;
        RECT 31.000 233.100 31.300 233.800 ;
        RECT 32.600 233.100 33.000 234.800 ;
        RECT 35.300 234.800 37.800 235.100 ;
        RECT 35.300 234.700 35.700 234.800 ;
        RECT 36.600 234.700 37.000 234.800 ;
        RECT 36.100 234.200 36.500 234.300 ;
        RECT 39.800 234.200 40.100 235.800 ;
        RECT 43.000 235.600 43.400 239.900 ;
        RECT 41.300 235.300 43.400 235.600 ;
        RECT 41.300 235.200 41.700 235.300 ;
        RECT 42.100 234.900 42.500 235.000 ;
        RECT 40.600 234.600 42.500 234.900 ;
        RECT 40.600 234.500 41.000 234.600 ;
        RECT 33.400 233.400 33.800 234.200 ;
        RECT 34.600 233.900 40.100 234.200 ;
        RECT 34.600 233.800 35.400 233.900 ;
        RECT 28.600 233.000 30.600 233.100 ;
        RECT 28.600 231.100 29.000 233.000 ;
        RECT 30.200 231.100 30.600 233.000 ;
        RECT 31.000 231.100 31.400 233.100 ;
        RECT 32.100 232.800 33.000 233.100 ;
        RECT 32.100 231.100 32.500 232.800 ;
        RECT 34.200 231.100 34.600 233.500 ;
        RECT 36.700 232.800 37.000 233.900 ;
        RECT 37.400 233.800 37.800 233.900 ;
        RECT 39.500 233.800 39.900 233.900 ;
        RECT 43.000 233.600 43.400 235.300 ;
        RECT 41.500 233.300 43.400 233.600 ;
        RECT 41.500 233.200 41.900 233.300 ;
        RECT 35.800 232.100 36.200 232.500 ;
        RECT 36.600 232.400 37.000 232.800 ;
        RECT 37.500 232.700 37.900 232.800 ;
        RECT 37.500 232.400 38.900 232.700 ;
        RECT 38.600 232.100 38.900 232.400 ;
        RECT 40.600 232.100 41.000 232.500 ;
        RECT 35.800 231.800 36.800 232.100 ;
        RECT 36.400 231.100 36.800 231.800 ;
        RECT 38.600 231.100 39.000 232.100 ;
        RECT 40.600 231.800 41.300 232.100 ;
        RECT 40.700 231.100 41.300 231.800 ;
        RECT 43.000 231.100 43.400 233.300 ;
        RECT 45.400 235.600 45.800 239.900 ;
        RECT 47.500 237.900 48.100 239.900 ;
        RECT 49.800 237.900 50.200 239.900 ;
        RECT 52.000 238.200 52.400 239.900 ;
        RECT 52.000 237.900 53.000 238.200 ;
        RECT 47.800 237.500 48.200 237.900 ;
        RECT 49.900 237.600 50.200 237.900 ;
        RECT 49.500 237.300 51.300 237.600 ;
        RECT 52.600 237.500 53.000 237.900 ;
        RECT 49.500 237.200 49.900 237.300 ;
        RECT 50.900 237.200 51.300 237.300 ;
        RECT 47.400 236.600 48.100 237.000 ;
        RECT 47.800 236.100 48.100 236.600 ;
        RECT 48.900 236.500 50.000 236.800 ;
        RECT 48.900 236.400 49.300 236.500 ;
        RECT 47.800 235.800 49.000 236.100 ;
        RECT 45.400 235.300 47.500 235.600 ;
        RECT 45.400 233.600 45.800 235.300 ;
        RECT 47.100 235.200 47.500 235.300 ;
        RECT 46.300 234.900 46.700 235.000 ;
        RECT 46.300 234.600 48.200 234.900 ;
        RECT 47.800 234.500 48.200 234.600 ;
        RECT 48.700 234.200 49.000 235.800 ;
        RECT 49.700 235.900 50.000 236.500 ;
        RECT 50.300 236.500 50.700 236.600 ;
        RECT 52.600 236.500 53.000 236.600 ;
        RECT 50.300 236.200 53.000 236.500 ;
        RECT 49.700 235.700 52.100 235.900 ;
        RECT 54.200 235.700 54.600 239.900 ;
        RECT 55.000 237.100 55.400 237.200 ;
        RECT 55.800 237.100 56.200 239.900 ;
        RECT 55.000 236.800 56.200 237.100 ;
        RECT 49.700 235.600 54.600 235.700 ;
        RECT 51.700 235.500 54.600 235.600 ;
        RECT 51.800 235.400 54.600 235.500 ;
        RECT 51.000 235.100 51.400 235.200 ;
        RECT 51.000 234.800 53.500 235.100 ;
        RECT 51.800 234.700 52.200 234.800 ;
        RECT 53.100 234.700 53.500 234.800 ;
        RECT 52.300 234.200 52.700 234.300 ;
        RECT 48.700 233.900 54.200 234.200 ;
        RECT 48.900 233.800 49.300 233.900 ;
        RECT 45.400 233.300 47.300 233.600 ;
        RECT 45.400 231.100 45.800 233.300 ;
        RECT 46.900 233.200 47.300 233.300 ;
        RECT 51.800 232.800 52.100 233.900 ;
        RECT 53.400 233.800 54.200 233.900 ;
        RECT 50.900 232.700 51.300 232.800 ;
        RECT 47.800 232.100 48.200 232.500 ;
        RECT 49.900 232.400 51.300 232.700 ;
        RECT 51.800 232.400 52.200 232.800 ;
        RECT 49.900 232.100 50.200 232.400 ;
        RECT 52.600 232.100 53.000 232.500 ;
        RECT 47.500 231.800 48.200 232.100 ;
        RECT 47.500 231.100 48.100 231.800 ;
        RECT 49.800 231.100 50.200 232.100 ;
        RECT 52.000 231.800 53.000 232.100 ;
        RECT 52.000 231.100 52.400 231.800 ;
        RECT 54.200 231.100 54.600 233.500 ;
        RECT 55.000 233.400 55.400 234.200 ;
        RECT 55.800 233.100 56.200 236.800 ;
        RECT 57.800 236.800 58.200 237.200 ;
        RECT 56.600 235.800 57.000 236.600 ;
        RECT 57.800 236.200 58.100 236.800 ;
        RECT 58.500 236.200 58.900 239.900 ;
        RECT 57.400 235.900 58.100 236.200 ;
        RECT 58.400 235.900 58.900 236.200 ;
        RECT 57.400 235.800 57.800 235.900 ;
        RECT 56.600 235.100 57.000 235.200 ;
        RECT 58.400 235.100 58.700 235.900 ;
        RECT 60.600 235.700 61.000 239.900 ;
        RECT 62.800 238.200 63.200 239.900 ;
        RECT 62.200 237.900 63.200 238.200 ;
        RECT 65.000 237.900 65.400 239.900 ;
        RECT 67.100 237.900 67.700 239.900 ;
        RECT 62.200 237.500 62.600 237.900 ;
        RECT 65.000 237.600 65.300 237.900 ;
        RECT 63.900 237.300 65.700 237.600 ;
        RECT 67.000 237.500 67.400 237.900 ;
        RECT 63.900 237.200 64.300 237.300 ;
        RECT 65.300 237.200 65.700 237.300 ;
        RECT 69.400 237.100 69.800 239.900 ;
        RECT 70.200 237.100 70.600 237.200 ;
        RECT 62.200 236.500 62.600 236.600 ;
        RECT 64.500 236.500 64.900 236.600 ;
        RECT 62.200 236.200 64.900 236.500 ;
        RECT 65.200 236.500 66.300 236.800 ;
        RECT 65.200 235.900 65.500 236.500 ;
        RECT 65.900 236.400 66.300 236.500 ;
        RECT 67.100 236.600 67.800 237.000 ;
        RECT 69.400 236.800 70.600 237.100 ;
        RECT 67.100 236.100 67.400 236.600 ;
        RECT 63.100 235.700 65.500 235.900 ;
        RECT 60.600 235.600 65.500 235.700 ;
        RECT 66.200 235.800 67.400 236.100 ;
        RECT 60.600 235.500 63.500 235.600 ;
        RECT 60.600 235.400 63.400 235.500 ;
        RECT 56.600 234.800 58.700 235.100 ;
        RECT 58.400 234.200 58.700 234.800 ;
        RECT 59.000 234.400 59.400 235.200 ;
        RECT 63.800 235.100 64.200 235.200 ;
        RECT 61.700 234.800 64.200 235.100 ;
        RECT 61.700 234.700 62.100 234.800 ;
        RECT 62.500 234.200 62.900 234.300 ;
        RECT 66.200 234.200 66.500 235.800 ;
        RECT 69.400 235.600 69.800 236.800 ;
        RECT 67.700 235.300 69.800 235.600 ;
        RECT 67.700 235.200 68.100 235.300 ;
        RECT 68.500 234.900 68.900 235.000 ;
        RECT 67.000 234.600 68.900 234.900 ;
        RECT 67.000 234.500 67.400 234.600 ;
        RECT 57.400 233.800 58.700 234.200 ;
        RECT 59.800 234.100 60.200 234.200 ;
        RECT 59.400 233.800 60.200 234.100 ;
        RECT 61.000 233.900 66.500 234.200 ;
        RECT 61.000 233.800 61.800 233.900 ;
        RECT 57.500 233.100 57.800 233.800 ;
        RECT 59.400 233.600 59.800 233.800 ;
        RECT 58.300 233.100 60.100 233.300 ;
        RECT 55.800 232.800 56.700 233.100 ;
        RECT 56.300 231.100 56.700 232.800 ;
        RECT 57.400 231.100 57.800 233.100 ;
        RECT 58.200 233.000 60.200 233.100 ;
        RECT 58.200 231.100 58.600 233.000 ;
        RECT 59.800 231.100 60.200 233.000 ;
        RECT 60.600 231.100 61.000 233.500 ;
        RECT 63.100 233.200 63.400 233.900 ;
        RECT 65.900 233.800 66.300 233.900 ;
        RECT 69.400 233.600 69.800 235.300 ;
        RECT 71.000 235.100 71.400 239.900 ;
        RECT 73.700 237.200 74.100 239.900 ;
        RECT 73.000 236.800 73.400 237.200 ;
        RECT 73.700 236.800 74.600 237.200 ;
        RECT 71.800 235.800 72.200 236.600 ;
        RECT 73.000 236.200 73.300 236.800 ;
        RECT 73.700 236.200 74.100 236.800 ;
        RECT 72.600 235.900 73.300 236.200 ;
        RECT 73.600 235.900 74.100 236.200 ;
        RECT 72.600 235.800 73.000 235.900 ;
        RECT 72.600 235.100 72.900 235.800 ;
        RECT 71.000 234.800 72.900 235.100 ;
        RECT 67.900 233.300 69.800 233.600 ;
        RECT 70.200 233.400 70.600 234.200 ;
        RECT 67.900 233.200 68.300 233.300 ;
        RECT 62.200 232.100 62.600 232.500 ;
        RECT 63.000 232.400 63.400 233.200 ;
        RECT 63.900 232.700 64.300 232.800 ;
        RECT 63.900 232.400 65.300 232.700 ;
        RECT 65.000 232.100 65.300 232.400 ;
        RECT 67.000 232.100 67.400 232.500 ;
        RECT 62.200 231.800 63.200 232.100 ;
        RECT 62.800 231.100 63.200 231.800 ;
        RECT 65.000 231.100 65.400 232.100 ;
        RECT 67.000 231.800 67.700 232.100 ;
        RECT 67.100 231.100 67.700 231.800 ;
        RECT 69.400 231.100 69.800 233.300 ;
        RECT 71.000 233.100 71.400 234.800 ;
        RECT 73.600 234.200 73.900 235.900 ;
        RECT 75.800 235.600 76.200 239.900 ;
        RECT 77.900 237.900 78.500 239.900 ;
        RECT 80.200 237.900 80.600 239.900 ;
        RECT 82.400 238.200 82.800 239.900 ;
        RECT 82.400 237.900 83.400 238.200 ;
        RECT 78.200 237.500 78.600 237.900 ;
        RECT 80.300 237.600 80.600 237.900 ;
        RECT 79.900 237.300 81.700 237.600 ;
        RECT 83.000 237.500 83.400 237.900 ;
        RECT 79.900 237.200 80.300 237.300 ;
        RECT 81.300 237.200 81.700 237.300 ;
        RECT 77.800 236.600 78.500 237.000 ;
        RECT 78.200 236.100 78.500 236.600 ;
        RECT 79.300 236.500 80.400 236.800 ;
        RECT 79.300 236.400 79.700 236.500 ;
        RECT 78.200 235.800 79.400 236.100 ;
        RECT 75.800 235.300 77.900 235.600 ;
        RECT 74.200 234.400 74.600 235.200 ;
        RECT 72.600 233.800 73.900 234.200 ;
        RECT 75.000 234.100 75.400 234.200 ;
        RECT 74.600 233.800 75.400 234.100 ;
        RECT 72.700 233.100 73.000 233.800 ;
        RECT 74.600 233.600 75.000 233.800 ;
        RECT 75.800 233.600 76.200 235.300 ;
        RECT 77.500 235.200 77.900 235.300 ;
        RECT 76.700 234.900 77.100 235.000 ;
        RECT 76.700 234.600 78.600 234.900 ;
        RECT 78.200 234.500 78.600 234.600 ;
        RECT 79.100 234.200 79.400 235.800 ;
        RECT 80.100 235.900 80.400 236.500 ;
        RECT 80.700 236.500 81.100 236.600 ;
        RECT 83.000 236.500 83.400 236.600 ;
        RECT 80.700 236.200 83.400 236.500 ;
        RECT 80.100 235.700 82.500 235.900 ;
        RECT 84.600 235.700 85.000 239.900 ;
        RECT 85.400 236.200 85.800 239.900 ;
        RECT 87.000 236.400 87.400 239.900 ;
        RECT 85.400 235.900 86.700 236.200 ;
        RECT 87.000 235.900 87.500 236.400 ;
        RECT 90.200 236.200 90.600 239.900 ;
        RECT 80.100 235.600 85.000 235.700 ;
        RECT 82.100 235.500 85.000 235.600 ;
        RECT 82.200 235.400 85.000 235.500 ;
        RECT 81.400 235.100 81.800 235.200 ;
        RECT 81.400 234.800 83.900 235.100 ;
        RECT 85.400 234.800 85.900 235.200 ;
        RECT 82.200 234.700 82.600 234.800 ;
        RECT 83.500 234.700 83.900 234.800 ;
        RECT 85.500 234.400 85.900 234.800 ;
        RECT 86.400 234.900 86.700 235.900 ;
        RECT 86.400 234.500 86.900 234.900 ;
        RECT 82.700 234.200 83.100 234.300 ;
        RECT 79.100 233.900 84.600 234.200 ;
        RECT 79.300 233.800 79.700 233.900 ;
        RECT 75.800 233.300 77.700 233.600 ;
        RECT 73.500 233.100 75.300 233.300 ;
        RECT 71.000 232.800 71.900 233.100 ;
        RECT 71.500 231.100 71.900 232.800 ;
        RECT 72.600 231.100 73.000 233.100 ;
        RECT 73.400 233.000 75.400 233.100 ;
        RECT 73.400 231.100 73.800 233.000 ;
        RECT 75.000 231.100 75.400 233.000 ;
        RECT 75.800 231.100 76.200 233.300 ;
        RECT 77.300 233.200 77.700 233.300 ;
        RECT 82.200 232.800 82.500 233.900 ;
        RECT 83.800 233.800 84.600 233.900 ;
        RECT 86.400 233.700 86.700 234.500 ;
        RECT 87.200 234.200 87.500 235.900 ;
        RECT 89.500 235.900 90.600 236.200 ;
        RECT 89.500 235.600 89.800 235.900 ;
        RECT 89.200 235.200 89.800 235.600 ;
        RECT 91.800 235.600 92.200 239.900 ;
        RECT 93.400 235.600 93.800 239.900 ;
        RECT 95.000 235.600 95.400 239.900 ;
        RECT 96.600 235.600 97.000 239.900 ;
        RECT 99.800 235.700 100.200 239.900 ;
        RECT 102.000 238.200 102.400 239.900 ;
        RECT 101.400 237.900 102.400 238.200 ;
        RECT 104.200 237.900 104.600 239.900 ;
        RECT 106.300 237.900 106.900 239.900 ;
        RECT 101.400 237.500 101.800 237.900 ;
        RECT 104.200 237.600 104.500 237.900 ;
        RECT 103.100 237.300 104.900 237.600 ;
        RECT 106.200 237.500 106.600 237.900 ;
        RECT 103.100 237.200 103.500 237.300 ;
        RECT 104.500 237.200 104.900 237.300 ;
        RECT 101.400 236.500 101.800 236.600 ;
        RECT 103.700 236.500 104.100 236.600 ;
        RECT 101.400 236.200 104.100 236.500 ;
        RECT 104.400 236.500 105.500 236.800 ;
        RECT 104.400 235.900 104.700 236.500 ;
        RECT 105.100 236.400 105.500 236.500 ;
        RECT 106.300 236.600 107.000 237.000 ;
        RECT 106.300 236.100 106.600 236.600 ;
        RECT 102.300 235.700 104.700 235.900 ;
        RECT 99.800 235.600 104.700 235.700 ;
        RECT 105.400 235.800 106.600 236.100 ;
        RECT 91.800 235.200 92.700 235.600 ;
        RECT 93.400 235.200 94.500 235.600 ;
        RECT 95.000 235.200 96.100 235.600 ;
        RECT 96.600 235.200 97.800 235.600 ;
        RECT 99.800 235.500 102.700 235.600 ;
        RECT 99.800 235.400 102.600 235.500 ;
        RECT 87.000 233.800 87.500 234.200 ;
        RECT 81.300 232.700 81.700 232.800 ;
        RECT 78.200 232.100 78.600 232.500 ;
        RECT 80.300 232.400 81.700 232.700 ;
        RECT 82.200 232.400 82.600 232.800 ;
        RECT 80.300 232.100 80.600 232.400 ;
        RECT 83.000 232.100 83.400 232.500 ;
        RECT 77.900 231.800 78.600 232.100 ;
        RECT 77.900 231.100 78.500 231.800 ;
        RECT 80.200 231.100 80.600 232.100 ;
        RECT 82.400 231.800 83.400 232.100 ;
        RECT 82.400 231.100 82.800 231.800 ;
        RECT 84.600 231.100 85.000 233.500 ;
        RECT 85.400 233.400 86.700 233.700 ;
        RECT 85.400 231.100 85.800 233.400 ;
        RECT 87.200 233.100 87.500 233.800 ;
        RECT 89.500 233.700 89.800 235.200 ;
        RECT 90.200 234.400 90.600 235.200 ;
        RECT 92.300 234.500 92.700 235.200 ;
        RECT 94.100 234.500 94.500 235.200 ;
        RECT 95.700 234.500 96.100 235.200 ;
        RECT 91.000 234.100 91.900 234.500 ;
        RECT 92.300 234.100 93.600 234.500 ;
        RECT 94.100 234.100 95.300 234.500 ;
        RECT 95.700 234.100 97.000 234.500 ;
        RECT 97.400 234.100 97.800 235.200 ;
        RECT 103.000 235.100 103.400 235.200 ;
        RECT 104.600 235.100 105.000 235.200 ;
        RECT 100.900 234.800 105.000 235.100 ;
        RECT 100.900 234.700 101.300 234.800 ;
        RECT 101.700 234.200 102.100 234.300 ;
        RECT 105.400 234.200 105.700 235.800 ;
        RECT 108.600 235.600 109.000 239.900 ;
        RECT 110.700 236.200 111.100 239.900 ;
        RECT 111.400 236.800 111.800 237.200 ;
        RECT 111.500 236.200 111.800 236.800 ;
        RECT 110.700 235.900 111.200 236.200 ;
        RECT 111.500 235.900 112.200 236.200 ;
        RECT 106.900 235.300 109.000 235.600 ;
        RECT 106.900 235.200 107.300 235.300 ;
        RECT 107.700 234.900 108.100 235.000 ;
        RECT 106.200 234.600 108.100 234.900 ;
        RECT 106.200 234.500 106.600 234.600 ;
        RECT 98.200 234.100 98.600 234.200 ;
        RECT 91.000 233.800 91.400 234.100 ;
        RECT 92.300 233.800 92.700 234.100 ;
        RECT 94.100 233.800 94.500 234.100 ;
        RECT 95.700 233.800 96.100 234.100 ;
        RECT 97.400 233.800 98.600 234.100 ;
        RECT 100.200 233.900 105.700 234.200 ;
        RECT 100.200 233.800 101.000 233.900 ;
        RECT 89.500 233.400 90.600 233.700 ;
        RECT 87.000 232.800 87.500 233.100 ;
        RECT 87.000 231.100 87.400 232.800 ;
        RECT 90.200 231.100 90.600 233.400 ;
        RECT 91.800 233.400 92.700 233.800 ;
        RECT 93.400 233.400 94.500 233.800 ;
        RECT 95.000 233.400 96.100 233.800 ;
        RECT 96.600 233.400 97.800 233.800 ;
        RECT 91.800 231.100 92.200 233.400 ;
        RECT 93.400 231.100 93.800 233.400 ;
        RECT 95.000 231.100 95.400 233.400 ;
        RECT 96.600 231.100 97.000 233.400 ;
        RECT 99.800 231.100 100.200 233.500 ;
        RECT 102.300 232.800 102.600 233.900 ;
        RECT 105.100 233.800 105.500 233.900 ;
        RECT 108.600 233.600 109.000 235.300 ;
        RECT 110.900 235.200 111.200 235.900 ;
        RECT 111.800 235.800 112.200 235.900 ;
        RECT 113.400 235.600 113.800 239.900 ;
        RECT 115.000 235.600 115.400 239.900 ;
        RECT 113.400 235.200 115.400 235.600 ;
        RECT 116.600 235.700 117.000 239.900 ;
        RECT 118.800 238.200 119.200 239.900 ;
        RECT 118.200 237.900 119.200 238.200 ;
        RECT 121.000 237.900 121.400 239.900 ;
        RECT 123.100 237.900 123.700 239.900 ;
        RECT 118.200 237.500 118.600 237.900 ;
        RECT 121.000 237.600 121.300 237.900 ;
        RECT 119.900 237.300 121.700 237.600 ;
        RECT 123.000 237.500 123.400 237.900 ;
        RECT 119.900 237.200 120.300 237.300 ;
        RECT 121.300 237.200 121.700 237.300 ;
        RECT 125.400 237.100 125.800 239.900 ;
        RECT 126.200 237.100 126.600 237.200 ;
        RECT 118.200 236.500 118.600 236.600 ;
        RECT 120.500 236.500 120.900 236.600 ;
        RECT 118.200 236.200 120.900 236.500 ;
        RECT 121.200 236.500 122.300 236.800 ;
        RECT 121.200 235.900 121.500 236.500 ;
        RECT 121.900 236.400 122.300 236.500 ;
        RECT 123.100 236.600 123.800 237.000 ;
        RECT 125.400 236.800 126.600 237.100 ;
        RECT 123.100 236.100 123.400 236.600 ;
        RECT 119.100 235.700 121.500 235.900 ;
        RECT 116.600 235.600 121.500 235.700 ;
        RECT 122.200 235.800 123.400 236.100 ;
        RECT 116.600 235.500 119.500 235.600 ;
        RECT 116.600 235.400 119.400 235.500 ;
        RECT 110.200 234.400 110.600 235.200 ;
        RECT 110.900 234.800 111.400 235.200 ;
        RECT 110.900 234.200 111.200 234.800 ;
        RECT 109.400 234.100 109.800 234.200 ;
        RECT 109.400 233.800 110.200 234.100 ;
        RECT 110.900 233.800 112.200 234.200 ;
        RECT 113.400 233.800 113.800 235.200 ;
        RECT 119.800 235.100 120.200 235.200 ;
        RECT 117.700 234.800 120.200 235.100 ;
        RECT 117.700 234.700 118.100 234.800 ;
        RECT 118.500 234.200 118.900 234.300 ;
        RECT 122.200 234.200 122.500 235.800 ;
        RECT 125.400 235.600 125.800 236.800 ;
        RECT 123.700 235.300 125.800 235.600 ;
        RECT 123.700 235.200 124.100 235.300 ;
        RECT 124.500 234.900 124.900 235.000 ;
        RECT 123.000 234.600 124.900 234.900 ;
        RECT 123.000 234.500 123.400 234.600 ;
        RECT 117.000 233.900 122.500 234.200 ;
        RECT 117.000 233.800 117.800 233.900 ;
        RECT 109.800 233.600 110.200 233.800 ;
        RECT 107.100 233.300 109.000 233.600 ;
        RECT 107.100 233.200 107.500 233.300 ;
        RECT 101.400 232.100 101.800 232.500 ;
        RECT 102.200 232.400 102.600 232.800 ;
        RECT 103.100 232.700 103.500 232.800 ;
        RECT 103.100 232.400 104.500 232.700 ;
        RECT 104.200 232.100 104.500 232.400 ;
        RECT 106.200 232.100 106.600 232.500 ;
        RECT 101.400 231.800 102.400 232.100 ;
        RECT 102.000 231.100 102.400 231.800 ;
        RECT 104.200 231.100 104.600 232.100 ;
        RECT 106.200 231.800 106.900 232.100 ;
        RECT 106.300 231.100 106.900 231.800 ;
        RECT 108.600 231.100 109.000 233.300 ;
        RECT 109.500 233.100 111.300 233.300 ;
        RECT 111.800 233.100 112.100 233.800 ;
        RECT 113.400 233.400 115.400 233.800 ;
        RECT 109.400 233.000 111.400 233.100 ;
        RECT 109.400 231.100 109.800 233.000 ;
        RECT 111.000 231.100 111.400 233.000 ;
        RECT 111.800 231.100 112.200 233.100 ;
        RECT 113.400 231.100 113.800 233.400 ;
        RECT 115.000 231.100 115.400 233.400 ;
        RECT 116.600 231.100 117.000 233.500 ;
        RECT 119.100 232.800 119.400 233.900 ;
        RECT 121.900 233.800 122.300 233.900 ;
        RECT 125.400 233.600 125.800 235.300 ;
        RECT 127.000 235.100 127.400 239.900 ;
        RECT 129.000 236.800 129.400 237.200 ;
        RECT 127.800 235.800 128.200 236.600 ;
        RECT 129.000 236.200 129.300 236.800 ;
        RECT 129.700 236.200 130.100 239.900 ;
        RECT 128.600 235.900 129.300 236.200 ;
        RECT 129.600 235.900 130.100 236.200 ;
        RECT 133.100 236.200 133.500 239.900 ;
        RECT 133.800 236.800 134.200 237.200 ;
        RECT 133.900 236.200 134.200 236.800 ;
        RECT 133.100 235.900 133.600 236.200 ;
        RECT 133.900 235.900 134.600 236.200 ;
        RECT 128.600 235.800 129.000 235.900 ;
        RECT 128.600 235.100 128.900 235.800 ;
        RECT 127.000 234.800 128.900 235.100 ;
        RECT 123.900 233.300 125.800 233.600 ;
        RECT 126.200 233.400 126.600 234.200 ;
        RECT 123.900 233.200 124.300 233.300 ;
        RECT 118.200 232.100 118.600 232.500 ;
        RECT 119.000 232.400 119.400 232.800 ;
        RECT 119.900 232.700 120.300 232.800 ;
        RECT 119.900 232.400 121.300 232.700 ;
        RECT 121.000 232.100 121.300 232.400 ;
        RECT 123.000 232.100 123.400 232.500 ;
        RECT 118.200 231.800 119.200 232.100 ;
        RECT 118.800 231.100 119.200 231.800 ;
        RECT 121.000 231.100 121.400 232.100 ;
        RECT 123.000 231.800 123.700 232.100 ;
        RECT 123.100 231.100 123.700 231.800 ;
        RECT 125.400 231.100 125.800 233.300 ;
        RECT 127.000 233.100 127.400 234.800 ;
        RECT 129.600 234.200 129.900 235.900 ;
        RECT 130.200 234.400 130.600 235.200 ;
        RECT 132.600 234.400 133.000 235.200 ;
        RECT 133.300 234.200 133.600 235.900 ;
        RECT 134.200 235.800 134.600 235.900 ;
        RECT 135.000 235.800 135.400 236.600 ;
        RECT 134.200 235.100 134.500 235.800 ;
        RECT 135.800 235.100 136.200 239.900 ;
        RECT 137.400 235.700 137.800 239.900 ;
        RECT 139.600 238.200 140.000 239.900 ;
        RECT 139.000 237.900 140.000 238.200 ;
        RECT 141.800 237.900 142.200 239.900 ;
        RECT 143.900 237.900 144.500 239.900 ;
        RECT 139.000 237.500 139.400 237.900 ;
        RECT 141.800 237.600 142.100 237.900 ;
        RECT 140.700 237.300 142.500 237.600 ;
        RECT 143.800 237.500 144.200 237.900 ;
        RECT 140.700 237.200 141.100 237.300 ;
        RECT 142.100 237.200 142.500 237.300 ;
        RECT 139.000 236.500 139.400 236.600 ;
        RECT 141.300 236.500 141.700 236.600 ;
        RECT 139.000 236.200 141.700 236.500 ;
        RECT 142.000 236.500 143.100 236.800 ;
        RECT 142.000 235.900 142.300 236.500 ;
        RECT 142.700 236.400 143.100 236.500 ;
        RECT 143.900 236.600 144.600 237.000 ;
        RECT 143.900 236.100 144.200 236.600 ;
        RECT 139.900 235.700 142.300 235.900 ;
        RECT 137.400 235.600 142.300 235.700 ;
        RECT 143.000 235.800 144.200 236.100 ;
        RECT 137.400 235.500 140.300 235.600 ;
        RECT 137.400 235.400 140.200 235.500 ;
        RECT 140.600 235.100 141.000 235.200 ;
        RECT 142.200 235.100 142.600 235.200 ;
        RECT 134.200 234.800 136.200 235.100 ;
        RECT 127.800 234.100 128.200 234.200 ;
        RECT 128.600 234.100 129.900 234.200 ;
        RECT 131.000 234.100 131.400 234.200 ;
        RECT 131.800 234.100 132.200 234.200 ;
        RECT 127.800 233.800 129.900 234.100 ;
        RECT 130.600 233.800 132.600 234.100 ;
        RECT 133.300 233.800 134.600 234.200 ;
        RECT 128.700 233.100 129.000 233.800 ;
        RECT 130.600 233.600 131.000 233.800 ;
        RECT 132.200 233.600 132.600 233.800 ;
        RECT 129.500 233.100 131.300 233.300 ;
        RECT 131.900 233.100 133.700 233.300 ;
        RECT 134.200 233.100 134.500 233.800 ;
        RECT 135.800 233.100 136.200 234.800 ;
        RECT 138.500 234.800 142.600 235.100 ;
        RECT 138.500 234.700 138.900 234.800 ;
        RECT 139.300 234.200 139.700 234.300 ;
        RECT 143.000 234.200 143.300 235.800 ;
        RECT 146.200 235.600 146.600 239.900 ;
        RECT 147.000 236.200 147.400 239.900 ;
        RECT 148.600 236.200 149.000 239.900 ;
        RECT 147.000 235.900 149.000 236.200 ;
        RECT 149.400 235.900 149.800 239.900 ;
        RECT 152.100 236.300 152.500 239.900 ;
        RECT 152.100 235.900 153.000 236.300 ;
        RECT 155.800 236.200 156.200 239.900 ;
        RECT 155.100 235.900 156.200 236.200 ;
        RECT 157.900 236.200 158.300 239.900 ;
        RECT 158.600 236.800 159.000 237.200 ;
        RECT 158.700 236.200 159.000 236.800 ;
        RECT 157.900 235.900 158.400 236.200 ;
        RECT 158.700 235.900 159.400 236.200 ;
        RECT 144.500 235.300 146.600 235.600 ;
        RECT 144.500 235.200 144.900 235.300 ;
        RECT 145.300 234.900 145.700 235.000 ;
        RECT 143.800 234.600 145.700 234.900 ;
        RECT 143.800 234.500 144.200 234.600 ;
        RECT 136.600 233.400 137.000 234.200 ;
        RECT 137.800 233.900 143.300 234.200 ;
        RECT 137.800 233.800 138.600 233.900 ;
        RECT 127.000 232.800 127.900 233.100 ;
        RECT 127.500 231.100 127.900 232.800 ;
        RECT 128.600 231.100 129.000 233.100 ;
        RECT 129.400 233.000 131.400 233.100 ;
        RECT 129.400 231.100 129.800 233.000 ;
        RECT 131.000 231.100 131.400 233.000 ;
        RECT 131.800 233.000 133.800 233.100 ;
        RECT 131.800 231.100 132.200 233.000 ;
        RECT 133.400 231.100 133.800 233.000 ;
        RECT 134.200 231.100 134.600 233.100 ;
        RECT 135.300 232.800 136.200 233.100 ;
        RECT 135.300 231.100 135.700 232.800 ;
        RECT 137.400 231.100 137.800 233.500 ;
        RECT 139.900 232.800 140.200 233.900 ;
        RECT 140.600 233.800 141.000 233.900 ;
        RECT 142.700 233.800 143.100 233.900 ;
        RECT 146.200 233.600 146.600 235.300 ;
        RECT 147.400 235.200 147.800 235.400 ;
        RECT 149.400 235.200 149.700 235.900 ;
        RECT 147.000 234.900 147.800 235.200 ;
        RECT 148.600 234.900 149.800 235.200 ;
        RECT 147.000 234.800 147.400 234.900 ;
        RECT 147.800 233.800 148.200 234.600 ;
        RECT 144.700 233.300 146.600 233.600 ;
        RECT 144.700 233.200 145.100 233.300 ;
        RECT 139.000 232.100 139.400 232.500 ;
        RECT 139.800 232.400 140.200 232.800 ;
        RECT 140.700 232.700 141.100 232.800 ;
        RECT 140.700 232.400 142.100 232.700 ;
        RECT 141.800 232.100 142.100 232.400 ;
        RECT 143.800 232.100 144.200 232.500 ;
        RECT 139.000 231.800 140.000 232.100 ;
        RECT 139.600 231.100 140.000 231.800 ;
        RECT 141.800 231.100 142.200 232.100 ;
        RECT 143.800 231.800 144.500 232.100 ;
        RECT 143.900 231.100 144.500 231.800 ;
        RECT 146.200 231.100 146.600 233.300 ;
        RECT 148.600 233.100 148.900 234.900 ;
        RECT 149.400 234.800 149.800 234.900 ;
        RECT 151.800 234.800 152.200 235.600 ;
        RECT 152.600 234.200 152.900 235.900 ;
        RECT 155.100 235.600 155.400 235.900 ;
        RECT 154.800 235.200 155.400 235.600 ;
        RECT 152.600 233.800 153.000 234.200 ;
        RECT 149.400 233.100 149.800 233.200 ;
        RECT 152.600 233.100 152.900 233.800 ;
        RECT 155.100 233.700 155.400 235.200 ;
        RECT 155.800 234.400 156.200 235.200 ;
        RECT 156.600 235.100 157.000 235.200 ;
        RECT 157.400 235.100 157.800 235.200 ;
        RECT 156.600 234.800 157.800 235.100 ;
        RECT 157.400 234.400 157.800 234.800 ;
        RECT 158.100 234.200 158.400 235.900 ;
        RECT 159.000 235.800 159.400 235.900 ;
        RECT 159.800 235.800 160.200 236.600 ;
        RECT 159.000 235.100 159.300 235.800 ;
        RECT 160.600 235.100 161.000 239.900 ;
        RECT 161.400 237.100 161.800 237.200 ;
        RECT 162.200 237.100 162.600 239.900 ;
        RECT 164.300 237.900 164.900 239.900 ;
        RECT 166.600 237.900 167.000 239.900 ;
        RECT 168.800 238.200 169.200 239.900 ;
        RECT 168.800 237.900 169.800 238.200 ;
        RECT 164.600 237.500 165.000 237.900 ;
        RECT 166.700 237.600 167.000 237.900 ;
        RECT 166.300 237.300 168.100 237.600 ;
        RECT 169.400 237.500 169.800 237.900 ;
        RECT 166.300 237.200 166.700 237.300 ;
        RECT 167.700 237.200 168.100 237.300 ;
        RECT 161.400 236.800 162.600 237.100 ;
        RECT 159.000 234.800 161.000 235.100 ;
        RECT 156.600 234.100 157.000 234.200 ;
        RECT 158.100 234.100 159.400 234.200 ;
        RECT 159.800 234.100 160.200 234.200 ;
        RECT 156.600 233.800 157.400 234.100 ;
        RECT 158.100 233.800 160.200 234.100 ;
        RECT 155.100 233.400 156.200 233.700 ;
        RECT 157.000 233.600 157.400 233.800 ;
        RECT 148.600 231.100 149.000 233.100 ;
        RECT 149.400 232.800 152.900 233.100 ;
        RECT 149.300 232.400 149.700 232.800 ;
        RECT 152.600 232.100 152.900 232.800 ;
        RECT 153.400 232.400 153.800 233.200 ;
        RECT 152.600 231.100 153.000 232.100 ;
        RECT 155.800 231.100 156.200 233.400 ;
        RECT 156.700 233.100 158.500 233.300 ;
        RECT 159.000 233.100 159.300 233.800 ;
        RECT 160.600 233.100 161.000 234.800 ;
        RECT 162.200 235.600 162.600 236.800 ;
        RECT 164.200 236.600 164.900 237.000 ;
        RECT 164.600 236.100 164.900 236.600 ;
        RECT 165.700 236.500 166.800 236.800 ;
        RECT 165.700 236.400 166.100 236.500 ;
        RECT 164.600 235.800 165.800 236.100 ;
        RECT 162.200 235.300 164.300 235.600 ;
        RECT 161.400 233.400 161.800 234.200 ;
        RECT 162.200 233.600 162.600 235.300 ;
        RECT 163.900 235.200 164.300 235.300 ;
        RECT 163.100 234.900 163.500 235.000 ;
        RECT 163.100 234.600 165.000 234.900 ;
        RECT 164.600 234.500 165.000 234.600 ;
        RECT 165.500 234.200 165.800 235.800 ;
        RECT 166.500 235.900 166.800 236.500 ;
        RECT 167.100 236.500 167.500 236.600 ;
        RECT 169.400 236.500 169.800 236.600 ;
        RECT 167.100 236.200 169.800 236.500 ;
        RECT 166.500 235.700 168.900 235.900 ;
        RECT 171.000 235.700 171.400 239.900 ;
        RECT 166.500 235.600 171.400 235.700 ;
        RECT 168.500 235.500 171.400 235.600 ;
        RECT 168.600 235.400 171.400 235.500 ;
        RECT 171.800 235.600 172.200 239.900 ;
        RECT 173.900 237.900 174.500 239.900 ;
        RECT 176.200 237.900 176.600 239.900 ;
        RECT 178.400 238.200 178.800 239.900 ;
        RECT 178.400 237.900 179.400 238.200 ;
        RECT 174.200 237.500 174.600 237.900 ;
        RECT 176.300 237.600 176.600 237.900 ;
        RECT 175.900 237.300 177.700 237.600 ;
        RECT 179.000 237.500 179.400 237.900 ;
        RECT 175.900 237.200 176.300 237.300 ;
        RECT 177.300 237.200 177.700 237.300 ;
        RECT 173.800 236.600 174.500 237.000 ;
        RECT 174.200 236.100 174.500 236.600 ;
        RECT 175.300 236.500 176.400 236.800 ;
        RECT 175.300 236.400 175.700 236.500 ;
        RECT 174.200 235.800 175.400 236.100 ;
        RECT 171.800 235.300 173.900 235.600 ;
        RECT 167.800 235.100 168.200 235.200 ;
        RECT 167.800 234.800 170.300 235.100 ;
        RECT 169.900 234.700 170.300 234.800 ;
        RECT 169.100 234.200 169.500 234.300 ;
        RECT 165.500 233.900 171.000 234.200 ;
        RECT 165.700 233.800 166.100 233.900 ;
        RECT 156.600 233.000 158.600 233.100 ;
        RECT 156.600 231.100 157.000 233.000 ;
        RECT 158.200 231.100 158.600 233.000 ;
        RECT 159.000 231.100 159.400 233.100 ;
        RECT 160.100 232.800 161.000 233.100 ;
        RECT 162.200 233.300 164.100 233.600 ;
        RECT 160.100 231.100 160.500 232.800 ;
        RECT 162.200 231.100 162.600 233.300 ;
        RECT 163.700 233.200 164.100 233.300 ;
        RECT 168.600 232.800 168.900 233.900 ;
        RECT 170.200 233.800 171.000 233.900 ;
        RECT 171.800 233.600 172.200 235.300 ;
        RECT 173.500 235.200 173.900 235.300 ;
        RECT 172.700 234.900 173.100 235.000 ;
        RECT 172.700 234.600 174.600 234.900 ;
        RECT 174.200 234.500 174.600 234.600 ;
        RECT 175.100 234.200 175.400 235.800 ;
        RECT 176.100 235.900 176.400 236.500 ;
        RECT 176.700 236.500 177.100 236.600 ;
        RECT 179.000 236.500 179.400 236.600 ;
        RECT 176.700 236.200 179.400 236.500 ;
        RECT 176.100 235.700 178.500 235.900 ;
        RECT 180.600 235.700 181.000 239.900 ;
        RECT 176.100 235.600 181.000 235.700 ;
        RECT 178.100 235.500 181.000 235.600 ;
        RECT 178.200 235.400 181.000 235.500 ;
        RECT 181.400 235.700 181.800 239.900 ;
        RECT 183.600 238.200 184.000 239.900 ;
        RECT 183.000 237.900 184.000 238.200 ;
        RECT 185.800 237.900 186.200 239.900 ;
        RECT 187.900 237.900 188.500 239.900 ;
        RECT 183.000 237.500 183.400 237.900 ;
        RECT 185.800 237.600 186.100 237.900 ;
        RECT 184.700 237.300 186.500 237.600 ;
        RECT 187.800 237.500 188.200 237.900 ;
        RECT 184.700 237.200 185.100 237.300 ;
        RECT 186.100 237.200 186.500 237.300 ;
        RECT 183.000 236.500 183.400 236.600 ;
        RECT 185.300 236.500 185.700 236.600 ;
        RECT 183.000 236.200 185.700 236.500 ;
        RECT 186.000 236.500 187.100 236.800 ;
        RECT 186.000 235.900 186.300 236.500 ;
        RECT 186.700 236.400 187.100 236.500 ;
        RECT 187.900 236.600 188.600 237.000 ;
        RECT 187.900 236.100 188.200 236.600 ;
        RECT 183.900 235.700 186.300 235.900 ;
        RECT 181.400 235.600 186.300 235.700 ;
        RECT 187.000 235.800 188.200 236.100 ;
        RECT 181.400 235.500 184.300 235.600 ;
        RECT 181.400 235.400 184.200 235.500 ;
        RECT 177.400 235.100 177.800 235.200 ;
        RECT 184.600 235.100 185.000 235.200 ;
        RECT 177.400 234.800 179.900 235.100 ;
        RECT 178.200 234.700 178.600 234.800 ;
        RECT 179.500 234.700 179.900 234.800 ;
        RECT 182.500 234.800 185.000 235.100 ;
        RECT 182.500 234.700 182.900 234.800 ;
        RECT 178.700 234.200 179.100 234.300 ;
        RECT 183.300 234.200 183.700 234.300 ;
        RECT 187.000 234.200 187.300 235.800 ;
        RECT 190.200 235.600 190.600 239.900 ;
        RECT 192.300 236.200 192.700 239.900 ;
        RECT 193.000 236.800 193.400 237.200 ;
        RECT 193.100 236.200 193.400 236.800 ;
        RECT 191.800 235.800 192.800 236.200 ;
        RECT 193.100 235.900 193.800 236.200 ;
        RECT 193.400 235.800 193.800 235.900 ;
        RECT 188.500 235.300 190.600 235.600 ;
        RECT 188.500 235.200 188.900 235.300 ;
        RECT 189.300 234.900 189.700 235.000 ;
        RECT 187.800 234.600 189.700 234.900 ;
        RECT 187.800 234.500 188.200 234.600 ;
        RECT 175.100 234.100 180.600 234.200 ;
        RECT 181.800 234.100 187.300 234.200 ;
        RECT 175.100 233.900 187.300 234.100 ;
        RECT 175.300 233.800 175.700 233.900 ;
        RECT 167.700 232.700 168.100 232.800 ;
        RECT 164.600 232.100 165.000 232.500 ;
        RECT 166.700 232.400 168.100 232.700 ;
        RECT 168.600 232.400 169.000 232.800 ;
        RECT 166.700 232.100 167.000 232.400 ;
        RECT 169.400 232.100 169.800 232.500 ;
        RECT 164.300 231.800 165.000 232.100 ;
        RECT 164.300 231.100 164.900 231.800 ;
        RECT 166.600 231.100 167.000 232.100 ;
        RECT 168.800 231.800 169.800 232.100 ;
        RECT 168.800 231.100 169.200 231.800 ;
        RECT 171.000 231.100 171.400 233.500 ;
        RECT 171.800 233.300 173.700 233.600 ;
        RECT 171.800 231.100 172.200 233.300 ;
        RECT 173.300 233.200 173.700 233.300 ;
        RECT 178.200 232.800 178.500 233.900 ;
        RECT 179.800 233.800 182.600 233.900 ;
        RECT 177.300 232.700 177.700 232.800 ;
        RECT 174.200 232.100 174.600 232.500 ;
        RECT 176.300 232.400 177.700 232.700 ;
        RECT 178.200 232.400 178.600 232.800 ;
        RECT 176.300 232.100 176.600 232.400 ;
        RECT 179.000 232.100 179.400 232.500 ;
        RECT 173.900 231.800 174.600 232.100 ;
        RECT 173.900 231.100 174.500 231.800 ;
        RECT 176.200 231.100 176.600 232.100 ;
        RECT 178.400 231.800 179.400 232.100 ;
        RECT 178.400 231.100 178.800 231.800 ;
        RECT 180.600 231.100 181.000 233.500 ;
        RECT 181.400 231.100 181.800 233.500 ;
        RECT 183.900 232.800 184.200 233.900 ;
        RECT 185.400 233.800 185.800 233.900 ;
        RECT 186.700 233.800 187.100 233.900 ;
        RECT 190.200 233.600 190.600 235.300 ;
        RECT 191.800 234.400 192.200 235.200 ;
        RECT 192.500 234.200 192.800 235.800 ;
        RECT 194.200 235.700 194.600 239.900 ;
        RECT 196.400 238.200 196.800 239.900 ;
        RECT 195.800 237.900 196.800 238.200 ;
        RECT 198.600 237.900 199.000 239.900 ;
        RECT 200.700 237.900 201.300 239.900 ;
        RECT 195.800 237.500 196.200 237.900 ;
        RECT 198.600 237.600 198.900 237.900 ;
        RECT 197.500 237.300 199.300 237.600 ;
        RECT 200.600 237.500 201.000 237.900 ;
        RECT 197.500 237.200 197.900 237.300 ;
        RECT 198.900 237.200 199.300 237.300 ;
        RECT 203.000 237.100 203.400 239.900 ;
        RECT 205.400 237.100 205.800 237.200 ;
        RECT 195.800 236.500 196.200 236.600 ;
        RECT 198.100 236.500 198.500 236.600 ;
        RECT 195.800 236.200 198.500 236.500 ;
        RECT 198.800 236.500 199.900 236.800 ;
        RECT 198.800 235.900 199.100 236.500 ;
        RECT 199.500 236.400 199.900 236.500 ;
        RECT 200.700 236.600 201.400 237.000 ;
        RECT 203.000 236.800 205.800 237.100 ;
        RECT 200.700 236.100 201.000 236.600 ;
        RECT 196.700 235.700 199.100 235.900 ;
        RECT 194.200 235.600 199.100 235.700 ;
        RECT 199.800 235.800 201.000 236.100 ;
        RECT 194.200 235.500 197.100 235.600 ;
        RECT 194.200 235.400 197.000 235.500 ;
        RECT 197.400 235.100 197.800 235.200 ;
        RECT 199.000 235.100 199.400 235.200 ;
        RECT 195.300 234.800 199.400 235.100 ;
        RECT 195.300 234.700 195.700 234.800 ;
        RECT 196.100 234.200 196.500 234.300 ;
        RECT 199.800 234.200 200.100 235.800 ;
        RECT 203.000 235.600 203.400 236.800 ;
        RECT 201.300 235.300 203.400 235.600 ;
        RECT 201.300 235.200 201.700 235.300 ;
        RECT 202.100 234.900 202.500 235.000 ;
        RECT 200.600 234.600 202.500 234.900 ;
        RECT 200.600 234.500 201.000 234.600 ;
        RECT 191.000 234.100 191.400 234.200 ;
        RECT 191.000 233.800 191.800 234.100 ;
        RECT 192.500 233.800 193.800 234.200 ;
        RECT 194.600 233.900 200.100 234.200 ;
        RECT 194.600 233.800 195.400 233.900 ;
        RECT 191.400 233.600 191.800 233.800 ;
        RECT 188.700 233.300 190.600 233.600 ;
        RECT 188.700 233.200 189.100 233.300 ;
        RECT 183.000 232.100 183.400 232.500 ;
        RECT 183.800 232.400 184.200 232.800 ;
        RECT 184.700 232.700 185.100 232.800 ;
        RECT 184.700 232.400 186.100 232.700 ;
        RECT 185.800 232.100 186.100 232.400 ;
        RECT 187.800 232.100 188.200 232.500 ;
        RECT 183.000 231.800 184.000 232.100 ;
        RECT 183.600 231.100 184.000 231.800 ;
        RECT 185.800 231.100 186.200 232.100 ;
        RECT 187.800 231.800 188.500 232.100 ;
        RECT 187.900 231.100 188.500 231.800 ;
        RECT 190.200 231.100 190.600 233.300 ;
        RECT 191.100 233.100 192.900 233.300 ;
        RECT 193.400 233.100 193.700 233.800 ;
        RECT 191.000 233.000 193.000 233.100 ;
        RECT 191.000 231.100 191.400 233.000 ;
        RECT 192.600 231.100 193.000 233.000 ;
        RECT 193.400 231.100 193.800 233.100 ;
        RECT 194.200 231.100 194.600 233.500 ;
        RECT 196.700 232.800 197.000 233.900 ;
        RECT 198.200 233.800 198.600 233.900 ;
        RECT 199.500 233.800 199.900 233.900 ;
        RECT 203.000 233.600 203.400 235.300 ;
        RECT 206.200 235.100 206.600 239.900 ;
        RECT 208.200 236.800 208.600 237.200 ;
        RECT 207.000 235.800 207.400 236.600 ;
        RECT 208.200 236.200 208.500 236.800 ;
        RECT 208.900 236.200 209.300 239.900 ;
        RECT 207.800 235.900 208.500 236.200 ;
        RECT 208.800 235.900 209.300 236.200 ;
        RECT 207.800 235.800 208.200 235.900 ;
        RECT 207.800 235.100 208.100 235.800 ;
        RECT 208.800 235.200 209.100 235.900 ;
        RECT 211.000 235.700 211.400 239.900 ;
        RECT 213.200 238.200 213.600 239.900 ;
        RECT 212.600 237.900 213.600 238.200 ;
        RECT 215.400 237.900 215.800 239.900 ;
        RECT 217.500 237.900 218.100 239.900 ;
        RECT 212.600 237.500 213.000 237.900 ;
        RECT 215.400 237.600 215.700 237.900 ;
        RECT 214.300 237.300 216.100 237.600 ;
        RECT 217.400 237.500 217.800 237.900 ;
        RECT 214.300 237.200 214.700 237.300 ;
        RECT 215.700 237.200 216.100 237.300 ;
        RECT 212.600 236.500 213.000 236.600 ;
        RECT 214.900 236.500 215.300 236.600 ;
        RECT 212.600 236.200 215.300 236.500 ;
        RECT 215.600 236.500 216.700 236.800 ;
        RECT 215.600 235.900 215.900 236.500 ;
        RECT 216.300 236.400 216.700 236.500 ;
        RECT 217.500 236.600 218.200 237.000 ;
        RECT 217.500 236.100 217.800 236.600 ;
        RECT 213.500 235.700 215.900 235.900 ;
        RECT 211.000 235.600 215.900 235.700 ;
        RECT 216.600 235.800 217.800 236.100 ;
        RECT 211.000 235.500 213.900 235.600 ;
        RECT 211.000 235.400 213.800 235.500 ;
        RECT 206.200 234.800 208.100 235.100 ;
        RECT 208.600 234.800 209.100 235.200 ;
        RECT 201.500 233.300 203.400 233.600 ;
        RECT 205.400 233.400 205.800 234.200 ;
        RECT 201.500 233.200 201.900 233.300 ;
        RECT 195.800 232.100 196.200 232.500 ;
        RECT 196.600 232.400 197.000 232.800 ;
        RECT 197.500 232.700 197.900 232.800 ;
        RECT 197.500 232.400 198.900 232.700 ;
        RECT 198.600 232.100 198.900 232.400 ;
        RECT 200.600 232.100 201.000 232.500 ;
        RECT 195.800 231.800 196.800 232.100 ;
        RECT 196.400 231.100 196.800 231.800 ;
        RECT 198.600 231.100 199.000 232.100 ;
        RECT 200.600 231.800 201.300 232.100 ;
        RECT 200.700 231.100 201.300 231.800 ;
        RECT 203.000 231.100 203.400 233.300 ;
        RECT 206.200 233.100 206.600 234.800 ;
        RECT 208.800 234.200 209.100 234.800 ;
        RECT 209.400 234.400 209.800 235.200 ;
        RECT 214.200 235.100 214.600 235.200 ;
        RECT 212.100 234.800 214.600 235.100 ;
        RECT 212.100 234.700 212.500 234.800 ;
        RECT 213.400 234.700 213.800 234.800 ;
        RECT 212.900 234.200 213.300 234.300 ;
        RECT 216.600 234.200 216.900 235.800 ;
        RECT 219.800 235.600 220.200 239.900 ;
        RECT 220.600 235.800 221.000 236.600 ;
        RECT 218.100 235.300 220.200 235.600 ;
        RECT 218.100 235.200 218.500 235.300 ;
        RECT 218.900 234.900 219.300 235.000 ;
        RECT 217.400 234.600 219.300 234.900 ;
        RECT 217.400 234.500 217.800 234.600 ;
        RECT 207.800 233.800 209.100 234.200 ;
        RECT 210.200 234.100 210.600 234.200 ;
        RECT 209.800 233.800 210.600 234.100 ;
        RECT 211.400 233.900 216.900 234.200 ;
        RECT 211.400 233.800 212.200 233.900 ;
        RECT 207.900 233.100 208.200 233.800 ;
        RECT 209.800 233.600 210.200 233.800 ;
        RECT 208.700 233.100 210.500 233.300 ;
        RECT 206.200 232.800 207.100 233.100 ;
        RECT 206.700 231.100 207.100 232.800 ;
        RECT 207.800 231.100 208.200 233.100 ;
        RECT 208.600 233.000 210.600 233.100 ;
        RECT 208.600 231.100 209.000 233.000 ;
        RECT 210.200 231.100 210.600 233.000 ;
        RECT 211.000 231.100 211.400 233.500 ;
        RECT 213.500 232.800 213.800 233.900 ;
        RECT 214.200 233.800 214.600 233.900 ;
        RECT 216.300 233.800 216.700 233.900 ;
        RECT 219.800 233.600 220.200 235.300 ;
        RECT 218.300 233.300 220.200 233.600 ;
        RECT 218.300 233.200 218.700 233.300 ;
        RECT 212.600 232.100 213.000 232.500 ;
        RECT 213.400 232.400 213.800 232.800 ;
        RECT 214.300 232.700 214.700 232.800 ;
        RECT 214.300 232.400 215.700 232.700 ;
        RECT 215.400 232.100 215.700 232.400 ;
        RECT 217.400 232.100 217.800 232.500 ;
        RECT 212.600 231.800 213.600 232.100 ;
        RECT 213.200 231.100 213.600 231.800 ;
        RECT 215.400 231.100 215.800 232.100 ;
        RECT 217.400 231.800 218.100 232.100 ;
        RECT 217.500 231.100 218.100 231.800 ;
        RECT 219.800 231.100 220.200 233.300 ;
        RECT 221.400 233.100 221.800 239.900 ;
        RECT 223.000 235.700 223.400 239.900 ;
        RECT 225.200 238.200 225.600 239.900 ;
        RECT 224.600 237.900 225.600 238.200 ;
        RECT 227.400 237.900 227.800 239.900 ;
        RECT 229.500 237.900 230.100 239.900 ;
        RECT 224.600 237.500 225.000 237.900 ;
        RECT 227.400 237.600 227.700 237.900 ;
        RECT 226.300 237.300 228.100 237.600 ;
        RECT 229.400 237.500 229.800 237.900 ;
        RECT 226.300 237.200 226.700 237.300 ;
        RECT 227.700 237.200 228.100 237.300 ;
        RECT 224.600 236.500 225.000 236.600 ;
        RECT 226.900 236.500 227.300 236.600 ;
        RECT 224.600 236.200 227.300 236.500 ;
        RECT 227.600 236.500 228.700 236.800 ;
        RECT 227.600 235.900 227.900 236.500 ;
        RECT 228.300 236.400 228.700 236.500 ;
        RECT 229.500 236.600 230.200 237.000 ;
        RECT 229.500 236.100 229.800 236.600 ;
        RECT 225.500 235.700 227.900 235.900 ;
        RECT 223.000 235.600 227.900 235.700 ;
        RECT 228.600 235.800 229.800 236.100 ;
        RECT 223.000 235.500 225.900 235.600 ;
        RECT 223.000 235.400 225.800 235.500 ;
        RECT 226.200 235.100 226.600 235.200 ;
        RECT 224.100 234.800 226.600 235.100 ;
        RECT 224.100 234.700 224.500 234.800 ;
        RECT 224.900 234.200 225.300 234.300 ;
        RECT 228.600 234.200 228.900 235.800 ;
        RECT 231.800 235.600 232.200 239.900 ;
        RECT 230.100 235.300 232.200 235.600 ;
        RECT 232.600 235.700 233.000 239.900 ;
        RECT 234.800 238.200 235.200 239.900 ;
        RECT 234.200 237.900 235.200 238.200 ;
        RECT 237.000 237.900 237.400 239.900 ;
        RECT 239.100 237.900 239.700 239.900 ;
        RECT 234.200 237.500 234.600 237.900 ;
        RECT 237.000 237.600 237.300 237.900 ;
        RECT 235.900 237.300 237.700 237.600 ;
        RECT 239.000 237.500 239.400 237.900 ;
        RECT 235.900 237.200 236.300 237.300 ;
        RECT 237.300 237.200 237.700 237.300 ;
        RECT 234.200 236.500 234.600 236.600 ;
        RECT 236.500 236.500 236.900 236.600 ;
        RECT 234.200 236.200 236.900 236.500 ;
        RECT 237.200 236.500 238.300 236.800 ;
        RECT 237.200 235.900 237.500 236.500 ;
        RECT 237.900 236.400 238.300 236.500 ;
        RECT 239.100 236.600 239.800 237.000 ;
        RECT 239.100 236.100 239.400 236.600 ;
        RECT 235.100 235.700 237.500 235.900 ;
        RECT 232.600 235.600 237.500 235.700 ;
        RECT 238.200 235.800 239.400 236.100 ;
        RECT 232.600 235.500 235.500 235.600 ;
        RECT 232.600 235.400 235.400 235.500 ;
        RECT 230.100 235.200 230.500 235.300 ;
        RECT 230.900 234.900 231.300 235.000 ;
        RECT 229.400 234.600 231.300 234.900 ;
        RECT 229.400 234.500 229.800 234.600 ;
        RECT 222.200 233.400 222.600 234.200 ;
        RECT 223.400 233.900 228.900 234.200 ;
        RECT 223.400 233.800 224.200 233.900 ;
        RECT 220.900 232.800 221.800 233.100 ;
        RECT 220.900 232.200 221.300 232.800 ;
        RECT 220.900 231.800 221.800 232.200 ;
        RECT 220.900 231.100 221.300 231.800 ;
        RECT 223.000 231.100 223.400 233.500 ;
        RECT 225.500 232.800 225.800 233.900 ;
        RECT 228.300 233.800 228.700 233.900 ;
        RECT 231.800 233.600 232.200 235.300 ;
        RECT 235.800 235.100 236.200 235.200 ;
        RECT 233.700 234.800 236.200 235.100 ;
        RECT 233.700 234.700 234.100 234.800 ;
        RECT 234.500 234.200 234.900 234.300 ;
        RECT 238.200 234.200 238.500 235.800 ;
        RECT 241.400 235.600 241.800 239.900 ;
        RECT 239.700 235.300 241.800 235.600 ;
        RECT 239.700 235.200 240.100 235.300 ;
        RECT 240.500 234.900 240.900 235.000 ;
        RECT 239.000 234.600 240.900 234.900 ;
        RECT 239.000 234.500 239.400 234.600 ;
        RECT 233.000 233.900 238.500 234.200 ;
        RECT 233.000 233.800 233.800 233.900 ;
        RECT 230.300 233.300 232.200 233.600 ;
        RECT 230.300 233.200 230.700 233.300 ;
        RECT 224.600 232.100 225.000 232.500 ;
        RECT 225.400 232.400 225.800 232.800 ;
        RECT 226.300 232.700 226.700 232.800 ;
        RECT 226.300 232.400 227.700 232.700 ;
        RECT 227.400 232.100 227.700 232.400 ;
        RECT 229.400 232.100 229.800 232.500 ;
        RECT 224.600 231.800 225.600 232.100 ;
        RECT 225.200 231.100 225.600 231.800 ;
        RECT 227.400 231.100 227.800 232.100 ;
        RECT 229.400 231.800 230.100 232.100 ;
        RECT 229.500 231.100 230.100 231.800 ;
        RECT 231.800 231.100 232.200 233.300 ;
        RECT 232.600 231.100 233.000 233.500 ;
        RECT 235.100 232.800 235.400 233.900 ;
        RECT 237.900 233.800 238.300 233.900 ;
        RECT 241.400 233.600 241.800 235.300 ;
        RECT 239.900 233.300 241.800 233.600 ;
        RECT 239.900 233.200 240.300 233.300 ;
        RECT 234.200 232.100 234.600 232.500 ;
        RECT 235.000 232.400 235.400 232.800 ;
        RECT 235.900 232.700 236.300 232.800 ;
        RECT 235.900 232.400 237.300 232.700 ;
        RECT 237.000 232.100 237.300 232.400 ;
        RECT 239.000 232.100 239.400 232.500 ;
        RECT 234.200 231.800 235.200 232.100 ;
        RECT 234.800 231.100 235.200 231.800 ;
        RECT 237.000 231.100 237.400 232.100 ;
        RECT 239.000 231.800 239.700 232.100 ;
        RECT 239.100 231.100 239.700 231.800 ;
        RECT 241.400 231.100 241.800 233.300 ;
        RECT 243.000 235.600 243.400 239.900 ;
        RECT 244.600 235.600 245.000 239.900 ;
        RECT 247.500 236.200 247.900 239.900 ;
        RECT 248.200 236.800 248.600 237.200 ;
        RECT 248.300 236.200 248.600 236.800 ;
        RECT 247.500 235.900 248.000 236.200 ;
        RECT 248.300 235.900 249.000 236.200 ;
        RECT 243.000 235.200 245.000 235.600 ;
        RECT 243.000 233.800 243.400 235.200 ;
        RECT 247.000 234.400 247.400 235.200 ;
        RECT 247.700 234.200 248.000 235.900 ;
        RECT 248.600 235.800 249.000 235.900 ;
        RECT 249.400 235.800 249.800 236.600 ;
        RECT 248.600 235.100 248.900 235.800 ;
        RECT 250.200 235.100 250.600 239.900 ;
        RECT 248.600 234.800 250.600 235.100 ;
        RECT 246.200 234.100 246.600 234.200 ;
        RECT 246.200 233.800 247.000 234.100 ;
        RECT 247.700 233.800 249.000 234.200 ;
        RECT 243.000 233.400 245.000 233.800 ;
        RECT 246.600 233.600 247.000 233.800 ;
        RECT 243.000 231.100 243.400 233.400 ;
        RECT 244.600 231.100 245.000 233.400 ;
        RECT 246.300 233.100 248.100 233.300 ;
        RECT 248.600 233.100 248.900 233.800 ;
        RECT 250.200 233.100 250.600 234.800 ;
        RECT 251.000 233.400 251.400 234.200 ;
        RECT 246.200 233.000 248.200 233.100 ;
        RECT 246.200 231.100 246.600 233.000 ;
        RECT 247.800 231.100 248.200 233.000 ;
        RECT 248.600 231.100 249.000 233.100 ;
        RECT 249.700 232.800 250.600 233.100 ;
        RECT 249.700 231.100 250.100 232.800 ;
        RECT 0.600 227.700 1.000 229.900 ;
        RECT 2.700 229.200 3.300 229.900 ;
        RECT 2.700 228.900 3.400 229.200 ;
        RECT 5.000 228.900 5.400 229.900 ;
        RECT 7.200 229.200 7.600 229.900 ;
        RECT 7.200 228.900 8.200 229.200 ;
        RECT 3.000 228.500 3.400 228.900 ;
        RECT 5.100 228.600 5.400 228.900 ;
        RECT 5.100 228.300 6.500 228.600 ;
        RECT 6.100 228.200 6.500 228.300 ;
        RECT 7.000 228.200 7.400 228.600 ;
        RECT 7.800 228.500 8.200 228.900 ;
        RECT 2.100 227.700 2.500 227.800 ;
        RECT 0.600 227.400 2.500 227.700 ;
        RECT 0.600 225.700 1.000 227.400 ;
        RECT 4.100 227.100 4.500 227.200 ;
        RECT 7.000 227.100 7.300 228.200 ;
        RECT 9.400 227.500 9.800 229.900 ;
        RECT 11.000 227.600 11.400 229.900 ;
        RECT 12.600 227.600 13.000 229.900 ;
        RECT 14.200 227.600 14.600 229.900 ;
        RECT 15.800 227.600 16.200 229.900 ;
        RECT 17.400 228.000 17.800 229.900 ;
        RECT 19.000 228.000 19.400 229.900 ;
        RECT 17.400 227.900 19.400 228.000 ;
        RECT 19.800 227.900 20.200 229.900 ;
        RECT 20.900 228.200 21.300 229.900 ;
        RECT 20.900 227.900 21.800 228.200 ;
        RECT 17.500 227.700 19.300 227.900 ;
        RECT 10.200 227.200 11.400 227.600 ;
        RECT 11.900 227.200 13.000 227.600 ;
        RECT 13.500 227.200 14.600 227.600 ;
        RECT 15.300 227.200 16.200 227.600 ;
        RECT 17.800 227.200 18.200 227.400 ;
        RECT 19.800 227.200 20.100 227.900 ;
        RECT 8.600 227.100 9.400 227.200 ;
        RECT 3.900 226.800 9.400 227.100 ;
        RECT 3.000 226.400 3.400 226.500 ;
        RECT 1.500 226.100 3.400 226.400 ;
        RECT 1.500 226.000 1.900 226.100 ;
        RECT 2.300 225.700 2.700 225.800 ;
        RECT 0.600 225.400 2.700 225.700 ;
        RECT 0.600 221.100 1.000 225.400 ;
        RECT 3.900 225.200 4.200 226.800 ;
        RECT 7.500 226.700 7.900 226.800 ;
        RECT 8.300 226.200 8.700 226.300 ;
        RECT 4.600 226.100 5.000 226.200 ;
        RECT 6.200 226.100 8.700 226.200 ;
        RECT 4.600 225.900 8.700 226.100 ;
        RECT 4.600 225.800 6.600 225.900 ;
        RECT 10.200 225.800 10.600 227.200 ;
        RECT 11.900 226.900 12.300 227.200 ;
        RECT 13.500 226.900 13.900 227.200 ;
        RECT 15.300 226.900 15.700 227.200 ;
        RECT 16.600 226.900 17.000 227.200 ;
        RECT 11.000 226.500 12.300 226.900 ;
        RECT 12.700 226.500 13.900 226.900 ;
        RECT 14.400 226.500 15.700 226.900 ;
        RECT 16.100 226.500 17.000 226.900 ;
        RECT 17.400 226.900 18.200 227.200 ;
        RECT 17.400 226.800 17.800 226.900 ;
        RECT 18.900 226.800 20.200 227.200 ;
        RECT 11.900 225.800 12.300 226.500 ;
        RECT 13.500 225.800 13.900 226.500 ;
        RECT 15.300 225.800 15.700 226.500 ;
        RECT 18.200 225.800 18.600 226.600 ;
        RECT 7.000 225.500 9.800 225.600 ;
        RECT 6.900 225.400 9.800 225.500 ;
        RECT 10.200 225.400 11.400 225.800 ;
        RECT 11.900 225.400 13.000 225.800 ;
        RECT 13.500 225.400 14.600 225.800 ;
        RECT 15.300 225.400 16.200 225.800 ;
        RECT 3.000 224.900 4.200 225.200 ;
        RECT 4.900 225.300 9.800 225.400 ;
        RECT 4.900 225.100 7.300 225.300 ;
        RECT 3.000 224.400 3.300 224.900 ;
        RECT 2.600 224.000 3.300 224.400 ;
        RECT 4.100 224.500 4.500 224.600 ;
        RECT 4.900 224.500 5.200 225.100 ;
        RECT 4.100 224.200 5.200 224.500 ;
        RECT 5.500 224.500 8.200 224.800 ;
        RECT 5.500 224.400 5.900 224.500 ;
        RECT 7.800 224.400 8.200 224.500 ;
        RECT 4.700 223.700 5.100 223.800 ;
        RECT 6.100 223.700 6.500 223.800 ;
        RECT 3.000 223.100 3.400 223.500 ;
        RECT 4.700 223.400 6.500 223.700 ;
        RECT 5.100 223.100 5.400 223.400 ;
        RECT 7.800 223.100 8.200 223.500 ;
        RECT 2.700 221.100 3.300 223.100 ;
        RECT 5.000 221.100 5.400 223.100 ;
        RECT 7.200 222.800 8.200 223.100 ;
        RECT 7.200 221.100 7.600 222.800 ;
        RECT 9.400 221.100 9.800 225.300 ;
        RECT 11.000 221.100 11.400 225.400 ;
        RECT 12.600 221.100 13.000 225.400 ;
        RECT 14.200 221.100 14.600 225.400 ;
        RECT 15.800 221.100 16.200 225.400 ;
        RECT 18.900 225.100 19.200 226.800 ;
        RECT 21.400 226.100 21.800 227.900 ;
        RECT 22.200 226.800 22.600 227.600 ;
        RECT 23.000 227.500 23.400 229.900 ;
        RECT 25.200 229.200 25.600 229.900 ;
        RECT 24.600 228.900 25.600 229.200 ;
        RECT 27.400 228.900 27.800 229.900 ;
        RECT 29.500 229.200 30.100 229.900 ;
        RECT 29.400 228.900 30.100 229.200 ;
        RECT 24.600 228.500 25.000 228.900 ;
        RECT 27.400 228.600 27.700 228.900 ;
        RECT 25.400 228.200 25.800 228.600 ;
        RECT 26.300 228.300 27.700 228.600 ;
        RECT 29.400 228.500 29.800 228.900 ;
        RECT 26.300 228.200 26.700 228.300 ;
        RECT 23.400 227.100 24.200 227.200 ;
        RECT 25.500 227.100 25.800 228.200 ;
        RECT 30.300 227.700 30.700 227.800 ;
        RECT 31.800 227.700 32.200 229.900 ;
        RECT 30.300 227.400 32.200 227.700 ;
        RECT 28.300 227.100 28.700 227.200 ;
        RECT 23.400 226.800 28.900 227.100 ;
        RECT 24.900 226.700 25.300 226.800 ;
        RECT 19.800 225.800 21.800 226.100 ;
        RECT 24.100 226.200 24.500 226.300 ;
        RECT 25.400 226.200 25.800 226.300 ;
        RECT 28.600 226.200 28.900 226.800 ;
        RECT 29.400 226.400 29.800 226.500 ;
        RECT 24.100 225.900 26.600 226.200 ;
        RECT 26.200 225.800 26.600 225.900 ;
        RECT 28.600 225.800 29.000 226.200 ;
        RECT 29.400 226.100 31.300 226.400 ;
        RECT 30.900 226.000 31.300 226.100 ;
        RECT 19.800 225.200 20.100 225.800 ;
        RECT 19.800 225.100 20.200 225.200 ;
        RECT 18.700 224.800 19.200 225.100 ;
        RECT 19.500 224.800 20.200 225.100 ;
        RECT 18.700 221.100 19.100 224.800 ;
        RECT 19.500 224.200 19.800 224.800 ;
        RECT 20.600 224.400 21.000 225.200 ;
        RECT 19.400 223.800 19.800 224.200 ;
        RECT 21.400 221.100 21.800 225.800 ;
        RECT 23.000 225.500 25.800 225.600 ;
        RECT 23.000 225.400 25.900 225.500 ;
        RECT 23.000 225.300 27.900 225.400 ;
        RECT 23.000 221.100 23.400 225.300 ;
        RECT 25.500 225.100 27.900 225.300 ;
        RECT 24.600 224.500 27.300 224.800 ;
        RECT 24.600 224.400 25.000 224.500 ;
        RECT 26.900 224.400 27.300 224.500 ;
        RECT 27.600 224.500 27.900 225.100 ;
        RECT 28.600 225.200 28.900 225.800 ;
        RECT 30.100 225.700 30.500 225.800 ;
        RECT 31.800 225.700 32.200 227.400 ;
        RECT 32.600 228.500 33.000 229.500 ;
        RECT 32.600 227.400 32.900 228.500 ;
        RECT 34.700 228.000 35.100 229.500 ;
        RECT 37.400 228.000 37.800 229.900 ;
        RECT 39.000 228.000 39.400 229.900 ;
        RECT 34.700 227.700 35.500 228.000 ;
        RECT 37.400 227.900 39.400 228.000 ;
        RECT 39.800 227.900 40.200 229.900 ;
        RECT 40.900 228.200 41.300 229.900 ;
        RECT 40.900 227.900 41.800 228.200 ;
        RECT 37.500 227.700 39.300 227.900 ;
        RECT 35.100 227.500 35.500 227.700 ;
        RECT 32.600 227.100 34.700 227.400 ;
        RECT 34.200 226.900 34.700 227.100 ;
        RECT 35.200 227.200 35.500 227.500 ;
        RECT 37.800 227.200 38.200 227.400 ;
        RECT 39.800 227.200 40.100 227.900 ;
        RECT 32.600 225.800 33.000 226.600 ;
        RECT 33.400 225.800 33.800 226.600 ;
        RECT 34.200 226.500 34.900 226.900 ;
        RECT 35.200 226.800 36.200 227.200 ;
        RECT 36.600 227.100 37.000 227.200 ;
        RECT 37.400 227.100 38.200 227.200 ;
        RECT 36.600 226.900 38.200 227.100 ;
        RECT 38.900 227.100 40.200 227.200 ;
        RECT 40.600 227.100 41.000 227.200 ;
        RECT 36.600 226.800 37.800 226.900 ;
        RECT 38.900 226.800 41.000 227.100 ;
        RECT 30.100 225.400 32.200 225.700 ;
        RECT 34.200 225.500 34.500 226.500 ;
        RECT 35.200 226.200 35.500 226.800 ;
        RECT 35.000 225.800 35.500 226.200 ;
        RECT 28.600 224.900 29.800 225.200 ;
        RECT 28.300 224.500 28.700 224.600 ;
        RECT 27.600 224.200 28.700 224.500 ;
        RECT 29.500 224.400 29.800 224.900 ;
        RECT 29.500 224.000 30.200 224.400 ;
        RECT 26.300 223.700 26.700 223.800 ;
        RECT 27.700 223.700 28.100 223.800 ;
        RECT 24.600 223.100 25.000 223.500 ;
        RECT 26.300 223.400 28.100 223.700 ;
        RECT 27.400 223.100 27.700 223.400 ;
        RECT 29.400 223.100 29.800 223.500 ;
        RECT 24.600 222.800 25.600 223.100 ;
        RECT 25.200 221.100 25.600 222.800 ;
        RECT 27.400 221.100 27.800 223.100 ;
        RECT 29.500 221.100 30.100 223.100 ;
        RECT 31.800 221.100 32.200 225.400 ;
        RECT 32.600 225.200 34.500 225.500 ;
        RECT 32.600 223.500 32.900 225.200 ;
        RECT 35.200 224.900 35.500 225.800 ;
        RECT 35.800 225.400 36.200 226.200 ;
        RECT 38.200 225.800 38.600 226.600 ;
        RECT 38.900 225.100 39.200 226.800 ;
        RECT 41.400 226.100 41.800 227.900 ;
        RECT 42.200 226.800 42.600 227.600 ;
        RECT 43.000 227.500 43.400 229.900 ;
        RECT 45.200 229.200 45.600 229.900 ;
        RECT 44.600 228.900 45.600 229.200 ;
        RECT 47.400 228.900 47.800 229.900 ;
        RECT 49.500 229.200 50.100 229.900 ;
        RECT 49.400 228.900 50.100 229.200 ;
        RECT 44.600 228.500 45.000 228.900 ;
        RECT 47.400 228.600 47.700 228.900 ;
        RECT 45.400 228.200 45.800 228.600 ;
        RECT 46.300 228.300 47.700 228.600 ;
        RECT 49.400 228.500 49.800 228.900 ;
        RECT 46.300 228.200 46.700 228.300 ;
        RECT 43.400 227.100 44.200 227.200 ;
        RECT 45.500 227.100 45.800 228.200 ;
        RECT 50.300 227.700 50.700 227.800 ;
        RECT 51.800 227.700 52.200 229.900 ;
        RECT 50.300 227.400 52.200 227.700 ;
        RECT 48.300 227.100 48.700 227.200 ;
        RECT 43.400 226.800 48.900 227.100 ;
        RECT 44.900 226.700 45.300 226.800 ;
        RECT 39.800 225.800 41.800 226.100 ;
        RECT 44.100 226.200 44.500 226.300 ;
        RECT 45.400 226.200 45.800 226.300 ;
        RECT 44.100 225.900 46.600 226.200 ;
        RECT 46.200 225.800 46.600 225.900 ;
        RECT 39.800 225.200 40.100 225.800 ;
        RECT 39.800 225.100 40.200 225.200 ;
        RECT 34.700 224.600 35.500 224.900 ;
        RECT 38.700 224.800 39.200 225.100 ;
        RECT 39.500 224.800 40.200 225.100 ;
        RECT 32.600 221.500 33.000 223.500 ;
        RECT 34.700 221.100 35.100 224.600 ;
        RECT 38.700 221.100 39.100 224.800 ;
        RECT 39.500 224.200 39.800 224.800 ;
        RECT 40.600 224.400 41.000 225.200 ;
        RECT 39.400 223.800 39.800 224.200 ;
        RECT 41.400 221.100 41.800 225.800 ;
        RECT 43.000 225.500 45.800 225.600 ;
        RECT 43.000 225.400 45.900 225.500 ;
        RECT 43.000 225.300 47.900 225.400 ;
        RECT 43.000 221.100 43.400 225.300 ;
        RECT 45.500 225.100 47.900 225.300 ;
        RECT 44.600 224.500 47.300 224.800 ;
        RECT 44.600 224.400 45.000 224.500 ;
        RECT 46.900 224.400 47.300 224.500 ;
        RECT 47.600 224.500 47.900 225.100 ;
        RECT 48.600 225.200 48.900 226.800 ;
        RECT 49.400 226.400 49.800 226.500 ;
        RECT 49.400 226.100 51.300 226.400 ;
        RECT 50.900 226.000 51.300 226.100 ;
        RECT 50.100 225.700 50.500 225.800 ;
        RECT 51.800 225.700 52.200 227.400 ;
        RECT 54.200 228.500 54.600 229.500 ;
        RECT 54.200 227.400 54.500 228.500 ;
        RECT 56.300 228.000 56.700 229.500 ;
        RECT 59.000 228.500 59.400 229.500 ;
        RECT 56.300 227.700 57.100 228.000 ;
        RECT 56.700 227.500 57.100 227.700 ;
        RECT 54.200 227.100 56.300 227.400 ;
        RECT 55.800 226.900 56.300 227.100 ;
        RECT 56.800 227.200 57.100 227.500 ;
        RECT 59.000 227.400 59.300 228.500 ;
        RECT 61.100 228.000 61.500 229.500 ;
        RECT 63.800 228.500 64.200 229.500 ;
        RECT 61.100 227.700 61.900 228.000 ;
        RECT 61.500 227.500 61.900 227.700 ;
        RECT 54.200 225.800 54.600 226.600 ;
        RECT 55.000 225.800 55.400 226.600 ;
        RECT 55.800 226.500 56.500 226.900 ;
        RECT 56.800 226.800 57.800 227.200 ;
        RECT 59.000 227.100 61.100 227.400 ;
        RECT 60.600 226.900 61.100 227.100 ;
        RECT 61.600 227.200 61.900 227.500 ;
        RECT 63.800 227.400 64.100 228.500 ;
        RECT 65.900 228.000 66.300 229.500 ;
        RECT 65.900 227.700 66.700 228.000 ;
        RECT 66.300 227.500 66.700 227.700 ;
        RECT 50.100 225.400 52.200 225.700 ;
        RECT 55.800 225.500 56.100 226.500 ;
        RECT 48.600 224.900 49.800 225.200 ;
        RECT 48.300 224.500 48.700 224.600 ;
        RECT 47.600 224.200 48.700 224.500 ;
        RECT 49.500 224.400 49.800 224.900 ;
        RECT 49.500 224.000 50.200 224.400 ;
        RECT 46.300 223.700 46.700 223.800 ;
        RECT 47.700 223.700 48.100 223.800 ;
        RECT 44.600 223.100 45.000 223.500 ;
        RECT 46.300 223.400 48.100 223.700 ;
        RECT 47.400 223.100 47.700 223.400 ;
        RECT 49.400 223.100 49.800 223.500 ;
        RECT 44.600 222.800 45.600 223.100 ;
        RECT 45.200 221.100 45.600 222.800 ;
        RECT 47.400 221.100 47.800 223.100 ;
        RECT 49.500 221.100 50.100 223.100 ;
        RECT 51.800 221.100 52.200 225.400 ;
        RECT 54.200 225.200 56.100 225.500 ;
        RECT 54.200 223.500 54.500 225.200 ;
        RECT 56.800 224.900 57.100 226.800 ;
        RECT 57.400 226.100 57.800 226.200 ;
        RECT 58.200 226.100 58.600 226.200 ;
        RECT 57.400 225.800 58.600 226.100 ;
        RECT 59.000 225.800 59.400 226.600 ;
        RECT 59.800 225.800 60.200 226.600 ;
        RECT 60.600 226.500 61.300 226.900 ;
        RECT 61.600 226.800 62.600 227.200 ;
        RECT 63.800 227.100 65.900 227.400 ;
        RECT 65.400 226.900 65.900 227.100 ;
        RECT 66.400 227.200 66.700 227.500 ;
        RECT 69.400 227.600 69.800 229.900 ;
        RECT 71.000 227.600 71.400 229.900 ;
        RECT 72.600 227.600 73.000 229.900 ;
        RECT 74.200 227.600 74.600 229.900 ;
        RECT 75.800 227.700 76.200 229.900 ;
        RECT 77.900 229.200 78.500 229.900 ;
        RECT 77.900 228.900 78.600 229.200 ;
        RECT 80.200 228.900 80.600 229.900 ;
        RECT 82.400 229.200 82.800 229.900 ;
        RECT 82.400 228.900 83.400 229.200 ;
        RECT 78.200 228.500 78.600 228.900 ;
        RECT 80.300 228.600 80.600 228.900 ;
        RECT 80.300 228.300 81.700 228.600 ;
        RECT 81.300 228.200 81.700 228.300 ;
        RECT 82.200 228.200 82.600 228.600 ;
        RECT 83.000 228.500 83.400 228.900 ;
        RECT 77.300 227.700 77.700 227.800 ;
        RECT 69.400 227.200 70.300 227.600 ;
        RECT 71.000 227.200 72.100 227.600 ;
        RECT 72.600 227.200 73.700 227.600 ;
        RECT 74.200 227.200 75.400 227.600 ;
        RECT 57.400 225.400 57.800 225.800 ;
        RECT 60.600 225.500 60.900 226.500 ;
        RECT 56.300 224.600 57.100 224.900 ;
        RECT 59.000 225.200 60.900 225.500 ;
        RECT 54.200 221.500 54.600 223.500 ;
        RECT 56.300 221.100 56.700 224.600 ;
        RECT 59.000 223.500 59.300 225.200 ;
        RECT 61.600 224.900 61.900 226.800 ;
        RECT 62.200 225.400 62.600 226.200 ;
        RECT 63.800 225.800 64.200 226.600 ;
        RECT 64.600 225.800 65.000 226.600 ;
        RECT 65.400 226.500 66.100 226.900 ;
        RECT 66.400 226.800 67.400 227.200 ;
        RECT 68.600 226.900 69.000 227.200 ;
        RECT 69.900 226.900 70.300 227.200 ;
        RECT 71.700 226.900 72.100 227.200 ;
        RECT 73.300 226.900 73.700 227.200 ;
        RECT 65.400 225.500 65.700 226.500 ;
        RECT 61.100 224.600 61.900 224.900 ;
        RECT 63.800 225.200 65.700 225.500 ;
        RECT 59.000 221.500 59.400 223.500 ;
        RECT 61.100 222.200 61.500 224.600 ;
        RECT 63.800 223.500 64.100 225.200 ;
        RECT 66.400 224.900 66.700 226.800 ;
        RECT 68.600 226.500 69.500 226.900 ;
        RECT 69.900 226.500 71.200 226.900 ;
        RECT 71.700 226.500 72.900 226.900 ;
        RECT 73.300 226.500 74.600 226.900 ;
        RECT 67.000 226.100 67.400 226.200 ;
        RECT 67.800 226.100 68.200 226.200 ;
        RECT 67.000 225.800 68.200 226.100 ;
        RECT 69.900 225.800 70.300 226.500 ;
        RECT 71.700 225.800 72.100 226.500 ;
        RECT 73.300 225.800 73.700 226.500 ;
        RECT 75.000 225.800 75.400 227.200 ;
        RECT 67.000 225.400 67.400 225.800 ;
        RECT 69.400 225.400 70.300 225.800 ;
        RECT 71.000 225.400 72.100 225.800 ;
        RECT 72.600 225.400 73.700 225.800 ;
        RECT 74.200 225.400 75.400 225.800 ;
        RECT 75.800 227.400 77.700 227.700 ;
        RECT 75.800 225.700 76.200 227.400 ;
        RECT 79.300 227.100 79.700 227.200 ;
        RECT 82.200 227.100 82.500 228.200 ;
        RECT 84.600 227.500 85.000 229.900 ;
        RECT 86.700 228.200 87.100 229.900 ;
        RECT 86.200 227.900 87.100 228.200 ;
        RECT 87.800 227.900 88.200 229.900 ;
        RECT 88.600 228.000 89.000 229.900 ;
        RECT 90.200 228.000 90.600 229.900 ;
        RECT 92.900 228.000 93.300 229.500 ;
        RECT 95.000 228.500 95.400 229.500 ;
        RECT 88.600 227.900 90.600 228.000 ;
        RECT 83.800 227.100 84.600 227.200 ;
        RECT 79.100 226.800 84.600 227.100 ;
        RECT 85.400 226.800 85.800 227.600 ;
        RECT 78.200 226.400 78.600 226.500 ;
        RECT 76.700 226.100 78.600 226.400 ;
        RECT 79.100 226.200 79.400 226.800 ;
        RECT 82.700 226.700 83.100 226.800 ;
        RECT 82.200 226.200 82.600 226.300 ;
        RECT 83.500 226.200 83.900 226.300 ;
        RECT 76.700 226.000 77.100 226.100 ;
        RECT 79.000 225.800 79.400 226.200 ;
        RECT 81.400 225.900 83.900 226.200 ;
        RECT 81.400 225.800 81.800 225.900 ;
        RECT 77.500 225.700 77.900 225.800 ;
        RECT 75.800 225.400 77.900 225.700 ;
        RECT 65.900 224.600 66.700 224.900 ;
        RECT 61.100 221.800 61.800 222.200 ;
        RECT 61.100 221.100 61.500 221.800 ;
        RECT 63.800 221.500 64.200 223.500 ;
        RECT 65.900 222.200 66.300 224.600 ;
        RECT 65.900 221.800 66.600 222.200 ;
        RECT 65.900 221.100 66.300 221.800 ;
        RECT 69.400 221.100 69.800 225.400 ;
        RECT 71.000 221.100 71.400 225.400 ;
        RECT 72.600 221.100 73.000 225.400 ;
        RECT 74.200 221.100 74.600 225.400 ;
        RECT 75.800 221.100 76.200 225.400 ;
        RECT 79.100 225.200 79.400 225.800 ;
        RECT 82.200 225.500 85.000 225.600 ;
        RECT 82.100 225.400 85.000 225.500 ;
        RECT 78.200 224.900 79.400 225.200 ;
        RECT 80.100 225.300 85.000 225.400 ;
        RECT 80.100 225.100 82.500 225.300 ;
        RECT 78.200 224.400 78.500 224.900 ;
        RECT 77.800 224.000 78.500 224.400 ;
        RECT 79.300 224.500 79.700 224.600 ;
        RECT 80.100 224.500 80.400 225.100 ;
        RECT 79.300 224.200 80.400 224.500 ;
        RECT 80.700 224.500 83.400 224.800 ;
        RECT 80.700 224.400 81.100 224.500 ;
        RECT 83.000 224.400 83.400 224.500 ;
        RECT 79.900 223.700 80.300 223.800 ;
        RECT 81.300 223.700 81.700 223.800 ;
        RECT 78.200 223.100 78.600 223.500 ;
        RECT 79.900 223.400 81.700 223.700 ;
        RECT 80.300 223.100 80.600 223.400 ;
        RECT 83.000 223.100 83.400 223.500 ;
        RECT 77.900 221.100 78.500 223.100 ;
        RECT 80.200 221.100 80.600 223.100 ;
        RECT 82.400 222.800 83.400 223.100 ;
        RECT 82.400 221.100 82.800 222.800 ;
        RECT 84.600 221.100 85.000 225.300 ;
        RECT 85.400 225.100 85.800 225.200 ;
        RECT 86.200 225.100 86.600 227.900 ;
        RECT 87.900 227.200 88.200 227.900 ;
        RECT 88.700 227.700 90.500 227.900 ;
        RECT 92.500 227.700 93.300 228.000 ;
        RECT 92.500 227.500 92.900 227.700 ;
        RECT 89.800 227.200 90.200 227.400 ;
        RECT 92.500 227.200 92.800 227.500 ;
        RECT 95.100 227.400 95.400 228.500 ;
        RECT 87.800 226.800 89.100 227.200 ;
        RECT 89.800 226.900 90.600 227.200 ;
        RECT 90.200 226.800 90.600 226.900 ;
        RECT 91.800 226.800 92.800 227.200 ;
        RECT 93.300 227.100 95.400 227.400 ;
        RECT 97.400 227.700 97.800 229.900 ;
        RECT 99.500 229.200 100.100 229.900 ;
        RECT 99.500 228.900 100.200 229.200 ;
        RECT 101.800 228.900 102.200 229.900 ;
        RECT 104.000 229.200 104.400 229.900 ;
        RECT 104.000 228.900 105.000 229.200 ;
        RECT 99.800 228.500 100.200 228.900 ;
        RECT 101.900 228.600 102.200 228.900 ;
        RECT 101.900 228.300 103.300 228.600 ;
        RECT 102.900 228.200 103.300 228.300 ;
        RECT 103.800 228.200 104.200 228.600 ;
        RECT 104.600 228.500 105.000 228.900 ;
        RECT 100.600 227.800 101.000 228.200 ;
        RECT 98.900 227.700 99.300 227.800 ;
        RECT 97.400 227.400 99.300 227.700 ;
        RECT 93.300 226.900 93.800 227.100 ;
        RECT 87.000 226.100 87.400 226.200 ;
        RECT 88.800 226.100 89.100 226.800 ;
        RECT 87.000 225.800 89.100 226.100 ;
        RECT 89.400 226.100 89.800 226.600 ;
        RECT 91.000 226.100 91.400 226.200 ;
        RECT 89.400 225.800 91.400 226.100 ;
        RECT 85.400 224.800 86.600 225.100 ;
        RECT 86.200 221.100 86.600 224.800 ;
        RECT 87.000 224.400 87.400 225.200 ;
        RECT 87.800 225.100 88.200 225.200 ;
        RECT 88.800 225.100 89.100 225.800 ;
        RECT 91.800 225.400 92.200 226.200 ;
        RECT 87.800 224.800 88.500 225.100 ;
        RECT 88.800 224.800 89.300 225.100 ;
        RECT 88.200 224.200 88.500 224.800 ;
        RECT 88.200 223.800 88.600 224.200 ;
        RECT 88.900 221.100 89.300 224.800 ;
        RECT 92.500 224.900 92.800 226.800 ;
        RECT 93.100 226.500 93.800 226.900 ;
        RECT 93.500 225.500 93.800 226.500 ;
        RECT 94.200 225.800 94.600 226.600 ;
        RECT 95.000 225.800 95.400 226.600 ;
        RECT 97.400 225.700 97.800 227.400 ;
        RECT 100.600 227.200 100.900 227.800 ;
        RECT 103.800 227.200 104.100 228.200 ;
        RECT 106.200 227.500 106.600 229.900 ;
        RECT 107.000 228.000 107.400 229.900 ;
        RECT 108.600 228.000 109.000 229.900 ;
        RECT 107.000 227.900 109.000 228.000 ;
        RECT 109.400 227.900 109.800 229.900 ;
        RECT 111.500 228.200 111.900 229.900 ;
        RECT 111.000 227.900 111.900 228.200 ;
        RECT 112.600 227.900 113.000 229.900 ;
        RECT 113.400 228.000 113.800 229.900 ;
        RECT 115.000 228.000 115.400 229.900 ;
        RECT 116.600 228.900 117.000 229.900 ;
        RECT 113.400 227.900 115.400 228.000 ;
        RECT 107.100 227.700 108.900 227.900 ;
        RECT 107.400 227.200 107.800 227.400 ;
        RECT 109.400 227.200 109.700 227.900 ;
        RECT 100.600 227.100 101.300 227.200 ;
        RECT 103.800 227.100 104.200 227.200 ;
        RECT 105.400 227.100 106.200 227.200 ;
        RECT 100.600 226.800 106.200 227.100 ;
        RECT 107.000 226.900 107.800 227.200 ;
        RECT 107.000 226.800 107.400 226.900 ;
        RECT 108.500 226.800 109.800 227.200 ;
        RECT 110.200 226.800 110.600 227.600 ;
        RECT 99.800 226.400 100.200 226.500 ;
        RECT 98.300 226.100 100.200 226.400 ;
        RECT 98.300 226.000 98.700 226.100 ;
        RECT 99.100 225.700 99.500 225.800 ;
        RECT 93.500 225.200 95.400 225.500 ;
        RECT 92.500 224.600 93.300 224.900 ;
        RECT 92.900 222.200 93.300 224.600 ;
        RECT 95.100 223.500 95.400 225.200 ;
        RECT 92.900 221.800 93.800 222.200 ;
        RECT 92.900 221.100 93.300 221.800 ;
        RECT 95.000 221.500 95.400 223.500 ;
        RECT 97.400 225.400 99.500 225.700 ;
        RECT 97.400 221.100 97.800 225.400 ;
        RECT 100.700 225.200 101.000 226.800 ;
        RECT 104.300 226.700 104.700 226.800 ;
        RECT 105.100 226.200 105.500 226.300 ;
        RECT 103.000 225.900 105.500 226.200 ;
        RECT 103.000 225.800 103.400 225.900 ;
        RECT 107.800 225.800 108.200 226.600 ;
        RECT 108.500 226.100 108.800 226.800 ;
        RECT 109.400 226.100 109.800 226.200 ;
        RECT 108.500 225.800 109.800 226.100 ;
        RECT 103.800 225.500 106.600 225.600 ;
        RECT 103.700 225.400 106.600 225.500 ;
        RECT 99.800 224.900 101.000 225.200 ;
        RECT 101.700 225.300 106.600 225.400 ;
        RECT 101.700 225.100 104.100 225.300 ;
        RECT 99.800 224.400 100.100 224.900 ;
        RECT 99.400 224.000 100.100 224.400 ;
        RECT 100.900 224.500 101.300 224.600 ;
        RECT 101.700 224.500 102.000 225.100 ;
        RECT 100.900 224.200 102.000 224.500 ;
        RECT 102.300 224.500 105.000 224.800 ;
        RECT 102.300 224.400 102.700 224.500 ;
        RECT 104.600 224.400 105.000 224.500 ;
        RECT 101.500 223.700 101.900 223.800 ;
        RECT 102.900 223.700 103.300 223.800 ;
        RECT 99.800 223.100 100.200 223.500 ;
        RECT 101.500 223.400 103.300 223.700 ;
        RECT 101.900 223.100 102.200 223.400 ;
        RECT 104.600 223.100 105.000 223.500 ;
        RECT 99.500 221.100 100.100 223.100 ;
        RECT 101.800 221.100 102.200 223.100 ;
        RECT 104.000 222.800 105.000 223.100 ;
        RECT 104.000 221.100 104.400 222.800 ;
        RECT 106.200 221.100 106.600 225.300 ;
        RECT 108.500 225.100 108.800 225.800 ;
        RECT 109.400 225.100 109.800 225.200 ;
        RECT 111.000 225.100 111.400 227.900 ;
        RECT 112.700 227.200 113.000 227.900 ;
        RECT 113.500 227.700 115.300 227.900 ;
        RECT 115.800 227.800 116.200 228.600 ;
        RECT 116.700 228.100 117.000 228.900 ;
        RECT 118.300 228.200 118.700 228.600 ;
        RECT 118.200 228.100 118.600 228.200 ;
        RECT 116.600 227.800 118.600 228.100 ;
        RECT 119.000 227.900 119.400 229.900 ;
        RECT 121.700 229.200 122.100 229.900 ;
        RECT 121.400 228.800 122.100 229.200 ;
        RECT 121.700 228.200 122.100 228.800 ;
        RECT 121.700 227.900 122.600 228.200 ;
        RECT 125.700 228.000 126.100 229.500 ;
        RECT 127.800 228.500 128.200 229.500 ;
        RECT 114.600 227.200 115.000 227.400 ;
        RECT 116.700 227.200 117.000 227.800 ;
        RECT 112.600 226.800 113.900 227.200 ;
        RECT 114.600 226.900 115.400 227.200 ;
        RECT 115.000 226.800 115.400 226.900 ;
        RECT 116.600 226.800 117.000 227.200 ;
        RECT 108.300 224.800 108.800 225.100 ;
        RECT 109.100 224.800 111.400 225.100 ;
        RECT 108.300 221.100 108.700 224.800 ;
        RECT 109.100 224.200 109.400 224.800 ;
        RECT 109.000 223.800 109.400 224.200 ;
        RECT 111.000 221.100 111.400 224.800 ;
        RECT 111.800 224.400 112.200 225.200 ;
        RECT 112.600 225.100 113.000 225.200 ;
        RECT 113.600 225.100 113.900 226.800 ;
        RECT 114.200 226.100 114.600 226.600 ;
        RECT 115.000 226.100 115.400 226.200 ;
        RECT 114.200 225.800 115.400 226.100 ;
        RECT 116.700 225.100 117.000 226.800 ;
        RECT 117.400 225.400 117.800 226.200 ;
        RECT 118.200 226.100 118.600 226.200 ;
        RECT 119.100 226.100 119.400 227.900 ;
        RECT 119.800 226.400 120.200 227.200 ;
        RECT 120.600 226.100 121.000 226.200 ;
        RECT 118.200 225.800 119.400 226.100 ;
        RECT 120.200 225.800 121.000 226.100 ;
        RECT 118.300 225.100 118.600 225.800 ;
        RECT 120.200 225.600 120.600 225.800 ;
        RECT 112.600 224.800 113.300 225.100 ;
        RECT 113.600 224.800 114.100 225.100 ;
        RECT 113.000 224.200 113.300 224.800 ;
        RECT 113.000 223.800 113.400 224.200 ;
        RECT 113.700 222.200 114.100 224.800 ;
        RECT 116.600 224.700 117.500 225.100 ;
        RECT 113.700 221.800 114.600 222.200 ;
        RECT 113.700 221.100 114.100 221.800 ;
        RECT 117.100 221.100 117.500 224.700 ;
        RECT 118.200 221.100 118.600 225.100 ;
        RECT 119.000 224.800 121.000 225.100 ;
        RECT 119.000 221.100 119.400 224.800 ;
        RECT 120.600 221.100 121.000 224.800 ;
        RECT 121.400 224.400 121.800 225.200 ;
        RECT 122.200 221.100 122.600 227.900 ;
        RECT 125.300 227.700 126.100 228.000 ;
        RECT 123.000 226.800 123.400 227.600 ;
        RECT 125.300 227.500 125.700 227.700 ;
        RECT 125.300 227.200 125.600 227.500 ;
        RECT 127.900 227.400 128.200 228.500 ;
        RECT 123.800 227.100 124.200 227.200 ;
        RECT 124.600 227.100 125.600 227.200 ;
        RECT 123.800 226.800 125.600 227.100 ;
        RECT 126.100 227.100 128.200 227.400 ;
        RECT 128.600 227.700 129.000 229.900 ;
        RECT 130.700 229.200 131.300 229.900 ;
        RECT 130.700 228.900 131.400 229.200 ;
        RECT 133.000 228.900 133.400 229.900 ;
        RECT 135.200 229.200 135.600 229.900 ;
        RECT 135.200 228.900 136.200 229.200 ;
        RECT 131.000 228.500 131.400 228.900 ;
        RECT 133.100 228.600 133.400 228.900 ;
        RECT 133.100 228.300 134.500 228.600 ;
        RECT 134.100 228.200 134.500 228.300 ;
        RECT 135.000 228.200 135.400 228.600 ;
        RECT 135.800 228.500 136.200 228.900 ;
        RECT 130.100 227.700 130.500 227.800 ;
        RECT 128.600 227.400 130.500 227.700 ;
        RECT 126.100 226.900 126.600 227.100 ;
        RECT 123.000 226.100 123.300 226.800 ;
        RECT 124.600 226.100 125.000 226.200 ;
        RECT 123.000 225.800 125.000 226.100 ;
        RECT 124.600 225.400 125.000 225.800 ;
        RECT 125.300 224.900 125.600 226.800 ;
        RECT 125.900 226.500 126.600 226.900 ;
        RECT 126.300 225.500 126.600 226.500 ;
        RECT 127.000 225.800 127.400 226.600 ;
        RECT 127.800 225.800 128.200 226.600 ;
        RECT 128.600 225.700 129.000 227.400 ;
        RECT 132.100 227.100 132.500 227.200 ;
        RECT 135.000 227.100 135.300 228.200 ;
        RECT 137.400 227.500 137.800 229.900 ;
        RECT 138.200 228.000 138.600 229.900 ;
        RECT 139.800 228.000 140.200 229.900 ;
        RECT 138.200 227.900 140.200 228.000 ;
        RECT 140.600 227.900 141.000 229.900 ;
        RECT 142.700 228.200 143.100 229.900 ;
        RECT 142.200 227.900 143.100 228.200 ;
        RECT 145.700 228.000 146.100 229.500 ;
        RECT 147.800 228.500 148.200 229.500 ;
        RECT 138.300 227.700 140.100 227.900 ;
        RECT 138.600 227.200 139.000 227.400 ;
        RECT 140.600 227.200 140.900 227.900 ;
        RECT 136.600 227.100 137.400 227.200 ;
        RECT 131.900 226.800 137.400 227.100 ;
        RECT 138.200 226.900 139.000 227.200 ;
        RECT 138.200 226.800 138.600 226.900 ;
        RECT 139.700 226.800 141.000 227.200 ;
        RECT 141.400 226.800 141.800 227.600 ;
        RECT 131.000 226.400 131.400 226.500 ;
        RECT 129.500 226.100 131.400 226.400 ;
        RECT 129.500 226.000 129.900 226.100 ;
        RECT 130.300 225.700 130.700 225.800 ;
        RECT 126.300 225.200 128.200 225.500 ;
        RECT 125.300 224.600 126.100 224.900 ;
        RECT 125.700 221.100 126.100 224.600 ;
        RECT 127.900 223.500 128.200 225.200 ;
        RECT 127.800 221.500 128.200 223.500 ;
        RECT 128.600 225.400 130.700 225.700 ;
        RECT 128.600 221.100 129.000 225.400 ;
        RECT 131.900 225.200 132.200 226.800 ;
        RECT 135.500 226.700 135.900 226.800 ;
        RECT 135.000 226.200 135.400 226.300 ;
        RECT 136.300 226.200 136.700 226.300 ;
        RECT 134.200 225.900 136.700 226.200 ;
        RECT 134.200 225.800 134.600 225.900 ;
        RECT 139.000 225.800 139.400 226.600 ;
        RECT 135.000 225.500 137.800 225.600 ;
        RECT 134.900 225.400 137.800 225.500 ;
        RECT 131.000 224.900 132.200 225.200 ;
        RECT 132.900 225.300 137.800 225.400 ;
        RECT 132.900 225.100 135.300 225.300 ;
        RECT 131.000 224.400 131.300 224.900 ;
        RECT 130.600 224.000 131.300 224.400 ;
        RECT 132.100 224.500 132.500 224.600 ;
        RECT 132.900 224.500 133.200 225.100 ;
        RECT 132.100 224.200 133.200 224.500 ;
        RECT 133.500 224.500 136.200 224.800 ;
        RECT 133.500 224.400 133.900 224.500 ;
        RECT 135.800 224.400 136.200 224.500 ;
        RECT 132.700 223.700 133.100 223.800 ;
        RECT 134.100 223.700 134.500 223.800 ;
        RECT 131.000 223.100 131.400 223.500 ;
        RECT 132.700 223.400 134.500 223.700 ;
        RECT 133.100 223.100 133.400 223.400 ;
        RECT 135.800 223.100 136.200 223.500 ;
        RECT 130.700 221.100 131.300 223.100 ;
        RECT 133.000 221.100 133.400 223.100 ;
        RECT 135.200 222.800 136.200 223.100 ;
        RECT 135.200 221.100 135.600 222.800 ;
        RECT 137.400 221.100 137.800 225.300 ;
        RECT 139.700 225.200 140.000 226.800 ;
        RECT 139.000 224.800 140.000 225.200 ;
        RECT 140.600 225.100 141.000 225.200 ;
        RECT 142.200 225.100 142.600 227.900 ;
        RECT 145.300 227.700 146.100 228.000 ;
        RECT 145.300 227.500 145.700 227.700 ;
        RECT 145.300 227.200 145.600 227.500 ;
        RECT 147.900 227.400 148.200 228.500 ;
        RECT 144.600 226.800 145.600 227.200 ;
        RECT 146.100 227.100 148.200 227.400 ;
        RECT 150.200 227.700 150.600 229.900 ;
        RECT 152.300 229.200 152.900 229.900 ;
        RECT 152.300 228.900 153.000 229.200 ;
        RECT 154.600 228.900 155.000 229.900 ;
        RECT 156.800 229.200 157.200 229.900 ;
        RECT 156.800 228.900 157.800 229.200 ;
        RECT 152.600 228.500 153.000 228.900 ;
        RECT 154.700 228.600 155.000 228.900 ;
        RECT 154.700 228.300 156.100 228.600 ;
        RECT 155.700 228.200 156.100 228.300 ;
        RECT 156.600 228.200 157.000 228.600 ;
        RECT 157.400 228.500 157.800 228.900 ;
        RECT 151.700 227.700 152.100 227.800 ;
        RECT 150.200 227.400 152.100 227.700 ;
        RECT 146.100 226.900 146.600 227.100 ;
        RECT 144.600 225.400 145.000 226.200 ;
        RECT 140.300 224.800 142.600 225.100 ;
        RECT 139.500 221.100 139.900 224.800 ;
        RECT 140.300 224.200 140.600 224.800 ;
        RECT 140.200 223.800 140.600 224.200 ;
        RECT 142.200 221.100 142.600 224.800 ;
        RECT 143.000 224.400 143.400 225.200 ;
        RECT 145.300 224.900 145.600 226.800 ;
        RECT 145.900 226.500 146.600 226.900 ;
        RECT 146.300 225.500 146.600 226.500 ;
        RECT 147.000 225.800 147.400 226.600 ;
        RECT 147.800 226.100 148.200 226.600 ;
        RECT 148.600 226.100 149.000 226.200 ;
        RECT 147.800 225.800 149.000 226.100 ;
        RECT 150.200 225.700 150.600 227.400 ;
        RECT 153.700 227.100 154.100 227.200 ;
        RECT 156.600 227.100 156.900 228.200 ;
        RECT 159.000 227.500 159.400 229.900 ;
        RECT 161.400 227.800 161.800 229.900 ;
        RECT 163.800 228.900 164.200 229.900 ;
        RECT 162.100 228.200 162.500 228.600 ;
        RECT 162.200 228.100 162.600 228.200 ;
        RECT 163.800 228.100 164.100 228.900 ;
        RECT 162.200 227.800 164.100 228.100 ;
        RECT 164.600 227.800 165.000 228.600 ;
        RECT 158.200 227.100 159.000 227.200 ;
        RECT 153.500 226.800 159.000 227.100 ;
        RECT 152.600 226.400 153.000 226.500 ;
        RECT 151.100 226.100 153.000 226.400 ;
        RECT 151.100 226.000 151.500 226.100 ;
        RECT 151.900 225.700 152.300 225.800 ;
        RECT 146.300 225.200 148.200 225.500 ;
        RECT 145.300 224.600 146.100 224.900 ;
        RECT 145.700 222.200 146.100 224.600 ;
        RECT 147.900 223.500 148.200 225.200 ;
        RECT 145.400 221.800 146.100 222.200 ;
        RECT 145.700 221.100 146.100 221.800 ;
        RECT 147.800 221.500 148.200 223.500 ;
        RECT 150.200 225.400 152.300 225.700 ;
        RECT 150.200 221.100 150.600 225.400 ;
        RECT 153.500 225.200 153.800 226.800 ;
        RECT 157.100 226.700 157.500 226.800 ;
        RECT 160.600 226.400 161.000 227.200 ;
        RECT 157.900 226.200 158.300 226.300 ;
        RECT 155.000 226.100 155.400 226.200 ;
        RECT 155.800 226.100 158.300 226.200 ;
        RECT 155.000 225.900 158.300 226.100 ;
        RECT 159.800 226.100 160.200 226.200 ;
        RECT 161.400 226.100 161.700 227.800 ;
        RECT 163.800 227.200 164.100 227.800 ;
        RECT 166.200 227.600 166.600 229.900 ;
        RECT 167.800 227.600 168.200 229.900 ;
        RECT 169.400 227.600 169.800 229.900 ;
        RECT 171.000 227.600 171.400 229.900 ;
        RECT 165.400 227.200 166.600 227.600 ;
        RECT 167.100 227.200 168.200 227.600 ;
        RECT 168.700 227.200 169.800 227.600 ;
        RECT 170.500 227.200 171.400 227.600 ;
        RECT 172.600 227.500 173.000 229.900 ;
        RECT 174.800 229.200 175.200 229.900 ;
        RECT 174.200 228.900 175.200 229.200 ;
        RECT 177.000 228.900 177.400 229.900 ;
        RECT 179.100 229.200 179.700 229.900 ;
        RECT 179.000 228.900 179.700 229.200 ;
        RECT 174.200 228.500 174.600 228.900 ;
        RECT 177.000 228.600 177.300 228.900 ;
        RECT 175.000 228.200 175.400 228.600 ;
        RECT 175.900 228.300 177.300 228.600 ;
        RECT 179.000 228.500 179.400 228.900 ;
        RECT 175.900 228.200 176.300 228.300 ;
        RECT 163.800 226.800 164.200 227.200 ;
        RECT 162.200 226.100 162.600 226.200 ;
        RECT 155.000 225.800 156.200 225.900 ;
        RECT 159.800 225.800 160.600 226.100 ;
        RECT 161.400 225.800 162.600 226.100 ;
        RECT 160.200 225.600 160.600 225.800 ;
        RECT 156.600 225.500 159.400 225.600 ;
        RECT 156.500 225.400 159.400 225.500 ;
        RECT 152.600 224.900 153.800 225.200 ;
        RECT 154.500 225.300 159.400 225.400 ;
        RECT 154.500 225.100 156.900 225.300 ;
        RECT 152.600 224.400 152.900 224.900 ;
        RECT 152.200 224.000 152.900 224.400 ;
        RECT 153.700 224.500 154.100 224.600 ;
        RECT 154.500 224.500 154.800 225.100 ;
        RECT 153.700 224.200 154.800 224.500 ;
        RECT 155.100 224.500 157.800 224.800 ;
        RECT 155.100 224.400 155.500 224.500 ;
        RECT 157.400 224.400 157.800 224.500 ;
        RECT 154.300 223.700 154.700 223.800 ;
        RECT 155.700 223.700 156.100 223.800 ;
        RECT 152.600 223.100 153.000 223.500 ;
        RECT 154.300 223.400 156.100 223.700 ;
        RECT 154.700 223.100 155.000 223.400 ;
        RECT 157.400 223.100 157.800 223.500 ;
        RECT 152.300 221.100 152.900 223.100 ;
        RECT 154.600 221.100 155.000 223.100 ;
        RECT 156.800 222.800 157.800 223.100 ;
        RECT 156.800 221.100 157.200 222.800 ;
        RECT 159.000 221.100 159.400 225.300 ;
        RECT 162.200 225.100 162.500 225.800 ;
        RECT 163.000 225.400 163.400 226.200 ;
        RECT 163.800 225.100 164.100 226.800 ;
        RECT 165.400 225.800 165.800 227.200 ;
        RECT 167.100 226.900 167.500 227.200 ;
        RECT 168.700 226.900 169.100 227.200 ;
        RECT 170.500 226.900 170.900 227.200 ;
        RECT 171.800 227.100 172.200 227.200 ;
        RECT 173.000 227.100 173.800 227.200 ;
        RECT 175.100 227.100 175.400 228.200 ;
        RECT 179.900 227.700 180.300 227.800 ;
        RECT 181.400 227.700 181.800 229.900 ;
        RECT 179.900 227.400 181.800 227.700 ;
        RECT 175.800 227.100 176.200 227.200 ;
        RECT 177.900 227.100 178.300 227.200 ;
        RECT 171.800 226.900 178.500 227.100 ;
        RECT 166.200 226.500 167.500 226.900 ;
        RECT 167.900 226.500 169.100 226.900 ;
        RECT 169.600 226.500 170.900 226.900 ;
        RECT 171.300 226.800 178.500 226.900 ;
        RECT 171.300 226.500 172.200 226.800 ;
        RECT 174.500 226.700 174.900 226.800 ;
        RECT 167.100 225.800 167.500 226.500 ;
        RECT 168.700 225.800 169.100 226.500 ;
        RECT 170.500 225.800 170.900 226.500 ;
        RECT 173.700 226.200 174.100 226.300 ;
        RECT 175.000 226.200 175.400 226.300 ;
        RECT 173.700 225.900 176.200 226.200 ;
        RECT 175.800 225.800 176.200 225.900 ;
        RECT 165.400 225.400 166.600 225.800 ;
        RECT 167.100 225.400 168.200 225.800 ;
        RECT 168.700 225.400 169.800 225.800 ;
        RECT 170.500 225.400 171.400 225.800 ;
        RECT 159.800 224.800 161.800 225.100 ;
        RECT 159.800 221.100 160.200 224.800 ;
        RECT 161.400 221.100 161.800 224.800 ;
        RECT 162.200 221.100 162.600 225.100 ;
        RECT 163.300 224.700 164.200 225.100 ;
        RECT 163.300 221.100 163.700 224.700 ;
        RECT 166.200 221.100 166.600 225.400 ;
        RECT 167.800 221.100 168.200 225.400 ;
        RECT 169.400 221.100 169.800 225.400 ;
        RECT 171.000 221.100 171.400 225.400 ;
        RECT 172.600 225.500 175.400 225.600 ;
        RECT 172.600 225.400 175.500 225.500 ;
        RECT 172.600 225.300 177.500 225.400 ;
        RECT 172.600 221.100 173.000 225.300 ;
        RECT 175.100 225.100 177.500 225.300 ;
        RECT 174.200 224.500 176.900 224.800 ;
        RECT 174.200 224.400 174.600 224.500 ;
        RECT 176.500 224.400 176.900 224.500 ;
        RECT 177.200 224.500 177.500 225.100 ;
        RECT 178.200 225.200 178.500 226.800 ;
        RECT 179.000 226.400 179.400 226.500 ;
        RECT 179.000 226.100 180.900 226.400 ;
        RECT 180.500 226.000 180.900 226.100 ;
        RECT 179.700 225.700 180.100 225.800 ;
        RECT 181.400 225.700 181.800 227.400 ;
        RECT 182.200 228.500 182.600 229.500 ;
        RECT 182.200 227.400 182.500 228.500 ;
        RECT 184.300 228.000 184.700 229.500 ;
        RECT 188.900 228.200 189.300 229.500 ;
        RECT 191.000 228.500 191.400 229.500 ;
        RECT 188.900 228.000 189.800 228.200 ;
        RECT 184.300 227.700 185.100 228.000 ;
        RECT 184.700 227.500 185.100 227.700 ;
        RECT 182.200 227.100 184.300 227.400 ;
        RECT 183.800 226.900 184.300 227.100 ;
        RECT 184.800 227.200 185.100 227.500 ;
        RECT 188.500 227.800 189.800 228.000 ;
        RECT 188.500 227.700 189.300 227.800 ;
        RECT 188.500 227.500 188.900 227.700 ;
        RECT 188.500 227.200 188.800 227.500 ;
        RECT 191.100 227.400 191.400 228.500 ;
        RECT 182.200 225.800 182.600 226.600 ;
        RECT 183.000 225.800 183.400 226.600 ;
        RECT 183.800 226.500 184.500 226.900 ;
        RECT 184.800 226.800 185.800 227.200 ;
        RECT 187.800 226.800 188.800 227.200 ;
        RECT 189.300 227.100 191.400 227.400 ;
        RECT 191.800 228.500 192.200 229.500 ;
        RECT 191.800 227.400 192.100 228.500 ;
        RECT 193.900 228.000 194.300 229.500 ;
        RECT 196.600 228.000 197.000 229.900 ;
        RECT 198.200 228.000 198.600 229.900 ;
        RECT 193.900 227.700 194.700 228.000 ;
        RECT 196.600 227.900 198.600 228.000 ;
        RECT 199.000 227.900 199.400 229.900 ;
        RECT 200.100 228.200 200.500 229.900 ;
        RECT 205.100 229.200 205.500 229.900 ;
        RECT 204.600 228.800 205.500 229.200 ;
        RECT 205.100 228.200 205.500 228.800 ;
        RECT 200.100 227.900 201.000 228.200 ;
        RECT 196.700 227.700 198.500 227.900 ;
        RECT 194.300 227.500 194.700 227.700 ;
        RECT 191.800 227.100 193.900 227.400 ;
        RECT 189.300 226.900 189.800 227.100 ;
        RECT 179.700 225.400 181.800 225.700 ;
        RECT 183.800 225.500 184.100 226.500 ;
        RECT 178.200 224.900 179.400 225.200 ;
        RECT 177.900 224.500 178.300 224.600 ;
        RECT 177.200 224.200 178.300 224.500 ;
        RECT 179.100 224.400 179.400 224.900 ;
        RECT 179.100 224.000 179.800 224.400 ;
        RECT 175.900 223.700 176.300 223.800 ;
        RECT 177.300 223.700 177.700 223.800 ;
        RECT 174.200 223.100 174.600 223.500 ;
        RECT 175.900 223.400 177.700 223.700 ;
        RECT 177.000 223.100 177.300 223.400 ;
        RECT 179.000 223.100 179.400 223.500 ;
        RECT 174.200 222.800 175.200 223.100 ;
        RECT 174.800 221.100 175.200 222.800 ;
        RECT 177.000 221.100 177.400 223.100 ;
        RECT 179.100 221.100 179.700 223.100 ;
        RECT 181.400 221.100 181.800 225.400 ;
        RECT 182.200 225.200 184.100 225.500 ;
        RECT 182.200 223.500 182.500 225.200 ;
        RECT 184.800 224.900 185.100 226.800 ;
        RECT 185.400 226.100 185.800 226.200 ;
        RECT 186.200 226.100 186.600 226.200 ;
        RECT 185.400 225.800 186.600 226.100 ;
        RECT 185.400 225.400 185.800 225.800 ;
        RECT 187.800 225.400 188.200 226.200 ;
        RECT 184.300 224.600 185.100 224.900 ;
        RECT 188.500 224.900 188.800 226.800 ;
        RECT 189.100 226.500 189.800 226.900 ;
        RECT 193.400 226.900 193.900 227.100 ;
        RECT 194.400 227.200 194.700 227.500 ;
        RECT 197.000 227.200 197.400 227.400 ;
        RECT 199.000 227.200 199.300 227.900 ;
        RECT 189.500 225.500 189.800 226.500 ;
        RECT 190.200 225.800 190.600 226.600 ;
        RECT 191.000 225.800 191.400 226.600 ;
        RECT 191.800 225.800 192.200 226.600 ;
        RECT 192.600 225.800 193.000 226.600 ;
        RECT 193.400 226.500 194.100 226.900 ;
        RECT 194.400 226.800 195.400 227.200 ;
        RECT 195.800 227.100 196.200 227.200 ;
        RECT 196.600 227.100 197.400 227.200 ;
        RECT 195.800 226.900 197.400 227.100 ;
        RECT 195.800 226.800 197.000 226.900 ;
        RECT 198.100 226.800 199.400 227.200 ;
        RECT 193.400 225.500 193.700 226.500 ;
        RECT 189.500 225.200 191.400 225.500 ;
        RECT 188.500 224.600 189.300 224.900 ;
        RECT 182.200 221.500 182.600 223.500 ;
        RECT 184.300 222.200 184.700 224.600 ;
        RECT 184.300 221.800 185.000 222.200 ;
        RECT 184.300 221.100 184.700 221.800 ;
        RECT 188.900 221.100 189.300 224.600 ;
        RECT 191.100 223.500 191.400 225.200 ;
        RECT 191.000 221.500 191.400 223.500 ;
        RECT 191.800 225.200 193.700 225.500 ;
        RECT 191.800 223.500 192.100 225.200 ;
        RECT 194.400 224.900 194.700 226.800 ;
        RECT 195.000 225.400 195.400 226.200 ;
        RECT 197.400 225.800 197.800 226.600 ;
        RECT 198.100 225.100 198.400 226.800 ;
        RECT 200.600 226.100 201.000 227.900 ;
        RECT 204.600 227.900 205.500 228.200 ;
        RECT 201.400 226.800 201.800 227.600 ;
        RECT 203.800 226.800 204.200 227.600 ;
        RECT 199.000 225.800 201.000 226.100 ;
        RECT 199.000 225.200 199.300 225.800 ;
        RECT 199.000 225.100 199.400 225.200 ;
        RECT 193.900 224.600 194.700 224.900 ;
        RECT 197.900 224.800 198.400 225.100 ;
        RECT 198.700 224.800 199.400 225.100 ;
        RECT 191.800 221.500 192.200 223.500 ;
        RECT 193.900 222.200 194.300 224.600 ;
        RECT 193.400 221.800 194.300 222.200 ;
        RECT 193.900 221.100 194.300 221.800 ;
        RECT 197.900 221.100 198.300 224.800 ;
        RECT 198.700 224.200 199.000 224.800 ;
        RECT 199.800 224.400 200.200 225.200 ;
        RECT 198.600 223.800 199.000 224.200 ;
        RECT 200.600 221.100 201.000 225.800 ;
        RECT 204.600 221.100 205.000 227.900 ;
        RECT 206.200 227.500 206.600 229.900 ;
        RECT 208.400 229.200 208.800 229.900 ;
        RECT 207.800 228.900 208.800 229.200 ;
        RECT 210.600 228.900 211.000 229.900 ;
        RECT 212.700 229.200 213.300 229.900 ;
        RECT 212.600 228.900 213.300 229.200 ;
        RECT 207.800 228.500 208.200 228.900 ;
        RECT 210.600 228.600 210.900 228.900 ;
        RECT 208.600 228.200 209.000 228.600 ;
        RECT 209.500 228.300 210.900 228.600 ;
        RECT 212.600 228.500 213.000 228.900 ;
        RECT 209.500 228.200 209.900 228.300 ;
        RECT 206.600 227.100 207.400 227.200 ;
        RECT 208.700 227.100 209.000 228.200 ;
        RECT 213.500 227.700 213.900 227.800 ;
        RECT 215.000 227.700 215.400 229.900 ;
        RECT 213.500 227.400 215.400 227.700 ;
        RECT 210.200 227.100 210.600 227.200 ;
        RECT 211.500 227.100 211.900 227.200 ;
        RECT 206.600 226.800 212.100 227.100 ;
        RECT 208.100 226.700 208.500 226.800 ;
        RECT 207.300 226.200 207.700 226.300 ;
        RECT 208.600 226.200 209.000 226.300 ;
        RECT 207.300 225.900 209.800 226.200 ;
        RECT 209.400 225.800 209.800 225.900 ;
        RECT 206.200 225.500 209.000 225.600 ;
        RECT 206.200 225.400 209.100 225.500 ;
        RECT 206.200 225.300 211.100 225.400 ;
        RECT 205.400 224.400 205.800 225.200 ;
        RECT 206.200 221.100 206.600 225.300 ;
        RECT 208.700 225.100 211.100 225.300 ;
        RECT 207.800 224.500 210.500 224.800 ;
        RECT 207.800 224.400 208.200 224.500 ;
        RECT 210.100 224.400 210.500 224.500 ;
        RECT 210.800 224.500 211.100 225.100 ;
        RECT 211.800 225.200 212.100 226.800 ;
        RECT 212.600 226.400 213.000 226.500 ;
        RECT 212.600 226.100 214.500 226.400 ;
        RECT 214.100 226.000 214.500 226.100 ;
        RECT 213.300 225.700 213.700 225.800 ;
        RECT 215.000 225.700 215.400 227.400 ;
        RECT 215.800 228.500 216.200 229.500 ;
        RECT 215.800 227.400 216.100 228.500 ;
        RECT 217.900 228.000 218.300 229.500 ;
        RECT 222.500 228.000 222.900 229.500 ;
        RECT 224.600 228.500 225.000 229.500 ;
        RECT 217.900 227.700 218.700 228.000 ;
        RECT 218.300 227.500 218.700 227.700 ;
        RECT 215.800 227.100 217.900 227.400 ;
        RECT 217.400 226.900 217.900 227.100 ;
        RECT 218.400 227.200 218.700 227.500 ;
        RECT 222.100 227.700 222.900 228.000 ;
        RECT 222.100 227.500 222.500 227.700 ;
        RECT 222.100 227.200 222.400 227.500 ;
        RECT 224.700 227.400 225.000 228.500 ;
        RECT 225.400 228.000 225.800 229.900 ;
        RECT 227.000 228.000 227.400 229.900 ;
        RECT 225.400 227.900 227.400 228.000 ;
        RECT 227.800 227.900 228.200 229.900 ;
        RECT 228.900 228.200 229.300 229.900 ;
        RECT 228.900 227.900 229.800 228.200 ;
        RECT 225.500 227.700 227.300 227.900 ;
        RECT 215.800 225.800 216.200 226.600 ;
        RECT 216.600 225.800 217.000 226.600 ;
        RECT 217.400 226.500 218.100 226.900 ;
        RECT 218.400 226.800 219.400 227.200 ;
        RECT 221.400 226.800 222.400 227.200 ;
        RECT 222.900 227.100 225.000 227.400 ;
        RECT 225.800 227.200 226.200 227.400 ;
        RECT 227.800 227.200 228.100 227.900 ;
        RECT 222.900 226.900 223.400 227.100 ;
        RECT 213.300 225.400 215.400 225.700 ;
        RECT 217.400 225.500 217.700 226.500 ;
        RECT 211.800 224.900 213.000 225.200 ;
        RECT 211.500 224.500 211.900 224.600 ;
        RECT 210.800 224.200 211.900 224.500 ;
        RECT 212.700 224.400 213.000 224.900 ;
        RECT 212.700 224.000 213.400 224.400 ;
        RECT 209.500 223.700 209.900 223.800 ;
        RECT 210.900 223.700 211.300 223.800 ;
        RECT 207.800 223.100 208.200 223.500 ;
        RECT 209.500 223.400 211.300 223.700 ;
        RECT 210.600 223.100 210.900 223.400 ;
        RECT 212.600 223.100 213.000 223.500 ;
        RECT 207.800 222.800 208.800 223.100 ;
        RECT 208.400 221.100 208.800 222.800 ;
        RECT 210.600 221.100 211.000 223.100 ;
        RECT 212.700 221.100 213.300 223.100 ;
        RECT 215.000 221.100 215.400 225.400 ;
        RECT 215.800 225.200 217.700 225.500 ;
        RECT 215.800 223.500 216.100 225.200 ;
        RECT 218.400 224.900 218.700 226.800 ;
        RECT 219.000 225.400 219.400 226.200 ;
        RECT 220.600 226.100 221.000 226.200 ;
        RECT 221.400 226.100 221.800 226.200 ;
        RECT 220.600 225.800 221.800 226.100 ;
        RECT 221.400 225.400 221.800 225.800 ;
        RECT 217.900 224.600 218.700 224.900 ;
        RECT 222.100 224.900 222.400 226.800 ;
        RECT 222.700 226.500 223.400 226.900 ;
        RECT 225.400 226.900 226.200 227.200 ;
        RECT 226.900 227.100 228.200 227.200 ;
        RECT 228.600 227.100 229.000 227.200 ;
        RECT 225.400 226.800 225.800 226.900 ;
        RECT 226.900 226.800 229.000 227.100 ;
        RECT 223.100 225.500 223.400 226.500 ;
        RECT 223.800 225.800 224.200 226.600 ;
        RECT 224.600 225.800 225.000 226.600 ;
        RECT 226.200 225.800 226.600 226.600 ;
        RECT 223.100 225.200 225.000 225.500 ;
        RECT 222.100 224.600 222.900 224.900 ;
        RECT 215.800 221.500 216.200 223.500 ;
        RECT 217.900 222.200 218.300 224.600 ;
        RECT 217.900 221.800 218.600 222.200 ;
        RECT 217.900 221.100 218.300 221.800 ;
        RECT 222.500 221.100 222.900 224.600 ;
        RECT 224.700 223.500 225.000 225.200 ;
        RECT 226.900 225.100 227.200 226.800 ;
        RECT 229.400 226.100 229.800 227.900 ;
        RECT 231.000 227.700 231.400 229.900 ;
        RECT 233.100 229.200 233.700 229.900 ;
        RECT 233.100 228.900 233.800 229.200 ;
        RECT 235.400 228.900 235.800 229.900 ;
        RECT 237.600 229.200 238.000 229.900 ;
        RECT 237.600 228.900 238.600 229.200 ;
        RECT 233.400 228.500 233.800 228.900 ;
        RECT 235.500 228.600 235.800 228.900 ;
        RECT 235.500 228.300 236.900 228.600 ;
        RECT 236.500 228.200 236.900 228.300 ;
        RECT 237.400 228.200 237.800 228.600 ;
        RECT 238.200 228.500 238.600 228.900 ;
        RECT 232.500 227.700 232.900 227.800 ;
        RECT 227.800 225.800 229.800 226.100 ;
        RECT 230.200 227.100 230.600 227.600 ;
        RECT 231.000 227.400 232.900 227.700 ;
        RECT 231.000 227.100 231.400 227.400 ;
        RECT 234.500 227.100 234.900 227.200 ;
        RECT 237.400 227.100 237.700 228.200 ;
        RECT 239.800 227.500 240.200 229.900 ;
        RECT 240.600 227.700 241.000 229.900 ;
        RECT 242.700 229.200 243.300 229.900 ;
        RECT 242.700 228.900 243.400 229.200 ;
        RECT 245.000 228.900 245.400 229.900 ;
        RECT 247.200 229.200 247.600 229.900 ;
        RECT 247.200 228.900 248.200 229.200 ;
        RECT 243.000 228.500 243.400 228.900 ;
        RECT 245.100 228.600 245.400 228.900 ;
        RECT 245.100 228.300 246.500 228.600 ;
        RECT 246.100 228.200 246.500 228.300 ;
        RECT 247.000 228.200 247.400 228.600 ;
        RECT 247.800 228.500 248.200 228.900 ;
        RECT 242.100 227.700 242.500 227.800 ;
        RECT 240.600 227.400 242.500 227.700 ;
        RECT 239.000 227.100 239.800 227.200 ;
        RECT 230.200 226.800 231.400 227.100 ;
        RECT 230.200 226.200 230.500 226.800 ;
        RECT 230.200 225.800 230.600 226.200 ;
        RECT 227.800 225.200 228.100 225.800 ;
        RECT 227.800 225.100 228.200 225.200 ;
        RECT 224.600 221.500 225.000 223.500 ;
        RECT 226.700 224.800 227.200 225.100 ;
        RECT 227.500 224.800 228.200 225.100 ;
        RECT 226.700 221.100 227.100 224.800 ;
        RECT 227.500 224.200 227.800 224.800 ;
        RECT 228.600 224.400 229.000 225.200 ;
        RECT 227.400 223.800 227.800 224.200 ;
        RECT 229.400 221.100 229.800 225.800 ;
        RECT 231.000 225.700 231.400 226.800 ;
        RECT 234.300 226.800 239.800 227.100 ;
        RECT 233.400 226.400 233.800 226.500 ;
        RECT 231.900 226.100 233.800 226.400 ;
        RECT 231.900 226.000 232.300 226.100 ;
        RECT 232.700 225.700 233.100 225.800 ;
        RECT 231.000 225.400 233.100 225.700 ;
        RECT 231.000 221.100 231.400 225.400 ;
        RECT 234.300 225.200 234.600 226.800 ;
        RECT 237.900 226.700 238.300 226.800 ;
        RECT 238.700 226.200 239.100 226.300 ;
        RECT 236.600 225.900 239.100 226.200 ;
        RECT 236.600 225.800 237.000 225.900 ;
        RECT 240.600 225.700 241.000 227.400 ;
        RECT 244.100 227.100 244.500 227.200 ;
        RECT 247.000 227.100 247.300 228.200 ;
        RECT 249.400 227.500 249.800 229.900 ;
        RECT 248.600 227.100 249.400 227.200 ;
        RECT 243.900 226.800 249.400 227.100 ;
        RECT 243.000 226.400 243.400 226.500 ;
        RECT 241.500 226.100 243.400 226.400 ;
        RECT 243.900 226.200 244.200 226.800 ;
        RECT 247.500 226.700 247.900 226.800 ;
        RECT 247.000 226.200 247.400 226.300 ;
        RECT 248.300 226.200 248.700 226.300 ;
        RECT 241.500 226.000 241.900 226.100 ;
        RECT 243.800 225.800 244.200 226.200 ;
        RECT 246.200 225.900 248.700 226.200 ;
        RECT 246.200 225.800 246.600 225.900 ;
        RECT 242.300 225.700 242.700 225.800 ;
        RECT 237.400 225.500 240.200 225.600 ;
        RECT 237.300 225.400 240.200 225.500 ;
        RECT 233.400 224.900 234.600 225.200 ;
        RECT 235.300 225.300 240.200 225.400 ;
        RECT 235.300 225.100 237.700 225.300 ;
        RECT 233.400 224.400 233.700 224.900 ;
        RECT 233.000 224.000 233.700 224.400 ;
        RECT 234.500 224.500 234.900 224.600 ;
        RECT 235.300 224.500 235.600 225.100 ;
        RECT 234.500 224.200 235.600 224.500 ;
        RECT 235.900 224.500 238.600 224.800 ;
        RECT 235.900 224.400 236.300 224.500 ;
        RECT 238.200 224.400 238.600 224.500 ;
        RECT 235.100 223.700 235.500 223.800 ;
        RECT 236.500 223.700 236.900 223.800 ;
        RECT 233.400 223.100 233.800 223.500 ;
        RECT 235.100 223.400 236.900 223.700 ;
        RECT 235.500 223.100 235.800 223.400 ;
        RECT 238.200 223.100 238.600 223.500 ;
        RECT 233.100 221.100 233.700 223.100 ;
        RECT 235.400 221.100 235.800 223.100 ;
        RECT 237.600 222.800 238.600 223.100 ;
        RECT 237.600 221.100 238.000 222.800 ;
        RECT 239.800 221.100 240.200 225.300 ;
        RECT 240.600 225.400 242.700 225.700 ;
        RECT 240.600 221.100 241.000 225.400 ;
        RECT 243.900 225.200 244.200 225.800 ;
        RECT 247.000 225.500 249.800 225.600 ;
        RECT 246.900 225.400 249.800 225.500 ;
        RECT 243.000 224.900 244.200 225.200 ;
        RECT 244.900 225.300 249.800 225.400 ;
        RECT 244.900 225.100 247.300 225.300 ;
        RECT 243.000 224.400 243.300 224.900 ;
        RECT 242.600 224.000 243.300 224.400 ;
        RECT 244.100 224.500 244.500 224.600 ;
        RECT 244.900 224.500 245.200 225.100 ;
        RECT 244.100 224.200 245.200 224.500 ;
        RECT 245.500 224.500 248.200 224.800 ;
        RECT 245.500 224.400 245.900 224.500 ;
        RECT 247.800 224.400 248.200 224.500 ;
        RECT 244.700 223.700 245.100 223.800 ;
        RECT 246.100 223.700 246.500 223.800 ;
        RECT 243.000 223.100 243.400 223.500 ;
        RECT 244.700 223.400 246.500 223.700 ;
        RECT 245.100 223.100 245.400 223.400 ;
        RECT 247.800 223.100 248.200 223.500 ;
        RECT 242.700 221.100 243.300 223.100 ;
        RECT 245.000 221.100 245.400 223.100 ;
        RECT 247.200 222.800 248.200 223.100 ;
        RECT 247.200 221.100 247.600 222.800 ;
        RECT 249.400 221.100 249.800 225.300 ;
        RECT 0.600 215.600 1.000 219.900 ;
        RECT 2.700 217.900 3.300 219.900 ;
        RECT 5.000 217.900 5.400 219.900 ;
        RECT 7.200 218.200 7.600 219.900 ;
        RECT 7.200 217.900 8.200 218.200 ;
        RECT 3.000 217.500 3.400 217.900 ;
        RECT 5.100 217.600 5.400 217.900 ;
        RECT 4.700 217.300 6.500 217.600 ;
        RECT 7.800 217.500 8.200 217.900 ;
        RECT 4.700 217.200 5.100 217.300 ;
        RECT 6.100 217.200 6.500 217.300 ;
        RECT 2.600 216.600 3.300 217.000 ;
        RECT 3.000 216.100 3.300 216.600 ;
        RECT 4.100 216.500 5.200 216.800 ;
        RECT 4.100 216.400 4.500 216.500 ;
        RECT 3.000 215.800 4.200 216.100 ;
        RECT 0.600 215.300 2.700 215.600 ;
        RECT 0.600 213.600 1.000 215.300 ;
        RECT 2.300 215.200 2.700 215.300 ;
        RECT 1.500 214.900 1.900 215.000 ;
        RECT 1.500 214.600 3.400 214.900 ;
        RECT 3.000 214.500 3.400 214.600 ;
        RECT 3.900 214.200 4.200 215.800 ;
        RECT 4.900 215.900 5.200 216.500 ;
        RECT 5.500 216.500 5.900 216.600 ;
        RECT 7.800 216.500 8.200 216.600 ;
        RECT 5.500 216.200 8.200 216.500 ;
        RECT 4.900 215.700 7.300 215.900 ;
        RECT 9.400 215.700 9.800 219.900 ;
        RECT 11.500 216.200 11.900 219.900 ;
        RECT 12.200 216.800 12.600 217.200 ;
        RECT 12.300 216.200 12.600 216.800 ;
        RECT 11.500 215.900 12.000 216.200 ;
        RECT 12.300 215.900 13.000 216.200 ;
        RECT 4.900 215.600 9.800 215.700 ;
        RECT 6.900 215.500 9.800 215.600 ;
        RECT 7.000 215.400 9.800 215.500 ;
        RECT 11.700 215.200 12.000 215.900 ;
        RECT 12.600 215.800 13.000 215.900 ;
        RECT 13.400 215.800 13.800 216.600 ;
        RECT 6.200 215.100 6.600 215.200 ;
        RECT 6.200 214.800 8.700 215.100 ;
        RECT 7.000 214.700 7.400 214.800 ;
        RECT 8.300 214.700 8.700 214.800 ;
        RECT 11.000 214.400 11.400 215.200 ;
        RECT 11.700 214.800 12.200 215.200 ;
        RECT 12.600 215.100 12.900 215.800 ;
        RECT 14.200 215.100 14.600 219.900 ;
        RECT 15.800 215.700 16.200 219.900 ;
        RECT 18.000 218.200 18.400 219.900 ;
        RECT 17.400 217.900 18.400 218.200 ;
        RECT 20.200 217.900 20.600 219.900 ;
        RECT 22.300 217.900 22.900 219.900 ;
        RECT 17.400 217.500 17.800 217.900 ;
        RECT 20.200 217.600 20.500 217.900 ;
        RECT 19.100 217.300 20.900 217.600 ;
        RECT 22.200 217.500 22.600 217.900 ;
        RECT 19.100 217.200 19.500 217.300 ;
        RECT 20.500 217.200 20.900 217.300 ;
        RECT 17.400 216.500 17.800 216.600 ;
        RECT 19.700 216.500 20.100 216.600 ;
        RECT 17.400 216.200 20.100 216.500 ;
        RECT 20.400 216.500 21.500 216.800 ;
        RECT 20.400 215.900 20.700 216.500 ;
        RECT 21.100 216.400 21.500 216.500 ;
        RECT 22.300 216.600 23.000 217.000 ;
        RECT 22.300 216.100 22.600 216.600 ;
        RECT 18.300 215.700 20.700 215.900 ;
        RECT 15.800 215.600 20.700 215.700 ;
        RECT 21.400 215.800 22.600 216.100 ;
        RECT 15.800 215.500 18.700 215.600 ;
        RECT 15.800 215.400 18.600 215.500 ;
        RECT 19.000 215.100 19.400 215.200 ;
        RECT 12.600 214.800 14.600 215.100 ;
        RECT 7.500 214.200 7.900 214.300 ;
        RECT 11.700 214.200 12.000 214.800 ;
        RECT 3.900 213.900 9.400 214.200 ;
        RECT 4.100 213.800 4.500 213.900 ;
        RECT 0.600 213.300 2.500 213.600 ;
        RECT 0.600 211.100 1.000 213.300 ;
        RECT 2.100 213.200 2.500 213.300 ;
        RECT 7.000 212.800 7.300 213.900 ;
        RECT 8.600 213.800 9.400 213.900 ;
        RECT 10.200 214.100 10.600 214.200 ;
        RECT 10.200 213.800 11.000 214.100 ;
        RECT 11.700 213.800 13.000 214.200 ;
        RECT 10.600 213.600 11.000 213.800 ;
        RECT 6.100 212.700 6.500 212.800 ;
        RECT 3.000 212.100 3.400 212.500 ;
        RECT 5.100 212.400 6.500 212.700 ;
        RECT 7.000 212.400 7.400 212.800 ;
        RECT 5.100 212.100 5.400 212.400 ;
        RECT 7.800 212.100 8.200 212.500 ;
        RECT 2.700 211.800 3.400 212.100 ;
        RECT 2.700 211.100 3.300 211.800 ;
        RECT 5.000 211.100 5.400 212.100 ;
        RECT 7.200 211.800 8.200 212.100 ;
        RECT 7.200 211.100 7.600 211.800 ;
        RECT 9.400 211.100 9.800 213.500 ;
        RECT 10.300 213.100 12.100 213.300 ;
        RECT 12.600 213.100 12.900 213.800 ;
        RECT 14.200 213.100 14.600 214.800 ;
        RECT 16.900 214.800 19.400 215.100 ;
        RECT 16.900 214.700 17.300 214.800 ;
        RECT 18.200 214.700 18.600 214.800 ;
        RECT 17.700 214.200 18.100 214.300 ;
        RECT 21.400 214.200 21.700 215.800 ;
        RECT 24.600 215.600 25.000 219.900 ;
        RECT 27.300 216.400 27.700 219.900 ;
        RECT 29.400 217.500 29.800 219.500 ;
        RECT 26.900 216.100 27.700 216.400 ;
        RECT 22.900 215.300 25.000 215.600 ;
        RECT 22.900 215.200 23.300 215.300 ;
        RECT 23.700 214.900 24.100 215.000 ;
        RECT 22.200 214.600 24.100 214.900 ;
        RECT 22.200 214.500 22.600 214.600 ;
        RECT 15.000 213.400 15.400 214.200 ;
        RECT 16.200 213.900 21.700 214.200 ;
        RECT 16.200 213.800 17.000 213.900 ;
        RECT 10.200 213.000 12.200 213.100 ;
        RECT 10.200 211.100 10.600 213.000 ;
        RECT 11.800 211.100 12.200 213.000 ;
        RECT 12.600 211.100 13.000 213.100 ;
        RECT 13.700 212.800 14.600 213.100 ;
        RECT 13.700 211.100 14.100 212.800 ;
        RECT 15.800 211.100 16.200 213.500 ;
        RECT 18.300 212.800 18.600 213.900 ;
        RECT 21.100 213.800 21.500 213.900 ;
        RECT 24.600 213.600 25.000 215.300 ;
        RECT 25.400 215.100 25.800 215.200 ;
        RECT 26.200 215.100 26.600 215.600 ;
        RECT 25.400 214.800 26.600 215.100 ;
        RECT 26.900 214.200 27.200 216.100 ;
        RECT 29.500 215.800 29.800 217.500 ;
        RECT 30.500 216.300 30.900 219.900 ;
        RECT 30.500 215.900 31.400 216.300 ;
        RECT 32.600 215.900 33.000 219.900 ;
        RECT 33.400 216.200 33.800 219.900 ;
        RECT 35.000 216.200 35.400 219.900 ;
        RECT 33.400 215.900 35.400 216.200 ;
        RECT 27.900 215.500 29.800 215.800 ;
        RECT 27.900 214.500 28.200 215.500 ;
        RECT 26.200 213.800 27.200 214.200 ;
        RECT 27.500 214.100 28.200 214.500 ;
        RECT 28.600 214.400 29.000 215.200 ;
        RECT 29.400 214.400 29.800 215.200 ;
        RECT 30.200 214.800 30.600 215.600 ;
        RECT 23.100 213.300 25.000 213.600 ;
        RECT 23.100 213.200 23.500 213.300 ;
        RECT 17.400 212.100 17.800 212.500 ;
        RECT 18.200 212.400 18.600 212.800 ;
        RECT 19.100 212.700 19.500 212.800 ;
        RECT 19.100 212.400 20.500 212.700 ;
        RECT 20.200 212.100 20.500 212.400 ;
        RECT 22.200 212.100 22.600 212.500 ;
        RECT 17.400 211.800 18.400 212.100 ;
        RECT 18.000 211.100 18.400 211.800 ;
        RECT 20.200 211.100 20.600 212.100 ;
        RECT 22.200 211.800 22.900 212.100 ;
        RECT 22.300 211.100 22.900 211.800 ;
        RECT 24.600 211.100 25.000 213.300 ;
        RECT 26.900 213.500 27.200 213.800 ;
        RECT 27.700 213.900 28.200 214.100 ;
        RECT 31.000 214.200 31.300 215.900 ;
        RECT 32.700 215.200 33.000 215.900 ;
        RECT 35.800 215.600 36.200 219.900 ;
        RECT 37.900 217.900 38.500 219.900 ;
        RECT 40.200 217.900 40.600 219.900 ;
        RECT 42.400 218.200 42.800 219.900 ;
        RECT 42.400 217.900 43.400 218.200 ;
        RECT 38.200 217.500 38.600 217.900 ;
        RECT 40.300 217.600 40.600 217.900 ;
        RECT 39.900 217.300 41.700 217.600 ;
        RECT 43.000 217.500 43.400 217.900 ;
        RECT 39.900 217.200 40.300 217.300 ;
        RECT 41.300 217.200 41.700 217.300 ;
        RECT 37.400 217.000 38.100 217.200 ;
        RECT 37.400 216.800 38.500 217.000 ;
        RECT 37.800 216.600 38.500 216.800 ;
        RECT 38.200 216.100 38.500 216.600 ;
        RECT 39.300 216.500 40.400 216.800 ;
        RECT 39.300 216.400 39.700 216.500 ;
        RECT 38.200 215.800 39.400 216.100 ;
        RECT 34.600 215.200 35.000 215.400 ;
        RECT 35.800 215.300 37.900 215.600 ;
        RECT 32.600 214.900 33.800 215.200 ;
        RECT 34.600 214.900 35.400 215.200 ;
        RECT 32.600 214.800 33.000 214.900 ;
        RECT 31.000 214.100 31.400 214.200 ;
        RECT 27.700 213.600 29.800 213.900 ;
        RECT 26.900 213.300 27.300 213.500 ;
        RECT 26.900 213.000 27.700 213.300 ;
        RECT 27.300 212.200 27.700 213.000 ;
        RECT 29.500 212.500 29.800 213.600 ;
        RECT 27.300 211.800 28.200 212.200 ;
        RECT 27.300 211.500 27.700 211.800 ;
        RECT 29.400 211.500 29.800 212.500 ;
        RECT 31.000 213.800 32.900 214.100 ;
        RECT 31.000 212.100 31.300 213.800 ;
        RECT 32.600 213.200 32.900 213.800 ;
        RECT 31.800 212.400 32.200 213.200 ;
        RECT 32.600 212.800 33.000 213.200 ;
        RECT 33.500 213.100 33.800 214.900 ;
        RECT 35.000 214.800 35.400 214.900 ;
        RECT 34.200 213.800 34.600 214.600 ;
        RECT 32.700 212.400 33.100 212.800 ;
        RECT 31.000 211.100 31.400 212.100 ;
        RECT 33.400 211.100 33.800 213.100 ;
        RECT 35.800 213.600 36.200 215.300 ;
        RECT 37.500 215.200 37.900 215.300 ;
        RECT 39.100 215.100 39.400 215.800 ;
        RECT 40.100 215.900 40.400 216.500 ;
        RECT 40.700 216.500 41.100 216.600 ;
        RECT 43.000 216.500 43.400 216.600 ;
        RECT 40.700 216.200 43.400 216.500 ;
        RECT 40.100 215.700 42.500 215.900 ;
        RECT 44.600 215.700 45.000 219.900 ;
        RECT 47.000 216.200 47.400 219.900 ;
        RECT 40.100 215.600 45.000 215.700 ;
        RECT 46.300 215.900 47.400 216.200 ;
        RECT 46.300 215.600 46.600 215.900 ;
        RECT 42.100 215.500 45.000 215.600 ;
        RECT 42.200 215.400 45.000 215.500 ;
        RECT 46.000 215.200 46.600 215.600 ;
        RECT 49.400 215.600 49.800 219.900 ;
        RECT 51.500 217.900 52.100 219.900 ;
        RECT 53.800 217.900 54.200 219.900 ;
        RECT 56.000 218.200 56.400 219.900 ;
        RECT 56.000 217.900 57.000 218.200 ;
        RECT 51.800 217.500 52.200 217.900 ;
        RECT 53.900 217.600 54.200 217.900 ;
        RECT 53.500 217.300 55.300 217.600 ;
        RECT 56.600 217.500 57.000 217.900 ;
        RECT 53.500 217.200 53.900 217.300 ;
        RECT 54.900 217.200 55.300 217.300 ;
        RECT 51.400 216.600 52.100 217.000 ;
        RECT 51.800 216.100 52.100 216.600 ;
        RECT 52.900 216.500 54.000 216.800 ;
        RECT 52.900 216.400 53.300 216.500 ;
        RECT 51.800 215.800 53.000 216.100 ;
        RECT 49.400 215.300 51.500 215.600 ;
        RECT 39.800 215.100 40.200 215.200 ;
        RECT 36.700 214.900 37.100 215.000 ;
        RECT 36.700 214.600 38.600 214.900 ;
        RECT 39.000 214.800 40.200 215.100 ;
        RECT 41.400 215.100 41.800 215.200 ;
        RECT 41.400 214.800 43.900 215.100 ;
        RECT 38.200 214.500 38.600 214.600 ;
        RECT 39.100 214.200 39.400 214.800 ;
        RECT 43.500 214.700 43.900 214.800 ;
        RECT 42.700 214.200 43.100 214.300 ;
        RECT 39.100 213.900 44.600 214.200 ;
        RECT 39.300 213.800 39.700 213.900 ;
        RECT 35.800 213.300 37.700 213.600 ;
        RECT 35.800 211.100 36.200 213.300 ;
        RECT 37.300 213.200 37.700 213.300 ;
        RECT 42.200 212.800 42.500 213.900 ;
        RECT 43.800 213.800 44.600 213.900 ;
        RECT 46.300 213.700 46.600 215.200 ;
        RECT 47.000 215.100 47.400 215.200 ;
        RECT 49.400 215.100 49.800 215.300 ;
        RECT 51.100 215.200 51.500 215.300 ;
        RECT 52.700 215.200 53.000 215.800 ;
        RECT 53.700 215.900 54.000 216.500 ;
        RECT 54.300 216.500 54.700 216.600 ;
        RECT 56.600 216.500 57.000 216.600 ;
        RECT 54.300 216.200 57.000 216.500 ;
        RECT 53.700 215.700 56.100 215.900 ;
        RECT 58.200 215.700 58.600 219.900 ;
        RECT 53.700 215.600 58.600 215.700 ;
        RECT 55.700 215.500 58.600 215.600 ;
        RECT 55.800 215.400 58.600 215.500 ;
        RECT 59.000 215.600 59.400 219.900 ;
        RECT 61.100 217.900 61.700 219.900 ;
        RECT 63.400 217.900 63.800 219.900 ;
        RECT 65.600 218.200 66.000 219.900 ;
        RECT 65.600 217.900 66.600 218.200 ;
        RECT 61.400 217.500 61.800 217.900 ;
        RECT 63.500 217.600 63.800 217.900 ;
        RECT 63.100 217.300 64.900 217.600 ;
        RECT 66.200 217.500 66.600 217.900 ;
        RECT 63.100 217.200 63.500 217.300 ;
        RECT 64.500 217.200 64.900 217.300 ;
        RECT 61.000 216.600 61.700 217.000 ;
        RECT 61.400 216.100 61.700 216.600 ;
        RECT 62.500 216.500 63.600 216.800 ;
        RECT 62.500 216.400 62.900 216.500 ;
        RECT 61.400 215.800 62.600 216.100 ;
        RECT 59.000 215.300 61.100 215.600 ;
        RECT 47.000 214.800 49.800 215.100 ;
        RECT 47.000 214.400 47.400 214.800 ;
        RECT 41.300 212.700 41.700 212.800 ;
        RECT 38.200 212.100 38.600 212.500 ;
        RECT 40.300 212.400 41.700 212.700 ;
        RECT 42.200 212.400 42.600 212.800 ;
        RECT 40.300 212.100 40.600 212.400 ;
        RECT 43.000 212.100 43.400 212.500 ;
        RECT 37.900 211.800 38.600 212.100 ;
        RECT 37.900 211.100 38.500 211.800 ;
        RECT 40.200 211.100 40.600 212.100 ;
        RECT 42.400 211.800 43.400 212.100 ;
        RECT 42.400 211.100 42.800 211.800 ;
        RECT 44.600 211.100 45.000 213.500 ;
        RECT 46.300 213.400 47.400 213.700 ;
        RECT 47.000 211.100 47.400 213.400 ;
        RECT 49.400 213.600 49.800 214.800 ;
        RECT 50.300 214.900 50.700 215.000 ;
        RECT 50.300 214.600 52.200 214.900 ;
        RECT 52.600 214.800 53.000 215.200 ;
        RECT 55.000 215.100 55.400 215.200 ;
        RECT 55.000 214.800 57.500 215.100 ;
        RECT 51.800 214.500 52.200 214.600 ;
        RECT 52.700 214.200 53.000 214.800 ;
        RECT 55.800 214.700 56.200 214.800 ;
        RECT 57.100 214.700 57.500 214.800 ;
        RECT 56.300 214.200 56.700 214.300 ;
        RECT 52.700 213.900 58.200 214.200 ;
        RECT 52.900 213.800 53.300 213.900 ;
        RECT 49.400 213.300 51.300 213.600 ;
        RECT 49.400 211.100 49.800 213.300 ;
        RECT 50.900 213.200 51.300 213.300 ;
        RECT 55.800 212.800 56.100 213.900 ;
        RECT 57.400 213.800 58.200 213.900 ;
        RECT 59.000 213.600 59.400 215.300 ;
        RECT 60.700 215.200 61.100 215.300 ;
        RECT 62.300 215.200 62.600 215.800 ;
        RECT 63.300 215.900 63.600 216.500 ;
        RECT 63.900 216.500 64.300 216.600 ;
        RECT 66.200 216.500 66.600 216.600 ;
        RECT 63.900 216.200 66.600 216.500 ;
        RECT 63.300 215.700 65.700 215.900 ;
        RECT 67.800 215.700 68.200 219.900 ;
        RECT 69.700 217.200 70.100 219.900 ;
        RECT 69.000 216.800 69.400 217.200 ;
        RECT 69.700 216.800 70.600 217.200 ;
        RECT 69.000 216.200 69.300 216.800 ;
        RECT 69.700 216.200 70.100 216.800 ;
        RECT 68.600 215.900 69.300 216.200 ;
        RECT 69.600 215.900 70.100 216.200 ;
        RECT 71.800 216.200 72.200 219.900 ;
        RECT 73.400 216.200 73.800 219.900 ;
        RECT 71.800 215.900 73.800 216.200 ;
        RECT 74.200 215.900 74.600 219.900 ;
        RECT 75.000 216.200 75.400 219.900 ;
        RECT 76.600 216.400 77.000 219.900 ;
        RECT 79.000 216.400 79.400 219.900 ;
        RECT 75.000 215.900 76.300 216.200 ;
        RECT 76.600 215.900 77.100 216.400 ;
        RECT 68.600 215.800 69.000 215.900 ;
        RECT 63.300 215.600 68.200 215.700 ;
        RECT 65.300 215.500 68.200 215.600 ;
        RECT 65.400 215.400 68.200 215.500 ;
        RECT 59.900 214.900 60.300 215.000 ;
        RECT 59.900 214.600 61.800 214.900 ;
        RECT 62.200 214.800 62.600 215.200 ;
        RECT 64.600 215.100 65.000 215.200 ;
        RECT 64.600 214.800 67.100 215.100 ;
        RECT 61.400 214.500 61.800 214.600 ;
        RECT 62.300 214.200 62.600 214.800 ;
        RECT 65.400 214.700 65.800 214.800 ;
        RECT 66.700 214.700 67.100 214.800 ;
        RECT 65.900 214.200 66.300 214.300 ;
        RECT 69.600 214.200 69.900 215.900 ;
        RECT 72.200 215.200 72.600 215.400 ;
        RECT 74.200 215.200 74.500 215.900 ;
        RECT 70.200 214.400 70.600 215.200 ;
        RECT 71.800 214.900 72.600 215.200 ;
        RECT 73.400 214.900 74.600 215.200 ;
        RECT 71.800 214.800 72.200 214.900 ;
        RECT 62.300 213.900 67.800 214.200 ;
        RECT 62.500 213.800 62.900 213.900 ;
        RECT 54.900 212.700 55.300 212.800 ;
        RECT 51.800 212.100 52.200 212.500 ;
        RECT 53.900 212.400 55.300 212.700 ;
        RECT 55.800 212.400 56.200 212.800 ;
        RECT 53.900 212.100 54.200 212.400 ;
        RECT 56.600 212.100 57.000 212.500 ;
        RECT 51.500 211.800 52.200 212.100 ;
        RECT 51.500 211.100 52.100 211.800 ;
        RECT 53.800 211.100 54.200 212.100 ;
        RECT 56.000 211.800 57.000 212.100 ;
        RECT 56.000 211.100 56.400 211.800 ;
        RECT 58.200 211.100 58.600 213.500 ;
        RECT 59.000 213.300 60.900 213.600 ;
        RECT 59.000 211.100 59.400 213.300 ;
        RECT 60.500 213.200 60.900 213.300 ;
        RECT 65.400 212.800 65.700 213.900 ;
        RECT 67.000 213.800 67.800 213.900 ;
        RECT 68.600 213.800 69.900 214.200 ;
        RECT 71.000 214.100 71.400 214.200 ;
        RECT 70.600 213.800 71.400 214.100 ;
        RECT 72.600 213.800 73.000 214.600 ;
        RECT 64.500 212.700 64.900 212.800 ;
        RECT 61.400 212.100 61.800 212.500 ;
        RECT 63.500 212.400 64.900 212.700 ;
        RECT 65.400 212.400 65.800 212.800 ;
        RECT 63.500 212.100 63.800 212.400 ;
        RECT 66.200 212.100 66.600 212.500 ;
        RECT 61.100 211.800 61.800 212.100 ;
        RECT 61.100 211.100 61.700 211.800 ;
        RECT 63.400 211.100 63.800 212.100 ;
        RECT 65.600 211.800 66.600 212.100 ;
        RECT 65.600 211.100 66.000 211.800 ;
        RECT 67.800 211.100 68.200 213.500 ;
        RECT 68.700 213.100 69.000 213.800 ;
        RECT 70.600 213.600 71.000 213.800 ;
        RECT 69.500 213.100 71.300 213.300 ;
        RECT 73.400 213.100 73.700 214.900 ;
        RECT 74.200 214.800 74.600 214.900 ;
        RECT 75.000 214.800 75.500 215.200 ;
        RECT 75.100 214.400 75.500 214.800 ;
        RECT 76.000 214.900 76.300 215.900 ;
        RECT 76.000 214.500 76.500 214.900 ;
        RECT 76.000 213.700 76.300 214.500 ;
        RECT 76.800 214.200 77.100 215.900 ;
        RECT 78.900 215.900 79.400 216.400 ;
        RECT 80.600 216.200 81.000 219.900 ;
        RECT 79.700 215.900 81.000 216.200 ;
        RECT 78.900 214.200 79.200 215.900 ;
        RECT 79.700 214.900 80.000 215.900 ;
        RECT 81.400 215.700 81.800 219.900 ;
        RECT 83.600 218.200 84.000 219.900 ;
        RECT 83.000 217.900 84.000 218.200 ;
        RECT 85.800 217.900 86.200 219.900 ;
        RECT 87.900 217.900 88.500 219.900 ;
        RECT 83.000 217.500 83.400 217.900 ;
        RECT 85.800 217.600 86.100 217.900 ;
        RECT 84.700 217.300 86.500 217.600 ;
        RECT 87.800 217.500 88.200 217.900 ;
        RECT 84.700 217.200 85.100 217.300 ;
        RECT 86.100 217.200 86.500 217.300 ;
        RECT 83.000 216.500 83.400 216.600 ;
        RECT 85.300 216.500 85.700 216.600 ;
        RECT 83.000 216.200 85.700 216.500 ;
        RECT 86.000 216.500 87.100 216.800 ;
        RECT 86.000 215.900 86.300 216.500 ;
        RECT 86.700 216.400 87.100 216.500 ;
        RECT 87.900 216.600 88.600 217.000 ;
        RECT 87.900 216.100 88.200 216.600 ;
        RECT 83.900 215.700 86.300 215.900 ;
        RECT 81.400 215.600 86.300 215.700 ;
        RECT 87.000 215.800 88.200 216.100 ;
        RECT 81.400 215.500 84.300 215.600 ;
        RECT 81.400 215.400 84.200 215.500 ;
        RECT 79.500 214.500 80.000 214.900 ;
        RECT 76.600 213.800 77.100 214.200 ;
        RECT 78.200 214.100 78.600 214.200 ;
        RECT 78.900 214.100 79.400 214.200 ;
        RECT 78.200 213.800 79.400 214.100 ;
        RECT 75.000 213.400 76.300 213.700 ;
        RECT 68.600 211.100 69.000 213.100 ;
        RECT 69.400 213.000 71.400 213.100 ;
        RECT 69.400 211.100 69.800 213.000 ;
        RECT 71.000 211.100 71.400 213.000 ;
        RECT 73.400 211.100 73.800 213.100 ;
        RECT 74.200 212.800 74.600 213.200 ;
        RECT 74.100 212.400 74.500 212.800 ;
        RECT 75.000 211.100 75.400 213.400 ;
        RECT 76.800 213.100 77.100 213.800 ;
        RECT 76.600 212.800 77.100 213.100 ;
        RECT 78.900 213.100 79.200 213.800 ;
        RECT 79.700 213.700 80.000 214.500 ;
        RECT 80.500 214.800 81.000 215.200 ;
        RECT 84.600 215.100 85.000 215.200 ;
        RECT 82.500 214.800 85.000 215.100 ;
        RECT 80.500 214.400 80.900 214.800 ;
        RECT 82.500 214.700 82.900 214.800 ;
        RECT 83.300 214.200 83.700 214.300 ;
        RECT 87.000 214.200 87.300 215.800 ;
        RECT 90.200 215.600 90.600 219.900 ;
        RECT 92.300 216.200 92.700 219.900 ;
        RECT 93.000 216.800 93.400 217.200 ;
        RECT 93.100 216.200 93.400 216.800 ;
        RECT 91.800 215.800 92.800 216.200 ;
        RECT 93.100 216.100 93.800 216.200 ;
        RECT 95.000 216.100 95.400 219.900 ;
        RECT 93.100 215.900 95.400 216.100 ;
        RECT 93.400 215.800 95.400 215.900 ;
        RECT 95.800 215.800 96.200 216.600 ;
        RECT 98.500 216.400 98.900 219.900 ;
        RECT 100.600 217.500 101.000 219.500 ;
        RECT 98.100 216.100 98.900 216.400 ;
        RECT 88.500 215.300 90.600 215.600 ;
        RECT 88.500 215.200 88.900 215.300 ;
        RECT 89.300 214.900 89.700 215.000 ;
        RECT 87.800 214.600 89.700 214.900 ;
        RECT 87.800 214.500 88.200 214.600 ;
        RECT 81.800 213.900 87.300 214.200 ;
        RECT 81.800 213.800 82.600 213.900 ;
        RECT 83.800 213.800 84.200 213.900 ;
        RECT 86.700 213.800 87.100 213.900 ;
        RECT 79.700 213.400 81.000 213.700 ;
        RECT 78.900 212.800 79.400 213.100 ;
        RECT 76.600 211.100 77.000 212.800 ;
        RECT 79.000 211.100 79.400 212.800 ;
        RECT 80.600 211.100 81.000 213.400 ;
        RECT 81.400 211.100 81.800 213.500 ;
        RECT 83.900 212.800 84.200 213.800 ;
        RECT 90.200 213.600 90.600 215.300 ;
        RECT 91.800 214.400 92.200 215.200 ;
        RECT 92.500 214.200 92.800 215.800 ;
        RECT 91.000 214.100 91.400 214.200 ;
        RECT 91.000 213.800 91.800 214.100 ;
        RECT 92.500 213.800 93.800 214.200 ;
        RECT 91.400 213.600 91.800 213.800 ;
        RECT 88.700 213.300 90.600 213.600 ;
        RECT 88.700 213.200 89.100 213.300 ;
        RECT 83.000 212.100 83.400 212.500 ;
        RECT 83.800 212.400 84.200 212.800 ;
        RECT 84.700 212.700 85.100 212.800 ;
        RECT 84.700 212.400 86.100 212.700 ;
        RECT 85.800 212.100 86.100 212.400 ;
        RECT 87.800 212.100 88.200 212.500 ;
        RECT 83.000 211.800 84.000 212.100 ;
        RECT 83.600 211.100 84.000 211.800 ;
        RECT 85.800 211.100 86.200 212.100 ;
        RECT 87.800 211.800 88.500 212.100 ;
        RECT 87.900 211.100 88.500 211.800 ;
        RECT 90.200 211.100 90.600 213.300 ;
        RECT 91.100 213.100 92.900 213.300 ;
        RECT 93.400 213.100 93.700 213.800 ;
        RECT 94.200 213.400 94.600 214.200 ;
        RECT 95.000 213.100 95.400 215.800 ;
        RECT 96.600 215.100 97.000 215.200 ;
        RECT 97.400 215.100 97.800 215.600 ;
        RECT 96.600 214.800 97.800 215.100 ;
        RECT 98.100 214.200 98.400 216.100 ;
        RECT 100.700 215.800 101.000 217.500 ;
        RECT 103.400 216.800 103.800 217.200 ;
        RECT 103.400 216.200 103.700 216.800 ;
        RECT 104.100 216.200 104.500 219.900 ;
        RECT 102.200 216.100 102.600 216.200 ;
        RECT 103.000 216.100 103.700 216.200 ;
        RECT 102.200 215.900 103.700 216.100 ;
        RECT 104.000 215.900 104.500 216.200 ;
        RECT 102.200 215.800 103.400 215.900 ;
        RECT 99.100 215.500 101.000 215.800 ;
        RECT 99.100 214.500 99.400 215.500 ;
        RECT 97.400 213.800 98.400 214.200 ;
        RECT 98.700 214.100 99.400 214.500 ;
        RECT 99.800 214.400 100.200 215.200 ;
        RECT 100.600 215.100 101.000 215.200 ;
        RECT 101.400 215.100 101.800 215.200 ;
        RECT 100.600 214.800 101.800 215.100 ;
        RECT 100.600 214.400 101.000 214.800 ;
        RECT 104.000 214.200 104.300 215.900 ;
        RECT 104.600 214.400 105.000 215.200 ;
        RECT 106.200 214.800 106.600 215.200 ;
        RECT 106.200 214.200 106.500 214.800 ;
        RECT 98.100 213.500 98.400 213.800 ;
        RECT 98.900 213.900 99.400 214.100 ;
        RECT 98.900 213.600 101.000 213.900 ;
        RECT 103.000 213.800 104.300 214.200 ;
        RECT 105.400 214.100 105.800 214.200 ;
        RECT 105.000 213.800 105.800 214.100 ;
        RECT 98.100 213.300 98.500 213.500 ;
        RECT 91.000 213.000 93.000 213.100 ;
        RECT 91.000 211.100 91.400 213.000 ;
        RECT 92.600 211.100 93.000 213.000 ;
        RECT 93.400 211.100 93.800 213.100 ;
        RECT 95.000 212.800 95.900 213.100 ;
        RECT 98.100 213.000 98.900 213.300 ;
        RECT 95.500 211.100 95.900 212.800 ;
        RECT 98.500 212.200 98.900 213.000 ;
        RECT 100.700 212.500 101.000 213.600 ;
        RECT 103.100 213.100 103.400 213.800 ;
        RECT 105.000 213.600 105.400 213.800 ;
        RECT 106.200 213.400 106.600 214.200 ;
        RECT 103.900 213.100 105.700 213.300 ;
        RECT 107.000 213.100 107.400 219.900 ;
        RECT 107.800 215.800 108.200 216.600 ;
        RECT 108.600 215.600 109.000 219.900 ;
        RECT 110.700 217.900 111.300 219.900 ;
        RECT 113.000 217.900 113.400 219.900 ;
        RECT 115.200 218.200 115.600 219.900 ;
        RECT 115.200 217.900 116.200 218.200 ;
        RECT 111.000 217.500 111.400 217.900 ;
        RECT 113.100 217.600 113.400 217.900 ;
        RECT 112.700 217.300 114.500 217.600 ;
        RECT 115.800 217.500 116.200 217.900 ;
        RECT 112.700 217.200 113.100 217.300 ;
        RECT 114.100 217.200 114.500 217.300 ;
        RECT 110.600 216.600 111.300 217.000 ;
        RECT 111.000 216.100 111.300 216.600 ;
        RECT 112.100 216.500 113.200 216.800 ;
        RECT 112.100 216.400 112.500 216.500 ;
        RECT 111.000 215.800 112.200 216.100 ;
        RECT 108.600 215.300 110.700 215.600 ;
        RECT 108.600 213.600 109.000 215.300 ;
        RECT 110.300 215.200 110.700 215.300 ;
        RECT 109.500 214.900 109.900 215.000 ;
        RECT 109.500 214.600 111.400 214.900 ;
        RECT 111.000 214.500 111.400 214.600 ;
        RECT 111.900 214.200 112.200 215.800 ;
        RECT 112.900 215.900 113.200 216.500 ;
        RECT 113.500 216.500 113.900 216.600 ;
        RECT 115.800 216.500 116.200 216.600 ;
        RECT 113.500 216.200 116.200 216.500 ;
        RECT 112.900 215.700 115.300 215.900 ;
        RECT 117.400 215.700 117.800 219.900 ;
        RECT 112.900 215.600 117.800 215.700 ;
        RECT 114.900 215.500 117.800 215.600 ;
        RECT 115.000 215.400 117.800 215.500 ;
        RECT 114.200 215.100 114.600 215.200 ;
        RECT 114.200 214.800 116.700 215.100 ;
        RECT 116.300 214.700 116.700 214.800 ;
        RECT 115.500 214.200 115.900 214.300 ;
        RECT 111.800 213.900 117.400 214.200 ;
        RECT 111.800 213.800 112.500 213.900 ;
        RECT 108.600 213.300 110.500 213.600 ;
        RECT 98.200 211.800 98.900 212.200 ;
        RECT 98.500 211.500 98.900 211.800 ;
        RECT 100.600 211.500 101.000 212.500 ;
        RECT 103.000 211.100 103.400 213.100 ;
        RECT 103.800 213.000 105.800 213.100 ;
        RECT 103.800 211.100 104.200 213.000 ;
        RECT 105.400 211.100 105.800 213.000 ;
        RECT 107.000 212.800 107.900 213.100 ;
        RECT 107.500 211.100 107.900 212.800 ;
        RECT 108.600 211.100 109.000 213.300 ;
        RECT 110.100 213.200 110.500 213.300 ;
        RECT 115.000 212.800 115.300 213.900 ;
        RECT 116.600 213.800 117.400 213.900 ;
        RECT 114.100 212.700 114.500 212.800 ;
        RECT 111.000 212.100 111.400 212.500 ;
        RECT 113.100 212.400 114.500 212.700 ;
        RECT 115.000 212.400 115.400 212.800 ;
        RECT 113.100 212.100 113.400 212.400 ;
        RECT 115.800 212.100 116.200 212.500 ;
        RECT 110.700 211.800 111.400 212.100 ;
        RECT 110.700 211.100 111.300 211.800 ;
        RECT 113.000 211.100 113.400 212.100 ;
        RECT 115.200 211.800 116.200 212.100 ;
        RECT 115.200 211.100 115.600 211.800 ;
        RECT 117.400 211.100 117.800 213.500 ;
        RECT 119.000 213.100 119.400 219.900 ;
        RECT 120.600 217.100 121.000 219.900 ;
        RECT 122.700 217.900 123.300 219.900 ;
        RECT 125.000 217.900 125.400 219.900 ;
        RECT 127.200 218.200 127.600 219.900 ;
        RECT 127.200 217.900 128.200 218.200 ;
        RECT 123.000 217.500 123.400 217.900 ;
        RECT 125.100 217.600 125.400 217.900 ;
        RECT 124.700 217.300 126.500 217.600 ;
        RECT 127.800 217.500 128.200 217.900 ;
        RECT 124.700 217.200 125.100 217.300 ;
        RECT 126.100 217.200 126.500 217.300 ;
        RECT 119.800 216.800 121.000 217.100 ;
        RECT 119.800 215.800 120.200 216.800 ;
        RECT 120.600 215.600 121.000 216.800 ;
        RECT 122.600 216.600 123.300 217.000 ;
        RECT 123.000 216.100 123.300 216.600 ;
        RECT 124.100 216.500 125.200 216.800 ;
        RECT 124.100 216.400 124.500 216.500 ;
        RECT 123.000 215.800 124.200 216.100 ;
        RECT 120.600 215.300 122.700 215.600 ;
        RECT 120.600 213.600 121.000 215.300 ;
        RECT 122.300 215.200 122.700 215.300 ;
        RECT 123.900 215.100 124.200 215.800 ;
        RECT 124.900 215.900 125.200 216.500 ;
        RECT 125.500 216.500 125.900 216.600 ;
        RECT 127.800 216.500 128.200 216.600 ;
        RECT 125.500 216.200 128.200 216.500 ;
        RECT 124.900 215.700 127.300 215.900 ;
        RECT 129.400 215.700 129.800 219.900 ;
        RECT 131.500 216.200 131.900 219.900 ;
        RECT 132.200 216.800 132.600 217.200 ;
        RECT 132.300 216.200 132.600 216.800 ;
        RECT 131.500 215.900 132.000 216.200 ;
        RECT 132.300 215.900 133.000 216.200 ;
        RECT 124.900 215.600 129.800 215.700 ;
        RECT 126.900 215.500 129.800 215.600 ;
        RECT 127.000 215.400 129.800 215.500 ;
        RECT 124.600 215.100 125.000 215.200 ;
        RECT 121.500 214.900 121.900 215.000 ;
        RECT 121.500 214.600 123.400 214.900 ;
        RECT 123.800 214.800 125.000 215.100 ;
        RECT 126.200 215.100 126.600 215.200 ;
        RECT 126.200 214.800 128.700 215.100 ;
        RECT 123.000 214.500 123.400 214.600 ;
        RECT 123.900 214.200 124.200 214.800 ;
        RECT 128.300 214.700 128.700 214.800 ;
        RECT 131.000 214.400 131.400 215.200 ;
        RECT 127.500 214.200 127.900 214.300 ;
        RECT 131.700 214.200 132.000 215.900 ;
        RECT 132.600 215.800 133.000 215.900 ;
        RECT 133.400 215.800 133.800 216.600 ;
        RECT 132.600 215.100 132.900 215.800 ;
        RECT 134.200 215.100 134.600 219.900 ;
        RECT 135.800 215.700 136.200 219.900 ;
        RECT 138.000 218.200 138.400 219.900 ;
        RECT 137.400 217.900 138.400 218.200 ;
        RECT 140.200 217.900 140.600 219.900 ;
        RECT 142.300 217.900 142.900 219.900 ;
        RECT 137.400 217.500 137.800 217.900 ;
        RECT 140.200 217.600 140.500 217.900 ;
        RECT 139.100 217.300 140.900 217.600 ;
        RECT 142.200 217.500 142.600 217.900 ;
        RECT 139.100 217.200 139.500 217.300 ;
        RECT 140.500 217.200 140.900 217.300 ;
        RECT 137.400 216.500 137.800 216.600 ;
        RECT 139.700 216.500 140.100 216.600 ;
        RECT 137.400 216.200 140.100 216.500 ;
        RECT 140.400 216.500 141.500 216.800 ;
        RECT 140.400 215.900 140.700 216.500 ;
        RECT 141.100 216.400 141.500 216.500 ;
        RECT 142.300 216.600 143.000 217.000 ;
        RECT 142.300 216.100 142.600 216.600 ;
        RECT 138.300 215.700 140.700 215.900 ;
        RECT 135.800 215.600 140.700 215.700 ;
        RECT 141.400 215.800 142.600 216.100 ;
        RECT 135.800 215.500 138.700 215.600 ;
        RECT 135.800 215.400 138.600 215.500 ;
        RECT 139.000 215.100 139.400 215.200 ;
        RECT 132.600 214.800 134.600 215.100 ;
        RECT 123.900 213.900 129.400 214.200 ;
        RECT 124.100 213.800 124.500 213.900 ;
        RECT 120.600 213.300 122.500 213.600 ;
        RECT 119.000 212.800 119.900 213.100 ;
        RECT 119.500 212.200 119.900 212.800 ;
        RECT 119.500 211.800 120.200 212.200 ;
        RECT 119.500 211.100 119.900 211.800 ;
        RECT 120.600 211.100 121.000 213.300 ;
        RECT 122.100 213.200 122.500 213.300 ;
        RECT 127.000 212.800 127.300 213.900 ;
        RECT 128.600 213.800 129.400 213.900 ;
        RECT 130.200 214.100 130.600 214.200 ;
        RECT 131.700 214.100 133.000 214.200 ;
        RECT 133.400 214.100 133.800 214.200 ;
        RECT 130.200 213.800 131.000 214.100 ;
        RECT 131.700 213.800 133.800 214.100 ;
        RECT 130.600 213.600 131.000 213.800 ;
        RECT 126.100 212.700 126.500 212.800 ;
        RECT 123.000 212.100 123.400 212.500 ;
        RECT 125.100 212.400 126.500 212.700 ;
        RECT 127.000 212.400 127.400 212.800 ;
        RECT 125.100 212.100 125.400 212.400 ;
        RECT 127.800 212.100 128.200 212.500 ;
        RECT 122.700 211.800 123.400 212.100 ;
        RECT 122.700 211.100 123.300 211.800 ;
        RECT 125.000 211.100 125.400 212.100 ;
        RECT 127.200 211.800 128.200 212.100 ;
        RECT 127.200 211.100 127.600 211.800 ;
        RECT 129.400 211.100 129.800 213.500 ;
        RECT 130.300 213.100 132.100 213.300 ;
        RECT 132.600 213.100 132.900 213.800 ;
        RECT 134.200 213.100 134.600 214.800 ;
        RECT 136.900 214.800 139.400 215.100 ;
        RECT 136.900 214.700 137.300 214.800 ;
        RECT 138.200 214.700 138.600 214.800 ;
        RECT 137.700 214.200 138.100 214.300 ;
        RECT 141.400 214.200 141.700 215.800 ;
        RECT 144.600 215.600 145.000 219.900 ;
        RECT 142.900 215.300 145.000 215.600 ;
        RECT 142.900 215.200 143.300 215.300 ;
        RECT 143.700 214.900 144.100 215.000 ;
        RECT 142.200 214.600 144.100 214.900 ;
        RECT 142.200 214.500 142.600 214.600 ;
        RECT 135.000 213.400 135.400 214.200 ;
        RECT 136.200 213.900 141.700 214.200 ;
        RECT 136.200 213.800 137.000 213.900 ;
        RECT 130.200 213.000 132.200 213.100 ;
        RECT 130.200 211.100 130.600 213.000 ;
        RECT 131.800 211.100 132.200 213.000 ;
        RECT 132.600 211.100 133.000 213.100 ;
        RECT 133.700 212.800 134.600 213.100 ;
        RECT 133.700 211.100 134.100 212.800 ;
        RECT 135.800 211.100 136.200 213.500 ;
        RECT 138.300 212.800 138.600 213.900 ;
        RECT 141.100 213.800 141.500 213.900 ;
        RECT 144.600 213.600 145.000 215.300 ;
        RECT 143.100 213.300 145.000 213.600 ;
        RECT 143.100 213.200 143.500 213.300 ;
        RECT 137.400 212.100 137.800 212.500 ;
        RECT 138.200 212.400 138.600 212.800 ;
        RECT 139.100 212.700 139.500 212.800 ;
        RECT 139.100 212.400 140.500 212.700 ;
        RECT 140.200 212.100 140.500 212.400 ;
        RECT 142.200 212.100 142.600 212.500 ;
        RECT 137.400 211.800 138.400 212.100 ;
        RECT 138.000 211.100 138.400 211.800 ;
        RECT 140.200 211.100 140.600 212.100 ;
        RECT 142.200 211.800 142.900 212.100 ;
        RECT 142.300 211.100 142.900 211.800 ;
        RECT 144.600 211.100 145.000 213.300 ;
        RECT 145.400 215.600 145.800 219.900 ;
        RECT 147.500 217.900 148.100 219.900 ;
        RECT 149.800 217.900 150.200 219.900 ;
        RECT 152.000 218.200 152.400 219.900 ;
        RECT 152.000 217.900 153.000 218.200 ;
        RECT 147.800 217.500 148.200 217.900 ;
        RECT 149.900 217.600 150.200 217.900 ;
        RECT 149.500 217.300 151.300 217.600 ;
        RECT 152.600 217.500 153.000 217.900 ;
        RECT 149.500 217.200 149.900 217.300 ;
        RECT 150.900 217.200 151.300 217.300 ;
        RECT 147.400 216.600 148.100 217.000 ;
        RECT 147.800 216.100 148.100 216.600 ;
        RECT 148.900 216.500 150.000 216.800 ;
        RECT 148.900 216.400 149.300 216.500 ;
        RECT 147.800 215.800 149.000 216.100 ;
        RECT 145.400 215.300 147.500 215.600 ;
        RECT 145.400 213.600 145.800 215.300 ;
        RECT 147.100 215.200 147.500 215.300 ;
        RECT 146.300 214.900 146.700 215.000 ;
        RECT 146.300 214.600 148.200 214.900 ;
        RECT 147.800 214.500 148.200 214.600 ;
        RECT 148.700 214.200 149.000 215.800 ;
        RECT 149.700 215.900 150.000 216.500 ;
        RECT 150.300 216.500 150.700 216.600 ;
        RECT 152.600 216.500 153.000 216.600 ;
        RECT 150.300 216.200 153.000 216.500 ;
        RECT 149.700 215.700 152.100 215.900 ;
        RECT 154.200 215.700 154.600 219.900 ;
        RECT 157.900 216.200 158.300 219.900 ;
        RECT 158.600 216.800 159.000 217.200 ;
        RECT 158.700 216.200 159.000 216.800 ;
        RECT 157.900 215.900 158.400 216.200 ;
        RECT 158.700 215.900 159.400 216.200 ;
        RECT 149.700 215.600 154.600 215.700 ;
        RECT 151.700 215.500 154.600 215.600 ;
        RECT 151.800 215.400 154.600 215.500 ;
        RECT 151.000 215.100 151.400 215.200 ;
        RECT 151.000 214.800 153.500 215.100 ;
        RECT 153.100 214.700 153.500 214.800 ;
        RECT 157.400 214.400 157.800 215.200 ;
        RECT 152.300 214.200 152.700 214.300 ;
        RECT 158.100 214.200 158.400 215.900 ;
        RECT 159.000 215.800 159.400 215.900 ;
        RECT 159.800 215.800 160.200 216.600 ;
        RECT 159.000 215.100 159.300 215.800 ;
        RECT 160.600 215.100 161.000 219.900 ;
        RECT 163.500 216.200 163.900 219.900 ;
        RECT 164.200 216.800 164.600 217.200 ;
        RECT 164.300 216.200 164.600 216.800 ;
        RECT 163.500 215.900 164.000 216.200 ;
        RECT 164.300 215.900 165.000 216.200 ;
        RECT 159.000 214.800 161.000 215.100 ;
        RECT 148.700 213.900 154.200 214.200 ;
        RECT 148.900 213.800 149.300 213.900 ;
        RECT 145.400 213.300 147.300 213.600 ;
        RECT 145.400 211.100 145.800 213.300 ;
        RECT 146.900 213.200 147.300 213.300 ;
        RECT 151.800 212.800 152.100 213.900 ;
        RECT 153.400 213.800 154.200 213.900 ;
        RECT 156.600 214.100 157.000 214.200 ;
        RECT 156.600 213.800 157.400 214.100 ;
        RECT 158.100 213.800 159.400 214.200 ;
        RECT 157.000 213.600 157.400 213.800 ;
        RECT 150.900 212.700 151.300 212.800 ;
        RECT 147.800 212.100 148.200 212.500 ;
        RECT 149.900 212.400 151.300 212.700 ;
        RECT 151.800 212.400 152.200 212.800 ;
        RECT 149.900 212.100 150.200 212.400 ;
        RECT 152.600 212.100 153.000 212.500 ;
        RECT 147.500 211.800 148.200 212.100 ;
        RECT 147.500 211.100 148.100 211.800 ;
        RECT 149.800 211.100 150.200 212.100 ;
        RECT 152.000 211.800 153.000 212.100 ;
        RECT 152.000 211.100 152.400 211.800 ;
        RECT 154.200 211.100 154.600 213.500 ;
        RECT 156.700 213.100 158.500 213.300 ;
        RECT 159.000 213.100 159.300 213.800 ;
        RECT 160.600 213.100 161.000 214.800 ;
        RECT 163.000 214.400 163.400 215.200 ;
        RECT 163.700 214.200 164.000 215.900 ;
        RECT 164.600 215.800 165.000 215.900 ;
        RECT 165.400 215.800 165.800 216.600 ;
        RECT 164.600 215.100 164.900 215.800 ;
        RECT 166.200 215.100 166.600 219.900 ;
        RECT 167.800 215.700 168.200 219.900 ;
        RECT 170.000 218.200 170.400 219.900 ;
        RECT 169.400 217.900 170.400 218.200 ;
        RECT 172.200 217.900 172.600 219.900 ;
        RECT 174.300 217.900 174.900 219.900 ;
        RECT 169.400 217.500 169.800 217.900 ;
        RECT 172.200 217.600 172.500 217.900 ;
        RECT 171.100 217.300 172.900 217.600 ;
        RECT 174.200 217.500 174.600 217.900 ;
        RECT 171.100 217.200 171.500 217.300 ;
        RECT 172.500 217.200 172.900 217.300 ;
        RECT 169.400 216.500 169.800 216.600 ;
        RECT 171.700 216.500 172.100 216.600 ;
        RECT 169.400 216.200 172.100 216.500 ;
        RECT 172.400 216.500 173.500 216.800 ;
        RECT 172.400 215.900 172.700 216.500 ;
        RECT 173.100 216.400 173.500 216.500 ;
        RECT 174.300 216.600 175.000 217.000 ;
        RECT 174.300 216.100 174.600 216.600 ;
        RECT 170.300 215.700 172.700 215.900 ;
        RECT 167.800 215.600 172.700 215.700 ;
        RECT 173.400 215.800 174.600 216.100 ;
        RECT 167.800 215.500 170.700 215.600 ;
        RECT 167.800 215.400 170.600 215.500 ;
        RECT 171.000 215.100 171.400 215.200 ;
        RECT 164.600 214.800 166.600 215.100 ;
        RECT 161.400 213.400 161.800 214.200 ;
        RECT 162.200 214.100 162.600 214.200 ;
        RECT 163.700 214.100 165.000 214.200 ;
        RECT 165.400 214.100 165.800 214.200 ;
        RECT 162.200 213.800 163.000 214.100 ;
        RECT 163.700 213.800 165.800 214.100 ;
        RECT 162.600 213.600 163.000 213.800 ;
        RECT 162.300 213.100 164.100 213.300 ;
        RECT 164.600 213.100 164.900 213.800 ;
        RECT 166.200 213.100 166.600 214.800 ;
        RECT 168.900 214.800 171.400 215.100 ;
        RECT 168.900 214.700 169.300 214.800 ;
        RECT 170.200 214.700 170.600 214.800 ;
        RECT 169.700 214.200 170.100 214.300 ;
        RECT 173.400 214.200 173.700 215.800 ;
        RECT 176.600 215.600 177.000 219.900 ;
        RECT 178.200 216.400 178.600 219.900 ;
        RECT 174.900 215.300 177.000 215.600 ;
        RECT 174.900 215.200 175.300 215.300 ;
        RECT 175.700 214.900 176.100 215.000 ;
        RECT 174.200 214.600 176.100 214.900 ;
        RECT 174.200 214.500 174.600 214.600 ;
        RECT 167.000 213.400 167.400 214.200 ;
        RECT 168.200 213.900 173.700 214.200 ;
        RECT 168.200 213.800 169.000 213.900 ;
        RECT 156.600 213.000 158.600 213.100 ;
        RECT 156.600 211.100 157.000 213.000 ;
        RECT 158.200 211.100 158.600 213.000 ;
        RECT 159.000 211.100 159.400 213.100 ;
        RECT 160.100 212.800 161.000 213.100 ;
        RECT 162.200 213.000 164.200 213.100 ;
        RECT 160.100 211.100 160.500 212.800 ;
        RECT 162.200 211.100 162.600 213.000 ;
        RECT 163.800 211.100 164.200 213.000 ;
        RECT 164.600 211.100 165.000 213.100 ;
        RECT 165.700 212.800 166.600 213.100 ;
        RECT 165.700 211.100 166.100 212.800 ;
        RECT 167.800 211.100 168.200 213.500 ;
        RECT 170.300 212.800 170.600 213.900 ;
        RECT 173.100 213.800 173.500 213.900 ;
        RECT 176.600 213.600 177.000 215.300 ;
        RECT 175.100 213.300 177.000 213.600 ;
        RECT 175.100 213.200 175.500 213.300 ;
        RECT 169.400 212.100 169.800 212.500 ;
        RECT 170.200 212.400 170.600 212.800 ;
        RECT 171.100 212.700 171.500 212.800 ;
        RECT 171.100 212.400 172.500 212.700 ;
        RECT 172.200 212.100 172.500 212.400 ;
        RECT 174.200 212.100 174.600 212.500 ;
        RECT 169.400 211.800 170.400 212.100 ;
        RECT 170.000 211.100 170.400 211.800 ;
        RECT 172.200 211.100 172.600 212.100 ;
        RECT 174.200 211.800 174.900 212.100 ;
        RECT 174.300 211.100 174.900 211.800 ;
        RECT 176.600 211.100 177.000 213.300 ;
        RECT 178.100 215.900 178.600 216.400 ;
        RECT 179.800 216.200 180.200 219.900 ;
        RECT 178.900 215.900 180.200 216.200 ;
        RECT 178.100 214.200 178.400 215.900 ;
        RECT 178.900 214.900 179.200 215.900 ;
        RECT 178.700 214.500 179.200 214.900 ;
        RECT 178.100 213.800 178.600 214.200 ;
        RECT 178.100 213.100 178.400 213.800 ;
        RECT 178.900 213.700 179.200 214.500 ;
        RECT 179.700 214.800 180.200 215.200 ;
        RECT 179.700 214.400 180.100 214.800 ;
        RECT 178.900 213.400 180.200 213.700 ;
        RECT 178.100 212.800 178.600 213.100 ;
        RECT 178.200 211.100 178.600 212.800 ;
        RECT 179.800 211.100 180.200 213.400 ;
        RECT 181.400 213.100 181.800 219.900 ;
        RECT 183.000 217.100 183.400 219.900 ;
        RECT 185.100 217.900 185.700 219.900 ;
        RECT 187.400 217.900 187.800 219.900 ;
        RECT 189.600 218.200 190.000 219.900 ;
        RECT 189.600 217.900 190.600 218.200 ;
        RECT 185.400 217.500 185.800 217.900 ;
        RECT 187.500 217.600 187.800 217.900 ;
        RECT 187.100 217.300 188.900 217.600 ;
        RECT 190.200 217.500 190.600 217.900 ;
        RECT 187.100 217.200 187.500 217.300 ;
        RECT 188.500 217.200 188.900 217.300 ;
        RECT 182.200 216.800 183.400 217.100 ;
        RECT 182.200 215.800 182.600 216.800 ;
        RECT 183.000 215.600 183.400 216.800 ;
        RECT 185.000 216.600 185.700 217.000 ;
        RECT 185.400 216.100 185.700 216.600 ;
        RECT 186.500 216.500 187.600 216.800 ;
        RECT 186.500 216.400 186.900 216.500 ;
        RECT 185.400 215.800 186.600 216.100 ;
        RECT 183.000 215.300 185.100 215.600 ;
        RECT 183.000 213.600 183.400 215.300 ;
        RECT 184.700 215.200 185.100 215.300 ;
        RECT 183.900 214.900 184.300 215.000 ;
        RECT 183.900 214.600 185.800 214.900 ;
        RECT 185.400 214.500 185.800 214.600 ;
        RECT 186.300 214.200 186.600 215.800 ;
        RECT 187.300 215.900 187.600 216.500 ;
        RECT 187.900 216.500 188.300 216.600 ;
        RECT 190.200 216.500 190.600 216.600 ;
        RECT 187.900 216.200 190.600 216.500 ;
        RECT 187.300 215.700 189.700 215.900 ;
        RECT 191.800 215.700 192.200 219.900 ;
        RECT 187.300 215.600 192.200 215.700 ;
        RECT 189.300 215.500 192.200 215.600 ;
        RECT 189.400 215.400 192.200 215.500 ;
        RECT 193.400 215.600 193.800 219.900 ;
        RECT 195.000 215.600 195.400 219.900 ;
        RECT 196.600 215.600 197.000 219.900 ;
        RECT 198.200 215.600 198.600 219.900 ;
        RECT 199.800 216.200 200.200 219.900 ;
        RECT 201.400 216.400 201.800 219.900 ;
        RECT 199.800 215.900 201.100 216.200 ;
        RECT 201.400 215.900 201.900 216.400 ;
        RECT 205.900 216.200 206.300 219.900 ;
        RECT 206.600 216.800 207.000 217.200 ;
        RECT 206.700 216.200 207.000 216.800 ;
        RECT 205.900 215.900 206.400 216.200 ;
        RECT 206.700 215.900 207.400 216.200 ;
        RECT 193.400 215.200 194.300 215.600 ;
        RECT 195.000 215.200 196.100 215.600 ;
        RECT 196.600 215.200 197.700 215.600 ;
        RECT 198.200 215.200 199.400 215.600 ;
        RECT 187.800 215.100 188.200 215.200 ;
        RECT 188.600 215.100 189.000 215.200 ;
        RECT 187.800 214.800 191.100 215.100 ;
        RECT 190.700 214.700 191.100 214.800 ;
        RECT 193.900 214.500 194.300 215.200 ;
        RECT 195.700 214.500 196.100 215.200 ;
        RECT 197.300 214.500 197.700 215.200 ;
        RECT 189.900 214.200 190.300 214.300 ;
        RECT 186.300 213.900 191.800 214.200 ;
        RECT 186.500 213.800 186.900 213.900 ;
        RECT 188.600 213.800 189.000 213.900 ;
        RECT 183.000 213.300 184.900 213.600 ;
        RECT 181.400 212.800 182.300 213.100 ;
        RECT 181.900 212.200 182.300 212.800 ;
        RECT 181.900 211.800 182.600 212.200 ;
        RECT 181.900 211.100 182.300 211.800 ;
        RECT 183.000 211.100 183.400 213.300 ;
        RECT 184.500 213.200 184.900 213.300 ;
        RECT 189.400 212.800 189.700 213.900 ;
        RECT 191.000 213.800 191.800 213.900 ;
        RECT 193.900 214.100 195.200 214.500 ;
        RECT 195.700 214.100 196.900 214.500 ;
        RECT 197.300 214.100 198.600 214.500 ;
        RECT 193.900 213.800 194.300 214.100 ;
        RECT 195.700 213.800 196.100 214.100 ;
        RECT 197.300 213.800 197.700 214.100 ;
        RECT 199.000 213.800 199.400 215.200 ;
        RECT 199.800 214.800 200.300 215.200 ;
        RECT 199.900 214.400 200.300 214.800 ;
        RECT 200.800 214.900 201.100 215.900 ;
        RECT 200.800 214.500 201.300 214.900 ;
        RECT 188.500 212.700 188.900 212.800 ;
        RECT 185.400 212.100 185.800 212.500 ;
        RECT 187.500 212.400 188.900 212.700 ;
        RECT 189.400 212.400 189.800 212.800 ;
        RECT 187.500 212.100 187.800 212.400 ;
        RECT 190.200 212.100 190.600 212.500 ;
        RECT 185.100 211.800 185.800 212.100 ;
        RECT 185.100 211.100 185.700 211.800 ;
        RECT 187.400 211.100 187.800 212.100 ;
        RECT 189.600 211.800 190.600 212.100 ;
        RECT 189.600 211.100 190.000 211.800 ;
        RECT 191.800 211.100 192.200 213.500 ;
        RECT 193.400 213.400 194.300 213.800 ;
        RECT 195.000 213.400 196.100 213.800 ;
        RECT 196.600 213.400 197.700 213.800 ;
        RECT 198.200 213.400 199.400 213.800 ;
        RECT 200.800 213.700 201.100 214.500 ;
        RECT 201.600 214.200 201.900 215.900 ;
        RECT 201.400 214.100 201.900 214.200 ;
        RECT 204.600 214.800 205.000 215.200 ;
        RECT 204.600 214.200 204.900 214.800 ;
        RECT 205.400 214.400 205.800 215.200 ;
        RECT 206.100 214.200 206.400 215.900 ;
        RECT 207.000 215.800 207.400 215.900 ;
        RECT 207.800 215.800 208.200 216.600 ;
        RECT 207.000 215.100 207.300 215.800 ;
        RECT 208.600 215.100 209.000 219.900 ;
        RECT 211.000 215.600 211.400 219.900 ;
        RECT 212.600 215.600 213.000 219.900 ;
        RECT 214.200 215.600 214.600 219.900 ;
        RECT 215.800 215.600 216.200 219.900 ;
        RECT 217.400 215.800 217.800 216.600 ;
        RECT 218.200 216.100 218.600 219.900 ;
        RECT 220.200 216.800 220.600 217.200 ;
        RECT 220.200 216.200 220.500 216.800 ;
        RECT 220.900 216.200 221.300 219.900 ;
        RECT 219.800 216.100 220.500 216.200 ;
        RECT 218.200 215.900 220.500 216.100 ;
        RECT 218.200 215.800 220.200 215.900 ;
        RECT 220.800 215.800 221.800 216.200 ;
        RECT 211.000 215.200 211.900 215.600 ;
        RECT 212.600 215.200 213.700 215.600 ;
        RECT 214.200 215.200 215.300 215.600 ;
        RECT 215.800 215.200 217.000 215.600 ;
        RECT 207.000 214.800 209.000 215.100 ;
        RECT 204.600 214.100 205.000 214.200 ;
        RECT 206.100 214.100 207.400 214.200 ;
        RECT 207.800 214.100 208.200 214.200 ;
        RECT 201.400 213.800 205.400 214.100 ;
        RECT 206.100 213.800 208.200 214.100 ;
        RECT 199.800 213.400 201.100 213.700 ;
        RECT 193.400 211.100 193.800 213.400 ;
        RECT 195.000 211.100 195.400 213.400 ;
        RECT 196.600 211.100 197.000 213.400 ;
        RECT 198.200 211.100 198.600 213.400 ;
        RECT 199.800 211.100 200.200 213.400 ;
        RECT 201.600 213.100 201.900 213.800 ;
        RECT 205.000 213.600 205.400 213.800 ;
        RECT 204.700 213.100 206.500 213.300 ;
        RECT 207.000 213.100 207.300 213.800 ;
        RECT 208.600 213.100 209.000 214.800 ;
        RECT 211.500 214.500 211.900 215.200 ;
        RECT 213.300 214.500 213.700 215.200 ;
        RECT 214.900 214.500 215.300 215.200 ;
        RECT 209.400 213.400 209.800 214.200 ;
        RECT 210.200 214.100 211.100 214.500 ;
        RECT 211.500 214.100 212.800 214.500 ;
        RECT 213.300 214.100 214.500 214.500 ;
        RECT 214.900 214.100 216.200 214.500 ;
        RECT 210.200 213.800 210.600 214.100 ;
        RECT 211.500 213.800 211.900 214.100 ;
        RECT 213.300 213.800 213.700 214.100 ;
        RECT 214.900 213.800 215.300 214.100 ;
        RECT 216.600 213.800 217.000 215.200 ;
        RECT 211.000 213.400 211.900 213.800 ;
        RECT 212.600 213.400 213.700 213.800 ;
        RECT 214.200 213.400 215.300 213.800 ;
        RECT 215.800 213.400 217.000 213.800 ;
        RECT 201.400 212.800 201.900 213.100 ;
        RECT 204.600 213.000 206.600 213.100 ;
        RECT 201.400 211.100 201.800 212.800 ;
        RECT 204.600 211.100 205.000 213.000 ;
        RECT 206.200 211.100 206.600 213.000 ;
        RECT 207.000 211.100 207.400 213.100 ;
        RECT 208.100 212.800 209.000 213.100 ;
        RECT 208.100 211.100 208.500 212.800 ;
        RECT 211.000 211.100 211.400 213.400 ;
        RECT 212.600 211.100 213.000 213.400 ;
        RECT 214.200 211.100 214.600 213.400 ;
        RECT 215.800 211.100 216.200 213.400 ;
        RECT 218.200 213.100 218.600 215.800 ;
        RECT 220.800 214.200 221.100 215.800 ;
        RECT 223.000 215.700 223.400 219.900 ;
        RECT 225.200 218.200 225.600 219.900 ;
        RECT 224.600 217.900 225.600 218.200 ;
        RECT 227.400 217.900 227.800 219.900 ;
        RECT 229.500 217.900 230.100 219.900 ;
        RECT 224.600 217.500 225.000 217.900 ;
        RECT 227.400 217.600 227.700 217.900 ;
        RECT 226.300 217.300 228.100 217.600 ;
        RECT 229.400 217.500 229.800 217.900 ;
        RECT 226.300 217.200 226.700 217.300 ;
        RECT 227.700 217.200 228.100 217.300 ;
        RECT 224.600 216.500 225.000 216.600 ;
        RECT 226.900 216.500 227.300 216.600 ;
        RECT 224.600 216.200 227.300 216.500 ;
        RECT 227.600 216.500 228.700 216.800 ;
        RECT 227.600 215.900 227.900 216.500 ;
        RECT 228.300 216.400 228.700 216.500 ;
        RECT 229.500 216.600 230.200 217.000 ;
        RECT 229.500 216.100 229.800 216.600 ;
        RECT 225.500 215.700 227.900 215.900 ;
        RECT 223.000 215.600 227.900 215.700 ;
        RECT 228.600 215.800 229.800 216.100 ;
        RECT 223.000 215.500 225.900 215.600 ;
        RECT 223.000 215.400 225.800 215.500 ;
        RECT 221.400 214.400 221.800 215.200 ;
        RECT 226.200 215.100 226.600 215.200 ;
        RECT 224.100 214.800 226.600 215.100 ;
        RECT 224.100 214.700 224.500 214.800 ;
        RECT 225.400 214.700 225.800 214.800 ;
        RECT 224.900 214.200 225.300 214.300 ;
        RECT 228.600 214.200 228.900 215.800 ;
        RECT 231.800 215.600 232.200 219.900 ;
        RECT 233.000 216.800 233.400 217.200 ;
        RECT 233.000 216.200 233.300 216.800 ;
        RECT 233.700 216.200 234.100 219.900 ;
        RECT 232.600 215.900 233.300 216.200 ;
        RECT 233.600 215.900 234.100 216.200 ;
        RECT 232.600 215.800 233.000 215.900 ;
        RECT 230.100 215.300 232.200 215.600 ;
        RECT 230.100 215.200 230.500 215.300 ;
        RECT 230.900 214.900 231.300 215.000 ;
        RECT 229.400 214.600 231.300 214.900 ;
        RECT 229.400 214.500 229.800 214.600 ;
        RECT 219.000 213.400 219.400 214.200 ;
        RECT 219.800 213.800 221.100 214.200 ;
        RECT 222.200 214.100 222.600 214.200 ;
        RECT 221.800 213.800 222.600 214.100 ;
        RECT 223.400 213.900 228.900 214.200 ;
        RECT 223.400 213.800 224.200 213.900 ;
        RECT 219.900 213.100 220.200 213.800 ;
        RECT 221.800 213.600 222.200 213.800 ;
        RECT 220.700 213.100 222.500 213.300 ;
        RECT 217.700 212.800 218.600 213.100 ;
        RECT 217.700 211.100 218.100 212.800 ;
        RECT 219.800 211.100 220.200 213.100 ;
        RECT 220.600 213.000 222.600 213.100 ;
        RECT 220.600 211.100 221.000 213.000 ;
        RECT 222.200 211.100 222.600 213.000 ;
        RECT 223.000 211.100 223.400 213.500 ;
        RECT 225.500 212.800 225.800 213.900 ;
        RECT 228.300 213.800 228.700 213.900 ;
        RECT 231.800 213.600 232.200 215.300 ;
        RECT 233.600 214.200 233.900 215.900 ;
        RECT 234.200 214.400 234.600 215.200 ;
        RECT 236.600 215.100 237.000 219.900 ;
        RECT 239.300 219.200 239.700 219.900 ;
        RECT 239.300 218.800 240.200 219.200 ;
        RECT 238.600 216.800 239.000 217.200 ;
        RECT 237.400 215.800 237.800 216.600 ;
        RECT 238.600 216.200 238.900 216.800 ;
        RECT 239.300 216.200 239.700 218.800 ;
        RECT 238.200 215.900 238.900 216.200 ;
        RECT 239.200 215.900 239.700 216.200 ;
        RECT 238.200 215.800 238.600 215.900 ;
        RECT 238.200 215.100 238.500 215.800 ;
        RECT 236.600 214.800 238.500 215.100 ;
        RECT 232.600 213.800 233.900 214.200 ;
        RECT 235.000 214.100 235.400 214.200 ;
        RECT 234.600 213.800 235.400 214.100 ;
        RECT 230.300 213.300 232.200 213.600 ;
        RECT 230.300 213.200 230.700 213.300 ;
        RECT 224.600 212.100 225.000 212.500 ;
        RECT 225.400 212.400 225.800 212.800 ;
        RECT 226.300 212.700 226.700 212.800 ;
        RECT 226.300 212.400 227.700 212.700 ;
        RECT 227.400 212.100 227.700 212.400 ;
        RECT 229.400 212.100 229.800 212.500 ;
        RECT 224.600 211.800 225.600 212.100 ;
        RECT 225.200 211.100 225.600 211.800 ;
        RECT 227.400 211.100 227.800 212.100 ;
        RECT 229.400 211.800 230.100 212.100 ;
        RECT 229.500 211.100 230.100 211.800 ;
        RECT 231.800 211.100 232.200 213.300 ;
        RECT 232.700 213.100 233.000 213.800 ;
        RECT 234.600 213.600 235.000 213.800 ;
        RECT 235.800 213.400 236.200 214.200 ;
        RECT 233.500 213.100 235.300 213.300 ;
        RECT 236.600 213.100 237.000 214.800 ;
        RECT 239.200 214.200 239.500 215.900 ;
        RECT 241.400 215.600 241.800 219.900 ;
        RECT 243.500 217.900 244.100 219.900 ;
        RECT 245.800 217.900 246.200 219.900 ;
        RECT 248.000 218.200 248.400 219.900 ;
        RECT 248.000 217.900 249.000 218.200 ;
        RECT 243.800 217.500 244.200 217.900 ;
        RECT 245.900 217.600 246.200 217.900 ;
        RECT 245.500 217.300 247.300 217.600 ;
        RECT 248.600 217.500 249.000 217.900 ;
        RECT 245.500 217.200 245.900 217.300 ;
        RECT 246.900 217.200 247.300 217.300 ;
        RECT 243.400 216.600 244.100 217.000 ;
        RECT 243.800 216.100 244.100 216.600 ;
        RECT 244.900 216.500 246.000 216.800 ;
        RECT 244.900 216.400 245.300 216.500 ;
        RECT 243.800 215.800 245.000 216.100 ;
        RECT 241.400 215.300 243.500 215.600 ;
        RECT 239.800 214.400 240.200 215.200 ;
        RECT 238.200 213.800 239.500 214.200 ;
        RECT 240.600 214.100 241.000 214.200 ;
        RECT 240.200 213.800 241.000 214.100 ;
        RECT 238.300 213.100 238.600 213.800 ;
        RECT 240.200 213.600 240.600 213.800 ;
        RECT 241.400 213.600 241.800 215.300 ;
        RECT 243.100 215.200 243.500 215.300 ;
        RECT 244.700 215.200 245.000 215.800 ;
        RECT 245.700 215.900 246.000 216.500 ;
        RECT 246.300 216.500 246.700 216.600 ;
        RECT 248.600 216.500 249.000 216.600 ;
        RECT 246.300 216.200 249.000 216.500 ;
        RECT 245.700 215.700 248.100 215.900 ;
        RECT 250.200 215.700 250.600 219.900 ;
        RECT 245.700 215.600 250.600 215.700 ;
        RECT 247.700 215.500 250.600 215.600 ;
        RECT 247.800 215.400 250.600 215.500 ;
        RECT 242.300 214.900 242.700 215.000 ;
        RECT 242.300 214.600 244.200 214.900 ;
        RECT 244.600 214.800 245.000 215.200 ;
        RECT 247.000 215.100 247.400 215.200 ;
        RECT 247.000 214.800 249.500 215.100 ;
        RECT 243.800 214.500 244.200 214.600 ;
        RECT 244.700 214.200 245.000 214.800 ;
        RECT 247.800 214.700 248.200 214.800 ;
        RECT 249.100 214.700 249.500 214.800 ;
        RECT 248.300 214.200 248.700 214.300 ;
        RECT 244.700 213.900 250.200 214.200 ;
        RECT 244.900 213.800 245.300 213.900 ;
        RECT 241.400 213.300 243.300 213.600 ;
        RECT 239.100 213.100 240.900 213.300 ;
        RECT 232.600 211.100 233.000 213.100 ;
        RECT 233.400 213.000 235.400 213.100 ;
        RECT 233.400 211.100 233.800 213.000 ;
        RECT 235.000 211.100 235.400 213.000 ;
        RECT 236.600 212.800 237.500 213.100 ;
        RECT 237.100 211.100 237.500 212.800 ;
        RECT 238.200 211.100 238.600 213.100 ;
        RECT 239.000 213.000 241.000 213.100 ;
        RECT 239.000 211.100 239.400 213.000 ;
        RECT 240.600 211.100 241.000 213.000 ;
        RECT 241.400 211.100 241.800 213.300 ;
        RECT 242.900 213.200 243.300 213.300 ;
        RECT 247.800 212.800 248.100 213.900 ;
        RECT 249.400 213.800 250.200 213.900 ;
        RECT 246.900 212.700 247.300 212.800 ;
        RECT 243.800 212.100 244.200 212.500 ;
        RECT 245.900 212.400 247.300 212.700 ;
        RECT 247.800 212.400 248.200 212.800 ;
        RECT 245.900 212.100 246.200 212.400 ;
        RECT 248.600 212.100 249.000 212.500 ;
        RECT 243.500 211.800 244.200 212.100 ;
        RECT 243.500 211.100 244.100 211.800 ;
        RECT 245.800 211.100 246.200 212.100 ;
        RECT 248.000 211.800 249.000 212.100 ;
        RECT 248.000 211.100 248.400 211.800 ;
        RECT 250.200 211.100 250.600 213.500 ;
        RECT 0.600 207.700 1.000 209.900 ;
        RECT 2.700 209.200 3.300 209.900 ;
        RECT 2.700 208.900 3.400 209.200 ;
        RECT 5.000 208.900 5.400 209.900 ;
        RECT 7.200 209.200 7.600 209.900 ;
        RECT 7.200 208.900 8.200 209.200 ;
        RECT 3.000 208.500 3.400 208.900 ;
        RECT 5.100 208.600 5.400 208.900 ;
        RECT 5.100 208.300 6.500 208.600 ;
        RECT 6.100 208.200 6.500 208.300 ;
        RECT 7.000 208.200 7.400 208.600 ;
        RECT 7.800 208.500 8.200 208.900 ;
        RECT 2.100 207.700 2.500 207.800 ;
        RECT 0.600 207.400 2.500 207.700 ;
        RECT 0.600 205.700 1.000 207.400 ;
        RECT 4.100 207.100 4.500 207.200 ;
        RECT 7.000 207.100 7.300 208.200 ;
        RECT 9.400 207.500 9.800 209.900 ;
        RECT 10.200 208.000 10.600 209.900 ;
        RECT 11.800 208.000 12.200 209.900 ;
        RECT 10.200 207.900 12.200 208.000 ;
        RECT 12.600 207.900 13.000 209.900 ;
        RECT 13.700 208.200 14.100 209.900 ;
        RECT 13.700 207.900 14.600 208.200 ;
        RECT 15.800 208.000 16.200 209.900 ;
        RECT 17.400 208.000 17.800 209.900 ;
        RECT 15.800 207.900 17.800 208.000 ;
        RECT 18.200 207.900 18.600 209.900 ;
        RECT 19.300 208.200 19.700 209.900 ;
        RECT 21.400 208.500 21.800 209.500 ;
        RECT 19.300 207.900 20.200 208.200 ;
        RECT 10.300 207.700 12.100 207.900 ;
        RECT 10.600 207.200 11.000 207.400 ;
        RECT 12.600 207.200 12.900 207.900 ;
        RECT 8.600 207.100 9.400 207.200 ;
        RECT 3.900 206.800 9.400 207.100 ;
        RECT 10.200 206.900 11.000 207.200 ;
        RECT 10.200 206.800 10.600 206.900 ;
        RECT 11.700 206.800 13.000 207.200 ;
        RECT 3.000 206.400 3.400 206.500 ;
        RECT 1.500 206.100 3.400 206.400 ;
        RECT 1.500 206.000 1.900 206.100 ;
        RECT 2.300 205.700 2.700 205.800 ;
        RECT 0.600 205.400 2.700 205.700 ;
        RECT 0.600 201.100 1.000 205.400 ;
        RECT 3.900 205.200 4.200 206.800 ;
        RECT 7.500 206.700 7.900 206.800 ;
        RECT 7.000 206.200 7.400 206.300 ;
        RECT 8.300 206.200 8.700 206.300 ;
        RECT 6.200 205.900 8.700 206.200 ;
        RECT 6.200 205.800 6.600 205.900 ;
        RECT 11.000 205.800 11.400 206.600 ;
        RECT 11.700 206.200 12.000 206.800 ;
        RECT 11.700 205.800 12.200 206.200 ;
        RECT 14.200 206.100 14.600 207.900 ;
        RECT 15.900 207.700 17.700 207.900 ;
        RECT 15.000 206.800 15.400 207.600 ;
        RECT 16.200 207.200 16.600 207.400 ;
        RECT 18.200 207.200 18.500 207.900 ;
        RECT 15.800 206.900 16.600 207.200 ;
        RECT 15.800 206.800 16.200 206.900 ;
        RECT 17.300 206.800 18.600 207.200 ;
        RECT 12.600 205.800 14.600 206.100 ;
        RECT 16.600 205.800 17.000 206.600 ;
        RECT 7.000 205.500 9.800 205.600 ;
        RECT 6.900 205.400 9.800 205.500 ;
        RECT 3.000 204.900 4.200 205.200 ;
        RECT 4.900 205.300 9.800 205.400 ;
        RECT 4.900 205.100 7.300 205.300 ;
        RECT 3.000 204.400 3.300 204.900 ;
        RECT 2.600 204.000 3.300 204.400 ;
        RECT 4.100 204.500 4.500 204.600 ;
        RECT 4.900 204.500 5.200 205.100 ;
        RECT 4.100 204.200 5.200 204.500 ;
        RECT 5.500 204.500 8.200 204.800 ;
        RECT 5.500 204.400 5.900 204.500 ;
        RECT 7.800 204.400 8.200 204.500 ;
        RECT 4.700 203.700 5.100 203.800 ;
        RECT 6.100 203.700 6.500 203.800 ;
        RECT 3.000 203.100 3.400 203.500 ;
        RECT 4.700 203.400 6.500 203.700 ;
        RECT 5.100 203.100 5.400 203.400 ;
        RECT 7.800 203.100 8.200 203.500 ;
        RECT 2.700 201.100 3.300 203.100 ;
        RECT 5.000 201.100 5.400 203.100 ;
        RECT 7.200 202.800 8.200 203.100 ;
        RECT 7.200 201.100 7.600 202.800 ;
        RECT 9.400 201.100 9.800 205.300 ;
        RECT 11.700 205.100 12.000 205.800 ;
        RECT 12.600 205.200 12.900 205.800 ;
        RECT 12.600 205.100 13.000 205.200 ;
        RECT 11.500 204.800 12.000 205.100 ;
        RECT 12.300 204.800 13.000 205.100 ;
        RECT 11.500 201.100 11.900 204.800 ;
        RECT 12.300 204.200 12.600 204.800 ;
        RECT 13.400 204.400 13.800 205.200 ;
        RECT 12.200 203.800 12.600 204.200 ;
        RECT 14.200 201.100 14.600 205.800 ;
        RECT 17.300 205.100 17.600 206.800 ;
        RECT 19.800 206.100 20.200 207.900 ;
        RECT 20.600 206.800 21.000 207.600 ;
        RECT 21.400 207.400 21.700 208.500 ;
        RECT 23.500 208.000 23.900 209.500 ;
        RECT 23.500 207.700 24.300 208.000 ;
        RECT 23.900 207.500 24.300 207.700 ;
        RECT 21.400 207.100 23.500 207.400 ;
        RECT 23.000 206.900 23.500 207.100 ;
        RECT 24.000 207.200 24.300 207.500 ;
        RECT 26.200 207.700 26.600 209.900 ;
        RECT 28.300 209.200 28.900 209.900 ;
        RECT 28.300 208.900 29.000 209.200 ;
        RECT 30.600 208.900 31.000 209.900 ;
        RECT 32.800 209.200 33.200 209.900 ;
        RECT 32.800 208.900 33.800 209.200 ;
        RECT 28.600 208.500 29.000 208.900 ;
        RECT 30.700 208.600 31.000 208.900 ;
        RECT 30.700 208.300 32.100 208.600 ;
        RECT 31.700 208.200 32.100 208.300 ;
        RECT 32.600 208.200 33.000 208.600 ;
        RECT 33.400 208.500 33.800 208.900 ;
        RECT 27.800 207.800 28.200 208.200 ;
        RECT 27.700 207.700 28.200 207.800 ;
        RECT 26.200 207.400 28.200 207.700 ;
        RECT 18.200 205.800 20.200 206.100 ;
        RECT 21.400 205.800 21.800 206.600 ;
        RECT 22.200 205.800 22.600 206.600 ;
        RECT 23.000 206.500 23.700 206.900 ;
        RECT 24.000 206.800 25.000 207.200 ;
        RECT 18.200 205.200 18.500 205.800 ;
        RECT 18.200 205.100 18.600 205.200 ;
        RECT 17.100 204.800 17.600 205.100 ;
        RECT 17.900 204.800 18.600 205.100 ;
        RECT 17.100 201.100 17.500 204.800 ;
        RECT 17.900 204.200 18.200 204.800 ;
        RECT 19.000 204.400 19.400 205.200 ;
        RECT 17.800 203.800 18.200 204.200 ;
        RECT 19.800 201.100 20.200 205.800 ;
        RECT 23.000 205.500 23.300 206.500 ;
        RECT 21.400 205.200 23.300 205.500 ;
        RECT 21.400 203.500 21.700 205.200 ;
        RECT 24.000 204.900 24.300 206.800 ;
        RECT 24.600 206.100 25.000 206.200 ;
        RECT 26.200 206.100 26.600 207.400 ;
        RECT 29.700 207.100 30.100 207.200 ;
        RECT 32.600 207.100 32.900 208.200 ;
        RECT 35.000 207.500 35.400 209.900 ;
        RECT 37.100 208.200 37.500 209.900 ;
        RECT 36.600 207.900 37.500 208.200 ;
        RECT 38.200 207.900 38.600 209.900 ;
        RECT 39.000 208.000 39.400 209.900 ;
        RECT 40.600 208.000 41.000 209.900 ;
        RECT 39.000 207.900 41.000 208.000 ;
        RECT 34.200 207.100 35.000 207.200 ;
        RECT 29.500 206.800 35.000 207.100 ;
        RECT 35.800 206.800 36.200 207.600 ;
        RECT 28.600 206.400 29.000 206.500 ;
        RECT 24.600 205.800 26.600 206.100 ;
        RECT 27.100 206.100 29.000 206.400 ;
        RECT 29.500 206.200 29.800 206.800 ;
        RECT 33.100 206.700 33.500 206.800 ;
        RECT 32.600 206.200 33.000 206.300 ;
        RECT 33.900 206.200 34.300 206.300 ;
        RECT 27.100 206.000 27.500 206.100 ;
        RECT 29.400 205.800 29.800 206.200 ;
        RECT 31.800 205.900 34.300 206.200 ;
        RECT 36.600 206.100 37.000 207.900 ;
        RECT 38.300 207.200 38.600 207.900 ;
        RECT 39.100 207.700 40.900 207.900 ;
        RECT 41.400 207.500 41.800 209.900 ;
        RECT 43.600 209.200 44.000 209.900 ;
        RECT 43.000 208.900 44.000 209.200 ;
        RECT 45.800 208.900 46.200 209.900 ;
        RECT 47.900 209.200 48.500 209.900 ;
        RECT 47.800 208.900 48.500 209.200 ;
        RECT 43.000 208.500 43.400 208.900 ;
        RECT 45.800 208.600 46.100 208.900 ;
        RECT 43.800 208.200 44.200 208.600 ;
        RECT 44.700 208.300 46.100 208.600 ;
        RECT 47.800 208.500 48.200 208.900 ;
        RECT 44.700 208.200 45.100 208.300 ;
        RECT 40.200 207.200 40.600 207.400 ;
        RECT 43.900 207.200 44.200 208.200 ;
        RECT 48.700 207.700 49.100 207.800 ;
        RECT 50.200 207.700 50.600 209.900 ;
        RECT 52.900 208.200 53.300 209.900 ;
        RECT 52.900 207.900 53.800 208.200 ;
        RECT 48.700 207.400 50.600 207.700 ;
        RECT 38.200 206.800 39.500 207.200 ;
        RECT 40.200 206.900 41.000 207.200 ;
        RECT 40.600 206.800 41.000 206.900 ;
        RECT 41.800 207.100 42.600 207.200 ;
        RECT 43.800 207.100 44.200 207.200 ;
        RECT 46.700 207.100 47.100 207.200 ;
        RECT 41.800 206.800 47.300 207.100 ;
        RECT 39.200 206.200 39.500 206.800 ;
        RECT 43.300 206.700 43.700 206.800 ;
        RECT 31.800 205.800 32.200 205.900 ;
        RECT 36.600 205.800 38.500 206.100 ;
        RECT 39.000 205.800 39.500 206.200 ;
        RECT 39.800 206.100 40.200 206.600 ;
        RECT 42.500 206.200 42.900 206.300 ;
        RECT 40.600 206.100 41.000 206.200 ;
        RECT 39.800 205.800 41.000 206.100 ;
        RECT 42.500 205.900 45.000 206.200 ;
        RECT 44.600 205.800 45.000 205.900 ;
        RECT 24.600 205.400 25.000 205.800 ;
        RECT 26.200 205.700 26.600 205.800 ;
        RECT 27.900 205.700 28.300 205.800 ;
        RECT 26.200 205.400 28.300 205.700 ;
        RECT 23.500 204.600 24.300 204.900 ;
        RECT 21.400 201.500 21.800 203.500 ;
        RECT 23.500 202.200 23.900 204.600 ;
        RECT 23.500 201.800 24.200 202.200 ;
        RECT 23.500 201.100 23.900 201.800 ;
        RECT 26.200 201.100 26.600 205.400 ;
        RECT 29.500 205.200 29.800 205.800 ;
        RECT 32.600 205.500 35.400 205.600 ;
        RECT 32.500 205.400 35.400 205.500 ;
        RECT 28.600 204.900 29.800 205.200 ;
        RECT 30.500 205.300 35.400 205.400 ;
        RECT 30.500 205.100 32.900 205.300 ;
        RECT 28.600 204.400 28.900 204.900 ;
        RECT 28.200 204.000 28.900 204.400 ;
        RECT 29.700 204.500 30.100 204.600 ;
        RECT 30.500 204.500 30.800 205.100 ;
        RECT 29.700 204.200 30.800 204.500 ;
        RECT 31.100 204.500 33.800 204.800 ;
        RECT 31.100 204.400 31.500 204.500 ;
        RECT 33.400 204.400 33.800 204.500 ;
        RECT 30.300 203.700 30.700 203.800 ;
        RECT 31.700 203.700 32.100 203.800 ;
        RECT 28.600 203.100 29.000 203.500 ;
        RECT 30.300 203.400 32.100 203.700 ;
        RECT 30.700 203.100 31.000 203.400 ;
        RECT 33.400 203.100 33.800 203.500 ;
        RECT 28.300 201.100 28.900 203.100 ;
        RECT 30.600 201.100 31.000 203.100 ;
        RECT 32.800 202.800 33.800 203.100 ;
        RECT 32.800 201.100 33.200 202.800 ;
        RECT 35.000 201.100 35.400 205.300 ;
        RECT 36.600 201.100 37.000 205.800 ;
        RECT 38.200 205.200 38.500 205.800 ;
        RECT 37.400 204.400 37.800 205.200 ;
        RECT 38.200 205.100 38.600 205.200 ;
        RECT 39.200 205.100 39.500 205.800 ;
        RECT 41.400 205.500 44.200 205.600 ;
        RECT 41.400 205.400 44.300 205.500 ;
        RECT 41.400 205.300 46.300 205.400 ;
        RECT 38.200 204.800 38.900 205.100 ;
        RECT 39.200 204.800 39.700 205.100 ;
        RECT 38.600 204.200 38.900 204.800 ;
        RECT 38.600 203.800 39.000 204.200 ;
        RECT 39.300 201.100 39.700 204.800 ;
        RECT 41.400 201.100 41.800 205.300 ;
        RECT 43.900 205.100 46.300 205.300 ;
        RECT 43.000 204.500 45.700 204.800 ;
        RECT 43.000 204.400 43.400 204.500 ;
        RECT 45.300 204.400 45.700 204.500 ;
        RECT 46.000 204.500 46.300 205.100 ;
        RECT 47.000 205.200 47.300 206.800 ;
        RECT 47.800 206.400 48.200 206.500 ;
        RECT 47.800 206.100 49.700 206.400 ;
        RECT 49.300 206.000 49.700 206.100 ;
        RECT 48.500 205.700 48.900 205.800 ;
        RECT 50.200 205.700 50.600 207.400 ;
        RECT 48.500 205.400 50.600 205.700 ;
        RECT 47.000 204.900 48.200 205.200 ;
        RECT 46.700 204.500 47.100 204.600 ;
        RECT 46.000 204.200 47.100 204.500 ;
        RECT 47.900 204.400 48.200 204.900 ;
        RECT 47.900 204.000 48.600 204.400 ;
        RECT 44.700 203.700 45.100 203.800 ;
        RECT 46.100 203.700 46.500 203.800 ;
        RECT 43.000 203.100 43.400 203.500 ;
        RECT 44.700 203.400 46.500 203.700 ;
        RECT 45.800 203.100 46.100 203.400 ;
        RECT 47.800 203.100 48.200 203.500 ;
        RECT 43.000 202.800 44.000 203.100 ;
        RECT 43.600 201.100 44.000 202.800 ;
        RECT 45.800 201.100 46.200 203.100 ;
        RECT 47.900 201.100 48.500 203.100 ;
        RECT 50.200 201.100 50.600 205.400 ;
        RECT 53.400 206.100 53.800 207.900 ;
        RECT 56.600 207.900 57.000 209.900 ;
        RECT 57.300 208.200 57.700 208.600 ;
        RECT 55.800 206.400 56.200 207.200 ;
        RECT 55.000 206.100 55.400 206.200 ;
        RECT 56.600 206.100 56.900 207.900 ;
        RECT 57.400 207.800 57.800 208.200 ;
        RECT 60.100 208.000 60.500 209.500 ;
        RECT 62.200 208.500 62.600 209.500 ;
        RECT 59.700 207.700 60.500 208.000 ;
        RECT 59.700 207.500 60.100 207.700 ;
        RECT 59.700 207.200 60.000 207.500 ;
        RECT 62.300 207.400 62.600 208.500 ;
        RECT 64.300 209.200 64.700 209.900 ;
        RECT 64.300 208.800 65.000 209.200 ;
        RECT 64.300 208.200 64.700 208.800 ;
        RECT 63.800 207.900 64.700 208.200 ;
        RECT 59.000 206.800 60.000 207.200 ;
        RECT 60.500 207.100 62.600 207.400 ;
        RECT 60.500 206.900 61.000 207.100 ;
        RECT 57.400 206.100 57.800 206.200 ;
        RECT 53.400 205.800 55.800 206.100 ;
        RECT 56.600 205.800 57.800 206.100 ;
        RECT 58.200 206.100 58.600 206.200 ;
        RECT 59.000 206.100 59.400 206.200 ;
        RECT 58.200 205.800 59.400 206.100 ;
        RECT 51.000 205.100 51.400 205.200 ;
        RECT 52.600 205.100 53.000 205.200 ;
        RECT 51.000 204.800 53.000 205.100 ;
        RECT 52.600 204.400 53.000 204.800 ;
        RECT 53.400 201.100 53.800 205.800 ;
        RECT 55.400 205.600 55.800 205.800 ;
        RECT 57.400 205.100 57.700 205.800 ;
        RECT 59.000 205.400 59.400 205.800 ;
        RECT 55.000 204.800 57.000 205.100 ;
        RECT 55.000 201.100 55.400 204.800 ;
        RECT 56.600 201.100 57.000 204.800 ;
        RECT 57.400 201.100 57.800 205.100 ;
        RECT 59.700 204.900 60.000 206.800 ;
        RECT 60.300 206.500 61.000 206.900 ;
        RECT 63.000 206.800 63.400 207.600 ;
        RECT 60.700 205.500 61.000 206.500 ;
        RECT 61.400 205.800 61.800 206.600 ;
        RECT 62.200 205.800 62.600 206.600 ;
        RECT 60.700 205.200 62.600 205.500 ;
        RECT 59.700 204.600 60.500 204.900 ;
        RECT 60.100 202.200 60.500 204.600 ;
        RECT 62.300 203.500 62.600 205.200 ;
        RECT 60.100 201.800 61.000 202.200 ;
        RECT 60.100 201.100 60.500 201.800 ;
        RECT 62.200 201.500 62.600 203.500 ;
        RECT 63.800 201.100 64.200 207.900 ;
        RECT 65.400 207.700 65.800 209.900 ;
        RECT 67.500 209.200 68.100 209.900 ;
        RECT 67.500 208.900 68.200 209.200 ;
        RECT 69.800 208.900 70.200 209.900 ;
        RECT 72.000 209.200 72.400 209.900 ;
        RECT 72.000 208.900 73.000 209.200 ;
        RECT 67.800 208.500 68.200 208.900 ;
        RECT 69.900 208.600 70.200 208.900 ;
        RECT 69.900 208.300 71.300 208.600 ;
        RECT 70.900 208.200 71.300 208.300 ;
        RECT 71.800 208.200 72.200 208.600 ;
        RECT 72.600 208.500 73.000 208.900 ;
        RECT 66.900 207.700 67.300 207.800 ;
        RECT 65.400 207.400 67.300 207.700 ;
        RECT 65.400 205.700 65.800 207.400 ;
        RECT 68.900 207.100 69.300 207.200 ;
        RECT 71.800 207.100 72.100 208.200 ;
        RECT 74.200 207.500 74.600 209.900 ;
        RECT 75.800 208.800 76.200 209.900 ;
        RECT 75.000 207.800 75.400 208.600 ;
        RECT 75.000 207.200 75.300 207.800 ;
        RECT 75.900 207.200 76.200 208.800 ;
        RECT 78.700 208.200 79.100 209.900 ;
        RECT 78.200 207.900 79.100 208.200 ;
        RECT 73.400 207.100 74.200 207.200 ;
        RECT 68.700 206.800 74.200 207.100 ;
        RECT 75.000 206.800 75.400 207.200 ;
        RECT 75.800 206.800 76.200 207.200 ;
        RECT 77.400 206.800 77.800 207.600 ;
        RECT 67.800 206.400 68.200 206.500 ;
        RECT 66.300 206.100 68.200 206.400 ;
        RECT 68.700 206.200 69.000 206.800 ;
        RECT 72.300 206.700 72.700 206.800 ;
        RECT 71.800 206.200 72.200 206.300 ;
        RECT 73.100 206.200 73.500 206.300 ;
        RECT 66.300 206.000 66.700 206.100 ;
        RECT 68.600 205.800 69.000 206.200 ;
        RECT 71.000 205.900 73.500 206.200 ;
        RECT 71.000 205.800 71.400 205.900 ;
        RECT 67.100 205.700 67.500 205.800 ;
        RECT 65.400 205.400 67.500 205.700 ;
        RECT 64.600 204.400 65.000 205.200 ;
        RECT 65.400 201.100 65.800 205.400 ;
        RECT 67.000 204.800 67.400 205.400 ;
        RECT 68.700 205.200 69.000 205.800 ;
        RECT 71.800 205.500 74.600 205.600 ;
        RECT 71.700 205.400 74.600 205.500 ;
        RECT 67.800 204.900 69.000 205.200 ;
        RECT 69.700 205.300 74.600 205.400 ;
        RECT 69.700 205.100 72.100 205.300 ;
        RECT 67.800 204.400 68.100 204.900 ;
        RECT 67.400 204.000 68.100 204.400 ;
        RECT 68.900 204.500 69.300 204.600 ;
        RECT 69.700 204.500 70.000 205.100 ;
        RECT 68.900 204.200 70.000 204.500 ;
        RECT 70.300 204.500 73.000 204.800 ;
        RECT 70.300 204.400 70.700 204.500 ;
        RECT 72.600 204.400 73.000 204.500 ;
        RECT 69.500 203.700 69.900 203.800 ;
        RECT 70.900 203.700 71.300 203.800 ;
        RECT 67.800 203.100 68.200 203.500 ;
        RECT 69.500 203.400 71.300 203.700 ;
        RECT 69.900 203.100 70.200 203.400 ;
        RECT 72.600 203.100 73.000 203.500 ;
        RECT 67.500 201.100 68.100 203.100 ;
        RECT 69.800 201.100 70.200 203.100 ;
        RECT 72.000 202.800 73.000 203.100 ;
        RECT 72.000 201.100 72.400 202.800 ;
        RECT 74.200 201.100 74.600 205.300 ;
        RECT 75.900 205.100 76.200 206.800 ;
        RECT 76.600 205.400 77.000 206.200 ;
        RECT 75.800 204.700 76.700 205.100 ;
        RECT 76.300 201.100 76.700 204.700 ;
        RECT 78.200 201.100 78.600 207.900 ;
        RECT 79.800 207.500 80.200 209.900 ;
        RECT 82.000 209.200 82.400 209.900 ;
        RECT 81.400 208.900 82.400 209.200 ;
        RECT 84.200 208.900 84.600 209.900 ;
        RECT 86.300 209.200 86.900 209.900 ;
        RECT 86.200 208.900 86.900 209.200 ;
        RECT 81.400 208.500 81.800 208.900 ;
        RECT 84.200 208.600 84.500 208.900 ;
        RECT 82.200 208.200 82.600 208.600 ;
        RECT 83.100 208.300 84.500 208.600 ;
        RECT 86.200 208.500 86.600 208.900 ;
        RECT 83.100 208.200 83.500 208.300 ;
        RECT 80.200 207.100 81.000 207.200 ;
        RECT 82.300 207.100 82.600 208.200 ;
        RECT 87.100 207.700 87.500 207.800 ;
        RECT 88.600 207.700 89.000 209.900 ;
        RECT 87.100 207.400 89.000 207.700 ;
        RECT 83.000 207.100 83.400 207.200 ;
        RECT 85.100 207.100 85.500 207.200 ;
        RECT 80.200 206.800 85.700 207.100 ;
        RECT 81.700 206.700 82.100 206.800 ;
        RECT 80.900 206.200 81.300 206.300 ;
        RECT 82.200 206.200 82.600 206.300 ;
        RECT 80.900 205.900 83.400 206.200 ;
        RECT 83.000 205.800 83.400 205.900 ;
        RECT 79.800 205.500 82.600 205.600 ;
        RECT 79.800 205.400 82.700 205.500 ;
        RECT 79.800 205.300 84.700 205.400 ;
        RECT 79.000 204.400 79.400 205.200 ;
        RECT 79.800 201.100 80.200 205.300 ;
        RECT 82.300 205.100 84.700 205.300 ;
        RECT 81.400 204.500 84.100 204.800 ;
        RECT 81.400 204.400 81.800 204.500 ;
        RECT 83.700 204.400 84.100 204.500 ;
        RECT 84.400 204.500 84.700 205.100 ;
        RECT 85.400 205.200 85.700 206.800 ;
        RECT 86.200 206.400 86.600 206.500 ;
        RECT 86.200 206.100 88.100 206.400 ;
        RECT 87.700 206.000 88.100 206.100 ;
        RECT 86.900 205.700 87.300 205.800 ;
        RECT 88.600 205.700 89.000 207.400 ;
        RECT 89.400 208.500 89.800 209.500 ;
        RECT 89.400 207.400 89.700 208.500 ;
        RECT 91.500 208.000 91.900 209.500 ;
        RECT 96.100 208.000 96.500 209.500 ;
        RECT 98.200 208.500 98.600 209.500 ;
        RECT 91.500 207.700 92.300 208.000 ;
        RECT 91.900 207.500 92.300 207.700 ;
        RECT 89.400 207.100 91.500 207.400 ;
        RECT 91.000 206.900 91.500 207.100 ;
        RECT 92.000 207.200 92.300 207.500 ;
        RECT 95.700 207.700 96.500 208.000 ;
        RECT 95.700 207.500 96.100 207.700 ;
        RECT 95.700 207.200 96.000 207.500 ;
        RECT 98.300 207.400 98.600 208.500 ;
        RECT 101.900 209.200 102.300 209.900 ;
        RECT 101.900 208.800 102.600 209.200 ;
        RECT 101.900 208.200 102.300 208.800 ;
        RECT 101.400 207.900 102.300 208.200 ;
        RECT 89.400 205.800 89.800 206.600 ;
        RECT 90.200 205.800 90.600 206.600 ;
        RECT 91.000 206.500 91.700 206.900 ;
        RECT 92.000 206.800 93.000 207.200 ;
        RECT 95.000 206.800 96.000 207.200 ;
        RECT 96.500 207.100 98.600 207.400 ;
        RECT 96.500 206.900 97.000 207.100 ;
        RECT 86.900 205.400 89.000 205.700 ;
        RECT 91.000 205.500 91.300 206.500 ;
        RECT 85.400 204.900 86.600 205.200 ;
        RECT 85.100 204.500 85.500 204.600 ;
        RECT 84.400 204.200 85.500 204.500 ;
        RECT 86.300 204.400 86.600 204.900 ;
        RECT 86.300 204.000 87.000 204.400 ;
        RECT 83.100 203.700 83.500 203.800 ;
        RECT 84.500 203.700 84.900 203.800 ;
        RECT 81.400 203.100 81.800 203.500 ;
        RECT 83.100 203.400 84.900 203.700 ;
        RECT 84.200 203.100 84.500 203.400 ;
        RECT 86.200 203.100 86.600 203.500 ;
        RECT 81.400 202.800 82.400 203.100 ;
        RECT 82.000 201.100 82.400 202.800 ;
        RECT 84.200 201.100 84.600 203.100 ;
        RECT 86.300 201.100 86.900 203.100 ;
        RECT 88.600 201.100 89.000 205.400 ;
        RECT 89.400 205.200 91.300 205.500 ;
        RECT 89.400 203.500 89.700 205.200 ;
        RECT 92.000 204.900 92.300 206.800 ;
        RECT 92.600 206.100 93.000 206.200 ;
        RECT 94.200 206.100 94.600 206.200 ;
        RECT 92.600 205.800 94.600 206.100 ;
        RECT 92.600 205.400 93.000 205.800 ;
        RECT 95.000 205.400 95.400 206.200 ;
        RECT 91.500 204.600 92.300 204.900 ;
        RECT 95.700 204.900 96.000 206.800 ;
        RECT 96.300 206.500 97.000 206.900 ;
        RECT 100.600 206.800 101.000 207.600 ;
        RECT 96.700 205.500 97.000 206.500 ;
        RECT 97.400 205.800 97.800 206.600 ;
        RECT 98.200 205.800 98.600 206.600 ;
        RECT 96.700 205.200 98.600 205.500 ;
        RECT 95.700 204.600 96.500 204.900 ;
        RECT 89.400 201.500 89.800 203.500 ;
        RECT 91.500 202.200 91.900 204.600 ;
        RECT 96.100 202.200 96.500 204.600 ;
        RECT 98.300 203.500 98.600 205.200 ;
        RECT 91.500 201.800 92.200 202.200 ;
        RECT 95.800 201.800 96.500 202.200 ;
        RECT 91.500 201.100 91.900 201.800 ;
        RECT 96.100 201.100 96.500 201.800 ;
        RECT 98.200 201.500 98.600 203.500 ;
        RECT 101.400 201.100 101.800 207.900 ;
        RECT 103.000 207.700 103.400 209.900 ;
        RECT 105.100 209.200 105.700 209.900 ;
        RECT 105.100 208.900 105.800 209.200 ;
        RECT 107.400 208.900 107.800 209.900 ;
        RECT 109.600 209.200 110.000 209.900 ;
        RECT 109.600 208.900 110.600 209.200 ;
        RECT 105.400 208.500 105.800 208.900 ;
        RECT 107.500 208.600 107.800 208.900 ;
        RECT 107.500 208.300 108.900 208.600 ;
        RECT 108.500 208.200 108.900 208.300 ;
        RECT 109.400 208.200 109.800 208.600 ;
        RECT 110.200 208.500 110.600 208.900 ;
        RECT 104.500 207.700 104.900 207.800 ;
        RECT 103.000 207.400 104.900 207.700 ;
        RECT 103.000 205.700 103.400 207.400 ;
        RECT 106.500 207.100 106.900 207.200 ;
        RECT 109.400 207.100 109.700 208.200 ;
        RECT 111.800 207.500 112.200 209.900 ;
        RECT 112.600 208.500 113.000 209.500 ;
        RECT 112.600 207.400 112.900 208.500 ;
        RECT 114.700 208.000 115.100 209.500 ;
        RECT 114.700 207.700 115.500 208.000 ;
        RECT 115.100 207.500 115.500 207.700 ;
        RECT 111.000 207.100 111.800 207.200 ;
        RECT 112.600 207.100 114.700 207.400 ;
        RECT 106.300 206.800 111.800 207.100 ;
        RECT 114.200 206.900 114.700 207.100 ;
        RECT 115.200 207.200 115.500 207.500 ;
        RECT 117.400 207.600 117.800 209.900 ;
        RECT 119.000 208.200 119.400 209.900 ;
        RECT 119.000 207.900 119.500 208.200 ;
        RECT 117.400 207.300 118.700 207.600 ;
        RECT 105.400 206.400 105.800 206.500 ;
        RECT 103.900 206.100 105.800 206.400 ;
        RECT 103.900 206.000 104.300 206.100 ;
        RECT 104.700 205.700 105.100 205.800 ;
        RECT 103.000 205.400 105.100 205.700 ;
        RECT 102.200 204.400 102.600 205.200 ;
        RECT 103.000 201.100 103.400 205.400 ;
        RECT 106.300 205.200 106.600 206.800 ;
        RECT 109.900 206.700 110.300 206.800 ;
        RECT 110.700 206.200 111.100 206.300 ;
        RECT 107.800 206.100 108.200 206.200 ;
        RECT 108.600 206.100 111.100 206.200 ;
        RECT 107.800 205.900 111.100 206.100 ;
        RECT 107.800 205.800 109.000 205.900 ;
        RECT 112.600 205.800 113.000 206.600 ;
        RECT 113.400 205.800 113.800 206.600 ;
        RECT 114.200 206.500 114.900 206.900 ;
        RECT 115.200 206.800 116.200 207.200 ;
        RECT 109.400 205.500 112.200 205.600 ;
        RECT 114.200 205.500 114.500 206.500 ;
        RECT 109.300 205.400 112.200 205.500 ;
        RECT 105.400 204.900 106.600 205.200 ;
        RECT 107.300 205.300 112.200 205.400 ;
        RECT 107.300 205.100 109.700 205.300 ;
        RECT 105.400 204.400 105.700 204.900 ;
        RECT 105.000 204.000 105.700 204.400 ;
        RECT 106.500 204.500 106.900 204.600 ;
        RECT 107.300 204.500 107.600 205.100 ;
        RECT 106.500 204.200 107.600 204.500 ;
        RECT 107.900 204.500 110.600 204.800 ;
        RECT 107.900 204.400 108.300 204.500 ;
        RECT 110.200 204.400 110.600 204.500 ;
        RECT 107.100 203.700 107.500 203.800 ;
        RECT 108.500 203.700 108.900 203.800 ;
        RECT 105.400 203.100 105.800 203.500 ;
        RECT 107.100 203.400 108.900 203.700 ;
        RECT 107.500 203.100 107.800 203.400 ;
        RECT 110.200 203.100 110.600 203.500 ;
        RECT 105.100 201.100 105.700 203.100 ;
        RECT 107.400 201.100 107.800 203.100 ;
        RECT 109.600 202.800 110.600 203.100 ;
        RECT 109.600 201.100 110.000 202.800 ;
        RECT 111.800 201.100 112.200 205.300 ;
        RECT 112.600 205.200 114.500 205.500 ;
        RECT 112.600 203.500 112.900 205.200 ;
        RECT 115.200 204.900 115.500 206.800 ;
        RECT 117.500 206.200 117.900 206.600 ;
        RECT 115.800 205.400 116.200 206.200 ;
        RECT 117.400 205.800 117.900 206.200 ;
        RECT 118.400 206.500 118.700 207.300 ;
        RECT 119.200 207.200 119.500 207.900 ;
        RECT 122.200 207.900 122.600 209.900 ;
        RECT 122.900 208.200 123.300 208.600 ;
        RECT 123.800 208.500 124.200 209.500 ;
        RECT 119.000 206.800 119.500 207.200 ;
        RECT 118.400 206.100 118.900 206.500 ;
        RECT 118.400 205.100 118.700 206.100 ;
        RECT 119.200 205.100 119.500 206.800 ;
        RECT 121.400 206.400 121.800 207.200 ;
        RECT 119.800 206.100 120.200 206.200 ;
        RECT 120.600 206.100 121.000 206.200 ;
        RECT 122.200 206.100 122.500 207.900 ;
        RECT 123.000 207.800 123.400 208.200 ;
        RECT 123.800 207.400 124.100 208.500 ;
        RECT 125.900 208.000 126.300 209.500 ;
        RECT 125.900 207.700 126.700 208.000 ;
        RECT 126.300 207.500 126.700 207.700 ;
        RECT 123.800 207.100 125.900 207.400 ;
        RECT 125.400 206.900 125.900 207.100 ;
        RECT 126.400 207.200 126.700 207.500 ;
        RECT 128.600 207.700 129.000 209.900 ;
        RECT 130.700 209.200 131.300 209.900 ;
        RECT 130.700 208.900 131.400 209.200 ;
        RECT 133.000 208.900 133.400 209.900 ;
        RECT 135.200 209.200 135.600 209.900 ;
        RECT 135.200 208.900 136.200 209.200 ;
        RECT 131.000 208.500 131.400 208.900 ;
        RECT 133.100 208.600 133.400 208.900 ;
        RECT 133.100 208.300 134.500 208.600 ;
        RECT 134.100 208.200 134.500 208.300 ;
        RECT 135.000 208.200 135.400 208.600 ;
        RECT 135.800 208.500 136.200 208.900 ;
        RECT 130.100 207.700 130.500 207.800 ;
        RECT 128.600 207.400 130.500 207.700 ;
        RECT 123.000 206.100 123.400 206.200 ;
        RECT 119.800 205.800 121.400 206.100 ;
        RECT 122.200 205.800 123.400 206.100 ;
        RECT 123.800 205.800 124.200 206.600 ;
        RECT 124.600 205.800 125.000 206.600 ;
        RECT 125.400 206.500 126.100 206.900 ;
        RECT 126.400 206.800 127.400 207.200 ;
        RECT 121.000 205.600 121.400 205.800 ;
        RECT 123.000 205.100 123.300 205.800 ;
        RECT 125.400 205.500 125.700 206.500 ;
        RECT 123.800 205.200 125.700 205.500 ;
        RECT 114.700 204.600 115.500 204.900 ;
        RECT 117.400 204.800 118.700 205.100 ;
        RECT 112.600 201.500 113.000 203.500 ;
        RECT 114.700 202.200 115.100 204.600 ;
        RECT 114.700 201.800 115.400 202.200 ;
        RECT 114.700 201.100 115.100 201.800 ;
        RECT 117.400 201.100 117.800 204.800 ;
        RECT 119.000 204.600 119.500 205.100 ;
        RECT 120.600 204.800 122.600 205.100 ;
        RECT 119.000 201.100 119.400 204.600 ;
        RECT 120.600 201.100 121.000 204.800 ;
        RECT 122.200 201.100 122.600 204.800 ;
        RECT 123.000 201.100 123.400 205.100 ;
        RECT 123.800 203.500 124.100 205.200 ;
        RECT 126.400 204.900 126.700 206.800 ;
        RECT 127.000 205.400 127.400 206.200 ;
        RECT 128.600 205.700 129.000 207.400 ;
        RECT 132.100 207.100 132.500 207.200 ;
        RECT 135.000 207.100 135.300 208.200 ;
        RECT 137.400 207.500 137.800 209.900 ;
        RECT 139.000 208.900 139.400 209.900 ;
        RECT 138.200 207.800 138.600 208.600 ;
        RECT 139.100 208.100 139.400 208.900 ;
        RECT 140.700 208.200 141.100 208.600 ;
        RECT 140.600 208.100 141.000 208.200 ;
        RECT 139.000 207.800 141.000 208.100 ;
        RECT 141.400 207.900 141.800 209.900 ;
        RECT 139.100 207.200 139.400 207.800 ;
        RECT 136.600 207.100 137.400 207.200 ;
        RECT 131.900 206.800 137.400 207.100 ;
        RECT 139.000 206.800 139.400 207.200 ;
        RECT 131.000 206.400 131.400 206.500 ;
        RECT 129.500 206.100 131.400 206.400 ;
        RECT 129.500 206.000 129.900 206.100 ;
        RECT 130.300 205.700 130.700 205.800 ;
        RECT 128.600 205.400 130.700 205.700 ;
        RECT 125.900 204.600 126.700 204.900 ;
        RECT 123.800 201.500 124.200 203.500 ;
        RECT 125.900 202.200 126.300 204.600 ;
        RECT 125.900 201.800 126.600 202.200 ;
        RECT 125.900 201.100 126.300 201.800 ;
        RECT 128.600 201.100 129.000 205.400 ;
        RECT 131.900 205.200 132.200 206.800 ;
        RECT 135.500 206.700 135.900 206.800 ;
        RECT 135.000 206.200 135.400 206.300 ;
        RECT 136.300 206.200 136.700 206.300 ;
        RECT 134.200 205.900 136.700 206.200 ;
        RECT 134.200 205.800 134.600 205.900 ;
        RECT 135.000 205.500 137.800 205.600 ;
        RECT 134.900 205.400 137.800 205.500 ;
        RECT 131.000 204.900 132.200 205.200 ;
        RECT 132.900 205.300 137.800 205.400 ;
        RECT 132.900 205.100 135.300 205.300 ;
        RECT 131.000 204.400 131.300 204.900 ;
        RECT 130.600 204.000 131.300 204.400 ;
        RECT 132.100 204.500 132.500 204.600 ;
        RECT 132.900 204.500 133.200 205.100 ;
        RECT 132.100 204.200 133.200 204.500 ;
        RECT 133.500 204.500 136.200 204.800 ;
        RECT 133.500 204.400 133.900 204.500 ;
        RECT 135.800 204.400 136.200 204.500 ;
        RECT 132.700 203.700 133.100 203.800 ;
        RECT 134.100 203.700 134.500 203.800 ;
        RECT 131.000 203.100 131.400 203.500 ;
        RECT 132.700 203.400 134.500 203.700 ;
        RECT 133.100 203.100 133.400 203.400 ;
        RECT 135.800 203.100 136.200 203.500 ;
        RECT 130.700 201.100 131.300 203.100 ;
        RECT 133.000 201.100 133.400 203.100 ;
        RECT 135.200 202.800 136.200 203.100 ;
        RECT 135.200 201.100 135.600 202.800 ;
        RECT 137.400 201.100 137.800 205.300 ;
        RECT 139.100 205.100 139.400 206.800 ;
        RECT 139.800 205.400 140.200 206.200 ;
        RECT 140.600 206.100 141.000 206.200 ;
        RECT 141.500 206.100 141.800 207.900 ;
        RECT 144.600 208.800 145.000 209.900 ;
        RECT 144.600 207.200 144.900 208.800 ;
        RECT 145.400 207.800 145.800 208.600 ;
        RECT 146.300 208.200 146.700 208.600 ;
        RECT 146.200 207.800 146.600 208.200 ;
        RECT 147.000 207.900 147.400 209.900 ;
        RECT 142.200 206.400 142.600 207.200 ;
        RECT 144.600 206.800 145.000 207.200 ;
        RECT 143.000 206.100 143.400 206.200 ;
        RECT 140.600 205.800 141.800 206.100 ;
        RECT 142.600 205.800 143.400 206.100 ;
        RECT 140.700 205.100 141.000 205.800 ;
        RECT 142.600 205.600 143.000 205.800 ;
        RECT 143.800 205.400 144.200 206.200 ;
        RECT 144.600 205.100 144.900 206.800 ;
        RECT 146.200 206.100 146.600 206.200 ;
        RECT 147.100 206.100 147.400 207.900 ;
        RECT 151.000 207.500 151.400 209.900 ;
        RECT 153.200 209.200 153.600 209.900 ;
        RECT 152.600 208.900 153.600 209.200 ;
        RECT 155.400 208.900 155.800 209.900 ;
        RECT 157.500 209.200 158.100 209.900 ;
        RECT 157.400 208.900 158.100 209.200 ;
        RECT 152.600 208.500 153.000 208.900 ;
        RECT 155.400 208.600 155.700 208.900 ;
        RECT 153.400 208.200 153.800 208.600 ;
        RECT 154.300 208.300 155.700 208.600 ;
        RECT 157.400 208.500 157.800 208.900 ;
        RECT 154.300 208.200 154.700 208.300 ;
        RECT 147.800 206.400 148.200 207.200 ;
        RECT 150.200 207.100 150.600 207.200 ;
        RECT 151.400 207.100 152.200 207.200 ;
        RECT 153.500 207.100 153.800 208.200 ;
        RECT 158.300 207.700 158.700 207.800 ;
        RECT 159.800 207.700 160.200 209.900 ;
        RECT 158.300 207.400 160.200 207.700 ;
        RECT 156.300 207.100 156.700 207.200 ;
        RECT 150.200 206.800 156.900 207.100 ;
        RECT 152.900 206.700 153.300 206.800 ;
        RECT 152.100 206.200 152.500 206.300 ;
        RECT 156.600 206.200 156.900 206.800 ;
        RECT 157.400 206.400 157.800 206.500 ;
        RECT 148.600 206.100 149.000 206.200 ;
        RECT 146.200 205.800 147.400 206.100 ;
        RECT 148.200 205.800 149.000 206.100 ;
        RECT 152.100 205.900 154.600 206.200 ;
        RECT 154.200 205.800 154.600 205.900 ;
        RECT 156.600 205.800 157.000 206.200 ;
        RECT 157.400 206.100 159.300 206.400 ;
        RECT 158.900 206.000 159.300 206.100 ;
        RECT 146.300 205.100 146.600 205.800 ;
        RECT 148.200 205.600 148.600 205.800 ;
        RECT 151.000 205.500 153.800 205.600 ;
        RECT 151.000 205.400 153.900 205.500 ;
        RECT 151.000 205.300 155.900 205.400 ;
        RECT 139.000 204.700 139.900 205.100 ;
        RECT 139.500 201.100 139.900 204.700 ;
        RECT 140.600 201.100 141.000 205.100 ;
        RECT 141.400 204.800 143.400 205.100 ;
        RECT 141.400 201.100 141.800 204.800 ;
        RECT 143.000 201.100 143.400 204.800 ;
        RECT 144.100 204.700 145.000 205.100 ;
        RECT 144.100 201.100 144.500 204.700 ;
        RECT 146.200 201.100 146.600 205.100 ;
        RECT 147.000 204.800 149.000 205.100 ;
        RECT 147.000 201.100 147.400 204.800 ;
        RECT 148.600 201.100 149.000 204.800 ;
        RECT 151.000 201.100 151.400 205.300 ;
        RECT 153.500 205.100 155.900 205.300 ;
        RECT 152.600 204.500 155.300 204.800 ;
        RECT 152.600 204.400 153.000 204.500 ;
        RECT 154.900 204.400 155.300 204.500 ;
        RECT 155.600 204.500 155.900 205.100 ;
        RECT 156.600 205.200 156.900 205.800 ;
        RECT 158.100 205.700 158.500 205.800 ;
        RECT 159.800 205.700 160.200 207.400 ;
        RECT 160.600 208.500 161.000 209.500 ;
        RECT 160.600 207.400 160.900 208.500 ;
        RECT 162.700 208.000 163.100 209.500 ;
        RECT 165.400 208.000 165.800 209.900 ;
        RECT 167.000 208.000 167.400 209.900 ;
        RECT 162.700 207.700 163.500 208.000 ;
        RECT 165.400 207.900 167.400 208.000 ;
        RECT 167.800 207.900 168.200 209.900 ;
        RECT 168.900 208.200 169.300 209.900 ;
        RECT 168.900 207.900 169.800 208.200 ;
        RECT 165.500 207.700 167.300 207.900 ;
        RECT 163.100 207.500 163.500 207.700 ;
        RECT 160.600 207.100 162.700 207.400 ;
        RECT 162.200 206.900 162.700 207.100 ;
        RECT 163.200 207.200 163.500 207.500 ;
        RECT 165.800 207.200 166.200 207.400 ;
        RECT 167.800 207.200 168.100 207.900 ;
        RECT 160.600 205.800 161.000 206.600 ;
        RECT 161.400 205.800 161.800 206.600 ;
        RECT 162.200 206.500 162.900 206.900 ;
        RECT 163.200 206.800 164.200 207.200 ;
        RECT 165.400 206.900 166.200 207.200 ;
        RECT 166.900 207.100 168.200 207.200 ;
        RECT 168.600 207.100 169.000 207.200 ;
        RECT 165.400 206.800 165.800 206.900 ;
        RECT 166.900 206.800 169.000 207.100 ;
        RECT 158.100 205.400 160.200 205.700 ;
        RECT 162.200 205.500 162.500 206.500 ;
        RECT 156.600 204.900 157.800 205.200 ;
        RECT 156.300 204.500 156.700 204.600 ;
        RECT 155.600 204.200 156.700 204.500 ;
        RECT 157.500 204.400 157.800 204.900 ;
        RECT 157.500 204.000 158.200 204.400 ;
        RECT 154.300 203.700 154.700 203.800 ;
        RECT 155.700 203.700 156.100 203.800 ;
        RECT 152.600 203.100 153.000 203.500 ;
        RECT 154.300 203.400 156.100 203.700 ;
        RECT 155.400 203.100 155.700 203.400 ;
        RECT 157.400 203.100 157.800 203.500 ;
        RECT 152.600 202.800 153.600 203.100 ;
        RECT 153.200 201.100 153.600 202.800 ;
        RECT 155.400 201.100 155.800 203.100 ;
        RECT 157.500 201.100 158.100 203.100 ;
        RECT 159.800 201.100 160.200 205.400 ;
        RECT 160.600 205.200 162.500 205.500 ;
        RECT 160.600 203.500 160.900 205.200 ;
        RECT 163.200 204.900 163.500 206.800 ;
        RECT 163.800 205.400 164.200 206.200 ;
        RECT 166.200 205.800 166.600 206.600 ;
        RECT 166.900 205.100 167.200 206.800 ;
        RECT 169.400 206.100 169.800 207.900 ;
        RECT 170.200 206.800 170.600 207.600 ;
        RECT 171.000 207.500 171.400 209.900 ;
        RECT 173.200 209.200 173.600 209.900 ;
        RECT 172.600 208.900 173.600 209.200 ;
        RECT 175.400 208.900 175.800 209.900 ;
        RECT 177.500 209.200 178.100 209.900 ;
        RECT 177.400 208.900 178.100 209.200 ;
        RECT 172.600 208.500 173.000 208.900 ;
        RECT 175.400 208.600 175.700 208.900 ;
        RECT 173.400 208.200 173.800 208.600 ;
        RECT 174.300 208.300 175.700 208.600 ;
        RECT 177.400 208.500 177.800 208.900 ;
        RECT 174.300 208.200 174.700 208.300 ;
        RECT 171.400 207.100 172.200 207.200 ;
        RECT 173.500 207.100 173.800 208.200 ;
        RECT 178.300 207.700 178.700 207.800 ;
        RECT 179.800 207.700 180.200 209.900 ;
        RECT 180.700 208.200 181.100 208.600 ;
        RECT 180.600 207.800 181.000 208.200 ;
        RECT 181.400 207.900 181.800 209.900 ;
        RECT 185.700 208.000 186.100 209.500 ;
        RECT 187.800 208.500 188.200 209.500 ;
        RECT 178.300 207.400 180.200 207.700 ;
        RECT 176.300 207.100 176.700 207.200 ;
        RECT 171.400 206.800 176.900 207.100 ;
        RECT 172.900 206.700 173.300 206.800 ;
        RECT 167.800 205.800 169.800 206.100 ;
        RECT 172.100 206.200 172.500 206.300 ;
        RECT 173.400 206.200 173.800 206.300 ;
        RECT 172.100 205.900 174.600 206.200 ;
        RECT 174.200 205.800 174.600 205.900 ;
        RECT 167.800 205.200 168.100 205.800 ;
        RECT 167.800 205.100 168.200 205.200 ;
        RECT 162.700 204.600 163.500 204.900 ;
        RECT 166.700 204.800 167.200 205.100 ;
        RECT 167.500 204.800 168.200 205.100 ;
        RECT 160.600 201.500 161.000 203.500 ;
        RECT 162.700 202.200 163.100 204.600 ;
        RECT 162.700 201.800 163.400 202.200 ;
        RECT 162.700 201.100 163.100 201.800 ;
        RECT 166.700 201.100 167.100 204.800 ;
        RECT 167.500 204.200 167.800 204.800 ;
        RECT 168.600 204.400 169.000 205.200 ;
        RECT 167.400 203.800 167.800 204.200 ;
        RECT 169.400 201.100 169.800 205.800 ;
        RECT 171.000 205.500 173.800 205.600 ;
        RECT 171.000 205.400 173.900 205.500 ;
        RECT 171.000 205.300 175.900 205.400 ;
        RECT 171.000 201.100 171.400 205.300 ;
        RECT 173.500 205.100 175.900 205.300 ;
        RECT 172.600 204.500 175.300 204.800 ;
        RECT 172.600 204.400 173.000 204.500 ;
        RECT 174.900 204.400 175.300 204.500 ;
        RECT 175.600 204.500 175.900 205.100 ;
        RECT 176.600 205.200 176.900 206.800 ;
        RECT 177.400 206.400 177.800 206.500 ;
        RECT 177.400 206.100 179.300 206.400 ;
        RECT 178.900 206.000 179.300 206.100 ;
        RECT 178.100 205.700 178.500 205.800 ;
        RECT 179.800 205.700 180.200 207.400 ;
        RECT 180.600 206.100 181.000 206.200 ;
        RECT 181.500 206.100 181.800 207.900 ;
        RECT 185.300 207.700 186.100 208.000 ;
        RECT 185.300 207.500 185.700 207.700 ;
        RECT 185.300 207.200 185.600 207.500 ;
        RECT 187.900 207.400 188.200 208.500 ;
        RECT 190.500 208.000 190.900 209.500 ;
        RECT 192.600 208.500 193.000 209.500 ;
        RECT 182.200 207.100 182.600 207.200 ;
        RECT 183.800 207.100 184.200 207.200 ;
        RECT 182.200 206.800 184.200 207.100 ;
        RECT 184.600 206.800 185.600 207.200 ;
        RECT 186.100 207.100 188.200 207.400 ;
        RECT 190.100 207.700 190.900 208.000 ;
        RECT 190.100 207.500 190.500 207.700 ;
        RECT 190.100 207.200 190.400 207.500 ;
        RECT 192.700 207.400 193.000 208.500 ;
        RECT 186.100 206.900 186.600 207.100 ;
        RECT 182.200 206.400 182.600 206.800 ;
        RECT 183.000 206.100 183.400 206.200 ;
        RECT 180.600 205.800 181.800 206.100 ;
        RECT 182.600 205.800 183.400 206.100 ;
        RECT 178.100 205.400 180.200 205.700 ;
        RECT 176.600 204.900 177.800 205.200 ;
        RECT 176.300 204.500 176.700 204.600 ;
        RECT 175.600 204.200 176.700 204.500 ;
        RECT 177.500 204.400 177.800 204.900 ;
        RECT 177.500 204.000 178.200 204.400 ;
        RECT 174.300 203.700 174.700 203.800 ;
        RECT 175.700 203.700 176.100 203.800 ;
        RECT 172.600 203.100 173.000 203.500 ;
        RECT 174.300 203.400 176.100 203.700 ;
        RECT 175.400 203.100 175.700 203.400 ;
        RECT 177.400 203.100 177.800 203.500 ;
        RECT 172.600 202.800 173.600 203.100 ;
        RECT 173.200 201.100 173.600 202.800 ;
        RECT 175.400 201.100 175.800 203.100 ;
        RECT 177.500 201.100 178.100 203.100 ;
        RECT 179.800 201.100 180.200 205.400 ;
        RECT 180.700 205.100 181.000 205.800 ;
        RECT 182.600 205.600 183.000 205.800 ;
        RECT 184.600 205.400 185.000 206.200 ;
        RECT 180.600 201.100 181.000 205.100 ;
        RECT 181.400 204.800 183.400 205.100 ;
        RECT 181.400 201.100 181.800 204.800 ;
        RECT 183.000 201.100 183.400 204.800 ;
        RECT 185.300 204.900 185.600 206.800 ;
        RECT 185.900 206.500 186.600 206.900 ;
        RECT 189.400 206.800 190.400 207.200 ;
        RECT 190.900 207.100 193.000 207.400 ;
        RECT 194.200 208.800 194.600 209.900 ;
        RECT 194.200 207.200 194.500 208.800 ;
        RECT 195.000 207.800 195.400 208.600 ;
        RECT 195.900 208.200 196.300 208.600 ;
        RECT 195.800 207.800 196.200 208.200 ;
        RECT 196.600 207.900 197.000 209.900 ;
        RECT 199.000 208.000 199.400 209.900 ;
        RECT 200.600 208.000 201.000 209.900 ;
        RECT 199.000 207.900 201.000 208.000 ;
        RECT 201.400 207.900 201.800 209.900 ;
        RECT 202.200 209.100 202.600 209.200 ;
        RECT 203.800 209.100 204.200 209.900 ;
        RECT 202.200 208.800 204.200 209.100 ;
        RECT 205.900 209.200 206.500 209.900 ;
        RECT 205.900 208.900 206.600 209.200 ;
        RECT 208.200 208.900 208.600 209.900 ;
        RECT 210.400 209.200 210.800 209.900 ;
        RECT 210.400 208.900 211.400 209.200 ;
        RECT 195.000 207.200 195.300 207.800 ;
        RECT 190.900 206.900 191.400 207.100 ;
        RECT 186.300 205.500 186.600 206.500 ;
        RECT 187.000 205.800 187.400 206.600 ;
        RECT 187.800 205.800 188.200 206.600 ;
        RECT 188.600 206.100 189.000 206.200 ;
        RECT 189.400 206.100 189.800 206.200 ;
        RECT 188.600 205.800 189.800 206.100 ;
        RECT 186.300 205.200 188.200 205.500 ;
        RECT 189.400 205.400 189.800 205.800 ;
        RECT 185.300 204.600 186.100 204.900 ;
        RECT 185.700 202.200 186.100 204.600 ;
        RECT 187.900 203.500 188.200 205.200 ;
        RECT 190.100 204.900 190.400 206.800 ;
        RECT 190.700 206.500 191.400 206.900 ;
        RECT 194.200 206.800 194.600 207.200 ;
        RECT 195.000 206.800 195.400 207.200 ;
        RECT 191.100 205.500 191.400 206.500 ;
        RECT 191.800 205.800 192.200 206.600 ;
        RECT 192.600 205.800 193.000 206.600 ;
        RECT 191.100 205.200 193.000 205.500 ;
        RECT 193.400 205.400 193.800 206.200 ;
        RECT 190.100 204.600 190.900 204.900 ;
        RECT 185.700 201.800 186.600 202.200 ;
        RECT 185.700 201.100 186.100 201.800 ;
        RECT 187.800 201.500 188.200 203.500 ;
        RECT 190.500 201.100 190.900 204.600 ;
        RECT 192.700 203.500 193.000 205.200 ;
        RECT 194.200 205.100 194.500 206.800 ;
        RECT 196.700 206.200 197.000 207.900 ;
        RECT 199.100 207.700 200.900 207.900 ;
        RECT 199.400 207.200 199.800 207.400 ;
        RECT 201.400 207.200 201.700 207.900 ;
        RECT 203.800 207.700 204.200 208.800 ;
        RECT 206.200 208.500 206.600 208.900 ;
        RECT 208.300 208.600 208.600 208.900 ;
        RECT 208.300 208.300 209.700 208.600 ;
        RECT 209.300 208.200 209.700 208.300 ;
        RECT 210.200 208.200 210.600 208.600 ;
        RECT 211.000 208.500 211.400 208.900 ;
        RECT 205.300 207.700 205.700 207.800 ;
        RECT 203.800 207.400 205.700 207.700 ;
        RECT 197.400 206.400 197.800 207.200 ;
        RECT 199.000 207.100 199.800 207.200 ;
        RECT 198.200 206.900 199.800 207.100 ;
        RECT 198.200 206.800 199.400 206.900 ;
        RECT 200.500 206.800 201.800 207.200 ;
        RECT 195.800 206.100 196.200 206.200 ;
        RECT 196.600 206.100 197.000 206.200 ;
        RECT 198.200 206.200 198.500 206.800 ;
        RECT 198.200 206.100 198.600 206.200 ;
        RECT 195.800 205.800 197.000 206.100 ;
        RECT 197.800 205.800 198.600 206.100 ;
        RECT 199.800 205.800 200.200 206.600 ;
        RECT 195.900 205.100 196.200 205.800 ;
        RECT 197.800 205.600 198.200 205.800 ;
        RECT 200.500 205.100 200.800 206.800 ;
        RECT 203.800 205.700 204.200 207.400 ;
        RECT 207.300 207.100 207.700 207.200 ;
        RECT 209.400 207.100 209.800 207.200 ;
        RECT 210.200 207.100 210.500 208.200 ;
        RECT 212.600 207.500 213.000 209.900 ;
        RECT 214.200 207.600 214.600 209.900 ;
        RECT 215.800 207.600 216.200 209.900 ;
        RECT 217.400 207.600 217.800 209.900 ;
        RECT 219.000 207.600 219.400 209.900 ;
        RECT 222.500 208.000 222.900 209.500 ;
        RECT 224.600 208.500 225.000 209.500 ;
        RECT 213.400 207.200 214.600 207.600 ;
        RECT 215.100 207.200 216.200 207.600 ;
        RECT 216.700 207.200 217.800 207.600 ;
        RECT 218.500 207.200 219.400 207.600 ;
        RECT 222.100 207.700 222.900 208.000 ;
        RECT 222.100 207.500 222.500 207.700 ;
        RECT 222.100 207.200 222.400 207.500 ;
        RECT 224.700 207.400 225.000 208.500 ;
        RECT 211.800 207.100 212.600 207.200 ;
        RECT 207.100 206.800 212.600 207.100 ;
        RECT 206.200 206.400 206.600 206.500 ;
        RECT 204.700 206.100 206.600 206.400 ;
        RECT 204.700 206.000 205.100 206.100 ;
        RECT 205.500 205.700 205.900 205.800 ;
        RECT 203.800 205.400 205.900 205.700 ;
        RECT 201.400 205.100 201.800 205.200 ;
        RECT 192.600 201.500 193.000 203.500 ;
        RECT 193.700 204.700 194.600 205.100 ;
        RECT 193.700 201.100 194.100 204.700 ;
        RECT 195.800 201.100 196.200 205.100 ;
        RECT 196.600 204.800 198.600 205.100 ;
        RECT 196.600 201.100 197.000 204.800 ;
        RECT 198.200 201.100 198.600 204.800 ;
        RECT 200.300 204.800 200.800 205.100 ;
        RECT 201.100 204.800 201.800 205.100 ;
        RECT 200.300 202.200 200.700 204.800 ;
        RECT 201.100 204.200 201.400 204.800 ;
        RECT 201.000 203.800 201.400 204.200 ;
        RECT 199.800 201.800 200.700 202.200 ;
        RECT 200.300 201.100 200.700 201.800 ;
        RECT 203.800 201.100 204.200 205.400 ;
        RECT 207.100 205.200 207.400 206.800 ;
        RECT 210.700 206.700 211.100 206.800 ;
        RECT 211.500 206.200 211.900 206.300 ;
        RECT 208.600 206.100 209.000 206.200 ;
        RECT 209.400 206.100 211.900 206.200 ;
        RECT 208.600 205.900 211.900 206.100 ;
        RECT 208.600 205.800 209.800 205.900 ;
        RECT 213.400 205.800 213.800 207.200 ;
        RECT 215.100 206.900 215.500 207.200 ;
        RECT 216.700 206.900 217.100 207.200 ;
        RECT 218.500 206.900 218.900 207.200 ;
        RECT 219.800 206.900 220.200 207.200 ;
        RECT 214.200 206.500 215.500 206.900 ;
        RECT 215.900 206.500 217.100 206.900 ;
        RECT 217.600 206.500 218.900 206.900 ;
        RECT 219.300 206.500 220.200 206.900 ;
        RECT 221.400 206.800 222.400 207.200 ;
        RECT 222.900 207.100 225.000 207.400 ;
        RECT 225.400 208.500 225.800 209.500 ;
        RECT 225.400 207.400 225.700 208.500 ;
        RECT 227.500 208.000 227.900 209.500 ;
        RECT 231.500 209.200 231.900 209.900 ;
        RECT 231.500 208.800 232.200 209.200 ;
        RECT 231.500 208.200 231.900 208.800 ;
        RECT 227.500 207.700 228.300 208.000 ;
        RECT 227.900 207.500 228.300 207.700 ;
        RECT 231.000 207.900 231.900 208.200 ;
        RECT 225.400 207.100 227.500 207.400 ;
        RECT 222.900 206.900 223.400 207.100 ;
        RECT 215.100 205.800 215.500 206.500 ;
        RECT 216.700 205.800 217.100 206.500 ;
        RECT 218.500 205.800 218.900 206.500 ;
        RECT 210.200 205.500 213.000 205.600 ;
        RECT 210.100 205.400 213.000 205.500 ;
        RECT 213.400 205.400 214.600 205.800 ;
        RECT 215.100 205.400 216.200 205.800 ;
        RECT 216.700 205.400 217.800 205.800 ;
        RECT 218.500 205.400 219.400 205.800 ;
        RECT 221.400 205.400 221.800 206.200 ;
        RECT 206.200 204.900 207.400 205.200 ;
        RECT 208.100 205.300 213.000 205.400 ;
        RECT 208.100 205.100 210.500 205.300 ;
        RECT 206.200 204.400 206.500 204.900 ;
        RECT 205.800 204.000 206.500 204.400 ;
        RECT 207.300 204.500 207.700 204.600 ;
        RECT 208.100 204.500 208.400 205.100 ;
        RECT 207.300 204.200 208.400 204.500 ;
        RECT 208.700 204.500 211.400 204.800 ;
        RECT 208.700 204.400 209.100 204.500 ;
        RECT 211.000 204.400 211.400 204.500 ;
        RECT 207.900 203.700 208.300 203.800 ;
        RECT 209.300 203.700 209.700 203.800 ;
        RECT 206.200 203.100 206.600 203.500 ;
        RECT 207.900 203.400 209.700 203.700 ;
        RECT 208.300 203.100 208.600 203.400 ;
        RECT 211.000 203.100 211.400 203.500 ;
        RECT 205.900 201.100 206.500 203.100 ;
        RECT 208.200 201.100 208.600 203.100 ;
        RECT 210.400 202.800 211.400 203.100 ;
        RECT 210.400 201.100 210.800 202.800 ;
        RECT 212.600 201.100 213.000 205.300 ;
        RECT 214.200 201.100 214.600 205.400 ;
        RECT 215.800 201.100 216.200 205.400 ;
        RECT 217.400 201.100 217.800 205.400 ;
        RECT 219.000 201.100 219.400 205.400 ;
        RECT 222.100 204.900 222.400 206.800 ;
        RECT 222.700 206.500 223.400 206.900 ;
        RECT 227.000 206.900 227.500 207.100 ;
        RECT 228.000 207.200 228.300 207.500 ;
        RECT 223.100 205.500 223.400 206.500 ;
        RECT 223.800 205.800 224.200 206.600 ;
        RECT 224.600 205.800 225.000 206.600 ;
        RECT 225.400 205.800 225.800 206.600 ;
        RECT 226.200 205.800 226.600 206.600 ;
        RECT 227.000 206.500 227.700 206.900 ;
        RECT 228.000 206.800 229.000 207.200 ;
        RECT 229.400 207.100 229.800 207.200 ;
        RECT 230.200 207.100 230.600 207.600 ;
        RECT 229.400 206.800 230.600 207.100 ;
        RECT 227.000 205.500 227.300 206.500 ;
        RECT 223.100 205.200 225.000 205.500 ;
        RECT 222.100 204.600 222.900 204.900 ;
        RECT 222.500 202.200 222.900 204.600 ;
        RECT 224.700 203.500 225.000 205.200 ;
        RECT 222.200 201.800 222.900 202.200 ;
        RECT 222.500 201.100 222.900 201.800 ;
        RECT 224.600 201.500 225.000 203.500 ;
        RECT 225.400 205.200 227.300 205.500 ;
        RECT 225.400 203.500 225.700 205.200 ;
        RECT 228.000 204.900 228.300 206.800 ;
        RECT 228.600 205.400 229.000 206.200 ;
        RECT 227.500 204.600 228.300 204.900 ;
        RECT 225.400 201.500 225.800 203.500 ;
        RECT 227.500 202.200 227.900 204.600 ;
        RECT 227.000 201.800 227.900 202.200 ;
        RECT 227.500 201.100 227.900 201.800 ;
        RECT 231.000 201.100 231.400 207.900 ;
        RECT 232.600 207.700 233.000 209.900 ;
        RECT 234.700 209.200 235.300 209.900 ;
        RECT 234.700 208.900 235.400 209.200 ;
        RECT 237.000 208.900 237.400 209.900 ;
        RECT 239.200 209.200 239.600 209.900 ;
        RECT 239.200 208.900 240.200 209.200 ;
        RECT 235.000 208.500 235.400 208.900 ;
        RECT 237.100 208.600 237.400 208.900 ;
        RECT 237.100 208.300 238.500 208.600 ;
        RECT 238.100 208.200 238.500 208.300 ;
        RECT 239.000 207.800 239.400 208.600 ;
        RECT 239.800 208.500 240.200 208.900 ;
        RECT 234.100 207.700 234.500 207.800 ;
        RECT 232.600 207.400 234.500 207.700 ;
        RECT 232.600 205.700 233.000 207.400 ;
        RECT 236.100 207.100 236.500 207.200 ;
        RECT 239.000 207.100 239.300 207.800 ;
        RECT 241.400 207.500 241.800 209.900 ;
        RECT 243.500 208.200 243.900 209.900 ;
        RECT 245.400 208.900 245.800 209.900 ;
        RECT 243.000 207.900 243.900 208.200 ;
        RECT 240.600 207.100 241.400 207.200 ;
        RECT 235.900 206.800 241.400 207.100 ;
        RECT 242.200 206.800 242.600 207.600 ;
        RECT 235.000 206.400 235.400 206.500 ;
        RECT 233.500 206.100 235.400 206.400 ;
        RECT 233.500 206.000 233.900 206.100 ;
        RECT 234.300 205.700 234.700 205.800 ;
        RECT 232.600 205.400 234.700 205.700 ;
        RECT 231.800 204.400 232.200 205.200 ;
        RECT 232.600 201.100 233.000 205.400 ;
        RECT 235.900 205.200 236.200 206.800 ;
        RECT 239.500 206.700 239.900 206.800 ;
        RECT 240.300 206.200 240.700 206.300 ;
        RECT 236.600 206.100 237.000 206.200 ;
        RECT 238.200 206.100 240.700 206.200 ;
        RECT 236.600 205.900 240.700 206.100 ;
        RECT 236.600 205.800 238.600 205.900 ;
        RECT 239.000 205.500 241.800 205.600 ;
        RECT 238.900 205.400 241.800 205.500 ;
        RECT 235.000 204.900 236.200 205.200 ;
        RECT 236.900 205.300 241.800 205.400 ;
        RECT 236.900 205.100 239.300 205.300 ;
        RECT 235.000 204.400 235.300 204.900 ;
        RECT 234.600 204.000 235.300 204.400 ;
        RECT 236.100 204.500 236.500 204.600 ;
        RECT 236.900 204.500 237.200 205.100 ;
        RECT 236.100 204.200 237.200 204.500 ;
        RECT 237.500 204.500 240.200 204.800 ;
        RECT 237.500 204.400 237.900 204.500 ;
        RECT 239.800 204.400 240.200 204.500 ;
        RECT 236.700 203.700 237.100 203.800 ;
        RECT 238.100 203.700 238.500 203.800 ;
        RECT 235.000 203.100 235.400 203.500 ;
        RECT 236.700 203.400 238.500 203.700 ;
        RECT 237.100 203.100 237.400 203.400 ;
        RECT 239.800 203.100 240.200 203.500 ;
        RECT 234.700 201.100 235.300 203.100 ;
        RECT 237.000 201.100 237.400 203.100 ;
        RECT 239.200 202.800 240.200 203.100 ;
        RECT 239.200 201.100 239.600 202.800 ;
        RECT 241.400 201.100 241.800 205.300 ;
        RECT 243.000 201.100 243.400 207.900 ;
        RECT 244.600 207.800 245.000 208.600 ;
        RECT 245.500 208.100 245.800 208.900 ;
        RECT 246.200 208.100 246.600 208.200 ;
        RECT 245.400 207.800 246.600 208.100 ;
        RECT 248.600 207.900 249.000 209.900 ;
        RECT 249.300 208.200 249.700 208.600 ;
        RECT 245.500 207.200 245.800 207.800 ;
        RECT 245.400 206.800 245.800 207.200 ;
        RECT 247.800 207.100 248.200 207.200 ;
        RECT 243.800 204.400 244.200 205.200 ;
        RECT 245.500 205.100 245.800 206.800 ;
        RECT 246.200 206.800 248.200 207.100 ;
        RECT 246.200 206.200 246.500 206.800 ;
        RECT 247.800 206.400 248.200 206.800 ;
        RECT 246.200 205.400 246.600 206.200 ;
        RECT 247.000 206.100 247.400 206.200 ;
        RECT 248.600 206.100 248.900 207.900 ;
        RECT 249.400 207.800 249.800 208.200 ;
        RECT 249.400 206.100 249.800 206.200 ;
        RECT 247.000 205.800 247.800 206.100 ;
        RECT 248.600 205.800 249.800 206.100 ;
        RECT 247.400 205.600 247.800 205.800 ;
        RECT 249.400 205.100 249.700 205.800 ;
        RECT 245.400 204.700 246.300 205.100 ;
        RECT 245.900 201.100 246.300 204.700 ;
        RECT 247.000 204.800 249.000 205.100 ;
        RECT 247.000 201.100 247.400 204.800 ;
        RECT 248.600 201.100 249.000 204.800 ;
        RECT 249.400 201.100 249.800 205.100 ;
        RECT 0.600 195.600 1.000 199.900 ;
        RECT 2.700 197.900 3.300 199.900 ;
        RECT 5.000 197.900 5.400 199.900 ;
        RECT 7.200 198.200 7.600 199.900 ;
        RECT 7.200 197.900 8.200 198.200 ;
        RECT 3.000 197.500 3.400 197.900 ;
        RECT 5.100 197.600 5.400 197.900 ;
        RECT 4.700 197.300 6.500 197.600 ;
        RECT 7.800 197.500 8.200 197.900 ;
        RECT 4.700 197.200 5.100 197.300 ;
        RECT 6.100 197.200 6.500 197.300 ;
        RECT 2.600 196.600 3.300 197.000 ;
        RECT 3.000 196.100 3.300 196.600 ;
        RECT 4.100 196.500 5.200 196.800 ;
        RECT 4.100 196.400 4.500 196.500 ;
        RECT 3.000 195.800 4.200 196.100 ;
        RECT 0.600 195.300 2.700 195.600 ;
        RECT 0.600 193.600 1.000 195.300 ;
        RECT 2.300 195.200 2.700 195.300 ;
        RECT 1.500 194.900 1.900 195.000 ;
        RECT 1.500 194.600 3.400 194.900 ;
        RECT 3.000 194.500 3.400 194.600 ;
        RECT 3.900 194.200 4.200 195.800 ;
        RECT 4.900 195.900 5.200 196.500 ;
        RECT 5.500 196.500 5.900 196.600 ;
        RECT 7.800 196.500 8.200 196.600 ;
        RECT 5.500 196.200 8.200 196.500 ;
        RECT 4.900 195.700 7.300 195.900 ;
        RECT 9.400 195.700 9.800 199.900 ;
        RECT 4.900 195.600 9.800 195.700 ;
        RECT 6.900 195.500 9.800 195.600 ;
        RECT 7.000 195.400 9.800 195.500 ;
        RECT 10.200 195.700 10.600 199.900 ;
        RECT 12.400 198.200 12.800 199.900 ;
        RECT 11.800 197.900 12.800 198.200 ;
        RECT 14.600 197.900 15.000 199.900 ;
        RECT 16.700 197.900 17.300 199.900 ;
        RECT 11.800 197.500 12.200 197.900 ;
        RECT 14.600 197.600 14.900 197.900 ;
        RECT 13.500 197.300 15.300 197.600 ;
        RECT 16.600 197.500 17.000 197.900 ;
        RECT 13.500 197.200 13.900 197.300 ;
        RECT 14.900 197.200 15.300 197.300 ;
        RECT 11.800 196.500 12.200 196.600 ;
        RECT 14.100 196.500 14.500 196.600 ;
        RECT 11.800 196.200 14.500 196.500 ;
        RECT 14.800 196.500 15.900 196.800 ;
        RECT 14.800 195.900 15.100 196.500 ;
        RECT 15.500 196.400 15.900 196.500 ;
        RECT 16.700 196.600 17.400 197.000 ;
        RECT 16.700 196.100 17.000 196.600 ;
        RECT 12.700 195.700 15.100 195.900 ;
        RECT 10.200 195.600 15.100 195.700 ;
        RECT 15.800 195.800 17.000 196.100 ;
        RECT 10.200 195.500 13.100 195.600 ;
        RECT 10.200 195.400 13.000 195.500 ;
        RECT 4.600 195.100 5.000 195.200 ;
        RECT 6.200 195.100 6.600 195.200 ;
        RECT 13.400 195.100 13.800 195.200 ;
        RECT 4.600 194.800 8.700 195.100 ;
        RECT 8.300 194.700 8.700 194.800 ;
        RECT 11.300 194.800 13.800 195.100 ;
        RECT 11.300 194.700 11.700 194.800 ;
        RECT 12.600 194.700 13.000 194.800 ;
        RECT 7.500 194.200 7.900 194.300 ;
        RECT 12.100 194.200 12.500 194.300 ;
        RECT 15.800 194.200 16.100 195.800 ;
        RECT 19.000 195.600 19.400 199.900 ;
        RECT 20.600 195.600 21.000 199.900 ;
        RECT 22.200 195.600 22.600 199.900 ;
        RECT 23.800 195.600 24.200 199.900 ;
        RECT 25.400 195.600 25.800 199.900 ;
        RECT 17.300 195.300 19.400 195.600 ;
        RECT 17.300 195.200 17.700 195.300 ;
        RECT 18.100 194.900 18.500 195.000 ;
        RECT 16.600 194.600 18.500 194.900 ;
        RECT 16.600 194.500 17.000 194.600 ;
        RECT 3.900 194.100 9.400 194.200 ;
        RECT 10.600 194.100 16.100 194.200 ;
        RECT 3.900 193.900 16.100 194.100 ;
        RECT 4.100 193.800 4.500 193.900 ;
        RECT 0.600 193.300 2.500 193.600 ;
        RECT 0.600 191.100 1.000 193.300 ;
        RECT 2.100 193.200 2.500 193.300 ;
        RECT 7.000 192.800 7.300 193.900 ;
        RECT 8.600 193.800 11.400 193.900 ;
        RECT 6.100 192.700 6.500 192.800 ;
        RECT 3.000 192.100 3.400 192.500 ;
        RECT 5.100 192.400 6.500 192.700 ;
        RECT 7.000 192.400 7.400 192.800 ;
        RECT 5.100 192.100 5.400 192.400 ;
        RECT 7.800 192.100 8.200 192.500 ;
        RECT 2.700 191.800 3.400 192.100 ;
        RECT 2.700 191.100 3.300 191.800 ;
        RECT 5.000 191.100 5.400 192.100 ;
        RECT 7.200 191.800 8.200 192.100 ;
        RECT 7.200 191.100 7.600 191.800 ;
        RECT 9.400 191.100 9.800 193.500 ;
        RECT 10.200 191.100 10.600 193.500 ;
        RECT 12.700 192.800 13.000 193.900 ;
        RECT 14.200 193.800 14.600 193.900 ;
        RECT 15.500 193.800 15.900 193.900 ;
        RECT 19.000 193.600 19.400 195.300 ;
        RECT 17.500 193.300 19.400 193.600 ;
        RECT 19.800 195.200 21.000 195.600 ;
        RECT 21.500 195.200 22.600 195.600 ;
        RECT 23.100 195.200 24.200 195.600 ;
        RECT 24.900 195.200 25.800 195.600 ;
        RECT 19.800 193.800 20.200 195.200 ;
        RECT 21.500 194.500 21.900 195.200 ;
        RECT 23.100 194.500 23.500 195.200 ;
        RECT 24.900 194.500 25.300 195.200 ;
        RECT 20.600 194.100 21.900 194.500 ;
        RECT 22.300 194.100 23.500 194.500 ;
        RECT 24.000 194.100 25.300 194.500 ;
        RECT 27.800 195.100 28.200 199.900 ;
        RECT 29.800 196.800 30.200 197.200 ;
        RECT 28.600 195.800 29.000 196.600 ;
        RECT 29.800 196.200 30.100 196.800 ;
        RECT 30.500 196.200 30.900 199.900 ;
        RECT 29.400 195.900 30.100 196.200 ;
        RECT 29.400 195.800 29.800 195.900 ;
        RECT 30.400 195.800 31.400 196.200 ;
        RECT 29.400 195.100 29.700 195.800 ;
        RECT 27.800 194.800 29.700 195.100 ;
        RECT 21.500 193.800 21.900 194.100 ;
        RECT 23.100 193.800 23.500 194.100 ;
        RECT 24.900 193.800 25.300 194.100 ;
        RECT 19.800 193.400 21.000 193.800 ;
        RECT 21.500 193.400 22.600 193.800 ;
        RECT 23.100 193.400 24.200 193.800 ;
        RECT 24.900 193.400 25.800 193.800 ;
        RECT 27.000 193.400 27.400 194.200 ;
        RECT 17.500 193.200 17.900 193.300 ;
        RECT 11.800 192.100 12.200 192.500 ;
        RECT 12.600 192.400 13.000 192.800 ;
        RECT 13.500 192.700 13.900 192.800 ;
        RECT 13.500 192.400 14.900 192.700 ;
        RECT 14.600 192.100 14.900 192.400 ;
        RECT 16.600 192.100 17.000 192.500 ;
        RECT 11.800 191.800 12.800 192.100 ;
        RECT 12.400 191.100 12.800 191.800 ;
        RECT 14.600 191.100 15.000 192.100 ;
        RECT 16.600 191.800 17.300 192.100 ;
        RECT 16.700 191.100 17.300 191.800 ;
        RECT 19.000 191.100 19.400 193.300 ;
        RECT 20.600 191.100 21.000 193.400 ;
        RECT 22.200 191.100 22.600 193.400 ;
        RECT 23.800 191.100 24.200 193.400 ;
        RECT 25.400 191.100 25.800 193.400 ;
        RECT 27.800 193.100 28.200 194.800 ;
        RECT 30.400 194.200 30.700 195.800 ;
        RECT 32.600 195.700 33.000 199.900 ;
        RECT 34.800 198.200 35.200 199.900 ;
        RECT 34.200 197.900 35.200 198.200 ;
        RECT 37.000 197.900 37.400 199.900 ;
        RECT 39.100 197.900 39.700 199.900 ;
        RECT 34.200 197.500 34.600 197.900 ;
        RECT 37.000 197.600 37.300 197.900 ;
        RECT 35.900 197.300 37.700 197.600 ;
        RECT 39.000 197.500 39.400 197.900 ;
        RECT 35.900 197.200 36.300 197.300 ;
        RECT 37.300 197.200 37.700 197.300 ;
        RECT 39.500 197.000 40.200 197.200 ;
        RECT 39.100 196.800 40.200 197.000 ;
        RECT 34.200 196.500 34.600 196.600 ;
        RECT 36.500 196.500 36.900 196.600 ;
        RECT 34.200 196.200 36.900 196.500 ;
        RECT 37.200 196.500 38.300 196.800 ;
        RECT 37.200 195.900 37.500 196.500 ;
        RECT 37.900 196.400 38.300 196.500 ;
        RECT 39.100 196.600 39.800 196.800 ;
        RECT 39.100 196.100 39.400 196.600 ;
        RECT 35.100 195.700 37.500 195.900 ;
        RECT 32.600 195.600 37.500 195.700 ;
        RECT 38.200 195.800 39.400 196.100 ;
        RECT 32.600 195.500 35.500 195.600 ;
        RECT 32.600 195.400 35.400 195.500 ;
        RECT 31.000 194.400 31.400 195.200 ;
        RECT 35.800 195.100 36.200 195.200 ;
        RECT 33.700 194.800 36.200 195.100 ;
        RECT 33.700 194.700 34.100 194.800 ;
        RECT 35.000 194.700 35.400 194.800 ;
        RECT 34.500 194.200 34.900 194.300 ;
        RECT 38.200 194.200 38.500 195.800 ;
        RECT 41.400 195.600 41.800 199.900 ;
        RECT 43.000 196.400 43.400 199.900 ;
        RECT 39.700 195.300 41.800 195.600 ;
        RECT 39.700 195.200 40.100 195.300 ;
        RECT 40.500 194.900 40.900 195.000 ;
        RECT 39.000 194.600 40.900 194.900 ;
        RECT 39.000 194.500 39.400 194.600 ;
        RECT 29.400 193.800 30.700 194.200 ;
        RECT 31.800 194.100 32.200 194.200 ;
        RECT 31.400 193.800 32.200 194.100 ;
        RECT 33.000 193.900 38.500 194.200 ;
        RECT 33.000 193.800 33.800 193.900 ;
        RECT 29.500 193.100 29.800 193.800 ;
        RECT 31.400 193.600 31.800 193.800 ;
        RECT 30.300 193.100 32.100 193.300 ;
        RECT 27.800 192.800 28.700 193.100 ;
        RECT 28.300 191.100 28.700 192.800 ;
        RECT 29.400 191.100 29.800 193.100 ;
        RECT 30.200 193.000 32.200 193.100 ;
        RECT 30.200 191.100 30.600 193.000 ;
        RECT 31.800 191.100 32.200 193.000 ;
        RECT 32.600 191.100 33.000 193.500 ;
        RECT 35.100 192.800 35.400 193.900 ;
        RECT 37.900 193.800 38.300 193.900 ;
        RECT 41.400 193.600 41.800 195.300 ;
        RECT 39.900 193.300 41.800 193.600 ;
        RECT 39.900 193.200 40.300 193.300 ;
        RECT 34.200 192.100 34.600 192.500 ;
        RECT 35.000 192.400 35.400 192.800 ;
        RECT 35.900 192.700 36.300 192.800 ;
        RECT 35.900 192.400 37.300 192.700 ;
        RECT 37.000 192.100 37.300 192.400 ;
        RECT 39.000 192.100 39.400 192.500 ;
        RECT 34.200 191.800 35.200 192.100 ;
        RECT 34.800 191.100 35.200 191.800 ;
        RECT 37.000 191.100 37.400 192.100 ;
        RECT 39.000 191.800 39.700 192.100 ;
        RECT 39.100 191.100 39.700 191.800 ;
        RECT 41.400 191.100 41.800 193.300 ;
        RECT 42.900 195.900 43.400 196.400 ;
        RECT 44.600 196.200 45.000 199.900 ;
        RECT 43.700 195.900 45.000 196.200 ;
        RECT 45.400 197.500 45.800 199.500 ;
        RECT 42.900 194.200 43.200 195.900 ;
        RECT 43.700 194.900 44.000 195.900 ;
        RECT 45.400 195.800 45.700 197.500 ;
        RECT 47.500 196.400 47.900 199.900 ;
        RECT 51.800 197.500 52.200 199.500 ;
        RECT 47.500 196.100 48.300 196.400 ;
        RECT 45.400 195.500 47.300 195.800 ;
        RECT 43.500 194.500 44.000 194.900 ;
        RECT 42.900 193.800 43.400 194.200 ;
        RECT 42.900 193.100 43.200 193.800 ;
        RECT 43.700 193.700 44.000 194.500 ;
        RECT 44.500 194.800 45.000 195.200 ;
        RECT 44.500 194.400 44.900 194.800 ;
        RECT 45.400 194.400 45.800 195.200 ;
        RECT 46.200 194.400 46.600 195.200 ;
        RECT 47.000 194.500 47.300 195.500 ;
        RECT 47.000 194.100 47.700 194.500 ;
        RECT 48.000 194.200 48.300 196.100 ;
        RECT 51.800 195.800 52.100 197.500 ;
        RECT 53.900 196.400 54.300 199.900 ;
        RECT 53.900 196.100 54.700 196.400 ;
        RECT 48.600 194.800 49.000 195.600 ;
        RECT 51.800 195.500 53.700 195.800 ;
        RECT 51.800 194.400 52.200 195.200 ;
        RECT 52.600 194.400 53.000 195.200 ;
        RECT 53.400 194.500 53.700 195.500 ;
        RECT 48.000 194.100 49.000 194.200 ;
        RECT 51.000 194.100 51.400 194.200 ;
        RECT 47.000 193.900 47.500 194.100 ;
        RECT 43.700 193.400 45.000 193.700 ;
        RECT 42.900 192.800 43.400 193.100 ;
        RECT 43.000 191.100 43.400 192.800 ;
        RECT 44.600 191.100 45.000 193.400 ;
        RECT 45.400 193.600 47.500 193.900 ;
        RECT 48.000 193.800 51.400 194.100 ;
        RECT 53.400 194.100 54.100 194.500 ;
        RECT 54.400 194.200 54.700 196.100 ;
        RECT 55.000 194.800 55.400 195.600 ;
        RECT 57.400 195.100 57.800 199.900 ;
        RECT 59.400 196.800 59.800 197.200 ;
        RECT 58.200 195.800 58.600 196.600 ;
        RECT 59.400 196.200 59.700 196.800 ;
        RECT 60.100 196.200 60.500 199.900 ;
        RECT 63.500 199.200 63.900 199.900 ;
        RECT 63.000 198.800 63.900 199.200 ;
        RECT 59.000 195.900 59.700 196.200 ;
        RECT 60.000 195.900 60.500 196.200 ;
        RECT 63.500 196.200 63.900 198.800 ;
        RECT 64.200 196.800 64.600 197.200 ;
        RECT 64.300 196.200 64.600 196.800 ;
        RECT 65.400 196.200 65.800 199.900 ;
        RECT 67.000 199.600 69.000 199.900 ;
        RECT 67.000 196.200 67.400 199.600 ;
        RECT 63.500 195.900 64.000 196.200 ;
        RECT 64.300 195.900 65.000 196.200 ;
        RECT 65.400 195.900 67.400 196.200 ;
        RECT 59.000 195.800 59.400 195.900 ;
        RECT 59.000 195.100 59.300 195.800 ;
        RECT 57.400 194.800 59.300 195.100 ;
        RECT 53.400 193.900 53.900 194.100 ;
        RECT 45.400 192.500 45.700 193.600 ;
        RECT 48.000 193.500 48.300 193.800 ;
        RECT 47.900 193.300 48.300 193.500 ;
        RECT 47.500 193.000 48.300 193.300 ;
        RECT 51.800 193.600 53.900 193.900 ;
        RECT 54.400 193.800 55.400 194.200 ;
        RECT 55.800 194.100 56.200 194.200 ;
        RECT 56.600 194.100 57.000 194.200 ;
        RECT 55.800 193.800 57.000 194.100 ;
        RECT 45.400 191.500 45.800 192.500 ;
        RECT 47.500 191.500 47.900 193.000 ;
        RECT 51.800 192.500 52.100 193.600 ;
        RECT 54.400 193.500 54.700 193.800 ;
        RECT 54.300 193.300 54.700 193.500 ;
        RECT 56.600 193.400 57.000 193.800 ;
        RECT 53.900 193.000 54.700 193.300 ;
        RECT 57.400 193.100 57.800 194.800 ;
        RECT 60.000 194.200 60.300 195.900 ;
        RECT 60.600 194.400 61.000 195.200 ;
        RECT 63.000 194.400 63.400 195.200 ;
        RECT 63.700 194.200 64.000 195.900 ;
        RECT 64.600 195.800 65.000 195.900 ;
        RECT 67.800 195.800 68.200 199.300 ;
        RECT 68.600 195.900 69.000 199.600 ;
        RECT 69.400 195.800 69.800 196.600 ;
        RECT 67.800 195.600 68.100 195.800 ;
        RECT 65.800 195.200 66.200 195.400 ;
        RECT 67.100 195.300 68.100 195.600 ;
        RECT 67.100 195.200 67.400 195.300 ;
        RECT 64.600 195.100 65.000 195.200 ;
        RECT 65.400 195.100 66.200 195.200 ;
        RECT 64.600 194.900 66.200 195.100 ;
        RECT 64.600 194.800 65.800 194.900 ;
        RECT 67.000 194.800 67.400 195.200 ;
        RECT 68.600 194.800 69.000 195.600 ;
        RECT 69.400 195.100 69.800 195.200 ;
        RECT 70.200 195.100 70.600 199.900 ;
        RECT 72.600 196.400 73.000 199.900 ;
        RECT 69.400 194.800 70.600 195.100 ;
        RECT 59.000 193.800 60.300 194.200 ;
        RECT 61.400 194.100 61.800 194.200 ;
        RECT 61.000 193.800 61.800 194.100 ;
        RECT 62.200 194.100 62.600 194.200 ;
        RECT 62.200 193.800 63.000 194.100 ;
        RECT 63.700 193.800 65.000 194.200 ;
        RECT 65.400 194.100 65.800 194.200 ;
        RECT 66.200 194.100 66.600 194.600 ;
        RECT 65.400 193.800 66.600 194.100 ;
        RECT 59.100 193.100 59.400 193.800 ;
        RECT 61.000 193.600 61.400 193.800 ;
        RECT 62.600 193.600 63.000 193.800 ;
        RECT 59.900 193.100 61.700 193.300 ;
        RECT 62.300 193.100 64.100 193.300 ;
        RECT 64.600 193.100 64.900 193.800 ;
        RECT 67.100 193.100 67.400 194.800 ;
        RECT 67.700 194.400 68.100 194.800 ;
        RECT 67.800 194.200 68.100 194.400 ;
        RECT 67.800 193.800 68.200 194.200 ;
        RECT 70.200 193.100 70.600 194.800 ;
        RECT 72.500 195.900 73.000 196.400 ;
        RECT 74.200 196.200 74.600 199.900 ;
        RECT 73.300 195.900 74.600 196.200 ;
        RECT 75.000 196.200 75.400 199.900 ;
        RECT 76.600 196.400 77.000 199.900 ;
        RECT 79.300 199.200 79.700 199.900 ;
        RECT 79.300 198.800 80.200 199.200 ;
        RECT 78.600 196.800 79.000 197.200 ;
        RECT 75.000 195.900 76.300 196.200 ;
        RECT 76.600 195.900 77.100 196.400 ;
        RECT 78.600 196.200 78.900 196.800 ;
        RECT 79.300 196.200 79.700 198.800 ;
        RECT 72.500 194.200 72.800 195.900 ;
        RECT 73.300 194.900 73.600 195.900 ;
        RECT 73.100 194.500 73.600 194.900 ;
        RECT 71.000 194.100 71.400 194.200 ;
        RECT 71.800 194.100 72.200 194.200 ;
        RECT 71.000 193.800 72.200 194.100 ;
        RECT 72.500 193.800 73.000 194.200 ;
        RECT 71.000 193.400 71.400 193.800 ;
        RECT 51.800 191.500 52.200 192.500 ;
        RECT 53.900 192.200 54.300 193.000 ;
        RECT 57.400 192.800 58.300 193.100 ;
        RECT 53.900 191.800 54.600 192.200 ;
        RECT 53.900 191.500 54.300 191.800 ;
        RECT 57.900 191.100 58.300 192.800 ;
        RECT 59.000 191.100 59.400 193.100 ;
        RECT 59.800 193.000 61.800 193.100 ;
        RECT 59.800 191.100 60.200 193.000 ;
        RECT 61.400 191.100 61.800 193.000 ;
        RECT 62.200 193.000 64.200 193.100 ;
        RECT 62.200 191.100 62.600 193.000 ;
        RECT 63.800 191.100 64.200 193.000 ;
        RECT 64.600 191.100 65.000 193.100 ;
        RECT 66.900 191.100 67.700 193.100 ;
        RECT 69.700 192.800 70.600 193.100 ;
        RECT 72.500 193.200 72.800 193.800 ;
        RECT 73.300 193.700 73.600 194.500 ;
        RECT 74.100 195.100 74.600 195.200 ;
        RECT 75.000 195.100 75.500 195.200 ;
        RECT 74.100 194.800 75.500 195.100 ;
        RECT 74.100 194.400 74.500 194.800 ;
        RECT 75.100 194.400 75.500 194.800 ;
        RECT 76.000 194.900 76.300 195.900 ;
        RECT 76.000 194.500 76.500 194.900 ;
        RECT 76.000 193.700 76.300 194.500 ;
        RECT 76.800 194.200 77.100 195.900 ;
        RECT 78.200 195.900 78.900 196.200 ;
        RECT 79.200 195.900 79.700 196.200 ;
        RECT 78.200 195.800 78.600 195.900 ;
        RECT 76.600 194.100 77.100 194.200 ;
        RECT 77.400 194.800 77.800 195.200 ;
        RECT 77.400 194.100 77.700 194.800 ;
        RECT 79.200 194.200 79.500 195.900 ;
        RECT 81.400 195.600 81.800 199.900 ;
        RECT 83.500 197.900 84.100 199.900 ;
        RECT 85.800 197.900 86.200 199.900 ;
        RECT 88.000 198.200 88.400 199.900 ;
        RECT 88.000 197.900 89.000 198.200 ;
        RECT 83.800 197.500 84.200 197.900 ;
        RECT 85.900 197.600 86.200 197.900 ;
        RECT 85.500 197.300 87.300 197.600 ;
        RECT 88.600 197.500 89.000 197.900 ;
        RECT 85.500 197.200 85.900 197.300 ;
        RECT 86.900 197.200 87.300 197.300 ;
        RECT 83.000 197.000 83.700 197.200 ;
        RECT 83.000 196.800 84.100 197.000 ;
        RECT 83.400 196.600 84.100 196.800 ;
        RECT 83.800 196.100 84.100 196.600 ;
        RECT 84.900 196.500 86.000 196.800 ;
        RECT 84.900 196.400 85.300 196.500 ;
        RECT 83.800 195.800 85.000 196.100 ;
        RECT 81.400 195.300 83.500 195.600 ;
        RECT 79.800 194.400 80.200 195.200 ;
        RECT 76.600 193.800 77.700 194.100 ;
        RECT 78.200 193.800 79.500 194.200 ;
        RECT 80.600 194.100 81.000 194.200 ;
        RECT 80.200 193.800 81.000 194.100 ;
        RECT 73.300 193.400 74.600 193.700 ;
        RECT 72.500 192.800 73.000 193.200 ;
        RECT 69.700 191.100 70.100 192.800 ;
        RECT 72.600 191.100 73.000 192.800 ;
        RECT 74.200 191.100 74.600 193.400 ;
        RECT 75.000 193.400 76.300 193.700 ;
        RECT 75.000 191.100 75.400 193.400 ;
        RECT 76.800 193.100 77.100 193.800 ;
        RECT 78.300 193.100 78.600 193.800 ;
        RECT 80.200 193.600 80.600 193.800 ;
        RECT 81.400 193.600 81.800 195.300 ;
        RECT 83.100 195.200 83.500 195.300 ;
        RECT 82.300 194.900 82.700 195.000 ;
        RECT 82.300 194.600 84.200 194.900 ;
        RECT 83.800 194.500 84.200 194.600 ;
        RECT 84.700 194.200 85.000 195.800 ;
        RECT 85.700 195.900 86.000 196.500 ;
        RECT 86.300 196.500 86.700 196.600 ;
        RECT 88.600 196.500 89.000 196.600 ;
        RECT 86.300 196.200 89.000 196.500 ;
        RECT 85.700 195.700 88.100 195.900 ;
        RECT 90.200 195.700 90.600 199.900 ;
        RECT 92.900 196.400 93.300 199.900 ;
        RECT 95.000 197.500 95.400 199.500 ;
        RECT 85.700 195.600 90.600 195.700 ;
        RECT 92.500 196.100 93.300 196.400 ;
        RECT 87.700 195.500 90.600 195.600 ;
        RECT 87.800 195.400 90.600 195.500 ;
        RECT 87.000 195.100 87.400 195.200 ;
        RECT 87.000 194.800 89.500 195.100 ;
        RECT 91.800 194.800 92.200 195.600 ;
        RECT 87.800 194.700 88.200 194.800 ;
        RECT 89.100 194.700 89.500 194.800 ;
        RECT 88.300 194.200 88.700 194.300 ;
        RECT 92.500 194.200 92.800 196.100 ;
        RECT 95.100 195.800 95.400 197.500 ;
        RECT 97.100 196.200 97.500 199.900 ;
        RECT 97.800 196.800 98.200 197.200 ;
        RECT 97.900 196.200 98.200 196.800 ;
        RECT 97.100 195.900 97.600 196.200 ;
        RECT 97.900 196.100 98.600 196.200 ;
        RECT 99.000 196.100 99.400 196.200 ;
        RECT 97.900 195.900 99.400 196.100 ;
        RECT 93.500 195.500 95.400 195.800 ;
        RECT 93.500 194.500 93.800 195.500 ;
        RECT 84.700 193.900 90.200 194.200 ;
        RECT 84.900 193.800 85.300 193.900 ;
        RECT 81.400 193.300 83.300 193.600 ;
        RECT 79.100 193.100 80.900 193.300 ;
        RECT 76.600 192.800 77.100 193.100 ;
        RECT 76.600 191.100 77.000 192.800 ;
        RECT 78.200 191.100 78.600 193.100 ;
        RECT 79.000 193.000 81.000 193.100 ;
        RECT 79.000 191.100 79.400 193.000 ;
        RECT 80.600 191.100 81.000 193.000 ;
        RECT 81.400 191.100 81.800 193.300 ;
        RECT 82.900 193.200 83.300 193.300 ;
        RECT 87.800 192.800 88.100 193.900 ;
        RECT 89.400 193.800 90.200 193.900 ;
        RECT 91.800 193.800 92.800 194.200 ;
        RECT 93.100 194.100 93.800 194.500 ;
        RECT 94.200 194.400 94.600 195.200 ;
        RECT 95.000 194.400 95.400 195.200 ;
        RECT 96.600 194.400 97.000 195.200 ;
        RECT 97.300 195.100 97.600 195.900 ;
        RECT 98.200 195.800 99.400 195.900 ;
        RECT 100.600 195.800 101.000 196.600 ;
        RECT 99.800 195.100 100.200 195.200 ;
        RECT 97.300 194.800 100.200 195.100 ;
        RECT 97.300 194.200 97.600 194.800 ;
        RECT 92.500 193.500 92.800 193.800 ;
        RECT 93.300 193.900 93.800 194.100 ;
        RECT 95.800 194.100 96.200 194.200 ;
        RECT 93.300 193.600 95.400 193.900 ;
        RECT 95.800 193.800 96.600 194.100 ;
        RECT 97.300 193.800 98.600 194.200 ;
        RECT 99.000 194.100 99.400 194.200 ;
        RECT 101.400 194.100 101.800 199.900 ;
        RECT 103.000 195.600 103.400 199.900 ;
        RECT 105.100 197.900 105.700 199.900 ;
        RECT 107.400 197.900 107.800 199.900 ;
        RECT 109.600 198.200 110.000 199.900 ;
        RECT 109.600 197.900 110.600 198.200 ;
        RECT 105.400 197.500 105.800 197.900 ;
        RECT 107.500 197.600 107.800 197.900 ;
        RECT 107.100 197.300 108.900 197.600 ;
        RECT 110.200 197.500 110.600 197.900 ;
        RECT 107.100 197.200 107.500 197.300 ;
        RECT 108.500 197.200 108.900 197.300 ;
        RECT 105.000 196.600 105.700 197.000 ;
        RECT 105.400 196.100 105.700 196.600 ;
        RECT 106.500 196.500 107.600 196.800 ;
        RECT 106.500 196.400 106.900 196.500 ;
        RECT 105.400 195.800 106.600 196.100 ;
        RECT 103.000 195.300 105.100 195.600 ;
        RECT 99.000 193.800 101.800 194.100 ;
        RECT 96.200 193.600 96.600 193.800 ;
        RECT 86.900 192.700 87.300 192.800 ;
        RECT 83.800 192.100 84.200 192.500 ;
        RECT 85.900 192.400 87.300 192.700 ;
        RECT 87.800 192.400 88.200 192.800 ;
        RECT 85.900 192.100 86.200 192.400 ;
        RECT 88.600 192.100 89.000 192.500 ;
        RECT 83.500 191.800 84.200 192.100 ;
        RECT 83.500 191.100 84.100 191.800 ;
        RECT 85.800 191.100 86.200 192.100 ;
        RECT 88.000 191.800 89.000 192.100 ;
        RECT 88.000 191.100 88.400 191.800 ;
        RECT 90.200 191.100 90.600 193.500 ;
        RECT 92.500 193.300 92.900 193.500 ;
        RECT 92.500 193.000 93.300 193.300 ;
        RECT 92.900 192.200 93.300 193.000 ;
        RECT 95.100 192.500 95.400 193.600 ;
        RECT 95.900 193.100 97.700 193.300 ;
        RECT 98.200 193.100 98.500 193.800 ;
        RECT 101.400 193.100 101.800 193.800 ;
        RECT 102.200 194.100 102.600 194.200 ;
        RECT 103.000 194.100 103.400 195.300 ;
        RECT 104.700 195.200 105.100 195.300 ;
        RECT 103.900 194.900 104.300 195.000 ;
        RECT 103.900 194.600 105.800 194.900 ;
        RECT 105.400 194.500 105.800 194.600 ;
        RECT 106.300 194.200 106.600 195.800 ;
        RECT 107.300 195.900 107.600 196.500 ;
        RECT 107.900 196.500 108.300 196.600 ;
        RECT 110.200 196.500 110.600 196.600 ;
        RECT 107.900 196.200 110.600 196.500 ;
        RECT 107.300 195.700 109.700 195.900 ;
        RECT 111.800 195.700 112.200 199.900 ;
        RECT 114.500 196.400 114.900 199.900 ;
        RECT 116.600 197.500 117.000 199.500 ;
        RECT 107.300 195.600 112.200 195.700 ;
        RECT 114.100 196.100 114.900 196.400 ;
        RECT 109.300 195.500 112.200 195.600 ;
        RECT 109.400 195.400 112.200 195.500 ;
        RECT 108.600 195.100 109.000 195.200 ;
        RECT 108.600 194.800 111.100 195.100 ;
        RECT 113.400 194.800 113.800 195.600 ;
        RECT 110.700 194.700 111.100 194.800 ;
        RECT 109.900 194.200 110.300 194.300 ;
        RECT 114.100 194.200 114.400 196.100 ;
        RECT 116.700 195.800 117.000 197.500 ;
        RECT 115.100 195.500 117.000 195.800 ;
        RECT 117.400 195.600 117.800 199.900 ;
        RECT 119.500 197.900 120.100 199.900 ;
        RECT 121.800 197.900 122.200 199.900 ;
        RECT 124.000 198.200 124.400 199.900 ;
        RECT 124.000 197.900 125.000 198.200 ;
        RECT 119.800 197.500 120.200 197.900 ;
        RECT 121.900 197.600 122.200 197.900 ;
        RECT 121.500 197.300 123.300 197.600 ;
        RECT 124.600 197.500 125.000 197.900 ;
        RECT 121.500 197.200 121.900 197.300 ;
        RECT 122.900 197.200 123.300 197.300 ;
        RECT 119.400 196.600 120.100 197.000 ;
        RECT 119.800 196.100 120.100 196.600 ;
        RECT 120.900 196.500 122.000 196.800 ;
        RECT 120.900 196.400 121.300 196.500 ;
        RECT 119.800 195.800 121.000 196.100 ;
        RECT 115.100 194.500 115.400 195.500 ;
        RECT 117.400 195.300 119.500 195.600 ;
        RECT 102.200 193.800 103.400 194.100 ;
        RECT 102.200 193.400 102.600 193.800 ;
        RECT 103.000 193.600 103.400 193.800 ;
        RECT 106.200 193.900 111.800 194.200 ;
        RECT 106.200 193.800 106.900 193.900 ;
        RECT 92.600 191.800 93.300 192.200 ;
        RECT 92.900 191.500 93.300 191.800 ;
        RECT 95.000 191.500 95.400 192.500 ;
        RECT 95.800 193.000 97.800 193.100 ;
        RECT 95.800 191.100 96.200 193.000 ;
        RECT 97.400 191.100 97.800 193.000 ;
        RECT 98.200 191.100 98.600 193.100 ;
        RECT 100.900 192.800 101.800 193.100 ;
        RECT 103.000 193.300 104.900 193.600 ;
        RECT 100.900 191.100 101.300 192.800 ;
        RECT 103.000 191.100 103.400 193.300 ;
        RECT 104.500 193.200 104.900 193.300 ;
        RECT 106.200 193.200 106.500 193.800 ;
        RECT 106.200 192.800 106.600 193.200 ;
        RECT 109.400 192.800 109.700 193.900 ;
        RECT 111.000 193.800 111.800 193.900 ;
        RECT 113.400 193.800 114.400 194.200 ;
        RECT 114.700 194.100 115.400 194.500 ;
        RECT 115.800 194.400 116.200 195.200 ;
        RECT 116.600 194.400 117.000 195.200 ;
        RECT 114.100 193.500 114.400 193.800 ;
        RECT 114.900 193.900 115.400 194.100 ;
        RECT 114.900 193.600 117.000 193.900 ;
        RECT 108.500 192.700 108.900 192.800 ;
        RECT 105.400 192.100 105.800 192.500 ;
        RECT 107.500 192.400 108.900 192.700 ;
        RECT 109.400 192.400 109.800 192.800 ;
        RECT 107.500 192.100 107.800 192.400 ;
        RECT 110.200 192.100 110.600 192.500 ;
        RECT 105.100 191.800 105.800 192.100 ;
        RECT 105.100 191.100 105.700 191.800 ;
        RECT 107.400 191.100 107.800 192.100 ;
        RECT 109.600 191.800 110.600 192.100 ;
        RECT 109.600 191.100 110.000 191.800 ;
        RECT 111.800 191.100 112.200 193.500 ;
        RECT 114.100 193.300 114.500 193.500 ;
        RECT 114.100 193.200 114.900 193.300 ;
        RECT 114.100 193.000 115.400 193.200 ;
        RECT 114.500 192.800 115.400 193.000 ;
        RECT 114.500 191.500 114.900 192.800 ;
        RECT 116.700 192.500 117.000 193.600 ;
        RECT 116.600 191.500 117.000 192.500 ;
        RECT 117.400 193.600 117.800 195.300 ;
        RECT 119.100 195.200 119.500 195.300 ;
        RECT 120.700 195.200 121.000 195.800 ;
        RECT 121.700 195.900 122.000 196.500 ;
        RECT 122.300 196.500 122.700 196.600 ;
        RECT 124.600 196.500 125.000 196.600 ;
        RECT 122.300 196.200 125.000 196.500 ;
        RECT 121.700 195.700 124.100 195.900 ;
        RECT 126.200 195.700 126.600 199.900 ;
        RECT 128.900 196.400 129.300 199.900 ;
        RECT 131.000 197.500 131.400 199.500 ;
        RECT 121.700 195.600 126.600 195.700 ;
        RECT 128.500 196.100 129.300 196.400 ;
        RECT 123.700 195.500 126.600 195.600 ;
        RECT 123.800 195.400 126.600 195.500 ;
        RECT 118.300 194.900 118.700 195.000 ;
        RECT 118.300 194.600 120.200 194.900 ;
        RECT 120.600 194.800 121.000 195.200 ;
        RECT 123.000 195.100 123.400 195.200 ;
        RECT 123.000 194.800 125.500 195.100 ;
        RECT 127.800 194.800 128.200 195.600 ;
        RECT 119.800 194.500 120.200 194.600 ;
        RECT 120.700 194.200 121.000 194.800 ;
        RECT 123.800 194.700 124.200 194.800 ;
        RECT 125.100 194.700 125.500 194.800 ;
        RECT 124.300 194.200 124.700 194.300 ;
        RECT 128.500 194.200 128.800 196.100 ;
        RECT 131.100 195.800 131.400 197.500 ;
        RECT 133.700 196.400 134.100 199.900 ;
        RECT 135.800 197.500 136.200 199.500 ;
        RECT 129.500 195.500 131.400 195.800 ;
        RECT 133.300 196.100 134.100 196.400 ;
        RECT 129.500 194.500 129.800 195.500 ;
        RECT 120.700 194.100 126.200 194.200 ;
        RECT 127.000 194.100 127.400 194.200 ;
        RECT 120.700 193.900 127.400 194.100 ;
        RECT 120.900 193.800 121.300 193.900 ;
        RECT 117.400 193.300 119.300 193.600 ;
        RECT 117.400 191.100 117.800 193.300 ;
        RECT 118.900 193.200 119.300 193.300 ;
        RECT 123.800 192.800 124.100 193.900 ;
        RECT 125.400 193.800 127.400 193.900 ;
        RECT 127.800 193.800 128.800 194.200 ;
        RECT 129.100 194.100 129.800 194.500 ;
        RECT 130.200 194.400 130.600 195.200 ;
        RECT 131.000 194.400 131.400 195.200 ;
        RECT 132.600 194.800 133.000 195.600 ;
        RECT 133.300 194.200 133.600 196.100 ;
        RECT 135.900 195.800 136.200 197.500 ;
        RECT 136.600 196.200 137.000 199.900 ;
        RECT 138.200 199.600 140.200 199.900 ;
        RECT 138.200 196.200 138.600 199.600 ;
        RECT 136.600 195.900 138.600 196.200 ;
        RECT 139.000 195.900 139.400 199.300 ;
        RECT 139.800 195.900 140.200 199.600 ;
        RECT 142.500 196.400 142.900 199.900 ;
        RECT 144.600 197.500 145.000 199.500 ;
        RECT 142.100 196.100 142.900 196.400 ;
        RECT 134.300 195.500 136.200 195.800 ;
        RECT 139.000 195.600 139.300 195.900 ;
        RECT 134.300 194.500 134.600 195.500 ;
        RECT 137.000 195.200 137.400 195.400 ;
        RECT 138.300 195.300 139.300 195.600 ;
        RECT 138.300 195.200 138.600 195.300 ;
        RECT 128.500 193.500 128.800 193.800 ;
        RECT 129.300 193.900 129.800 194.100 ;
        RECT 131.800 194.100 132.200 194.200 ;
        RECT 132.600 194.100 133.600 194.200 ;
        RECT 133.900 194.100 134.600 194.500 ;
        RECT 135.000 194.400 135.400 195.200 ;
        RECT 135.800 194.400 136.200 195.200 ;
        RECT 136.600 194.900 137.400 195.200 ;
        RECT 136.600 194.800 137.000 194.900 ;
        RECT 138.200 194.800 138.600 195.200 ;
        RECT 139.800 194.800 140.200 195.600 ;
        RECT 141.400 194.800 141.800 195.600 ;
        RECT 129.300 193.600 131.400 193.900 ;
        RECT 131.800 193.800 133.600 194.100 ;
        RECT 122.900 192.700 123.300 192.800 ;
        RECT 119.800 192.100 120.200 192.500 ;
        RECT 121.900 192.400 123.300 192.700 ;
        RECT 123.800 192.400 124.200 192.800 ;
        RECT 121.900 192.100 122.200 192.400 ;
        RECT 124.600 192.100 125.000 192.500 ;
        RECT 119.500 191.800 120.200 192.100 ;
        RECT 119.500 191.100 120.100 191.800 ;
        RECT 121.800 191.100 122.200 192.100 ;
        RECT 124.000 191.800 125.000 192.100 ;
        RECT 124.000 191.100 124.400 191.800 ;
        RECT 126.200 191.100 126.600 193.500 ;
        RECT 128.500 193.300 128.900 193.500 ;
        RECT 128.500 193.000 129.300 193.300 ;
        RECT 128.900 192.200 129.300 193.000 ;
        RECT 131.100 192.500 131.400 193.600 ;
        RECT 133.300 193.500 133.600 193.800 ;
        RECT 134.100 193.900 134.600 194.100 ;
        RECT 134.100 193.600 136.200 193.900 ;
        RECT 137.400 193.800 137.800 194.600 ;
        RECT 133.300 193.300 133.700 193.500 ;
        RECT 133.300 193.000 134.100 193.300 ;
        RECT 128.900 191.800 129.800 192.200 ;
        RECT 128.900 191.500 129.300 191.800 ;
        RECT 131.000 191.500 131.400 192.500 ;
        RECT 133.700 191.500 134.100 193.000 ;
        RECT 135.900 192.500 136.200 193.600 ;
        RECT 138.300 193.100 138.600 194.800 ;
        RECT 138.900 194.400 139.300 194.800 ;
        RECT 139.000 194.200 139.300 194.400 ;
        RECT 142.100 194.200 142.400 196.100 ;
        RECT 144.700 195.800 145.000 197.500 ;
        RECT 146.700 196.200 147.100 199.900 ;
        RECT 147.400 196.800 147.800 197.200 ;
        RECT 147.500 196.200 147.800 196.800 ;
        RECT 146.700 195.900 147.200 196.200 ;
        RECT 147.500 195.900 148.200 196.200 ;
        RECT 143.100 195.500 145.000 195.800 ;
        RECT 143.100 194.500 143.400 195.500 ;
        RECT 139.000 194.100 139.400 194.200 ;
        RECT 141.400 194.100 142.400 194.200 ;
        RECT 142.700 194.100 143.400 194.500 ;
        RECT 143.800 194.400 144.200 195.200 ;
        RECT 144.600 194.400 145.000 195.200 ;
        RECT 146.200 194.400 146.600 195.200 ;
        RECT 146.900 194.200 147.200 195.900 ;
        RECT 147.800 195.800 148.200 195.900 ;
        RECT 150.200 195.700 150.600 199.900 ;
        RECT 152.400 198.200 152.800 199.900 ;
        RECT 151.800 197.900 152.800 198.200 ;
        RECT 154.600 197.900 155.000 199.900 ;
        RECT 156.700 197.900 157.300 199.900 ;
        RECT 151.800 197.500 152.200 197.900 ;
        RECT 154.600 197.600 154.900 197.900 ;
        RECT 153.500 197.300 155.300 197.600 ;
        RECT 156.600 197.500 157.000 197.900 ;
        RECT 153.500 197.200 153.900 197.300 ;
        RECT 154.900 197.200 155.300 197.300 ;
        RECT 151.800 196.500 152.200 196.600 ;
        RECT 154.100 196.500 154.500 196.600 ;
        RECT 151.800 196.200 154.500 196.500 ;
        RECT 154.800 196.500 155.900 196.800 ;
        RECT 154.800 195.900 155.100 196.500 ;
        RECT 155.500 196.400 155.900 196.500 ;
        RECT 156.700 196.600 157.400 197.000 ;
        RECT 156.700 196.100 157.000 196.600 ;
        RECT 152.700 195.700 155.100 195.900 ;
        RECT 150.200 195.600 155.100 195.700 ;
        RECT 155.800 195.800 157.000 196.100 ;
        RECT 150.200 195.500 153.100 195.600 ;
        RECT 150.200 195.400 153.000 195.500 ;
        RECT 153.400 195.100 153.800 195.200 ;
        RECT 151.300 194.800 153.800 195.100 ;
        RECT 151.300 194.700 151.700 194.800 ;
        RECT 152.600 194.700 153.000 194.800 ;
        RECT 152.100 194.200 152.500 194.300 ;
        RECT 155.800 194.200 156.100 195.800 ;
        RECT 159.000 195.600 159.400 199.900 ;
        RECT 157.300 195.300 159.400 195.600 ;
        RECT 157.300 195.200 157.700 195.300 ;
        RECT 158.100 194.900 158.500 195.000 ;
        RECT 156.600 194.600 158.500 194.900 ;
        RECT 156.600 194.500 157.000 194.600 ;
        RECT 139.000 193.800 142.400 194.100 ;
        RECT 142.100 193.500 142.400 193.800 ;
        RECT 142.900 193.900 143.400 194.100 ;
        RECT 145.400 194.100 145.800 194.200 ;
        RECT 146.900 194.100 148.200 194.200 ;
        RECT 148.600 194.100 149.000 194.200 ;
        RECT 142.900 193.600 145.000 193.900 ;
        RECT 145.400 193.800 146.200 194.100 ;
        RECT 146.900 193.800 149.000 194.100 ;
        RECT 150.600 193.900 156.200 194.200 ;
        RECT 150.600 193.800 151.400 193.900 ;
        RECT 145.800 193.600 146.200 193.800 ;
        RECT 142.100 193.300 142.500 193.500 ;
        RECT 135.800 191.500 136.200 192.500 ;
        RECT 138.100 192.200 138.900 193.100 ;
        RECT 142.100 193.000 142.900 193.300 ;
        RECT 138.100 191.800 139.400 192.200 ;
        RECT 138.100 191.100 138.900 191.800 ;
        RECT 142.500 191.500 142.900 193.000 ;
        RECT 144.700 192.500 145.000 193.600 ;
        RECT 145.500 193.100 147.300 193.300 ;
        RECT 147.800 193.100 148.100 193.800 ;
        RECT 144.600 191.500 145.000 192.500 ;
        RECT 145.400 193.000 147.400 193.100 ;
        RECT 145.400 191.100 145.800 193.000 ;
        RECT 147.000 191.100 147.400 193.000 ;
        RECT 147.800 191.100 148.200 193.100 ;
        RECT 150.200 191.100 150.600 193.500 ;
        RECT 152.700 192.800 153.000 193.900 ;
        RECT 153.400 193.800 153.800 193.900 ;
        RECT 155.500 193.800 156.200 193.900 ;
        RECT 159.000 193.600 159.400 195.300 ;
        RECT 157.500 193.300 159.400 193.600 ;
        RECT 157.500 193.200 157.900 193.300 ;
        RECT 151.800 192.100 152.200 192.500 ;
        RECT 152.600 192.400 153.000 192.800 ;
        RECT 153.500 192.700 153.900 192.800 ;
        RECT 153.500 192.400 154.900 192.700 ;
        RECT 154.600 192.100 154.900 192.400 ;
        RECT 156.600 192.100 157.000 192.500 ;
        RECT 151.800 191.800 152.800 192.100 ;
        RECT 152.400 191.100 152.800 191.800 ;
        RECT 154.600 191.100 155.000 192.100 ;
        RECT 156.600 191.800 157.300 192.100 ;
        RECT 156.700 191.100 157.300 191.800 ;
        RECT 159.000 191.100 159.400 193.300 ;
        RECT 159.800 195.600 160.200 199.900 ;
        RECT 161.900 197.900 162.500 199.900 ;
        RECT 164.200 197.900 164.600 199.900 ;
        RECT 166.400 198.200 166.800 199.900 ;
        RECT 166.400 197.900 167.400 198.200 ;
        RECT 162.200 197.500 162.600 197.900 ;
        RECT 164.300 197.600 164.600 197.900 ;
        RECT 163.900 197.300 165.700 197.600 ;
        RECT 167.000 197.500 167.400 197.900 ;
        RECT 163.900 197.200 164.300 197.300 ;
        RECT 165.300 197.200 165.700 197.300 ;
        RECT 161.400 197.000 162.100 197.200 ;
        RECT 161.400 196.800 162.500 197.000 ;
        RECT 161.800 196.600 162.500 196.800 ;
        RECT 162.200 196.100 162.500 196.600 ;
        RECT 163.300 196.500 164.400 196.800 ;
        RECT 163.300 196.400 163.700 196.500 ;
        RECT 162.200 195.800 163.400 196.100 ;
        RECT 159.800 195.300 161.900 195.600 ;
        RECT 159.800 193.600 160.200 195.300 ;
        RECT 161.500 195.200 161.900 195.300 ;
        RECT 160.700 194.900 161.100 195.000 ;
        RECT 160.700 194.600 162.600 194.900 ;
        RECT 162.200 194.500 162.600 194.600 ;
        RECT 163.100 194.200 163.400 195.800 ;
        RECT 164.100 195.900 164.400 196.500 ;
        RECT 164.700 196.500 165.100 196.600 ;
        RECT 167.000 196.500 167.400 196.600 ;
        RECT 164.700 196.200 167.400 196.500 ;
        RECT 164.100 195.700 166.500 195.900 ;
        RECT 168.600 195.700 169.000 199.900 ;
        RECT 164.100 195.600 169.000 195.700 ;
        RECT 166.100 195.500 169.000 195.600 ;
        RECT 166.200 195.400 169.000 195.500 ;
        RECT 165.400 195.100 165.800 195.200 ;
        RECT 170.200 195.100 170.600 199.900 ;
        RECT 172.900 198.200 173.300 199.900 ;
        RECT 172.900 197.800 173.800 198.200 ;
        RECT 172.200 196.800 172.600 197.200 ;
        RECT 171.000 195.800 171.400 196.600 ;
        RECT 172.200 196.200 172.500 196.800 ;
        RECT 172.900 196.200 173.300 197.800 ;
        RECT 171.800 195.900 172.500 196.200 ;
        RECT 172.800 195.900 173.300 196.200 ;
        RECT 171.800 195.800 172.200 195.900 ;
        RECT 171.800 195.100 172.100 195.800 ;
        RECT 165.400 194.800 167.900 195.100 ;
        RECT 166.200 194.700 166.600 194.800 ;
        RECT 167.500 194.700 167.900 194.800 ;
        RECT 170.200 194.800 172.100 195.100 ;
        RECT 166.700 194.200 167.100 194.300 ;
        RECT 163.100 193.900 168.600 194.200 ;
        RECT 163.300 193.800 163.700 193.900 ;
        RECT 159.800 193.300 161.700 193.600 ;
        RECT 159.800 191.100 160.200 193.300 ;
        RECT 161.300 193.200 161.700 193.300 ;
        RECT 166.200 192.800 166.500 193.900 ;
        RECT 167.800 193.800 168.600 193.900 ;
        RECT 165.300 192.700 165.700 192.800 ;
        RECT 162.200 192.100 162.600 192.500 ;
        RECT 164.300 192.400 165.700 192.700 ;
        RECT 166.200 192.400 166.600 192.800 ;
        RECT 164.300 192.100 164.600 192.400 ;
        RECT 167.000 192.100 167.400 192.500 ;
        RECT 161.900 191.800 162.600 192.100 ;
        RECT 161.900 191.100 162.500 191.800 ;
        RECT 164.200 191.100 164.600 192.100 ;
        RECT 166.400 191.800 167.400 192.100 ;
        RECT 166.400 191.100 166.800 191.800 ;
        RECT 168.600 191.100 169.000 193.500 ;
        RECT 169.400 193.400 169.800 194.200 ;
        RECT 170.200 193.100 170.600 194.800 ;
        RECT 172.800 194.200 173.100 195.900 ;
        RECT 175.800 195.600 176.200 199.900 ;
        RECT 177.400 195.600 177.800 199.900 ;
        RECT 179.000 195.600 179.400 199.900 ;
        RECT 180.600 195.600 181.000 199.900 ;
        RECT 183.300 199.200 183.700 199.900 ;
        RECT 183.300 198.800 184.200 199.200 ;
        RECT 182.600 196.800 183.000 197.200 ;
        RECT 182.600 196.200 182.900 196.800 ;
        RECT 183.300 196.200 183.700 198.800 ;
        RECT 182.200 195.900 182.900 196.200 ;
        RECT 183.200 195.900 183.700 196.200 ;
        RECT 182.200 195.800 182.600 195.900 ;
        RECT 175.000 195.200 176.200 195.600 ;
        RECT 176.700 195.200 177.800 195.600 ;
        RECT 178.300 195.200 179.400 195.600 ;
        RECT 180.100 195.200 181.000 195.600 ;
        RECT 173.400 194.400 173.800 195.200 ;
        RECT 171.800 193.800 173.100 194.200 ;
        RECT 174.200 194.100 174.600 194.200 ;
        RECT 173.800 193.800 174.600 194.100 ;
        RECT 175.000 193.800 175.400 195.200 ;
        RECT 176.700 194.500 177.100 195.200 ;
        RECT 178.300 194.500 178.700 195.200 ;
        RECT 180.100 194.500 180.500 195.200 ;
        RECT 175.800 194.100 177.100 194.500 ;
        RECT 177.500 194.100 178.700 194.500 ;
        RECT 179.200 194.100 180.500 194.500 ;
        RECT 183.200 194.200 183.500 195.900 ;
        RECT 185.400 195.800 185.800 196.600 ;
        RECT 183.800 195.100 184.200 195.200 ;
        RECT 186.200 195.100 186.600 199.900 ;
        RECT 187.800 199.600 189.800 199.900 ;
        RECT 187.800 195.900 188.200 199.600 ;
        RECT 188.600 195.800 189.000 199.300 ;
        RECT 189.400 196.200 189.800 199.600 ;
        RECT 191.000 196.200 191.400 199.900 ;
        RECT 189.400 195.900 191.400 196.200 ;
        RECT 191.800 197.500 192.200 199.500 ;
        RECT 188.700 195.600 189.000 195.800 ;
        RECT 191.800 195.800 192.100 197.500 ;
        RECT 193.900 196.400 194.300 199.900 ;
        RECT 198.500 196.400 198.900 199.900 ;
        RECT 200.600 197.500 201.000 199.500 ;
        RECT 193.900 196.100 194.700 196.400 ;
        RECT 183.800 194.800 186.600 195.100 ;
        RECT 187.800 194.800 188.200 195.600 ;
        RECT 188.700 195.300 189.700 195.600 ;
        RECT 191.800 195.500 193.700 195.800 ;
        RECT 189.400 195.200 189.700 195.300 ;
        RECT 190.600 195.200 191.000 195.400 ;
        RECT 189.400 194.800 189.800 195.200 ;
        RECT 190.600 194.900 191.400 195.200 ;
        RECT 191.000 194.800 191.400 194.900 ;
        RECT 183.800 194.400 184.200 194.800 ;
        RECT 176.700 193.800 177.100 194.100 ;
        RECT 178.300 193.800 178.700 194.100 ;
        RECT 180.100 193.800 180.500 194.100 ;
        RECT 182.200 193.800 183.500 194.200 ;
        RECT 184.600 194.100 185.000 194.200 ;
        RECT 184.200 193.800 185.000 194.100 ;
        RECT 171.900 193.100 172.200 193.800 ;
        RECT 173.800 193.600 174.200 193.800 ;
        RECT 175.000 193.400 176.200 193.800 ;
        RECT 176.700 193.400 177.800 193.800 ;
        RECT 178.300 193.400 179.400 193.800 ;
        RECT 180.100 193.400 181.000 193.800 ;
        RECT 172.700 193.100 174.500 193.300 ;
        RECT 170.200 192.800 171.100 193.100 ;
        RECT 170.700 191.100 171.100 192.800 ;
        RECT 171.800 191.100 172.200 193.100 ;
        RECT 172.600 193.000 174.600 193.100 ;
        RECT 172.600 191.100 173.000 193.000 ;
        RECT 174.200 191.100 174.600 193.000 ;
        RECT 175.800 191.100 176.200 193.400 ;
        RECT 177.400 191.100 177.800 193.400 ;
        RECT 179.000 191.100 179.400 193.400 ;
        RECT 180.600 191.100 181.000 193.400 ;
        RECT 182.300 193.100 182.600 193.800 ;
        RECT 184.200 193.600 184.600 193.800 ;
        RECT 183.100 193.100 184.900 193.300 ;
        RECT 186.200 193.100 186.600 194.800 ;
        RECT 188.700 194.400 189.100 194.800 ;
        RECT 188.700 194.200 189.000 194.400 ;
        RECT 187.000 193.400 187.400 194.200 ;
        RECT 188.600 193.800 189.000 194.200 ;
        RECT 189.400 193.100 189.700 194.800 ;
        RECT 190.200 193.800 190.600 194.600 ;
        RECT 191.800 194.400 192.200 195.200 ;
        RECT 192.600 194.400 193.000 195.200 ;
        RECT 193.400 194.500 193.700 195.500 ;
        RECT 193.400 194.100 194.100 194.500 ;
        RECT 194.400 194.200 194.700 196.100 ;
        RECT 198.100 196.100 198.900 196.400 ;
        RECT 195.000 194.800 195.400 195.600 ;
        RECT 197.400 194.800 197.800 195.600 ;
        RECT 198.100 194.200 198.400 196.100 ;
        RECT 200.700 195.800 201.000 197.500 ;
        RECT 199.100 195.500 201.000 195.800 ;
        RECT 203.000 195.600 203.400 199.900 ;
        RECT 205.100 197.900 205.700 199.900 ;
        RECT 207.400 197.900 207.800 199.900 ;
        RECT 209.600 198.200 210.000 199.900 ;
        RECT 209.600 197.900 210.600 198.200 ;
        RECT 205.400 197.500 205.800 197.900 ;
        RECT 207.500 197.600 207.800 197.900 ;
        RECT 207.100 197.300 208.900 197.600 ;
        RECT 210.200 197.500 210.600 197.900 ;
        RECT 207.100 197.200 207.500 197.300 ;
        RECT 208.500 197.200 208.900 197.300 ;
        RECT 205.000 196.600 205.700 197.000 ;
        RECT 205.400 196.100 205.700 196.600 ;
        RECT 206.500 196.500 207.600 196.800 ;
        RECT 206.500 196.400 206.900 196.500 ;
        RECT 205.400 195.800 206.600 196.100 ;
        RECT 199.100 194.500 199.400 195.500 ;
        RECT 203.000 195.300 205.100 195.600 ;
        RECT 193.400 193.900 193.900 194.100 ;
        RECT 191.800 193.600 193.900 193.900 ;
        RECT 194.400 193.800 195.400 194.200 ;
        RECT 195.800 194.100 196.200 194.200 ;
        RECT 197.400 194.100 198.400 194.200 ;
        RECT 198.700 194.100 199.400 194.500 ;
        RECT 199.800 194.400 200.200 195.200 ;
        RECT 200.600 194.400 201.000 195.200 ;
        RECT 195.800 193.800 198.400 194.100 ;
        RECT 182.200 191.100 182.600 193.100 ;
        RECT 183.000 193.000 185.000 193.100 ;
        RECT 183.000 191.100 183.400 193.000 ;
        RECT 184.600 191.100 185.000 193.000 ;
        RECT 185.700 192.800 186.600 193.100 ;
        RECT 185.700 191.100 186.100 192.800 ;
        RECT 189.100 191.100 189.900 193.100 ;
        RECT 191.800 192.500 192.100 193.600 ;
        RECT 194.400 193.500 194.700 193.800 ;
        RECT 194.300 193.300 194.700 193.500 ;
        RECT 193.900 193.000 194.700 193.300 ;
        RECT 198.100 193.500 198.400 193.800 ;
        RECT 198.900 193.900 199.400 194.100 ;
        RECT 198.900 193.600 201.000 193.900 ;
        RECT 198.100 193.300 198.500 193.500 ;
        RECT 198.100 193.000 198.900 193.300 ;
        RECT 191.800 191.500 192.200 192.500 ;
        RECT 193.900 192.200 194.300 193.000 ;
        RECT 193.400 191.800 194.300 192.200 ;
        RECT 193.900 191.500 194.300 191.800 ;
        RECT 198.500 191.500 198.900 193.000 ;
        RECT 200.700 192.500 201.000 193.600 ;
        RECT 200.600 191.500 201.000 192.500 ;
        RECT 203.000 193.600 203.400 195.300 ;
        RECT 204.700 195.200 205.100 195.300 ;
        RECT 203.900 194.900 204.300 195.000 ;
        RECT 203.900 194.600 205.800 194.900 ;
        RECT 205.400 194.500 205.800 194.600 ;
        RECT 206.300 194.200 206.600 195.800 ;
        RECT 207.300 195.900 207.600 196.500 ;
        RECT 207.900 196.500 208.300 196.600 ;
        RECT 210.200 196.500 210.600 196.600 ;
        RECT 207.900 196.200 210.600 196.500 ;
        RECT 207.300 195.700 209.700 195.900 ;
        RECT 211.800 195.700 212.200 199.900 ;
        RECT 213.900 196.200 214.300 199.900 ;
        RECT 214.600 196.800 215.000 197.200 ;
        RECT 214.700 196.200 215.000 196.800 ;
        RECT 217.100 196.200 217.500 199.900 ;
        RECT 217.800 196.800 218.200 197.200 ;
        RECT 217.900 196.200 218.200 196.800 ;
        RECT 213.400 195.800 214.400 196.200 ;
        RECT 214.700 195.900 215.400 196.200 ;
        RECT 217.100 195.900 217.600 196.200 ;
        RECT 217.900 195.900 218.600 196.200 ;
        RECT 215.000 195.800 215.400 195.900 ;
        RECT 207.300 195.600 212.200 195.700 ;
        RECT 209.300 195.500 212.200 195.600 ;
        RECT 209.400 195.400 212.200 195.500 ;
        RECT 208.600 195.100 209.000 195.200 ;
        RECT 208.600 194.800 211.100 195.100 ;
        RECT 210.700 194.700 211.100 194.800 ;
        RECT 213.400 194.400 213.800 195.200 ;
        RECT 209.900 194.200 210.300 194.300 ;
        RECT 214.100 194.200 214.400 195.800 ;
        RECT 216.600 194.400 217.000 195.200 ;
        RECT 217.300 194.200 217.600 195.900 ;
        RECT 218.200 195.800 218.600 195.900 ;
        RECT 219.000 195.800 219.400 196.600 ;
        RECT 218.200 195.100 218.500 195.800 ;
        RECT 219.800 195.100 220.200 199.900 ;
        RECT 220.600 197.100 221.000 197.200 ;
        RECT 221.400 197.100 221.800 199.900 ;
        RECT 223.500 197.900 224.100 199.900 ;
        RECT 225.800 197.900 226.200 199.900 ;
        RECT 228.000 198.200 228.400 199.900 ;
        RECT 228.000 197.900 229.000 198.200 ;
        RECT 223.800 197.500 224.200 197.900 ;
        RECT 225.900 197.600 226.200 197.900 ;
        RECT 225.500 197.300 227.300 197.600 ;
        RECT 228.600 197.500 229.000 197.900 ;
        RECT 225.500 197.200 225.900 197.300 ;
        RECT 226.900 197.200 227.300 197.300 ;
        RECT 220.600 196.800 221.800 197.100 ;
        RECT 218.200 194.800 220.200 195.100 ;
        RECT 206.300 193.900 211.800 194.200 ;
        RECT 206.500 193.800 206.900 193.900 ;
        RECT 209.400 193.800 209.800 193.900 ;
        RECT 211.000 193.800 211.800 193.900 ;
        RECT 212.600 194.100 213.000 194.200 ;
        RECT 212.600 193.800 213.400 194.100 ;
        RECT 214.100 193.800 215.400 194.200 ;
        RECT 215.800 194.100 216.200 194.200 ;
        RECT 217.300 194.100 218.600 194.200 ;
        RECT 219.000 194.100 219.400 194.200 ;
        RECT 215.800 193.800 216.600 194.100 ;
        RECT 217.300 193.800 219.400 194.100 ;
        RECT 203.000 193.300 204.900 193.600 ;
        RECT 203.000 191.100 203.400 193.300 ;
        RECT 204.500 193.200 204.900 193.300 ;
        RECT 209.400 192.800 209.700 193.800 ;
        RECT 213.000 193.600 213.400 193.800 ;
        RECT 208.500 192.700 208.900 192.800 ;
        RECT 205.400 192.100 205.800 192.500 ;
        RECT 207.500 192.400 208.900 192.700 ;
        RECT 209.400 192.400 209.800 192.800 ;
        RECT 207.500 192.100 207.800 192.400 ;
        RECT 210.200 192.100 210.600 192.500 ;
        RECT 205.100 191.800 205.800 192.100 ;
        RECT 205.100 191.100 205.700 191.800 ;
        RECT 207.400 191.100 207.800 192.100 ;
        RECT 209.600 191.800 210.600 192.100 ;
        RECT 209.600 191.100 210.000 191.800 ;
        RECT 211.800 191.100 212.200 193.500 ;
        RECT 212.700 193.100 214.500 193.300 ;
        RECT 215.000 193.100 215.300 193.800 ;
        RECT 216.200 193.600 216.600 193.800 ;
        RECT 215.900 193.100 217.700 193.300 ;
        RECT 218.200 193.100 218.500 193.800 ;
        RECT 219.800 193.100 220.200 194.800 ;
        RECT 221.400 195.600 221.800 196.800 ;
        RECT 223.400 196.600 224.100 197.000 ;
        RECT 223.800 196.100 224.100 196.600 ;
        RECT 224.900 196.500 226.000 196.800 ;
        RECT 224.900 196.400 225.300 196.500 ;
        RECT 223.800 195.800 225.000 196.100 ;
        RECT 221.400 195.300 223.500 195.600 ;
        RECT 220.600 193.400 221.000 194.200 ;
        RECT 221.400 193.600 221.800 195.300 ;
        RECT 223.100 195.200 223.500 195.300 ;
        RECT 224.700 195.200 225.000 195.800 ;
        RECT 225.700 195.900 226.000 196.500 ;
        RECT 226.300 196.500 226.700 196.600 ;
        RECT 228.600 196.500 229.000 196.600 ;
        RECT 226.300 196.200 229.000 196.500 ;
        RECT 225.700 195.700 228.100 195.900 ;
        RECT 230.200 195.700 230.600 199.900 ;
        RECT 232.300 196.200 232.700 199.900 ;
        RECT 233.000 196.800 233.400 197.200 ;
        RECT 233.100 196.200 233.400 196.800 ;
        RECT 232.300 195.900 232.800 196.200 ;
        RECT 233.100 195.900 233.800 196.200 ;
        RECT 225.700 195.600 230.600 195.700 ;
        RECT 227.700 195.500 230.600 195.600 ;
        RECT 227.800 195.400 230.600 195.500 ;
        RECT 222.300 194.900 222.700 195.000 ;
        RECT 222.300 194.600 224.200 194.900 ;
        RECT 224.600 194.800 225.000 195.200 ;
        RECT 227.000 195.100 227.400 195.200 ;
        RECT 227.000 194.800 229.500 195.100 ;
        RECT 223.800 194.500 224.200 194.600 ;
        RECT 224.700 194.200 225.000 194.800 ;
        RECT 229.100 194.700 229.500 194.800 ;
        RECT 231.800 194.400 232.200 195.200 ;
        RECT 228.300 194.200 228.700 194.300 ;
        RECT 232.500 194.200 232.800 195.900 ;
        RECT 233.400 195.800 233.800 195.900 ;
        RECT 234.200 195.600 234.600 199.900 ;
        RECT 236.300 197.900 236.900 199.900 ;
        RECT 238.600 197.900 239.000 199.900 ;
        RECT 240.800 198.200 241.200 199.900 ;
        RECT 240.800 197.900 241.800 198.200 ;
        RECT 236.600 197.500 237.000 197.900 ;
        RECT 238.700 197.600 239.000 197.900 ;
        RECT 238.300 197.300 240.100 197.600 ;
        RECT 241.400 197.500 241.800 197.900 ;
        RECT 238.300 197.200 238.700 197.300 ;
        RECT 239.700 197.200 240.100 197.300 ;
        RECT 236.200 196.600 236.900 197.000 ;
        RECT 236.600 196.100 236.900 196.600 ;
        RECT 237.700 196.500 238.800 196.800 ;
        RECT 237.700 196.400 238.100 196.500 ;
        RECT 236.600 195.800 237.800 196.100 ;
        RECT 234.200 195.300 236.300 195.600 ;
        RECT 224.700 193.900 230.200 194.200 ;
        RECT 224.900 193.800 225.300 193.900 ;
        RECT 212.600 193.000 214.600 193.100 ;
        RECT 212.600 191.100 213.000 193.000 ;
        RECT 214.200 191.100 214.600 193.000 ;
        RECT 215.000 191.100 215.400 193.100 ;
        RECT 215.800 193.000 217.800 193.100 ;
        RECT 215.800 191.100 216.200 193.000 ;
        RECT 217.400 191.100 217.800 193.000 ;
        RECT 218.200 191.100 218.600 193.100 ;
        RECT 219.300 192.800 220.200 193.100 ;
        RECT 221.400 193.300 223.300 193.600 ;
        RECT 219.300 191.100 219.700 192.800 ;
        RECT 221.400 191.100 221.800 193.300 ;
        RECT 222.900 193.200 223.300 193.300 ;
        RECT 227.800 192.800 228.100 193.900 ;
        RECT 229.400 193.800 230.200 193.900 ;
        RECT 231.000 194.100 231.400 194.200 ;
        RECT 231.000 193.800 231.800 194.100 ;
        RECT 232.500 193.800 233.800 194.200 ;
        RECT 231.400 193.600 231.800 193.800 ;
        RECT 226.900 192.700 227.300 192.800 ;
        RECT 223.800 192.100 224.200 192.500 ;
        RECT 225.900 192.400 227.300 192.700 ;
        RECT 227.800 192.400 228.200 192.800 ;
        RECT 225.900 192.100 226.200 192.400 ;
        RECT 228.600 192.100 229.000 192.500 ;
        RECT 223.500 191.800 224.200 192.100 ;
        RECT 223.500 191.100 224.100 191.800 ;
        RECT 225.800 191.100 226.200 192.100 ;
        RECT 228.000 191.800 229.000 192.100 ;
        RECT 228.000 191.100 228.400 191.800 ;
        RECT 230.200 191.100 230.600 193.500 ;
        RECT 231.100 193.100 232.900 193.300 ;
        RECT 233.400 193.100 233.700 193.800 ;
        RECT 234.200 193.600 234.600 195.300 ;
        RECT 235.900 195.200 236.300 195.300 ;
        RECT 235.100 194.900 235.500 195.000 ;
        RECT 235.100 194.600 237.000 194.900 ;
        RECT 236.600 194.500 237.000 194.600 ;
        RECT 237.500 194.200 237.800 195.800 ;
        RECT 238.500 195.900 238.800 196.500 ;
        RECT 239.100 196.500 239.500 196.600 ;
        RECT 241.400 196.500 241.800 196.600 ;
        RECT 239.100 196.200 241.800 196.500 ;
        RECT 238.500 195.700 240.900 195.900 ;
        RECT 243.000 195.700 243.400 199.900 ;
        RECT 244.200 196.800 244.600 197.200 ;
        RECT 244.200 196.200 244.500 196.800 ;
        RECT 244.900 196.200 245.300 199.900 ;
        RECT 243.800 195.900 244.500 196.200 ;
        RECT 244.800 195.900 245.300 196.200 ;
        RECT 247.000 196.200 247.400 199.900 ;
        RECT 248.600 196.400 249.000 199.900 ;
        RECT 247.000 195.900 248.300 196.200 ;
        RECT 248.600 195.900 249.100 196.400 ;
        RECT 243.800 195.800 244.200 195.900 ;
        RECT 238.500 195.600 243.400 195.700 ;
        RECT 240.500 195.500 243.400 195.600 ;
        RECT 240.600 195.400 243.400 195.500 ;
        RECT 239.000 195.100 239.400 195.200 ;
        RECT 239.800 195.100 240.200 195.200 ;
        RECT 239.000 194.800 242.300 195.100 ;
        RECT 241.900 194.700 242.300 194.800 ;
        RECT 241.100 194.200 241.500 194.300 ;
        RECT 244.800 194.200 245.100 195.900 ;
        RECT 245.400 194.400 245.800 195.200 ;
        RECT 247.000 194.800 247.500 195.200 ;
        RECT 247.100 194.400 247.500 194.800 ;
        RECT 248.000 194.900 248.300 195.900 ;
        RECT 248.000 194.500 248.500 194.900 ;
        RECT 237.500 193.900 243.000 194.200 ;
        RECT 237.700 193.800 238.100 193.900 ;
        RECT 234.200 193.300 236.100 193.600 ;
        RECT 231.000 193.000 233.000 193.100 ;
        RECT 231.000 191.100 231.400 193.000 ;
        RECT 232.600 191.100 233.000 193.000 ;
        RECT 233.400 191.100 233.800 193.100 ;
        RECT 234.200 191.100 234.600 193.300 ;
        RECT 235.700 193.200 236.100 193.300 ;
        RECT 240.600 193.200 240.900 193.900 ;
        RECT 242.200 193.800 243.000 193.900 ;
        RECT 243.800 193.800 245.100 194.200 ;
        RECT 246.200 194.100 246.600 194.200 ;
        RECT 245.800 193.800 246.600 194.100 ;
        RECT 239.700 192.700 240.100 192.800 ;
        RECT 236.600 192.100 237.000 192.500 ;
        RECT 238.700 192.400 240.100 192.700 ;
        RECT 240.600 192.400 241.000 193.200 ;
        RECT 238.700 192.100 239.000 192.400 ;
        RECT 241.400 192.100 241.800 192.500 ;
        RECT 236.300 191.800 237.000 192.100 ;
        RECT 236.300 191.100 236.900 191.800 ;
        RECT 238.600 191.100 239.000 192.100 ;
        RECT 240.800 191.800 241.800 192.100 ;
        RECT 240.800 191.100 241.200 191.800 ;
        RECT 243.000 191.100 243.400 193.500 ;
        RECT 243.900 193.100 244.200 193.800 ;
        RECT 245.800 193.600 246.200 193.800 ;
        RECT 248.000 193.700 248.300 194.500 ;
        RECT 248.800 194.200 249.100 195.900 ;
        RECT 248.600 193.800 249.100 194.200 ;
        RECT 247.000 193.400 248.300 193.700 ;
        RECT 244.700 193.100 246.500 193.300 ;
        RECT 243.800 191.100 244.200 193.100 ;
        RECT 244.600 193.000 246.600 193.100 ;
        RECT 244.600 191.100 245.000 193.000 ;
        RECT 246.200 191.100 246.600 193.000 ;
        RECT 247.000 191.100 247.400 193.400 ;
        RECT 248.800 193.100 249.100 193.800 ;
        RECT 248.600 192.800 249.100 193.100 ;
        RECT 248.600 191.100 249.000 192.800 ;
        RECT 1.900 188.200 2.300 189.900 ;
        RECT 1.400 187.900 2.300 188.200 ;
        RECT 3.000 187.900 3.400 189.900 ;
        RECT 3.800 188.000 4.200 189.900 ;
        RECT 5.400 188.000 5.800 189.900 ;
        RECT 3.800 187.900 5.800 188.000 ;
        RECT 6.200 188.000 6.600 189.900 ;
        RECT 7.800 188.000 8.200 189.900 ;
        RECT 6.200 187.900 8.200 188.000 ;
        RECT 8.600 187.900 9.000 189.900 ;
        RECT 9.700 188.200 10.100 189.900 ;
        RECT 9.700 187.900 10.600 188.200 ;
        RECT 13.700 188.000 14.100 189.500 ;
        RECT 15.800 188.500 16.200 189.500 ;
        RECT 0.600 186.800 1.000 187.600 ;
        RECT 1.400 186.100 1.800 187.900 ;
        RECT 3.100 187.200 3.400 187.900 ;
        RECT 3.900 187.700 5.700 187.900 ;
        RECT 6.300 187.700 8.100 187.900 ;
        RECT 5.000 187.200 5.400 187.400 ;
        RECT 6.600 187.200 7.000 187.400 ;
        RECT 8.600 187.200 8.900 187.900 ;
        RECT 3.000 186.800 4.300 187.200 ;
        RECT 5.000 187.100 5.800 187.200 ;
        RECT 6.200 187.100 7.000 187.200 ;
        RECT 5.000 186.900 7.000 187.100 ;
        RECT 5.400 186.800 6.600 186.900 ;
        RECT 7.700 186.800 9.000 187.200 ;
        RECT 1.400 185.800 3.300 186.100 ;
        RECT 1.400 181.100 1.800 185.800 ;
        RECT 3.000 185.200 3.300 185.800 ;
        RECT 2.200 184.400 2.600 185.200 ;
        RECT 3.000 185.100 3.400 185.200 ;
        RECT 4.000 185.100 4.300 186.800 ;
        RECT 4.600 185.800 5.000 186.600 ;
        RECT 7.000 185.800 7.400 186.600 ;
        RECT 7.700 185.100 8.000 186.800 ;
        RECT 10.200 186.100 10.600 187.900 ;
        RECT 13.300 187.700 14.100 188.000 ;
        RECT 11.000 187.100 11.400 187.600 ;
        RECT 13.300 187.500 13.700 187.700 ;
        RECT 13.300 187.200 13.600 187.500 ;
        RECT 15.900 187.400 16.200 188.500 ;
        RECT 17.400 187.600 17.800 189.900 ;
        RECT 19.000 187.600 19.400 189.900 ;
        RECT 20.600 187.600 21.000 189.900 ;
        RECT 22.200 187.600 22.600 189.900 ;
        RECT 25.700 188.000 26.100 189.500 ;
        RECT 27.800 188.500 28.200 189.500 ;
        RECT 11.800 187.100 12.200 187.200 ;
        RECT 11.000 186.800 12.200 187.100 ;
        RECT 12.600 186.800 13.600 187.200 ;
        RECT 14.100 187.100 16.200 187.400 ;
        RECT 16.600 187.200 17.800 187.600 ;
        RECT 18.300 187.200 19.400 187.600 ;
        RECT 19.900 187.200 21.000 187.600 ;
        RECT 21.700 187.200 22.600 187.600 ;
        RECT 25.300 187.700 26.100 188.000 ;
        RECT 25.300 187.500 25.700 187.700 ;
        RECT 25.300 187.200 25.600 187.500 ;
        RECT 27.900 187.400 28.200 188.500 ;
        RECT 30.500 188.000 30.900 189.500 ;
        RECT 32.600 188.500 33.000 189.500 ;
        RECT 14.100 186.900 14.600 187.100 ;
        RECT 8.600 185.800 10.600 186.100 ;
        RECT 11.000 186.100 11.400 186.200 ;
        RECT 12.600 186.100 13.000 186.200 ;
        RECT 11.000 185.800 13.000 186.100 ;
        RECT 8.600 185.200 8.900 185.800 ;
        RECT 8.600 185.100 9.000 185.200 ;
        RECT 3.000 184.800 3.700 185.100 ;
        RECT 4.000 184.800 4.500 185.100 ;
        RECT 3.400 184.200 3.700 184.800 ;
        RECT 3.400 183.800 3.800 184.200 ;
        RECT 4.100 181.100 4.500 184.800 ;
        RECT 7.500 184.800 8.000 185.100 ;
        RECT 8.300 184.800 9.000 185.100 ;
        RECT 7.500 181.100 7.900 184.800 ;
        RECT 8.300 184.200 8.600 184.800 ;
        RECT 9.400 184.400 9.800 185.200 ;
        RECT 8.200 183.800 8.600 184.200 ;
        RECT 10.200 181.100 10.600 185.800 ;
        RECT 12.600 185.400 13.000 185.800 ;
        RECT 13.300 185.200 13.600 186.800 ;
        RECT 13.900 186.500 14.600 186.900 ;
        RECT 14.300 185.500 14.600 186.500 ;
        RECT 15.000 185.800 15.400 186.600 ;
        RECT 15.800 185.800 16.200 186.600 ;
        RECT 16.600 185.800 17.000 187.200 ;
        RECT 18.300 186.900 18.700 187.200 ;
        RECT 19.900 186.900 20.300 187.200 ;
        RECT 21.700 186.900 22.100 187.200 ;
        RECT 23.000 186.900 23.400 187.200 ;
        RECT 17.400 186.500 18.700 186.900 ;
        RECT 19.100 186.500 20.300 186.900 ;
        RECT 20.800 186.500 22.100 186.900 ;
        RECT 22.500 186.500 23.400 186.900 ;
        RECT 24.600 186.800 25.600 187.200 ;
        RECT 26.100 187.100 28.200 187.400 ;
        RECT 30.100 187.700 30.900 188.000 ;
        RECT 30.100 187.500 30.500 187.700 ;
        RECT 30.100 187.200 30.400 187.500 ;
        RECT 32.700 187.400 33.000 188.500 ;
        RECT 34.200 187.600 34.600 189.900 ;
        RECT 35.800 187.600 36.200 189.900 ;
        RECT 37.400 187.600 37.800 189.900 ;
        RECT 39.000 187.600 39.400 189.900 ;
        RECT 41.400 188.900 41.800 189.900 ;
        RECT 40.600 187.800 41.000 188.600 ;
        RECT 41.500 188.100 41.800 188.900 ;
        RECT 43.100 188.200 43.500 188.600 ;
        RECT 43.000 188.100 43.400 188.200 ;
        RECT 41.400 187.800 43.400 188.100 ;
        RECT 43.800 187.900 44.200 189.900 ;
        RECT 26.100 186.900 26.600 187.100 ;
        RECT 18.300 185.800 18.700 186.500 ;
        RECT 19.900 185.800 20.300 186.500 ;
        RECT 21.700 185.800 22.100 186.500 ;
        RECT 14.300 185.200 16.200 185.500 ;
        RECT 16.600 185.400 17.800 185.800 ;
        RECT 18.300 185.400 19.400 185.800 ;
        RECT 19.900 185.400 21.000 185.800 ;
        RECT 21.700 185.400 22.600 185.800 ;
        RECT 24.600 185.400 25.000 186.200 ;
        RECT 13.300 184.900 13.800 185.200 ;
        RECT 13.300 184.600 14.100 184.900 ;
        RECT 13.700 181.100 14.100 184.600 ;
        RECT 15.900 183.500 16.200 185.200 ;
        RECT 15.800 181.500 16.200 183.500 ;
        RECT 17.400 181.100 17.800 185.400 ;
        RECT 19.000 181.100 19.400 185.400 ;
        RECT 20.600 181.100 21.000 185.400 ;
        RECT 22.200 181.100 22.600 185.400 ;
        RECT 25.300 184.900 25.600 186.800 ;
        RECT 25.900 186.500 26.600 186.900 ;
        RECT 29.400 186.800 30.400 187.200 ;
        RECT 30.900 187.100 33.000 187.400 ;
        RECT 33.400 187.200 34.600 187.600 ;
        RECT 35.100 187.200 36.200 187.600 ;
        RECT 36.700 187.200 37.800 187.600 ;
        RECT 38.500 187.200 39.400 187.600 ;
        RECT 41.500 187.200 41.800 187.800 ;
        RECT 30.900 186.900 31.400 187.100 ;
        RECT 26.300 185.500 26.600 186.500 ;
        RECT 27.000 185.800 27.400 186.600 ;
        RECT 27.800 185.800 28.200 186.600 ;
        RECT 26.300 185.200 28.200 185.500 ;
        RECT 29.400 185.400 29.800 186.200 ;
        RECT 25.300 184.600 26.100 184.900 ;
        RECT 25.700 182.200 26.100 184.600 ;
        RECT 27.900 183.500 28.200 185.200 ;
        RECT 30.100 184.900 30.400 186.800 ;
        RECT 30.700 186.500 31.400 186.900 ;
        RECT 31.100 185.500 31.400 186.500 ;
        RECT 31.800 185.800 32.200 186.600 ;
        RECT 32.600 185.800 33.000 186.600 ;
        RECT 33.400 185.800 33.800 187.200 ;
        RECT 35.100 186.900 35.500 187.200 ;
        RECT 36.700 186.900 37.100 187.200 ;
        RECT 38.500 186.900 38.900 187.200 ;
        RECT 39.800 186.900 40.200 187.200 ;
        RECT 34.200 186.500 35.500 186.900 ;
        RECT 35.900 186.500 37.100 186.900 ;
        RECT 37.600 186.500 38.900 186.900 ;
        RECT 39.300 186.500 40.200 186.900 ;
        RECT 41.400 186.800 41.800 187.200 ;
        RECT 35.100 185.800 35.500 186.500 ;
        RECT 36.700 185.800 37.100 186.500 ;
        RECT 38.500 185.800 38.900 186.500 ;
        RECT 31.100 185.200 33.000 185.500 ;
        RECT 33.400 185.400 34.600 185.800 ;
        RECT 35.100 185.400 36.200 185.800 ;
        RECT 36.700 185.400 37.800 185.800 ;
        RECT 38.500 185.400 39.400 185.800 ;
        RECT 30.100 184.600 30.900 184.900 ;
        RECT 25.400 181.800 26.100 182.200 ;
        RECT 25.700 181.100 26.100 181.800 ;
        RECT 27.800 181.500 28.200 183.500 ;
        RECT 30.500 182.200 30.900 184.600 ;
        RECT 32.700 183.500 33.000 185.200 ;
        RECT 30.200 181.800 30.900 182.200 ;
        RECT 30.500 181.100 30.900 181.800 ;
        RECT 32.600 181.500 33.000 183.500 ;
        RECT 34.200 181.100 34.600 185.400 ;
        RECT 35.800 181.100 36.200 185.400 ;
        RECT 37.400 181.100 37.800 185.400 ;
        RECT 39.000 181.100 39.400 185.400 ;
        RECT 41.500 185.100 41.800 186.800 ;
        RECT 43.900 186.200 44.200 187.900 ;
        RECT 47.800 187.700 48.200 189.900 ;
        RECT 49.900 189.200 50.500 189.900 ;
        RECT 49.900 188.900 50.600 189.200 ;
        RECT 52.200 188.900 52.600 189.900 ;
        RECT 54.400 189.200 54.800 189.900 ;
        RECT 54.400 188.900 55.400 189.200 ;
        RECT 50.200 188.500 50.600 188.900 ;
        RECT 52.300 188.600 52.600 188.900 ;
        RECT 52.300 188.300 53.700 188.600 ;
        RECT 53.300 188.200 53.700 188.300 ;
        RECT 54.200 188.200 54.600 188.600 ;
        RECT 55.000 188.500 55.400 188.900 ;
        RECT 49.300 187.700 49.700 187.800 ;
        RECT 47.800 187.400 49.700 187.700 ;
        RECT 44.600 186.400 45.000 187.200 ;
        RECT 42.200 185.400 42.600 186.200 ;
        RECT 43.000 186.100 43.400 186.200 ;
        RECT 43.800 186.100 44.200 186.200 ;
        RECT 45.400 186.100 45.800 186.200 ;
        RECT 43.000 185.800 44.200 186.100 ;
        RECT 45.000 185.800 45.800 186.100 ;
        RECT 43.100 185.100 43.400 185.800 ;
        RECT 45.000 185.600 45.400 185.800 ;
        RECT 47.800 185.700 48.200 187.400 ;
        RECT 51.300 187.100 51.700 187.200 ;
        RECT 54.200 187.100 54.500 188.200 ;
        RECT 56.600 187.500 57.000 189.900 ;
        RECT 57.400 188.500 57.800 189.500 ;
        RECT 57.400 187.400 57.700 188.500 ;
        RECT 59.500 188.000 59.900 189.500 ;
        RECT 64.100 188.000 64.500 189.500 ;
        RECT 66.200 188.500 66.600 189.500 ;
        RECT 59.500 187.700 60.300 188.000 ;
        RECT 59.900 187.500 60.300 187.700 ;
        RECT 55.800 187.100 56.600 187.200 ;
        RECT 57.400 187.100 59.500 187.400 ;
        RECT 51.100 186.800 56.600 187.100 ;
        RECT 59.000 186.900 59.500 187.100 ;
        RECT 60.000 187.200 60.300 187.500 ;
        RECT 63.700 187.700 64.500 188.000 ;
        RECT 63.700 187.500 64.100 187.700 ;
        RECT 63.700 187.200 64.000 187.500 ;
        RECT 66.300 187.400 66.600 188.500 ;
        RECT 50.200 186.400 50.600 186.500 ;
        RECT 48.700 186.100 50.600 186.400 ;
        RECT 51.100 186.200 51.400 186.800 ;
        RECT 54.700 186.700 55.100 186.800 ;
        RECT 55.500 186.200 55.900 186.300 ;
        RECT 48.700 186.000 49.100 186.100 ;
        RECT 51.000 185.800 51.400 186.200 ;
        RECT 53.400 185.900 55.900 186.200 ;
        RECT 53.400 185.800 53.800 185.900 ;
        RECT 57.400 185.800 57.800 186.600 ;
        RECT 58.200 185.800 58.600 186.600 ;
        RECT 59.000 186.500 59.700 186.900 ;
        RECT 60.000 186.800 61.000 187.200 ;
        RECT 63.000 186.800 64.000 187.200 ;
        RECT 64.500 187.100 66.600 187.400 ;
        RECT 67.000 188.500 67.400 189.500 ;
        RECT 67.000 187.400 67.300 188.500 ;
        RECT 69.100 188.000 69.500 189.500 ;
        RECT 73.100 189.200 73.900 189.900 ;
        RECT 72.600 188.800 73.900 189.200 ;
        RECT 69.100 187.700 69.900 188.000 ;
        RECT 73.100 187.900 73.900 188.800 ;
        RECT 69.500 187.500 69.900 187.700 ;
        RECT 67.000 187.100 69.100 187.400 ;
        RECT 64.500 186.900 65.000 187.100 ;
        RECT 49.500 185.700 49.900 185.800 ;
        RECT 47.800 185.400 49.900 185.700 ;
        RECT 41.400 184.700 42.300 185.100 ;
        RECT 41.900 181.100 42.300 184.700 ;
        RECT 43.000 181.100 43.400 185.100 ;
        RECT 43.800 184.800 45.800 185.100 ;
        RECT 43.800 181.100 44.200 184.800 ;
        RECT 45.400 181.100 45.800 184.800 ;
        RECT 47.800 181.100 48.200 185.400 ;
        RECT 51.100 185.200 51.400 185.800 ;
        RECT 54.200 185.500 57.000 185.600 ;
        RECT 59.000 185.500 59.300 186.500 ;
        RECT 54.100 185.400 57.000 185.500 ;
        RECT 50.200 184.900 51.400 185.200 ;
        RECT 52.100 185.300 57.000 185.400 ;
        RECT 52.100 185.100 54.500 185.300 ;
        RECT 50.200 184.400 50.500 184.900 ;
        RECT 49.800 184.000 50.500 184.400 ;
        RECT 51.300 184.500 51.700 184.600 ;
        RECT 52.100 184.500 52.400 185.100 ;
        RECT 51.300 184.200 52.400 184.500 ;
        RECT 52.700 184.500 55.400 184.800 ;
        RECT 52.700 184.400 53.100 184.500 ;
        RECT 55.000 184.400 55.400 184.500 ;
        RECT 51.900 183.700 52.300 183.800 ;
        RECT 53.300 183.700 53.700 183.800 ;
        RECT 50.200 183.100 50.600 183.500 ;
        RECT 51.900 183.400 53.700 183.700 ;
        RECT 52.300 183.100 52.600 183.400 ;
        RECT 55.000 183.100 55.400 183.500 ;
        RECT 49.900 181.100 50.500 183.100 ;
        RECT 52.200 181.100 52.600 183.100 ;
        RECT 54.400 182.800 55.400 183.100 ;
        RECT 54.400 181.100 54.800 182.800 ;
        RECT 56.600 181.100 57.000 185.300 ;
        RECT 57.400 185.200 59.300 185.500 ;
        RECT 57.400 183.500 57.700 185.200 ;
        RECT 60.000 184.900 60.300 186.800 ;
        RECT 63.700 186.200 64.000 186.800 ;
        RECT 64.300 186.500 65.000 186.900 ;
        RECT 68.600 186.900 69.100 187.100 ;
        RECT 69.600 187.200 69.900 187.500 ;
        RECT 60.600 185.400 61.000 186.200 ;
        RECT 63.000 185.400 63.400 186.200 ;
        RECT 63.700 185.800 64.200 186.200 ;
        RECT 59.500 184.600 60.300 184.900 ;
        RECT 63.700 184.900 64.000 185.800 ;
        RECT 64.700 185.500 65.000 186.500 ;
        RECT 65.400 185.800 65.800 186.600 ;
        RECT 66.200 185.800 66.600 186.600 ;
        RECT 67.000 185.800 67.400 186.600 ;
        RECT 67.800 185.800 68.200 186.600 ;
        RECT 68.600 186.500 69.300 186.900 ;
        RECT 69.600 186.800 70.600 187.200 ;
        RECT 71.800 187.100 72.200 187.200 ;
        RECT 72.600 187.100 73.000 187.200 ;
        RECT 71.800 186.800 73.000 187.100 ;
        RECT 68.600 185.500 68.900 186.500 ;
        RECT 64.700 185.200 66.600 185.500 ;
        RECT 63.700 184.600 64.500 184.900 ;
        RECT 57.400 181.500 57.800 183.500 ;
        RECT 59.500 182.200 59.900 184.600 ;
        RECT 59.000 181.800 59.900 182.200 ;
        RECT 59.500 181.100 59.900 181.800 ;
        RECT 64.100 181.100 64.500 184.600 ;
        RECT 66.300 183.500 66.600 185.200 ;
        RECT 66.200 181.500 66.600 183.500 ;
        RECT 67.000 185.200 68.900 185.500 ;
        RECT 67.000 183.500 67.300 185.200 ;
        RECT 69.600 184.900 69.900 186.800 ;
        RECT 72.700 186.600 73.000 186.800 ;
        RECT 72.700 186.200 73.100 186.600 ;
        RECT 73.400 186.200 73.700 187.900 ;
        RECT 75.800 187.500 76.200 189.900 ;
        RECT 78.000 189.200 78.400 189.900 ;
        RECT 77.400 188.900 78.400 189.200 ;
        RECT 80.200 188.900 80.600 189.900 ;
        RECT 82.300 189.200 82.900 189.900 ;
        RECT 82.200 188.900 82.900 189.200 ;
        RECT 77.400 188.500 77.800 188.900 ;
        RECT 80.200 188.600 80.500 188.900 ;
        RECT 78.200 188.200 78.600 188.600 ;
        RECT 79.100 188.300 80.500 188.600 ;
        RECT 82.200 188.500 82.600 188.900 ;
        RECT 79.100 188.200 79.500 188.300 ;
        RECT 74.200 186.400 74.600 187.200 ;
        RECT 76.200 187.100 77.000 187.200 ;
        RECT 78.300 187.100 78.600 188.200 ;
        RECT 83.100 187.700 83.500 187.800 ;
        RECT 84.600 187.700 85.000 189.900 ;
        RECT 86.700 188.200 87.100 189.900 ;
        RECT 83.100 187.400 85.000 187.700 ;
        RECT 86.200 187.900 87.100 188.200 ;
        RECT 87.800 187.900 88.200 189.900 ;
        RECT 88.600 188.000 89.000 189.900 ;
        RECT 90.200 188.000 90.600 189.900 ;
        RECT 92.300 188.200 92.700 189.900 ;
        RECT 88.600 187.900 90.600 188.000 ;
        RECT 91.800 187.900 92.700 188.200 ;
        RECT 93.400 187.900 93.800 189.900 ;
        RECT 94.200 188.000 94.600 189.900 ;
        RECT 95.800 188.000 96.200 189.900 ;
        RECT 98.500 188.000 98.900 189.500 ;
        RECT 100.600 188.500 101.000 189.500 ;
        RECT 94.200 187.900 96.200 188.000 ;
        RECT 79.000 187.100 79.400 187.200 ;
        RECT 81.100 187.100 81.500 187.200 ;
        RECT 76.200 186.800 81.700 187.100 ;
        RECT 77.700 186.700 78.100 186.800 ;
        RECT 76.900 186.200 77.300 186.300 ;
        RECT 70.200 186.100 70.600 186.200 ;
        RECT 71.000 186.100 71.400 186.200 ;
        RECT 70.200 185.800 71.400 186.100 ;
        RECT 70.200 185.400 70.600 185.800 ;
        RECT 71.800 185.400 72.200 186.200 ;
        RECT 73.400 185.800 73.800 186.200 ;
        RECT 75.000 186.100 75.400 186.200 ;
        RECT 74.600 185.800 75.400 186.100 ;
        RECT 76.900 186.100 79.400 186.200 ;
        RECT 79.800 186.100 80.200 186.200 ;
        RECT 76.900 185.900 80.200 186.100 ;
        RECT 79.000 185.800 80.200 185.900 ;
        RECT 73.400 185.700 73.700 185.800 ;
        RECT 72.700 185.400 73.700 185.700 ;
        RECT 74.600 185.600 75.000 185.800 ;
        RECT 75.800 185.500 78.600 185.600 ;
        RECT 75.800 185.400 78.700 185.500 ;
        RECT 72.700 185.100 73.000 185.400 ;
        RECT 75.800 185.300 80.700 185.400 ;
        RECT 69.100 184.600 69.900 184.900 ;
        RECT 67.000 181.500 67.400 183.500 ;
        RECT 69.100 183.200 69.500 184.600 ;
        RECT 68.600 182.800 69.500 183.200 ;
        RECT 69.100 181.100 69.500 182.800 ;
        RECT 71.800 181.400 72.200 185.100 ;
        RECT 72.600 181.700 73.000 185.100 ;
        RECT 73.400 184.800 75.400 185.100 ;
        RECT 73.400 181.400 73.800 184.800 ;
        RECT 71.800 181.100 73.800 181.400 ;
        RECT 75.000 181.100 75.400 184.800 ;
        RECT 75.800 181.100 76.200 185.300 ;
        RECT 78.300 185.100 80.700 185.300 ;
        RECT 77.400 184.500 80.100 184.800 ;
        RECT 77.400 184.400 77.800 184.500 ;
        RECT 79.700 184.400 80.100 184.500 ;
        RECT 80.400 184.500 80.700 185.100 ;
        RECT 81.400 185.200 81.700 186.800 ;
        RECT 82.200 186.400 82.600 186.500 ;
        RECT 82.200 186.100 84.100 186.400 ;
        RECT 83.700 186.000 84.100 186.100 ;
        RECT 82.900 185.700 83.300 185.800 ;
        RECT 84.600 185.700 85.000 187.400 ;
        RECT 85.400 186.800 85.800 187.600 ;
        RECT 82.900 185.400 85.000 185.700 ;
        RECT 81.400 184.900 82.600 185.200 ;
        RECT 81.100 184.500 81.500 184.600 ;
        RECT 80.400 184.200 81.500 184.500 ;
        RECT 82.300 184.400 82.600 184.900 ;
        RECT 82.300 184.000 83.000 184.400 ;
        RECT 79.100 183.700 79.500 183.800 ;
        RECT 80.500 183.700 80.900 183.800 ;
        RECT 77.400 183.100 77.800 183.500 ;
        RECT 79.100 183.400 80.900 183.700 ;
        RECT 80.200 183.100 80.500 183.400 ;
        RECT 82.200 183.100 82.600 183.500 ;
        RECT 77.400 182.800 78.400 183.100 ;
        RECT 78.000 181.100 78.400 182.800 ;
        RECT 80.200 181.100 80.600 183.100 ;
        RECT 82.300 181.100 82.900 183.100 ;
        RECT 84.600 181.100 85.000 185.400 ;
        RECT 86.200 186.100 86.600 187.900 ;
        RECT 87.900 187.200 88.200 187.900 ;
        RECT 88.700 187.700 90.500 187.900 ;
        RECT 89.800 187.200 90.200 187.400 ;
        RECT 87.800 186.800 89.100 187.200 ;
        RECT 89.800 186.900 90.600 187.200 ;
        RECT 90.200 186.800 90.600 186.900 ;
        RECT 91.000 186.800 91.400 187.600 ;
        RECT 86.200 185.800 88.100 186.100 ;
        RECT 86.200 181.100 86.600 185.800 ;
        RECT 87.800 185.200 88.100 185.800 ;
        RECT 87.000 184.400 87.400 185.200 ;
        RECT 87.800 185.100 88.200 185.200 ;
        RECT 88.800 185.100 89.100 186.800 ;
        RECT 89.400 185.800 89.800 186.600 ;
        RECT 91.800 186.100 92.200 187.900 ;
        RECT 93.500 187.200 93.800 187.900 ;
        RECT 94.300 187.700 96.100 187.900 ;
        RECT 98.100 187.700 98.900 188.000 ;
        RECT 98.100 187.500 98.500 187.700 ;
        RECT 95.400 187.200 95.800 187.400 ;
        RECT 98.100 187.200 98.400 187.500 ;
        RECT 100.700 187.400 101.000 188.500 ;
        RECT 103.000 187.500 103.400 189.900 ;
        RECT 105.200 189.200 105.600 189.900 ;
        RECT 104.600 188.900 105.600 189.200 ;
        RECT 107.400 188.900 107.800 189.900 ;
        RECT 109.500 189.200 110.100 189.900 ;
        RECT 109.400 188.900 110.100 189.200 ;
        RECT 104.600 188.500 105.000 188.900 ;
        RECT 107.400 188.600 107.700 188.900 ;
        RECT 105.400 188.200 105.800 188.600 ;
        RECT 106.300 188.300 107.700 188.600 ;
        RECT 109.400 188.500 109.800 188.900 ;
        RECT 106.300 188.200 106.700 188.300 ;
        RECT 93.400 186.800 94.700 187.200 ;
        RECT 95.400 186.900 96.200 187.200 ;
        RECT 95.800 186.800 96.200 186.900 ;
        RECT 97.400 186.800 98.400 187.200 ;
        RECT 98.900 187.100 101.000 187.400 ;
        RECT 103.400 187.100 104.200 187.200 ;
        RECT 105.500 187.100 105.800 188.200 ;
        RECT 110.300 187.700 110.700 187.800 ;
        RECT 111.800 187.700 112.200 189.900 ;
        RECT 113.900 188.200 114.300 189.900 ;
        RECT 110.200 187.400 112.200 187.700 ;
        RECT 113.400 187.900 114.300 188.200 ;
        RECT 115.000 187.900 115.400 189.900 ;
        RECT 115.800 188.000 116.200 189.900 ;
        RECT 117.400 188.000 117.800 189.900 ;
        RECT 115.800 187.900 117.800 188.000 ;
        RECT 118.200 188.000 118.600 189.900 ;
        RECT 119.800 188.000 120.200 189.900 ;
        RECT 118.200 187.900 120.200 188.000 ;
        RECT 120.600 187.900 121.000 189.900 ;
        RECT 108.300 187.100 108.700 187.200 ;
        RECT 98.900 186.900 99.400 187.100 ;
        RECT 91.800 185.800 93.700 186.100 ;
        RECT 87.800 184.800 88.500 185.100 ;
        RECT 88.800 184.800 89.300 185.100 ;
        RECT 88.200 184.200 88.500 184.800 ;
        RECT 88.200 183.800 88.600 184.200 ;
        RECT 88.900 181.100 89.300 184.800 ;
        RECT 91.800 181.100 92.200 185.800 ;
        RECT 93.400 185.200 93.700 185.800 ;
        RECT 92.600 184.400 93.000 185.200 ;
        RECT 93.400 185.100 93.800 185.200 ;
        RECT 94.400 185.100 94.700 186.800 ;
        RECT 95.000 185.800 95.400 186.600 ;
        RECT 96.600 186.100 97.000 186.200 ;
        RECT 97.400 186.100 97.800 186.200 ;
        RECT 96.600 185.800 97.800 186.100 ;
        RECT 97.400 185.400 97.800 185.800 ;
        RECT 93.400 184.800 94.100 185.100 ;
        RECT 94.400 184.800 94.900 185.100 ;
        RECT 93.800 184.200 94.100 184.800 ;
        RECT 93.800 183.800 94.200 184.200 ;
        RECT 94.500 181.100 94.900 184.800 ;
        RECT 98.100 184.900 98.400 186.800 ;
        RECT 98.700 186.500 99.400 186.900 ;
        RECT 103.400 186.800 108.900 187.100 ;
        RECT 110.200 186.800 110.600 187.400 ;
        RECT 111.800 187.100 112.200 187.400 ;
        RECT 112.600 187.100 113.000 187.600 ;
        RECT 111.800 186.800 113.000 187.100 ;
        RECT 104.900 186.700 105.300 186.800 ;
        RECT 99.100 185.500 99.400 186.500 ;
        RECT 99.800 185.800 100.200 186.600 ;
        RECT 100.600 186.100 101.000 186.600 ;
        RECT 104.100 186.200 104.500 186.300 ;
        RECT 101.400 186.100 101.800 186.200 ;
        RECT 100.600 185.800 101.800 186.100 ;
        RECT 104.100 185.900 106.600 186.200 ;
        RECT 106.200 185.800 106.600 185.900 ;
        RECT 103.000 185.500 105.800 185.600 ;
        RECT 99.100 185.200 101.000 185.500 ;
        RECT 98.100 184.600 98.900 184.900 ;
        RECT 98.500 182.200 98.900 184.600 ;
        RECT 100.700 183.500 101.000 185.200 ;
        RECT 98.200 181.800 98.900 182.200 ;
        RECT 98.500 181.100 98.900 181.800 ;
        RECT 100.600 181.500 101.000 183.500 ;
        RECT 103.000 185.400 105.900 185.500 ;
        RECT 103.000 185.300 107.900 185.400 ;
        RECT 103.000 181.100 103.400 185.300 ;
        RECT 105.500 185.100 107.900 185.300 ;
        RECT 104.600 184.500 107.300 184.800 ;
        RECT 104.600 184.400 105.000 184.500 ;
        RECT 106.900 184.400 107.300 184.500 ;
        RECT 107.600 184.500 107.900 185.100 ;
        RECT 108.600 185.200 108.900 186.800 ;
        RECT 109.400 186.400 109.800 186.500 ;
        RECT 109.400 186.100 111.300 186.400 ;
        RECT 110.900 186.000 111.300 186.100 ;
        RECT 110.100 185.700 110.500 185.800 ;
        RECT 111.800 185.700 112.200 186.800 ;
        RECT 110.100 185.400 112.200 185.700 ;
        RECT 108.600 184.900 109.800 185.200 ;
        RECT 108.300 184.500 108.700 184.600 ;
        RECT 107.600 184.200 108.700 184.500 ;
        RECT 109.500 184.400 109.800 184.900 ;
        RECT 109.500 184.000 110.200 184.400 ;
        RECT 106.300 183.700 106.700 183.800 ;
        RECT 107.700 183.700 108.100 183.800 ;
        RECT 104.600 183.100 105.000 183.500 ;
        RECT 106.300 183.400 108.100 183.700 ;
        RECT 107.400 183.100 107.700 183.400 ;
        RECT 109.400 183.100 109.800 183.500 ;
        RECT 104.600 182.800 105.600 183.100 ;
        RECT 105.200 181.100 105.600 182.800 ;
        RECT 107.400 181.100 107.800 183.100 ;
        RECT 109.500 181.100 110.100 183.100 ;
        RECT 111.800 181.100 112.200 185.400 ;
        RECT 113.400 186.100 113.800 187.900 ;
        RECT 115.100 187.200 115.400 187.900 ;
        RECT 115.900 187.700 117.700 187.900 ;
        RECT 118.300 187.700 120.100 187.900 ;
        RECT 117.000 187.200 117.400 187.400 ;
        RECT 118.600 187.200 119.000 187.400 ;
        RECT 120.600 187.200 120.900 187.900 ;
        RECT 121.400 187.700 121.800 189.900 ;
        RECT 123.500 189.200 124.100 189.900 ;
        RECT 123.500 188.900 124.200 189.200 ;
        RECT 125.800 188.900 126.200 189.900 ;
        RECT 128.000 189.200 128.400 189.900 ;
        RECT 128.000 188.900 129.000 189.200 ;
        RECT 123.800 188.500 124.200 188.900 ;
        RECT 125.900 188.600 126.200 188.900 ;
        RECT 125.900 188.300 127.300 188.600 ;
        RECT 126.900 188.200 127.300 188.300 ;
        RECT 127.800 188.200 128.200 188.600 ;
        RECT 128.600 188.500 129.000 188.900 ;
        RECT 122.900 187.700 123.300 187.800 ;
        RECT 121.400 187.400 123.300 187.700 ;
        RECT 114.200 187.100 114.600 187.200 ;
        RECT 115.000 187.100 116.300 187.200 ;
        RECT 114.200 186.800 116.300 187.100 ;
        RECT 117.000 187.100 117.800 187.200 ;
        RECT 118.200 187.100 119.000 187.200 ;
        RECT 117.000 186.900 119.000 187.100 ;
        RECT 117.400 186.800 118.600 186.900 ;
        RECT 119.700 186.800 121.000 187.200 ;
        RECT 113.400 185.800 115.300 186.100 ;
        RECT 113.400 181.100 113.800 185.800 ;
        RECT 115.000 185.200 115.300 185.800 ;
        RECT 114.200 184.400 114.600 185.200 ;
        RECT 115.000 185.100 115.400 185.200 ;
        RECT 116.000 185.100 116.300 186.800 ;
        RECT 116.600 186.100 117.000 186.600 ;
        RECT 118.200 186.100 118.600 186.200 ;
        RECT 116.600 185.800 118.600 186.100 ;
        RECT 119.000 185.800 119.400 186.600 ;
        RECT 119.700 186.100 120.000 186.800 ;
        RECT 120.600 186.100 121.000 186.200 ;
        RECT 119.700 185.800 121.000 186.100 ;
        RECT 119.700 185.100 120.000 185.800 ;
        RECT 121.400 185.700 121.800 187.400 ;
        RECT 124.900 187.100 125.300 187.200 ;
        RECT 127.000 187.100 127.400 187.200 ;
        RECT 127.800 187.100 128.100 188.200 ;
        RECT 130.200 187.500 130.600 189.900 ;
        RECT 131.000 188.000 131.400 189.900 ;
        RECT 132.600 188.000 133.000 189.900 ;
        RECT 131.000 187.900 133.000 188.000 ;
        RECT 133.400 187.900 133.800 189.900 ;
        RECT 131.100 187.700 132.900 187.900 ;
        RECT 131.400 187.200 131.800 187.400 ;
        RECT 133.400 187.200 133.700 187.900 ;
        RECT 135.000 187.600 135.400 189.900 ;
        RECT 136.600 187.600 137.000 189.900 ;
        RECT 138.200 187.600 138.600 189.900 ;
        RECT 139.800 187.600 140.200 189.900 ;
        RECT 142.200 188.900 142.600 189.900 ;
        RECT 141.400 187.800 141.800 188.600 ;
        RECT 142.300 188.100 142.600 188.900 ;
        RECT 143.900 188.200 144.300 188.600 ;
        RECT 143.800 188.100 144.200 188.200 ;
        RECT 142.200 187.800 144.200 188.100 ;
        RECT 144.600 187.900 145.000 189.900 ;
        RECT 147.300 189.200 147.700 189.900 ;
        RECT 147.000 188.800 147.700 189.200 ;
        RECT 147.300 188.200 147.700 188.800 ;
        RECT 147.300 187.900 148.200 188.200 ;
        RECT 152.500 187.900 153.300 189.900 ;
        RECT 134.200 187.200 135.400 187.600 ;
        RECT 135.900 187.200 137.000 187.600 ;
        RECT 137.500 187.200 138.600 187.600 ;
        RECT 139.300 187.200 140.200 187.600 ;
        RECT 142.300 187.200 142.600 187.800 ;
        RECT 129.400 187.100 130.200 187.200 ;
        RECT 124.700 186.800 130.200 187.100 ;
        RECT 131.000 186.900 131.800 187.200 ;
        RECT 131.000 186.800 131.400 186.900 ;
        RECT 132.500 186.800 133.800 187.200 ;
        RECT 123.800 186.400 124.200 186.500 ;
        RECT 122.300 186.100 124.200 186.400 ;
        RECT 122.300 186.000 122.700 186.100 ;
        RECT 123.100 185.700 123.500 185.800 ;
        RECT 121.400 185.400 123.500 185.700 ;
        RECT 120.600 185.100 121.000 185.200 ;
        RECT 115.000 184.800 115.700 185.100 ;
        RECT 116.000 184.800 116.500 185.100 ;
        RECT 115.400 184.200 115.700 184.800 ;
        RECT 115.400 183.800 115.800 184.200 ;
        RECT 116.100 181.100 116.500 184.800 ;
        RECT 119.500 184.800 120.000 185.100 ;
        RECT 120.300 184.800 121.000 185.100 ;
        RECT 119.500 181.100 119.900 184.800 ;
        RECT 120.300 184.200 120.600 184.800 ;
        RECT 120.200 183.800 120.600 184.200 ;
        RECT 121.400 181.100 121.800 185.400 ;
        RECT 124.700 185.200 125.000 186.800 ;
        RECT 128.300 186.700 128.700 186.800 ;
        RECT 129.100 186.200 129.500 186.300 ;
        RECT 126.200 186.100 126.600 186.200 ;
        RECT 127.000 186.100 129.500 186.200 ;
        RECT 126.200 185.900 129.500 186.100 ;
        RECT 126.200 185.800 127.400 185.900 ;
        RECT 131.800 185.800 132.200 186.600 ;
        RECT 127.800 185.500 130.600 185.600 ;
        RECT 127.700 185.400 130.600 185.500 ;
        RECT 123.800 184.900 125.000 185.200 ;
        RECT 125.700 185.300 130.600 185.400 ;
        RECT 125.700 185.100 128.100 185.300 ;
        RECT 123.800 184.400 124.100 184.900 ;
        RECT 123.400 184.000 124.100 184.400 ;
        RECT 124.900 184.500 125.300 184.600 ;
        RECT 125.700 184.500 126.000 185.100 ;
        RECT 124.900 184.200 126.000 184.500 ;
        RECT 126.300 184.500 129.000 184.800 ;
        RECT 126.300 184.400 126.700 184.500 ;
        RECT 128.600 184.400 129.000 184.500 ;
        RECT 125.500 183.700 125.900 183.800 ;
        RECT 126.900 183.700 127.300 183.800 ;
        RECT 123.800 183.100 124.200 183.500 ;
        RECT 125.500 183.400 127.300 183.700 ;
        RECT 125.900 183.100 126.200 183.400 ;
        RECT 128.600 183.100 129.000 183.500 ;
        RECT 123.500 181.100 124.100 183.100 ;
        RECT 125.800 181.100 126.200 183.100 ;
        RECT 128.000 182.800 129.000 183.100 ;
        RECT 128.000 181.100 128.400 182.800 ;
        RECT 130.200 181.100 130.600 185.300 ;
        RECT 132.500 185.100 132.800 186.800 ;
        RECT 134.200 185.800 134.600 187.200 ;
        RECT 135.900 186.900 136.300 187.200 ;
        RECT 137.500 186.900 137.900 187.200 ;
        RECT 139.300 186.900 139.700 187.200 ;
        RECT 140.600 186.900 141.000 187.200 ;
        RECT 135.000 186.500 136.300 186.900 ;
        RECT 136.700 186.500 137.900 186.900 ;
        RECT 138.400 186.500 139.700 186.900 ;
        RECT 140.100 186.500 141.000 186.900 ;
        RECT 142.200 186.800 142.600 187.200 ;
        RECT 135.900 185.800 136.300 186.500 ;
        RECT 137.500 185.800 137.900 186.500 ;
        RECT 139.300 185.800 139.700 186.500 ;
        RECT 134.200 185.400 135.400 185.800 ;
        RECT 135.900 185.400 137.000 185.800 ;
        RECT 137.500 185.400 138.600 185.800 ;
        RECT 139.300 185.400 140.200 185.800 ;
        RECT 133.400 185.100 133.800 185.200 ;
        RECT 132.300 184.800 132.800 185.100 ;
        RECT 133.100 184.800 133.800 185.100 ;
        RECT 132.300 181.100 132.700 184.800 ;
        RECT 133.100 184.200 133.400 184.800 ;
        RECT 133.000 183.800 133.400 184.200 ;
        RECT 135.000 181.100 135.400 185.400 ;
        RECT 136.600 181.100 137.000 185.400 ;
        RECT 138.200 181.100 138.600 185.400 ;
        RECT 139.800 181.100 140.200 185.400 ;
        RECT 142.300 185.100 142.600 186.800 ;
        RECT 143.000 185.400 143.400 186.200 ;
        RECT 143.800 186.100 144.200 186.200 ;
        RECT 144.700 186.100 145.000 187.900 ;
        RECT 145.400 186.400 145.800 187.200 ;
        RECT 146.200 186.100 146.600 186.200 ;
        RECT 143.800 185.800 145.000 186.100 ;
        RECT 145.800 185.800 146.600 186.100 ;
        RECT 143.900 185.100 144.200 185.800 ;
        RECT 145.800 185.600 146.200 185.800 ;
        RECT 142.200 184.700 143.100 185.100 ;
        RECT 142.700 181.100 143.100 184.700 ;
        RECT 143.800 181.100 144.200 185.100 ;
        RECT 144.600 184.800 146.600 185.100 ;
        RECT 144.600 181.100 145.000 184.800 ;
        RECT 146.200 181.100 146.600 184.800 ;
        RECT 147.000 184.400 147.400 185.200 ;
        RECT 147.800 181.100 148.200 187.900 ;
        RECT 148.600 186.800 149.000 187.600 ;
        RECT 151.800 186.400 152.200 187.200 ;
        RECT 152.700 186.200 153.000 187.900 ;
        RECT 155.000 187.600 155.400 189.900 ;
        RECT 156.600 188.200 157.000 189.900 ;
        RECT 158.500 189.200 158.900 189.900 ;
        RECT 158.200 188.800 158.900 189.200 ;
        RECT 158.500 188.200 158.900 188.800 ;
        RECT 161.900 188.200 162.300 189.900 ;
        RECT 156.600 187.900 157.100 188.200 ;
        RECT 158.500 187.900 159.400 188.200 ;
        RECT 155.000 187.300 156.300 187.600 ;
        RECT 153.400 186.800 153.800 187.200 ;
        RECT 153.400 186.600 153.700 186.800 ;
        RECT 153.300 186.200 153.700 186.600 ;
        RECT 155.100 186.200 155.500 186.600 ;
        RECT 151.000 186.100 151.400 186.200 ;
        RECT 151.000 185.800 151.800 186.100 ;
        RECT 152.600 185.800 153.000 186.200 ;
        RECT 151.400 185.600 151.800 185.800 ;
        RECT 152.700 185.700 153.000 185.800 ;
        RECT 152.700 185.400 153.700 185.700 ;
        RECT 154.200 185.400 154.600 186.200 ;
        RECT 155.000 185.800 155.500 186.200 ;
        RECT 156.000 186.500 156.300 187.300 ;
        RECT 156.800 187.200 157.100 187.900 ;
        RECT 156.600 187.100 157.100 187.200 ;
        RECT 156.600 186.800 158.500 187.100 ;
        RECT 156.000 186.100 156.500 186.500 ;
        RECT 153.400 185.100 153.700 185.400 ;
        RECT 156.000 185.100 156.300 186.100 ;
        RECT 156.800 185.100 157.100 186.800 ;
        RECT 158.200 186.200 158.500 186.800 ;
        RECT 158.200 185.800 158.600 186.200 ;
        RECT 151.000 184.800 153.000 185.100 ;
        RECT 151.000 181.100 151.400 184.800 ;
        RECT 152.600 181.400 153.000 184.800 ;
        RECT 153.400 181.700 153.800 185.100 ;
        RECT 154.200 181.400 154.600 185.100 ;
        RECT 152.600 181.100 154.600 181.400 ;
        RECT 155.000 184.800 156.300 185.100 ;
        RECT 155.000 181.100 155.400 184.800 ;
        RECT 156.600 184.600 157.100 185.100 ;
        RECT 156.600 181.100 157.000 184.600 ;
        RECT 158.200 184.400 158.600 185.200 ;
        RECT 159.000 181.100 159.400 187.900 ;
        RECT 161.400 187.900 162.300 188.200 ;
        RECT 163.000 188.000 163.400 189.900 ;
        RECT 164.600 188.000 165.000 189.900 ;
        RECT 163.000 187.900 165.000 188.000 ;
        RECT 165.400 187.900 165.800 189.900 ;
        RECT 159.800 186.800 160.200 187.600 ;
        RECT 160.600 186.800 161.000 187.600 ;
        RECT 161.400 181.100 161.800 187.900 ;
        RECT 163.100 187.700 164.900 187.900 ;
        RECT 163.400 187.200 163.800 187.400 ;
        RECT 165.400 187.200 165.700 187.900 ;
        RECT 166.200 187.700 166.600 189.900 ;
        RECT 168.300 189.200 168.900 189.900 ;
        RECT 168.300 188.900 169.000 189.200 ;
        RECT 170.600 188.900 171.000 189.900 ;
        RECT 172.800 189.200 173.200 189.900 ;
        RECT 172.800 188.900 173.800 189.200 ;
        RECT 168.600 188.500 169.000 188.900 ;
        RECT 170.700 188.600 171.000 188.900 ;
        RECT 170.700 188.300 172.100 188.600 ;
        RECT 171.700 188.200 172.100 188.300 ;
        RECT 172.600 188.200 173.000 188.600 ;
        RECT 173.400 188.500 173.800 188.900 ;
        RECT 167.700 187.700 168.100 187.800 ;
        RECT 166.200 187.400 168.100 187.700 ;
        RECT 163.000 186.900 163.800 187.200 ;
        RECT 163.000 186.800 163.400 186.900 ;
        RECT 164.500 186.800 165.800 187.200 ;
        RECT 163.800 186.100 164.200 186.600 ;
        RECT 162.200 185.800 164.200 186.100 ;
        RECT 162.200 185.200 162.500 185.800 ;
        RECT 162.200 183.800 162.600 185.200 ;
        RECT 164.500 185.100 164.800 186.800 ;
        RECT 166.200 185.700 166.600 187.400 ;
        RECT 169.700 187.100 170.100 187.200 ;
        RECT 171.800 187.100 172.200 187.200 ;
        RECT 172.600 187.100 172.900 188.200 ;
        RECT 175.000 187.500 175.400 189.900 ;
        RECT 175.800 188.500 176.200 189.500 ;
        RECT 175.800 187.400 176.100 188.500 ;
        RECT 177.900 188.000 178.300 189.500 ;
        RECT 180.600 188.000 181.000 189.900 ;
        RECT 182.200 188.000 182.600 189.900 ;
        RECT 177.900 187.700 178.700 188.000 ;
        RECT 180.600 187.900 182.600 188.000 ;
        RECT 183.000 187.900 183.400 189.900 ;
        RECT 184.100 188.200 184.500 189.900 ;
        RECT 187.500 189.200 188.300 189.900 ;
        RECT 187.000 188.800 188.300 189.200 ;
        RECT 184.100 187.900 185.000 188.200 ;
        RECT 187.500 187.900 188.300 188.800 ;
        RECT 180.700 187.700 182.500 187.900 ;
        RECT 178.300 187.500 178.700 187.700 ;
        RECT 174.200 187.100 175.000 187.200 ;
        RECT 175.800 187.100 177.900 187.400 ;
        RECT 169.500 186.800 175.000 187.100 ;
        RECT 177.400 186.900 177.900 187.100 ;
        RECT 178.400 187.200 178.700 187.500 ;
        RECT 181.000 187.200 181.400 187.400 ;
        RECT 183.000 187.200 183.300 187.900 ;
        RECT 168.600 186.400 169.000 186.500 ;
        RECT 167.100 186.100 169.000 186.400 ;
        RECT 167.100 186.000 167.500 186.100 ;
        RECT 167.900 185.700 168.300 185.800 ;
        RECT 166.200 185.400 168.300 185.700 ;
        RECT 165.400 185.100 165.800 185.200 ;
        RECT 164.300 184.800 164.800 185.100 ;
        RECT 165.100 184.800 165.800 185.100 ;
        RECT 164.300 181.100 164.700 184.800 ;
        RECT 165.100 184.200 165.400 184.800 ;
        RECT 165.000 183.800 165.400 184.200 ;
        RECT 166.200 181.100 166.600 185.400 ;
        RECT 169.500 185.200 169.800 186.800 ;
        RECT 173.100 186.700 173.500 186.800 ;
        RECT 173.900 186.200 174.300 186.300 ;
        RECT 170.200 186.100 170.600 186.200 ;
        RECT 171.800 186.100 174.300 186.200 ;
        RECT 170.200 185.900 174.300 186.100 ;
        RECT 170.200 185.800 172.200 185.900 ;
        RECT 175.800 185.800 176.200 186.600 ;
        RECT 176.600 185.800 177.000 186.600 ;
        RECT 177.400 186.500 178.100 186.900 ;
        RECT 178.400 186.800 179.400 187.200 ;
        RECT 180.600 186.900 181.400 187.200 ;
        RECT 182.100 187.100 183.400 187.200 ;
        RECT 183.800 187.100 184.200 187.200 ;
        RECT 180.600 186.800 181.000 186.900 ;
        RECT 182.100 186.800 184.200 187.100 ;
        RECT 172.600 185.500 175.400 185.600 ;
        RECT 177.400 185.500 177.700 186.500 ;
        RECT 172.500 185.400 175.400 185.500 ;
        RECT 168.600 184.900 169.800 185.200 ;
        RECT 170.500 185.300 175.400 185.400 ;
        RECT 170.500 185.100 172.900 185.300 ;
        RECT 168.600 184.400 168.900 184.900 ;
        RECT 168.200 184.200 168.900 184.400 ;
        RECT 169.700 184.500 170.100 184.600 ;
        RECT 170.500 184.500 170.800 185.100 ;
        RECT 169.700 184.200 170.800 184.500 ;
        RECT 171.100 184.500 173.800 184.800 ;
        RECT 171.100 184.400 171.500 184.500 ;
        RECT 173.400 184.400 173.800 184.500 ;
        RECT 167.800 184.000 168.900 184.200 ;
        RECT 167.800 183.800 168.500 184.000 ;
        RECT 170.300 183.700 170.700 183.800 ;
        RECT 171.700 183.700 172.100 183.800 ;
        RECT 168.600 183.100 169.000 183.500 ;
        RECT 170.300 183.400 172.100 183.700 ;
        RECT 170.700 183.100 171.000 183.400 ;
        RECT 173.400 183.100 173.800 183.500 ;
        RECT 168.300 181.100 168.900 183.100 ;
        RECT 170.600 181.100 171.000 183.100 ;
        RECT 172.800 182.800 173.800 183.100 ;
        RECT 172.800 181.100 173.200 182.800 ;
        RECT 175.000 181.100 175.400 185.300 ;
        RECT 175.800 185.200 177.700 185.500 ;
        RECT 175.800 183.500 176.100 185.200 ;
        RECT 178.400 184.900 178.700 186.800 ;
        RECT 179.000 185.400 179.400 186.200 ;
        RECT 181.400 185.800 181.800 186.600 ;
        RECT 182.100 185.100 182.400 186.800 ;
        RECT 184.600 186.100 185.000 187.900 ;
        RECT 185.400 187.100 185.800 187.600 ;
        RECT 186.200 187.100 186.600 187.200 ;
        RECT 185.400 186.800 186.600 187.100 ;
        RECT 187.000 186.800 187.400 187.200 ;
        RECT 187.100 186.600 187.400 186.800 ;
        RECT 187.100 186.200 187.500 186.600 ;
        RECT 187.800 186.200 188.100 187.900 ;
        RECT 190.200 187.700 190.600 189.900 ;
        RECT 192.300 189.200 192.900 189.900 ;
        RECT 192.300 188.900 193.000 189.200 ;
        RECT 194.600 188.900 195.000 189.900 ;
        RECT 196.800 189.200 197.200 189.900 ;
        RECT 196.800 188.900 197.800 189.200 ;
        RECT 192.600 188.500 193.000 188.900 ;
        RECT 194.700 188.600 195.000 188.900 ;
        RECT 194.700 188.300 196.100 188.600 ;
        RECT 195.700 188.200 196.100 188.300 ;
        RECT 196.600 188.200 197.000 188.600 ;
        RECT 197.400 188.500 197.800 188.900 ;
        RECT 191.700 187.700 192.100 187.800 ;
        RECT 190.200 187.400 192.100 187.700 ;
        RECT 188.600 186.400 189.000 187.200 ;
        RECT 183.000 185.800 185.000 186.100 ;
        RECT 183.000 185.200 183.300 185.800 ;
        RECT 183.000 185.100 183.400 185.200 ;
        RECT 177.900 184.600 178.700 184.900 ;
        RECT 181.900 184.800 182.400 185.100 ;
        RECT 182.700 184.800 183.400 185.100 ;
        RECT 175.800 181.500 176.200 183.500 ;
        RECT 177.900 183.200 178.300 184.600 ;
        RECT 177.400 182.800 178.300 183.200 ;
        RECT 177.900 181.100 178.300 182.800 ;
        RECT 181.900 181.100 182.300 184.800 ;
        RECT 182.700 184.200 183.000 184.800 ;
        RECT 183.800 184.400 184.200 185.200 ;
        RECT 182.600 183.800 183.000 184.200 ;
        RECT 184.600 181.100 185.000 185.800 ;
        RECT 186.200 185.400 186.600 186.200 ;
        RECT 187.800 185.800 188.200 186.200 ;
        RECT 189.400 186.100 189.800 186.200 ;
        RECT 189.000 185.800 189.800 186.100 ;
        RECT 187.800 185.700 188.100 185.800 ;
        RECT 187.100 185.400 188.100 185.700 ;
        RECT 189.000 185.600 189.400 185.800 ;
        RECT 190.200 185.700 190.600 187.400 ;
        RECT 193.700 187.100 194.100 187.200 ;
        RECT 196.600 187.100 196.900 188.200 ;
        RECT 199.000 187.500 199.400 189.900 ;
        RECT 200.100 189.200 200.500 189.900 ;
        RECT 200.100 188.800 201.000 189.200 ;
        RECT 203.000 189.100 203.400 189.200 ;
        RECT 203.800 189.100 204.200 189.900 ;
        RECT 203.000 188.800 204.200 189.100 ;
        RECT 205.900 189.200 206.500 189.900 ;
        RECT 205.900 188.900 206.600 189.200 ;
        RECT 208.200 188.900 208.600 189.900 ;
        RECT 210.400 189.200 210.800 189.900 ;
        RECT 210.400 188.900 211.400 189.200 ;
        RECT 200.100 188.200 200.500 188.800 ;
        RECT 200.100 187.900 201.000 188.200 ;
        RECT 198.200 187.100 199.000 187.200 ;
        RECT 193.500 186.800 199.000 187.100 ;
        RECT 192.600 186.400 193.000 186.500 ;
        RECT 191.100 186.100 193.000 186.400 ;
        RECT 191.100 186.000 191.500 186.100 ;
        RECT 191.900 185.700 192.300 185.800 ;
        RECT 190.200 185.400 192.300 185.700 ;
        RECT 187.100 185.100 187.400 185.400 ;
        RECT 186.200 181.400 186.600 185.100 ;
        RECT 187.000 181.700 187.400 185.100 ;
        RECT 187.800 184.800 189.800 185.100 ;
        RECT 187.800 181.400 188.200 184.800 ;
        RECT 186.200 181.100 188.200 181.400 ;
        RECT 189.400 181.100 189.800 184.800 ;
        RECT 190.200 181.100 190.600 185.400 ;
        RECT 193.500 185.200 193.800 186.800 ;
        RECT 197.100 186.700 197.500 186.800 ;
        RECT 197.900 186.200 198.300 186.300 ;
        RECT 195.800 185.900 198.300 186.200 ;
        RECT 195.800 185.800 196.200 185.900 ;
        RECT 196.600 185.500 199.400 185.600 ;
        RECT 196.500 185.400 199.400 185.500 ;
        RECT 192.600 184.900 193.800 185.200 ;
        RECT 194.500 185.300 199.400 185.400 ;
        RECT 194.500 185.100 196.900 185.300 ;
        RECT 192.600 184.400 192.900 184.900 ;
        RECT 192.200 184.200 192.900 184.400 ;
        RECT 193.700 184.500 194.100 184.600 ;
        RECT 194.500 184.500 194.800 185.100 ;
        RECT 193.700 184.200 194.800 184.500 ;
        RECT 195.100 184.500 197.800 184.800 ;
        RECT 195.100 184.400 195.500 184.500 ;
        RECT 197.400 184.400 197.800 184.500 ;
        RECT 191.800 184.000 192.900 184.200 ;
        RECT 191.800 183.800 192.500 184.000 ;
        RECT 194.300 183.700 194.700 183.800 ;
        RECT 195.700 183.700 196.100 183.800 ;
        RECT 192.600 183.100 193.000 183.500 ;
        RECT 194.300 183.400 196.100 183.700 ;
        RECT 194.700 183.100 195.000 183.400 ;
        RECT 197.400 183.100 197.800 183.500 ;
        RECT 192.300 181.100 192.900 183.100 ;
        RECT 194.600 181.100 195.000 183.100 ;
        RECT 196.800 182.800 197.800 183.100 ;
        RECT 196.800 181.100 197.200 182.800 ;
        RECT 199.000 181.100 199.400 185.300 ;
        RECT 199.800 184.400 200.200 185.200 ;
        RECT 200.600 181.100 201.000 187.900 ;
        RECT 203.800 187.700 204.200 188.800 ;
        RECT 206.200 188.500 206.600 188.900 ;
        RECT 208.300 188.600 208.600 188.900 ;
        RECT 208.300 188.300 209.700 188.600 ;
        RECT 209.300 188.200 209.700 188.300 ;
        RECT 210.200 188.200 210.600 188.600 ;
        RECT 211.000 188.500 211.400 188.900 ;
        RECT 207.000 187.800 207.400 188.200 ;
        RECT 205.300 187.700 205.700 187.800 ;
        RECT 201.400 187.100 201.800 187.600 ;
        RECT 203.800 187.400 205.700 187.700 ;
        RECT 203.000 187.100 203.400 187.200 ;
        RECT 201.400 186.800 203.400 187.100 ;
        RECT 203.800 185.700 204.200 187.400 ;
        RECT 207.000 187.200 207.300 187.800 ;
        RECT 207.000 187.100 207.700 187.200 ;
        RECT 210.200 187.100 210.500 188.200 ;
        RECT 212.600 187.500 213.000 189.900 ;
        RECT 214.700 189.200 215.100 189.900 ;
        RECT 214.700 188.800 215.400 189.200 ;
        RECT 214.700 188.200 215.100 188.800 ;
        RECT 214.200 187.900 215.100 188.200 ;
        RECT 215.800 188.500 216.200 189.500 ;
        RECT 211.800 187.100 212.600 187.200 ;
        RECT 207.000 186.800 212.600 187.100 ;
        RECT 213.400 186.800 213.800 187.600 ;
        RECT 206.200 186.400 206.600 186.500 ;
        RECT 204.700 186.100 206.600 186.400 ;
        RECT 204.700 186.000 205.100 186.100 ;
        RECT 205.500 185.700 205.900 185.800 ;
        RECT 203.800 185.400 205.900 185.700 ;
        RECT 203.800 181.100 204.200 185.400 ;
        RECT 207.100 185.200 207.400 186.800 ;
        RECT 210.700 186.700 211.100 186.800 ;
        RECT 211.500 186.200 211.900 186.300 ;
        RECT 207.800 186.100 208.200 186.200 ;
        RECT 209.400 186.100 211.900 186.200 ;
        RECT 207.800 185.900 211.900 186.100 ;
        RECT 207.800 185.800 209.800 185.900 ;
        RECT 210.200 185.500 213.000 185.600 ;
        RECT 210.100 185.400 213.000 185.500 ;
        RECT 206.200 184.900 207.400 185.200 ;
        RECT 208.100 185.300 213.000 185.400 ;
        RECT 208.100 185.100 210.500 185.300 ;
        RECT 206.200 184.400 206.500 184.900 ;
        RECT 205.800 184.000 206.500 184.400 ;
        RECT 207.300 184.500 207.700 184.600 ;
        RECT 208.100 184.500 208.400 185.100 ;
        RECT 207.300 184.200 208.400 184.500 ;
        RECT 208.700 184.500 211.400 184.800 ;
        RECT 208.700 184.400 209.100 184.500 ;
        RECT 211.000 184.400 211.400 184.500 ;
        RECT 207.900 183.700 208.300 183.800 ;
        RECT 209.300 183.700 209.700 183.800 ;
        RECT 206.200 183.100 206.600 183.500 ;
        RECT 207.900 183.400 209.700 183.700 ;
        RECT 208.300 183.100 208.600 183.400 ;
        RECT 211.000 183.100 211.400 183.500 ;
        RECT 205.900 181.100 206.500 183.100 ;
        RECT 208.200 181.100 208.600 183.100 ;
        RECT 210.400 182.800 211.400 183.100 ;
        RECT 210.400 181.100 210.800 182.800 ;
        RECT 212.600 181.100 213.000 185.300 ;
        RECT 214.200 181.100 214.600 187.900 ;
        RECT 215.800 187.400 216.100 188.500 ;
        RECT 217.900 188.000 218.300 189.500 ;
        RECT 222.500 188.000 222.900 189.500 ;
        RECT 224.600 188.500 225.000 189.500 ;
        RECT 217.900 187.700 218.700 188.000 ;
        RECT 218.300 187.500 218.700 187.700 ;
        RECT 215.800 187.100 217.900 187.400 ;
        RECT 217.400 186.900 217.900 187.100 ;
        RECT 218.400 187.200 218.700 187.500 ;
        RECT 222.100 187.700 222.900 188.000 ;
        RECT 222.100 187.500 222.500 187.700 ;
        RECT 222.100 187.200 222.400 187.500 ;
        RECT 224.700 187.400 225.000 188.500 ;
        RECT 225.400 188.000 225.800 189.900 ;
        RECT 227.000 188.000 227.400 189.900 ;
        RECT 225.400 187.900 227.400 188.000 ;
        RECT 227.800 187.900 228.200 189.900 ;
        RECT 228.900 188.200 229.300 189.900 ;
        RECT 228.900 187.900 229.800 188.200 ;
        RECT 225.500 187.700 227.300 187.900 ;
        RECT 215.800 185.800 216.200 186.600 ;
        RECT 216.600 185.800 217.000 186.600 ;
        RECT 217.400 186.500 218.100 186.900 ;
        RECT 218.400 186.800 219.400 187.200 ;
        RECT 219.800 187.100 220.200 187.200 ;
        RECT 221.400 187.100 222.400 187.200 ;
        RECT 219.800 186.800 222.400 187.100 ;
        RECT 222.900 187.100 225.000 187.400 ;
        RECT 225.800 187.200 226.200 187.400 ;
        RECT 227.800 187.200 228.100 187.900 ;
        RECT 222.900 186.900 223.400 187.100 ;
        RECT 217.400 185.500 217.700 186.500 ;
        RECT 215.800 185.200 217.700 185.500 ;
        RECT 215.000 184.400 215.400 185.200 ;
        RECT 215.800 183.500 216.100 185.200 ;
        RECT 218.400 184.900 218.700 186.800 ;
        RECT 219.000 186.100 219.400 186.200 ;
        RECT 220.600 186.100 221.000 186.200 ;
        RECT 219.000 185.800 221.000 186.100 ;
        RECT 219.000 185.400 219.400 185.800 ;
        RECT 221.400 185.400 221.800 186.200 ;
        RECT 217.900 184.600 218.700 184.900 ;
        RECT 222.100 184.900 222.400 186.800 ;
        RECT 222.700 186.500 223.400 186.900 ;
        RECT 225.400 186.900 226.200 187.200 ;
        RECT 226.900 187.100 228.200 187.200 ;
        RECT 228.600 187.100 229.000 187.200 ;
        RECT 225.400 186.800 225.800 186.900 ;
        RECT 226.900 186.800 229.000 187.100 ;
        RECT 223.100 185.500 223.400 186.500 ;
        RECT 223.800 185.800 224.200 186.600 ;
        RECT 224.600 185.800 225.000 186.600 ;
        RECT 226.200 185.800 226.600 186.600 ;
        RECT 223.100 185.200 225.000 185.500 ;
        RECT 222.100 184.600 222.900 184.900 ;
        RECT 215.800 181.500 216.200 183.500 ;
        RECT 217.900 182.200 218.300 184.600 ;
        RECT 217.400 181.800 218.300 182.200 ;
        RECT 217.900 181.100 218.300 181.800 ;
        RECT 222.500 181.100 222.900 184.600 ;
        RECT 224.700 183.500 225.000 185.200 ;
        RECT 226.900 185.100 227.200 186.800 ;
        RECT 229.400 186.100 229.800 187.900 ;
        RECT 230.200 186.800 230.600 187.600 ;
        RECT 231.000 187.500 231.400 189.900 ;
        RECT 233.200 189.200 233.600 189.900 ;
        RECT 232.600 188.900 233.600 189.200 ;
        RECT 235.400 188.900 235.800 189.900 ;
        RECT 237.500 189.200 238.100 189.900 ;
        RECT 237.400 188.900 238.100 189.200 ;
        RECT 232.600 188.500 233.000 188.900 ;
        RECT 235.400 188.600 235.700 188.900 ;
        RECT 233.400 187.800 233.800 188.600 ;
        RECT 234.300 188.300 235.700 188.600 ;
        RECT 237.400 188.500 237.800 188.900 ;
        RECT 234.300 188.200 234.700 188.300 ;
        RECT 231.400 187.100 232.200 187.200 ;
        RECT 233.500 187.100 233.800 187.800 ;
        RECT 238.300 187.700 238.700 187.800 ;
        RECT 239.800 187.700 240.200 189.900 ;
        RECT 238.300 187.400 240.200 187.700 ;
        RECT 241.400 187.600 241.800 189.900 ;
        RECT 243.000 187.600 243.400 189.900 ;
        RECT 244.600 187.600 245.000 189.900 ;
        RECT 246.200 187.600 246.600 189.900 ;
        RECT 248.600 188.200 249.000 189.900 ;
        RECT 236.300 187.100 236.700 187.200 ;
        RECT 231.400 186.800 236.900 187.100 ;
        RECT 232.900 186.700 233.300 186.800 ;
        RECT 227.800 185.800 229.800 186.100 ;
        RECT 232.100 186.200 232.500 186.300 ;
        RECT 233.400 186.200 233.800 186.300 ;
        RECT 232.100 185.900 234.600 186.200 ;
        RECT 234.200 185.800 234.600 185.900 ;
        RECT 227.800 185.200 228.100 185.800 ;
        RECT 227.800 185.100 228.200 185.200 ;
        RECT 224.600 181.500 225.000 183.500 ;
        RECT 226.700 184.800 227.200 185.100 ;
        RECT 227.500 184.800 228.200 185.100 ;
        RECT 226.700 181.100 227.100 184.800 ;
        RECT 227.500 184.200 227.800 184.800 ;
        RECT 228.600 184.400 229.000 185.200 ;
        RECT 227.400 183.800 227.800 184.200 ;
        RECT 229.400 181.100 229.800 185.800 ;
        RECT 231.000 185.500 233.800 185.600 ;
        RECT 231.000 185.400 233.900 185.500 ;
        RECT 231.000 185.300 235.900 185.400 ;
        RECT 231.000 181.100 231.400 185.300 ;
        RECT 233.500 185.100 235.900 185.300 ;
        RECT 232.600 184.500 235.300 184.800 ;
        RECT 232.600 184.400 233.000 184.500 ;
        RECT 234.900 184.400 235.300 184.500 ;
        RECT 235.600 184.500 235.900 185.100 ;
        RECT 236.600 185.200 236.900 186.800 ;
        RECT 237.400 186.400 237.800 186.500 ;
        RECT 237.400 186.100 239.300 186.400 ;
        RECT 238.900 186.000 239.300 186.100 ;
        RECT 238.100 185.700 238.500 185.800 ;
        RECT 239.800 185.700 240.200 187.400 ;
        RECT 238.100 185.400 240.200 185.700 ;
        RECT 240.600 187.200 241.800 187.600 ;
        RECT 242.300 187.200 243.400 187.600 ;
        RECT 243.900 187.200 245.000 187.600 ;
        RECT 245.700 187.200 246.600 187.600 ;
        RECT 248.500 187.900 249.000 188.200 ;
        RECT 248.500 187.200 248.800 187.900 ;
        RECT 250.200 187.600 250.600 189.900 ;
        RECT 249.300 187.300 250.600 187.600 ;
        RECT 240.600 185.800 241.000 187.200 ;
        RECT 242.300 186.900 242.700 187.200 ;
        RECT 243.900 186.900 244.300 187.200 ;
        RECT 245.700 186.900 246.100 187.200 ;
        RECT 241.400 186.500 242.700 186.900 ;
        RECT 243.100 186.500 244.300 186.900 ;
        RECT 244.800 186.500 246.100 186.900 ;
        RECT 242.300 185.800 242.700 186.500 ;
        RECT 243.900 185.800 244.300 186.500 ;
        RECT 245.700 185.800 246.100 186.500 ;
        RECT 248.500 186.800 249.000 187.200 ;
        RECT 240.600 185.400 241.800 185.800 ;
        RECT 242.300 185.400 243.400 185.800 ;
        RECT 243.900 185.400 245.000 185.800 ;
        RECT 245.700 185.400 246.600 185.800 ;
        RECT 236.600 184.900 237.800 185.200 ;
        RECT 236.300 184.500 236.700 184.600 ;
        RECT 235.600 184.200 236.700 184.500 ;
        RECT 237.500 184.400 237.800 184.900 ;
        RECT 237.500 184.000 238.200 184.400 ;
        RECT 234.300 183.700 234.700 183.800 ;
        RECT 235.700 183.700 236.100 183.800 ;
        RECT 232.600 183.100 233.000 183.500 ;
        RECT 234.300 183.400 236.100 183.700 ;
        RECT 235.400 183.100 235.700 183.400 ;
        RECT 237.400 183.100 237.800 183.500 ;
        RECT 232.600 182.800 233.600 183.100 ;
        RECT 233.200 181.100 233.600 182.800 ;
        RECT 235.400 181.100 235.800 183.100 ;
        RECT 237.500 181.100 238.100 183.100 ;
        RECT 239.800 181.100 240.200 185.400 ;
        RECT 241.400 181.100 241.800 185.400 ;
        RECT 243.000 181.100 243.400 185.400 ;
        RECT 244.600 181.100 245.000 185.400 ;
        RECT 246.200 181.100 246.600 185.400 ;
        RECT 248.500 185.100 248.800 186.800 ;
        RECT 249.300 186.500 249.600 187.300 ;
        RECT 249.100 186.100 249.600 186.500 ;
        RECT 249.300 185.100 249.600 186.100 ;
        RECT 250.100 186.200 250.500 186.600 ;
        RECT 250.100 185.800 250.600 186.200 ;
        RECT 248.500 184.600 249.000 185.100 ;
        RECT 249.300 184.800 250.600 185.100 ;
        RECT 248.600 181.100 249.000 184.600 ;
        RECT 250.200 181.100 250.600 184.800 ;
        RECT 0.600 175.600 1.000 179.900 ;
        RECT 2.700 177.900 3.300 179.900 ;
        RECT 5.000 177.900 5.400 179.900 ;
        RECT 7.200 178.200 7.600 179.900 ;
        RECT 7.200 177.900 8.200 178.200 ;
        RECT 3.000 177.500 3.400 177.900 ;
        RECT 5.100 177.600 5.400 177.900 ;
        RECT 4.700 177.300 6.500 177.600 ;
        RECT 7.800 177.500 8.200 177.900 ;
        RECT 4.700 177.200 5.100 177.300 ;
        RECT 6.100 177.200 6.500 177.300 ;
        RECT 2.600 176.600 3.300 177.000 ;
        RECT 3.000 176.100 3.300 176.600 ;
        RECT 4.100 176.500 5.200 176.800 ;
        RECT 4.100 176.400 4.500 176.500 ;
        RECT 3.000 175.800 4.200 176.100 ;
        RECT 0.600 175.300 2.700 175.600 ;
        RECT 0.600 173.600 1.000 175.300 ;
        RECT 2.300 175.200 2.700 175.300 ;
        RECT 1.500 174.900 1.900 175.000 ;
        RECT 1.500 174.600 3.400 174.900 ;
        RECT 3.000 174.500 3.400 174.600 ;
        RECT 3.900 174.200 4.200 175.800 ;
        RECT 4.900 175.900 5.200 176.500 ;
        RECT 5.500 176.500 5.900 176.600 ;
        RECT 7.800 176.500 8.200 176.600 ;
        RECT 5.500 176.200 8.200 176.500 ;
        RECT 4.900 175.700 7.300 175.900 ;
        RECT 9.400 175.700 9.800 179.900 ;
        RECT 10.600 176.800 11.000 177.200 ;
        RECT 10.600 176.200 10.900 176.800 ;
        RECT 11.300 176.200 11.700 179.900 ;
        RECT 10.200 175.900 10.900 176.200 ;
        RECT 11.200 175.900 11.700 176.200 ;
        RECT 10.200 175.800 10.600 175.900 ;
        RECT 4.900 175.600 9.800 175.700 ;
        RECT 6.900 175.500 9.800 175.600 ;
        RECT 7.000 175.400 9.800 175.500 ;
        RECT 11.200 175.200 11.500 175.900 ;
        RECT 13.400 175.800 13.800 176.600 ;
        RECT 6.200 175.100 6.600 175.200 ;
        RECT 6.200 174.800 8.700 175.100 ;
        RECT 11.000 174.800 11.500 175.200 ;
        RECT 7.000 174.700 7.400 174.800 ;
        RECT 8.300 174.700 8.700 174.800 ;
        RECT 7.500 174.200 7.900 174.300 ;
        RECT 11.200 174.200 11.500 174.800 ;
        RECT 11.800 175.100 12.200 175.200 ;
        RECT 13.400 175.100 13.700 175.800 ;
        RECT 11.800 174.800 13.700 175.100 ;
        RECT 11.800 174.400 12.200 174.800 ;
        RECT 3.900 173.900 9.400 174.200 ;
        RECT 4.100 173.800 4.500 173.900 ;
        RECT 0.600 173.300 2.500 173.600 ;
        RECT 0.600 171.100 1.000 173.300 ;
        RECT 2.100 173.200 2.500 173.300 ;
        RECT 7.000 172.800 7.300 173.900 ;
        RECT 8.600 173.800 9.400 173.900 ;
        RECT 10.200 173.800 11.500 174.200 ;
        RECT 12.600 174.100 13.000 174.200 ;
        RECT 12.200 173.800 13.000 174.100 ;
        RECT 13.400 174.100 13.800 174.200 ;
        RECT 14.200 174.100 14.600 179.900 ;
        RECT 13.400 173.800 14.600 174.100 ;
        RECT 6.100 172.700 6.500 172.800 ;
        RECT 3.000 172.100 3.400 172.500 ;
        RECT 5.100 172.400 6.500 172.700 ;
        RECT 7.000 172.400 7.400 172.800 ;
        RECT 5.100 172.100 5.400 172.400 ;
        RECT 7.800 172.100 8.200 172.500 ;
        RECT 2.700 171.800 3.400 172.100 ;
        RECT 2.700 171.100 3.300 171.800 ;
        RECT 5.000 171.100 5.400 172.100 ;
        RECT 7.200 171.800 8.200 172.100 ;
        RECT 7.200 171.100 7.600 171.800 ;
        RECT 9.400 171.100 9.800 173.500 ;
        RECT 10.300 173.100 10.600 173.800 ;
        RECT 12.200 173.600 12.600 173.800 ;
        RECT 11.100 173.100 12.900 173.300 ;
        RECT 14.200 173.100 14.600 173.800 ;
        RECT 15.000 173.400 15.400 174.200 ;
        RECT 15.800 173.400 16.200 174.200 ;
        RECT 10.200 171.100 10.600 173.100 ;
        RECT 11.000 173.000 13.000 173.100 ;
        RECT 11.000 171.100 11.400 173.000 ;
        RECT 12.600 171.100 13.000 173.000 ;
        RECT 13.700 172.800 14.600 173.100 ;
        RECT 16.600 173.100 17.000 179.900 ;
        RECT 17.400 175.800 17.800 176.600 ;
        RECT 19.500 176.200 19.900 179.900 ;
        RECT 20.200 176.800 20.600 177.200 ;
        RECT 20.300 176.200 20.600 176.800 ;
        RECT 19.500 175.900 20.000 176.200 ;
        RECT 20.300 175.900 21.000 176.200 ;
        RECT 19.000 174.400 19.400 175.200 ;
        RECT 19.700 174.200 20.000 175.900 ;
        RECT 20.600 175.800 21.000 175.900 ;
        RECT 21.400 175.800 21.800 176.600 ;
        RECT 20.600 175.100 20.900 175.800 ;
        RECT 22.200 175.100 22.600 179.900 ;
        RECT 23.800 175.700 24.200 179.900 ;
        RECT 26.000 178.200 26.400 179.900 ;
        RECT 25.400 177.900 26.400 178.200 ;
        RECT 28.200 177.900 28.600 179.900 ;
        RECT 30.300 177.900 30.900 179.900 ;
        RECT 25.400 177.500 25.800 177.900 ;
        RECT 28.200 177.600 28.500 177.900 ;
        RECT 27.100 177.300 28.900 177.600 ;
        RECT 30.200 177.500 30.600 177.900 ;
        RECT 27.100 177.200 27.500 177.300 ;
        RECT 28.500 177.200 28.900 177.300 ;
        RECT 25.400 176.500 25.800 176.600 ;
        RECT 27.700 176.500 28.100 176.600 ;
        RECT 25.400 176.200 28.100 176.500 ;
        RECT 28.400 176.500 29.500 176.800 ;
        RECT 28.400 175.900 28.700 176.500 ;
        RECT 29.100 176.400 29.500 176.500 ;
        RECT 30.300 176.600 31.000 177.000 ;
        RECT 30.300 176.100 30.600 176.600 ;
        RECT 26.300 175.700 28.700 175.900 ;
        RECT 23.800 175.600 28.700 175.700 ;
        RECT 29.400 175.800 30.600 176.100 ;
        RECT 23.800 175.500 26.700 175.600 ;
        RECT 23.800 175.400 26.600 175.500 ;
        RECT 27.000 175.100 27.400 175.200 ;
        RECT 20.600 174.800 22.600 175.100 ;
        RECT 18.200 174.100 18.600 174.200 ;
        RECT 19.700 174.100 21.000 174.200 ;
        RECT 21.400 174.100 21.800 174.200 ;
        RECT 18.200 173.800 19.000 174.100 ;
        RECT 19.700 173.800 21.800 174.100 ;
        RECT 18.600 173.600 19.000 173.800 ;
        RECT 18.300 173.100 20.100 173.300 ;
        RECT 20.600 173.100 20.900 173.800 ;
        RECT 22.200 173.100 22.600 174.800 ;
        RECT 24.900 174.800 27.400 175.100 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 29.400 175.100 29.700 175.800 ;
        RECT 32.600 175.600 33.000 179.900 ;
        RECT 30.900 175.300 33.000 175.600 ;
        RECT 30.900 175.200 31.300 175.300 ;
        RECT 28.600 174.800 29.700 175.100 ;
        RECT 31.700 174.900 32.100 175.000 ;
        RECT 24.900 174.700 25.300 174.800 ;
        RECT 26.200 174.700 26.600 174.800 ;
        RECT 25.700 174.200 26.100 174.300 ;
        RECT 29.400 174.200 29.700 174.800 ;
        RECT 30.200 174.600 32.100 174.900 ;
        RECT 30.200 174.500 30.600 174.600 ;
        RECT 23.000 173.400 23.400 174.200 ;
        RECT 24.200 173.900 29.700 174.200 ;
        RECT 24.200 173.800 25.000 173.900 ;
        RECT 16.600 172.800 17.500 173.100 ;
        RECT 13.700 171.100 14.100 172.800 ;
        RECT 17.100 172.200 17.500 172.800 ;
        RECT 18.200 173.000 20.200 173.100 ;
        RECT 17.100 171.800 17.800 172.200 ;
        RECT 17.100 171.100 17.500 171.800 ;
        RECT 18.200 171.100 18.600 173.000 ;
        RECT 19.800 171.100 20.200 173.000 ;
        RECT 20.600 171.100 21.000 173.100 ;
        RECT 21.700 172.800 22.600 173.100 ;
        RECT 21.700 171.100 22.100 172.800 ;
        RECT 23.800 171.100 24.200 173.500 ;
        RECT 26.300 172.800 26.600 173.900 ;
        RECT 29.100 173.800 29.500 173.900 ;
        RECT 32.600 173.600 33.000 175.300 ;
        RECT 31.100 173.300 33.000 173.600 ;
        RECT 31.100 173.200 31.500 173.300 ;
        RECT 25.400 172.100 25.800 172.500 ;
        RECT 26.200 172.400 26.600 172.800 ;
        RECT 27.100 172.700 27.500 172.800 ;
        RECT 27.100 172.400 28.500 172.700 ;
        RECT 28.200 172.100 28.500 172.400 ;
        RECT 30.200 172.100 30.600 172.500 ;
        RECT 25.400 171.800 26.400 172.100 ;
        RECT 26.000 171.100 26.400 171.800 ;
        RECT 28.200 171.100 28.600 172.100 ;
        RECT 30.200 171.800 30.900 172.100 ;
        RECT 30.300 171.100 30.900 171.800 ;
        RECT 32.600 171.100 33.000 173.300 ;
        RECT 33.400 175.600 33.800 179.900 ;
        RECT 35.500 177.900 36.100 179.900 ;
        RECT 37.800 177.900 38.200 179.900 ;
        RECT 40.000 178.200 40.400 179.900 ;
        RECT 40.000 177.900 41.000 178.200 ;
        RECT 35.800 177.500 36.200 177.900 ;
        RECT 37.900 177.600 38.200 177.900 ;
        RECT 37.500 177.300 39.300 177.600 ;
        RECT 40.600 177.500 41.000 177.900 ;
        RECT 37.500 177.200 37.900 177.300 ;
        RECT 38.900 177.200 39.300 177.300 ;
        RECT 35.400 176.600 36.100 177.000 ;
        RECT 35.800 176.100 36.100 176.600 ;
        RECT 36.900 176.500 38.000 176.800 ;
        RECT 36.900 176.400 37.300 176.500 ;
        RECT 35.800 175.800 37.000 176.100 ;
        RECT 33.400 175.300 35.500 175.600 ;
        RECT 33.400 173.600 33.800 175.300 ;
        RECT 35.100 175.200 35.500 175.300 ;
        RECT 36.700 175.200 37.000 175.800 ;
        RECT 37.700 175.900 38.000 176.500 ;
        RECT 38.300 176.500 38.700 176.600 ;
        RECT 40.600 176.500 41.000 176.600 ;
        RECT 38.300 176.200 41.000 176.500 ;
        RECT 37.700 175.700 40.100 175.900 ;
        RECT 42.200 175.700 42.600 179.900 ;
        RECT 43.400 176.800 43.800 177.200 ;
        RECT 43.400 176.200 43.700 176.800 ;
        RECT 44.100 176.200 44.500 179.900 ;
        RECT 43.000 175.900 43.700 176.200 ;
        RECT 44.000 175.900 44.500 176.200 ;
        RECT 47.800 177.500 48.200 179.500 ;
        RECT 43.000 175.800 43.400 175.900 ;
        RECT 37.700 175.600 42.600 175.700 ;
        RECT 39.700 175.500 42.600 175.600 ;
        RECT 39.800 175.400 42.600 175.500 ;
        RECT 44.000 175.200 44.300 175.900 ;
        RECT 47.800 175.800 48.100 177.500 ;
        RECT 49.900 176.400 50.300 179.900 ;
        RECT 49.900 176.100 50.700 176.400 ;
        RECT 47.800 175.500 49.700 175.800 ;
        RECT 34.300 174.900 34.700 175.000 ;
        RECT 34.300 174.600 36.200 174.900 ;
        RECT 36.600 174.800 37.000 175.200 ;
        RECT 39.000 175.100 39.400 175.200 ;
        RECT 39.000 174.800 41.500 175.100 ;
        RECT 43.800 174.800 44.300 175.200 ;
        RECT 35.800 174.500 36.200 174.600 ;
        RECT 36.700 174.200 37.000 174.800 ;
        RECT 39.800 174.700 40.200 174.800 ;
        RECT 41.100 174.700 41.500 174.800 ;
        RECT 40.300 174.200 40.700 174.300 ;
        RECT 44.000 174.200 44.300 174.800 ;
        RECT 44.600 174.400 45.000 175.200 ;
        RECT 47.800 174.400 48.200 175.200 ;
        RECT 48.600 174.400 49.000 175.200 ;
        RECT 49.400 174.500 49.700 175.500 ;
        RECT 36.700 173.900 42.200 174.200 ;
        RECT 36.900 173.800 37.300 173.900 ;
        RECT 33.400 173.300 35.300 173.600 ;
        RECT 33.400 171.100 33.800 173.300 ;
        RECT 34.900 173.200 35.300 173.300 ;
        RECT 39.800 172.800 40.100 173.900 ;
        RECT 41.400 173.800 42.200 173.900 ;
        RECT 43.000 173.800 44.300 174.200 ;
        RECT 45.400 174.100 45.800 174.200 ;
        RECT 45.000 173.800 45.800 174.100 ;
        RECT 49.400 174.100 50.100 174.500 ;
        RECT 50.400 174.200 50.700 176.100 ;
        RECT 52.600 175.800 53.000 176.600 ;
        RECT 51.000 175.100 51.400 175.600 ;
        RECT 51.800 175.100 52.200 175.200 ;
        RECT 51.000 174.800 52.200 175.100 ;
        RECT 50.400 174.100 51.400 174.200 ;
        RECT 52.600 174.100 53.000 174.200 ;
        RECT 49.400 173.900 49.900 174.100 ;
        RECT 38.900 172.700 39.300 172.800 ;
        RECT 35.800 172.100 36.200 172.500 ;
        RECT 37.900 172.400 39.300 172.700 ;
        RECT 39.800 172.400 40.200 172.800 ;
        RECT 37.900 172.100 38.200 172.400 ;
        RECT 40.600 172.100 41.000 172.500 ;
        RECT 35.500 171.800 36.200 172.100 ;
        RECT 35.500 171.100 36.100 171.800 ;
        RECT 37.800 171.100 38.200 172.100 ;
        RECT 40.000 171.800 41.000 172.100 ;
        RECT 40.000 171.100 40.400 171.800 ;
        RECT 42.200 171.100 42.600 173.500 ;
        RECT 43.100 173.100 43.400 173.800 ;
        RECT 45.000 173.600 45.400 173.800 ;
        RECT 47.800 173.600 49.900 173.900 ;
        RECT 50.400 173.800 53.000 174.100 ;
        RECT 43.900 173.100 45.700 173.300 ;
        RECT 43.000 171.100 43.400 173.100 ;
        RECT 43.800 173.000 45.800 173.100 ;
        RECT 43.800 171.100 44.200 173.000 ;
        RECT 45.400 171.100 45.800 173.000 ;
        RECT 47.800 172.500 48.100 173.600 ;
        RECT 50.400 173.500 50.700 173.800 ;
        RECT 50.300 173.300 50.700 173.500 ;
        RECT 49.900 173.000 50.700 173.300 ;
        RECT 53.400 173.100 53.800 179.900 ;
        RECT 55.000 176.200 55.400 179.900 ;
        RECT 56.600 179.600 58.600 179.900 ;
        RECT 56.600 176.200 57.000 179.600 ;
        RECT 55.000 175.900 57.000 176.200 ;
        RECT 57.400 175.900 57.800 179.300 ;
        RECT 58.200 175.900 58.600 179.600 ;
        RECT 57.400 175.600 57.700 175.900 ;
        RECT 55.400 175.200 55.800 175.400 ;
        RECT 56.700 175.300 57.700 175.600 ;
        RECT 56.700 175.200 57.000 175.300 ;
        RECT 55.000 174.900 55.800 175.200 ;
        RECT 55.000 174.800 55.400 174.900 ;
        RECT 56.600 174.800 57.000 175.200 ;
        RECT 58.200 174.800 58.600 175.600 ;
        RECT 59.800 175.100 60.200 179.900 ;
        RECT 61.800 176.800 62.200 177.200 ;
        RECT 60.600 175.800 61.000 176.600 ;
        RECT 61.800 176.200 62.100 176.800 ;
        RECT 62.500 176.200 62.900 179.900 ;
        RECT 61.400 175.900 62.100 176.200 ;
        RECT 61.400 175.800 61.800 175.900 ;
        RECT 62.400 175.800 63.400 176.200 ;
        RECT 61.400 175.100 61.700 175.800 ;
        RECT 59.800 174.800 61.700 175.100 ;
        RECT 54.200 173.400 54.600 174.200 ;
        RECT 55.000 174.100 55.400 174.200 ;
        RECT 55.800 174.100 56.200 174.600 ;
        RECT 56.700 174.200 57.000 174.800 ;
        RECT 57.300 174.400 57.700 174.800 ;
        RECT 55.000 173.800 56.200 174.100 ;
        RECT 56.600 173.800 57.000 174.200 ;
        RECT 57.400 174.200 57.700 174.400 ;
        RECT 57.400 173.800 57.800 174.200 ;
        RECT 56.700 173.100 57.000 173.800 ;
        RECT 59.000 173.400 59.400 174.200 ;
        RECT 59.800 173.100 60.200 174.800 ;
        RECT 62.400 174.200 62.700 175.800 ;
        RECT 64.600 175.600 65.000 179.900 ;
        RECT 66.700 177.900 67.300 179.900 ;
        RECT 69.000 177.900 69.400 179.900 ;
        RECT 71.200 178.200 71.600 179.900 ;
        RECT 71.200 177.900 72.200 178.200 ;
        RECT 67.000 177.500 67.400 177.900 ;
        RECT 69.100 177.600 69.400 177.900 ;
        RECT 68.700 177.300 70.500 177.600 ;
        RECT 71.800 177.500 72.200 177.900 ;
        RECT 68.700 177.200 69.100 177.300 ;
        RECT 70.100 177.200 70.500 177.300 ;
        RECT 66.600 176.600 67.300 177.000 ;
        RECT 67.000 176.100 67.300 176.600 ;
        RECT 68.100 176.500 69.200 176.800 ;
        RECT 68.100 176.400 68.500 176.500 ;
        RECT 67.000 175.800 68.200 176.100 ;
        RECT 64.600 175.300 66.700 175.600 ;
        RECT 63.000 174.400 63.400 175.200 ;
        RECT 61.400 173.800 62.700 174.200 ;
        RECT 63.800 174.100 64.200 174.200 ;
        RECT 63.400 173.800 64.200 174.100 ;
        RECT 61.500 173.100 61.800 173.800 ;
        RECT 63.400 173.600 63.800 173.800 ;
        RECT 64.600 173.600 65.000 175.300 ;
        RECT 66.300 175.200 66.700 175.300 ;
        RECT 65.500 174.900 65.900 175.000 ;
        RECT 65.500 174.600 67.400 174.900 ;
        RECT 67.000 174.500 67.400 174.600 ;
        RECT 67.900 174.200 68.200 175.800 ;
        RECT 68.900 175.900 69.200 176.500 ;
        RECT 69.500 176.500 69.900 176.600 ;
        RECT 71.800 176.500 72.200 176.600 ;
        RECT 69.500 176.200 72.200 176.500 ;
        RECT 68.900 175.700 71.300 175.900 ;
        RECT 73.400 175.700 73.800 179.900 ;
        RECT 76.100 176.400 76.500 179.900 ;
        RECT 78.200 177.500 78.600 179.500 ;
        RECT 68.900 175.600 73.800 175.700 ;
        RECT 75.700 176.100 76.500 176.400 ;
        RECT 70.900 175.500 73.800 175.600 ;
        RECT 71.000 175.400 73.800 175.500 ;
        RECT 70.200 175.100 70.600 175.200 ;
        RECT 74.200 175.100 74.600 175.200 ;
        RECT 75.000 175.100 75.400 175.600 ;
        RECT 70.200 174.800 72.700 175.100 ;
        RECT 74.200 174.800 75.400 175.100 ;
        RECT 72.300 174.700 72.700 174.800 ;
        RECT 71.500 174.200 71.900 174.300 ;
        RECT 75.700 174.200 76.000 176.100 ;
        RECT 78.300 175.800 78.600 177.500 ;
        RECT 76.700 175.500 78.600 175.800 ;
        RECT 79.000 175.700 79.400 179.900 ;
        RECT 81.200 178.200 81.600 179.900 ;
        RECT 80.600 177.900 81.600 178.200 ;
        RECT 83.400 177.900 83.800 179.900 ;
        RECT 85.500 177.900 86.100 179.900 ;
        RECT 80.600 177.500 81.000 177.900 ;
        RECT 83.400 177.600 83.700 177.900 ;
        RECT 82.300 177.300 84.100 177.600 ;
        RECT 85.400 177.500 85.800 177.900 ;
        RECT 82.300 177.200 82.700 177.300 ;
        RECT 83.700 177.200 84.100 177.300 ;
        RECT 80.600 176.500 81.000 176.600 ;
        RECT 82.900 176.500 83.300 176.600 ;
        RECT 80.600 176.200 83.300 176.500 ;
        RECT 83.600 176.500 84.700 176.800 ;
        RECT 83.600 175.900 83.900 176.500 ;
        RECT 84.300 176.400 84.700 176.500 ;
        RECT 85.500 176.600 86.200 177.000 ;
        RECT 85.500 176.100 85.800 176.600 ;
        RECT 81.500 175.700 83.900 175.900 ;
        RECT 79.000 175.600 83.900 175.700 ;
        RECT 84.600 175.800 85.800 176.100 ;
        RECT 79.000 175.500 81.900 175.600 ;
        RECT 76.700 174.500 77.000 175.500 ;
        RECT 79.000 175.400 81.800 175.500 ;
        RECT 67.900 173.900 73.400 174.200 ;
        RECT 68.100 173.800 68.500 173.900 ;
        RECT 64.600 173.300 66.500 173.600 ;
        RECT 62.300 173.100 64.100 173.300 ;
        RECT 47.800 171.500 48.200 172.500 ;
        RECT 49.900 171.500 50.300 173.000 ;
        RECT 52.900 172.800 53.800 173.100 ;
        RECT 52.900 171.100 53.300 172.800 ;
        RECT 56.500 171.100 57.300 173.100 ;
        RECT 59.800 172.800 60.700 173.100 ;
        RECT 60.300 171.100 60.700 172.800 ;
        RECT 61.400 171.100 61.800 173.100 ;
        RECT 62.200 173.000 64.200 173.100 ;
        RECT 62.200 171.100 62.600 173.000 ;
        RECT 63.800 171.100 64.200 173.000 ;
        RECT 64.600 171.100 65.000 173.300 ;
        RECT 66.100 173.200 66.500 173.300 ;
        RECT 71.000 173.200 71.300 173.900 ;
        RECT 72.600 173.800 73.400 173.900 ;
        RECT 75.000 173.800 76.000 174.200 ;
        RECT 76.300 174.100 77.000 174.500 ;
        RECT 77.400 174.400 77.800 175.200 ;
        RECT 78.200 174.400 78.600 175.200 ;
        RECT 82.200 175.100 82.600 175.200 ;
        RECT 80.100 174.800 82.600 175.100 ;
        RECT 80.100 174.700 80.500 174.800 ;
        RECT 81.400 174.700 81.800 174.800 ;
        RECT 80.900 174.200 81.300 174.300 ;
        RECT 84.600 174.200 84.900 175.800 ;
        RECT 87.800 175.600 88.200 179.900 ;
        RECT 90.500 176.400 90.900 179.900 ;
        RECT 92.600 177.500 93.000 179.500 ;
        RECT 90.100 176.100 90.900 176.400 ;
        RECT 86.100 175.300 88.200 175.600 ;
        RECT 86.100 175.200 86.500 175.300 ;
        RECT 87.800 175.100 88.200 175.300 ;
        RECT 89.400 175.100 89.800 175.600 ;
        RECT 86.900 174.900 87.300 175.000 ;
        RECT 85.400 174.600 87.300 174.900 ;
        RECT 87.800 174.800 89.800 175.100 ;
        RECT 85.400 174.500 85.800 174.600 ;
        RECT 75.700 173.500 76.000 173.800 ;
        RECT 76.500 173.900 77.000 174.100 ;
        RECT 79.400 173.900 84.900 174.200 ;
        RECT 76.500 173.600 78.600 173.900 ;
        RECT 79.400 173.800 80.200 173.900 ;
        RECT 70.100 172.700 70.500 172.800 ;
        RECT 67.000 172.100 67.400 172.500 ;
        RECT 69.100 172.400 70.500 172.700 ;
        RECT 71.000 172.400 71.400 173.200 ;
        RECT 69.100 172.100 69.400 172.400 ;
        RECT 71.800 172.100 72.200 172.500 ;
        RECT 66.700 171.800 67.400 172.100 ;
        RECT 66.700 171.100 67.300 171.800 ;
        RECT 69.000 171.100 69.400 172.100 ;
        RECT 71.200 171.800 72.200 172.100 ;
        RECT 71.200 171.100 71.600 171.800 ;
        RECT 73.400 171.100 73.800 173.500 ;
        RECT 75.700 173.300 76.100 173.500 ;
        RECT 75.700 173.000 76.500 173.300 ;
        RECT 76.100 171.500 76.500 173.000 ;
        RECT 78.300 172.500 78.600 173.600 ;
        RECT 78.200 171.500 78.600 172.500 ;
        RECT 79.000 171.100 79.400 173.500 ;
        RECT 81.500 172.800 81.800 173.900 ;
        RECT 84.300 173.800 84.700 173.900 ;
        RECT 87.800 173.600 88.200 174.800 ;
        RECT 90.100 174.200 90.400 176.100 ;
        RECT 92.700 175.800 93.000 177.500 ;
        RECT 95.300 176.400 95.700 179.900 ;
        RECT 97.400 177.500 97.800 179.500 ;
        RECT 91.100 175.500 93.000 175.800 ;
        RECT 94.900 176.100 95.700 176.400 ;
        RECT 91.100 174.500 91.400 175.500 ;
        RECT 88.600 174.100 89.000 174.200 ;
        RECT 89.400 174.100 90.400 174.200 ;
        RECT 90.700 174.100 91.400 174.500 ;
        RECT 91.800 174.400 92.200 175.200 ;
        RECT 92.600 174.400 93.000 175.200 ;
        RECT 94.200 174.800 94.600 175.600 ;
        RECT 94.900 174.200 95.200 176.100 ;
        RECT 97.500 175.800 97.800 177.500 ;
        RECT 101.700 176.400 102.100 179.900 ;
        RECT 103.800 177.500 104.200 179.500 ;
        RECT 95.900 175.500 97.800 175.800 ;
        RECT 101.300 176.100 102.100 176.400 ;
        RECT 95.900 174.500 96.200 175.500 ;
        RECT 88.600 173.800 90.400 174.100 ;
        RECT 86.300 173.300 88.200 173.600 ;
        RECT 86.300 173.200 86.700 173.300 ;
        RECT 80.600 172.100 81.000 172.500 ;
        RECT 81.400 172.400 81.800 172.800 ;
        RECT 82.300 172.700 82.700 172.800 ;
        RECT 82.300 172.400 83.700 172.700 ;
        RECT 83.400 172.100 83.700 172.400 ;
        RECT 85.400 172.100 85.800 172.500 ;
        RECT 80.600 171.800 81.600 172.100 ;
        RECT 81.200 171.100 81.600 171.800 ;
        RECT 83.400 171.100 83.800 172.100 ;
        RECT 85.400 171.800 86.100 172.100 ;
        RECT 85.500 171.100 86.100 171.800 ;
        RECT 87.800 171.100 88.200 173.300 ;
        RECT 90.100 173.500 90.400 173.800 ;
        RECT 90.900 173.900 91.400 174.100 ;
        RECT 90.900 173.600 93.000 173.900 ;
        RECT 94.200 173.800 95.200 174.200 ;
        RECT 95.500 174.100 96.200 174.500 ;
        RECT 96.600 174.400 97.000 175.200 ;
        RECT 97.400 174.400 97.800 175.200 ;
        RECT 100.600 174.800 101.000 175.600 ;
        RECT 101.300 174.200 101.600 176.100 ;
        RECT 103.900 175.800 104.200 177.500 ;
        RECT 102.300 175.500 104.200 175.800 ;
        RECT 104.600 175.600 105.000 179.900 ;
        RECT 106.700 177.900 107.300 179.900 ;
        RECT 109.000 177.900 109.400 179.900 ;
        RECT 111.200 178.200 111.600 179.900 ;
        RECT 111.200 177.900 112.200 178.200 ;
        RECT 107.000 177.500 107.400 177.900 ;
        RECT 109.100 177.600 109.400 177.900 ;
        RECT 108.700 177.300 110.500 177.600 ;
        RECT 111.800 177.500 112.200 177.900 ;
        RECT 108.700 177.200 109.100 177.300 ;
        RECT 110.100 177.200 110.500 177.300 ;
        RECT 106.600 176.600 107.300 177.000 ;
        RECT 107.000 176.100 107.300 176.600 ;
        RECT 108.100 176.500 109.200 176.800 ;
        RECT 108.100 176.400 108.500 176.500 ;
        RECT 107.000 175.800 108.200 176.100 ;
        RECT 102.300 174.500 102.600 175.500 ;
        RECT 104.600 175.300 106.700 175.600 ;
        RECT 90.100 173.300 90.500 173.500 ;
        RECT 90.100 173.000 90.900 173.300 ;
        RECT 90.500 171.500 90.900 173.000 ;
        RECT 92.700 172.500 93.000 173.600 ;
        RECT 94.900 173.500 95.200 173.800 ;
        RECT 95.700 173.900 96.200 174.100 ;
        RECT 98.200 174.100 98.600 174.200 ;
        RECT 100.600 174.100 101.600 174.200 ;
        RECT 101.900 174.100 102.600 174.500 ;
        RECT 103.000 174.400 103.400 175.200 ;
        RECT 103.800 174.400 104.200 175.200 ;
        RECT 95.700 173.600 97.800 173.900 ;
        RECT 98.200 173.800 101.600 174.100 ;
        RECT 94.900 173.300 95.300 173.500 ;
        RECT 94.900 173.000 95.700 173.300 ;
        RECT 92.600 171.500 93.000 172.500 ;
        RECT 95.300 172.200 95.700 173.000 ;
        RECT 97.500 172.500 97.800 173.600 ;
        RECT 101.300 173.500 101.600 173.800 ;
        RECT 102.100 173.900 102.600 174.100 ;
        RECT 102.100 173.600 104.200 173.900 ;
        RECT 101.300 173.300 101.700 173.500 ;
        RECT 101.300 173.000 102.100 173.300 ;
        RECT 95.000 171.800 95.700 172.200 ;
        RECT 95.300 171.500 95.700 171.800 ;
        RECT 97.400 171.500 97.800 172.500 ;
        RECT 101.700 171.500 102.100 173.000 ;
        RECT 103.900 172.500 104.200 173.600 ;
        RECT 103.800 171.500 104.200 172.500 ;
        RECT 104.600 173.600 105.000 175.300 ;
        RECT 106.300 175.200 106.700 175.300 ;
        RECT 105.500 174.900 105.900 175.000 ;
        RECT 105.500 174.600 107.400 174.900 ;
        RECT 107.000 174.500 107.400 174.600 ;
        RECT 107.900 174.200 108.200 175.800 ;
        RECT 108.900 175.900 109.200 176.500 ;
        RECT 109.500 176.500 109.900 176.600 ;
        RECT 111.800 176.500 112.200 176.600 ;
        RECT 109.500 176.200 112.200 176.500 ;
        RECT 108.900 175.700 111.300 175.900 ;
        RECT 113.400 175.700 113.800 179.900 ;
        RECT 108.900 175.600 113.800 175.700 ;
        RECT 110.900 175.500 113.800 175.600 ;
        RECT 111.000 175.400 113.800 175.500 ;
        RECT 110.200 175.100 110.600 175.200 ;
        RECT 115.000 175.100 115.400 179.900 ;
        RECT 117.000 176.800 117.400 177.200 ;
        RECT 115.800 175.800 116.200 176.600 ;
        RECT 117.000 176.200 117.300 176.800 ;
        RECT 117.700 176.200 118.100 179.900 ;
        RECT 116.600 175.900 117.300 176.200 ;
        RECT 117.600 175.900 118.100 176.200 ;
        RECT 116.600 175.800 117.000 175.900 ;
        RECT 116.600 175.100 116.900 175.800 ;
        RECT 110.200 174.800 112.700 175.100 ;
        RECT 111.000 174.700 111.400 174.800 ;
        RECT 112.300 174.700 112.700 174.800 ;
        RECT 115.000 174.800 116.900 175.100 ;
        RECT 111.500 174.200 111.900 174.300 ;
        RECT 107.900 173.900 113.400 174.200 ;
        RECT 108.100 173.800 109.000 173.900 ;
        RECT 104.600 173.300 106.500 173.600 ;
        RECT 104.600 171.100 105.000 173.300 ;
        RECT 106.100 173.200 106.500 173.300 ;
        RECT 111.000 172.800 111.300 173.900 ;
        RECT 112.600 173.800 113.400 173.900 ;
        RECT 110.100 172.700 110.500 172.800 ;
        RECT 107.000 172.100 107.400 172.500 ;
        RECT 109.100 172.400 110.500 172.700 ;
        RECT 111.000 172.400 111.400 172.800 ;
        RECT 109.100 172.100 109.400 172.400 ;
        RECT 111.800 172.100 112.200 172.500 ;
        RECT 106.700 171.800 107.400 172.100 ;
        RECT 106.700 171.100 107.300 171.800 ;
        RECT 109.000 171.100 109.400 172.100 ;
        RECT 111.200 171.800 112.200 172.100 ;
        RECT 111.200 171.100 111.600 171.800 ;
        RECT 113.400 171.100 113.800 173.500 ;
        RECT 114.200 173.400 114.600 174.200 ;
        RECT 115.000 173.100 115.400 174.800 ;
        RECT 117.600 174.200 117.900 175.900 ;
        RECT 119.800 175.800 120.200 176.600 ;
        RECT 118.200 174.400 118.600 175.200 ;
        RECT 115.800 174.100 116.200 174.200 ;
        RECT 116.600 174.100 117.900 174.200 ;
        RECT 119.000 174.100 119.400 174.200 ;
        RECT 115.800 173.800 117.900 174.100 ;
        RECT 118.600 173.800 119.400 174.100 ;
        RECT 116.700 173.100 117.000 173.800 ;
        RECT 118.600 173.600 119.000 173.800 ;
        RECT 117.500 173.100 119.300 173.300 ;
        RECT 120.600 173.100 121.000 179.900 ;
        RECT 123.000 176.400 123.400 179.900 ;
        RECT 122.900 175.900 123.400 176.400 ;
        RECT 124.600 176.200 125.000 179.900 ;
        RECT 127.300 176.400 127.700 179.900 ;
        RECT 129.400 177.500 129.800 179.500 ;
        RECT 123.700 175.900 125.000 176.200 ;
        RECT 126.900 176.100 127.700 176.400 ;
        RECT 122.900 174.200 123.200 175.900 ;
        RECT 123.700 174.900 124.000 175.900 ;
        RECT 123.500 174.500 124.000 174.900 ;
        RECT 121.400 173.400 121.800 174.200 ;
        RECT 122.900 173.800 123.400 174.200 ;
        RECT 115.000 172.800 115.900 173.100 ;
        RECT 115.500 171.100 115.900 172.800 ;
        RECT 116.600 171.100 117.000 173.100 ;
        RECT 117.400 173.000 119.400 173.100 ;
        RECT 117.400 171.100 117.800 173.000 ;
        RECT 119.000 171.100 119.400 173.000 ;
        RECT 120.100 172.800 121.000 173.100 ;
        RECT 122.900 173.100 123.200 173.800 ;
        RECT 123.700 173.700 124.000 174.500 ;
        RECT 124.500 175.100 125.000 175.200 ;
        RECT 125.400 175.100 125.800 175.200 ;
        RECT 124.500 174.800 125.800 175.100 ;
        RECT 126.200 174.800 126.600 175.600 ;
        RECT 124.500 174.400 124.900 174.800 ;
        RECT 126.900 174.200 127.200 176.100 ;
        RECT 129.500 175.800 129.800 177.500 ;
        RECT 130.200 176.200 130.600 179.900 ;
        RECT 131.800 179.600 133.800 179.900 ;
        RECT 131.800 176.200 132.200 179.600 ;
        RECT 130.200 175.900 132.200 176.200 ;
        RECT 132.600 175.900 133.000 179.300 ;
        RECT 133.400 175.900 133.800 179.600 ;
        RECT 136.100 176.400 136.500 179.900 ;
        RECT 138.200 177.500 138.600 179.500 ;
        RECT 135.700 176.100 136.500 176.400 ;
        RECT 127.900 175.500 129.800 175.800 ;
        RECT 132.600 175.600 132.900 175.900 ;
        RECT 127.900 174.500 128.200 175.500 ;
        RECT 130.600 175.200 131.000 175.400 ;
        RECT 131.900 175.300 132.900 175.600 ;
        RECT 131.900 175.200 132.200 175.300 ;
        RECT 126.200 173.800 127.200 174.200 ;
        RECT 127.500 174.100 128.200 174.500 ;
        RECT 128.600 174.400 129.000 175.200 ;
        RECT 129.400 174.400 129.800 175.200 ;
        RECT 130.200 174.900 131.000 175.200 ;
        RECT 130.200 174.800 130.600 174.900 ;
        RECT 131.800 174.800 132.200 175.200 ;
        RECT 133.400 174.800 133.800 175.600 ;
        RECT 135.000 174.800 135.400 175.600 ;
        RECT 123.700 173.400 125.000 173.700 ;
        RECT 122.900 172.800 123.400 173.100 ;
        RECT 120.100 171.100 120.500 172.800 ;
        RECT 123.000 171.100 123.400 172.800 ;
        RECT 124.600 171.100 125.000 173.400 ;
        RECT 126.900 173.500 127.200 173.800 ;
        RECT 127.700 173.900 128.200 174.100 ;
        RECT 127.700 173.600 129.800 173.900 ;
        RECT 131.000 173.800 131.400 174.600 ;
        RECT 126.900 173.300 127.300 173.500 ;
        RECT 126.900 173.200 127.700 173.300 ;
        RECT 126.900 173.000 128.200 173.200 ;
        RECT 127.300 172.800 128.200 173.000 ;
        RECT 127.300 171.500 127.700 172.800 ;
        RECT 129.500 172.500 129.800 173.600 ;
        RECT 131.900 173.100 132.200 174.800 ;
        RECT 132.500 174.400 132.900 174.800 ;
        RECT 132.600 174.200 132.900 174.400 ;
        RECT 135.700 174.200 136.000 176.100 ;
        RECT 138.300 175.800 138.600 177.500 ;
        RECT 140.900 179.200 141.300 179.900 ;
        RECT 140.900 178.800 141.800 179.200 ;
        RECT 140.900 176.400 141.300 178.800 ;
        RECT 143.000 177.500 143.400 179.500 ;
        RECT 136.700 175.500 138.600 175.800 ;
        RECT 140.500 176.100 141.300 176.400 ;
        RECT 136.700 174.500 137.000 175.500 ;
        RECT 132.600 174.100 133.000 174.200 ;
        RECT 135.000 174.100 136.000 174.200 ;
        RECT 136.300 174.100 137.000 174.500 ;
        RECT 137.400 174.400 137.800 175.200 ;
        RECT 138.200 174.400 138.600 175.200 ;
        RECT 139.800 174.800 140.200 175.600 ;
        RECT 140.500 174.200 140.800 176.100 ;
        RECT 143.100 175.800 143.400 177.500 ;
        RECT 145.700 176.400 146.100 179.900 ;
        RECT 147.800 177.500 148.200 179.500 ;
        RECT 141.500 175.500 143.400 175.800 ;
        RECT 145.300 176.100 146.100 176.400 ;
        RECT 141.500 174.500 141.800 175.500 ;
        RECT 132.600 173.800 136.000 174.100 ;
        RECT 135.700 173.500 136.000 173.800 ;
        RECT 136.500 173.900 137.000 174.100 ;
        RECT 136.500 173.600 138.600 173.900 ;
        RECT 139.800 173.800 140.800 174.200 ;
        RECT 141.100 174.100 141.800 174.500 ;
        RECT 142.200 174.400 142.600 175.200 ;
        RECT 143.000 174.400 143.400 175.200 ;
        RECT 143.800 174.800 144.200 175.200 ;
        RECT 144.600 174.800 145.000 175.600 ;
        RECT 135.700 173.300 136.100 173.500 ;
        RECT 129.400 171.500 129.800 172.500 ;
        RECT 131.700 171.100 132.500 173.100 ;
        RECT 135.700 173.000 136.500 173.300 ;
        RECT 136.100 171.500 136.500 173.000 ;
        RECT 138.300 172.500 138.600 173.600 ;
        RECT 140.500 173.500 140.800 173.800 ;
        RECT 141.300 173.900 141.800 174.100 ;
        RECT 143.800 174.100 144.100 174.800 ;
        RECT 145.300 174.200 145.600 176.100 ;
        RECT 147.900 175.800 148.200 177.500 ;
        RECT 146.300 175.500 148.200 175.800 ;
        RECT 146.300 174.500 146.600 175.500 ;
        RECT 144.600 174.100 145.600 174.200 ;
        RECT 145.900 174.100 146.600 174.500 ;
        RECT 147.000 174.400 147.400 175.200 ;
        RECT 147.800 174.400 148.200 175.200 ;
        RECT 149.400 175.100 149.800 179.900 ;
        RECT 153.000 176.800 153.400 177.200 ;
        RECT 150.200 175.800 150.600 176.600 ;
        RECT 153.000 176.200 153.300 176.800 ;
        RECT 153.700 176.200 154.100 179.900 ;
        RECT 152.600 175.900 153.300 176.200 ;
        RECT 152.600 175.800 153.000 175.900 ;
        RECT 153.600 175.800 154.600 176.200 ;
        RECT 152.600 175.100 152.900 175.800 ;
        RECT 149.400 174.800 152.900 175.100 ;
        RECT 141.300 173.600 143.400 173.900 ;
        RECT 143.800 173.800 145.600 174.100 ;
        RECT 140.500 173.300 140.900 173.500 ;
        RECT 140.500 173.000 141.300 173.300 ;
        RECT 138.200 171.500 138.600 172.500 ;
        RECT 140.900 171.500 141.300 173.000 ;
        RECT 143.100 172.500 143.400 173.600 ;
        RECT 145.300 173.500 145.600 173.800 ;
        RECT 146.100 173.900 146.600 174.100 ;
        RECT 146.100 173.600 148.200 173.900 ;
        RECT 145.300 173.300 145.700 173.500 ;
        RECT 145.300 173.000 146.100 173.300 ;
        RECT 143.000 171.500 143.400 172.500 ;
        RECT 145.700 171.500 146.100 173.000 ;
        RECT 147.900 172.500 148.200 173.600 ;
        RECT 148.600 173.400 149.000 174.200 ;
        RECT 149.400 173.100 149.800 174.800 ;
        RECT 153.600 174.200 153.900 175.800 ;
        RECT 155.800 175.600 156.200 179.900 ;
        RECT 157.900 177.900 158.500 179.900 ;
        RECT 160.200 177.900 160.600 179.900 ;
        RECT 162.400 178.200 162.800 179.900 ;
        RECT 162.400 177.900 163.400 178.200 ;
        RECT 158.200 177.500 158.600 177.900 ;
        RECT 160.300 177.600 160.600 177.900 ;
        RECT 159.900 177.300 161.700 177.600 ;
        RECT 163.000 177.500 163.400 177.900 ;
        RECT 159.900 177.200 160.300 177.300 ;
        RECT 161.300 177.200 161.700 177.300 ;
        RECT 157.800 176.600 158.500 177.000 ;
        RECT 158.200 176.100 158.500 176.600 ;
        RECT 159.300 176.500 160.400 176.800 ;
        RECT 159.300 176.400 159.700 176.500 ;
        RECT 158.200 175.800 159.400 176.100 ;
        RECT 155.800 175.300 157.900 175.600 ;
        RECT 154.200 174.400 154.600 175.200 ;
        RECT 152.600 173.800 153.900 174.200 ;
        RECT 155.000 174.100 155.400 174.200 ;
        RECT 154.600 173.800 155.400 174.100 ;
        RECT 152.700 173.100 153.000 173.800 ;
        RECT 154.600 173.600 155.000 173.800 ;
        RECT 155.800 173.600 156.200 175.300 ;
        RECT 157.500 175.200 157.900 175.300 ;
        RECT 159.100 175.200 159.400 175.800 ;
        RECT 160.100 175.900 160.400 176.500 ;
        RECT 160.700 176.500 161.100 176.600 ;
        RECT 163.000 176.500 163.400 176.600 ;
        RECT 160.700 176.200 163.400 176.500 ;
        RECT 160.100 175.700 162.500 175.900 ;
        RECT 164.600 175.700 165.000 179.900 ;
        RECT 167.300 176.400 167.700 179.900 ;
        RECT 169.400 177.500 169.800 179.500 ;
        RECT 160.100 175.600 165.000 175.700 ;
        RECT 166.900 176.100 167.700 176.400 ;
        RECT 162.100 175.500 165.000 175.600 ;
        RECT 162.200 175.400 165.000 175.500 ;
        RECT 156.700 174.900 157.100 175.000 ;
        RECT 156.700 174.600 158.600 174.900 ;
        RECT 159.000 174.800 159.400 175.200 ;
        RECT 161.400 175.100 161.800 175.200 ;
        RECT 161.400 174.800 163.900 175.100 ;
        RECT 166.200 174.800 166.600 175.600 ;
        RECT 158.200 174.500 158.600 174.600 ;
        RECT 159.100 174.200 159.400 174.800 ;
        RECT 163.500 174.700 163.900 174.800 ;
        RECT 162.700 174.200 163.100 174.300 ;
        RECT 166.900 174.200 167.200 176.100 ;
        RECT 169.500 175.800 169.800 177.500 ;
        RECT 167.900 175.500 169.800 175.800 ;
        RECT 167.900 174.500 168.200 175.500 ;
        RECT 159.100 173.900 164.600 174.200 ;
        RECT 159.300 173.800 159.700 173.900 ;
        RECT 155.800 173.300 157.700 173.600 ;
        RECT 153.500 173.100 155.300 173.300 ;
        RECT 149.400 172.800 150.300 173.100 ;
        RECT 147.800 171.500 148.200 172.500 ;
        RECT 149.900 171.100 150.300 172.800 ;
        RECT 152.600 171.100 153.000 173.100 ;
        RECT 153.400 173.000 155.400 173.100 ;
        RECT 153.400 171.100 153.800 173.000 ;
        RECT 155.000 171.100 155.400 173.000 ;
        RECT 155.800 171.100 156.200 173.300 ;
        RECT 157.300 173.200 157.700 173.300 ;
        RECT 162.200 172.800 162.500 173.900 ;
        RECT 163.800 173.800 164.600 173.900 ;
        RECT 165.400 174.100 165.800 174.200 ;
        RECT 166.200 174.100 167.200 174.200 ;
        RECT 167.500 174.100 168.200 174.500 ;
        RECT 168.600 174.400 169.000 175.200 ;
        RECT 169.400 174.400 169.800 175.200 ;
        RECT 171.000 175.100 171.400 179.900 ;
        RECT 173.700 177.200 174.100 179.900 ;
        RECT 173.000 176.800 173.400 177.200 ;
        RECT 173.700 176.800 174.600 177.200 ;
        RECT 171.800 175.800 172.200 176.600 ;
        RECT 173.000 176.200 173.300 176.800 ;
        RECT 173.700 176.200 174.100 176.800 ;
        RECT 172.600 175.900 173.300 176.200 ;
        RECT 173.600 175.900 174.100 176.200 ;
        RECT 172.600 175.800 173.000 175.900 ;
        RECT 172.600 175.100 172.900 175.800 ;
        RECT 171.000 174.800 172.900 175.100 ;
        RECT 165.400 173.800 167.200 174.100 ;
        RECT 166.900 173.500 167.200 173.800 ;
        RECT 167.700 173.900 168.200 174.100 ;
        RECT 167.700 173.600 169.800 173.900 ;
        RECT 161.300 172.700 161.700 172.800 ;
        RECT 158.200 172.100 158.600 172.500 ;
        RECT 160.300 172.400 161.700 172.700 ;
        RECT 162.200 172.400 162.600 172.800 ;
        RECT 160.300 172.100 160.600 172.400 ;
        RECT 163.000 172.100 163.400 172.500 ;
        RECT 157.900 171.800 158.600 172.100 ;
        RECT 157.900 171.100 158.500 171.800 ;
        RECT 160.200 171.100 160.600 172.100 ;
        RECT 162.400 171.800 163.400 172.100 ;
        RECT 162.400 171.100 162.800 171.800 ;
        RECT 164.600 171.100 165.000 173.500 ;
        RECT 166.900 173.300 167.300 173.500 ;
        RECT 166.900 173.000 167.700 173.300 ;
        RECT 167.300 171.500 167.700 173.000 ;
        RECT 169.500 172.500 169.800 173.600 ;
        RECT 170.200 173.400 170.600 174.200 ;
        RECT 171.000 173.100 171.400 174.800 ;
        RECT 173.600 174.200 173.900 175.900 ;
        RECT 175.800 175.600 176.200 179.900 ;
        RECT 177.900 177.900 178.500 179.900 ;
        RECT 180.200 177.900 180.600 179.900 ;
        RECT 182.400 178.200 182.800 179.900 ;
        RECT 182.400 177.900 183.400 178.200 ;
        RECT 178.200 177.500 178.600 177.900 ;
        RECT 180.300 177.600 180.600 177.900 ;
        RECT 179.900 177.300 181.700 177.600 ;
        RECT 183.000 177.500 183.400 177.900 ;
        RECT 179.900 177.200 180.300 177.300 ;
        RECT 181.300 177.200 181.700 177.300 ;
        RECT 177.400 177.000 178.100 177.200 ;
        RECT 177.400 176.800 178.500 177.000 ;
        RECT 177.800 176.600 178.500 176.800 ;
        RECT 178.200 176.100 178.500 176.600 ;
        RECT 179.300 176.500 180.400 176.800 ;
        RECT 179.300 176.400 179.700 176.500 ;
        RECT 178.200 175.800 179.400 176.100 ;
        RECT 175.800 175.300 177.900 175.600 ;
        RECT 174.200 174.400 174.600 175.200 ;
        RECT 172.600 173.800 173.900 174.200 ;
        RECT 175.000 174.100 175.400 174.200 ;
        RECT 174.600 173.800 175.400 174.100 ;
        RECT 172.700 173.100 173.000 173.800 ;
        RECT 174.600 173.600 175.000 173.800 ;
        RECT 175.800 173.600 176.200 175.300 ;
        RECT 177.500 175.200 177.900 175.300 ;
        RECT 176.700 174.900 177.100 175.000 ;
        RECT 176.700 174.600 178.600 174.900 ;
        RECT 178.200 174.500 178.600 174.600 ;
        RECT 179.100 174.200 179.400 175.800 ;
        RECT 180.100 175.900 180.400 176.500 ;
        RECT 180.700 176.500 181.100 176.600 ;
        RECT 183.000 176.500 183.400 176.600 ;
        RECT 180.700 176.200 183.400 176.500 ;
        RECT 180.100 175.700 182.500 175.900 ;
        RECT 184.600 175.700 185.000 179.900 ;
        RECT 185.400 176.200 185.800 179.900 ;
        RECT 187.000 176.400 187.400 179.900 ;
        RECT 185.400 175.900 186.700 176.200 ;
        RECT 187.000 175.900 187.500 176.400 ;
        RECT 180.100 175.600 185.000 175.700 ;
        RECT 182.100 175.500 185.000 175.600 ;
        RECT 182.200 175.400 185.000 175.500 ;
        RECT 180.600 175.100 181.000 175.200 ;
        RECT 181.400 175.100 181.800 175.200 ;
        RECT 180.600 174.800 183.900 175.100 ;
        RECT 185.400 174.800 185.900 175.200 ;
        RECT 183.500 174.700 183.900 174.800 ;
        RECT 185.500 174.400 185.900 174.800 ;
        RECT 186.400 174.900 186.700 175.900 ;
        RECT 186.400 174.500 186.900 174.900 ;
        RECT 182.700 174.200 183.100 174.300 ;
        RECT 179.100 173.900 184.600 174.200 ;
        RECT 179.300 173.800 179.700 173.900 ;
        RECT 175.800 173.300 177.700 173.600 ;
        RECT 173.500 173.100 175.300 173.300 ;
        RECT 171.000 172.800 171.900 173.100 ;
        RECT 169.400 171.500 169.800 172.500 ;
        RECT 171.500 171.100 171.900 172.800 ;
        RECT 172.600 171.100 173.000 173.100 ;
        RECT 173.400 173.000 175.400 173.100 ;
        RECT 173.400 171.100 173.800 173.000 ;
        RECT 175.000 171.100 175.400 173.000 ;
        RECT 175.800 171.100 176.200 173.300 ;
        RECT 177.300 173.200 177.700 173.300 ;
        RECT 182.200 172.800 182.500 173.900 ;
        RECT 183.800 173.800 184.600 173.900 ;
        RECT 186.400 173.700 186.700 174.500 ;
        RECT 187.200 174.200 187.500 175.900 ;
        RECT 188.600 175.700 189.000 179.900 ;
        RECT 190.800 178.200 191.200 179.900 ;
        RECT 190.200 177.900 191.200 178.200 ;
        RECT 193.000 177.900 193.400 179.900 ;
        RECT 195.100 177.900 195.700 179.900 ;
        RECT 190.200 177.500 190.600 177.900 ;
        RECT 193.000 177.600 193.300 177.900 ;
        RECT 191.900 177.300 193.700 177.600 ;
        RECT 195.000 177.500 195.400 177.900 ;
        RECT 191.900 177.200 192.300 177.300 ;
        RECT 193.300 177.200 193.700 177.300 ;
        RECT 190.200 176.500 190.600 176.600 ;
        RECT 192.500 176.500 192.900 176.600 ;
        RECT 190.200 176.200 192.900 176.500 ;
        RECT 193.200 176.500 194.300 176.800 ;
        RECT 193.200 175.900 193.500 176.500 ;
        RECT 193.900 176.400 194.300 176.500 ;
        RECT 195.100 176.600 195.800 177.000 ;
        RECT 195.100 176.100 195.400 176.600 ;
        RECT 191.100 175.700 193.500 175.900 ;
        RECT 188.600 175.600 193.500 175.700 ;
        RECT 194.200 175.800 195.400 176.100 ;
        RECT 188.600 175.500 191.500 175.600 ;
        RECT 188.600 175.400 191.400 175.500 ;
        RECT 191.800 175.100 192.200 175.200 ;
        RECT 192.600 175.100 193.000 175.200 ;
        RECT 189.700 174.800 193.000 175.100 ;
        RECT 189.700 174.700 190.100 174.800 ;
        RECT 190.500 174.200 190.900 174.300 ;
        RECT 194.200 174.200 194.500 175.800 ;
        RECT 197.400 175.600 197.800 179.900 ;
        RECT 195.700 175.300 197.800 175.600 ;
        RECT 198.200 177.500 198.600 179.500 ;
        RECT 200.300 179.200 200.700 179.900 ;
        RECT 199.800 178.800 200.700 179.200 ;
        RECT 198.200 175.800 198.500 177.500 ;
        RECT 200.300 176.400 200.700 178.800 ;
        RECT 204.600 179.600 206.600 179.900 ;
        RECT 200.300 176.100 201.100 176.400 ;
        RECT 198.200 175.500 200.100 175.800 ;
        RECT 195.700 175.200 196.100 175.300 ;
        RECT 196.500 174.900 196.900 175.000 ;
        RECT 195.000 174.600 196.900 174.900 ;
        RECT 195.000 174.500 195.400 174.600 ;
        RECT 187.000 173.800 187.500 174.200 ;
        RECT 189.000 173.900 194.500 174.200 ;
        RECT 189.000 173.800 189.800 173.900 ;
        RECT 181.300 172.700 181.700 172.800 ;
        RECT 178.200 172.100 178.600 172.500 ;
        RECT 180.300 172.400 181.700 172.700 ;
        RECT 182.200 172.400 182.600 172.800 ;
        RECT 180.300 172.100 180.600 172.400 ;
        RECT 183.000 172.100 183.400 172.500 ;
        RECT 177.900 171.800 178.600 172.100 ;
        RECT 177.900 171.100 178.500 171.800 ;
        RECT 180.200 171.100 180.600 172.100 ;
        RECT 182.400 171.800 183.400 172.100 ;
        RECT 182.400 171.100 182.800 171.800 ;
        RECT 184.600 171.100 185.000 173.500 ;
        RECT 185.400 173.400 186.700 173.700 ;
        RECT 185.400 171.100 185.800 173.400 ;
        RECT 187.200 173.100 187.500 173.800 ;
        RECT 187.000 172.800 187.500 173.100 ;
        RECT 187.000 171.100 187.400 172.800 ;
        RECT 188.600 171.100 189.000 173.500 ;
        RECT 191.100 172.800 191.400 173.900 ;
        RECT 191.800 173.800 192.200 173.900 ;
        RECT 193.900 173.800 194.300 173.900 ;
        RECT 197.400 173.600 197.800 175.300 ;
        RECT 198.200 174.400 198.600 175.200 ;
        RECT 199.000 174.400 199.400 175.200 ;
        RECT 199.800 174.500 200.100 175.500 ;
        RECT 199.800 174.100 200.500 174.500 ;
        RECT 200.800 174.200 201.100 176.100 ;
        RECT 204.600 175.900 205.000 179.600 ;
        RECT 205.400 175.900 205.800 179.300 ;
        RECT 206.200 176.200 206.600 179.600 ;
        RECT 207.800 176.200 208.200 179.900 ;
        RECT 206.200 175.900 208.200 176.200 ;
        RECT 209.900 176.200 210.300 179.900 ;
        RECT 210.600 176.800 211.000 177.200 ;
        RECT 210.700 176.200 211.000 176.800 ;
        RECT 209.900 175.900 210.400 176.200 ;
        RECT 210.700 175.900 211.400 176.200 ;
        RECT 205.500 175.600 205.800 175.900 ;
        RECT 201.400 174.800 201.800 175.600 ;
        RECT 204.600 174.800 205.000 175.600 ;
        RECT 205.500 175.300 206.500 175.600 ;
        RECT 206.200 175.200 206.500 175.300 ;
        RECT 207.400 175.200 207.800 175.400 ;
        RECT 210.100 175.200 210.400 175.900 ;
        RECT 211.000 175.800 211.400 175.900 ;
        RECT 211.800 175.600 212.200 179.900 ;
        RECT 213.900 177.900 214.500 179.900 ;
        RECT 216.200 177.900 216.600 179.900 ;
        RECT 218.400 178.200 218.800 179.900 ;
        RECT 218.400 177.900 219.400 178.200 ;
        RECT 214.200 177.500 214.600 177.900 ;
        RECT 216.300 177.600 216.600 177.900 ;
        RECT 215.900 177.300 217.700 177.600 ;
        RECT 219.000 177.500 219.400 177.900 ;
        RECT 215.900 177.200 216.300 177.300 ;
        RECT 217.300 177.200 217.700 177.300 ;
        RECT 213.800 176.600 214.500 177.000 ;
        RECT 214.200 176.100 214.500 176.600 ;
        RECT 215.300 176.500 216.400 176.800 ;
        RECT 215.300 176.400 215.700 176.500 ;
        RECT 214.200 175.800 215.400 176.100 ;
        RECT 211.800 175.300 213.900 175.600 ;
        RECT 206.200 174.800 206.600 175.200 ;
        RECT 207.400 174.900 208.200 175.200 ;
        RECT 207.800 174.800 208.200 174.900 ;
        RECT 205.500 174.400 205.900 174.800 ;
        RECT 205.500 174.200 205.800 174.400 ;
        RECT 199.800 173.900 200.300 174.100 ;
        RECT 195.900 173.300 197.800 173.600 ;
        RECT 195.900 173.200 196.300 173.300 ;
        RECT 190.200 172.100 190.600 172.500 ;
        RECT 191.000 172.400 191.400 172.800 ;
        RECT 191.900 172.700 192.300 172.800 ;
        RECT 191.900 172.400 193.300 172.700 ;
        RECT 193.000 172.100 193.300 172.400 ;
        RECT 195.000 172.100 195.400 172.500 ;
        RECT 190.200 171.800 191.200 172.100 ;
        RECT 190.800 171.100 191.200 171.800 ;
        RECT 193.000 171.100 193.400 172.100 ;
        RECT 195.000 171.800 195.700 172.100 ;
        RECT 195.100 171.100 195.700 171.800 ;
        RECT 197.400 171.100 197.800 173.300 ;
        RECT 198.200 173.600 200.300 173.900 ;
        RECT 200.800 173.800 201.800 174.200 ;
        RECT 205.400 173.800 205.800 174.200 ;
        RECT 198.200 172.500 198.500 173.600 ;
        RECT 200.800 173.500 201.100 173.800 ;
        RECT 200.700 173.300 201.100 173.500 ;
        RECT 200.300 173.000 201.100 173.300 ;
        RECT 206.200 173.100 206.500 174.800 ;
        RECT 207.000 173.800 207.400 174.600 ;
        RECT 209.400 174.400 209.800 175.200 ;
        RECT 210.100 174.800 210.600 175.200 ;
        RECT 210.100 174.200 210.400 174.800 ;
        RECT 208.600 174.100 209.000 174.200 ;
        RECT 208.600 173.800 209.400 174.100 ;
        RECT 210.100 173.800 211.400 174.200 ;
        RECT 209.000 173.600 209.400 173.800 ;
        RECT 208.700 173.100 210.500 173.300 ;
        RECT 211.000 173.100 211.300 173.800 ;
        RECT 211.800 173.600 212.200 175.300 ;
        RECT 213.500 175.200 213.900 175.300 ;
        RECT 212.700 174.900 213.100 175.000 ;
        RECT 212.700 174.600 214.600 174.900 ;
        RECT 214.200 174.500 214.600 174.600 ;
        RECT 215.100 174.200 215.400 175.800 ;
        RECT 216.100 175.900 216.400 176.500 ;
        RECT 216.700 176.500 217.100 176.600 ;
        RECT 219.000 176.500 219.400 176.600 ;
        RECT 216.700 176.200 219.400 176.500 ;
        RECT 216.100 175.700 218.500 175.900 ;
        RECT 220.600 175.700 221.000 179.900 ;
        RECT 223.300 176.400 223.700 179.900 ;
        RECT 225.400 177.500 225.800 179.500 ;
        RECT 216.100 175.600 221.000 175.700 ;
        RECT 222.900 176.100 223.700 176.400 ;
        RECT 218.100 175.500 221.000 175.600 ;
        RECT 218.200 175.400 221.000 175.500 ;
        RECT 215.800 175.100 216.200 175.200 ;
        RECT 217.400 175.100 217.800 175.200 ;
        RECT 215.800 174.800 219.900 175.100 ;
        RECT 222.200 174.800 222.600 175.600 ;
        RECT 219.500 174.700 219.900 174.800 ;
        RECT 218.700 174.200 219.100 174.300 ;
        RECT 222.900 174.200 223.200 176.100 ;
        RECT 225.500 175.800 225.800 177.500 ;
        RECT 223.900 175.500 225.800 175.800 ;
        RECT 226.200 177.500 226.600 179.500 ;
        RECT 226.200 175.800 226.500 177.500 ;
        RECT 228.300 176.400 228.700 179.900 ;
        RECT 232.900 176.400 233.300 179.900 ;
        RECT 235.000 177.500 235.400 179.500 ;
        RECT 228.300 176.100 229.100 176.400 ;
        RECT 226.200 175.500 228.100 175.800 ;
        RECT 223.900 174.500 224.200 175.500 ;
        RECT 215.100 173.900 220.600 174.200 ;
        RECT 215.300 173.800 215.700 173.900 ;
        RECT 211.800 173.300 213.700 173.600 ;
        RECT 198.200 171.500 198.600 172.500 ;
        RECT 200.300 171.500 200.700 173.000 ;
        RECT 205.900 172.200 206.700 173.100 ;
        RECT 205.400 171.800 206.700 172.200 ;
        RECT 205.900 171.100 206.700 171.800 ;
        RECT 208.600 173.000 210.600 173.100 ;
        RECT 208.600 171.100 209.000 173.000 ;
        RECT 210.200 171.100 210.600 173.000 ;
        RECT 211.000 171.100 211.400 173.100 ;
        RECT 211.800 171.100 212.200 173.300 ;
        RECT 213.300 173.200 213.700 173.300 ;
        RECT 218.200 173.200 218.500 173.900 ;
        RECT 219.800 173.800 220.600 173.900 ;
        RECT 221.400 174.100 221.800 174.200 ;
        RECT 222.200 174.100 223.200 174.200 ;
        RECT 223.500 174.100 224.200 174.500 ;
        RECT 224.600 174.400 225.000 175.200 ;
        RECT 225.400 174.400 225.800 175.200 ;
        RECT 226.200 174.400 226.600 175.200 ;
        RECT 227.000 174.400 227.400 175.200 ;
        RECT 227.800 174.500 228.100 175.500 ;
        RECT 221.400 173.800 223.200 174.100 ;
        RECT 222.900 173.500 223.200 173.800 ;
        RECT 223.700 173.900 224.200 174.100 ;
        RECT 227.800 174.100 228.500 174.500 ;
        RECT 228.800 174.200 229.100 176.100 ;
        RECT 232.500 176.100 233.300 176.400 ;
        RECT 229.400 175.100 229.800 175.600 ;
        RECT 230.200 175.100 230.600 175.200 ;
        RECT 229.400 174.800 230.600 175.100 ;
        RECT 231.800 174.800 232.200 175.600 ;
        RECT 232.500 174.200 232.800 176.100 ;
        RECT 235.100 175.800 235.400 177.500 ;
        RECT 233.500 175.500 235.400 175.800 ;
        RECT 233.500 174.500 233.800 175.500 ;
        RECT 227.800 173.900 228.300 174.100 ;
        RECT 223.700 173.600 225.800 173.900 ;
        RECT 217.300 172.700 217.700 172.800 ;
        RECT 214.200 172.100 214.600 172.500 ;
        RECT 216.300 172.400 217.700 172.700 ;
        RECT 218.200 172.400 218.600 173.200 ;
        RECT 216.300 172.100 216.600 172.400 ;
        RECT 219.000 172.100 219.400 172.500 ;
        RECT 213.900 171.800 214.600 172.100 ;
        RECT 213.900 171.100 214.500 171.800 ;
        RECT 216.200 171.100 216.600 172.100 ;
        RECT 218.400 171.800 219.400 172.100 ;
        RECT 218.400 171.100 218.800 171.800 ;
        RECT 220.600 171.100 221.000 173.500 ;
        RECT 222.900 173.300 223.300 173.500 ;
        RECT 222.900 173.000 223.700 173.300 ;
        RECT 223.300 171.500 223.700 173.000 ;
        RECT 225.500 172.500 225.800 173.600 ;
        RECT 225.400 171.500 225.800 172.500 ;
        RECT 226.200 173.600 228.300 173.900 ;
        RECT 228.800 173.800 229.800 174.200 ;
        RECT 231.000 174.100 231.400 174.200 ;
        RECT 231.800 174.100 232.800 174.200 ;
        RECT 233.100 174.100 233.800 174.500 ;
        RECT 234.200 174.400 234.600 175.200 ;
        RECT 235.000 174.400 235.400 175.200 ;
        RECT 231.000 173.800 232.800 174.100 ;
        RECT 226.200 172.500 226.500 173.600 ;
        RECT 228.800 173.500 229.100 173.800 ;
        RECT 228.700 173.300 229.100 173.500 ;
        RECT 228.300 173.200 229.100 173.300 ;
        RECT 227.800 173.000 229.100 173.200 ;
        RECT 232.500 173.500 232.800 173.800 ;
        RECT 233.300 173.900 233.800 174.100 ;
        RECT 233.300 173.600 235.400 173.900 ;
        RECT 232.500 173.300 232.900 173.500 ;
        RECT 232.500 173.000 233.300 173.300 ;
        RECT 227.800 172.800 228.700 173.000 ;
        RECT 226.200 171.500 226.600 172.500 ;
        RECT 228.300 171.500 228.700 172.800 ;
        RECT 232.900 171.500 233.300 173.000 ;
        RECT 235.100 172.500 235.400 173.600 ;
        RECT 235.800 173.400 236.200 174.200 ;
        RECT 236.600 173.100 237.000 179.900 ;
        RECT 237.400 175.800 237.800 176.600 ;
        RECT 238.200 175.600 238.600 179.900 ;
        RECT 240.300 177.900 240.900 179.900 ;
        RECT 242.600 177.900 243.000 179.900 ;
        RECT 244.800 178.200 245.200 179.900 ;
        RECT 244.800 177.900 245.800 178.200 ;
        RECT 240.600 177.500 241.000 177.900 ;
        RECT 242.700 177.600 243.000 177.900 ;
        RECT 242.300 177.300 244.100 177.600 ;
        RECT 245.400 177.500 245.800 177.900 ;
        RECT 242.300 177.200 242.700 177.300 ;
        RECT 243.700 177.200 244.100 177.300 ;
        RECT 240.200 176.600 240.900 177.000 ;
        RECT 240.600 176.100 240.900 176.600 ;
        RECT 241.700 176.500 242.800 176.800 ;
        RECT 241.700 176.400 242.100 176.500 ;
        RECT 240.600 175.800 241.800 176.100 ;
        RECT 238.200 175.300 240.300 175.600 ;
        RECT 238.200 173.600 238.600 175.300 ;
        RECT 239.900 175.200 240.300 175.300 ;
        RECT 241.500 175.100 241.800 175.800 ;
        RECT 242.500 175.900 242.800 176.500 ;
        RECT 243.100 176.500 243.500 176.600 ;
        RECT 245.400 176.500 245.800 176.600 ;
        RECT 243.100 176.200 245.800 176.500 ;
        RECT 242.500 175.700 244.900 175.900 ;
        RECT 247.000 175.700 247.400 179.900 ;
        RECT 249.100 176.200 249.500 179.900 ;
        RECT 249.800 176.800 250.200 177.200 ;
        RECT 249.900 176.200 250.200 176.800 ;
        RECT 248.600 175.800 249.600 176.200 ;
        RECT 249.900 175.900 250.600 176.200 ;
        RECT 250.200 175.800 250.600 175.900 ;
        RECT 242.500 175.600 247.400 175.700 ;
        RECT 244.500 175.500 247.400 175.600 ;
        RECT 244.600 175.400 247.400 175.500 ;
        RECT 242.200 175.100 242.600 175.200 ;
        RECT 239.100 174.900 239.500 175.000 ;
        RECT 239.100 174.600 241.000 174.900 ;
        RECT 241.400 174.800 242.600 175.100 ;
        RECT 243.800 175.100 244.200 175.200 ;
        RECT 243.800 174.800 246.300 175.100 ;
        RECT 240.600 174.500 241.000 174.600 ;
        RECT 241.500 174.200 241.800 174.800 ;
        RECT 244.600 174.700 245.000 174.800 ;
        RECT 245.900 174.700 246.300 174.800 ;
        RECT 248.600 174.400 249.000 175.200 ;
        RECT 245.100 174.200 245.500 174.300 ;
        RECT 249.300 174.200 249.600 175.800 ;
        RECT 241.500 173.900 247.000 174.200 ;
        RECT 241.700 173.800 242.100 173.900 ;
        RECT 238.200 173.300 240.100 173.600 ;
        RECT 236.600 172.800 237.500 173.100 ;
        RECT 235.000 171.500 235.400 172.500 ;
        RECT 237.100 172.200 237.500 172.800 ;
        RECT 236.600 171.800 237.500 172.200 ;
        RECT 237.100 171.100 237.500 171.800 ;
        RECT 238.200 171.100 238.600 173.300 ;
        RECT 239.700 173.200 240.100 173.300 ;
        RECT 244.600 172.800 244.900 173.900 ;
        RECT 246.200 173.800 247.000 173.900 ;
        RECT 247.800 174.100 248.200 174.200 ;
        RECT 247.800 173.800 248.600 174.100 ;
        RECT 249.300 173.800 250.600 174.200 ;
        RECT 248.200 173.600 248.600 173.800 ;
        RECT 243.700 172.700 244.100 172.800 ;
        RECT 240.600 172.100 241.000 172.500 ;
        RECT 242.700 172.400 244.100 172.700 ;
        RECT 244.600 172.400 245.000 172.800 ;
        RECT 242.700 172.100 243.000 172.400 ;
        RECT 245.400 172.100 245.800 172.500 ;
        RECT 240.300 171.800 241.000 172.100 ;
        RECT 240.300 171.100 240.900 171.800 ;
        RECT 242.600 171.100 243.000 172.100 ;
        RECT 244.800 171.800 245.800 172.100 ;
        RECT 244.800 171.100 245.200 171.800 ;
        RECT 247.000 171.100 247.400 173.500 ;
        RECT 247.900 173.100 249.700 173.300 ;
        RECT 250.200 173.100 250.500 173.800 ;
        RECT 247.800 173.000 249.800 173.100 ;
        RECT 247.800 171.100 248.200 173.000 ;
        RECT 249.400 171.100 249.800 173.000 ;
        RECT 250.200 171.100 250.600 173.100 ;
        RECT 1.400 167.600 1.800 169.900 ;
        RECT 3.000 167.600 3.400 169.900 ;
        RECT 4.600 167.600 5.000 169.900 ;
        RECT 6.200 167.600 6.600 169.900 ;
        RECT 0.600 167.200 1.800 167.600 ;
        RECT 2.300 167.200 3.400 167.600 ;
        RECT 3.900 167.200 5.000 167.600 ;
        RECT 5.700 167.200 6.600 167.600 ;
        RECT 7.800 167.500 8.200 169.900 ;
        RECT 10.000 169.200 10.400 169.900 ;
        RECT 9.400 168.900 10.400 169.200 ;
        RECT 12.200 168.900 12.600 169.900 ;
        RECT 14.300 169.200 14.900 169.900 ;
        RECT 14.200 168.900 14.900 169.200 ;
        RECT 9.400 168.500 9.800 168.900 ;
        RECT 12.200 168.600 12.500 168.900 ;
        RECT 10.200 168.200 10.600 168.600 ;
        RECT 11.100 168.300 12.500 168.600 ;
        RECT 14.200 168.500 14.600 168.900 ;
        RECT 11.100 168.200 11.500 168.300 ;
        RECT 0.600 165.800 1.000 167.200 ;
        RECT 2.300 166.900 2.700 167.200 ;
        RECT 3.900 166.900 4.300 167.200 ;
        RECT 5.700 166.900 6.100 167.200 ;
        RECT 7.000 167.100 7.400 167.200 ;
        RECT 8.200 167.100 9.000 167.200 ;
        RECT 10.300 167.100 10.600 168.200 ;
        RECT 15.100 167.700 15.500 167.800 ;
        RECT 16.600 167.700 17.000 169.900 ;
        RECT 17.400 167.900 17.800 169.900 ;
        RECT 18.200 168.000 18.600 169.900 ;
        RECT 19.800 168.000 20.200 169.900 ;
        RECT 18.200 167.900 20.200 168.000 ;
        RECT 15.100 167.400 17.000 167.700 ;
        RECT 11.800 167.100 12.200 167.200 ;
        RECT 13.100 167.100 13.500 167.200 ;
        RECT 7.000 166.900 13.700 167.100 ;
        RECT 1.400 166.500 2.700 166.900 ;
        RECT 3.100 166.500 4.300 166.900 ;
        RECT 4.800 166.500 6.100 166.900 ;
        RECT 6.500 166.800 13.700 166.900 ;
        RECT 6.500 166.500 7.400 166.800 ;
        RECT 9.700 166.700 10.100 166.800 ;
        RECT 2.300 165.800 2.700 166.500 ;
        RECT 3.900 165.800 4.300 166.500 ;
        RECT 5.700 165.800 6.100 166.500 ;
        RECT 8.900 166.200 9.300 166.300 ;
        RECT 8.900 165.900 11.400 166.200 ;
        RECT 11.000 165.800 11.400 165.900 ;
        RECT 0.600 165.400 1.800 165.800 ;
        RECT 2.300 165.400 3.400 165.800 ;
        RECT 3.900 165.400 5.000 165.800 ;
        RECT 5.700 165.400 6.600 165.800 ;
        RECT 1.400 161.100 1.800 165.400 ;
        RECT 3.000 161.100 3.400 165.400 ;
        RECT 4.600 161.100 5.000 165.400 ;
        RECT 6.200 161.100 6.600 165.400 ;
        RECT 7.800 165.500 10.600 165.600 ;
        RECT 7.800 165.400 10.700 165.500 ;
        RECT 7.800 165.300 12.700 165.400 ;
        RECT 7.800 161.100 8.200 165.300 ;
        RECT 10.300 165.100 12.700 165.300 ;
        RECT 9.400 164.500 12.100 164.800 ;
        RECT 9.400 164.400 9.800 164.500 ;
        RECT 11.700 164.400 12.100 164.500 ;
        RECT 12.400 164.500 12.700 165.100 ;
        RECT 13.400 165.200 13.700 166.800 ;
        RECT 14.200 166.400 14.600 166.500 ;
        RECT 14.200 166.100 16.100 166.400 ;
        RECT 15.700 166.000 16.100 166.100 ;
        RECT 14.900 165.700 15.300 165.800 ;
        RECT 16.600 165.700 17.000 167.400 ;
        RECT 17.500 167.200 17.800 167.900 ;
        RECT 18.300 167.700 20.100 167.900 ;
        RECT 20.600 167.500 21.000 169.900 ;
        RECT 22.800 169.200 23.200 169.900 ;
        RECT 22.200 168.900 23.200 169.200 ;
        RECT 25.000 168.900 25.400 169.900 ;
        RECT 27.100 169.200 27.700 169.900 ;
        RECT 27.000 168.900 27.700 169.200 ;
        RECT 22.200 168.500 22.600 168.900 ;
        RECT 25.000 168.600 25.300 168.900 ;
        RECT 23.000 167.800 23.400 168.600 ;
        RECT 23.900 168.300 25.300 168.600 ;
        RECT 27.000 168.500 27.400 168.900 ;
        RECT 23.900 168.200 24.300 168.300 ;
        RECT 19.400 167.200 19.800 167.400 ;
        RECT 17.400 166.800 18.700 167.200 ;
        RECT 19.400 166.900 20.200 167.200 ;
        RECT 19.800 166.800 20.200 166.900 ;
        RECT 21.000 167.100 21.800 167.200 ;
        RECT 23.100 167.100 23.400 167.800 ;
        RECT 27.900 167.700 28.300 167.800 ;
        RECT 29.400 167.700 29.800 169.900 ;
        RECT 31.500 168.200 31.900 169.900 ;
        RECT 27.900 167.400 29.800 167.700 ;
        RECT 31.000 167.900 31.900 168.200 ;
        RECT 32.600 167.900 33.000 169.900 ;
        RECT 33.400 168.000 33.800 169.900 ;
        RECT 35.000 168.000 35.400 169.900 ;
        RECT 37.700 168.000 38.100 169.500 ;
        RECT 39.800 168.500 40.200 169.500 ;
        RECT 33.400 167.900 35.400 168.000 ;
        RECT 25.900 167.100 26.300 167.200 ;
        RECT 21.000 166.800 26.500 167.100 ;
        RECT 14.900 165.400 17.000 165.700 ;
        RECT 13.400 164.900 14.600 165.200 ;
        RECT 13.100 164.500 13.500 164.600 ;
        RECT 12.400 164.200 13.500 164.500 ;
        RECT 14.300 164.400 14.600 164.900 ;
        RECT 14.300 164.000 15.000 164.400 ;
        RECT 11.100 163.700 11.500 163.800 ;
        RECT 12.500 163.700 12.900 163.800 ;
        RECT 9.400 163.100 9.800 163.500 ;
        RECT 11.100 163.400 12.900 163.700 ;
        RECT 12.200 163.100 12.500 163.400 ;
        RECT 14.200 163.100 14.600 163.500 ;
        RECT 9.400 162.800 10.400 163.100 ;
        RECT 10.000 161.100 10.400 162.800 ;
        RECT 12.200 161.100 12.600 163.100 ;
        RECT 14.300 161.100 14.900 163.100 ;
        RECT 16.600 161.100 17.000 165.400 ;
        RECT 17.400 165.100 17.800 165.200 ;
        RECT 18.400 165.100 18.700 166.800 ;
        RECT 22.500 166.700 22.900 166.800 ;
        RECT 19.000 165.800 19.400 166.600 ;
        RECT 21.700 166.200 22.100 166.300 ;
        RECT 21.700 166.100 24.200 166.200 ;
        RECT 25.400 166.100 25.800 166.200 ;
        RECT 21.700 165.900 25.800 166.100 ;
        RECT 23.800 165.800 25.800 165.900 ;
        RECT 20.600 165.500 23.400 165.600 ;
        RECT 20.600 165.400 23.500 165.500 ;
        RECT 20.600 165.300 25.500 165.400 ;
        RECT 17.400 164.800 18.100 165.100 ;
        RECT 18.400 164.800 18.900 165.100 ;
        RECT 17.800 164.200 18.100 164.800 ;
        RECT 18.500 164.200 18.900 164.800 ;
        RECT 17.800 163.800 18.200 164.200 ;
        RECT 18.500 163.800 19.400 164.200 ;
        RECT 18.500 161.100 18.900 163.800 ;
        RECT 20.600 161.100 21.000 165.300 ;
        RECT 23.100 165.100 25.500 165.300 ;
        RECT 22.200 164.500 24.900 164.800 ;
        RECT 22.200 164.400 22.600 164.500 ;
        RECT 24.500 164.400 24.900 164.500 ;
        RECT 25.200 164.500 25.500 165.100 ;
        RECT 26.200 165.200 26.500 166.800 ;
        RECT 27.000 166.400 27.400 166.500 ;
        RECT 27.000 166.100 28.900 166.400 ;
        RECT 28.500 166.000 28.900 166.100 ;
        RECT 27.700 165.700 28.100 165.800 ;
        RECT 29.400 165.700 29.800 167.400 ;
        RECT 30.200 166.800 30.600 167.600 ;
        RECT 27.700 165.400 29.800 165.700 ;
        RECT 26.200 164.900 27.400 165.200 ;
        RECT 25.900 164.500 26.300 164.600 ;
        RECT 25.200 164.200 26.300 164.500 ;
        RECT 27.100 164.400 27.400 164.900 ;
        RECT 27.100 164.000 27.800 164.400 ;
        RECT 23.900 163.700 24.300 163.800 ;
        RECT 25.300 163.700 25.700 163.800 ;
        RECT 22.200 163.100 22.600 163.500 ;
        RECT 23.900 163.400 25.700 163.700 ;
        RECT 25.000 163.100 25.300 163.400 ;
        RECT 27.000 163.100 27.400 163.500 ;
        RECT 22.200 162.800 23.200 163.100 ;
        RECT 22.800 161.100 23.200 162.800 ;
        RECT 25.000 161.100 25.400 163.100 ;
        RECT 27.100 161.100 27.700 163.100 ;
        RECT 29.400 161.100 29.800 165.400 ;
        RECT 31.000 166.100 31.400 167.900 ;
        RECT 32.700 167.200 33.000 167.900 ;
        RECT 33.500 167.700 35.300 167.900 ;
        RECT 37.300 167.700 38.100 168.000 ;
        RECT 37.300 167.500 37.700 167.700 ;
        RECT 34.600 167.200 35.000 167.400 ;
        RECT 37.300 167.200 37.600 167.500 ;
        RECT 39.900 167.400 40.200 168.500 ;
        RECT 41.900 169.200 42.300 169.900 ;
        RECT 41.900 168.800 42.600 169.200 ;
        RECT 41.900 168.200 42.300 168.800 ;
        RECT 41.400 167.900 42.300 168.200 ;
        RECT 44.900 168.200 45.300 169.500 ;
        RECT 47.000 168.500 47.400 169.500 ;
        RECT 44.900 168.000 45.800 168.200 ;
        RECT 32.600 166.800 33.900 167.200 ;
        RECT 34.600 166.900 35.400 167.200 ;
        RECT 35.000 166.800 35.400 166.900 ;
        RECT 36.600 166.800 37.600 167.200 ;
        RECT 38.100 167.100 40.200 167.400 ;
        RECT 38.100 166.900 38.600 167.100 ;
        RECT 31.000 165.800 32.900 166.100 ;
        RECT 31.000 161.100 31.400 165.800 ;
        RECT 32.600 165.200 32.900 165.800 ;
        RECT 31.800 164.400 32.200 165.200 ;
        RECT 32.600 165.100 33.000 165.200 ;
        RECT 33.600 165.100 33.900 166.800 ;
        RECT 34.200 165.800 34.600 166.600 ;
        RECT 35.800 166.100 36.200 166.200 ;
        RECT 36.600 166.100 37.000 166.200 ;
        RECT 35.800 165.800 37.000 166.100 ;
        RECT 36.600 165.400 37.000 165.800 ;
        RECT 32.600 164.800 33.300 165.100 ;
        RECT 33.600 164.800 34.100 165.100 ;
        RECT 33.000 164.200 33.300 164.800 ;
        RECT 33.000 163.800 33.400 164.200 ;
        RECT 33.700 161.100 34.100 164.800 ;
        RECT 37.300 164.900 37.600 166.800 ;
        RECT 37.900 166.500 38.600 166.900 ;
        RECT 40.600 166.800 41.000 167.600 ;
        RECT 38.300 165.500 38.600 166.500 ;
        RECT 39.000 165.800 39.400 166.600 ;
        RECT 39.800 165.800 40.200 166.600 ;
        RECT 40.600 166.200 40.900 166.800 ;
        RECT 40.600 165.800 41.000 166.200 ;
        RECT 38.300 165.200 40.200 165.500 ;
        RECT 37.300 164.600 38.100 164.900 ;
        RECT 37.700 164.200 38.100 164.600 ;
        RECT 37.700 163.800 38.600 164.200 ;
        RECT 37.700 161.100 38.100 163.800 ;
        RECT 39.900 163.500 40.200 165.200 ;
        RECT 39.800 161.500 40.200 163.500 ;
        RECT 41.400 161.100 41.800 167.900 ;
        RECT 44.500 167.800 45.800 168.000 ;
        RECT 44.500 167.700 45.300 167.800 ;
        RECT 44.500 167.500 44.900 167.700 ;
        RECT 44.500 167.200 44.800 167.500 ;
        RECT 47.100 167.400 47.400 168.500 ;
        RECT 50.700 167.900 51.500 169.900 ;
        RECT 43.800 166.800 44.800 167.200 ;
        RECT 45.300 167.100 47.400 167.400 ;
        RECT 45.300 166.900 45.800 167.100 ;
        RECT 43.800 165.400 44.200 166.200 ;
        RECT 42.200 164.400 42.600 165.200 ;
        RECT 44.500 164.900 44.800 166.800 ;
        RECT 45.100 166.500 45.800 166.900 ;
        RECT 50.200 166.800 50.600 167.200 ;
        RECT 50.300 166.600 50.600 166.800 ;
        RECT 45.500 165.500 45.800 166.500 ;
        RECT 46.200 165.800 46.600 166.600 ;
        RECT 47.000 165.800 47.400 166.600 ;
        RECT 50.300 166.200 50.700 166.600 ;
        RECT 51.000 166.200 51.300 167.900 ;
        RECT 53.400 167.500 53.800 169.900 ;
        RECT 55.600 169.200 56.000 169.900 ;
        RECT 55.000 168.900 56.000 169.200 ;
        RECT 57.800 168.900 58.200 169.900 ;
        RECT 59.900 169.200 60.500 169.900 ;
        RECT 59.800 168.900 60.500 169.200 ;
        RECT 55.000 168.500 55.400 168.900 ;
        RECT 57.800 168.600 58.100 168.900 ;
        RECT 55.800 167.800 56.200 168.600 ;
        RECT 56.700 168.300 58.100 168.600 ;
        RECT 59.800 168.500 60.200 168.900 ;
        RECT 56.700 168.200 57.100 168.300 ;
        RECT 51.800 166.400 52.200 167.200 ;
        RECT 53.800 167.100 54.600 167.200 ;
        RECT 55.900 167.100 56.200 167.800 ;
        RECT 60.700 167.700 61.100 167.800 ;
        RECT 62.200 167.700 62.600 169.900 ;
        RECT 63.000 168.000 63.400 169.900 ;
        RECT 64.600 168.000 65.000 169.900 ;
        RECT 63.000 167.900 65.000 168.000 ;
        RECT 65.400 167.900 65.800 169.900 ;
        RECT 66.500 168.200 66.900 169.900 ;
        RECT 68.600 168.500 69.000 169.500 ;
        RECT 70.700 169.200 71.100 169.500 ;
        RECT 70.200 168.800 71.100 169.200 ;
        RECT 66.500 167.900 67.400 168.200 ;
        RECT 63.100 167.700 64.900 167.900 ;
        RECT 60.700 167.400 62.600 167.700 ;
        RECT 58.700 167.100 59.100 167.200 ;
        RECT 53.800 166.800 59.300 167.100 ;
        RECT 55.300 166.700 55.700 166.800 ;
        RECT 54.500 166.200 54.900 166.300 ;
        RECT 47.800 166.100 48.200 166.200 ;
        RECT 49.400 166.100 49.800 166.200 ;
        RECT 47.800 165.800 49.800 166.100 ;
        RECT 45.500 165.200 47.400 165.500 ;
        RECT 49.400 165.400 49.800 165.800 ;
        RECT 51.000 165.800 51.400 166.200 ;
        RECT 52.600 166.100 53.000 166.200 ;
        RECT 52.200 165.800 53.000 166.100 ;
        RECT 54.500 165.900 57.000 166.200 ;
        RECT 56.600 165.800 57.000 165.900 ;
        RECT 51.000 165.700 51.300 165.800 ;
        RECT 50.300 165.400 51.300 165.700 ;
        RECT 52.200 165.600 52.600 165.800 ;
        RECT 53.400 165.500 56.200 165.600 ;
        RECT 53.400 165.400 56.300 165.500 ;
        RECT 44.500 164.600 45.300 164.900 ;
        RECT 44.900 161.100 45.300 164.600 ;
        RECT 47.100 163.500 47.400 165.200 ;
        RECT 50.300 165.100 50.600 165.400 ;
        RECT 53.400 165.300 58.300 165.400 ;
        RECT 47.000 161.500 47.400 163.500 ;
        RECT 49.400 161.400 49.800 165.100 ;
        RECT 50.200 161.700 50.600 165.100 ;
        RECT 51.000 164.800 53.000 165.100 ;
        RECT 51.000 161.400 51.400 164.800 ;
        RECT 49.400 161.100 51.400 161.400 ;
        RECT 52.600 161.100 53.000 164.800 ;
        RECT 53.400 161.100 53.800 165.300 ;
        RECT 55.900 165.100 58.300 165.300 ;
        RECT 55.000 164.500 57.700 164.800 ;
        RECT 55.000 164.400 55.400 164.500 ;
        RECT 57.300 164.400 57.700 164.500 ;
        RECT 58.000 164.500 58.300 165.100 ;
        RECT 59.000 165.200 59.300 166.800 ;
        RECT 59.800 166.400 60.200 166.500 ;
        RECT 59.800 166.100 61.700 166.400 ;
        RECT 61.300 166.000 61.700 166.100 ;
        RECT 60.500 165.700 60.900 165.800 ;
        RECT 62.200 165.700 62.600 167.400 ;
        RECT 63.400 167.200 63.800 167.400 ;
        RECT 65.400 167.200 65.700 167.900 ;
        RECT 63.000 166.900 63.800 167.200 ;
        RECT 63.000 166.800 63.400 166.900 ;
        RECT 64.500 166.800 65.800 167.200 ;
        RECT 63.800 165.800 64.200 166.600 ;
        RECT 60.500 165.400 62.600 165.700 ;
        RECT 59.000 164.900 60.200 165.200 ;
        RECT 58.700 164.500 59.100 164.600 ;
        RECT 58.000 164.200 59.100 164.500 ;
        RECT 59.900 164.400 60.200 164.900 ;
        RECT 59.900 164.000 60.600 164.400 ;
        RECT 56.700 163.700 57.100 163.800 ;
        RECT 58.100 163.700 58.500 163.800 ;
        RECT 55.000 163.100 55.400 163.500 ;
        RECT 56.700 163.400 58.500 163.700 ;
        RECT 57.800 163.100 58.100 163.400 ;
        RECT 59.800 163.100 60.200 163.500 ;
        RECT 55.000 162.800 56.000 163.100 ;
        RECT 55.600 161.100 56.000 162.800 ;
        RECT 57.800 161.100 58.200 163.100 ;
        RECT 59.900 161.100 60.500 163.100 ;
        RECT 62.200 161.100 62.600 165.400 ;
        RECT 64.500 165.200 64.800 166.800 ;
        RECT 67.000 166.100 67.400 167.900 ;
        RECT 67.800 166.800 68.200 167.600 ;
        RECT 68.600 167.400 68.900 168.500 ;
        RECT 70.700 168.000 71.100 168.800 ;
        RECT 75.300 168.000 75.700 169.500 ;
        RECT 77.400 168.500 77.800 169.500 ;
        RECT 70.700 167.700 71.500 168.000 ;
        RECT 71.100 167.500 71.500 167.700 ;
        RECT 68.600 167.100 70.700 167.400 ;
        RECT 70.200 166.900 70.700 167.100 ;
        RECT 71.200 167.200 71.500 167.500 ;
        RECT 74.900 167.700 75.700 168.000 ;
        RECT 74.900 167.500 75.300 167.700 ;
        RECT 74.900 167.200 75.200 167.500 ;
        RECT 77.500 167.400 77.800 168.500 ;
        RECT 78.200 168.000 78.600 169.900 ;
        RECT 79.800 168.000 80.200 169.900 ;
        RECT 78.200 167.900 80.200 168.000 ;
        RECT 80.600 167.900 81.000 169.900 ;
        RECT 81.700 168.200 82.100 169.900 ;
        RECT 81.700 167.900 82.600 168.200 ;
        RECT 85.100 167.900 85.900 169.900 ;
        RECT 78.300 167.700 80.100 167.900 ;
        RECT 63.800 164.800 64.800 165.200 ;
        RECT 65.400 165.800 67.400 166.100 ;
        RECT 68.600 165.800 69.000 166.600 ;
        RECT 69.400 165.800 69.800 166.600 ;
        RECT 70.200 166.500 70.900 166.900 ;
        RECT 71.200 166.800 72.200 167.200 ;
        RECT 74.200 166.800 75.200 167.200 ;
        RECT 75.700 167.100 77.800 167.400 ;
        RECT 78.600 167.200 79.000 167.400 ;
        RECT 80.600 167.200 80.900 167.900 ;
        RECT 75.700 166.900 76.200 167.100 ;
        RECT 65.400 165.200 65.700 165.800 ;
        RECT 65.400 165.100 65.800 165.200 ;
        RECT 65.100 164.800 65.800 165.100 ;
        RECT 64.300 161.100 64.700 164.800 ;
        RECT 65.100 164.200 65.400 164.800 ;
        RECT 66.200 164.400 66.600 165.200 ;
        RECT 65.000 163.800 65.400 164.200 ;
        RECT 67.000 161.100 67.400 165.800 ;
        RECT 70.200 165.500 70.500 166.500 ;
        RECT 68.600 165.200 70.500 165.500 ;
        RECT 68.600 163.500 68.900 165.200 ;
        RECT 71.200 164.900 71.500 166.800 ;
        RECT 71.800 166.100 72.200 166.200 ;
        RECT 72.600 166.100 73.000 166.200 ;
        RECT 71.800 165.800 73.000 166.100 ;
        RECT 73.400 166.100 73.800 166.200 ;
        RECT 74.200 166.100 74.600 166.200 ;
        RECT 73.400 165.800 74.600 166.100 ;
        RECT 71.800 165.400 72.200 165.800 ;
        RECT 74.200 165.400 74.600 165.800 ;
        RECT 70.700 164.600 71.500 164.900 ;
        RECT 74.900 164.900 75.200 166.800 ;
        RECT 75.500 166.500 76.200 166.900 ;
        RECT 78.200 166.900 79.000 167.200 ;
        RECT 79.700 167.100 81.000 167.200 ;
        RECT 81.400 167.100 81.800 167.200 ;
        RECT 78.200 166.800 78.600 166.900 ;
        RECT 79.700 166.800 81.800 167.100 ;
        RECT 75.900 165.500 76.200 166.500 ;
        RECT 76.600 165.800 77.000 166.600 ;
        RECT 77.400 165.800 77.800 166.600 ;
        RECT 79.000 165.800 79.400 166.600 ;
        RECT 75.900 165.200 77.800 165.500 ;
        RECT 74.900 164.600 75.700 164.900 ;
        RECT 68.600 161.500 69.000 163.500 ;
        RECT 70.700 161.100 71.100 164.600 ;
        RECT 75.300 161.100 75.700 164.600 ;
        RECT 77.500 163.500 77.800 165.200 ;
        RECT 79.700 165.100 80.000 166.800 ;
        RECT 82.200 166.100 82.600 167.900 ;
        RECT 83.000 167.100 83.400 167.600 ;
        RECT 83.800 167.100 84.200 167.200 ;
        RECT 83.000 166.800 84.200 167.100 ;
        RECT 84.600 166.800 85.000 167.200 ;
        RECT 84.700 166.600 85.000 166.800 ;
        RECT 84.700 166.200 85.100 166.600 ;
        RECT 85.400 166.200 85.700 167.900 ;
        RECT 87.800 167.700 88.200 169.900 ;
        RECT 89.900 169.200 90.500 169.900 ;
        RECT 89.900 168.900 90.600 169.200 ;
        RECT 92.200 168.900 92.600 169.900 ;
        RECT 94.400 169.200 94.800 169.900 ;
        RECT 94.400 168.900 95.400 169.200 ;
        RECT 90.200 168.500 90.600 168.900 ;
        RECT 92.300 168.600 92.600 168.900 ;
        RECT 92.300 168.300 93.700 168.600 ;
        RECT 93.300 168.200 93.700 168.300 ;
        RECT 94.200 168.200 94.600 168.600 ;
        RECT 95.000 168.500 95.400 168.900 ;
        RECT 89.300 167.700 89.700 167.800 ;
        RECT 87.800 167.400 89.700 167.700 ;
        RECT 86.200 166.400 86.600 167.200 ;
        RECT 80.600 165.800 82.600 166.100 ;
        RECT 80.600 165.200 80.900 165.800 ;
        RECT 80.600 165.100 81.000 165.200 ;
        RECT 77.400 161.500 77.800 163.500 ;
        RECT 79.500 164.800 80.000 165.100 ;
        RECT 80.300 164.800 81.000 165.100 ;
        RECT 79.500 161.100 79.900 164.800 ;
        RECT 80.300 164.200 80.600 164.800 ;
        RECT 81.400 164.400 81.800 165.200 ;
        RECT 80.200 163.800 80.600 164.200 ;
        RECT 82.200 161.100 82.600 165.800 ;
        RECT 83.800 165.400 84.200 166.200 ;
        RECT 85.400 165.800 85.800 166.200 ;
        RECT 87.000 166.100 87.400 166.200 ;
        RECT 86.600 165.800 87.400 166.100 ;
        RECT 85.400 165.700 85.700 165.800 ;
        RECT 84.700 165.400 85.700 165.700 ;
        RECT 86.600 165.600 87.000 165.800 ;
        RECT 87.800 165.700 88.200 167.400 ;
        RECT 91.300 167.100 91.700 167.200 ;
        RECT 94.200 167.100 94.500 168.200 ;
        RECT 96.600 167.500 97.000 169.900 ;
        RECT 98.700 168.200 99.100 169.900 ;
        RECT 98.200 167.900 99.100 168.200 ;
        RECT 101.400 167.900 101.800 169.900 ;
        RECT 102.200 168.000 102.600 169.900 ;
        RECT 103.800 168.000 104.200 169.900 ;
        RECT 102.200 167.900 104.200 168.000 ;
        RECT 95.800 167.100 96.600 167.200 ;
        RECT 91.100 166.800 96.600 167.100 ;
        RECT 97.400 166.800 97.800 167.600 ;
        RECT 90.200 166.400 90.600 166.500 ;
        RECT 88.700 166.100 90.600 166.400 ;
        RECT 88.700 166.000 89.100 166.100 ;
        RECT 89.500 165.700 89.900 165.800 ;
        RECT 87.800 165.400 89.900 165.700 ;
        RECT 84.700 165.100 85.000 165.400 ;
        RECT 83.800 161.400 84.200 165.100 ;
        RECT 84.600 161.700 85.000 165.100 ;
        RECT 85.400 164.800 87.400 165.100 ;
        RECT 85.400 161.400 85.800 164.800 ;
        RECT 83.800 161.100 85.800 161.400 ;
        RECT 87.000 161.100 87.400 164.800 ;
        RECT 87.800 161.100 88.200 165.400 ;
        RECT 91.100 165.200 91.400 166.800 ;
        RECT 94.700 166.700 95.100 166.800 ;
        RECT 94.200 166.200 94.600 166.300 ;
        RECT 95.500 166.200 95.900 166.300 ;
        RECT 93.400 165.900 95.900 166.200 ;
        RECT 98.200 166.100 98.600 167.900 ;
        RECT 101.500 167.200 101.800 167.900 ;
        RECT 102.300 167.700 104.100 167.900 ;
        RECT 104.600 167.500 105.000 169.900 ;
        RECT 106.800 169.200 107.200 169.900 ;
        RECT 106.200 168.900 107.200 169.200 ;
        RECT 109.000 168.900 109.400 169.900 ;
        RECT 111.100 169.200 111.700 169.900 ;
        RECT 111.000 168.900 111.700 169.200 ;
        RECT 106.200 168.500 106.600 168.900 ;
        RECT 109.000 168.600 109.300 168.900 ;
        RECT 107.000 168.200 107.400 168.600 ;
        RECT 107.900 168.300 109.300 168.600 ;
        RECT 111.000 168.500 111.400 168.900 ;
        RECT 107.900 168.200 108.300 168.300 ;
        RECT 103.400 167.200 103.800 167.400 ;
        RECT 101.400 166.800 102.700 167.200 ;
        RECT 103.400 166.900 104.200 167.200 ;
        RECT 103.800 166.800 104.200 166.900 ;
        RECT 105.000 167.100 105.800 167.200 ;
        RECT 107.100 167.100 107.400 168.200 ;
        RECT 111.900 167.700 112.300 167.800 ;
        RECT 113.400 167.700 113.800 169.900 ;
        RECT 114.200 168.000 114.600 169.900 ;
        RECT 115.800 168.000 116.200 169.900 ;
        RECT 114.200 167.900 116.200 168.000 ;
        RECT 116.600 167.900 117.000 169.900 ;
        RECT 117.700 168.200 118.100 169.900 ;
        RECT 121.700 169.200 122.100 169.500 ;
        RECT 121.700 168.800 122.600 169.200 ;
        RECT 117.700 167.900 118.600 168.200 ;
        RECT 121.700 168.000 122.100 168.800 ;
        RECT 123.800 168.500 124.200 169.500 ;
        RECT 114.300 167.700 116.100 167.900 ;
        RECT 111.900 167.400 113.800 167.700 ;
        RECT 108.600 167.100 109.000 167.200 ;
        RECT 109.900 167.100 110.300 167.200 ;
        RECT 105.000 166.800 110.500 167.100 ;
        RECT 93.400 165.800 93.800 165.900 ;
        RECT 98.200 165.800 101.700 166.100 ;
        RECT 94.200 165.500 97.000 165.600 ;
        RECT 94.100 165.400 97.000 165.500 ;
        RECT 90.200 164.900 91.400 165.200 ;
        RECT 92.100 165.300 97.000 165.400 ;
        RECT 92.100 165.100 94.500 165.300 ;
        RECT 90.200 164.400 90.500 164.900 ;
        RECT 89.800 164.000 90.500 164.400 ;
        RECT 91.300 164.500 91.700 164.600 ;
        RECT 92.100 164.500 92.400 165.100 ;
        RECT 91.300 164.200 92.400 164.500 ;
        RECT 92.700 164.500 95.400 164.800 ;
        RECT 92.700 164.400 93.100 164.500 ;
        RECT 95.000 164.400 95.400 164.500 ;
        RECT 91.900 163.700 92.300 163.800 ;
        RECT 93.300 163.700 93.700 163.800 ;
        RECT 90.200 163.100 90.600 163.500 ;
        RECT 91.900 163.400 93.700 163.700 ;
        RECT 92.300 163.100 92.600 163.400 ;
        RECT 95.000 163.100 95.400 163.500 ;
        RECT 89.900 161.100 90.500 163.100 ;
        RECT 92.200 161.100 92.600 163.100 ;
        RECT 94.400 162.800 95.400 163.100 ;
        RECT 94.400 161.100 94.800 162.800 ;
        RECT 96.600 161.100 97.000 165.300 ;
        RECT 98.200 161.100 98.600 165.800 ;
        RECT 101.400 165.200 101.700 165.800 ;
        RECT 99.000 164.400 99.400 165.200 ;
        RECT 101.400 165.100 101.800 165.200 ;
        RECT 102.400 165.100 102.700 166.800 ;
        RECT 106.500 166.700 106.900 166.800 ;
        RECT 103.000 165.800 103.400 166.600 ;
        RECT 105.700 166.200 106.100 166.300 ;
        RECT 105.700 165.900 108.200 166.200 ;
        RECT 107.800 165.800 108.200 165.900 ;
        RECT 104.600 165.500 107.400 165.600 ;
        RECT 104.600 165.400 107.500 165.500 ;
        RECT 104.600 165.300 109.500 165.400 ;
        RECT 101.400 164.800 102.100 165.100 ;
        RECT 102.400 164.800 102.900 165.100 ;
        RECT 101.800 164.200 102.100 164.800 ;
        RECT 101.800 163.800 102.200 164.200 ;
        RECT 102.500 161.100 102.900 164.800 ;
        RECT 104.600 161.100 105.000 165.300 ;
        RECT 107.100 165.100 109.500 165.300 ;
        RECT 106.200 164.500 108.900 164.800 ;
        RECT 106.200 164.400 106.600 164.500 ;
        RECT 108.500 164.400 108.900 164.500 ;
        RECT 109.200 164.500 109.500 165.100 ;
        RECT 110.200 165.200 110.500 166.800 ;
        RECT 111.000 166.400 111.400 166.500 ;
        RECT 111.000 166.100 112.900 166.400 ;
        RECT 112.500 166.000 112.900 166.100 ;
        RECT 111.700 165.700 112.100 165.800 ;
        RECT 113.400 165.700 113.800 167.400 ;
        RECT 114.600 167.200 115.000 167.400 ;
        RECT 116.600 167.200 116.900 167.900 ;
        RECT 114.200 166.900 115.000 167.200 ;
        RECT 114.200 166.800 114.600 166.900 ;
        RECT 115.700 166.800 117.000 167.200 ;
        RECT 114.200 166.100 114.600 166.200 ;
        RECT 115.000 166.100 115.400 166.600 ;
        RECT 114.200 165.800 115.400 166.100 ;
        RECT 115.700 166.200 116.000 166.800 ;
        RECT 115.700 165.800 116.200 166.200 ;
        RECT 118.200 166.100 118.600 167.900 ;
        RECT 121.300 167.700 122.100 168.000 ;
        RECT 119.000 167.100 119.400 167.600 ;
        RECT 121.300 167.500 121.700 167.700 ;
        RECT 121.300 167.200 121.600 167.500 ;
        RECT 123.900 167.400 124.200 168.500 ;
        RECT 125.900 168.200 126.300 169.900 ;
        RECT 125.400 167.900 126.300 168.200 ;
        RECT 127.000 167.900 127.400 169.900 ;
        RECT 127.800 168.000 128.200 169.900 ;
        RECT 129.400 168.000 129.800 169.900 ;
        RECT 127.800 167.900 129.800 168.000 ;
        RECT 130.500 169.200 130.900 169.900 ;
        RECT 130.500 168.800 131.400 169.200 ;
        RECT 130.500 168.200 130.900 168.800 ;
        RECT 130.500 167.900 131.400 168.200 ;
        RECT 119.000 166.800 120.100 167.100 ;
        RECT 120.600 166.800 121.600 167.200 ;
        RECT 122.100 167.100 124.200 167.400 ;
        RECT 122.100 166.900 122.600 167.100 ;
        RECT 116.600 165.800 118.600 166.100 ;
        RECT 119.800 166.100 120.100 166.800 ;
        RECT 120.600 166.100 121.000 166.200 ;
        RECT 119.800 165.800 121.000 166.100 ;
        RECT 111.700 165.400 113.800 165.700 ;
        RECT 110.200 164.900 111.400 165.200 ;
        RECT 109.900 164.500 110.300 164.600 ;
        RECT 109.200 164.200 110.300 164.500 ;
        RECT 111.100 164.400 111.400 164.900 ;
        RECT 111.100 164.200 111.800 164.400 ;
        RECT 111.100 164.000 112.200 164.200 ;
        RECT 111.500 163.800 112.200 164.000 ;
        RECT 107.900 163.700 108.300 163.800 ;
        RECT 109.300 163.700 109.700 163.800 ;
        RECT 106.200 163.100 106.600 163.500 ;
        RECT 107.900 163.400 109.700 163.700 ;
        RECT 109.000 163.100 109.300 163.400 ;
        RECT 111.000 163.100 111.400 163.500 ;
        RECT 106.200 162.800 107.200 163.100 ;
        RECT 106.800 161.100 107.200 162.800 ;
        RECT 109.000 161.100 109.400 163.100 ;
        RECT 111.100 161.100 111.700 163.100 ;
        RECT 113.400 161.100 113.800 165.400 ;
        RECT 115.700 165.100 116.000 165.800 ;
        RECT 116.600 165.200 116.900 165.800 ;
        RECT 116.600 165.100 117.000 165.200 ;
        RECT 115.500 164.800 116.000 165.100 ;
        RECT 116.300 164.800 117.000 165.100 ;
        RECT 115.500 161.100 115.900 164.800 ;
        RECT 116.300 164.200 116.600 164.800 ;
        RECT 117.400 164.400 117.800 165.200 ;
        RECT 116.200 163.800 116.600 164.200 ;
        RECT 118.200 161.100 118.600 165.800 ;
        RECT 120.600 165.400 121.000 165.800 ;
        RECT 121.300 164.900 121.600 166.800 ;
        RECT 121.900 166.500 122.600 166.900 ;
        RECT 124.600 166.800 125.000 167.600 ;
        RECT 122.300 165.500 122.600 166.500 ;
        RECT 123.000 165.800 123.400 166.600 ;
        RECT 123.800 165.800 124.200 166.600 ;
        RECT 125.400 166.100 125.800 167.900 ;
        RECT 127.100 167.200 127.400 167.900 ;
        RECT 127.900 167.700 129.700 167.900 ;
        RECT 129.000 167.200 129.400 167.400 ;
        RECT 127.000 166.800 128.300 167.200 ;
        RECT 129.000 166.900 129.800 167.200 ;
        RECT 129.400 166.800 129.800 166.900 ;
        RECT 125.400 165.800 127.300 166.100 ;
        RECT 122.300 165.200 124.200 165.500 ;
        RECT 121.300 164.600 122.100 164.900 ;
        RECT 121.700 161.100 122.100 164.600 ;
        RECT 123.900 163.500 124.200 165.200 ;
        RECT 123.800 161.500 124.200 163.500 ;
        RECT 125.400 161.100 125.800 165.800 ;
        RECT 127.000 165.200 127.300 165.800 ;
        RECT 128.000 165.200 128.300 166.800 ;
        RECT 128.600 165.800 129.000 166.600 ;
        RECT 126.200 164.400 126.600 165.200 ;
        RECT 127.000 165.100 127.400 165.200 ;
        RECT 127.000 164.800 127.700 165.100 ;
        RECT 128.000 164.800 129.000 165.200 ;
        RECT 127.400 164.200 127.700 164.800 ;
        RECT 127.400 163.800 127.800 164.200 ;
        RECT 128.100 161.100 128.500 164.800 ;
        RECT 130.200 164.400 130.600 165.200 ;
        RECT 131.000 161.100 131.400 167.900 ;
        RECT 132.600 167.700 133.000 169.900 ;
        RECT 134.700 169.200 135.300 169.900 ;
        RECT 134.700 168.900 135.400 169.200 ;
        RECT 137.000 168.900 137.400 169.900 ;
        RECT 139.200 169.200 139.600 169.900 ;
        RECT 139.200 168.900 140.200 169.200 ;
        RECT 135.000 168.500 135.400 168.900 ;
        RECT 137.100 168.600 137.400 168.900 ;
        RECT 137.100 168.300 138.500 168.600 ;
        RECT 138.100 168.200 138.500 168.300 ;
        RECT 139.000 168.200 139.400 168.600 ;
        RECT 139.800 168.500 140.200 168.900 ;
        RECT 134.100 167.700 134.500 167.800 ;
        RECT 131.800 166.800 132.200 167.600 ;
        RECT 132.600 167.400 134.500 167.700 ;
        RECT 132.600 165.700 133.000 167.400 ;
        RECT 136.100 167.100 136.500 167.200 ;
        RECT 137.400 167.100 137.800 167.200 ;
        RECT 139.000 167.100 139.300 168.200 ;
        RECT 141.400 167.500 141.800 169.900 ;
        RECT 142.200 168.000 142.600 169.900 ;
        RECT 143.800 168.000 144.200 169.900 ;
        RECT 142.200 167.900 144.200 168.000 ;
        RECT 144.600 167.900 145.000 169.900 ;
        RECT 142.300 167.700 144.100 167.900 ;
        RECT 142.600 167.200 143.000 167.400 ;
        RECT 144.600 167.200 144.900 167.900 ;
        RECT 145.400 167.700 145.800 169.900 ;
        RECT 147.500 169.200 148.100 169.900 ;
        RECT 147.500 168.900 148.200 169.200 ;
        RECT 149.800 168.900 150.200 169.900 ;
        RECT 152.000 169.200 152.400 169.900 ;
        RECT 152.000 168.900 153.000 169.200 ;
        RECT 147.800 168.500 148.200 168.900 ;
        RECT 149.900 168.600 150.200 168.900 ;
        RECT 149.900 168.300 151.300 168.600 ;
        RECT 150.900 168.200 151.300 168.300 ;
        RECT 151.800 167.800 152.200 168.600 ;
        RECT 152.600 168.500 153.000 168.900 ;
        RECT 146.900 167.700 147.300 167.800 ;
        RECT 145.400 167.400 147.300 167.700 ;
        RECT 140.600 167.100 141.400 167.200 ;
        RECT 135.900 166.800 141.400 167.100 ;
        RECT 142.200 166.900 143.000 167.200 ;
        RECT 142.200 166.800 142.600 166.900 ;
        RECT 143.700 166.800 145.000 167.200 ;
        RECT 135.000 166.400 135.400 166.500 ;
        RECT 133.500 166.100 135.400 166.400 ;
        RECT 133.500 166.000 133.900 166.100 ;
        RECT 134.300 165.700 134.700 165.800 ;
        RECT 132.600 165.400 134.700 165.700 ;
        RECT 132.600 161.100 133.000 165.400 ;
        RECT 135.900 165.200 136.200 166.800 ;
        RECT 139.500 166.700 139.900 166.800 ;
        RECT 140.300 166.200 140.700 166.300 ;
        RECT 138.200 165.900 140.700 166.200 ;
        RECT 142.200 166.100 142.600 166.200 ;
        RECT 143.000 166.100 143.400 166.600 ;
        RECT 138.200 165.800 138.600 165.900 ;
        RECT 142.200 165.800 143.400 166.100 ;
        RECT 139.000 165.500 141.800 165.600 ;
        RECT 138.900 165.400 141.800 165.500 ;
        RECT 135.000 164.900 136.200 165.200 ;
        RECT 136.900 165.300 141.800 165.400 ;
        RECT 136.900 165.100 139.300 165.300 ;
        RECT 135.000 164.400 135.300 164.900 ;
        RECT 134.600 164.000 135.300 164.400 ;
        RECT 136.100 164.500 136.500 164.600 ;
        RECT 136.900 164.500 137.200 165.100 ;
        RECT 136.100 164.200 137.200 164.500 ;
        RECT 137.500 164.500 140.200 164.800 ;
        RECT 137.500 164.400 137.900 164.500 ;
        RECT 139.800 164.400 140.200 164.500 ;
        RECT 136.700 163.700 137.100 163.800 ;
        RECT 138.100 163.700 138.500 163.800 ;
        RECT 135.000 163.100 135.400 163.500 ;
        RECT 136.700 163.400 138.500 163.700 ;
        RECT 137.100 163.100 137.400 163.400 ;
        RECT 139.800 163.100 140.200 163.500 ;
        RECT 134.700 161.100 135.300 163.100 ;
        RECT 137.000 161.100 137.400 163.100 ;
        RECT 139.200 162.800 140.200 163.100 ;
        RECT 139.200 161.100 139.600 162.800 ;
        RECT 141.400 161.100 141.800 165.300 ;
        RECT 143.700 165.100 144.000 166.800 ;
        RECT 145.400 165.700 145.800 167.400 ;
        RECT 148.900 167.100 149.300 167.200 ;
        RECT 151.800 167.100 152.100 167.800 ;
        RECT 154.200 167.500 154.600 169.900 ;
        RECT 156.600 168.500 157.000 169.500 ;
        RECT 156.600 167.400 156.900 168.500 ;
        RECT 158.700 168.000 159.100 169.500 ;
        RECT 158.700 167.700 159.500 168.000 ;
        RECT 162.700 167.900 163.500 169.900 ;
        RECT 165.400 168.000 165.800 169.900 ;
        RECT 167.000 168.000 167.400 169.900 ;
        RECT 165.400 167.900 167.400 168.000 ;
        RECT 167.800 167.900 168.200 169.900 ;
        RECT 168.900 168.200 169.300 169.900 ;
        RECT 171.000 168.500 171.400 169.500 ;
        RECT 168.900 167.900 169.800 168.200 ;
        RECT 159.100 167.500 159.500 167.700 ;
        RECT 153.400 167.100 154.200 167.200 ;
        RECT 156.600 167.100 158.700 167.400 ;
        RECT 148.700 166.800 154.200 167.100 ;
        RECT 158.200 166.900 158.700 167.100 ;
        RECT 159.200 167.200 159.500 167.500 ;
        RECT 159.200 167.100 160.200 167.200 ;
        RECT 162.200 167.100 162.600 167.200 ;
        RECT 147.800 166.400 148.200 166.500 ;
        RECT 146.300 166.100 148.200 166.400 ;
        RECT 146.300 166.000 146.700 166.100 ;
        RECT 147.100 165.700 147.500 165.800 ;
        RECT 145.400 165.400 147.500 165.700 ;
        RECT 144.600 165.100 145.000 165.200 ;
        RECT 143.500 164.800 144.000 165.100 ;
        RECT 144.300 164.800 145.000 165.100 ;
        RECT 143.500 161.100 143.900 164.800 ;
        RECT 144.300 164.200 144.600 164.800 ;
        RECT 144.200 163.800 144.600 164.200 ;
        RECT 145.400 161.100 145.800 165.400 ;
        RECT 148.700 165.200 149.000 166.800 ;
        RECT 152.300 166.700 152.700 166.800 ;
        RECT 153.100 166.200 153.500 166.300 ;
        RECT 150.200 166.100 150.600 166.200 ;
        RECT 151.000 166.100 153.500 166.200 ;
        RECT 150.200 165.900 153.500 166.100 ;
        RECT 150.200 165.800 151.400 165.900 ;
        RECT 156.600 165.800 157.000 166.600 ;
        RECT 157.400 165.800 157.800 166.600 ;
        RECT 158.200 166.500 158.900 166.900 ;
        RECT 159.200 166.800 162.600 167.100 ;
        RECT 151.800 165.500 154.600 165.600 ;
        RECT 158.200 165.500 158.500 166.500 ;
        RECT 151.700 165.400 154.600 165.500 ;
        RECT 147.800 164.900 149.000 165.200 ;
        RECT 149.700 165.300 154.600 165.400 ;
        RECT 149.700 165.100 152.100 165.300 ;
        RECT 147.800 164.400 148.100 164.900 ;
        RECT 147.400 164.000 148.100 164.400 ;
        RECT 148.900 164.500 149.300 164.600 ;
        RECT 149.700 164.500 150.000 165.100 ;
        RECT 148.900 164.200 150.000 164.500 ;
        RECT 150.300 164.500 153.000 164.800 ;
        RECT 150.300 164.400 150.700 164.500 ;
        RECT 152.600 164.400 153.000 164.500 ;
        RECT 149.500 163.700 149.900 163.800 ;
        RECT 150.900 163.700 151.300 163.800 ;
        RECT 147.800 163.100 148.200 163.500 ;
        RECT 149.500 163.400 151.300 163.700 ;
        RECT 149.900 163.100 150.200 163.400 ;
        RECT 152.600 163.100 153.000 163.500 ;
        RECT 147.500 161.100 148.100 163.100 ;
        RECT 149.800 161.100 150.200 163.100 ;
        RECT 152.000 162.800 153.000 163.100 ;
        RECT 152.000 161.100 152.400 162.800 ;
        RECT 154.200 161.100 154.600 165.300 ;
        RECT 156.600 165.200 158.500 165.500 ;
        RECT 156.600 163.500 156.900 165.200 ;
        RECT 159.200 164.900 159.500 166.800 ;
        RECT 162.300 166.600 162.600 166.800 ;
        RECT 162.300 166.200 162.700 166.600 ;
        RECT 163.000 166.200 163.300 167.900 ;
        RECT 165.500 167.700 167.300 167.900 ;
        RECT 165.800 167.200 166.200 167.400 ;
        RECT 167.800 167.200 168.100 167.900 ;
        RECT 163.800 166.400 164.200 167.200 ;
        RECT 165.400 166.900 166.200 167.200 ;
        RECT 165.400 166.800 165.800 166.900 ;
        RECT 166.900 166.800 168.200 167.200 ;
        RECT 159.800 165.400 160.200 166.200 ;
        RECT 161.400 165.400 161.800 166.200 ;
        RECT 163.000 165.800 163.400 166.200 ;
        RECT 164.600 166.100 165.000 166.200 ;
        RECT 164.200 165.800 165.000 166.100 ;
        RECT 165.400 166.100 165.800 166.200 ;
        RECT 166.200 166.100 166.600 166.600 ;
        RECT 165.400 165.800 166.600 166.100 ;
        RECT 163.000 165.700 163.300 165.800 ;
        RECT 162.300 165.400 163.300 165.700 ;
        RECT 164.200 165.600 164.600 165.800 ;
        RECT 162.300 165.100 162.600 165.400 ;
        RECT 166.900 165.100 167.200 166.800 ;
        RECT 169.400 166.100 169.800 167.900 ;
        RECT 170.200 166.800 170.600 167.600 ;
        RECT 171.000 167.400 171.300 168.500 ;
        RECT 173.100 168.000 173.500 169.500 ;
        RECT 175.800 168.500 176.200 169.500 ;
        RECT 177.900 169.200 178.300 169.500 ;
        RECT 177.400 168.800 178.300 169.200 ;
        RECT 173.100 167.700 173.900 168.000 ;
        RECT 173.500 167.500 173.900 167.700 ;
        RECT 171.000 167.100 173.100 167.400 ;
        RECT 172.600 166.900 173.100 167.100 ;
        RECT 173.600 167.200 173.900 167.500 ;
        RECT 175.800 167.400 176.100 168.500 ;
        RECT 177.900 168.000 178.300 168.800 ;
        RECT 180.900 169.200 181.300 169.900 ;
        RECT 180.900 168.800 181.800 169.200 ;
        RECT 180.900 168.200 181.300 168.800 ;
        RECT 177.900 167.700 178.700 168.000 ;
        RECT 180.900 167.900 181.800 168.200 ;
        RECT 178.300 167.500 178.700 167.700 ;
        RECT 173.600 167.100 174.600 167.200 ;
        RECT 175.000 167.100 175.400 167.200 ;
        RECT 175.800 167.100 177.900 167.400 ;
        RECT 167.800 165.800 169.800 166.100 ;
        RECT 171.000 165.800 171.400 166.600 ;
        RECT 171.800 165.800 172.200 166.600 ;
        RECT 172.600 166.500 173.300 166.900 ;
        RECT 173.600 166.800 175.400 167.100 ;
        RECT 177.400 166.900 177.900 167.100 ;
        RECT 178.400 167.200 178.700 167.500 ;
        RECT 167.800 165.200 168.100 165.800 ;
        RECT 167.800 165.100 168.200 165.200 ;
        RECT 158.700 164.600 159.500 164.900 ;
        RECT 156.600 161.500 157.000 163.500 ;
        RECT 158.700 161.100 159.100 164.600 ;
        RECT 161.400 161.400 161.800 165.100 ;
        RECT 162.200 161.700 162.600 165.100 ;
        RECT 163.000 164.800 165.000 165.100 ;
        RECT 163.000 161.400 163.400 164.800 ;
        RECT 161.400 161.100 163.400 161.400 ;
        RECT 164.600 161.100 165.000 164.800 ;
        RECT 166.700 164.800 167.200 165.100 ;
        RECT 167.500 164.800 168.200 165.100 ;
        RECT 166.700 161.100 167.100 164.800 ;
        RECT 167.500 164.200 167.800 164.800 ;
        RECT 168.600 164.400 169.000 165.200 ;
        RECT 167.400 163.800 167.800 164.200 ;
        RECT 169.400 161.100 169.800 165.800 ;
        RECT 172.600 165.500 172.900 166.500 ;
        RECT 171.000 165.200 172.900 165.500 ;
        RECT 171.000 163.500 171.300 165.200 ;
        RECT 173.600 164.900 173.900 166.800 ;
        RECT 174.200 165.400 174.600 166.200 ;
        RECT 175.800 165.800 176.200 166.600 ;
        RECT 176.600 165.800 177.000 166.600 ;
        RECT 177.400 166.500 178.100 166.900 ;
        RECT 178.400 166.800 179.400 167.200 ;
        RECT 177.400 165.500 177.700 166.500 ;
        RECT 173.100 164.600 173.900 164.900 ;
        RECT 175.800 165.200 177.700 165.500 ;
        RECT 171.000 161.500 171.400 163.500 ;
        RECT 173.100 161.100 173.500 164.600 ;
        RECT 175.800 163.500 176.100 165.200 ;
        RECT 178.400 164.900 178.700 166.800 ;
        RECT 179.000 166.100 179.400 166.200 ;
        RECT 179.800 166.100 180.200 166.200 ;
        RECT 179.000 165.800 180.200 166.100 ;
        RECT 179.000 165.400 179.400 165.800 ;
        RECT 177.900 164.600 178.700 164.900 ;
        RECT 175.800 161.500 176.200 163.500 ;
        RECT 177.900 161.100 178.300 164.600 ;
        RECT 180.600 164.400 181.000 165.200 ;
        RECT 181.400 161.100 181.800 167.900 ;
        RECT 183.000 167.700 183.400 169.900 ;
        RECT 185.100 169.200 185.700 169.900 ;
        RECT 185.100 168.900 185.800 169.200 ;
        RECT 187.400 168.900 187.800 169.900 ;
        RECT 189.600 169.200 190.000 169.900 ;
        RECT 189.600 168.900 190.600 169.200 ;
        RECT 185.400 168.500 185.800 168.900 ;
        RECT 187.500 168.600 187.800 168.900 ;
        RECT 187.500 168.300 188.900 168.600 ;
        RECT 188.500 168.200 188.900 168.300 ;
        RECT 189.400 168.200 189.800 168.600 ;
        RECT 190.200 168.500 190.600 168.900 ;
        RECT 184.500 167.700 184.900 167.800 ;
        RECT 182.200 166.800 182.600 167.600 ;
        RECT 183.000 167.400 184.900 167.700 ;
        RECT 183.000 165.700 183.400 167.400 ;
        RECT 189.400 167.200 189.700 168.200 ;
        RECT 191.800 167.500 192.200 169.900 ;
        RECT 192.600 168.000 193.000 169.900 ;
        RECT 194.200 168.000 194.600 169.900 ;
        RECT 192.600 167.900 194.600 168.000 ;
        RECT 195.000 167.900 195.400 169.900 ;
        RECT 196.100 168.200 196.500 169.900 ;
        RECT 198.200 168.500 198.600 169.500 ;
        RECT 200.300 169.200 200.700 169.500 ;
        RECT 200.300 168.800 201.000 169.200 ;
        RECT 196.100 167.900 197.000 168.200 ;
        RECT 192.700 167.700 194.500 167.900 ;
        RECT 193.000 167.200 193.400 167.400 ;
        RECT 195.000 167.200 195.300 167.900 ;
        RECT 186.500 167.100 186.900 167.200 ;
        RECT 189.400 167.100 189.800 167.200 ;
        RECT 191.000 167.100 191.800 167.200 ;
        RECT 186.300 166.800 191.800 167.100 ;
        RECT 192.600 166.900 193.400 167.200 ;
        RECT 192.600 166.800 193.000 166.900 ;
        RECT 194.100 166.800 195.400 167.200 ;
        RECT 185.400 166.400 185.800 166.500 ;
        RECT 183.900 166.100 185.800 166.400 ;
        RECT 183.900 166.000 184.300 166.100 ;
        RECT 184.700 165.700 185.100 165.800 ;
        RECT 183.000 165.400 185.100 165.700 ;
        RECT 183.000 161.100 183.400 165.400 ;
        RECT 186.300 165.200 186.600 166.800 ;
        RECT 189.900 166.700 190.300 166.800 ;
        RECT 190.700 166.200 191.100 166.300 ;
        RECT 187.000 166.100 187.400 166.200 ;
        RECT 188.600 166.100 191.100 166.200 ;
        RECT 187.000 165.900 191.100 166.100 ;
        RECT 187.000 165.800 189.000 165.900 ;
        RECT 193.400 165.800 193.800 166.600 ;
        RECT 189.400 165.500 192.200 165.600 ;
        RECT 189.300 165.400 192.200 165.500 ;
        RECT 185.400 164.900 186.600 165.200 ;
        RECT 187.300 165.300 192.200 165.400 ;
        RECT 187.300 165.100 189.700 165.300 ;
        RECT 185.400 164.400 185.700 164.900 ;
        RECT 185.000 164.000 185.700 164.400 ;
        RECT 186.500 164.500 186.900 164.600 ;
        RECT 187.300 164.500 187.600 165.100 ;
        RECT 186.500 164.200 187.600 164.500 ;
        RECT 187.900 164.500 190.600 164.800 ;
        RECT 187.900 164.400 188.300 164.500 ;
        RECT 190.200 164.400 190.600 164.500 ;
        RECT 187.100 163.700 187.500 163.800 ;
        RECT 188.500 163.700 188.900 163.800 ;
        RECT 185.400 163.100 185.800 163.500 ;
        RECT 187.100 163.400 188.900 163.700 ;
        RECT 187.500 163.100 187.800 163.400 ;
        RECT 190.200 163.100 190.600 163.500 ;
        RECT 185.100 161.100 185.700 163.100 ;
        RECT 187.400 161.100 187.800 163.100 ;
        RECT 189.600 162.800 190.600 163.100 ;
        RECT 189.600 161.100 190.000 162.800 ;
        RECT 191.800 161.100 192.200 165.300 ;
        RECT 194.100 165.100 194.400 166.800 ;
        RECT 196.600 166.100 197.000 167.900 ;
        RECT 197.400 166.800 197.800 167.600 ;
        RECT 198.200 167.400 198.500 168.500 ;
        RECT 200.300 168.000 200.700 168.800 ;
        RECT 204.600 168.500 205.000 169.500 ;
        RECT 200.300 167.700 201.100 168.000 ;
        RECT 200.700 167.500 201.100 167.700 ;
        RECT 198.200 167.100 200.300 167.400 ;
        RECT 199.800 166.900 200.300 167.100 ;
        RECT 200.800 167.200 201.100 167.500 ;
        RECT 204.600 167.400 204.900 168.500 ;
        RECT 206.700 168.200 207.100 169.500 ;
        RECT 210.700 169.200 211.100 169.900 ;
        RECT 210.700 168.800 211.400 169.200 ;
        RECT 210.700 168.200 211.100 168.800 ;
        RECT 213.100 168.200 213.500 169.900 ;
        RECT 206.200 168.000 207.100 168.200 ;
        RECT 206.200 167.800 207.500 168.000 ;
        RECT 206.700 167.700 207.500 167.800 ;
        RECT 207.100 167.500 207.500 167.700 ;
        RECT 210.200 167.900 211.100 168.200 ;
        RECT 212.600 167.900 213.500 168.200 ;
        RECT 195.000 165.800 197.000 166.100 ;
        RECT 198.200 165.800 198.600 166.600 ;
        RECT 199.000 165.800 199.400 166.600 ;
        RECT 199.800 166.500 200.500 166.900 ;
        RECT 200.800 166.800 201.800 167.200 ;
        RECT 204.600 167.100 206.700 167.400 ;
        RECT 206.200 166.900 206.700 167.100 ;
        RECT 207.200 167.200 207.500 167.500 ;
        RECT 195.000 165.200 195.300 165.800 ;
        RECT 195.000 165.100 195.400 165.200 ;
        RECT 193.900 164.800 194.400 165.100 ;
        RECT 194.700 164.800 195.400 165.100 ;
        RECT 193.900 161.100 194.300 164.800 ;
        RECT 194.700 164.200 195.000 164.800 ;
        RECT 195.800 164.400 196.200 165.200 ;
        RECT 194.600 163.800 195.000 164.200 ;
        RECT 196.600 161.100 197.000 165.800 ;
        RECT 199.800 165.500 200.100 166.500 ;
        RECT 198.200 165.200 200.100 165.500 ;
        RECT 198.200 163.500 198.500 165.200 ;
        RECT 200.800 164.900 201.100 166.800 ;
        RECT 201.400 165.400 201.800 166.200 ;
        RECT 204.600 165.800 205.000 166.600 ;
        RECT 205.400 165.800 205.800 166.600 ;
        RECT 206.200 166.500 206.900 166.900 ;
        RECT 207.200 166.800 208.200 167.200 ;
        RECT 208.600 167.100 209.000 167.200 ;
        RECT 209.400 167.100 209.800 167.600 ;
        RECT 208.600 166.800 209.800 167.100 ;
        RECT 206.200 165.500 206.500 166.500 ;
        RECT 200.300 164.600 201.100 164.900 ;
        RECT 204.600 165.200 206.500 165.500 ;
        RECT 198.200 161.500 198.600 163.500 ;
        RECT 200.300 161.100 200.700 164.600 ;
        RECT 204.600 163.500 204.900 165.200 ;
        RECT 207.200 164.900 207.500 166.800 ;
        RECT 207.800 166.100 208.200 166.200 ;
        RECT 207.800 165.800 209.700 166.100 ;
        RECT 207.800 165.400 208.200 165.800 ;
        RECT 206.700 164.600 207.500 164.900 ;
        RECT 209.400 165.200 209.700 165.800 ;
        RECT 209.400 164.800 209.800 165.200 ;
        RECT 204.600 161.500 205.000 163.500 ;
        RECT 206.700 161.100 207.100 164.600 ;
        RECT 210.200 161.100 210.600 167.900 ;
        RECT 211.800 166.800 212.200 167.600 ;
        RECT 212.600 166.100 213.000 167.900 ;
        RECT 214.200 167.800 214.600 169.900 ;
        RECT 215.000 168.000 215.400 169.900 ;
        RECT 216.600 168.000 217.000 169.900 ;
        RECT 215.000 167.900 217.000 168.000 ;
        RECT 214.300 167.200 214.600 167.800 ;
        RECT 215.100 167.700 216.900 167.900 ;
        RECT 217.400 167.700 217.800 169.900 ;
        RECT 219.500 169.200 220.100 169.900 ;
        RECT 219.500 168.900 220.200 169.200 ;
        RECT 221.800 168.900 222.200 169.900 ;
        RECT 224.000 169.200 224.400 169.900 ;
        RECT 224.000 168.900 225.000 169.200 ;
        RECT 219.800 168.500 220.200 168.900 ;
        RECT 221.900 168.600 222.200 168.900 ;
        RECT 221.900 168.300 223.300 168.600 ;
        RECT 222.900 168.200 223.300 168.300 ;
        RECT 223.800 168.200 224.200 168.600 ;
        RECT 224.600 168.500 225.000 168.900 ;
        RECT 218.900 167.700 219.300 167.800 ;
        RECT 217.400 167.400 219.300 167.700 ;
        RECT 216.200 167.200 216.600 167.400 ;
        RECT 214.200 166.800 215.500 167.200 ;
        RECT 216.200 166.900 217.000 167.200 ;
        RECT 216.600 166.800 217.000 166.900 ;
        RECT 212.600 165.800 214.500 166.100 ;
        RECT 211.000 164.400 211.400 165.200 ;
        RECT 212.600 161.100 213.000 165.800 ;
        RECT 214.200 165.200 214.500 165.800 ;
        RECT 213.400 164.400 213.800 165.200 ;
        RECT 214.200 165.100 214.600 165.200 ;
        RECT 215.200 165.100 215.500 166.800 ;
        RECT 215.800 165.800 216.200 166.600 ;
        RECT 217.400 165.700 217.800 167.400 ;
        RECT 220.900 167.100 221.300 167.200 ;
        RECT 223.800 167.100 224.100 168.200 ;
        RECT 226.200 167.500 226.600 169.900 ;
        RECT 227.800 167.600 228.200 169.900 ;
        RECT 229.400 167.600 229.800 169.900 ;
        RECT 231.000 167.600 231.400 169.900 ;
        RECT 232.600 167.600 233.000 169.900 ;
        RECT 227.000 167.200 228.200 167.600 ;
        RECT 228.700 167.200 229.800 167.600 ;
        RECT 230.300 167.200 231.400 167.600 ;
        RECT 232.100 167.200 233.000 167.600 ;
        RECT 234.200 167.700 234.600 169.900 ;
        RECT 236.300 169.200 236.900 169.900 ;
        RECT 236.300 168.900 237.000 169.200 ;
        RECT 238.600 168.900 239.000 169.900 ;
        RECT 240.800 169.200 241.200 169.900 ;
        RECT 240.800 168.900 241.800 169.200 ;
        RECT 236.600 168.500 237.000 168.900 ;
        RECT 238.700 168.600 239.000 168.900 ;
        RECT 238.700 168.300 240.100 168.600 ;
        RECT 239.700 168.200 240.100 168.300 ;
        RECT 240.600 168.200 241.000 168.600 ;
        RECT 241.400 168.500 241.800 168.900 ;
        RECT 237.400 167.800 237.800 168.200 ;
        RECT 235.700 167.700 236.100 167.800 ;
        RECT 234.200 167.400 236.100 167.700 ;
        RECT 225.400 167.100 226.200 167.200 ;
        RECT 220.700 166.800 226.200 167.100 ;
        RECT 219.800 166.400 220.200 166.500 ;
        RECT 218.300 166.100 220.200 166.400 ;
        RECT 218.300 166.000 218.700 166.100 ;
        RECT 219.100 165.700 219.500 165.800 ;
        RECT 217.400 165.400 219.500 165.700 ;
        RECT 214.200 164.800 214.900 165.100 ;
        RECT 215.200 164.800 215.700 165.100 ;
        RECT 214.600 164.200 214.900 164.800 ;
        RECT 214.600 163.800 215.000 164.200 ;
        RECT 215.300 161.100 215.700 164.800 ;
        RECT 217.400 161.100 217.800 165.400 ;
        RECT 220.700 165.200 221.000 166.800 ;
        RECT 224.300 166.700 224.700 166.800 ;
        RECT 225.100 166.200 225.500 166.300 ;
        RECT 221.400 166.100 221.800 166.200 ;
        RECT 223.000 166.100 225.500 166.200 ;
        RECT 221.400 165.900 225.500 166.100 ;
        RECT 221.400 165.800 223.400 165.900 ;
        RECT 227.000 165.800 227.400 167.200 ;
        RECT 228.700 166.900 229.100 167.200 ;
        RECT 230.300 166.900 230.700 167.200 ;
        RECT 232.100 166.900 232.500 167.200 ;
        RECT 233.400 166.900 233.800 167.200 ;
        RECT 227.800 166.500 229.100 166.900 ;
        RECT 229.500 166.500 230.700 166.900 ;
        RECT 231.200 166.500 232.500 166.900 ;
        RECT 232.900 166.500 233.800 166.900 ;
        RECT 228.700 165.800 229.100 166.500 ;
        RECT 230.300 165.800 230.700 166.500 ;
        RECT 232.100 165.800 232.500 166.500 ;
        RECT 223.800 165.500 226.600 165.600 ;
        RECT 223.700 165.400 226.600 165.500 ;
        RECT 227.000 165.400 228.200 165.800 ;
        RECT 228.700 165.400 229.800 165.800 ;
        RECT 230.300 165.400 231.400 165.800 ;
        RECT 232.100 165.400 233.000 165.800 ;
        RECT 219.800 164.900 221.000 165.200 ;
        RECT 221.700 165.300 226.600 165.400 ;
        RECT 221.700 165.100 224.100 165.300 ;
        RECT 219.800 164.400 220.100 164.900 ;
        RECT 219.400 164.000 220.100 164.400 ;
        RECT 220.900 164.500 221.300 164.600 ;
        RECT 221.700 164.500 222.000 165.100 ;
        RECT 220.900 164.200 222.000 164.500 ;
        RECT 222.300 164.500 225.000 164.800 ;
        RECT 222.300 164.400 222.700 164.500 ;
        RECT 224.600 164.400 225.000 164.500 ;
        RECT 221.500 163.700 221.900 163.800 ;
        RECT 222.900 163.700 223.300 163.800 ;
        RECT 219.800 163.100 220.200 163.500 ;
        RECT 221.500 163.400 223.300 163.700 ;
        RECT 221.900 163.100 222.200 163.400 ;
        RECT 224.600 163.100 225.000 163.500 ;
        RECT 219.500 161.100 220.100 163.100 ;
        RECT 221.800 161.100 222.200 163.100 ;
        RECT 224.000 162.800 225.000 163.100 ;
        RECT 224.000 161.100 224.400 162.800 ;
        RECT 226.200 161.100 226.600 165.300 ;
        RECT 227.800 161.100 228.200 165.400 ;
        RECT 229.400 161.100 229.800 165.400 ;
        RECT 231.000 161.100 231.400 165.400 ;
        RECT 232.600 161.100 233.000 165.400 ;
        RECT 234.200 165.700 234.600 167.400 ;
        RECT 237.400 167.200 237.700 167.800 ;
        RECT 237.400 167.100 238.100 167.200 ;
        RECT 240.600 167.100 240.900 168.200 ;
        RECT 243.000 167.500 243.400 169.900 ;
        RECT 244.600 168.200 245.000 169.900 ;
        RECT 244.500 167.900 245.000 168.200 ;
        RECT 244.500 167.200 244.800 167.900 ;
        RECT 246.200 167.600 246.600 169.900 ;
        RECT 247.000 167.800 247.400 169.900 ;
        RECT 247.800 168.000 248.200 169.900 ;
        RECT 249.400 168.000 249.800 169.900 ;
        RECT 247.800 167.900 249.800 168.000 ;
        RECT 245.300 167.300 246.600 167.600 ;
        RECT 242.200 167.100 243.000 167.200 ;
        RECT 237.400 166.800 243.000 167.100 ;
        RECT 244.500 166.800 245.000 167.200 ;
        RECT 236.600 166.400 237.000 166.500 ;
        RECT 235.100 166.100 237.000 166.400 ;
        RECT 235.100 166.000 235.500 166.100 ;
        RECT 235.900 165.700 236.300 165.800 ;
        RECT 234.200 165.400 236.300 165.700 ;
        RECT 234.200 161.100 234.600 165.400 ;
        RECT 237.500 165.200 237.800 166.800 ;
        RECT 241.100 166.700 241.500 166.800 ;
        RECT 240.600 166.200 241.000 166.300 ;
        RECT 241.900 166.200 242.300 166.300 ;
        RECT 239.800 165.900 242.300 166.200 ;
        RECT 239.800 165.800 240.200 165.900 ;
        RECT 240.600 165.500 243.400 165.600 ;
        RECT 240.500 165.400 243.400 165.500 ;
        RECT 236.600 164.900 237.800 165.200 ;
        RECT 238.500 165.300 243.400 165.400 ;
        RECT 238.500 165.100 240.900 165.300 ;
        RECT 236.600 164.400 236.900 164.900 ;
        RECT 236.200 164.000 236.900 164.400 ;
        RECT 237.700 164.500 238.100 164.600 ;
        RECT 238.500 164.500 238.800 165.100 ;
        RECT 237.700 164.200 238.800 164.500 ;
        RECT 239.100 164.500 241.800 164.800 ;
        RECT 239.100 164.400 239.500 164.500 ;
        RECT 241.400 164.400 241.800 164.500 ;
        RECT 238.300 163.700 238.700 163.800 ;
        RECT 239.700 163.700 240.100 163.800 ;
        RECT 236.600 163.100 237.000 163.500 ;
        RECT 238.300 163.400 240.100 163.700 ;
        RECT 238.700 163.100 239.000 163.400 ;
        RECT 241.400 163.100 241.800 163.500 ;
        RECT 236.300 161.100 236.900 163.100 ;
        RECT 238.600 161.100 239.000 163.100 ;
        RECT 240.800 162.800 241.800 163.100 ;
        RECT 240.800 161.100 241.200 162.800 ;
        RECT 243.000 161.100 243.400 165.300 ;
        RECT 244.500 165.100 244.800 166.800 ;
        RECT 245.300 166.500 245.600 167.300 ;
        RECT 247.100 167.200 247.400 167.800 ;
        RECT 247.900 167.700 249.700 167.900 ;
        RECT 249.000 167.200 249.400 167.400 ;
        RECT 247.000 166.800 248.300 167.200 ;
        RECT 249.000 166.900 249.800 167.200 ;
        RECT 249.400 166.800 249.800 166.900 ;
        RECT 245.100 166.100 245.600 166.500 ;
        RECT 245.300 165.100 245.600 166.100 ;
        RECT 246.100 166.200 246.500 166.600 ;
        RECT 246.100 165.800 246.600 166.200 ;
        RECT 247.000 165.100 247.400 165.200 ;
        RECT 248.000 165.100 248.300 166.800 ;
        RECT 248.600 165.800 249.000 166.600 ;
        RECT 244.500 164.600 245.000 165.100 ;
        RECT 245.300 164.800 246.600 165.100 ;
        RECT 247.000 164.800 247.700 165.100 ;
        RECT 248.000 164.800 248.500 165.100 ;
        RECT 244.600 161.100 245.000 164.600 ;
        RECT 246.200 161.100 246.600 164.800 ;
        RECT 247.400 164.200 247.700 164.800 ;
        RECT 247.400 163.800 247.800 164.200 ;
        RECT 248.100 161.100 248.500 164.800 ;
        RECT 0.600 155.700 1.000 159.900 ;
        RECT 2.800 158.200 3.200 159.900 ;
        RECT 2.200 157.900 3.200 158.200 ;
        RECT 5.000 157.900 5.400 159.900 ;
        RECT 7.100 157.900 7.700 159.900 ;
        RECT 2.200 157.500 2.600 157.900 ;
        RECT 5.000 157.600 5.300 157.900 ;
        RECT 3.900 157.300 5.700 157.600 ;
        RECT 7.000 157.500 7.400 157.900 ;
        RECT 3.900 157.200 4.300 157.300 ;
        RECT 5.300 157.200 5.700 157.300 ;
        RECT 9.400 157.100 9.800 159.900 ;
        RECT 10.200 157.100 10.600 157.200 ;
        RECT 2.200 156.500 2.600 156.600 ;
        RECT 4.500 156.500 4.900 156.600 ;
        RECT 2.200 156.200 4.900 156.500 ;
        RECT 5.200 156.500 6.300 156.800 ;
        RECT 5.200 155.900 5.500 156.500 ;
        RECT 5.900 156.400 6.300 156.500 ;
        RECT 7.100 156.600 7.800 157.000 ;
        RECT 9.400 156.800 10.600 157.100 ;
        RECT 7.100 156.100 7.400 156.600 ;
        RECT 3.100 155.700 5.500 155.900 ;
        RECT 0.600 155.600 5.500 155.700 ;
        RECT 6.200 155.800 7.400 156.100 ;
        RECT 0.600 155.500 3.500 155.600 ;
        RECT 0.600 155.400 3.400 155.500 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 4.600 155.100 5.000 155.200 ;
        RECT 1.700 154.800 5.000 155.100 ;
        RECT 1.700 154.700 2.100 154.800 ;
        RECT 2.500 154.200 2.900 154.300 ;
        RECT 6.200 154.200 6.500 155.800 ;
        RECT 9.400 155.600 9.800 156.800 ;
        RECT 7.700 155.300 9.800 155.600 ;
        RECT 7.700 155.200 8.100 155.300 ;
        RECT 8.500 154.900 8.900 155.000 ;
        RECT 7.000 154.600 8.900 154.900 ;
        RECT 7.000 154.500 7.400 154.600 ;
        RECT 1.000 153.900 6.500 154.200 ;
        RECT 1.000 153.800 1.800 153.900 ;
        RECT 0.600 151.100 1.000 153.500 ;
        RECT 3.100 152.800 3.400 153.900 ;
        RECT 5.900 153.800 6.300 153.900 ;
        RECT 9.400 153.600 9.800 155.300 ;
        RECT 11.000 155.100 11.400 159.900 ;
        RECT 13.000 156.800 13.400 157.200 ;
        RECT 11.800 155.800 12.200 156.600 ;
        RECT 13.000 156.200 13.300 156.800 ;
        RECT 13.700 156.200 14.100 159.900 ;
        RECT 17.700 156.400 18.100 159.900 ;
        RECT 19.800 157.500 20.200 159.500 ;
        RECT 12.600 155.900 13.300 156.200 ;
        RECT 13.600 155.900 14.100 156.200 ;
        RECT 17.300 156.100 18.100 156.400 ;
        RECT 12.600 155.800 13.000 155.900 ;
        RECT 12.600 155.100 12.900 155.800 ;
        RECT 13.600 155.200 13.900 155.900 ;
        RECT 11.000 154.800 12.900 155.100 ;
        RECT 13.400 154.800 13.900 155.200 ;
        RECT 7.900 153.300 9.800 153.600 ;
        RECT 10.200 153.400 10.600 154.200 ;
        RECT 7.900 153.200 8.300 153.300 ;
        RECT 2.200 152.100 2.600 152.500 ;
        RECT 3.000 152.400 3.400 152.800 ;
        RECT 3.900 152.700 4.300 152.800 ;
        RECT 3.900 152.400 5.300 152.700 ;
        RECT 5.000 152.100 5.300 152.400 ;
        RECT 7.000 152.100 7.400 152.500 ;
        RECT 2.200 151.800 3.200 152.100 ;
        RECT 2.800 151.100 3.200 151.800 ;
        RECT 5.000 151.100 5.400 152.100 ;
        RECT 7.000 151.800 7.700 152.100 ;
        RECT 7.100 151.100 7.700 151.800 ;
        RECT 9.400 151.100 9.800 153.300 ;
        RECT 11.000 153.100 11.400 154.800 ;
        RECT 13.600 154.200 13.900 154.800 ;
        RECT 14.200 154.400 14.600 155.200 ;
        RECT 15.800 155.100 16.200 155.200 ;
        RECT 16.600 155.100 17.000 155.600 ;
        RECT 15.800 154.800 17.000 155.100 ;
        RECT 17.300 154.200 17.600 156.100 ;
        RECT 19.900 155.800 20.200 157.500 ;
        RECT 21.900 156.200 22.300 159.900 ;
        RECT 22.600 156.800 23.000 157.200 ;
        RECT 22.700 156.200 23.000 156.800 ;
        RECT 21.900 155.900 22.400 156.200 ;
        RECT 22.700 155.900 23.400 156.200 ;
        RECT 18.300 155.500 20.200 155.800 ;
        RECT 18.300 154.500 18.600 155.500 ;
        RECT 12.600 153.800 13.900 154.200 ;
        RECT 15.000 154.100 15.400 154.200 ;
        RECT 14.600 153.800 15.400 154.100 ;
        RECT 16.600 153.800 17.600 154.200 ;
        RECT 17.900 154.100 18.600 154.500 ;
        RECT 19.000 154.400 19.400 155.200 ;
        RECT 19.800 154.400 20.200 155.200 ;
        RECT 21.400 154.400 21.800 155.200 ;
        RECT 22.100 154.200 22.400 155.900 ;
        RECT 23.000 155.800 23.400 155.900 ;
        RECT 23.800 155.800 24.200 156.600 ;
        RECT 23.000 155.100 23.300 155.800 ;
        RECT 24.600 155.100 25.000 159.900 ;
        RECT 23.000 154.800 25.000 155.100 ;
        RECT 12.700 153.100 13.000 153.800 ;
        RECT 14.600 153.600 15.000 153.800 ;
        RECT 17.300 153.500 17.600 153.800 ;
        RECT 18.100 153.900 18.600 154.100 ;
        RECT 20.600 154.100 21.000 154.200 ;
        RECT 18.100 153.600 20.200 153.900 ;
        RECT 20.600 153.800 21.400 154.100 ;
        RECT 22.100 153.800 23.400 154.200 ;
        RECT 21.000 153.600 21.400 153.800 ;
        RECT 17.300 153.300 17.700 153.500 ;
        RECT 13.500 153.100 15.300 153.300 ;
        RECT 11.000 152.800 11.900 153.100 ;
        RECT 11.500 151.100 11.900 152.800 ;
        RECT 12.600 151.100 13.000 153.100 ;
        RECT 13.400 153.000 15.400 153.100 ;
        RECT 17.300 153.000 18.100 153.300 ;
        RECT 13.400 151.100 13.800 153.000 ;
        RECT 15.000 151.100 15.400 153.000 ;
        RECT 17.700 152.200 18.100 153.000 ;
        RECT 19.900 152.500 20.200 153.600 ;
        RECT 20.700 153.100 22.500 153.300 ;
        RECT 23.000 153.200 23.300 153.800 ;
        RECT 17.700 151.800 18.600 152.200 ;
        RECT 17.700 151.500 18.100 151.800 ;
        RECT 19.800 151.500 20.200 152.500 ;
        RECT 20.600 153.000 22.600 153.100 ;
        RECT 20.600 151.100 21.000 153.000 ;
        RECT 22.200 151.100 22.600 153.000 ;
        RECT 23.000 151.100 23.400 153.200 ;
        RECT 24.600 153.100 25.000 154.800 ;
        RECT 26.200 155.600 26.600 159.900 ;
        RECT 28.300 157.900 28.900 159.900 ;
        RECT 30.600 157.900 31.000 159.900 ;
        RECT 32.800 158.200 33.200 159.900 ;
        RECT 32.800 157.900 33.800 158.200 ;
        RECT 28.600 157.500 29.000 157.900 ;
        RECT 30.700 157.600 31.000 157.900 ;
        RECT 30.300 157.300 32.100 157.600 ;
        RECT 33.400 157.500 33.800 157.900 ;
        RECT 30.300 157.200 30.700 157.300 ;
        RECT 31.700 157.200 32.100 157.300 ;
        RECT 28.200 156.600 28.900 157.000 ;
        RECT 28.600 156.100 28.900 156.600 ;
        RECT 29.700 156.500 30.800 156.800 ;
        RECT 29.700 156.400 30.100 156.500 ;
        RECT 28.600 155.800 29.800 156.100 ;
        RECT 26.200 155.300 28.300 155.600 ;
        RECT 25.400 153.400 25.800 154.200 ;
        RECT 26.200 153.600 26.600 155.300 ;
        RECT 27.900 155.200 28.300 155.300 ;
        RECT 27.100 154.900 27.500 155.000 ;
        RECT 27.100 154.600 29.000 154.900 ;
        RECT 28.600 154.500 29.000 154.600 ;
        RECT 29.500 154.200 29.800 155.800 ;
        RECT 30.500 155.900 30.800 156.500 ;
        RECT 31.100 156.500 31.500 156.600 ;
        RECT 33.400 156.500 33.800 156.600 ;
        RECT 31.100 156.200 33.800 156.500 ;
        RECT 30.500 155.700 32.900 155.900 ;
        RECT 35.000 155.700 35.400 159.900 ;
        RECT 36.100 159.200 36.500 159.900 ;
        RECT 38.500 159.200 38.900 159.900 ;
        RECT 36.100 158.800 37.000 159.200 ;
        RECT 38.500 158.800 39.400 159.200 ;
        RECT 36.100 156.300 36.500 158.800 ;
        RECT 38.500 156.300 38.900 158.800 ;
        RECT 36.100 155.900 37.000 156.300 ;
        RECT 38.500 155.900 39.400 156.300 ;
        RECT 30.500 155.600 35.400 155.700 ;
        RECT 32.500 155.500 35.400 155.600 ;
        RECT 32.600 155.400 35.400 155.500 ;
        RECT 30.200 155.100 30.600 155.200 ;
        RECT 31.800 155.100 32.200 155.200 ;
        RECT 30.200 154.800 34.300 155.100 ;
        RECT 35.800 154.800 36.200 155.600 ;
        RECT 33.900 154.700 34.300 154.800 ;
        RECT 33.100 154.200 33.500 154.300 ;
        RECT 36.600 154.200 36.900 155.900 ;
        RECT 37.400 155.100 37.800 155.200 ;
        RECT 38.200 155.100 38.600 155.600 ;
        RECT 37.400 154.800 38.600 155.100 ;
        RECT 39.000 154.200 39.300 155.900 ;
        RECT 29.500 153.900 35.000 154.200 ;
        RECT 29.700 153.800 30.100 153.900 ;
        RECT 24.100 152.800 25.000 153.100 ;
        RECT 26.200 153.300 28.100 153.600 ;
        RECT 24.100 151.100 24.500 152.800 ;
        RECT 26.200 151.100 26.600 153.300 ;
        RECT 27.700 153.200 28.100 153.300 ;
        RECT 32.600 152.800 32.900 153.900 ;
        RECT 34.200 153.800 35.000 153.900 ;
        RECT 36.600 153.800 37.000 154.200 ;
        RECT 39.000 153.800 39.400 154.200 ;
        RECT 31.700 152.700 32.100 152.800 ;
        RECT 28.600 152.100 29.000 152.500 ;
        RECT 30.700 152.400 32.100 152.700 ;
        RECT 32.600 152.400 33.000 152.800 ;
        RECT 30.700 152.100 31.000 152.400 ;
        RECT 33.400 152.100 33.800 152.500 ;
        RECT 28.300 151.800 29.000 152.100 ;
        RECT 28.300 151.100 28.900 151.800 ;
        RECT 30.600 151.100 31.000 152.100 ;
        RECT 32.800 151.800 33.800 152.100 ;
        RECT 32.800 151.100 33.200 151.800 ;
        RECT 35.000 151.100 35.400 153.500 ;
        RECT 36.600 152.200 36.900 153.800 ;
        RECT 39.000 152.200 39.300 153.800 ;
        RECT 39.800 153.100 40.200 153.200 ;
        RECT 40.600 153.100 41.000 159.900 ;
        RECT 44.100 159.200 44.500 159.900 ;
        RECT 44.100 158.800 45.000 159.200 ;
        RECT 44.100 156.400 44.500 158.800 ;
        RECT 46.200 157.500 46.600 159.500 ;
        RECT 43.700 156.100 44.500 156.400 ;
        RECT 42.200 155.100 42.600 155.200 ;
        RECT 43.000 155.100 43.400 155.600 ;
        RECT 42.200 154.800 43.400 155.100 ;
        RECT 43.700 154.200 44.000 156.100 ;
        RECT 46.300 155.800 46.600 157.500 ;
        RECT 47.300 156.300 47.700 159.900 ;
        RECT 51.300 159.200 51.700 159.900 ;
        RECT 51.300 158.800 52.200 159.200 ;
        RECT 51.300 156.300 51.700 158.800 ;
        RECT 47.300 155.900 48.200 156.300 ;
        RECT 51.300 155.900 52.200 156.300 ;
        RECT 44.700 155.500 46.600 155.800 ;
        RECT 44.700 154.500 45.000 155.500 ;
        RECT 43.000 153.800 44.000 154.200 ;
        RECT 44.300 154.100 45.000 154.500 ;
        RECT 45.400 154.400 45.800 155.200 ;
        RECT 46.200 154.400 46.600 155.200 ;
        RECT 47.000 154.800 47.400 155.600 ;
        RECT 39.800 152.800 41.000 153.100 ;
        RECT 43.700 153.500 44.000 153.800 ;
        RECT 44.500 153.900 45.000 154.100 ;
        RECT 47.800 154.200 48.100 155.900 ;
        RECT 49.400 155.100 49.800 155.200 ;
        RECT 51.000 155.100 51.400 155.600 ;
        RECT 49.400 154.800 51.400 155.100 ;
        RECT 51.800 154.200 52.100 155.900 ;
        RECT 53.400 155.600 53.800 159.900 ;
        RECT 55.500 157.900 56.100 159.900 ;
        RECT 57.800 157.900 58.200 159.900 ;
        RECT 60.000 158.200 60.400 159.900 ;
        RECT 60.000 157.900 61.000 158.200 ;
        RECT 55.800 157.500 56.200 157.900 ;
        RECT 57.900 157.600 58.200 157.900 ;
        RECT 57.500 157.300 59.300 157.600 ;
        RECT 60.600 157.500 61.000 157.900 ;
        RECT 57.500 157.200 57.900 157.300 ;
        RECT 58.900 157.200 59.300 157.300 ;
        RECT 55.400 156.600 56.100 157.000 ;
        RECT 55.800 156.100 56.100 156.600 ;
        RECT 56.900 156.500 58.000 156.800 ;
        RECT 56.900 156.400 57.300 156.500 ;
        RECT 55.800 155.800 57.000 156.100 ;
        RECT 53.400 155.300 55.500 155.600 ;
        RECT 47.800 154.100 48.200 154.200 ;
        RECT 51.000 154.100 51.400 154.200 ;
        RECT 44.500 153.600 46.600 153.900 ;
        RECT 43.700 153.300 44.100 153.500 ;
        RECT 43.700 153.000 44.500 153.300 ;
        RECT 39.800 152.400 40.200 152.800 ;
        RECT 36.600 151.100 37.000 152.200 ;
        RECT 39.000 151.100 39.400 152.200 ;
        RECT 40.600 151.100 41.000 152.800 ;
        RECT 44.100 151.500 44.500 153.000 ;
        RECT 46.300 152.500 46.600 153.600 ;
        RECT 46.200 151.500 46.600 152.500 ;
        RECT 47.800 153.800 51.400 154.100 ;
        RECT 51.800 153.800 52.200 154.200 ;
        RECT 47.800 152.100 48.100 153.800 ;
        RECT 48.600 152.400 49.000 153.200 ;
        RECT 51.800 152.100 52.100 153.800 ;
        RECT 53.400 153.600 53.800 155.300 ;
        RECT 55.100 155.200 55.500 155.300 ;
        RECT 56.700 155.200 57.000 155.800 ;
        RECT 57.700 155.900 58.000 156.500 ;
        RECT 58.300 156.500 58.700 156.600 ;
        RECT 60.600 156.500 61.000 156.600 ;
        RECT 58.300 156.200 61.000 156.500 ;
        RECT 57.700 155.700 60.100 155.900 ;
        RECT 62.200 155.700 62.600 159.900 ;
        RECT 57.700 155.600 62.600 155.700 ;
        RECT 59.700 155.500 62.600 155.600 ;
        RECT 59.800 155.400 62.600 155.500 ;
        RECT 54.300 154.900 54.700 155.000 ;
        RECT 54.300 154.600 56.200 154.900 ;
        RECT 56.600 154.800 57.000 155.200 ;
        RECT 59.000 155.100 59.400 155.200 ;
        RECT 63.800 155.100 64.200 159.900 ;
        RECT 65.800 156.800 66.200 157.200 ;
        RECT 64.600 155.800 65.000 156.600 ;
        RECT 65.800 156.200 66.100 156.800 ;
        RECT 66.500 156.200 66.900 159.900 ;
        RECT 65.400 155.900 66.100 156.200 ;
        RECT 66.400 155.900 66.900 156.200 ;
        RECT 65.400 155.800 65.800 155.900 ;
        RECT 65.400 155.100 65.700 155.800 ;
        RECT 66.400 155.200 66.700 155.900 ;
        RECT 69.400 155.600 69.800 159.900 ;
        RECT 71.000 155.600 71.400 159.900 ;
        RECT 72.600 155.600 73.000 159.900 ;
        RECT 74.200 155.600 74.600 159.900 ;
        RECT 77.100 156.200 77.500 159.900 ;
        RECT 77.800 156.800 78.200 157.200 ;
        RECT 77.900 156.200 78.200 156.800 ;
        RECT 77.100 155.900 77.600 156.200 ;
        RECT 77.900 156.100 78.600 156.200 ;
        RECT 79.800 156.100 80.200 159.900 ;
        RECT 77.900 155.900 80.200 156.100 ;
        RECT 69.400 155.200 70.300 155.600 ;
        RECT 71.000 155.200 72.100 155.600 ;
        RECT 72.600 155.200 73.700 155.600 ;
        RECT 74.200 155.200 75.400 155.600 ;
        RECT 59.000 154.800 61.500 155.100 ;
        RECT 55.800 154.500 56.200 154.600 ;
        RECT 56.700 154.200 57.000 154.800 ;
        RECT 59.800 154.700 60.200 154.800 ;
        RECT 61.100 154.700 61.500 154.800 ;
        RECT 63.800 154.800 65.700 155.100 ;
        RECT 66.200 154.800 66.700 155.200 ;
        RECT 60.300 154.200 60.700 154.300 ;
        RECT 55.000 153.600 55.400 154.200 ;
        RECT 56.700 153.900 62.200 154.200 ;
        RECT 56.900 153.800 57.300 153.900 ;
        RECT 53.400 153.300 55.400 153.600 ;
        RECT 47.800 151.100 48.200 152.100 ;
        RECT 51.800 151.100 52.200 152.100 ;
        RECT 53.400 151.100 53.800 153.300 ;
        RECT 54.900 153.200 55.300 153.300 ;
        RECT 59.800 152.800 60.100 153.900 ;
        RECT 61.400 153.800 62.200 153.900 ;
        RECT 58.900 152.700 59.300 152.800 ;
        RECT 55.800 152.100 56.200 152.500 ;
        RECT 57.900 152.400 59.300 152.700 ;
        RECT 59.800 152.400 60.200 152.800 ;
        RECT 57.900 152.100 58.200 152.400 ;
        RECT 60.600 152.100 61.000 152.500 ;
        RECT 55.500 151.800 56.200 152.100 ;
        RECT 55.500 151.100 56.100 151.800 ;
        RECT 57.800 151.100 58.200 152.100 ;
        RECT 60.000 151.800 61.000 152.100 ;
        RECT 60.000 151.100 60.400 151.800 ;
        RECT 62.200 151.100 62.600 153.500 ;
        RECT 63.000 153.400 63.400 154.200 ;
        RECT 63.800 153.100 64.200 154.800 ;
        RECT 66.400 154.200 66.700 154.800 ;
        RECT 67.000 154.400 67.400 155.200 ;
        RECT 69.900 154.500 70.300 155.200 ;
        RECT 71.700 154.500 72.100 155.200 ;
        RECT 73.300 154.500 73.700 155.200 ;
        RECT 65.400 153.800 66.700 154.200 ;
        RECT 67.800 154.100 68.200 154.200 ;
        RECT 67.400 153.800 68.200 154.100 ;
        RECT 68.600 154.100 69.500 154.500 ;
        RECT 69.900 154.100 71.200 154.500 ;
        RECT 71.700 154.100 72.900 154.500 ;
        RECT 73.300 154.100 74.600 154.500 ;
        RECT 68.600 153.800 69.000 154.100 ;
        RECT 69.900 153.800 70.300 154.100 ;
        RECT 71.700 153.800 72.100 154.100 ;
        RECT 73.300 153.800 73.700 154.100 ;
        RECT 75.000 153.800 75.400 155.200 ;
        RECT 76.600 154.400 77.000 155.200 ;
        RECT 77.300 155.100 77.600 155.900 ;
        RECT 78.200 155.800 80.200 155.900 ;
        RECT 80.600 155.800 81.000 156.600 ;
        RECT 78.200 155.100 78.600 155.200 ;
        RECT 77.300 154.800 78.600 155.100 ;
        RECT 77.300 154.200 77.600 154.800 ;
        RECT 75.800 154.100 76.200 154.200 ;
        RECT 75.800 153.800 76.600 154.100 ;
        RECT 77.300 153.800 78.600 154.200 ;
        RECT 65.500 153.100 65.800 153.800 ;
        RECT 67.400 153.600 67.800 153.800 ;
        RECT 69.400 153.400 70.300 153.800 ;
        RECT 71.000 153.400 72.100 153.800 ;
        RECT 72.600 153.400 73.700 153.800 ;
        RECT 74.200 153.400 75.400 153.800 ;
        RECT 76.200 153.600 76.600 153.800 ;
        RECT 66.300 153.100 68.100 153.300 ;
        RECT 63.800 152.800 64.700 153.100 ;
        RECT 64.300 151.100 64.700 152.800 ;
        RECT 65.400 151.100 65.800 153.100 ;
        RECT 66.200 153.000 68.200 153.100 ;
        RECT 66.200 151.100 66.600 153.000 ;
        RECT 67.800 151.100 68.200 153.000 ;
        RECT 69.400 151.100 69.800 153.400 ;
        RECT 71.000 151.100 71.400 153.400 ;
        RECT 72.600 151.100 73.000 153.400 ;
        RECT 74.200 151.100 74.600 153.400 ;
        RECT 75.900 153.100 77.700 153.300 ;
        RECT 78.200 153.100 78.500 153.800 ;
        RECT 79.000 153.400 79.400 154.200 ;
        RECT 79.800 153.100 80.200 155.800 ;
        RECT 81.400 155.600 81.800 159.900 ;
        RECT 83.500 157.900 84.100 159.900 ;
        RECT 85.800 157.900 86.200 159.900 ;
        RECT 88.000 158.200 88.400 159.900 ;
        RECT 88.000 157.900 89.000 158.200 ;
        RECT 83.800 157.500 84.200 157.900 ;
        RECT 85.900 157.600 86.200 157.900 ;
        RECT 85.500 157.300 87.300 157.600 ;
        RECT 88.600 157.500 89.000 157.900 ;
        RECT 85.500 157.200 85.900 157.300 ;
        RECT 86.900 157.200 87.300 157.300 ;
        RECT 83.400 156.600 84.100 157.000 ;
        RECT 83.800 156.100 84.100 156.600 ;
        RECT 84.900 156.500 86.000 156.800 ;
        RECT 84.900 156.400 85.300 156.500 ;
        RECT 83.800 155.800 85.000 156.100 ;
        RECT 81.400 155.300 83.500 155.600 ;
        RECT 81.400 153.600 81.800 155.300 ;
        RECT 83.100 155.200 83.500 155.300 ;
        RECT 84.700 155.200 85.000 155.800 ;
        RECT 85.700 155.900 86.000 156.500 ;
        RECT 86.300 156.500 86.700 156.600 ;
        RECT 88.600 156.500 89.000 156.600 ;
        RECT 86.300 156.200 89.000 156.500 ;
        RECT 85.700 155.700 88.100 155.900 ;
        RECT 90.200 155.700 90.600 159.900 ;
        RECT 91.000 156.200 91.400 159.900 ;
        RECT 93.400 156.200 93.800 159.900 ;
        RECT 95.000 156.200 95.400 159.900 ;
        RECT 91.000 155.900 92.100 156.200 ;
        RECT 93.400 155.900 95.400 156.200 ;
        RECT 95.800 155.900 96.200 159.900 ;
        RECT 96.900 156.300 97.300 159.900 ;
        RECT 96.900 155.900 97.800 156.300 ;
        RECT 100.600 156.200 101.000 159.900 ;
        RECT 102.200 156.200 102.600 159.900 ;
        RECT 100.600 155.900 102.600 156.200 ;
        RECT 103.000 155.900 103.400 159.900 ;
        RECT 104.100 156.300 104.500 159.900 ;
        RECT 104.100 155.900 105.000 156.300 ;
        RECT 106.200 156.200 106.600 159.900 ;
        RECT 107.800 156.200 108.200 159.900 ;
        RECT 106.200 155.900 108.200 156.200 ;
        RECT 108.600 155.900 109.000 159.900 ;
        RECT 109.700 156.300 110.100 159.900 ;
        RECT 109.700 155.900 110.600 156.300 ;
        RECT 85.700 155.600 90.600 155.700 ;
        RECT 87.700 155.500 90.600 155.600 ;
        RECT 87.800 155.400 90.600 155.500 ;
        RECT 91.800 155.600 92.100 155.900 ;
        RECT 91.800 155.200 92.400 155.600 ;
        RECT 93.800 155.200 94.200 155.400 ;
        RECT 95.800 155.200 96.100 155.900 ;
        RECT 82.300 154.900 82.700 155.000 ;
        RECT 82.300 154.600 84.200 154.900 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 87.000 155.100 87.400 155.200 ;
        RECT 87.000 154.800 89.500 155.100 ;
        RECT 83.800 154.500 84.200 154.600 ;
        RECT 84.700 154.200 85.000 154.800 ;
        RECT 89.100 154.700 89.500 154.800 ;
        RECT 91.000 154.400 91.400 155.200 ;
        RECT 88.300 154.200 88.700 154.300 ;
        RECT 84.700 153.900 90.200 154.200 ;
        RECT 84.900 153.800 85.300 153.900 ;
        RECT 81.400 153.300 83.300 153.600 ;
        RECT 75.800 153.000 77.800 153.100 ;
        RECT 75.800 151.100 76.200 153.000 ;
        RECT 77.400 151.100 77.800 153.000 ;
        RECT 78.200 151.100 78.600 153.100 ;
        RECT 79.800 152.800 80.700 153.100 ;
        RECT 80.300 151.100 80.700 152.800 ;
        RECT 81.400 151.100 81.800 153.300 ;
        RECT 82.900 153.200 83.300 153.300 ;
        RECT 87.800 152.800 88.100 153.900 ;
        RECT 89.400 153.800 90.200 153.900 ;
        RECT 91.800 153.700 92.100 155.200 ;
        RECT 93.400 154.900 94.200 155.200 ;
        RECT 95.000 154.900 96.200 155.200 ;
        RECT 93.400 154.800 93.800 154.900 ;
        RECT 94.200 153.800 94.600 154.600 ;
        RECT 86.900 152.700 87.300 152.800 ;
        RECT 83.800 152.100 84.200 152.500 ;
        RECT 85.900 152.400 87.300 152.700 ;
        RECT 87.800 152.400 88.200 152.800 ;
        RECT 85.900 152.100 86.200 152.400 ;
        RECT 88.600 152.100 89.000 152.500 ;
        RECT 83.500 151.800 84.200 152.100 ;
        RECT 83.500 151.100 84.100 151.800 ;
        RECT 85.800 151.100 86.200 152.100 ;
        RECT 88.000 151.800 89.000 152.100 ;
        RECT 88.000 151.100 88.400 151.800 ;
        RECT 90.200 151.100 90.600 153.500 ;
        RECT 91.000 153.400 92.100 153.700 ;
        RECT 91.000 151.100 91.400 153.400 ;
        RECT 95.000 153.100 95.300 154.900 ;
        RECT 95.800 154.800 96.200 154.900 ;
        RECT 96.600 154.800 97.000 155.600 ;
        RECT 97.400 154.200 97.700 155.900 ;
        RECT 101.000 155.200 101.400 155.400 ;
        RECT 103.000 155.200 103.300 155.900 ;
        RECT 100.600 154.900 101.400 155.200 ;
        RECT 102.200 154.900 103.400 155.200 ;
        RECT 100.600 154.800 101.000 154.900 ;
        RECT 97.400 153.800 97.800 154.200 ;
        RECT 101.400 153.800 101.800 154.600 ;
        RECT 95.800 153.100 96.200 153.200 ;
        RECT 97.400 153.100 97.700 153.800 ;
        RECT 95.000 151.100 95.400 153.100 ;
        RECT 95.800 152.800 97.700 153.100 ;
        RECT 95.700 152.400 96.100 152.800 ;
        RECT 97.400 152.100 97.700 152.800 ;
        RECT 98.200 153.100 98.600 153.200 ;
        RECT 99.800 153.100 100.200 153.200 ;
        RECT 98.200 152.800 100.200 153.100 ;
        RECT 102.200 153.100 102.500 154.900 ;
        RECT 103.000 154.800 103.400 154.900 ;
        RECT 103.800 154.800 104.200 155.600 ;
        RECT 104.600 154.200 104.900 155.900 ;
        RECT 106.600 155.200 107.000 155.400 ;
        RECT 108.600 155.200 108.900 155.900 ;
        RECT 106.200 154.900 107.000 155.200 ;
        RECT 107.800 154.900 109.000 155.200 ;
        RECT 106.200 154.800 106.600 154.900 ;
        RECT 104.600 153.800 105.000 154.200 ;
        RECT 107.000 153.800 107.400 154.600 ;
        RECT 103.000 153.100 103.400 153.200 ;
        RECT 104.600 153.100 104.900 153.800 ;
        RECT 98.200 152.400 98.600 152.800 ;
        RECT 97.400 151.100 97.800 152.100 ;
        RECT 102.200 151.100 102.600 153.100 ;
        RECT 103.000 152.800 104.900 153.100 ;
        RECT 102.900 152.400 103.300 152.800 ;
        RECT 104.600 152.100 104.900 152.800 ;
        RECT 105.400 152.400 105.800 153.200 ;
        RECT 107.800 153.100 108.100 154.900 ;
        RECT 108.600 154.800 109.000 154.900 ;
        RECT 109.400 154.800 109.800 155.600 ;
        RECT 110.200 154.200 110.500 155.900 ;
        RECT 110.200 153.800 110.600 154.200 ;
        RECT 108.600 153.100 109.000 153.200 ;
        RECT 110.200 153.100 110.500 153.800 ;
        RECT 104.600 151.100 105.000 152.100 ;
        RECT 107.800 151.100 108.200 153.100 ;
        RECT 108.600 152.800 110.500 153.100 ;
        RECT 108.500 152.400 108.900 152.800 ;
        RECT 110.200 152.100 110.500 152.800 ;
        RECT 111.000 152.400 111.400 153.200 ;
        RECT 110.200 151.100 110.600 152.100 ;
        RECT 112.600 151.100 113.000 159.900 ;
        RECT 114.200 155.700 114.600 159.900 ;
        RECT 116.400 158.200 116.800 159.900 ;
        RECT 115.800 157.900 116.800 158.200 ;
        RECT 118.600 157.900 119.000 159.900 ;
        RECT 120.700 157.900 121.300 159.900 ;
        RECT 115.800 157.500 116.200 157.900 ;
        RECT 118.600 157.600 118.900 157.900 ;
        RECT 117.500 157.300 119.300 157.600 ;
        RECT 120.600 157.500 121.000 157.900 ;
        RECT 117.500 157.200 117.900 157.300 ;
        RECT 118.900 157.200 119.300 157.300 ;
        RECT 123.000 157.100 123.400 159.900 ;
        RECT 123.800 157.100 124.200 157.200 ;
        RECT 115.800 156.500 116.200 156.600 ;
        RECT 118.100 156.500 118.500 156.600 ;
        RECT 115.800 156.200 118.500 156.500 ;
        RECT 118.800 156.500 119.900 156.800 ;
        RECT 118.800 155.900 119.100 156.500 ;
        RECT 119.500 156.400 119.900 156.500 ;
        RECT 120.700 156.600 121.400 157.000 ;
        RECT 123.000 156.800 124.200 157.100 ;
        RECT 120.700 156.100 121.000 156.600 ;
        RECT 116.700 155.700 119.100 155.900 ;
        RECT 114.200 155.600 119.100 155.700 ;
        RECT 119.800 155.800 121.000 156.100 ;
        RECT 114.200 155.500 117.100 155.600 ;
        RECT 114.200 155.400 117.000 155.500 ;
        RECT 117.400 155.100 117.800 155.200 ;
        RECT 115.300 154.800 117.800 155.100 ;
        RECT 115.300 154.700 115.700 154.800 ;
        RECT 116.100 154.200 116.500 154.300 ;
        RECT 119.800 154.200 120.100 155.800 ;
        RECT 123.000 155.600 123.400 156.800 ;
        RECT 121.300 155.300 123.400 155.600 ;
        RECT 121.300 155.200 121.700 155.300 ;
        RECT 122.100 154.900 122.500 155.000 ;
        RECT 120.600 154.600 122.500 154.900 ;
        RECT 120.600 154.500 121.000 154.600 ;
        RECT 114.600 153.900 120.100 154.200 ;
        RECT 114.600 153.800 115.400 153.900 ;
        RECT 114.200 151.100 114.600 153.500 ;
        RECT 116.700 152.800 117.000 153.900 ;
        RECT 119.500 153.800 119.900 153.900 ;
        RECT 123.000 153.600 123.400 155.300 ;
        RECT 124.600 155.100 125.000 159.900 ;
        RECT 126.600 156.800 127.000 157.200 ;
        RECT 125.400 155.800 125.800 156.600 ;
        RECT 126.600 156.200 126.900 156.800 ;
        RECT 127.300 156.200 127.700 159.900 ;
        RECT 126.200 155.900 126.900 156.200 ;
        RECT 127.200 155.900 127.700 156.200 ;
        RECT 129.400 157.500 129.800 159.500 ;
        RECT 131.500 159.200 131.900 159.900 ;
        RECT 131.000 158.800 131.900 159.200 ;
        RECT 126.200 155.800 126.600 155.900 ;
        RECT 126.200 155.100 126.500 155.800 ;
        RECT 124.600 154.800 126.500 155.100 ;
        RECT 121.500 153.300 123.400 153.600 ;
        RECT 123.800 153.400 124.200 154.200 ;
        RECT 121.500 153.200 121.900 153.300 ;
        RECT 115.800 152.100 116.200 152.500 ;
        RECT 116.600 152.400 117.000 152.800 ;
        RECT 117.500 152.700 117.900 152.800 ;
        RECT 117.500 152.400 118.900 152.700 ;
        RECT 118.600 152.100 118.900 152.400 ;
        RECT 120.600 152.100 121.000 152.500 ;
        RECT 115.800 151.800 116.800 152.100 ;
        RECT 116.400 151.100 116.800 151.800 ;
        RECT 118.600 151.100 119.000 152.100 ;
        RECT 120.600 151.800 121.300 152.100 ;
        RECT 120.700 151.100 121.300 151.800 ;
        RECT 123.000 151.100 123.400 153.300 ;
        RECT 124.600 153.100 125.000 154.800 ;
        RECT 127.200 154.200 127.500 155.900 ;
        RECT 129.400 155.800 129.700 157.500 ;
        RECT 131.500 156.400 131.900 158.800 ;
        RECT 131.500 156.100 132.300 156.400 ;
        RECT 129.400 155.500 131.300 155.800 ;
        RECT 127.800 154.400 128.200 155.200 ;
        RECT 129.400 154.400 129.800 155.200 ;
        RECT 130.200 154.400 130.600 155.200 ;
        RECT 131.000 154.500 131.300 155.500 ;
        RECT 125.400 154.100 125.800 154.200 ;
        RECT 126.200 154.100 127.500 154.200 ;
        RECT 128.600 154.100 129.000 154.200 ;
        RECT 125.400 153.800 127.500 154.100 ;
        RECT 128.200 153.800 129.000 154.100 ;
        RECT 131.000 154.100 131.700 154.500 ;
        RECT 132.000 154.200 132.300 156.100 ;
        RECT 134.200 155.700 134.600 159.900 ;
        RECT 136.400 158.200 136.800 159.900 ;
        RECT 135.800 157.900 136.800 158.200 ;
        RECT 138.600 157.900 139.000 159.900 ;
        RECT 140.700 157.900 141.300 159.900 ;
        RECT 135.800 157.500 136.200 157.900 ;
        RECT 138.600 157.600 138.900 157.900 ;
        RECT 137.500 157.300 139.300 157.600 ;
        RECT 140.600 157.500 141.000 157.900 ;
        RECT 137.500 157.200 137.900 157.300 ;
        RECT 138.900 157.200 139.300 157.300 ;
        RECT 135.800 156.500 136.200 156.600 ;
        RECT 138.100 156.500 138.500 156.600 ;
        RECT 135.800 156.200 138.500 156.500 ;
        RECT 138.800 156.500 139.900 156.800 ;
        RECT 138.800 155.900 139.100 156.500 ;
        RECT 139.500 156.400 139.900 156.500 ;
        RECT 140.700 156.600 141.400 157.000 ;
        RECT 140.700 156.100 141.000 156.600 ;
        RECT 136.700 155.700 139.100 155.900 ;
        RECT 134.200 155.600 139.100 155.700 ;
        RECT 139.800 155.800 141.000 156.100 ;
        RECT 132.600 154.800 133.000 155.600 ;
        RECT 134.200 155.500 137.100 155.600 ;
        RECT 134.200 155.400 137.000 155.500 ;
        RECT 139.800 155.200 140.100 155.800 ;
        RECT 143.000 155.600 143.400 159.900 ;
        RECT 143.800 155.800 144.200 156.600 ;
        RECT 141.300 155.300 143.400 155.600 ;
        RECT 141.300 155.200 141.700 155.300 ;
        RECT 137.400 155.100 137.800 155.200 ;
        RECT 138.200 155.100 138.600 155.200 ;
        RECT 135.300 154.800 138.600 155.100 ;
        RECT 139.800 154.800 140.200 155.200 ;
        RECT 142.100 154.900 142.500 155.000 ;
        RECT 135.300 154.700 135.700 154.800 ;
        RECT 136.100 154.200 136.500 154.300 ;
        RECT 139.800 154.200 140.100 154.800 ;
        RECT 140.600 154.600 142.500 154.900 ;
        RECT 140.600 154.500 141.000 154.600 ;
        RECT 131.000 153.900 131.500 154.100 ;
        RECT 126.300 153.100 126.600 153.800 ;
        RECT 128.200 153.600 128.600 153.800 ;
        RECT 129.400 153.600 131.500 153.900 ;
        RECT 132.000 153.800 133.000 154.200 ;
        RECT 134.600 153.900 140.100 154.200 ;
        RECT 134.600 153.800 135.400 153.900 ;
        RECT 127.100 153.100 128.900 153.300 ;
        RECT 124.600 152.800 125.500 153.100 ;
        RECT 125.100 151.100 125.500 152.800 ;
        RECT 126.200 151.100 126.600 153.100 ;
        RECT 127.000 153.000 129.000 153.100 ;
        RECT 127.000 151.100 127.400 153.000 ;
        RECT 128.600 151.100 129.000 153.000 ;
        RECT 129.400 152.500 129.700 153.600 ;
        RECT 132.000 153.500 132.300 153.800 ;
        RECT 131.900 153.300 132.300 153.500 ;
        RECT 131.500 153.000 132.300 153.300 ;
        RECT 129.400 151.500 129.800 152.500 ;
        RECT 131.500 151.500 131.900 153.000 ;
        RECT 134.200 151.100 134.600 153.500 ;
        RECT 136.700 152.800 137.000 153.900 ;
        RECT 137.400 153.800 137.800 153.900 ;
        RECT 139.500 153.800 139.900 153.900 ;
        RECT 143.000 153.600 143.400 155.300 ;
        RECT 141.500 153.300 143.400 153.600 ;
        RECT 141.500 153.200 141.900 153.300 ;
        RECT 135.800 152.100 136.200 152.500 ;
        RECT 136.600 152.400 137.000 152.800 ;
        RECT 137.500 152.700 137.900 152.800 ;
        RECT 137.500 152.400 138.900 152.700 ;
        RECT 138.600 152.100 138.900 152.400 ;
        RECT 140.600 152.100 141.000 152.500 ;
        RECT 135.800 151.800 136.800 152.100 ;
        RECT 136.400 151.100 136.800 151.800 ;
        RECT 138.600 151.100 139.000 152.100 ;
        RECT 140.600 151.800 141.300 152.100 ;
        RECT 140.700 151.100 141.300 151.800 ;
        RECT 143.000 151.100 143.400 153.300 ;
        RECT 144.600 153.100 145.000 159.900 ;
        RECT 145.400 153.400 145.800 154.200 ;
        RECT 146.200 153.400 146.600 154.200 ;
        RECT 144.100 152.800 145.000 153.100 ;
        RECT 147.000 153.100 147.400 159.900 ;
        RECT 152.100 159.200 152.500 159.900 ;
        RECT 152.100 158.800 153.000 159.200 ;
        RECT 147.800 155.800 148.200 156.600 ;
        RECT 152.100 156.400 152.500 158.800 ;
        RECT 154.200 157.500 154.600 159.500 ;
        RECT 151.700 156.100 152.500 156.400 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 151.000 155.100 151.400 155.600 ;
        RECT 147.800 154.800 151.400 155.100 ;
        RECT 151.700 154.200 152.000 156.100 ;
        RECT 154.300 155.800 154.600 157.500 ;
        RECT 156.300 156.200 156.700 159.900 ;
        RECT 157.000 156.800 157.400 157.200 ;
        RECT 157.100 156.200 157.400 156.800 ;
        RECT 156.300 155.900 156.800 156.200 ;
        RECT 157.100 155.900 157.800 156.200 ;
        RECT 152.700 155.500 154.600 155.800 ;
        RECT 152.700 154.500 153.000 155.500 ;
        RECT 151.000 153.800 152.000 154.200 ;
        RECT 152.300 154.100 153.000 154.500 ;
        RECT 153.400 154.400 153.800 155.200 ;
        RECT 154.200 154.400 154.600 155.200 ;
        RECT 155.800 154.400 156.200 155.200 ;
        RECT 156.500 154.200 156.800 155.900 ;
        RECT 157.400 155.800 157.800 155.900 ;
        RECT 158.200 155.800 158.600 156.600 ;
        RECT 157.400 155.100 157.700 155.800 ;
        RECT 159.000 155.100 159.400 159.900 ;
        RECT 159.800 157.100 160.200 157.200 ;
        RECT 160.600 157.100 161.000 159.900 ;
        RECT 162.700 157.900 163.300 159.900 ;
        RECT 165.000 157.900 165.400 159.900 ;
        RECT 167.200 158.200 167.600 159.900 ;
        RECT 167.200 157.900 168.200 158.200 ;
        RECT 163.000 157.500 163.400 157.900 ;
        RECT 165.100 157.600 165.400 157.900 ;
        RECT 164.700 157.300 166.500 157.600 ;
        RECT 167.800 157.500 168.200 157.900 ;
        RECT 164.700 157.200 165.100 157.300 ;
        RECT 166.100 157.200 166.500 157.300 ;
        RECT 159.800 156.800 161.000 157.100 ;
        RECT 157.400 154.800 159.400 155.100 ;
        RECT 151.700 153.500 152.000 153.800 ;
        RECT 152.500 153.900 153.000 154.100 ;
        RECT 155.000 154.100 155.400 154.200 ;
        RECT 156.500 154.100 157.800 154.200 ;
        RECT 158.200 154.100 158.600 154.200 ;
        RECT 152.500 153.600 154.600 153.900 ;
        RECT 155.000 153.800 155.800 154.100 ;
        RECT 156.500 153.800 158.600 154.100 ;
        RECT 155.400 153.600 155.800 153.800 ;
        RECT 151.700 153.300 152.100 153.500 ;
        RECT 147.000 152.800 147.900 153.100 ;
        RECT 151.700 153.000 152.500 153.300 ;
        RECT 144.100 151.100 144.500 152.800 ;
        RECT 147.500 152.200 147.900 152.800 ;
        RECT 147.500 151.800 148.200 152.200 ;
        RECT 147.500 151.100 147.900 151.800 ;
        RECT 152.100 151.500 152.500 153.000 ;
        RECT 154.300 152.500 154.600 153.600 ;
        RECT 155.100 153.100 156.900 153.300 ;
        RECT 157.400 153.100 157.700 153.800 ;
        RECT 159.000 153.100 159.400 154.800 ;
        RECT 160.600 155.600 161.000 156.800 ;
        RECT 162.600 156.600 163.300 157.000 ;
        RECT 163.000 156.100 163.300 156.600 ;
        RECT 164.100 156.500 165.200 156.800 ;
        RECT 164.100 156.400 164.500 156.500 ;
        RECT 163.000 155.800 164.200 156.100 ;
        RECT 160.600 155.300 162.700 155.600 ;
        RECT 159.800 153.400 160.200 154.200 ;
        RECT 160.600 153.600 161.000 155.300 ;
        RECT 162.300 155.200 162.700 155.300 ;
        RECT 161.500 154.900 161.900 155.000 ;
        RECT 161.500 154.600 163.400 154.900 ;
        RECT 163.000 154.500 163.400 154.600 ;
        RECT 163.900 154.200 164.200 155.800 ;
        RECT 164.900 155.900 165.200 156.500 ;
        RECT 165.500 156.500 165.900 156.600 ;
        RECT 167.800 156.500 168.200 156.600 ;
        RECT 165.500 156.200 168.200 156.500 ;
        RECT 164.900 155.700 167.300 155.900 ;
        RECT 169.400 155.700 169.800 159.900 ;
        RECT 164.900 155.600 169.800 155.700 ;
        RECT 166.900 155.500 169.800 155.600 ;
        RECT 167.000 155.400 169.800 155.500 ;
        RECT 166.200 155.100 166.600 155.200 ;
        RECT 166.200 154.800 168.700 155.100 ;
        RECT 168.300 154.700 168.700 154.800 ;
        RECT 167.500 154.200 167.900 154.300 ;
        RECT 163.900 153.900 169.400 154.200 ;
        RECT 164.100 153.800 164.500 153.900 ;
        RECT 154.200 151.500 154.600 152.500 ;
        RECT 155.000 153.000 157.000 153.100 ;
        RECT 155.000 151.100 155.400 153.000 ;
        RECT 156.600 151.100 157.000 153.000 ;
        RECT 157.400 151.100 157.800 153.100 ;
        RECT 158.500 152.800 159.400 153.100 ;
        RECT 160.600 153.300 162.500 153.600 ;
        RECT 158.500 151.100 158.900 152.800 ;
        RECT 160.600 151.100 161.000 153.300 ;
        RECT 162.100 153.200 162.500 153.300 ;
        RECT 167.000 152.800 167.300 153.900 ;
        RECT 168.600 153.800 169.400 153.900 ;
        RECT 166.100 152.700 166.500 152.800 ;
        RECT 163.000 152.100 163.400 152.500 ;
        RECT 165.100 152.400 166.500 152.700 ;
        RECT 167.000 152.400 167.400 152.800 ;
        RECT 165.100 152.100 165.400 152.400 ;
        RECT 167.800 152.100 168.200 152.500 ;
        RECT 162.700 151.800 163.400 152.100 ;
        RECT 162.700 151.100 163.300 151.800 ;
        RECT 165.000 151.100 165.400 152.100 ;
        RECT 167.200 151.800 168.200 152.100 ;
        RECT 167.200 151.100 167.600 151.800 ;
        RECT 169.400 151.100 169.800 153.500 ;
        RECT 170.200 153.400 170.600 154.200 ;
        RECT 171.000 153.100 171.400 159.900 ;
        RECT 171.800 155.800 172.200 156.600 ;
        RECT 173.900 156.200 174.300 159.900 ;
        RECT 174.600 156.800 175.000 157.200 ;
        RECT 174.700 156.200 175.000 156.800 ;
        RECT 173.900 155.900 174.400 156.200 ;
        RECT 174.700 155.900 175.400 156.200 ;
        RECT 173.400 154.400 173.800 155.200 ;
        RECT 174.100 154.200 174.400 155.900 ;
        RECT 175.000 155.800 175.400 155.900 ;
        RECT 175.800 155.800 176.200 156.600 ;
        RECT 175.000 155.100 175.300 155.800 ;
        RECT 176.600 155.100 177.000 159.900 ;
        RECT 178.200 157.500 178.600 159.500 ;
        RECT 180.300 159.200 180.700 159.900 ;
        RECT 179.800 158.800 180.700 159.200 ;
        RECT 178.200 155.800 178.500 157.500 ;
        RECT 180.300 156.400 180.700 158.800 ;
        RECT 180.300 156.100 181.100 156.400 ;
        RECT 178.200 155.500 180.100 155.800 ;
        RECT 175.000 154.800 177.000 155.100 ;
        RECT 172.600 154.100 173.000 154.200 ;
        RECT 172.600 153.800 173.400 154.100 ;
        RECT 174.100 153.800 175.400 154.200 ;
        RECT 173.000 153.600 173.400 153.800 ;
        RECT 172.700 153.100 174.500 153.300 ;
        RECT 175.000 153.100 175.300 153.800 ;
        RECT 176.600 153.100 177.000 154.800 ;
        RECT 178.200 154.400 178.600 155.200 ;
        RECT 179.000 154.400 179.400 155.200 ;
        RECT 179.800 154.500 180.100 155.500 ;
        RECT 177.400 153.400 177.800 154.200 ;
        RECT 179.800 154.100 180.500 154.500 ;
        RECT 180.800 154.200 181.100 156.100 ;
        RECT 183.000 155.600 183.400 159.900 ;
        RECT 185.100 157.900 185.700 159.900 ;
        RECT 187.400 157.900 187.800 159.900 ;
        RECT 189.600 158.200 190.000 159.900 ;
        RECT 189.600 157.900 190.600 158.200 ;
        RECT 185.400 157.500 185.800 157.900 ;
        RECT 187.500 157.600 187.800 157.900 ;
        RECT 187.100 157.300 188.900 157.600 ;
        RECT 190.200 157.500 190.600 157.900 ;
        RECT 187.100 157.200 187.500 157.300 ;
        RECT 188.500 157.200 188.900 157.300 ;
        RECT 185.000 156.600 185.700 157.000 ;
        RECT 185.400 156.100 185.700 156.600 ;
        RECT 186.500 156.500 187.600 156.800 ;
        RECT 186.500 156.400 186.900 156.500 ;
        RECT 185.400 155.800 186.600 156.100 ;
        RECT 181.400 155.100 181.800 155.600 ;
        RECT 183.000 155.300 185.100 155.600 ;
        RECT 182.200 155.100 182.600 155.200 ;
        RECT 181.400 154.800 182.600 155.100 ;
        RECT 179.800 153.900 180.300 154.100 ;
        RECT 178.200 153.600 180.300 153.900 ;
        RECT 180.800 153.800 181.800 154.200 ;
        RECT 171.000 152.800 171.900 153.100 ;
        RECT 171.500 152.200 171.900 152.800 ;
        RECT 172.600 153.000 174.600 153.100 ;
        RECT 171.500 151.800 172.200 152.200 ;
        RECT 171.500 151.100 171.900 151.800 ;
        RECT 172.600 151.100 173.000 153.000 ;
        RECT 174.200 151.100 174.600 153.000 ;
        RECT 175.000 151.100 175.400 153.100 ;
        RECT 176.100 152.800 177.000 153.100 ;
        RECT 176.100 151.100 176.500 152.800 ;
        RECT 178.200 152.500 178.500 153.600 ;
        RECT 180.800 153.500 181.100 153.800 ;
        RECT 180.700 153.300 181.100 153.500 ;
        RECT 180.300 153.000 181.100 153.300 ;
        RECT 183.000 153.600 183.400 155.300 ;
        RECT 184.700 155.200 185.100 155.300 ;
        RECT 183.900 154.900 184.300 155.000 ;
        RECT 183.900 154.600 185.800 154.900 ;
        RECT 185.400 154.500 185.800 154.600 ;
        RECT 186.300 154.200 186.600 155.800 ;
        RECT 187.300 155.900 187.600 156.500 ;
        RECT 187.900 156.500 188.300 156.600 ;
        RECT 190.200 156.500 190.600 156.600 ;
        RECT 187.900 156.200 190.600 156.500 ;
        RECT 187.300 155.700 189.700 155.900 ;
        RECT 191.800 155.700 192.200 159.900 ;
        RECT 187.300 155.600 192.200 155.700 ;
        RECT 189.300 155.500 192.200 155.600 ;
        RECT 189.400 155.400 192.200 155.500 ;
        RECT 188.600 155.100 189.000 155.200 ;
        RECT 193.400 155.100 193.800 159.900 ;
        RECT 195.400 156.800 195.800 157.200 ;
        RECT 194.200 155.800 194.600 156.600 ;
        RECT 195.400 156.200 195.700 156.800 ;
        RECT 196.100 156.200 196.500 159.900 ;
        RECT 195.000 155.900 195.700 156.200 ;
        RECT 196.000 155.900 196.500 156.200 ;
        RECT 199.500 156.200 199.900 159.900 ;
        RECT 200.200 156.800 200.600 157.200 ;
        RECT 200.300 156.200 200.600 156.800 ;
        RECT 199.500 155.900 200.000 156.200 ;
        RECT 200.300 156.100 201.000 156.200 ;
        RECT 201.400 156.100 201.800 156.200 ;
        RECT 200.300 155.900 201.800 156.100 ;
        RECT 195.000 155.800 195.400 155.900 ;
        RECT 195.000 155.100 195.300 155.800 ;
        RECT 196.000 155.200 196.300 155.900 ;
        RECT 188.600 154.800 191.100 155.100 ;
        RECT 190.700 154.700 191.100 154.800 ;
        RECT 193.400 154.800 195.300 155.100 ;
        RECT 195.800 154.800 196.300 155.200 ;
        RECT 189.900 154.200 190.300 154.300 ;
        RECT 186.300 153.900 191.800 154.200 ;
        RECT 186.500 153.800 186.900 153.900 ;
        RECT 189.400 153.800 189.800 153.900 ;
        RECT 191.000 153.800 191.800 153.900 ;
        RECT 183.000 153.300 184.900 153.600 ;
        RECT 178.200 151.500 178.600 152.500 ;
        RECT 180.300 151.500 180.700 153.000 ;
        RECT 183.000 151.100 183.400 153.300 ;
        RECT 184.500 153.200 184.900 153.300 ;
        RECT 189.400 152.800 189.700 153.800 ;
        RECT 188.500 152.700 188.900 152.800 ;
        RECT 185.400 152.100 185.800 152.500 ;
        RECT 187.500 152.400 188.900 152.700 ;
        RECT 189.400 152.400 189.800 152.800 ;
        RECT 187.500 152.100 187.800 152.400 ;
        RECT 190.200 152.100 190.600 152.500 ;
        RECT 185.100 151.800 185.800 152.100 ;
        RECT 185.100 151.100 185.700 151.800 ;
        RECT 187.400 151.100 187.800 152.100 ;
        RECT 189.600 151.800 190.600 152.100 ;
        RECT 189.600 151.100 190.000 151.800 ;
        RECT 191.800 151.100 192.200 153.500 ;
        RECT 192.600 153.400 193.000 154.200 ;
        RECT 193.400 153.100 193.800 154.800 ;
        RECT 196.000 154.200 196.300 154.800 ;
        RECT 196.600 154.400 197.000 155.200 ;
        RECT 199.000 154.400 199.400 155.200 ;
        RECT 199.700 155.100 200.000 155.900 ;
        RECT 200.600 155.800 201.800 155.900 ;
        RECT 203.000 155.800 203.400 156.600 ;
        RECT 202.200 155.100 202.600 155.200 ;
        RECT 199.700 154.800 202.600 155.100 ;
        RECT 199.700 154.200 200.000 154.800 ;
        RECT 195.000 153.800 196.300 154.200 ;
        RECT 197.400 154.100 197.800 154.200 ;
        RECT 198.200 154.100 198.600 154.200 ;
        RECT 197.000 153.800 199.000 154.100 ;
        RECT 199.700 153.800 201.000 154.200 ;
        RECT 201.400 154.100 201.800 154.200 ;
        RECT 203.800 154.100 204.200 159.900 ;
        RECT 205.400 155.600 205.800 159.900 ;
        RECT 207.500 157.900 208.100 159.900 ;
        RECT 209.800 157.900 210.200 159.900 ;
        RECT 212.000 158.200 212.400 159.900 ;
        RECT 212.000 157.900 213.000 158.200 ;
        RECT 207.800 157.500 208.200 157.900 ;
        RECT 209.900 157.600 210.200 157.900 ;
        RECT 209.500 157.300 211.300 157.600 ;
        RECT 212.600 157.500 213.000 157.900 ;
        RECT 209.500 157.200 209.900 157.300 ;
        RECT 210.900 157.200 211.300 157.300 ;
        RECT 207.000 157.000 207.700 157.200 ;
        RECT 207.000 156.800 208.100 157.000 ;
        RECT 207.400 156.600 208.100 156.800 ;
        RECT 207.800 156.100 208.100 156.600 ;
        RECT 208.900 156.500 210.000 156.800 ;
        RECT 208.900 156.400 209.300 156.500 ;
        RECT 207.800 155.800 209.000 156.100 ;
        RECT 205.400 155.300 207.500 155.600 ;
        RECT 201.400 153.800 204.200 154.100 ;
        RECT 195.100 153.100 195.400 153.800 ;
        RECT 197.000 153.600 197.400 153.800 ;
        RECT 198.600 153.600 199.000 153.800 ;
        RECT 195.900 153.100 197.700 153.300 ;
        RECT 198.300 153.100 200.100 153.300 ;
        RECT 200.600 153.100 200.900 153.800 ;
        RECT 203.800 153.100 204.200 153.800 ;
        RECT 204.600 153.400 205.000 154.200 ;
        RECT 205.400 153.600 205.800 155.300 ;
        RECT 207.100 155.200 207.500 155.300 ;
        RECT 206.300 154.900 206.700 155.000 ;
        RECT 206.300 154.600 208.200 154.900 ;
        RECT 207.800 154.500 208.200 154.600 ;
        RECT 208.700 154.200 209.000 155.800 ;
        RECT 209.700 155.900 210.000 156.500 ;
        RECT 210.300 156.500 210.700 156.600 ;
        RECT 212.600 156.500 213.000 156.600 ;
        RECT 210.300 156.200 213.000 156.500 ;
        RECT 209.700 155.700 212.100 155.900 ;
        RECT 214.200 155.700 214.600 159.900 ;
        RECT 209.700 155.600 214.600 155.700 ;
        RECT 211.700 155.500 214.600 155.600 ;
        RECT 211.800 155.400 214.600 155.500 ;
        RECT 215.000 155.600 215.400 159.900 ;
        RECT 217.100 157.900 217.700 159.900 ;
        RECT 219.400 157.900 219.800 159.900 ;
        RECT 221.600 158.200 222.000 159.900 ;
        RECT 221.600 157.900 222.600 158.200 ;
        RECT 217.400 157.500 217.800 157.900 ;
        RECT 219.500 157.600 219.800 157.900 ;
        RECT 219.100 157.300 220.900 157.600 ;
        RECT 222.200 157.500 222.600 157.900 ;
        RECT 219.100 157.200 219.500 157.300 ;
        RECT 220.500 157.200 220.900 157.300 ;
        RECT 217.000 156.600 217.700 157.000 ;
        RECT 217.400 156.100 217.700 156.600 ;
        RECT 218.500 156.500 219.600 156.800 ;
        RECT 218.500 156.400 218.900 156.500 ;
        RECT 217.400 155.800 218.600 156.100 ;
        RECT 215.000 155.300 217.100 155.600 ;
        RECT 210.200 155.100 210.600 155.200 ;
        RECT 211.000 155.100 211.400 155.200 ;
        RECT 210.200 154.800 213.500 155.100 ;
        RECT 213.100 154.700 213.500 154.800 ;
        RECT 212.300 154.200 212.700 154.300 ;
        RECT 208.700 153.900 214.200 154.200 ;
        RECT 208.900 153.800 209.300 153.900 ;
        RECT 193.400 152.800 194.300 153.100 ;
        RECT 193.900 151.100 194.300 152.800 ;
        RECT 195.000 151.100 195.400 153.100 ;
        RECT 195.800 153.000 197.800 153.100 ;
        RECT 195.800 151.100 196.200 153.000 ;
        RECT 197.400 151.100 197.800 153.000 ;
        RECT 198.200 153.000 200.200 153.100 ;
        RECT 198.200 151.100 198.600 153.000 ;
        RECT 199.800 151.100 200.200 153.000 ;
        RECT 200.600 151.100 201.000 153.100 ;
        RECT 203.300 152.800 204.200 153.100 ;
        RECT 205.400 153.300 207.300 153.600 ;
        RECT 203.300 151.100 203.700 152.800 ;
        RECT 205.400 151.100 205.800 153.300 ;
        RECT 206.900 153.200 207.300 153.300 ;
        RECT 211.800 152.800 212.100 153.900 ;
        RECT 213.400 153.800 214.200 153.900 ;
        RECT 215.000 153.600 215.400 155.300 ;
        RECT 216.700 155.200 217.100 155.300 ;
        RECT 215.900 154.900 216.300 155.000 ;
        RECT 215.900 154.600 217.800 154.900 ;
        RECT 217.400 154.500 217.800 154.600 ;
        RECT 218.300 154.200 218.600 155.800 ;
        RECT 219.300 155.900 219.600 156.500 ;
        RECT 219.900 156.500 220.300 156.600 ;
        RECT 222.200 156.500 222.600 156.600 ;
        RECT 219.900 156.200 222.600 156.500 ;
        RECT 219.300 155.700 221.700 155.900 ;
        RECT 223.800 155.700 224.200 159.900 ;
        RECT 219.300 155.600 224.200 155.700 ;
        RECT 221.300 155.500 224.200 155.600 ;
        RECT 221.400 155.400 224.200 155.500 ;
        RECT 225.400 155.600 225.800 159.900 ;
        RECT 227.000 155.600 227.400 159.900 ;
        RECT 228.600 155.600 229.000 159.900 ;
        RECT 230.200 155.600 230.600 159.900 ;
        RECT 233.100 156.200 233.500 159.900 ;
        RECT 233.800 156.800 234.200 157.200 ;
        RECT 233.900 156.200 234.200 156.800 ;
        RECT 233.100 155.900 233.600 156.200 ;
        RECT 233.900 155.900 234.600 156.200 ;
        RECT 225.400 155.200 226.300 155.600 ;
        RECT 227.000 155.200 228.100 155.600 ;
        RECT 228.600 155.200 229.700 155.600 ;
        RECT 230.200 155.200 231.400 155.600 ;
        RECT 220.600 155.100 221.000 155.200 ;
        RECT 220.600 154.800 223.100 155.100 ;
        RECT 222.700 154.700 223.100 154.800 ;
        RECT 225.900 154.500 226.300 155.200 ;
        RECT 227.700 154.500 228.100 155.200 ;
        RECT 229.300 154.500 229.700 155.200 ;
        RECT 221.900 154.200 222.300 154.300 ;
        RECT 218.300 153.900 223.800 154.200 ;
        RECT 218.500 153.800 218.900 153.900 ;
        RECT 210.900 152.700 211.300 152.800 ;
        RECT 207.800 152.100 208.200 152.500 ;
        RECT 209.900 152.400 211.300 152.700 ;
        RECT 211.800 152.400 212.200 152.800 ;
        RECT 209.900 152.100 210.200 152.400 ;
        RECT 212.600 152.100 213.000 152.500 ;
        RECT 207.500 151.800 208.200 152.100 ;
        RECT 207.500 151.100 208.100 151.800 ;
        RECT 209.800 151.100 210.200 152.100 ;
        RECT 212.000 151.800 213.000 152.100 ;
        RECT 212.000 151.100 212.400 151.800 ;
        RECT 214.200 151.100 214.600 153.500 ;
        RECT 215.000 153.300 216.900 153.600 ;
        RECT 215.000 151.100 215.400 153.300 ;
        RECT 216.500 153.200 216.900 153.300 ;
        RECT 221.400 152.800 221.700 153.900 ;
        RECT 223.000 153.800 223.800 153.900 ;
        RECT 225.900 154.100 227.200 154.500 ;
        RECT 227.700 154.100 228.900 154.500 ;
        RECT 229.300 154.100 230.600 154.500 ;
        RECT 225.900 153.800 226.300 154.100 ;
        RECT 227.700 153.800 228.100 154.100 ;
        RECT 229.300 153.800 229.700 154.100 ;
        RECT 231.000 153.800 231.400 155.200 ;
        RECT 232.600 154.400 233.000 155.200 ;
        RECT 233.300 154.200 233.600 155.900 ;
        RECT 234.200 155.800 234.600 155.900 ;
        RECT 235.000 155.800 235.400 156.600 ;
        RECT 234.200 155.100 234.500 155.800 ;
        RECT 235.800 155.100 236.200 159.900 ;
        RECT 236.600 157.100 237.000 157.200 ;
        RECT 237.400 157.100 237.800 159.900 ;
        RECT 239.500 157.900 240.100 159.900 ;
        RECT 241.800 157.900 242.200 159.900 ;
        RECT 244.000 158.200 244.400 159.900 ;
        RECT 244.000 157.900 245.000 158.200 ;
        RECT 239.800 157.500 240.200 157.900 ;
        RECT 241.900 157.600 242.200 157.900 ;
        RECT 241.500 157.300 243.300 157.600 ;
        RECT 244.600 157.500 245.000 157.900 ;
        RECT 241.500 157.200 241.900 157.300 ;
        RECT 242.900 157.200 243.300 157.300 ;
        RECT 236.600 156.800 237.800 157.100 ;
        RECT 234.200 154.800 236.200 155.100 ;
        RECT 231.800 154.100 232.200 154.200 ;
        RECT 233.300 154.100 234.600 154.200 ;
        RECT 235.000 154.100 235.400 154.200 ;
        RECT 231.800 153.800 232.600 154.100 ;
        RECT 233.300 153.800 235.400 154.100 ;
        RECT 220.500 152.700 220.900 152.800 ;
        RECT 217.400 152.100 217.800 152.500 ;
        RECT 219.500 152.400 220.900 152.700 ;
        RECT 221.400 152.400 221.800 152.800 ;
        RECT 219.500 152.100 219.800 152.400 ;
        RECT 222.200 152.100 222.600 152.500 ;
        RECT 217.100 151.800 217.800 152.100 ;
        RECT 217.100 151.100 217.700 151.800 ;
        RECT 219.400 151.100 219.800 152.100 ;
        RECT 221.600 151.800 222.600 152.100 ;
        RECT 221.600 151.100 222.000 151.800 ;
        RECT 223.800 151.100 224.200 153.500 ;
        RECT 225.400 153.400 226.300 153.800 ;
        RECT 227.000 153.400 228.100 153.800 ;
        RECT 228.600 153.400 229.700 153.800 ;
        RECT 230.200 153.400 231.400 153.800 ;
        RECT 232.200 153.600 232.600 153.800 ;
        RECT 225.400 151.100 225.800 153.400 ;
        RECT 227.000 151.100 227.400 153.400 ;
        RECT 228.600 151.100 229.000 153.400 ;
        RECT 230.200 151.100 230.600 153.400 ;
        RECT 231.900 153.100 233.700 153.300 ;
        RECT 234.200 153.100 234.500 153.800 ;
        RECT 235.800 153.100 236.200 154.800 ;
        RECT 237.400 155.600 237.800 156.800 ;
        RECT 239.400 156.600 240.100 157.000 ;
        RECT 239.800 156.100 240.100 156.600 ;
        RECT 240.900 156.500 242.000 156.800 ;
        RECT 240.900 156.400 241.300 156.500 ;
        RECT 239.800 155.800 241.000 156.100 ;
        RECT 237.400 155.300 239.500 155.600 ;
        RECT 236.600 153.400 237.000 154.200 ;
        RECT 237.400 153.600 237.800 155.300 ;
        RECT 239.100 155.200 239.500 155.300 ;
        RECT 238.300 154.900 238.700 155.000 ;
        RECT 238.300 154.600 240.200 154.900 ;
        RECT 239.800 154.500 240.200 154.600 ;
        RECT 240.700 154.200 241.000 155.800 ;
        RECT 241.700 155.900 242.000 156.500 ;
        RECT 242.300 156.500 242.700 156.600 ;
        RECT 244.600 156.500 245.000 156.600 ;
        RECT 242.300 156.200 245.000 156.500 ;
        RECT 241.700 155.700 244.100 155.900 ;
        RECT 246.200 155.700 246.600 159.900 ;
        RECT 248.300 156.300 248.700 159.900 ;
        RECT 247.800 155.900 248.700 156.300 ;
        RECT 241.700 155.600 246.600 155.700 ;
        RECT 243.700 155.500 246.600 155.600 ;
        RECT 243.800 155.400 246.600 155.500 ;
        RECT 243.000 155.100 243.400 155.200 ;
        RECT 243.000 154.800 245.500 155.100 ;
        RECT 245.100 154.700 245.500 154.800 ;
        RECT 244.300 154.200 244.700 154.300 ;
        RECT 247.900 154.200 248.200 155.900 ;
        RECT 248.600 154.800 249.000 155.600 ;
        RECT 240.700 153.900 246.200 154.200 ;
        RECT 240.900 153.800 241.300 153.900 ;
        RECT 231.800 153.000 233.800 153.100 ;
        RECT 231.800 151.100 232.200 153.000 ;
        RECT 233.400 151.100 233.800 153.000 ;
        RECT 234.200 151.100 234.600 153.100 ;
        RECT 235.300 152.800 236.200 153.100 ;
        RECT 237.400 153.300 239.300 153.600 ;
        RECT 235.300 151.100 235.700 152.800 ;
        RECT 237.400 151.100 237.800 153.300 ;
        RECT 238.900 153.200 239.300 153.300 ;
        RECT 243.800 152.800 244.100 153.900 ;
        RECT 245.400 153.800 246.200 153.900 ;
        RECT 247.800 153.800 248.200 154.200 ;
        RECT 248.600 154.100 249.000 154.200 ;
        RECT 249.400 154.100 249.800 154.200 ;
        RECT 248.600 153.800 249.800 154.100 ;
        RECT 242.900 152.700 243.300 152.800 ;
        RECT 239.800 152.100 240.200 152.500 ;
        RECT 241.900 152.400 243.300 152.700 ;
        RECT 243.800 152.400 244.200 152.800 ;
        RECT 241.900 152.100 242.200 152.400 ;
        RECT 244.600 152.100 245.000 152.500 ;
        RECT 239.500 151.800 240.200 152.100 ;
        RECT 239.500 151.100 240.100 151.800 ;
        RECT 241.800 151.100 242.200 152.100 ;
        RECT 244.000 151.800 245.000 152.100 ;
        RECT 244.000 151.100 244.400 151.800 ;
        RECT 246.200 151.100 246.600 153.500 ;
        RECT 247.000 152.400 247.400 153.200 ;
        RECT 247.900 152.200 248.200 153.800 ;
        RECT 249.400 153.400 249.800 153.800 ;
        RECT 250.200 153.100 250.600 159.900 ;
        RECT 251.000 156.100 251.400 156.600 ;
        RECT 251.800 156.100 252.200 156.200 ;
        RECT 251.000 155.800 252.200 156.100 ;
        RECT 250.200 152.800 251.100 153.100 ;
        RECT 250.700 152.200 251.100 152.800 ;
        RECT 247.800 151.100 248.200 152.200 ;
        RECT 250.200 151.800 251.100 152.200 ;
        RECT 250.700 151.100 251.100 151.800 ;
        RECT 0.600 147.500 1.000 149.900 ;
        RECT 2.800 149.200 3.200 149.900 ;
        RECT 2.200 148.900 3.200 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.100 149.200 7.700 149.900 ;
        RECT 7.000 148.900 7.700 149.200 ;
        RECT 2.200 148.500 2.600 148.900 ;
        RECT 5.000 148.600 5.300 148.900 ;
        RECT 3.000 148.200 3.400 148.600 ;
        RECT 3.900 148.300 5.300 148.600 ;
        RECT 7.000 148.500 7.400 148.900 ;
        RECT 3.900 148.200 4.300 148.300 ;
        RECT 1.000 147.100 1.800 147.200 ;
        RECT 3.100 147.100 3.400 148.200 ;
        RECT 7.900 147.700 8.300 147.800 ;
        RECT 9.400 147.700 9.800 149.900 ;
        RECT 11.500 148.200 11.900 149.900 ;
        RECT 7.900 147.400 9.800 147.700 ;
        RECT 11.000 147.900 11.900 148.200 ;
        RECT 12.600 147.900 13.000 149.900 ;
        RECT 13.400 148.000 13.800 149.900 ;
        RECT 15.000 148.000 15.400 149.900 ;
        RECT 13.400 147.900 15.400 148.000 ;
        RECT 5.900 147.100 6.300 147.200 ;
        RECT 1.000 146.800 6.500 147.100 ;
        RECT 2.500 146.700 2.900 146.800 ;
        RECT 1.700 146.200 2.100 146.300 ;
        RECT 1.700 145.900 4.200 146.200 ;
        RECT 3.800 145.800 4.200 145.900 ;
        RECT 5.400 146.100 5.800 146.200 ;
        RECT 6.200 146.100 6.500 146.800 ;
        RECT 7.000 146.400 7.400 146.500 ;
        RECT 7.000 146.100 8.900 146.400 ;
        RECT 5.400 145.800 6.500 146.100 ;
        RECT 8.500 146.000 8.900 146.100 ;
        RECT 0.600 145.500 3.400 145.600 ;
        RECT 0.600 145.400 3.500 145.500 ;
        RECT 0.600 145.300 5.500 145.400 ;
        RECT 0.600 141.100 1.000 145.300 ;
        RECT 3.100 145.100 5.500 145.300 ;
        RECT 2.200 144.500 4.900 144.800 ;
        RECT 2.200 144.400 2.600 144.500 ;
        RECT 4.500 144.400 4.900 144.500 ;
        RECT 5.200 144.500 5.500 145.100 ;
        RECT 6.200 145.200 6.500 145.800 ;
        RECT 7.700 145.700 8.100 145.800 ;
        RECT 9.400 145.700 9.800 147.400 ;
        RECT 10.200 146.800 10.600 147.600 ;
        RECT 7.700 145.400 9.800 145.700 ;
        RECT 6.200 144.900 7.400 145.200 ;
        RECT 5.900 144.500 6.300 144.600 ;
        RECT 5.200 144.200 6.300 144.500 ;
        RECT 7.100 144.400 7.400 144.900 ;
        RECT 7.100 144.000 7.800 144.400 ;
        RECT 9.400 144.100 9.800 145.400 ;
        RECT 11.000 146.100 11.400 147.900 ;
        RECT 12.700 147.200 13.000 147.900 ;
        RECT 13.500 147.700 15.300 147.900 ;
        RECT 15.800 147.500 16.200 149.900 ;
        RECT 18.000 149.200 18.400 149.900 ;
        RECT 17.400 148.900 18.400 149.200 ;
        RECT 20.200 148.900 20.600 149.900 ;
        RECT 22.300 149.200 22.900 149.900 ;
        RECT 22.200 148.900 22.900 149.200 ;
        RECT 17.400 148.500 17.800 148.900 ;
        RECT 20.200 148.600 20.500 148.900 ;
        RECT 18.200 148.200 18.600 148.600 ;
        RECT 19.100 148.300 20.500 148.600 ;
        RECT 22.200 148.500 22.600 148.900 ;
        RECT 19.100 148.200 19.500 148.300 ;
        RECT 14.600 147.200 15.000 147.400 ;
        RECT 11.800 147.100 12.200 147.200 ;
        RECT 12.600 147.100 13.900 147.200 ;
        RECT 11.800 146.800 13.900 147.100 ;
        RECT 14.600 146.900 15.400 147.200 ;
        RECT 15.000 146.800 15.400 146.900 ;
        RECT 16.200 147.100 17.000 147.200 ;
        RECT 18.300 147.100 18.600 148.200 ;
        RECT 23.100 147.700 23.500 147.800 ;
        RECT 24.600 147.700 25.000 149.900 ;
        RECT 25.400 148.000 25.800 149.900 ;
        RECT 27.000 148.000 27.400 149.900 ;
        RECT 25.400 147.900 27.400 148.000 ;
        RECT 27.800 147.900 28.200 149.900 ;
        RECT 28.900 148.200 29.300 149.900 ;
        RECT 28.900 147.900 29.800 148.200 ;
        RECT 25.500 147.700 27.300 147.900 ;
        RECT 23.100 147.400 25.000 147.700 ;
        RECT 21.100 147.100 21.500 147.200 ;
        RECT 16.200 146.800 21.700 147.100 ;
        RECT 11.000 145.800 12.900 146.100 ;
        RECT 10.200 144.100 10.600 144.200 ;
        RECT 9.400 143.800 10.600 144.100 ;
        RECT 3.900 143.700 4.300 143.800 ;
        RECT 5.300 143.700 5.700 143.800 ;
        RECT 2.200 143.100 2.600 143.500 ;
        RECT 3.900 143.400 5.700 143.700 ;
        RECT 5.000 143.100 5.300 143.400 ;
        RECT 7.000 143.100 7.400 143.500 ;
        RECT 2.200 142.800 3.200 143.100 ;
        RECT 2.800 141.100 3.200 142.800 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.100 141.100 7.700 143.100 ;
        RECT 9.400 141.100 9.800 143.800 ;
        RECT 11.000 141.100 11.400 145.800 ;
        RECT 12.600 145.200 12.900 145.800 ;
        RECT 11.800 144.400 12.200 145.200 ;
        RECT 12.600 145.100 13.000 145.200 ;
        RECT 13.600 145.100 13.900 146.800 ;
        RECT 17.700 146.700 18.100 146.800 ;
        RECT 14.200 145.800 14.600 146.600 ;
        RECT 16.900 146.200 17.300 146.300 ;
        RECT 16.900 146.100 19.400 146.200 ;
        RECT 19.800 146.100 20.200 146.200 ;
        RECT 16.900 145.900 20.200 146.100 ;
        RECT 19.000 145.800 20.200 145.900 ;
        RECT 15.800 145.500 18.600 145.600 ;
        RECT 15.800 145.400 18.700 145.500 ;
        RECT 15.800 145.300 20.700 145.400 ;
        RECT 12.600 144.800 13.300 145.100 ;
        RECT 13.600 144.800 14.100 145.100 ;
        RECT 13.000 144.200 13.300 144.800 ;
        RECT 13.000 143.800 13.400 144.200 ;
        RECT 13.700 141.100 14.100 144.800 ;
        RECT 15.800 141.100 16.200 145.300 ;
        RECT 18.300 145.100 20.700 145.300 ;
        RECT 17.400 144.500 20.100 144.800 ;
        RECT 17.400 144.400 17.800 144.500 ;
        RECT 19.700 144.400 20.100 144.500 ;
        RECT 20.400 144.500 20.700 145.100 ;
        RECT 21.400 145.200 21.700 146.800 ;
        RECT 22.200 146.400 22.600 146.500 ;
        RECT 22.200 146.100 24.100 146.400 ;
        RECT 23.700 146.000 24.100 146.100 ;
        RECT 22.900 145.700 23.300 145.800 ;
        RECT 24.600 145.700 25.000 147.400 ;
        RECT 25.800 147.200 26.200 147.400 ;
        RECT 27.800 147.200 28.100 147.900 ;
        RECT 25.400 146.900 26.200 147.200 ;
        RECT 25.400 146.800 25.800 146.900 ;
        RECT 26.900 146.800 28.200 147.200 ;
        RECT 26.200 145.800 26.600 146.600 ;
        RECT 26.900 146.200 27.200 146.800 ;
        RECT 26.900 145.800 27.400 146.200 ;
        RECT 29.400 146.100 29.800 147.900 ;
        RECT 30.200 146.800 30.600 147.600 ;
        RECT 27.800 145.800 29.800 146.100 ;
        RECT 22.900 145.400 25.000 145.700 ;
        RECT 21.400 144.900 22.600 145.200 ;
        RECT 21.100 144.500 21.500 144.600 ;
        RECT 20.400 144.200 21.500 144.500 ;
        RECT 22.300 144.400 22.600 144.900 ;
        RECT 22.300 144.000 23.000 144.400 ;
        RECT 19.100 143.700 19.500 143.800 ;
        RECT 20.500 143.700 20.900 143.800 ;
        RECT 17.400 143.100 17.800 143.500 ;
        RECT 19.100 143.400 20.900 143.700 ;
        RECT 20.200 143.100 20.500 143.400 ;
        RECT 22.200 143.100 22.600 143.500 ;
        RECT 17.400 142.800 18.400 143.100 ;
        RECT 18.000 141.100 18.400 142.800 ;
        RECT 20.200 141.100 20.600 143.100 ;
        RECT 22.300 141.100 22.900 143.100 ;
        RECT 24.600 141.100 25.000 145.400 ;
        RECT 26.900 145.100 27.200 145.800 ;
        RECT 27.800 145.200 28.100 145.800 ;
        RECT 27.800 145.100 28.200 145.200 ;
        RECT 26.700 144.800 27.200 145.100 ;
        RECT 27.500 144.800 28.200 145.100 ;
        RECT 26.700 141.100 27.100 144.800 ;
        RECT 27.500 144.200 27.800 144.800 ;
        RECT 28.600 144.400 29.000 145.200 ;
        RECT 27.400 143.800 27.800 144.200 ;
        RECT 29.400 141.100 29.800 145.800 ;
        RECT 31.800 146.100 32.200 149.900 ;
        RECT 33.900 149.200 34.300 149.900 ;
        RECT 35.300 149.200 35.700 149.900 ;
        RECT 33.400 148.800 34.300 149.200 ;
        RECT 35.000 148.800 35.700 149.200 ;
        RECT 33.900 148.200 34.300 148.800 ;
        RECT 33.400 147.900 34.300 148.200 ;
        RECT 35.300 148.200 35.700 148.800 ;
        RECT 35.300 147.900 36.200 148.200 ;
        RECT 31.800 145.800 32.900 146.100 ;
        RECT 31.800 141.100 32.200 145.800 ;
        RECT 32.600 145.200 32.900 145.800 ;
        RECT 32.600 144.800 33.000 145.200 ;
        RECT 33.400 141.100 33.800 147.900 ;
        RECT 34.200 145.100 34.600 145.200 ;
        RECT 35.000 145.100 35.400 145.200 ;
        RECT 34.200 144.800 35.400 145.100 ;
        RECT 34.200 144.400 34.600 144.800 ;
        RECT 35.000 144.400 35.400 144.800 ;
        RECT 35.800 141.100 36.200 147.900 ;
        RECT 36.600 147.100 37.000 147.600 ;
        RECT 37.400 147.100 37.800 149.900 ;
        RECT 40.900 148.000 41.300 149.500 ;
        RECT 43.000 148.500 43.400 149.500 ;
        RECT 40.500 147.700 41.300 148.000 ;
        RECT 40.500 147.500 40.900 147.700 ;
        RECT 40.500 147.200 40.800 147.500 ;
        RECT 43.100 147.400 43.400 148.500 ;
        RECT 45.100 148.200 45.500 149.900 ;
        RECT 47.500 148.200 47.900 149.900 ;
        RECT 51.000 148.900 51.400 149.900 ;
        RECT 36.600 146.800 37.800 147.100 ;
        RECT 39.800 146.800 40.800 147.200 ;
        RECT 41.300 147.100 43.400 147.400 ;
        RECT 44.600 147.900 45.500 148.200 ;
        RECT 47.000 147.900 47.900 148.200 ;
        RECT 44.600 147.100 45.000 147.900 ;
        RECT 45.400 147.100 45.800 147.200 ;
        RECT 41.300 146.900 41.800 147.100 ;
        RECT 37.400 141.100 37.800 146.800 ;
        RECT 39.800 145.400 40.200 146.200 ;
        RECT 40.500 144.900 40.800 146.800 ;
        RECT 41.100 146.500 41.800 146.900 ;
        RECT 44.600 146.800 45.800 147.100 ;
        RECT 41.500 145.500 41.800 146.500 ;
        RECT 42.200 145.800 42.600 146.600 ;
        RECT 43.000 145.800 43.400 146.600 ;
        RECT 41.500 145.200 43.400 145.500 ;
        RECT 40.500 144.600 41.300 144.900 ;
        RECT 40.900 142.200 41.300 144.600 ;
        RECT 43.100 143.500 43.400 145.200 ;
        RECT 40.900 141.800 41.800 142.200 ;
        RECT 40.900 141.100 41.300 141.800 ;
        RECT 43.000 141.500 43.400 143.500 ;
        RECT 44.600 141.100 45.000 146.800 ;
        RECT 47.000 141.100 47.400 147.900 ;
        RECT 51.100 147.200 51.400 148.900 ;
        RECT 53.400 148.900 53.800 149.900 ;
        RECT 53.400 147.200 53.700 148.900 ;
        RECT 55.800 148.800 56.200 149.900 ;
        RECT 58.200 148.900 58.600 149.900 ;
        RECT 54.200 147.800 54.600 148.600 ;
        RECT 54.200 147.200 54.500 147.800 ;
        RECT 55.900 147.200 56.200 148.800 ;
        RECT 56.600 148.100 57.000 148.200 ;
        RECT 57.400 148.100 57.800 148.600 ;
        RECT 56.600 147.800 57.800 148.100 ;
        RECT 58.300 147.800 58.600 148.900 ;
        RECT 59.800 147.900 60.200 149.900 ;
        RECT 58.300 147.500 59.500 147.800 ;
        RECT 51.000 146.800 51.400 147.200 ;
        RECT 47.800 144.400 48.200 145.200 ;
        RECT 51.100 145.100 51.400 146.800 ;
        RECT 51.800 146.800 52.200 147.200 ;
        RECT 53.400 146.800 53.800 147.200 ;
        RECT 54.200 146.800 54.600 147.200 ;
        RECT 55.800 146.800 56.200 147.200 ;
        RECT 58.200 146.800 58.700 147.200 ;
        RECT 51.800 146.200 52.100 146.800 ;
        RECT 51.800 146.100 52.200 146.200 ;
        RECT 52.600 146.100 53.000 146.200 ;
        RECT 51.800 145.800 53.000 146.100 ;
        RECT 51.800 145.400 52.200 145.800 ;
        RECT 52.600 145.400 53.000 145.800 ;
        RECT 53.400 145.100 53.700 146.800 ;
        RECT 55.900 145.100 56.200 146.800 ;
        RECT 58.400 146.400 58.800 146.800 ;
        RECT 56.600 145.400 57.000 146.200 ;
        RECT 59.200 146.000 59.500 147.500 ;
        RECT 59.900 147.100 60.200 147.900 ;
        RECT 61.400 147.600 61.800 149.900 ;
        RECT 63.000 147.600 63.400 149.900 ;
        RECT 60.600 147.100 61.000 147.600 ;
        RECT 61.400 147.200 63.400 147.600 ;
        RECT 64.600 147.500 65.000 149.900 ;
        RECT 66.800 149.200 67.200 149.900 ;
        RECT 66.200 148.900 67.200 149.200 ;
        RECT 69.000 148.900 69.400 149.900 ;
        RECT 71.100 149.200 71.700 149.900 ;
        RECT 71.000 148.900 71.700 149.200 ;
        RECT 66.200 148.500 66.600 148.900 ;
        RECT 69.000 148.600 69.300 148.900 ;
        RECT 67.000 148.200 67.400 148.600 ;
        RECT 67.900 148.300 69.300 148.600 ;
        RECT 71.000 148.500 71.400 148.900 ;
        RECT 67.900 148.200 68.300 148.300 ;
        RECT 59.800 146.800 61.000 147.100 ;
        RECT 59.900 146.200 60.200 146.800 ;
        RECT 59.100 145.700 59.500 146.000 ;
        RECT 59.800 145.800 60.200 146.200 ;
        RECT 63.000 145.800 63.400 147.200 ;
        RECT 65.000 147.100 65.800 147.200 ;
        RECT 67.100 147.100 67.400 148.200 ;
        RECT 71.900 147.700 72.300 147.800 ;
        RECT 73.400 147.700 73.800 149.900 ;
        RECT 74.300 148.200 74.700 148.600 ;
        RECT 74.200 147.800 74.600 148.200 ;
        RECT 75.000 147.900 75.400 149.900 ;
        RECT 77.700 148.200 78.100 149.900 ;
        RECT 77.700 147.900 78.600 148.200 ;
        RECT 71.900 147.400 73.800 147.700 ;
        RECT 68.600 147.100 69.000 147.200 ;
        RECT 69.900 147.100 70.300 147.200 ;
        RECT 65.000 146.800 70.500 147.100 ;
        RECT 66.500 146.700 66.900 146.800 ;
        RECT 65.700 146.200 66.100 146.300 ;
        RECT 65.700 145.900 68.200 146.200 ;
        RECT 67.800 145.800 68.200 145.900 ;
        RECT 57.400 145.600 59.500 145.700 ;
        RECT 57.400 145.400 59.400 145.600 ;
        RECT 51.000 144.700 51.900 145.100 ;
        RECT 51.500 142.200 51.900 144.700 ;
        RECT 52.900 144.700 53.800 145.100 ;
        RECT 55.800 144.700 56.700 145.100 ;
        RECT 52.900 142.200 53.300 144.700 ;
        RECT 51.500 141.800 52.200 142.200 ;
        RECT 52.900 141.800 53.800 142.200 ;
        RECT 51.500 141.100 51.900 141.800 ;
        RECT 52.900 141.100 53.300 141.800 ;
        RECT 56.300 141.100 56.700 144.700 ;
        RECT 57.400 141.100 57.800 145.400 ;
        RECT 59.900 145.100 60.200 145.800 ;
        RECT 59.500 144.800 60.200 145.100 ;
        RECT 61.400 145.400 63.400 145.800 ;
        RECT 59.500 141.100 59.900 144.800 ;
        RECT 61.400 141.100 61.800 145.400 ;
        RECT 63.000 141.100 63.400 145.400 ;
        RECT 64.600 145.500 67.400 145.600 ;
        RECT 64.600 145.400 67.500 145.500 ;
        RECT 64.600 145.300 69.500 145.400 ;
        RECT 64.600 141.100 65.000 145.300 ;
        RECT 67.100 145.100 69.500 145.300 ;
        RECT 66.200 144.500 68.900 144.800 ;
        RECT 66.200 144.400 66.600 144.500 ;
        RECT 68.500 144.400 68.900 144.500 ;
        RECT 69.200 144.500 69.500 145.100 ;
        RECT 70.200 145.200 70.500 146.800 ;
        RECT 71.000 146.400 71.400 146.500 ;
        RECT 71.000 146.100 72.900 146.400 ;
        RECT 72.500 146.000 72.900 146.100 ;
        RECT 71.700 145.700 72.100 145.800 ;
        RECT 73.400 145.700 73.800 147.400 ;
        RECT 75.100 146.200 75.400 147.900 ;
        RECT 75.800 146.400 76.200 147.200 ;
        RECT 74.200 146.100 74.600 146.200 ;
        RECT 75.000 146.100 75.400 146.200 ;
        RECT 76.600 146.100 77.000 146.200 ;
        RECT 78.200 146.100 78.600 147.900 ;
        RECT 74.200 145.800 75.400 146.100 ;
        RECT 76.200 145.800 78.600 146.100 ;
        RECT 71.700 145.400 73.800 145.700 ;
        RECT 70.200 144.900 71.400 145.200 ;
        RECT 69.900 144.500 70.300 144.600 ;
        RECT 69.200 144.200 70.300 144.500 ;
        RECT 71.100 144.400 71.400 144.900 ;
        RECT 71.100 144.000 71.800 144.400 ;
        RECT 67.900 143.700 68.300 143.800 ;
        RECT 69.300 143.700 69.700 143.800 ;
        RECT 66.200 143.100 66.600 143.500 ;
        RECT 67.900 143.400 69.700 143.700 ;
        RECT 69.000 143.100 69.300 143.400 ;
        RECT 71.000 143.100 71.400 143.500 ;
        RECT 66.200 142.800 67.200 143.100 ;
        RECT 66.800 141.100 67.200 142.800 ;
        RECT 69.000 141.100 69.400 143.100 ;
        RECT 71.100 141.100 71.700 143.100 ;
        RECT 73.400 141.100 73.800 145.400 ;
        RECT 74.300 145.100 74.600 145.800 ;
        RECT 76.200 145.600 76.600 145.800 ;
        RECT 74.200 141.100 74.600 145.100 ;
        RECT 75.000 144.800 77.000 145.100 ;
        RECT 75.000 141.100 75.400 144.800 ;
        RECT 76.600 141.100 77.000 144.800 ;
        RECT 77.400 144.400 77.800 145.200 ;
        RECT 78.200 141.100 78.600 145.800 ;
        RECT 79.800 147.700 80.200 149.900 ;
        RECT 81.900 149.200 82.500 149.900 ;
        RECT 81.900 148.900 82.600 149.200 ;
        RECT 84.200 148.900 84.600 149.900 ;
        RECT 86.400 149.200 86.800 149.900 ;
        RECT 86.400 148.900 87.400 149.200 ;
        RECT 82.200 148.500 82.600 148.900 ;
        RECT 84.300 148.600 84.600 148.900 ;
        RECT 84.300 148.300 85.700 148.600 ;
        RECT 85.300 148.200 85.700 148.300 ;
        RECT 86.200 148.200 86.600 148.600 ;
        RECT 87.000 148.500 87.400 148.900 ;
        RECT 81.300 147.700 81.700 147.800 ;
        RECT 79.800 147.400 81.700 147.700 ;
        RECT 79.800 145.700 80.200 147.400 ;
        RECT 86.200 147.200 86.500 148.200 ;
        RECT 88.600 147.500 89.000 149.900 ;
        RECT 90.200 147.600 90.600 149.900 ;
        RECT 91.800 147.600 92.200 149.900 ;
        RECT 93.400 147.600 93.800 149.900 ;
        RECT 95.000 147.600 95.400 149.900 ;
        RECT 90.200 147.200 91.100 147.600 ;
        RECT 91.800 147.200 92.900 147.600 ;
        RECT 93.400 147.200 94.500 147.600 ;
        RECT 95.000 147.200 96.200 147.600 ;
        RECT 98.200 147.500 98.600 149.900 ;
        RECT 100.400 149.200 100.800 149.900 ;
        RECT 99.800 148.900 100.800 149.200 ;
        RECT 102.600 148.900 103.000 149.900 ;
        RECT 104.700 149.200 105.300 149.900 ;
        RECT 104.600 148.900 105.300 149.200 ;
        RECT 99.800 148.500 100.200 148.900 ;
        RECT 102.600 148.600 102.900 148.900 ;
        RECT 100.600 148.200 101.000 148.600 ;
        RECT 101.500 148.300 102.900 148.600 ;
        RECT 104.600 148.500 105.000 148.900 ;
        RECT 101.500 148.200 101.900 148.300 ;
        RECT 83.300 147.100 83.700 147.200 ;
        RECT 86.200 147.100 86.600 147.200 ;
        RECT 87.800 147.100 88.600 147.200 ;
        RECT 83.100 146.800 88.600 147.100 ;
        RECT 89.400 146.900 89.800 147.200 ;
        RECT 90.700 146.900 91.100 147.200 ;
        RECT 92.500 146.900 92.900 147.200 ;
        RECT 94.100 146.900 94.500 147.200 ;
        RECT 82.200 146.400 82.600 146.500 ;
        RECT 80.700 146.100 82.600 146.400 ;
        RECT 80.700 146.000 81.100 146.100 ;
        RECT 81.500 145.700 81.900 145.800 ;
        RECT 79.800 145.400 81.900 145.700 ;
        RECT 79.800 141.100 80.200 145.400 ;
        RECT 83.100 145.200 83.400 146.800 ;
        RECT 86.700 146.700 87.100 146.800 ;
        RECT 89.400 146.500 90.300 146.900 ;
        RECT 90.700 146.500 92.000 146.900 ;
        RECT 92.500 146.500 93.700 146.900 ;
        RECT 94.100 146.500 95.400 146.900 ;
        RECT 87.500 146.200 87.900 146.300 ;
        RECT 85.400 145.900 87.900 146.200 ;
        RECT 85.400 145.800 85.800 145.900 ;
        RECT 90.700 145.800 91.100 146.500 ;
        RECT 92.500 145.800 92.900 146.500 ;
        RECT 94.100 145.800 94.500 146.500 ;
        RECT 95.800 145.800 96.200 147.200 ;
        RECT 98.600 147.100 99.400 147.200 ;
        RECT 100.700 147.100 101.000 148.200 ;
        RECT 105.500 147.700 105.900 147.800 ;
        RECT 107.000 147.700 107.400 149.900 ;
        RECT 105.500 147.400 107.400 147.700 ;
        RECT 107.800 147.500 108.200 149.900 ;
        RECT 110.000 149.200 110.400 149.900 ;
        RECT 109.400 148.900 110.400 149.200 ;
        RECT 112.200 148.900 112.600 149.900 ;
        RECT 114.300 149.200 114.900 149.900 ;
        RECT 114.200 148.900 114.900 149.200 ;
        RECT 109.400 148.500 109.800 148.900 ;
        RECT 112.200 148.600 112.500 148.900 ;
        RECT 110.200 148.200 110.600 148.600 ;
        RECT 111.100 148.300 112.500 148.600 ;
        RECT 114.200 148.500 114.600 148.900 ;
        RECT 111.100 148.200 111.500 148.300 ;
        RECT 103.500 147.100 103.900 147.200 ;
        RECT 98.600 146.800 104.100 147.100 ;
        RECT 100.100 146.700 100.500 146.800 ;
        RECT 99.300 146.200 99.700 146.300 ;
        RECT 100.600 146.200 101.000 146.300 ;
        RECT 99.300 145.900 101.800 146.200 ;
        RECT 101.400 145.800 101.800 145.900 ;
        RECT 86.200 145.500 89.000 145.600 ;
        RECT 86.100 145.400 89.000 145.500 ;
        RECT 82.200 144.900 83.400 145.200 ;
        RECT 84.100 145.300 89.000 145.400 ;
        RECT 84.100 145.100 86.500 145.300 ;
        RECT 82.200 144.400 82.500 144.900 ;
        RECT 81.800 144.000 82.500 144.400 ;
        RECT 83.300 144.500 83.700 144.600 ;
        RECT 84.100 144.500 84.400 145.100 ;
        RECT 83.300 144.200 84.400 144.500 ;
        RECT 84.700 144.500 87.400 144.800 ;
        RECT 84.700 144.400 85.100 144.500 ;
        RECT 87.000 144.400 87.400 144.500 ;
        RECT 83.900 143.700 84.300 143.800 ;
        RECT 85.300 143.700 85.700 143.800 ;
        RECT 82.200 143.100 82.600 143.500 ;
        RECT 83.900 143.400 85.700 143.700 ;
        RECT 84.300 143.100 84.600 143.400 ;
        RECT 87.000 143.100 87.400 143.500 ;
        RECT 81.900 141.100 82.500 143.100 ;
        RECT 84.200 141.100 84.600 143.100 ;
        RECT 86.400 142.800 87.400 143.100 ;
        RECT 86.400 141.100 86.800 142.800 ;
        RECT 88.600 141.100 89.000 145.300 ;
        RECT 90.200 145.400 91.100 145.800 ;
        RECT 91.800 145.400 92.900 145.800 ;
        RECT 93.400 145.400 94.500 145.800 ;
        RECT 95.000 145.400 96.200 145.800 ;
        RECT 98.200 145.500 101.000 145.600 ;
        RECT 98.200 145.400 101.100 145.500 ;
        RECT 90.200 141.100 90.600 145.400 ;
        RECT 91.800 141.100 92.200 145.400 ;
        RECT 93.400 141.100 93.800 145.400 ;
        RECT 95.000 141.100 95.400 145.400 ;
        RECT 98.200 145.300 103.100 145.400 ;
        RECT 98.200 141.100 98.600 145.300 ;
        RECT 100.700 145.100 103.100 145.300 ;
        RECT 99.800 144.500 102.500 144.800 ;
        RECT 99.800 144.400 100.200 144.500 ;
        RECT 102.100 144.400 102.500 144.500 ;
        RECT 102.800 144.500 103.100 145.100 ;
        RECT 103.800 145.200 104.100 146.800 ;
        RECT 104.600 146.400 105.000 146.500 ;
        RECT 104.600 146.100 106.500 146.400 ;
        RECT 106.100 146.000 106.500 146.100 ;
        RECT 105.300 145.700 105.700 145.800 ;
        RECT 107.000 145.700 107.400 147.400 ;
        RECT 108.200 147.100 109.000 147.200 ;
        RECT 110.300 147.100 110.600 148.200 ;
        RECT 115.100 147.700 115.500 147.800 ;
        RECT 116.600 147.700 117.000 149.900 ;
        RECT 115.100 147.400 117.000 147.700 ;
        RECT 113.100 147.100 113.500 147.200 ;
        RECT 108.200 146.800 113.700 147.100 ;
        RECT 109.700 146.700 110.100 146.800 ;
        RECT 108.900 146.200 109.300 146.300 ;
        RECT 110.200 146.200 110.600 146.300 ;
        RECT 108.900 145.900 111.400 146.200 ;
        RECT 111.000 145.800 111.400 145.900 ;
        RECT 105.300 145.400 107.400 145.700 ;
        RECT 103.800 144.900 105.000 145.200 ;
        RECT 103.500 144.500 103.900 144.600 ;
        RECT 102.800 144.200 103.900 144.500 ;
        RECT 104.700 144.400 105.000 144.900 ;
        RECT 104.700 144.000 105.400 144.400 ;
        RECT 101.500 143.700 101.900 143.800 ;
        RECT 102.900 143.700 103.300 143.800 ;
        RECT 99.800 143.100 100.200 143.500 ;
        RECT 101.500 143.400 103.300 143.700 ;
        RECT 102.600 143.100 102.900 143.400 ;
        RECT 104.600 143.100 105.000 143.500 ;
        RECT 99.800 142.800 100.800 143.100 ;
        RECT 100.400 141.100 100.800 142.800 ;
        RECT 102.600 141.100 103.000 143.100 ;
        RECT 104.700 141.100 105.300 143.100 ;
        RECT 107.000 141.100 107.400 145.400 ;
        RECT 107.800 145.500 110.600 145.600 ;
        RECT 107.800 145.400 110.700 145.500 ;
        RECT 107.800 145.300 112.700 145.400 ;
        RECT 107.800 141.100 108.200 145.300 ;
        RECT 110.300 145.100 112.700 145.300 ;
        RECT 109.400 144.500 112.100 144.800 ;
        RECT 109.400 144.400 109.800 144.500 ;
        RECT 111.700 144.400 112.100 144.500 ;
        RECT 112.400 144.500 112.700 145.100 ;
        RECT 113.400 145.200 113.700 146.800 ;
        RECT 114.200 146.400 114.600 146.500 ;
        RECT 114.200 146.100 116.100 146.400 ;
        RECT 115.700 146.000 116.100 146.100 ;
        RECT 114.900 145.700 115.300 145.800 ;
        RECT 116.600 145.700 117.000 147.400 ;
        RECT 117.400 148.500 117.800 149.500 ;
        RECT 117.400 147.400 117.700 148.500 ;
        RECT 119.500 148.000 119.900 149.500 ;
        RECT 119.500 147.700 120.300 148.000 ;
        RECT 119.900 147.500 120.300 147.700 ;
        RECT 122.200 147.500 122.600 149.900 ;
        RECT 124.400 149.200 124.800 149.900 ;
        RECT 123.800 148.900 124.800 149.200 ;
        RECT 126.600 148.900 127.000 149.900 ;
        RECT 128.700 149.200 129.300 149.900 ;
        RECT 128.600 148.900 129.300 149.200 ;
        RECT 123.800 148.500 124.200 148.900 ;
        RECT 126.600 148.600 126.900 148.900 ;
        RECT 124.600 148.200 125.000 148.600 ;
        RECT 125.500 148.300 126.900 148.600 ;
        RECT 128.600 148.500 129.000 148.900 ;
        RECT 125.500 148.200 125.900 148.300 ;
        RECT 117.400 147.100 119.500 147.400 ;
        RECT 119.000 146.900 119.500 147.100 ;
        RECT 120.000 147.200 120.300 147.500 ;
        RECT 117.400 145.800 117.800 146.600 ;
        RECT 118.200 145.800 118.600 146.600 ;
        RECT 119.000 146.500 119.700 146.900 ;
        RECT 120.000 146.800 121.000 147.200 ;
        RECT 122.600 147.100 123.400 147.200 ;
        RECT 124.700 147.100 125.000 148.200 ;
        RECT 129.500 147.700 129.900 147.800 ;
        RECT 131.000 147.700 131.400 149.900 ;
        RECT 133.700 148.000 134.100 149.500 ;
        RECT 135.800 148.500 136.200 149.500 ;
        RECT 129.500 147.400 131.400 147.700 ;
        RECT 127.500 147.100 127.900 147.200 ;
        RECT 122.600 146.800 128.100 147.100 ;
        RECT 114.900 145.400 117.000 145.700 ;
        RECT 119.000 145.500 119.300 146.500 ;
        RECT 113.400 144.900 114.600 145.200 ;
        RECT 113.100 144.500 113.500 144.600 ;
        RECT 112.400 144.200 113.500 144.500 ;
        RECT 114.300 144.400 114.600 144.900 ;
        RECT 114.300 144.000 115.000 144.400 ;
        RECT 111.100 143.700 111.500 143.800 ;
        RECT 112.500 143.700 112.900 143.800 ;
        RECT 109.400 143.100 109.800 143.500 ;
        RECT 111.100 143.400 112.900 143.700 ;
        RECT 112.200 143.100 112.500 143.400 ;
        RECT 114.200 143.100 114.600 143.500 ;
        RECT 109.400 142.800 110.400 143.100 ;
        RECT 110.000 141.100 110.400 142.800 ;
        RECT 112.200 141.100 112.600 143.100 ;
        RECT 114.300 141.100 114.900 143.100 ;
        RECT 116.600 141.100 117.000 145.400 ;
        RECT 117.400 145.200 119.300 145.500 ;
        RECT 117.400 143.500 117.700 145.200 ;
        RECT 120.000 144.900 120.300 146.800 ;
        RECT 124.100 146.700 124.500 146.800 ;
        RECT 123.300 146.200 123.700 146.300 ;
        RECT 124.600 146.200 125.000 146.300 ;
        RECT 120.600 146.100 121.000 146.200 ;
        RECT 121.400 146.100 121.800 146.200 ;
        RECT 120.600 145.800 121.800 146.100 ;
        RECT 123.300 145.900 125.800 146.200 ;
        RECT 125.400 145.800 125.800 145.900 ;
        RECT 120.600 145.400 121.000 145.800 ;
        RECT 122.200 145.500 125.000 145.600 ;
        RECT 122.200 145.400 125.100 145.500 ;
        RECT 119.500 144.600 120.300 144.900 ;
        RECT 122.200 145.300 127.100 145.400 ;
        RECT 117.400 141.500 117.800 143.500 ;
        RECT 119.500 142.200 119.900 144.600 ;
        RECT 119.000 141.800 119.900 142.200 ;
        RECT 119.500 141.100 119.900 141.800 ;
        RECT 122.200 141.100 122.600 145.300 ;
        RECT 124.700 145.100 127.100 145.300 ;
        RECT 123.800 144.500 126.500 144.800 ;
        RECT 123.800 144.400 124.200 144.500 ;
        RECT 126.100 144.400 126.500 144.500 ;
        RECT 126.800 144.500 127.100 145.100 ;
        RECT 127.800 145.200 128.100 146.800 ;
        RECT 128.600 146.400 129.000 146.500 ;
        RECT 128.600 146.100 130.500 146.400 ;
        RECT 130.100 146.000 130.500 146.100 ;
        RECT 129.300 145.700 129.700 145.800 ;
        RECT 131.000 145.700 131.400 147.400 ;
        RECT 133.300 147.700 134.100 148.000 ;
        RECT 133.300 147.500 133.700 147.700 ;
        RECT 133.300 147.200 133.600 147.500 ;
        RECT 135.900 147.400 136.200 148.500 ;
        RECT 132.600 146.800 133.600 147.200 ;
        RECT 134.100 147.100 136.200 147.400 ;
        RECT 136.600 147.700 137.000 149.900 ;
        RECT 138.700 149.200 139.300 149.900 ;
        RECT 138.700 148.900 139.400 149.200 ;
        RECT 141.000 148.900 141.400 149.900 ;
        RECT 143.200 149.200 143.600 149.900 ;
        RECT 143.200 148.900 144.200 149.200 ;
        RECT 139.000 148.500 139.400 148.900 ;
        RECT 141.100 148.600 141.400 148.900 ;
        RECT 141.100 148.300 142.500 148.600 ;
        RECT 142.100 148.200 142.500 148.300 ;
        RECT 143.000 148.200 143.400 148.600 ;
        RECT 143.800 148.500 144.200 148.900 ;
        RECT 138.100 147.700 138.500 147.800 ;
        RECT 136.600 147.400 138.500 147.700 ;
        RECT 134.100 146.900 134.600 147.100 ;
        RECT 129.300 145.400 131.400 145.700 ;
        RECT 132.600 145.400 133.000 146.200 ;
        RECT 127.800 144.900 129.000 145.200 ;
        RECT 127.500 144.500 127.900 144.600 ;
        RECT 126.800 144.200 127.900 144.500 ;
        RECT 128.700 144.400 129.000 144.900 ;
        RECT 128.700 144.000 129.400 144.400 ;
        RECT 125.500 143.700 125.900 143.800 ;
        RECT 126.900 143.700 127.300 143.800 ;
        RECT 123.800 143.100 124.200 143.500 ;
        RECT 125.500 143.400 127.300 143.700 ;
        RECT 126.600 143.100 126.900 143.400 ;
        RECT 128.600 143.100 129.000 143.500 ;
        RECT 123.800 142.800 124.800 143.100 ;
        RECT 124.400 141.100 124.800 142.800 ;
        RECT 126.600 141.100 127.000 143.100 ;
        RECT 128.700 141.100 129.300 143.100 ;
        RECT 131.000 141.100 131.400 145.400 ;
        RECT 133.300 144.900 133.600 146.800 ;
        RECT 133.900 146.500 134.600 146.900 ;
        RECT 134.300 145.500 134.600 146.500 ;
        RECT 135.000 145.800 135.400 146.600 ;
        RECT 135.800 145.800 136.200 146.600 ;
        RECT 136.600 145.700 137.000 147.400 ;
        RECT 140.100 147.100 140.500 147.200 ;
        RECT 143.000 147.100 143.300 148.200 ;
        RECT 145.400 147.500 145.800 149.900 ;
        RECT 146.200 148.000 146.600 149.900 ;
        RECT 147.800 148.000 148.200 149.900 ;
        RECT 146.200 147.900 148.200 148.000 ;
        RECT 148.600 147.900 149.000 149.900 ;
        RECT 150.700 148.200 151.100 149.900 ;
        RECT 150.200 147.900 151.100 148.200 ;
        RECT 153.400 147.900 153.800 149.900 ;
        RECT 154.200 148.000 154.600 149.900 ;
        RECT 155.800 148.000 156.200 149.900 ;
        RECT 154.200 147.900 156.200 148.000 ;
        RECT 156.600 148.000 157.000 149.900 ;
        RECT 158.200 148.000 158.600 149.900 ;
        RECT 156.600 147.900 158.600 148.000 ;
        RECT 159.000 147.900 159.400 149.900 ;
        RECT 160.100 148.200 160.500 149.900 ;
        RECT 160.100 147.900 161.000 148.200 ;
        RECT 146.300 147.700 148.100 147.900 ;
        RECT 146.600 147.200 147.000 147.400 ;
        RECT 148.600 147.200 148.900 147.900 ;
        RECT 144.600 147.100 145.400 147.200 ;
        RECT 139.900 146.800 145.400 147.100 ;
        RECT 146.200 146.900 147.000 147.200 ;
        RECT 146.200 146.800 146.600 146.900 ;
        RECT 147.700 146.800 149.000 147.200 ;
        RECT 149.400 146.800 149.800 147.600 ;
        RECT 139.000 146.400 139.400 146.500 ;
        RECT 137.500 146.100 139.400 146.400 ;
        RECT 139.900 146.200 140.200 146.800 ;
        RECT 143.500 146.700 143.900 146.800 ;
        RECT 143.000 146.200 143.400 146.300 ;
        RECT 144.300 146.200 144.700 146.300 ;
        RECT 137.500 146.000 137.900 146.100 ;
        RECT 139.800 145.800 140.200 146.200 ;
        RECT 142.200 145.900 144.700 146.200 ;
        RECT 142.200 145.800 142.600 145.900 ;
        RECT 147.000 145.800 147.400 146.600 ;
        RECT 138.300 145.700 138.700 145.800 ;
        RECT 134.300 145.200 136.200 145.500 ;
        RECT 133.300 144.600 134.100 144.900 ;
        RECT 133.700 142.200 134.100 144.600 ;
        RECT 135.900 143.500 136.200 145.200 ;
        RECT 133.400 141.800 134.100 142.200 ;
        RECT 133.700 141.100 134.100 141.800 ;
        RECT 135.800 141.500 136.200 143.500 ;
        RECT 136.600 145.400 138.700 145.700 ;
        RECT 136.600 141.100 137.000 145.400 ;
        RECT 139.900 145.200 140.200 145.800 ;
        RECT 143.000 145.500 145.800 145.600 ;
        RECT 142.900 145.400 145.800 145.500 ;
        RECT 139.000 144.900 140.200 145.200 ;
        RECT 140.900 145.300 145.800 145.400 ;
        RECT 140.900 145.100 143.300 145.300 ;
        RECT 139.000 144.400 139.300 144.900 ;
        RECT 138.600 144.000 139.300 144.400 ;
        RECT 140.100 144.500 140.500 144.600 ;
        RECT 140.900 144.500 141.200 145.100 ;
        RECT 140.100 144.200 141.200 144.500 ;
        RECT 141.500 144.500 144.200 144.800 ;
        RECT 141.500 144.400 141.900 144.500 ;
        RECT 143.800 144.400 144.200 144.500 ;
        RECT 140.700 143.700 141.100 143.800 ;
        RECT 142.100 143.700 142.500 143.800 ;
        RECT 139.000 143.100 139.400 143.500 ;
        RECT 140.700 143.400 142.500 143.700 ;
        RECT 141.100 143.100 141.400 143.400 ;
        RECT 143.800 143.100 144.200 143.500 ;
        RECT 138.700 141.100 139.300 143.100 ;
        RECT 141.000 141.100 141.400 143.100 ;
        RECT 143.200 142.800 144.200 143.100 ;
        RECT 143.200 141.100 143.600 142.800 ;
        RECT 145.400 141.100 145.800 145.300 ;
        RECT 147.700 145.100 148.000 146.800 ;
        RECT 148.600 146.200 148.900 146.800 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 148.600 145.100 149.000 145.200 ;
        RECT 150.200 145.100 150.600 147.900 ;
        RECT 153.500 147.200 153.800 147.900 ;
        RECT 154.300 147.700 156.100 147.900 ;
        RECT 156.700 147.700 158.500 147.900 ;
        RECT 155.400 147.200 155.800 147.400 ;
        RECT 157.000 147.200 157.400 147.400 ;
        RECT 159.000 147.200 159.300 147.900 ;
        RECT 153.400 146.800 154.700 147.200 ;
        RECT 155.400 146.900 156.200 147.200 ;
        RECT 155.800 146.800 156.200 146.900 ;
        RECT 156.600 146.900 157.400 147.200 ;
        RECT 158.100 147.100 159.400 147.200 ;
        RECT 159.800 147.100 160.200 147.200 ;
        RECT 156.600 146.800 157.000 146.900 ;
        RECT 158.100 146.800 160.200 147.100 ;
        RECT 147.500 144.800 148.000 145.100 ;
        RECT 148.300 144.800 150.600 145.100 ;
        RECT 147.500 141.100 147.900 144.800 ;
        RECT 148.300 144.200 148.600 144.800 ;
        RECT 148.200 143.800 148.600 144.200 ;
        RECT 150.200 141.100 150.600 144.800 ;
        RECT 151.000 144.400 151.400 145.200 ;
        RECT 153.400 145.100 153.800 145.200 ;
        RECT 154.400 145.100 154.700 146.800 ;
        RECT 155.000 145.800 155.400 146.600 ;
        RECT 155.800 146.100 156.200 146.200 ;
        RECT 157.400 146.100 157.800 146.600 ;
        RECT 155.800 145.800 157.800 146.100 ;
        RECT 158.100 145.100 158.400 146.800 ;
        RECT 160.600 146.100 161.000 147.900 ;
        RECT 161.400 146.800 161.800 147.600 ;
        RECT 162.200 147.500 162.600 149.900 ;
        RECT 164.400 149.200 164.800 149.900 ;
        RECT 163.800 148.900 164.800 149.200 ;
        RECT 166.600 148.900 167.000 149.900 ;
        RECT 168.700 149.200 169.300 149.900 ;
        RECT 168.600 148.900 169.300 149.200 ;
        RECT 163.800 148.500 164.200 148.900 ;
        RECT 166.600 148.600 166.900 148.900 ;
        RECT 164.600 148.200 165.000 148.600 ;
        RECT 165.500 148.300 166.900 148.600 ;
        RECT 168.600 148.500 169.000 148.900 ;
        RECT 165.500 148.200 165.900 148.300 ;
        RECT 162.600 147.100 163.400 147.200 ;
        RECT 164.700 147.100 165.000 148.200 ;
        RECT 169.500 147.700 169.900 147.800 ;
        RECT 171.000 147.700 171.400 149.900 ;
        RECT 171.800 147.900 172.200 149.900 ;
        RECT 172.600 148.000 173.000 149.900 ;
        RECT 174.200 148.000 174.600 149.900 ;
        RECT 172.600 147.900 174.600 148.000 ;
        RECT 169.500 147.400 171.400 147.700 ;
        RECT 167.500 147.100 167.900 147.200 ;
        RECT 162.600 146.800 168.100 147.100 ;
        RECT 164.100 146.700 164.500 146.800 ;
        RECT 159.000 145.800 161.000 146.100 ;
        RECT 163.300 146.200 163.700 146.300 ;
        RECT 164.600 146.200 165.000 146.300 ;
        RECT 167.800 146.200 168.100 146.800 ;
        RECT 168.600 146.400 169.000 146.500 ;
        RECT 163.300 145.900 165.800 146.200 ;
        RECT 165.400 145.800 165.800 145.900 ;
        RECT 167.800 145.800 168.200 146.200 ;
        RECT 168.600 146.100 170.500 146.400 ;
        RECT 170.100 146.000 170.500 146.100 ;
        RECT 159.000 145.200 159.300 145.800 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 153.400 144.800 154.100 145.100 ;
        RECT 154.400 144.800 154.900 145.100 ;
        RECT 153.800 144.200 154.100 144.800 ;
        RECT 153.800 143.800 154.200 144.200 ;
        RECT 154.500 141.100 154.900 144.800 ;
        RECT 157.900 144.800 158.400 145.100 ;
        RECT 158.700 144.800 159.400 145.100 ;
        RECT 157.900 141.100 158.300 144.800 ;
        RECT 158.700 144.200 159.000 144.800 ;
        RECT 159.800 144.400 160.200 145.200 ;
        RECT 158.600 143.800 159.000 144.200 ;
        RECT 160.600 141.100 161.000 145.800 ;
        RECT 162.200 145.500 165.000 145.600 ;
        RECT 162.200 145.400 165.100 145.500 ;
        RECT 162.200 145.300 167.100 145.400 ;
        RECT 162.200 141.100 162.600 145.300 ;
        RECT 164.700 145.100 167.100 145.300 ;
        RECT 163.800 144.500 166.500 144.800 ;
        RECT 163.800 144.400 164.200 144.500 ;
        RECT 166.100 144.400 166.500 144.500 ;
        RECT 166.800 144.500 167.100 145.100 ;
        RECT 167.800 145.200 168.100 145.800 ;
        RECT 169.300 145.700 169.700 145.800 ;
        RECT 171.000 145.700 171.400 147.400 ;
        RECT 171.900 147.200 172.200 147.900 ;
        RECT 172.700 147.700 174.500 147.900 ;
        RECT 175.000 147.700 175.400 149.900 ;
        RECT 177.100 149.200 177.700 149.900 ;
        RECT 177.100 148.900 177.800 149.200 ;
        RECT 179.400 148.900 179.800 149.900 ;
        RECT 181.600 149.200 182.000 149.900 ;
        RECT 181.600 148.900 182.600 149.200 ;
        RECT 177.400 148.500 177.800 148.900 ;
        RECT 179.500 148.600 179.800 148.900 ;
        RECT 179.500 148.300 180.900 148.600 ;
        RECT 180.500 148.200 180.900 148.300 ;
        RECT 181.400 148.200 181.800 148.600 ;
        RECT 182.200 148.500 182.600 148.900 ;
        RECT 176.500 147.700 176.900 147.800 ;
        RECT 175.000 147.400 176.900 147.700 ;
        RECT 173.800 147.200 174.200 147.400 ;
        RECT 171.800 146.800 173.100 147.200 ;
        RECT 173.800 146.900 174.600 147.200 ;
        RECT 174.200 146.800 174.600 146.900 ;
        RECT 172.800 146.200 173.100 146.800 ;
        RECT 172.600 145.800 173.100 146.200 ;
        RECT 173.400 145.800 173.800 146.600 ;
        RECT 169.300 145.400 171.400 145.700 ;
        RECT 167.800 144.900 169.000 145.200 ;
        RECT 167.500 144.500 167.900 144.600 ;
        RECT 166.800 144.200 167.900 144.500 ;
        RECT 168.700 144.400 169.000 144.900 ;
        RECT 168.700 144.000 169.400 144.400 ;
        RECT 165.500 143.700 165.900 143.800 ;
        RECT 166.900 143.700 167.300 143.800 ;
        RECT 163.800 143.100 164.200 143.500 ;
        RECT 165.500 143.400 167.300 143.700 ;
        RECT 166.600 143.100 166.900 143.400 ;
        RECT 168.600 143.100 169.000 143.500 ;
        RECT 163.800 142.800 164.800 143.100 ;
        RECT 164.400 141.100 164.800 142.800 ;
        RECT 166.600 141.100 167.000 143.100 ;
        RECT 168.700 141.100 169.300 143.100 ;
        RECT 171.000 141.100 171.400 145.400 ;
        RECT 171.800 145.100 172.200 145.200 ;
        RECT 172.800 145.100 173.100 145.800 ;
        RECT 175.000 145.700 175.400 147.400 ;
        RECT 178.500 147.100 179.400 147.200 ;
        RECT 181.400 147.100 181.700 148.200 ;
        RECT 183.800 147.500 184.200 149.900 ;
        RECT 185.400 147.600 185.800 149.900 ;
        RECT 187.000 147.600 187.400 149.900 ;
        RECT 188.600 147.600 189.000 149.900 ;
        RECT 190.200 147.600 190.600 149.900 ;
        RECT 184.600 147.200 185.800 147.600 ;
        RECT 186.300 147.200 187.400 147.600 ;
        RECT 187.900 147.200 189.000 147.600 ;
        RECT 189.700 147.200 190.600 147.600 ;
        RECT 191.800 148.500 192.200 149.500 ;
        RECT 191.800 147.400 192.100 148.500 ;
        RECT 193.900 148.000 194.300 149.500 ;
        RECT 196.600 148.000 197.000 149.900 ;
        RECT 198.200 148.000 198.600 149.900 ;
        RECT 193.900 147.700 194.700 148.000 ;
        RECT 196.600 147.900 198.600 148.000 ;
        RECT 199.000 147.900 199.400 149.900 ;
        RECT 200.100 148.200 200.500 149.900 ;
        RECT 203.800 148.500 204.200 149.500 ;
        RECT 200.100 147.900 201.000 148.200 ;
        RECT 196.700 147.700 198.500 147.900 ;
        RECT 194.300 147.500 194.700 147.700 ;
        RECT 183.000 147.100 183.800 147.200 ;
        RECT 178.300 146.800 183.800 147.100 ;
        RECT 177.400 146.400 177.800 146.500 ;
        RECT 175.900 146.100 177.800 146.400 ;
        RECT 175.900 146.000 176.300 146.100 ;
        RECT 176.700 145.700 177.100 145.800 ;
        RECT 175.000 145.400 177.100 145.700 ;
        RECT 171.800 144.800 172.500 145.100 ;
        RECT 172.800 144.800 173.300 145.100 ;
        RECT 172.200 144.200 172.500 144.800 ;
        RECT 172.200 143.800 172.600 144.200 ;
        RECT 172.900 141.100 173.300 144.800 ;
        RECT 175.000 141.100 175.400 145.400 ;
        RECT 178.300 145.200 178.600 146.800 ;
        RECT 181.900 146.700 182.300 146.800 ;
        RECT 182.700 146.200 183.100 146.300 ;
        RECT 179.800 146.100 180.200 146.200 ;
        RECT 180.600 146.100 183.100 146.200 ;
        RECT 179.800 145.900 183.100 146.100 ;
        RECT 179.800 145.800 181.000 145.900 ;
        RECT 184.600 145.800 185.000 147.200 ;
        RECT 186.300 146.900 186.700 147.200 ;
        RECT 187.900 146.900 188.300 147.200 ;
        RECT 189.700 146.900 190.100 147.200 ;
        RECT 191.800 147.100 193.900 147.400 ;
        RECT 185.400 146.500 186.700 146.900 ;
        RECT 187.100 146.500 188.300 146.900 ;
        RECT 188.800 146.500 190.100 146.900 ;
        RECT 193.400 146.900 193.900 147.100 ;
        RECT 194.400 147.200 194.700 147.500 ;
        RECT 197.000 147.200 197.400 147.400 ;
        RECT 199.000 147.200 199.300 147.900 ;
        RECT 186.300 145.800 186.700 146.500 ;
        RECT 187.900 145.800 188.300 146.500 ;
        RECT 189.700 145.800 190.100 146.500 ;
        RECT 191.800 145.800 192.200 146.600 ;
        RECT 192.600 145.800 193.000 146.600 ;
        RECT 193.400 146.500 194.100 146.900 ;
        RECT 194.400 146.800 195.400 147.200 ;
        RECT 195.800 147.100 196.200 147.200 ;
        RECT 196.600 147.100 197.400 147.200 ;
        RECT 195.800 146.900 197.400 147.100 ;
        RECT 198.100 147.100 199.400 147.200 ;
        RECT 199.800 147.100 200.200 147.200 ;
        RECT 195.800 146.800 197.000 146.900 ;
        RECT 198.100 146.800 200.200 147.100 ;
        RECT 181.400 145.500 184.200 145.600 ;
        RECT 181.300 145.400 184.200 145.500 ;
        RECT 184.600 145.400 185.800 145.800 ;
        RECT 186.300 145.400 187.400 145.800 ;
        RECT 187.900 145.400 189.000 145.800 ;
        RECT 189.700 145.400 190.600 145.800 ;
        RECT 193.400 145.500 193.700 146.500 ;
        RECT 177.400 144.900 178.600 145.200 ;
        RECT 179.300 145.300 184.200 145.400 ;
        RECT 179.300 145.100 181.700 145.300 ;
        RECT 177.400 144.400 177.700 144.900 ;
        RECT 177.000 144.000 177.700 144.400 ;
        RECT 178.500 144.500 178.900 144.600 ;
        RECT 179.300 144.500 179.600 145.100 ;
        RECT 178.500 144.200 179.600 144.500 ;
        RECT 179.900 144.500 182.600 144.800 ;
        RECT 179.900 144.400 180.300 144.500 ;
        RECT 182.200 144.400 182.600 144.500 ;
        RECT 179.100 143.700 179.500 143.800 ;
        RECT 180.500 143.700 180.900 143.800 ;
        RECT 177.400 143.100 177.800 143.500 ;
        RECT 179.100 143.400 180.900 143.700 ;
        RECT 179.500 143.100 179.800 143.400 ;
        RECT 182.200 143.100 182.600 143.500 ;
        RECT 177.100 141.100 177.700 143.100 ;
        RECT 179.400 141.100 179.800 143.100 ;
        RECT 181.600 142.800 182.600 143.100 ;
        RECT 181.600 141.100 182.000 142.800 ;
        RECT 183.800 141.100 184.200 145.300 ;
        RECT 185.400 141.100 185.800 145.400 ;
        RECT 187.000 141.100 187.400 145.400 ;
        RECT 188.600 141.100 189.000 145.400 ;
        RECT 190.200 141.100 190.600 145.400 ;
        RECT 191.800 145.200 193.700 145.500 ;
        RECT 191.800 143.500 192.100 145.200 ;
        RECT 194.400 144.900 194.700 146.800 ;
        RECT 195.000 145.400 195.400 146.200 ;
        RECT 197.400 145.800 197.800 146.600 ;
        RECT 198.100 145.100 198.400 146.800 ;
        RECT 200.600 146.100 201.000 147.900 ;
        RECT 201.400 147.100 201.800 147.600 ;
        RECT 203.800 147.400 204.100 148.500 ;
        RECT 205.900 148.200 206.300 149.500 ;
        RECT 205.400 148.000 206.300 148.200 ;
        RECT 205.400 147.800 206.700 148.000 ;
        RECT 205.900 147.700 206.700 147.800 ;
        RECT 206.300 147.500 206.700 147.700 ;
        RECT 202.200 147.100 202.600 147.200 ;
        RECT 203.800 147.100 205.900 147.400 ;
        RECT 201.400 146.800 202.600 147.100 ;
        RECT 205.400 146.900 205.900 147.100 ;
        RECT 206.400 147.200 206.700 147.500 ;
        RECT 208.600 147.700 209.000 149.900 ;
        RECT 210.700 149.200 211.300 149.900 ;
        RECT 210.700 148.900 211.400 149.200 ;
        RECT 213.000 148.900 213.400 149.900 ;
        RECT 215.200 149.200 215.600 149.900 ;
        RECT 215.200 148.900 216.200 149.200 ;
        RECT 211.000 148.500 211.400 148.900 ;
        RECT 213.100 148.600 213.400 148.900 ;
        RECT 213.100 148.300 214.500 148.600 ;
        RECT 214.100 148.200 214.500 148.300 ;
        RECT 215.000 148.200 215.400 148.600 ;
        RECT 215.800 148.500 216.200 148.900 ;
        RECT 210.100 147.700 210.500 147.800 ;
        RECT 208.600 147.400 210.500 147.700 ;
        RECT 199.000 145.800 201.000 146.100 ;
        RECT 203.800 145.800 204.200 146.600 ;
        RECT 204.600 145.800 205.000 146.600 ;
        RECT 205.400 146.500 206.100 146.900 ;
        RECT 206.400 146.800 207.400 147.200 ;
        RECT 199.000 145.200 199.300 145.800 ;
        RECT 199.000 145.100 199.400 145.200 ;
        RECT 193.900 144.600 194.700 144.900 ;
        RECT 197.900 144.800 198.400 145.100 ;
        RECT 198.700 144.800 199.400 145.100 ;
        RECT 191.800 141.500 192.200 143.500 ;
        RECT 193.900 142.200 194.300 144.600 ;
        RECT 193.400 141.800 194.300 142.200 ;
        RECT 193.900 141.100 194.300 141.800 ;
        RECT 197.900 141.100 198.300 144.800 ;
        RECT 198.700 144.200 199.000 144.800 ;
        RECT 199.800 144.400 200.200 145.200 ;
        RECT 198.600 143.800 199.000 144.200 ;
        RECT 200.600 141.100 201.000 145.800 ;
        RECT 205.400 145.500 205.700 146.500 ;
        RECT 203.800 145.200 205.700 145.500 ;
        RECT 203.800 143.500 204.100 145.200 ;
        RECT 206.400 144.900 206.700 146.800 ;
        RECT 207.000 145.400 207.400 146.200 ;
        RECT 208.600 145.700 209.000 147.400 ;
        RECT 212.100 147.100 212.500 147.200 ;
        RECT 215.000 147.100 215.300 148.200 ;
        RECT 217.400 147.500 217.800 149.900 ;
        RECT 220.100 149.200 220.500 149.500 ;
        RECT 219.800 148.800 220.500 149.200 ;
        RECT 220.100 148.000 220.500 148.800 ;
        RECT 222.200 148.500 222.600 149.500 ;
        RECT 219.700 147.700 220.500 148.000 ;
        RECT 219.700 147.500 220.100 147.700 ;
        RECT 219.700 147.200 220.000 147.500 ;
        RECT 222.300 147.400 222.600 148.500 ;
        RECT 224.300 148.200 224.700 149.900 ;
        RECT 223.800 147.900 224.700 148.200 ;
        RECT 225.400 147.900 225.800 149.900 ;
        RECT 226.200 148.000 226.600 149.900 ;
        RECT 227.800 148.000 228.200 149.900 ;
        RECT 226.200 147.900 228.200 148.000 ;
        RECT 216.600 147.100 217.400 147.200 ;
        RECT 211.900 146.800 217.400 147.100 ;
        RECT 219.000 146.800 220.000 147.200 ;
        RECT 220.500 147.100 222.600 147.400 ;
        RECT 220.500 146.900 221.000 147.100 ;
        RECT 211.000 146.400 211.400 146.500 ;
        RECT 209.500 146.100 211.400 146.400 ;
        RECT 209.500 146.000 209.900 146.100 ;
        RECT 210.300 145.700 210.700 145.800 ;
        RECT 208.600 145.400 210.700 145.700 ;
        RECT 205.900 144.600 206.700 144.900 ;
        RECT 203.800 141.500 204.200 143.500 ;
        RECT 205.900 141.100 206.300 144.600 ;
        RECT 208.600 141.100 209.000 145.400 ;
        RECT 211.900 145.200 212.200 146.800 ;
        RECT 215.500 146.700 215.900 146.800 ;
        RECT 216.300 146.200 216.700 146.300 ;
        RECT 214.200 145.900 216.700 146.200 ;
        RECT 214.200 145.800 214.600 145.900 ;
        RECT 215.000 145.500 217.800 145.600 ;
        RECT 214.900 145.400 217.800 145.500 ;
        RECT 219.000 145.400 219.400 146.200 ;
        RECT 211.000 144.900 212.200 145.200 ;
        RECT 212.900 145.300 217.800 145.400 ;
        RECT 212.900 145.100 215.300 145.300 ;
        RECT 211.000 144.400 211.300 144.900 ;
        RECT 210.600 144.000 211.300 144.400 ;
        RECT 212.100 144.500 212.500 144.600 ;
        RECT 212.900 144.500 213.200 145.100 ;
        RECT 212.100 144.200 213.200 144.500 ;
        RECT 213.500 144.500 216.200 144.800 ;
        RECT 213.500 144.400 213.900 144.500 ;
        RECT 215.800 144.400 216.200 144.500 ;
        RECT 212.700 143.700 213.100 143.800 ;
        RECT 214.100 143.700 214.500 143.800 ;
        RECT 211.000 143.100 211.400 143.500 ;
        RECT 212.700 143.400 214.500 143.700 ;
        RECT 213.100 143.100 213.400 143.400 ;
        RECT 215.800 143.100 216.200 143.500 ;
        RECT 210.700 141.100 211.300 143.100 ;
        RECT 213.000 141.100 213.400 143.100 ;
        RECT 215.200 142.800 216.200 143.100 ;
        RECT 215.200 141.100 215.600 142.800 ;
        RECT 217.400 141.100 217.800 145.300 ;
        RECT 219.700 144.900 220.000 146.800 ;
        RECT 220.300 146.500 221.000 146.900 ;
        RECT 223.000 146.800 223.400 147.600 ;
        RECT 220.700 145.500 221.000 146.500 ;
        RECT 221.400 145.800 221.800 146.600 ;
        RECT 222.200 145.800 222.600 146.600 ;
        RECT 223.000 146.200 223.300 146.800 ;
        RECT 223.000 145.800 223.400 146.200 ;
        RECT 223.800 146.100 224.200 147.900 ;
        RECT 225.500 147.200 225.800 147.900 ;
        RECT 226.300 147.700 228.100 147.900 ;
        RECT 228.600 147.700 229.000 149.900 ;
        RECT 230.700 149.200 231.300 149.900 ;
        RECT 230.700 148.900 231.400 149.200 ;
        RECT 233.000 148.900 233.400 149.900 ;
        RECT 235.200 149.200 235.600 149.900 ;
        RECT 235.200 148.900 236.200 149.200 ;
        RECT 231.000 148.500 231.400 148.900 ;
        RECT 233.100 148.600 233.400 148.900 ;
        RECT 233.100 148.300 234.500 148.600 ;
        RECT 234.100 148.200 234.500 148.300 ;
        RECT 235.000 148.200 235.400 148.600 ;
        RECT 235.800 148.500 236.200 148.900 ;
        RECT 230.100 147.700 230.500 147.800 ;
        RECT 228.600 147.400 230.500 147.700 ;
        RECT 227.400 147.200 227.800 147.400 ;
        RECT 225.400 146.800 226.700 147.200 ;
        RECT 227.400 146.900 228.200 147.200 ;
        RECT 227.800 146.800 228.200 146.900 ;
        RECT 223.800 145.800 225.700 146.100 ;
        RECT 220.700 145.200 222.600 145.500 ;
        RECT 219.700 144.600 220.500 144.900 ;
        RECT 220.100 141.100 220.500 144.600 ;
        RECT 222.300 143.500 222.600 145.200 ;
        RECT 222.200 141.500 222.600 143.500 ;
        RECT 223.800 141.100 224.200 145.800 ;
        RECT 225.400 145.200 225.700 145.800 ;
        RECT 226.400 145.200 226.700 146.800 ;
        RECT 227.000 146.100 227.400 146.600 ;
        RECT 227.800 146.100 228.200 146.200 ;
        RECT 227.000 145.800 228.200 146.100 ;
        RECT 228.600 145.700 229.000 147.400 ;
        RECT 231.800 147.100 232.500 147.200 ;
        RECT 235.000 147.100 235.300 148.200 ;
        RECT 237.400 147.500 237.800 149.900 ;
        RECT 238.200 148.000 238.600 149.900 ;
        RECT 239.800 148.000 240.200 149.900 ;
        RECT 238.200 147.900 240.200 148.000 ;
        RECT 240.600 147.900 241.000 149.900 ;
        RECT 238.300 147.700 240.100 147.900 ;
        RECT 238.600 147.200 239.000 147.400 ;
        RECT 240.600 147.200 240.900 147.900 ;
        RECT 241.400 147.500 241.800 149.900 ;
        RECT 243.600 149.200 244.000 149.900 ;
        RECT 243.000 148.900 244.000 149.200 ;
        RECT 245.800 148.900 246.200 149.900 ;
        RECT 247.900 149.200 248.500 149.900 ;
        RECT 247.800 148.900 248.500 149.200 ;
        RECT 243.000 148.500 243.400 148.900 ;
        RECT 245.800 148.600 246.100 148.900 ;
        RECT 243.800 148.200 244.200 148.600 ;
        RECT 244.700 148.300 246.100 148.600 ;
        RECT 247.800 148.500 248.200 148.900 ;
        RECT 244.700 148.200 245.100 148.300 ;
        RECT 243.900 147.200 244.200 148.200 ;
        RECT 248.700 147.700 249.100 147.800 ;
        RECT 250.200 147.700 250.600 149.900 ;
        RECT 248.700 147.400 250.600 147.700 ;
        RECT 236.600 147.100 237.400 147.200 ;
        RECT 231.800 146.800 237.400 147.100 ;
        RECT 238.200 146.900 239.000 147.200 ;
        RECT 238.200 146.800 238.600 146.900 ;
        RECT 239.700 146.800 241.000 147.200 ;
        RECT 241.800 147.100 242.600 147.200 ;
        RECT 243.800 147.100 244.200 147.200 ;
        RECT 246.700 147.100 247.100 147.200 ;
        RECT 241.800 146.800 247.300 147.100 ;
        RECT 231.000 146.400 231.400 146.500 ;
        RECT 229.500 146.100 231.400 146.400 ;
        RECT 229.500 146.000 229.900 146.100 ;
        RECT 230.300 145.700 230.700 145.800 ;
        RECT 228.600 145.400 230.700 145.700 ;
        RECT 224.600 144.400 225.000 145.200 ;
        RECT 225.400 145.100 225.800 145.200 ;
        RECT 225.400 144.800 226.100 145.100 ;
        RECT 226.400 144.800 227.400 145.200 ;
        RECT 225.800 144.200 226.100 144.800 ;
        RECT 225.800 143.800 226.200 144.200 ;
        RECT 226.500 141.100 226.900 144.800 ;
        RECT 228.600 141.100 229.000 145.400 ;
        RECT 231.900 145.200 232.200 146.800 ;
        RECT 235.500 146.700 235.900 146.800 ;
        RECT 236.300 146.200 236.700 146.300 ;
        RECT 234.200 145.900 236.700 146.200 ;
        RECT 234.200 145.800 234.600 145.900 ;
        RECT 239.000 145.800 239.400 146.600 ;
        RECT 235.000 145.500 237.800 145.600 ;
        RECT 234.900 145.400 237.800 145.500 ;
        RECT 231.000 144.900 232.200 145.200 ;
        RECT 232.900 145.300 237.800 145.400 ;
        RECT 232.900 145.100 235.300 145.300 ;
        RECT 231.000 144.400 231.300 144.900 ;
        RECT 230.600 144.000 231.300 144.400 ;
        RECT 232.100 144.500 232.500 144.600 ;
        RECT 232.900 144.500 233.200 145.100 ;
        RECT 232.100 144.200 233.200 144.500 ;
        RECT 233.500 144.500 236.200 144.800 ;
        RECT 233.500 144.400 233.900 144.500 ;
        RECT 235.800 144.400 236.200 144.500 ;
        RECT 232.700 143.700 233.100 143.800 ;
        RECT 234.100 143.700 234.500 143.800 ;
        RECT 231.000 143.100 231.400 143.500 ;
        RECT 232.700 143.400 234.500 143.700 ;
        RECT 233.100 143.100 233.400 143.400 ;
        RECT 235.800 143.100 236.200 143.500 ;
        RECT 230.700 141.100 231.300 143.100 ;
        RECT 233.000 141.100 233.400 143.100 ;
        RECT 235.200 142.800 236.200 143.100 ;
        RECT 235.200 141.100 235.600 142.800 ;
        RECT 237.400 141.100 237.800 145.300 ;
        RECT 239.700 145.100 240.000 146.800 ;
        RECT 243.300 146.700 243.700 146.800 ;
        RECT 242.500 146.200 242.900 146.300 ;
        RECT 242.500 145.900 245.000 146.200 ;
        RECT 244.600 145.800 245.000 145.900 ;
        RECT 241.400 145.500 244.200 145.600 ;
        RECT 241.400 145.400 244.300 145.500 ;
        RECT 241.400 145.300 246.300 145.400 ;
        RECT 240.600 145.100 241.000 145.200 ;
        RECT 239.500 144.800 240.000 145.100 ;
        RECT 240.300 144.800 241.000 145.100 ;
        RECT 239.500 141.100 239.900 144.800 ;
        RECT 240.300 144.200 240.600 144.800 ;
        RECT 240.200 143.800 240.600 144.200 ;
        RECT 241.400 141.100 241.800 145.300 ;
        RECT 243.900 145.100 246.300 145.300 ;
        RECT 243.000 144.500 245.700 144.800 ;
        RECT 243.000 144.400 243.400 144.500 ;
        RECT 245.300 144.400 245.700 144.500 ;
        RECT 246.000 144.500 246.300 145.100 ;
        RECT 247.000 145.200 247.300 146.800 ;
        RECT 247.800 146.400 248.200 146.500 ;
        RECT 247.800 146.100 249.700 146.400 ;
        RECT 249.300 146.000 249.700 146.100 ;
        RECT 248.500 145.700 248.900 145.800 ;
        RECT 250.200 145.700 250.600 147.400 ;
        RECT 248.500 145.400 250.600 145.700 ;
        RECT 247.000 144.900 248.200 145.200 ;
        RECT 246.700 144.500 247.100 144.600 ;
        RECT 246.000 144.200 247.100 144.500 ;
        RECT 247.900 144.400 248.200 144.900 ;
        RECT 247.900 144.000 248.600 144.400 ;
        RECT 244.700 143.700 245.100 143.800 ;
        RECT 246.100 143.700 246.500 143.800 ;
        RECT 243.000 143.100 243.400 143.500 ;
        RECT 244.700 143.400 246.500 143.700 ;
        RECT 245.800 143.100 246.100 143.400 ;
        RECT 247.800 143.100 248.200 143.500 ;
        RECT 243.000 142.800 244.000 143.100 ;
        RECT 243.600 141.100 244.000 142.800 ;
        RECT 245.800 141.100 246.200 143.100 ;
        RECT 247.900 141.100 248.500 143.100 ;
        RECT 250.200 141.100 250.600 145.400 ;
        RECT 1.400 135.600 1.800 139.900 ;
        RECT 3.000 135.600 3.400 139.900 ;
        RECT 1.400 135.200 3.400 135.600 ;
        RECT 4.600 135.700 5.000 139.900 ;
        RECT 6.800 138.200 7.200 139.900 ;
        RECT 6.200 137.900 7.200 138.200 ;
        RECT 9.000 137.900 9.400 139.900 ;
        RECT 11.100 137.900 11.700 139.900 ;
        RECT 6.200 137.500 6.600 137.900 ;
        RECT 9.000 137.600 9.300 137.900 ;
        RECT 7.900 137.300 9.700 137.600 ;
        RECT 11.000 137.500 11.400 137.900 ;
        RECT 7.900 137.200 8.300 137.300 ;
        RECT 9.300 137.200 9.700 137.300 ;
        RECT 6.200 136.500 6.600 136.600 ;
        RECT 8.500 136.500 8.900 136.600 ;
        RECT 6.200 136.200 8.900 136.500 ;
        RECT 9.200 136.500 10.300 136.800 ;
        RECT 9.200 135.900 9.500 136.500 ;
        RECT 9.900 136.400 10.300 136.500 ;
        RECT 11.100 136.600 11.800 137.000 ;
        RECT 11.100 136.100 11.400 136.600 ;
        RECT 7.100 135.700 9.500 135.900 ;
        RECT 4.600 135.600 9.500 135.700 ;
        RECT 10.200 135.800 11.400 136.100 ;
        RECT 4.600 135.500 7.500 135.600 ;
        RECT 4.600 135.400 7.400 135.500 ;
        RECT 3.000 133.800 3.400 135.200 ;
        RECT 7.800 135.100 8.200 135.200 ;
        RECT 5.700 134.800 8.200 135.100 ;
        RECT 5.700 134.700 6.100 134.800 ;
        RECT 6.500 134.200 6.900 134.300 ;
        RECT 10.200 134.200 10.500 135.800 ;
        RECT 13.400 135.600 13.800 139.900 ;
        RECT 15.500 136.200 15.900 139.900 ;
        RECT 16.200 136.800 16.600 137.200 ;
        RECT 16.300 136.200 16.600 136.800 ;
        RECT 15.500 135.900 16.000 136.200 ;
        RECT 16.300 135.900 17.000 136.200 ;
        RECT 11.700 135.300 13.800 135.600 ;
        RECT 11.700 135.200 12.100 135.300 ;
        RECT 12.500 134.900 12.900 135.000 ;
        RECT 11.000 134.600 12.900 134.900 ;
        RECT 11.000 134.500 11.400 134.600 ;
        RECT 5.000 133.900 10.500 134.200 ;
        RECT 5.000 133.800 5.800 133.900 ;
        RECT 1.400 133.400 3.400 133.800 ;
        RECT 1.400 131.100 1.800 133.400 ;
        RECT 3.000 131.100 3.400 133.400 ;
        RECT 4.600 131.100 5.000 133.500 ;
        RECT 7.100 132.800 7.400 133.900 ;
        RECT 9.900 133.800 10.300 133.900 ;
        RECT 13.400 133.600 13.800 135.300 ;
        RECT 15.700 135.200 16.000 135.900 ;
        RECT 16.600 135.800 17.000 135.900 ;
        RECT 17.400 135.800 17.800 136.600 ;
        RECT 15.000 134.400 15.400 135.200 ;
        RECT 15.700 134.800 16.200 135.200 ;
        RECT 16.600 135.100 16.900 135.800 ;
        RECT 18.200 135.100 18.600 139.900 ;
        RECT 19.800 135.800 20.200 136.600 ;
        RECT 16.600 134.800 18.600 135.100 ;
        RECT 15.700 134.200 16.000 134.800 ;
        RECT 14.200 134.100 14.600 134.200 ;
        RECT 14.200 133.800 15.000 134.100 ;
        RECT 15.700 133.800 17.000 134.200 ;
        RECT 14.600 133.600 15.000 133.800 ;
        RECT 11.900 133.300 13.800 133.600 ;
        RECT 11.900 133.200 12.300 133.300 ;
        RECT 6.200 132.100 6.600 132.500 ;
        RECT 7.000 132.400 7.400 132.800 ;
        RECT 7.900 132.700 8.300 132.800 ;
        RECT 7.900 132.400 9.300 132.700 ;
        RECT 9.000 132.100 9.300 132.400 ;
        RECT 11.000 132.100 11.400 132.500 ;
        RECT 6.200 131.800 7.200 132.100 ;
        RECT 6.800 131.100 7.200 131.800 ;
        RECT 9.000 131.100 9.400 132.100 ;
        RECT 11.000 131.800 11.700 132.100 ;
        RECT 11.100 131.100 11.700 131.800 ;
        RECT 13.400 131.100 13.800 133.300 ;
        RECT 14.300 133.100 16.100 133.300 ;
        RECT 16.600 133.100 16.900 133.800 ;
        RECT 18.200 133.100 18.600 134.800 ;
        RECT 19.000 133.400 19.400 134.200 ;
        RECT 20.600 133.100 21.000 139.900 ;
        RECT 22.200 137.500 22.600 139.500 ;
        RECT 22.200 135.800 22.500 137.500 ;
        RECT 24.300 137.200 24.700 139.900 ;
        RECT 24.300 136.800 25.000 137.200 ;
        RECT 24.300 136.400 24.700 136.800 ;
        RECT 24.300 136.100 25.100 136.400 ;
        RECT 22.200 135.500 24.100 135.800 ;
        RECT 21.400 135.100 21.800 135.200 ;
        RECT 22.200 135.100 22.600 135.200 ;
        RECT 21.400 134.800 22.600 135.100 ;
        RECT 22.200 134.400 22.600 134.800 ;
        RECT 23.000 134.400 23.400 135.200 ;
        RECT 23.800 134.500 24.100 135.500 ;
        RECT 21.400 133.400 21.800 134.200 ;
        RECT 23.800 134.100 24.500 134.500 ;
        RECT 24.800 134.200 25.100 136.100 ;
        RECT 27.000 136.200 27.400 139.900 ;
        RECT 28.600 136.400 29.000 139.900 ;
        RECT 27.000 135.900 28.300 136.200 ;
        RECT 28.600 135.900 29.100 136.400 ;
        RECT 25.400 134.800 25.800 135.600 ;
        RECT 27.000 134.800 27.500 135.200 ;
        RECT 27.100 134.400 27.500 134.800 ;
        RECT 28.000 134.900 28.300 135.900 ;
        RECT 28.000 134.500 28.500 134.900 ;
        RECT 23.800 133.900 24.300 134.100 ;
        RECT 22.200 133.600 24.300 133.900 ;
        RECT 24.800 133.800 25.800 134.200 ;
        RECT 14.200 133.000 16.200 133.100 ;
        RECT 14.200 131.100 14.600 133.000 ;
        RECT 15.800 131.100 16.200 133.000 ;
        RECT 16.600 131.100 17.000 133.100 ;
        RECT 17.700 132.800 18.600 133.100 ;
        RECT 20.100 132.800 21.000 133.100 ;
        RECT 17.700 131.100 18.100 132.800 ;
        RECT 20.100 132.200 20.500 132.800 ;
        RECT 19.800 131.800 20.500 132.200 ;
        RECT 20.100 131.100 20.500 131.800 ;
        RECT 22.200 132.500 22.500 133.600 ;
        RECT 24.800 133.500 25.100 133.800 ;
        RECT 28.000 133.700 28.300 134.500 ;
        RECT 28.800 134.200 29.100 135.900 ;
        RECT 31.000 135.600 31.400 139.900 ;
        RECT 32.600 135.600 33.000 139.900 ;
        RECT 34.200 135.600 34.600 139.900 ;
        RECT 35.800 135.600 36.200 139.900 ;
        RECT 39.300 139.200 39.700 139.900 ;
        RECT 39.300 138.800 40.200 139.200 ;
        RECT 39.300 136.400 39.700 138.800 ;
        RECT 41.400 137.500 41.800 139.500 ;
        RECT 38.900 136.100 39.700 136.400 ;
        RECT 31.000 135.200 31.900 135.600 ;
        RECT 32.600 135.200 33.700 135.600 ;
        RECT 34.200 135.200 35.300 135.600 ;
        RECT 35.800 135.200 37.000 135.600 ;
        RECT 31.500 134.500 31.900 135.200 ;
        RECT 33.300 134.500 33.700 135.200 ;
        RECT 34.900 134.500 35.300 135.200 ;
        RECT 28.600 134.100 29.100 134.200 ;
        RECT 29.400 134.100 29.800 134.200 ;
        RECT 28.600 133.800 29.800 134.100 ;
        RECT 31.500 134.100 32.800 134.500 ;
        RECT 33.300 134.100 34.500 134.500 ;
        RECT 34.900 134.100 36.200 134.500 ;
        RECT 31.500 133.800 31.900 134.100 ;
        RECT 33.300 133.800 33.700 134.100 ;
        RECT 34.900 133.800 35.300 134.100 ;
        RECT 36.600 133.800 37.000 135.200 ;
        RECT 37.400 135.100 37.800 135.200 ;
        RECT 38.200 135.100 38.600 135.600 ;
        RECT 37.400 134.800 38.600 135.100 ;
        RECT 38.900 134.200 39.200 136.100 ;
        RECT 41.500 135.800 41.800 137.500 ;
        RECT 42.200 136.200 42.600 139.900 ;
        RECT 43.800 139.600 45.800 139.900 ;
        RECT 43.800 136.200 44.200 139.600 ;
        RECT 42.200 135.900 44.200 136.200 ;
        RECT 44.600 135.900 45.000 139.300 ;
        RECT 45.400 135.900 45.800 139.600 ;
        RECT 47.800 137.500 48.200 139.500 ;
        RECT 39.900 135.500 41.800 135.800 ;
        RECT 44.600 135.600 44.900 135.900 ;
        RECT 47.800 135.800 48.100 137.500 ;
        RECT 49.900 136.400 50.300 139.900 ;
        RECT 49.900 136.100 50.700 136.400 ;
        RECT 39.900 134.500 40.200 135.500 ;
        RECT 42.600 135.200 43.000 135.400 ;
        RECT 43.900 135.300 44.900 135.600 ;
        RECT 43.900 135.200 44.200 135.300 ;
        RECT 38.200 133.800 39.200 134.200 ;
        RECT 39.500 134.100 40.200 134.500 ;
        RECT 40.600 134.400 41.000 135.200 ;
        RECT 41.400 134.400 41.800 135.200 ;
        RECT 42.200 134.900 43.000 135.200 ;
        RECT 42.200 134.800 42.600 134.900 ;
        RECT 43.800 134.800 44.200 135.200 ;
        RECT 45.400 134.800 45.800 135.600 ;
        RECT 47.800 135.500 49.700 135.800 ;
        RECT 24.700 133.300 25.100 133.500 ;
        RECT 24.300 133.000 25.100 133.300 ;
        RECT 27.000 133.400 28.300 133.700 ;
        RECT 22.200 131.500 22.600 132.500 ;
        RECT 24.300 131.500 24.700 133.000 ;
        RECT 27.000 131.100 27.400 133.400 ;
        RECT 28.800 133.100 29.100 133.800 ;
        RECT 28.600 132.800 29.100 133.100 ;
        RECT 31.000 133.400 31.900 133.800 ;
        RECT 32.600 133.400 33.700 133.800 ;
        RECT 34.200 133.400 35.300 133.800 ;
        RECT 35.800 133.400 37.000 133.800 ;
        RECT 38.900 133.500 39.200 133.800 ;
        RECT 39.700 133.900 40.200 134.100 ;
        RECT 39.700 133.600 41.800 133.900 ;
        RECT 43.000 133.800 43.400 134.600 ;
        RECT 28.600 131.100 29.000 132.800 ;
        RECT 31.000 131.100 31.400 133.400 ;
        RECT 32.600 131.100 33.000 133.400 ;
        RECT 34.200 131.100 34.600 133.400 ;
        RECT 35.800 131.100 36.200 133.400 ;
        RECT 38.900 133.300 39.300 133.500 ;
        RECT 38.900 133.000 39.700 133.300 ;
        RECT 39.300 131.500 39.700 133.000 ;
        RECT 41.500 132.500 41.800 133.600 ;
        RECT 43.900 133.100 44.200 134.800 ;
        RECT 44.500 134.400 44.900 134.800 ;
        RECT 47.800 134.400 48.200 135.200 ;
        RECT 48.600 134.400 49.000 135.200 ;
        RECT 49.400 134.500 49.700 135.500 ;
        RECT 44.600 134.200 44.900 134.400 ;
        RECT 44.600 133.800 45.000 134.200 ;
        RECT 49.400 134.100 50.100 134.500 ;
        RECT 50.400 134.200 50.700 136.100 ;
        RECT 52.600 135.600 53.000 139.900 ;
        RECT 54.700 137.900 55.300 139.900 ;
        RECT 57.000 137.900 57.400 139.900 ;
        RECT 59.200 138.200 59.600 139.900 ;
        RECT 59.200 137.900 60.200 138.200 ;
        RECT 55.000 137.500 55.400 137.900 ;
        RECT 57.100 137.600 57.400 137.900 ;
        RECT 56.700 137.300 58.500 137.600 ;
        RECT 59.800 137.500 60.200 137.900 ;
        RECT 56.700 137.200 57.100 137.300 ;
        RECT 58.100 137.200 58.500 137.300 ;
        RECT 54.600 136.600 55.300 137.000 ;
        RECT 55.000 136.100 55.300 136.600 ;
        RECT 56.100 136.500 57.200 136.800 ;
        RECT 56.100 136.400 56.500 136.500 ;
        RECT 55.000 135.800 56.200 136.100 ;
        RECT 51.000 134.800 51.400 135.600 ;
        RECT 52.600 135.300 54.700 135.600 ;
        RECT 50.400 134.100 51.400 134.200 ;
        RECT 51.800 134.100 52.200 134.200 ;
        RECT 49.400 133.900 49.900 134.100 ;
        RECT 47.800 133.600 49.900 133.900 ;
        RECT 50.400 133.800 52.200 134.100 ;
        RECT 41.400 131.500 41.800 132.500 ;
        RECT 43.700 131.100 44.500 133.100 ;
        RECT 47.800 132.500 48.100 133.600 ;
        RECT 50.400 133.500 50.700 133.800 ;
        RECT 50.300 133.300 50.700 133.500 ;
        RECT 49.900 133.000 50.700 133.300 ;
        RECT 52.600 133.600 53.000 135.300 ;
        RECT 54.300 135.200 54.700 135.300 ;
        RECT 53.500 134.900 53.900 135.000 ;
        RECT 53.500 134.600 55.400 134.900 ;
        RECT 55.000 134.500 55.400 134.600 ;
        RECT 55.900 134.200 56.200 135.800 ;
        RECT 56.900 135.900 57.200 136.500 ;
        RECT 57.500 136.500 57.900 136.600 ;
        RECT 59.800 136.500 60.200 136.600 ;
        RECT 57.500 136.200 60.200 136.500 ;
        RECT 56.900 135.700 59.300 135.900 ;
        RECT 61.400 135.700 61.800 139.900 ;
        RECT 62.200 136.200 62.600 139.900 ;
        RECT 63.800 139.600 65.800 139.900 ;
        RECT 63.800 136.200 64.200 139.600 ;
        RECT 62.200 135.900 64.200 136.200 ;
        RECT 64.600 135.900 65.000 139.300 ;
        RECT 65.400 135.900 65.800 139.600 ;
        RECT 56.900 135.600 61.800 135.700 ;
        RECT 64.600 135.600 64.900 135.900 ;
        RECT 58.900 135.500 61.800 135.600 ;
        RECT 59.000 135.400 61.800 135.500 ;
        RECT 62.600 135.200 63.000 135.400 ;
        RECT 63.900 135.300 64.900 135.600 ;
        RECT 63.900 135.200 64.200 135.300 ;
        RECT 58.200 135.100 58.600 135.200 ;
        RECT 58.200 134.800 60.700 135.100 ;
        RECT 62.200 134.900 63.000 135.200 ;
        RECT 62.200 134.800 62.600 134.900 ;
        RECT 63.800 134.800 64.200 135.200 ;
        RECT 65.400 135.100 65.800 135.600 ;
        RECT 66.200 135.100 66.600 135.200 ;
        RECT 65.400 134.800 66.600 135.100 ;
        RECT 60.300 134.700 60.700 134.800 ;
        RECT 59.500 134.200 59.900 134.300 ;
        RECT 55.900 133.900 61.400 134.200 ;
        RECT 56.100 133.800 56.500 133.900 ;
        RECT 52.600 133.300 54.500 133.600 ;
        RECT 47.800 131.500 48.200 132.500 ;
        RECT 49.900 131.500 50.300 133.000 ;
        RECT 52.600 131.100 53.000 133.300 ;
        RECT 54.100 133.200 54.500 133.300 ;
        RECT 59.000 132.800 59.300 133.900 ;
        RECT 60.600 133.800 61.400 133.900 ;
        RECT 63.000 133.800 63.400 134.600 ;
        RECT 58.100 132.700 58.500 132.800 ;
        RECT 55.000 132.100 55.400 132.500 ;
        RECT 57.100 132.400 58.500 132.700 ;
        RECT 59.000 132.400 59.400 132.800 ;
        RECT 57.100 132.100 57.400 132.400 ;
        RECT 59.800 132.100 60.200 132.500 ;
        RECT 54.700 131.800 55.400 132.100 ;
        RECT 54.700 131.100 55.300 131.800 ;
        RECT 57.000 131.100 57.400 132.100 ;
        RECT 59.200 131.800 60.200 132.100 ;
        RECT 59.200 131.100 59.600 131.800 ;
        RECT 61.400 131.100 61.800 133.500 ;
        RECT 63.900 133.200 64.200 134.800 ;
        RECT 64.500 134.400 64.900 134.800 ;
        RECT 64.600 134.200 64.900 134.400 ;
        RECT 64.600 133.800 65.000 134.200 ;
        RECT 65.400 134.100 65.800 134.200 ;
        RECT 66.200 134.100 66.600 134.200 ;
        RECT 65.400 133.800 66.600 134.100 ;
        RECT 66.200 133.400 66.600 133.800 ;
        RECT 67.000 134.100 67.400 139.900 ;
        RECT 69.900 139.200 70.300 139.900 ;
        RECT 69.400 138.800 70.300 139.200 ;
        RECT 67.800 135.800 68.200 136.600 ;
        RECT 69.900 136.200 70.300 138.800 ;
        RECT 70.600 136.800 71.000 137.200 ;
        RECT 70.700 136.200 71.000 136.800 ;
        RECT 71.800 136.200 72.200 139.900 ;
        RECT 73.400 136.400 73.800 139.900 ;
        RECT 75.000 137.500 75.400 139.500 ;
        RECT 69.900 135.900 70.400 136.200 ;
        RECT 70.700 135.900 71.400 136.200 ;
        RECT 71.800 135.900 73.100 136.200 ;
        RECT 69.400 134.400 69.800 135.200 ;
        RECT 70.100 134.200 70.400 135.900 ;
        RECT 71.000 135.800 71.400 135.900 ;
        RECT 71.000 135.100 71.400 135.200 ;
        RECT 71.800 135.100 72.300 135.200 ;
        RECT 71.000 134.800 72.300 135.100 ;
        RECT 71.900 134.400 72.300 134.800 ;
        RECT 72.800 134.900 73.100 135.900 ;
        RECT 73.400 135.800 73.900 136.400 ;
        RECT 72.800 134.500 73.300 134.900 ;
        RECT 68.600 134.100 69.000 134.200 ;
        RECT 67.000 133.800 69.400 134.100 ;
        RECT 70.100 133.800 71.400 134.200 ;
        RECT 63.900 133.100 65.000 133.200 ;
        RECT 63.700 132.800 65.000 133.100 ;
        RECT 67.000 133.100 67.400 133.800 ;
        RECT 69.000 133.600 69.400 133.800 ;
        RECT 68.700 133.100 70.500 133.300 ;
        RECT 71.000 133.100 71.300 133.800 ;
        RECT 72.800 133.700 73.100 134.500 ;
        RECT 73.600 134.200 73.900 135.800 ;
        RECT 75.000 135.800 75.300 137.500 ;
        RECT 77.100 136.400 77.500 139.900 ;
        RECT 77.100 136.100 77.900 136.400 ;
        RECT 75.000 135.500 76.900 135.800 ;
        RECT 75.000 134.400 75.400 135.200 ;
        RECT 75.800 134.400 76.200 135.200 ;
        RECT 76.600 134.500 76.900 135.500 ;
        RECT 73.400 133.800 73.900 134.200 ;
        RECT 76.600 134.100 77.300 134.500 ;
        RECT 77.600 134.200 77.900 136.100 ;
        RECT 78.200 134.800 78.600 135.600 ;
        RECT 79.000 134.800 79.400 135.200 ;
        RECT 80.600 135.100 81.000 139.900 ;
        RECT 83.300 139.200 83.700 139.900 ;
        RECT 83.300 138.800 84.200 139.200 ;
        RECT 82.600 136.800 83.000 137.200 ;
        RECT 81.400 135.800 81.800 136.600 ;
        RECT 82.600 136.200 82.900 136.800 ;
        RECT 83.300 136.200 83.700 138.800 ;
        RECT 82.200 135.900 82.900 136.200 ;
        RECT 83.200 135.900 83.700 136.200 ;
        RECT 86.700 136.200 87.100 139.900 ;
        RECT 87.400 136.800 87.800 137.200 ;
        RECT 87.500 136.200 87.800 136.800 ;
        RECT 86.700 135.900 87.200 136.200 ;
        RECT 87.500 135.900 88.200 136.200 ;
        RECT 82.200 135.800 82.600 135.900 ;
        RECT 82.200 135.100 82.500 135.800 ;
        RECT 80.600 134.800 82.500 135.100 ;
        RECT 76.600 133.900 77.100 134.100 ;
        RECT 71.800 133.400 73.100 133.700 ;
        RECT 67.000 132.800 67.900 133.100 ;
        RECT 63.700 131.100 64.500 132.800 ;
        RECT 67.500 131.100 67.900 132.800 ;
        RECT 68.600 133.000 70.600 133.100 ;
        RECT 68.600 131.100 69.000 133.000 ;
        RECT 70.200 131.100 70.600 133.000 ;
        RECT 71.000 131.100 71.400 133.100 ;
        RECT 71.800 131.100 72.200 133.400 ;
        RECT 73.600 133.100 73.900 133.800 ;
        RECT 73.400 132.800 73.900 133.100 ;
        RECT 75.000 133.600 77.100 133.900 ;
        RECT 77.600 133.800 78.600 134.200 ;
        RECT 79.000 134.100 79.300 134.800 ;
        RECT 79.800 134.100 80.200 134.200 ;
        RECT 79.000 133.800 80.200 134.100 ;
        RECT 73.400 131.100 73.800 132.800 ;
        RECT 75.000 132.500 75.300 133.600 ;
        RECT 77.600 133.500 77.900 133.800 ;
        RECT 77.500 133.300 77.900 133.500 ;
        RECT 79.800 133.400 80.200 133.800 ;
        RECT 77.100 133.000 77.900 133.300 ;
        RECT 80.600 133.100 81.000 134.800 ;
        RECT 83.200 134.200 83.500 135.900 ;
        RECT 83.800 134.400 84.200 135.200 ;
        RECT 86.200 134.400 86.600 135.200 ;
        RECT 86.900 134.200 87.200 135.900 ;
        RECT 87.800 135.800 88.200 135.900 ;
        RECT 88.600 135.800 89.000 136.600 ;
        RECT 87.800 135.100 88.100 135.800 ;
        RECT 89.400 135.100 89.800 139.900 ;
        RECT 91.000 135.700 91.400 139.900 ;
        RECT 93.200 138.200 93.600 139.900 ;
        RECT 92.600 137.900 93.600 138.200 ;
        RECT 95.400 137.900 95.800 139.900 ;
        RECT 97.500 137.900 98.100 139.900 ;
        RECT 92.600 137.500 93.000 137.900 ;
        RECT 95.400 137.600 95.700 137.900 ;
        RECT 94.300 137.300 96.100 137.600 ;
        RECT 97.400 137.500 97.800 137.900 ;
        RECT 94.300 137.200 94.700 137.300 ;
        RECT 95.700 137.200 96.100 137.300 ;
        RECT 92.600 136.500 93.000 136.600 ;
        RECT 94.900 136.500 95.300 136.600 ;
        RECT 92.600 136.200 95.300 136.500 ;
        RECT 95.600 136.500 96.700 136.800 ;
        RECT 95.600 135.900 95.900 136.500 ;
        RECT 96.300 136.400 96.700 136.500 ;
        RECT 97.500 136.600 98.200 137.000 ;
        RECT 97.500 136.100 97.800 136.600 ;
        RECT 93.500 135.700 95.900 135.900 ;
        RECT 91.000 135.600 95.900 135.700 ;
        RECT 96.600 135.800 97.800 136.100 ;
        RECT 91.000 135.500 93.900 135.600 ;
        RECT 91.000 135.400 93.800 135.500 ;
        RECT 94.200 135.100 94.600 135.200 ;
        RECT 87.800 134.800 89.800 135.100 ;
        RECT 82.200 133.800 83.500 134.200 ;
        RECT 84.600 134.100 85.000 134.200 ;
        RECT 84.200 133.800 85.000 134.100 ;
        RECT 85.400 134.100 85.800 134.200 ;
        RECT 86.900 134.100 88.200 134.200 ;
        RECT 88.600 134.100 89.000 134.200 ;
        RECT 85.400 133.800 86.200 134.100 ;
        RECT 86.900 133.800 89.000 134.100 ;
        RECT 82.300 133.100 82.600 133.800 ;
        RECT 84.200 133.600 84.600 133.800 ;
        RECT 85.800 133.600 86.200 133.800 ;
        RECT 83.100 133.100 84.900 133.300 ;
        RECT 85.500 133.100 87.300 133.300 ;
        RECT 87.800 133.100 88.100 133.800 ;
        RECT 89.400 133.100 89.800 134.800 ;
        RECT 92.100 134.800 94.600 135.100 ;
        RECT 95.800 135.100 96.200 135.200 ;
        RECT 96.600 135.100 96.900 135.800 ;
        RECT 99.800 135.600 100.200 139.900 ;
        RECT 98.100 135.300 100.200 135.600 ;
        RECT 102.200 135.700 102.600 139.900 ;
        RECT 104.400 138.200 104.800 139.900 ;
        RECT 103.800 137.900 104.800 138.200 ;
        RECT 106.600 137.900 107.000 139.900 ;
        RECT 108.700 137.900 109.300 139.900 ;
        RECT 103.800 137.500 104.200 137.900 ;
        RECT 106.600 137.600 106.900 137.900 ;
        RECT 105.500 137.300 107.300 137.600 ;
        RECT 108.600 137.500 109.000 137.900 ;
        RECT 105.500 137.200 105.900 137.300 ;
        RECT 106.900 137.200 107.300 137.300 ;
        RECT 111.000 137.100 111.400 139.900 ;
        RECT 111.800 137.100 112.200 137.200 ;
        RECT 103.800 136.500 104.200 136.600 ;
        RECT 106.100 136.500 106.500 136.600 ;
        RECT 103.800 136.200 106.500 136.500 ;
        RECT 106.800 136.500 107.900 136.800 ;
        RECT 106.800 135.900 107.100 136.500 ;
        RECT 107.500 136.400 107.900 136.500 ;
        RECT 108.700 136.600 109.400 137.000 ;
        RECT 111.000 136.800 112.200 137.100 ;
        RECT 108.700 136.100 109.000 136.600 ;
        RECT 104.700 135.700 107.100 135.900 ;
        RECT 102.200 135.600 107.100 135.700 ;
        RECT 107.800 135.800 109.000 136.100 ;
        RECT 102.200 135.500 105.100 135.600 ;
        RECT 102.200 135.400 105.000 135.500 ;
        RECT 98.100 135.200 98.500 135.300 ;
        RECT 95.800 134.800 96.900 135.100 ;
        RECT 98.900 134.900 99.300 135.000 ;
        RECT 92.100 134.700 92.500 134.800 ;
        RECT 93.400 134.700 93.800 134.800 ;
        RECT 92.900 134.200 93.300 134.300 ;
        RECT 96.600 134.200 96.900 134.800 ;
        RECT 97.400 134.600 99.300 134.900 ;
        RECT 97.400 134.500 97.800 134.600 ;
        RECT 90.200 133.400 90.600 134.200 ;
        RECT 91.400 133.900 96.900 134.200 ;
        RECT 91.400 133.800 92.200 133.900 ;
        RECT 75.000 131.500 75.400 132.500 ;
        RECT 77.100 132.200 77.500 133.000 ;
        RECT 80.600 132.800 81.500 133.100 ;
        RECT 76.600 131.800 77.500 132.200 ;
        RECT 77.100 131.500 77.500 131.800 ;
        RECT 81.100 131.100 81.500 132.800 ;
        RECT 82.200 131.100 82.600 133.100 ;
        RECT 83.000 133.000 85.000 133.100 ;
        RECT 83.000 131.100 83.400 133.000 ;
        RECT 84.600 131.100 85.000 133.000 ;
        RECT 85.400 133.000 87.400 133.100 ;
        RECT 85.400 131.100 85.800 133.000 ;
        RECT 87.000 131.100 87.400 133.000 ;
        RECT 87.800 131.100 88.200 133.100 ;
        RECT 88.900 132.800 89.800 133.100 ;
        RECT 88.900 131.100 89.300 132.800 ;
        RECT 91.000 131.100 91.400 133.500 ;
        RECT 93.500 132.800 93.800 133.900 ;
        RECT 96.300 133.800 96.700 133.900 ;
        RECT 99.800 133.600 100.200 135.300 ;
        RECT 105.400 135.100 105.800 135.200 ;
        RECT 103.300 134.800 105.800 135.100 ;
        RECT 103.300 134.700 103.700 134.800 ;
        RECT 104.100 134.200 104.500 134.300 ;
        RECT 107.800 134.200 108.100 135.800 ;
        RECT 111.000 135.600 111.400 136.800 ;
        RECT 109.300 135.300 111.400 135.600 ;
        RECT 109.300 135.200 109.700 135.300 ;
        RECT 110.100 134.900 110.500 135.000 ;
        RECT 108.600 134.600 110.500 134.900 ;
        RECT 108.600 134.500 109.000 134.600 ;
        RECT 102.600 133.900 108.100 134.200 ;
        RECT 102.600 133.800 103.400 133.900 ;
        RECT 104.600 133.800 105.000 133.900 ;
        RECT 107.500 133.800 107.900 133.900 ;
        RECT 98.300 133.300 100.200 133.600 ;
        RECT 98.300 133.200 98.700 133.300 ;
        RECT 92.600 132.100 93.000 132.500 ;
        RECT 93.400 132.400 93.800 132.800 ;
        RECT 94.300 132.700 94.700 132.800 ;
        RECT 94.300 132.400 95.700 132.700 ;
        RECT 95.400 132.100 95.700 132.400 ;
        RECT 97.400 132.100 97.800 132.500 ;
        RECT 92.600 131.800 93.600 132.100 ;
        RECT 93.200 131.100 93.600 131.800 ;
        RECT 95.400 131.100 95.800 132.100 ;
        RECT 97.400 131.800 98.100 132.100 ;
        RECT 97.500 131.100 98.100 131.800 ;
        RECT 99.800 131.100 100.200 133.300 ;
        RECT 102.200 131.100 102.600 133.500 ;
        RECT 104.700 132.800 105.000 133.800 ;
        RECT 111.000 133.600 111.400 135.300 ;
        RECT 112.600 135.100 113.000 139.900 ;
        RECT 114.600 136.800 115.000 137.200 ;
        RECT 113.400 135.800 113.800 136.600 ;
        RECT 114.600 136.200 114.900 136.800 ;
        RECT 115.300 136.200 115.700 139.900 ;
        RECT 119.300 136.400 119.700 139.900 ;
        RECT 121.400 137.500 121.800 139.500 ;
        RECT 114.200 135.900 114.900 136.200 ;
        RECT 115.200 135.900 115.700 136.200 ;
        RECT 118.900 136.100 119.700 136.400 ;
        RECT 114.200 135.800 114.600 135.900 ;
        RECT 114.200 135.100 114.500 135.800 ;
        RECT 112.600 134.800 114.500 135.100 ;
        RECT 109.500 133.300 111.400 133.600 ;
        RECT 111.800 133.400 112.200 134.200 ;
        RECT 109.500 133.200 109.900 133.300 ;
        RECT 103.800 132.100 104.200 132.500 ;
        RECT 104.600 132.400 105.000 132.800 ;
        RECT 105.500 132.700 105.900 132.800 ;
        RECT 105.500 132.400 106.900 132.700 ;
        RECT 106.600 132.100 106.900 132.400 ;
        RECT 108.600 132.100 109.000 132.500 ;
        RECT 103.800 131.800 104.800 132.100 ;
        RECT 104.400 131.100 104.800 131.800 ;
        RECT 106.600 131.100 107.000 132.100 ;
        RECT 108.600 131.800 109.300 132.100 ;
        RECT 108.700 131.100 109.300 131.800 ;
        RECT 111.000 131.100 111.400 133.300 ;
        RECT 112.600 133.100 113.000 134.800 ;
        RECT 115.200 134.200 115.500 135.900 ;
        RECT 115.800 134.400 116.200 135.200 ;
        RECT 118.200 134.800 118.600 135.600 ;
        RECT 118.900 134.200 119.200 136.100 ;
        RECT 121.500 135.800 121.800 137.500 ;
        RECT 119.900 135.500 121.800 135.800 ;
        RECT 119.900 134.500 120.200 135.500 ;
        RECT 113.400 134.100 113.800 134.200 ;
        RECT 114.200 134.100 115.500 134.200 ;
        RECT 116.600 134.100 117.000 134.200 ;
        RECT 113.400 133.800 115.500 134.100 ;
        RECT 116.200 133.800 117.000 134.100 ;
        RECT 118.200 133.800 119.200 134.200 ;
        RECT 119.500 134.100 120.200 134.500 ;
        RECT 120.600 134.400 121.000 135.200 ;
        RECT 121.400 134.400 121.800 135.200 ;
        RECT 123.000 135.100 123.400 139.900 ;
        RECT 125.000 136.800 125.400 137.200 ;
        RECT 123.800 135.800 124.200 136.600 ;
        RECT 125.000 136.200 125.300 136.800 ;
        RECT 125.700 136.200 126.100 139.900 ;
        RECT 124.600 135.900 125.300 136.200 ;
        RECT 125.600 135.900 126.100 136.200 ;
        RECT 124.600 135.800 125.000 135.900 ;
        RECT 124.600 135.100 124.900 135.800 ;
        RECT 123.000 134.800 124.900 135.100 ;
        RECT 114.300 133.100 114.600 133.800 ;
        RECT 116.200 133.600 116.600 133.800 ;
        RECT 118.900 133.500 119.200 133.800 ;
        RECT 119.700 133.900 120.200 134.100 ;
        RECT 119.700 133.600 121.800 133.900 ;
        RECT 118.900 133.300 119.300 133.500 ;
        RECT 115.100 133.100 116.900 133.300 ;
        RECT 112.600 132.800 113.500 133.100 ;
        RECT 113.100 131.100 113.500 132.800 ;
        RECT 114.200 131.100 114.600 133.100 ;
        RECT 115.000 133.000 117.000 133.100 ;
        RECT 118.900 133.000 119.700 133.300 ;
        RECT 115.000 131.100 115.400 133.000 ;
        RECT 116.600 131.100 117.000 133.000 ;
        RECT 119.300 132.200 119.700 133.000 ;
        RECT 121.500 132.500 121.800 133.600 ;
        RECT 122.200 133.400 122.600 134.200 ;
        RECT 123.000 133.100 123.400 134.800 ;
        RECT 125.600 134.200 125.900 135.900 ;
        RECT 127.800 135.600 128.200 139.900 ;
        RECT 129.900 137.900 130.500 139.900 ;
        RECT 132.200 137.900 132.600 139.900 ;
        RECT 134.400 138.200 134.800 139.900 ;
        RECT 134.400 137.900 135.400 138.200 ;
        RECT 130.200 137.500 130.600 137.900 ;
        RECT 132.300 137.600 132.600 137.900 ;
        RECT 131.900 137.300 133.700 137.600 ;
        RECT 135.000 137.500 135.400 137.900 ;
        RECT 131.900 137.200 132.300 137.300 ;
        RECT 133.300 137.200 133.700 137.300 ;
        RECT 129.800 136.600 130.500 137.000 ;
        RECT 130.200 136.100 130.500 136.600 ;
        RECT 131.300 136.500 132.400 136.800 ;
        RECT 131.300 136.400 131.700 136.500 ;
        RECT 130.200 135.800 131.400 136.100 ;
        RECT 127.800 135.300 129.900 135.600 ;
        RECT 126.200 134.400 126.600 135.200 ;
        RECT 124.600 133.800 125.900 134.200 ;
        RECT 127.000 134.100 127.400 134.200 ;
        RECT 126.600 133.800 127.400 134.100 ;
        RECT 124.700 133.100 125.000 133.800 ;
        RECT 126.600 133.600 127.000 133.800 ;
        RECT 127.800 133.600 128.200 135.300 ;
        RECT 129.500 135.200 129.900 135.300 ;
        RECT 128.700 134.900 129.100 135.000 ;
        RECT 128.700 134.600 130.600 134.900 ;
        RECT 130.200 134.500 130.600 134.600 ;
        RECT 131.100 134.200 131.400 135.800 ;
        RECT 132.100 135.900 132.400 136.500 ;
        RECT 132.700 136.500 133.100 136.600 ;
        RECT 135.000 136.500 135.400 136.600 ;
        RECT 132.700 136.200 135.400 136.500 ;
        RECT 132.100 135.700 134.500 135.900 ;
        RECT 136.600 135.700 137.000 139.900 ;
        RECT 132.100 135.600 137.000 135.700 ;
        RECT 134.100 135.500 137.000 135.600 ;
        RECT 134.200 135.400 137.000 135.500 ;
        RECT 137.400 135.700 137.800 139.900 ;
        RECT 139.600 138.200 140.000 139.900 ;
        RECT 139.000 137.900 140.000 138.200 ;
        RECT 141.800 137.900 142.200 139.900 ;
        RECT 143.900 137.900 144.500 139.900 ;
        RECT 139.000 137.500 139.400 137.900 ;
        RECT 141.800 137.600 142.100 137.900 ;
        RECT 140.700 137.300 142.500 137.600 ;
        RECT 143.800 137.500 144.200 137.900 ;
        RECT 140.700 137.200 141.100 137.300 ;
        RECT 142.100 137.200 142.500 137.300 ;
        RECT 146.200 137.100 146.600 139.900 ;
        RECT 147.000 137.100 147.400 137.200 ;
        RECT 139.000 136.500 139.400 136.600 ;
        RECT 141.300 136.500 141.700 136.600 ;
        RECT 139.000 136.200 141.700 136.500 ;
        RECT 142.000 136.500 143.100 136.800 ;
        RECT 142.000 135.900 142.300 136.500 ;
        RECT 142.700 136.400 143.100 136.500 ;
        RECT 143.900 136.600 144.600 137.000 ;
        RECT 146.200 136.800 147.400 137.100 ;
        RECT 143.900 136.100 144.200 136.600 ;
        RECT 139.900 135.700 142.300 135.900 ;
        RECT 137.400 135.600 142.300 135.700 ;
        RECT 143.000 135.800 144.200 136.100 ;
        RECT 137.400 135.500 140.300 135.600 ;
        RECT 137.400 135.400 140.200 135.500 ;
        RECT 133.400 135.100 133.800 135.200 ;
        RECT 140.600 135.100 141.000 135.200 ;
        RECT 142.200 135.100 142.600 135.200 ;
        RECT 133.400 134.800 135.900 135.100 ;
        RECT 135.500 134.700 135.900 134.800 ;
        RECT 138.500 134.800 142.600 135.100 ;
        RECT 138.500 134.700 138.900 134.800 ;
        RECT 134.700 134.200 135.100 134.300 ;
        RECT 139.300 134.200 139.700 134.300 ;
        RECT 143.000 134.200 143.300 135.800 ;
        RECT 146.200 135.600 146.600 136.800 ;
        RECT 144.500 135.300 146.600 135.600 ;
        RECT 144.500 135.200 144.900 135.300 ;
        RECT 145.300 134.900 145.700 135.000 ;
        RECT 143.800 134.600 145.700 134.900 ;
        RECT 143.800 134.500 144.200 134.600 ;
        RECT 131.100 133.900 136.600 134.200 ;
        RECT 131.300 133.800 131.700 133.900 ;
        RECT 127.800 133.300 129.700 133.600 ;
        RECT 125.500 133.100 127.300 133.300 ;
        RECT 123.000 132.800 123.900 133.100 ;
        RECT 119.000 131.800 119.700 132.200 ;
        RECT 119.300 131.500 119.700 131.800 ;
        RECT 121.400 131.500 121.800 132.500 ;
        RECT 123.500 131.100 123.900 132.800 ;
        RECT 124.600 131.100 125.000 133.100 ;
        RECT 125.400 133.000 127.400 133.100 ;
        RECT 125.400 131.100 125.800 133.000 ;
        RECT 127.000 131.100 127.400 133.000 ;
        RECT 127.800 131.100 128.200 133.300 ;
        RECT 129.300 133.200 129.700 133.300 ;
        RECT 134.200 133.200 134.500 133.900 ;
        RECT 135.800 133.800 136.600 133.900 ;
        RECT 137.800 133.900 143.300 134.200 ;
        RECT 137.800 133.800 138.600 133.900 ;
        RECT 133.300 132.700 133.700 132.800 ;
        RECT 130.200 132.100 130.600 132.500 ;
        RECT 132.300 132.400 133.700 132.700 ;
        RECT 134.200 132.400 134.600 133.200 ;
        RECT 132.300 132.100 132.600 132.400 ;
        RECT 135.000 132.100 135.400 132.500 ;
        RECT 129.900 131.800 130.600 132.100 ;
        RECT 129.900 131.100 130.500 131.800 ;
        RECT 132.200 131.100 132.600 132.100 ;
        RECT 134.400 131.800 135.400 132.100 ;
        RECT 134.400 131.100 134.800 131.800 ;
        RECT 136.600 131.100 137.000 133.500 ;
        RECT 137.400 131.100 137.800 133.500 ;
        RECT 139.900 132.800 140.200 133.900 ;
        RECT 142.700 133.800 143.100 133.900 ;
        RECT 146.200 133.600 146.600 135.300 ;
        RECT 144.700 133.300 146.600 133.600 ;
        RECT 147.000 133.400 147.400 134.200 ;
        RECT 144.700 133.200 145.100 133.300 ;
        RECT 139.000 132.100 139.400 132.500 ;
        RECT 139.800 132.400 140.200 132.800 ;
        RECT 140.700 132.700 141.100 132.800 ;
        RECT 140.700 132.400 142.100 132.700 ;
        RECT 141.800 132.100 142.100 132.400 ;
        RECT 143.800 132.100 144.200 132.500 ;
        RECT 139.000 131.800 140.000 132.100 ;
        RECT 139.600 131.100 140.000 131.800 ;
        RECT 141.800 131.100 142.200 132.100 ;
        RECT 143.800 131.800 144.500 132.100 ;
        RECT 143.900 131.100 144.500 131.800 ;
        RECT 146.200 131.100 146.600 133.300 ;
        RECT 147.800 133.100 148.200 139.900 ;
        RECT 148.600 135.800 149.000 136.600 ;
        RECT 152.900 136.400 153.300 139.900 ;
        RECT 155.000 137.500 155.400 139.500 ;
        RECT 152.500 136.100 153.300 136.400 ;
        RECT 148.600 135.100 149.000 135.200 ;
        RECT 151.800 135.100 152.200 135.600 ;
        RECT 148.600 134.800 152.200 135.100 ;
        RECT 152.500 134.200 152.800 136.100 ;
        RECT 155.100 135.800 155.400 137.500 ;
        RECT 153.500 135.500 155.400 135.800 ;
        RECT 155.800 135.700 156.200 139.900 ;
        RECT 158.000 138.200 158.400 139.900 ;
        RECT 157.400 137.900 158.400 138.200 ;
        RECT 160.200 137.900 160.600 139.900 ;
        RECT 162.300 137.900 162.900 139.900 ;
        RECT 157.400 137.500 157.800 137.900 ;
        RECT 160.200 137.600 160.500 137.900 ;
        RECT 159.100 137.300 160.900 137.600 ;
        RECT 162.200 137.500 162.600 137.900 ;
        RECT 159.100 137.200 159.500 137.300 ;
        RECT 160.500 137.200 160.900 137.300 ;
        RECT 157.400 136.500 157.800 136.600 ;
        RECT 159.700 136.500 160.100 136.600 ;
        RECT 157.400 136.200 160.100 136.500 ;
        RECT 160.400 136.500 161.500 136.800 ;
        RECT 160.400 135.900 160.700 136.500 ;
        RECT 161.100 136.400 161.500 136.500 ;
        RECT 162.300 136.600 163.000 137.000 ;
        RECT 162.300 136.100 162.600 136.600 ;
        RECT 158.300 135.700 160.700 135.900 ;
        RECT 155.800 135.600 160.700 135.700 ;
        RECT 161.400 135.800 162.600 136.100 ;
        RECT 155.800 135.500 158.700 135.600 ;
        RECT 153.500 134.500 153.800 135.500 ;
        RECT 155.800 135.400 158.600 135.500 ;
        RECT 151.800 133.800 152.800 134.200 ;
        RECT 153.100 134.100 153.800 134.500 ;
        RECT 154.200 134.400 154.600 135.200 ;
        RECT 155.000 134.400 155.400 135.200 ;
        RECT 159.000 135.100 159.400 135.200 ;
        RECT 156.900 134.800 159.400 135.100 ;
        RECT 156.900 134.700 157.300 134.800 ;
        RECT 157.700 134.200 158.100 134.300 ;
        RECT 161.400 134.200 161.700 135.800 ;
        RECT 164.600 135.600 165.000 139.900 ;
        RECT 162.900 135.300 165.000 135.600 ;
        RECT 165.400 137.500 165.800 139.500 ;
        RECT 165.400 135.800 165.700 137.500 ;
        RECT 167.500 136.400 167.900 139.900 ;
        RECT 167.500 136.100 168.300 136.400 ;
        RECT 167.800 135.800 168.300 136.100 ;
        RECT 165.400 135.500 167.300 135.800 ;
        RECT 162.900 135.200 163.300 135.300 ;
        RECT 163.700 134.900 164.100 135.000 ;
        RECT 162.200 134.600 164.100 134.900 ;
        RECT 162.200 134.500 162.600 134.600 ;
        RECT 152.500 133.500 152.800 133.800 ;
        RECT 153.300 133.900 153.800 134.100 ;
        RECT 156.200 133.900 161.700 134.200 ;
        RECT 153.300 133.600 155.400 133.900 ;
        RECT 156.200 133.800 157.000 133.900 ;
        RECT 152.500 133.300 152.900 133.500 ;
        RECT 147.800 132.800 148.700 133.100 ;
        RECT 152.500 133.000 153.300 133.300 ;
        RECT 148.300 132.200 148.700 132.800 ;
        RECT 147.800 131.800 148.700 132.200 ;
        RECT 148.300 131.100 148.700 131.800 ;
        RECT 152.900 132.200 153.300 133.000 ;
        RECT 155.100 132.500 155.400 133.600 ;
        RECT 152.900 131.800 153.800 132.200 ;
        RECT 152.900 131.500 153.300 131.800 ;
        RECT 155.000 131.500 155.400 132.500 ;
        RECT 155.800 131.100 156.200 133.500 ;
        RECT 158.300 132.800 158.600 133.900 ;
        RECT 161.100 133.800 161.500 133.900 ;
        RECT 164.600 133.600 165.000 135.300 ;
        RECT 165.400 134.400 165.800 135.200 ;
        RECT 166.200 134.400 166.600 135.200 ;
        RECT 167.000 134.500 167.300 135.500 ;
        RECT 167.000 134.100 167.700 134.500 ;
        RECT 168.000 134.200 168.300 135.800 ;
        RECT 168.600 135.100 169.000 135.600 ;
        RECT 171.000 135.100 171.400 139.900 ;
        RECT 173.000 136.800 173.400 137.200 ;
        RECT 171.800 135.800 172.200 136.600 ;
        RECT 173.000 136.200 173.300 136.800 ;
        RECT 173.700 136.200 174.100 139.900 ;
        RECT 172.600 135.900 173.300 136.200 ;
        RECT 173.600 135.900 174.100 136.200 ;
        RECT 175.800 137.500 176.200 139.500 ;
        RECT 172.600 135.800 173.000 135.900 ;
        RECT 172.600 135.100 172.900 135.800 ;
        RECT 168.600 134.800 169.700 135.100 ;
        RECT 167.000 133.900 167.500 134.100 ;
        RECT 163.100 133.300 165.000 133.600 ;
        RECT 163.100 133.200 163.500 133.300 ;
        RECT 157.400 132.100 157.800 132.500 ;
        RECT 158.200 132.400 158.600 132.800 ;
        RECT 159.100 132.700 159.500 132.800 ;
        RECT 159.100 132.400 160.500 132.700 ;
        RECT 160.200 132.100 160.500 132.400 ;
        RECT 162.200 132.100 162.600 132.500 ;
        RECT 157.400 131.800 158.400 132.100 ;
        RECT 158.000 131.100 158.400 131.800 ;
        RECT 160.200 131.100 160.600 132.100 ;
        RECT 162.200 131.800 162.900 132.100 ;
        RECT 162.300 131.100 162.900 131.800 ;
        RECT 164.600 131.100 165.000 133.300 ;
        RECT 165.400 133.600 167.500 133.900 ;
        RECT 168.000 133.800 169.000 134.200 ;
        RECT 169.400 134.100 169.700 134.800 ;
        RECT 171.000 134.800 172.900 135.100 ;
        RECT 170.200 134.100 170.600 134.200 ;
        RECT 169.400 133.800 170.600 134.100 ;
        RECT 165.400 132.500 165.700 133.600 ;
        RECT 168.000 133.500 168.300 133.800 ;
        RECT 167.900 133.300 168.300 133.500 ;
        RECT 170.200 133.400 170.600 133.800 ;
        RECT 167.500 133.000 168.300 133.300 ;
        RECT 171.000 133.100 171.400 134.800 ;
        RECT 173.600 134.200 173.900 135.900 ;
        RECT 175.800 135.800 176.100 137.500 ;
        RECT 177.900 136.400 178.300 139.900 ;
        RECT 180.600 139.600 182.600 139.900 ;
        RECT 177.900 136.100 178.700 136.400 ;
        RECT 175.800 135.500 177.700 135.800 ;
        RECT 174.200 134.400 174.600 135.200 ;
        RECT 175.800 134.400 176.200 135.200 ;
        RECT 176.600 134.400 177.000 135.200 ;
        RECT 177.400 134.500 177.700 135.500 ;
        RECT 171.800 134.100 172.200 134.200 ;
        RECT 172.600 134.100 173.900 134.200 ;
        RECT 175.000 134.100 175.400 134.200 ;
        RECT 171.800 133.800 173.900 134.100 ;
        RECT 174.600 133.800 175.400 134.100 ;
        RECT 177.400 134.100 178.100 134.500 ;
        RECT 178.400 134.200 178.700 136.100 ;
        RECT 180.600 135.900 181.000 139.600 ;
        RECT 181.400 135.900 181.800 139.300 ;
        RECT 182.200 136.200 182.600 139.600 ;
        RECT 183.800 136.200 184.200 139.900 ;
        RECT 182.200 135.900 184.200 136.200 ;
        RECT 181.500 135.600 181.800 135.900 ;
        RECT 184.600 135.800 185.000 136.600 ;
        RECT 179.000 134.800 179.400 135.600 ;
        RECT 180.600 134.800 181.000 135.600 ;
        RECT 181.500 135.300 182.500 135.600 ;
        RECT 182.200 135.200 182.500 135.300 ;
        RECT 183.400 135.200 183.800 135.400 ;
        RECT 182.200 134.800 182.600 135.200 ;
        RECT 183.400 134.900 184.200 135.200 ;
        RECT 183.800 134.800 184.200 134.900 ;
        RECT 181.500 134.400 181.900 134.800 ;
        RECT 181.500 134.200 181.800 134.400 ;
        RECT 178.400 134.100 179.400 134.200 ;
        RECT 181.400 134.100 181.800 134.200 ;
        RECT 177.400 133.900 177.900 134.100 ;
        RECT 172.700 133.100 173.000 133.800 ;
        RECT 174.600 133.600 175.000 133.800 ;
        RECT 175.800 133.600 177.900 133.900 ;
        RECT 178.400 133.800 181.800 134.100 ;
        RECT 173.500 133.100 175.300 133.300 ;
        RECT 165.400 131.500 165.800 132.500 ;
        RECT 167.500 131.500 167.900 133.000 ;
        RECT 171.000 132.800 171.900 133.100 ;
        RECT 171.500 131.100 171.900 132.800 ;
        RECT 172.600 131.100 173.000 133.100 ;
        RECT 173.400 133.000 175.400 133.100 ;
        RECT 173.400 131.100 173.800 133.000 ;
        RECT 175.000 131.100 175.400 133.000 ;
        RECT 175.800 132.500 176.100 133.600 ;
        RECT 178.400 133.500 178.700 133.800 ;
        RECT 178.300 133.300 178.700 133.500 ;
        RECT 177.900 133.000 178.700 133.300 ;
        RECT 182.200 133.100 182.500 134.800 ;
        RECT 183.000 133.800 183.400 134.600 ;
        RECT 185.400 133.100 185.800 139.900 ;
        RECT 187.000 136.200 187.400 139.900 ;
        RECT 188.600 136.400 189.000 139.900 ;
        RECT 192.100 136.400 192.500 139.900 ;
        RECT 194.200 137.500 194.600 139.500 ;
        RECT 187.000 135.900 188.300 136.200 ;
        RECT 188.600 135.900 189.100 136.400 ;
        RECT 187.000 134.800 187.500 135.200 ;
        RECT 187.100 134.400 187.500 134.800 ;
        RECT 188.000 134.900 188.300 135.900 ;
        RECT 188.000 134.500 188.500 134.900 ;
        RECT 186.200 133.400 186.600 134.200 ;
        RECT 188.000 133.700 188.300 134.500 ;
        RECT 188.800 134.200 189.100 135.900 ;
        RECT 191.700 136.100 192.500 136.400 ;
        RECT 191.000 134.800 191.400 135.600 ;
        RECT 191.700 134.200 192.000 136.100 ;
        RECT 194.300 135.800 194.600 137.500 ;
        RECT 196.300 136.200 196.700 139.900 ;
        RECT 197.000 136.800 197.400 137.200 ;
        RECT 197.100 136.200 197.400 136.800 ;
        RECT 196.300 135.900 196.800 136.200 ;
        RECT 197.100 135.900 197.800 136.200 ;
        RECT 192.700 135.500 194.600 135.800 ;
        RECT 192.700 134.500 193.000 135.500 ;
        RECT 188.600 133.800 189.100 134.200 ;
        RECT 189.400 134.100 189.800 134.200 ;
        RECT 191.000 134.100 192.000 134.200 ;
        RECT 192.300 134.100 193.000 134.500 ;
        RECT 193.400 134.400 193.800 135.200 ;
        RECT 194.200 134.400 194.600 135.200 ;
        RECT 195.800 134.400 196.200 135.200 ;
        RECT 196.500 134.200 196.800 135.900 ;
        RECT 197.400 135.800 197.800 135.900 ;
        RECT 198.200 135.800 198.600 136.600 ;
        RECT 197.400 135.100 197.700 135.800 ;
        RECT 199.000 135.100 199.400 139.900 ;
        RECT 201.400 137.100 201.800 137.200 ;
        RECT 202.200 137.100 202.600 139.900 ;
        RECT 204.300 137.900 204.900 139.900 ;
        RECT 206.600 137.900 207.000 139.900 ;
        RECT 208.800 138.200 209.200 139.900 ;
        RECT 208.800 137.900 209.800 138.200 ;
        RECT 204.600 137.500 205.000 137.900 ;
        RECT 206.700 137.600 207.000 137.900 ;
        RECT 206.300 137.300 208.100 137.600 ;
        RECT 209.400 137.500 209.800 137.900 ;
        RECT 206.300 137.200 206.700 137.300 ;
        RECT 207.700 137.200 208.100 137.300 ;
        RECT 201.400 136.800 202.600 137.100 ;
        RECT 197.400 134.800 199.400 135.100 ;
        RECT 189.400 133.800 192.000 134.100 ;
        RECT 187.000 133.400 188.300 133.700 ;
        RECT 175.800 131.500 176.200 132.500 ;
        RECT 177.900 131.500 178.300 133.000 ;
        RECT 181.900 131.100 182.700 133.100 ;
        RECT 184.900 132.800 185.800 133.100 ;
        RECT 184.900 132.200 185.300 132.800 ;
        RECT 184.600 131.800 185.300 132.200 ;
        RECT 184.900 131.100 185.300 131.800 ;
        RECT 187.000 131.100 187.400 133.400 ;
        RECT 188.800 133.100 189.100 133.800 ;
        RECT 188.600 132.800 189.100 133.100 ;
        RECT 191.700 133.500 192.000 133.800 ;
        RECT 192.500 133.900 193.000 134.100 ;
        RECT 195.000 134.100 195.400 134.200 ;
        RECT 196.500 134.100 197.800 134.200 ;
        RECT 198.200 134.100 198.600 134.200 ;
        RECT 192.500 133.600 194.600 133.900 ;
        RECT 195.000 133.800 195.800 134.100 ;
        RECT 196.500 133.800 198.600 134.100 ;
        RECT 195.400 133.600 195.800 133.800 ;
        RECT 191.700 133.300 192.100 133.500 ;
        RECT 191.700 133.000 192.500 133.300 ;
        RECT 188.600 131.100 189.000 132.800 ;
        RECT 192.100 131.500 192.500 133.000 ;
        RECT 194.300 132.500 194.600 133.600 ;
        RECT 195.100 133.100 196.900 133.300 ;
        RECT 197.400 133.100 197.700 133.800 ;
        RECT 199.000 133.100 199.400 134.800 ;
        RECT 202.200 135.600 202.600 136.800 ;
        RECT 204.200 136.600 204.900 137.000 ;
        RECT 204.600 136.100 204.900 136.600 ;
        RECT 205.700 136.500 206.800 136.800 ;
        RECT 205.700 136.400 206.100 136.500 ;
        RECT 204.600 135.800 205.800 136.100 ;
        RECT 202.200 135.300 204.300 135.600 ;
        RECT 199.800 134.100 200.200 134.200 ;
        RECT 201.400 134.100 201.800 134.200 ;
        RECT 199.800 133.800 201.800 134.100 ;
        RECT 199.800 133.400 200.200 133.800 ;
        RECT 202.200 133.600 202.600 135.300 ;
        RECT 203.900 135.200 204.300 135.300 ;
        RECT 203.100 134.900 203.500 135.000 ;
        RECT 203.100 134.600 205.000 134.900 ;
        RECT 204.600 134.500 205.000 134.600 ;
        RECT 205.500 134.200 205.800 135.800 ;
        RECT 206.500 135.900 206.800 136.500 ;
        RECT 207.100 136.500 207.500 136.600 ;
        RECT 209.400 136.500 209.800 136.600 ;
        RECT 207.100 136.200 209.800 136.500 ;
        RECT 206.500 135.700 208.900 135.900 ;
        RECT 211.000 135.700 211.400 139.900 ;
        RECT 206.500 135.600 211.400 135.700 ;
        RECT 208.500 135.500 211.400 135.600 ;
        RECT 208.600 135.400 211.400 135.500 ;
        RECT 207.800 135.100 208.200 135.200 ;
        RECT 212.600 135.100 213.000 139.900 ;
        RECT 214.600 136.800 215.000 137.200 ;
        RECT 213.400 135.800 213.800 136.600 ;
        RECT 214.600 136.200 214.900 136.800 ;
        RECT 215.300 136.200 215.700 139.900 ;
        RECT 214.200 135.900 214.900 136.200 ;
        RECT 215.200 135.900 215.700 136.200 ;
        RECT 214.200 135.800 214.600 135.900 ;
        RECT 214.200 135.100 214.500 135.800 ;
        RECT 215.200 135.200 215.500 135.900 ;
        RECT 217.400 135.600 217.800 139.900 ;
        RECT 219.500 137.900 220.100 139.900 ;
        RECT 221.800 137.900 222.200 139.900 ;
        RECT 224.000 138.200 224.400 139.900 ;
        RECT 224.000 137.900 225.000 138.200 ;
        RECT 219.800 137.500 220.200 137.900 ;
        RECT 221.900 137.600 222.200 137.900 ;
        RECT 221.500 137.300 223.300 137.600 ;
        RECT 224.600 137.500 225.000 137.900 ;
        RECT 221.500 137.200 221.900 137.300 ;
        RECT 222.900 137.200 223.300 137.300 ;
        RECT 219.000 137.000 219.700 137.200 ;
        RECT 219.000 136.800 220.100 137.000 ;
        RECT 219.400 136.600 220.100 136.800 ;
        RECT 219.800 136.100 220.100 136.600 ;
        RECT 220.900 136.500 222.000 136.800 ;
        RECT 220.900 136.400 221.300 136.500 ;
        RECT 219.800 135.800 221.000 136.100 ;
        RECT 217.400 135.300 219.500 135.600 ;
        RECT 207.800 134.800 210.300 135.100 ;
        RECT 209.900 134.700 210.300 134.800 ;
        RECT 212.600 134.800 214.500 135.100 ;
        RECT 215.000 134.800 215.500 135.200 ;
        RECT 209.100 134.200 209.500 134.300 ;
        RECT 205.500 133.900 211.000 134.200 ;
        RECT 205.700 133.800 206.100 133.900 ;
        RECT 207.000 133.800 207.400 133.900 ;
        RECT 194.200 131.500 194.600 132.500 ;
        RECT 195.000 133.000 197.000 133.100 ;
        RECT 195.000 131.100 195.400 133.000 ;
        RECT 196.600 131.100 197.000 133.000 ;
        RECT 197.400 131.100 197.800 133.100 ;
        RECT 198.500 132.800 199.400 133.100 ;
        RECT 202.200 133.300 204.100 133.600 ;
        RECT 198.500 131.100 198.900 132.800 ;
        RECT 202.200 131.100 202.600 133.300 ;
        RECT 203.700 133.200 204.100 133.300 ;
        RECT 208.600 132.800 208.900 133.900 ;
        RECT 210.200 133.800 211.000 133.900 ;
        RECT 207.700 132.700 208.100 132.800 ;
        RECT 204.600 132.100 205.000 132.500 ;
        RECT 206.700 132.400 208.100 132.700 ;
        RECT 208.600 132.400 209.000 132.800 ;
        RECT 206.700 132.100 207.000 132.400 ;
        RECT 209.400 132.100 209.800 132.500 ;
        RECT 204.300 131.800 205.000 132.100 ;
        RECT 204.300 131.100 204.900 131.800 ;
        RECT 206.600 131.100 207.000 132.100 ;
        RECT 208.800 131.800 209.800 132.100 ;
        RECT 208.800 131.100 209.200 131.800 ;
        RECT 211.000 131.100 211.400 133.500 ;
        RECT 211.800 133.400 212.200 134.200 ;
        RECT 212.600 133.100 213.000 134.800 ;
        RECT 215.200 134.200 215.500 134.800 ;
        RECT 215.800 134.400 216.200 135.200 ;
        RECT 214.200 133.800 215.500 134.200 ;
        RECT 216.600 134.100 217.000 134.200 ;
        RECT 216.200 133.800 217.000 134.100 ;
        RECT 214.300 133.100 214.600 133.800 ;
        RECT 216.200 133.600 216.600 133.800 ;
        RECT 217.400 133.600 217.800 135.300 ;
        RECT 219.100 135.200 219.500 135.300 ;
        RECT 218.300 134.900 218.700 135.000 ;
        RECT 218.300 134.600 220.200 134.900 ;
        RECT 219.800 134.500 220.200 134.600 ;
        RECT 220.700 134.200 221.000 135.800 ;
        RECT 221.700 135.900 222.000 136.500 ;
        RECT 222.300 136.500 222.700 136.600 ;
        RECT 224.600 136.500 225.000 136.600 ;
        RECT 222.300 136.200 225.000 136.500 ;
        RECT 221.700 135.700 224.100 135.900 ;
        RECT 226.200 135.700 226.600 139.900 ;
        RECT 221.700 135.600 226.600 135.700 ;
        RECT 223.700 135.500 226.600 135.600 ;
        RECT 223.800 135.400 226.600 135.500 ;
        RECT 227.000 135.600 227.400 139.900 ;
        RECT 229.100 137.900 229.700 139.900 ;
        RECT 231.400 137.900 231.800 139.900 ;
        RECT 233.600 138.200 234.000 139.900 ;
        RECT 233.600 137.900 234.600 138.200 ;
        RECT 229.400 137.500 229.800 137.900 ;
        RECT 231.500 137.600 231.800 137.900 ;
        RECT 231.100 137.300 232.900 137.600 ;
        RECT 234.200 137.500 234.600 137.900 ;
        RECT 231.100 137.200 231.500 137.300 ;
        RECT 232.500 137.200 232.900 137.300 ;
        RECT 229.000 136.600 229.700 137.000 ;
        RECT 229.400 136.100 229.700 136.600 ;
        RECT 230.500 136.500 231.600 136.800 ;
        RECT 230.500 136.400 230.900 136.500 ;
        RECT 229.400 135.800 230.600 136.100 ;
        RECT 227.000 135.300 229.100 135.600 ;
        RECT 223.000 135.100 223.400 135.200 ;
        RECT 223.000 134.800 225.500 135.100 ;
        RECT 225.100 134.700 225.500 134.800 ;
        RECT 224.300 134.200 224.700 134.300 ;
        RECT 220.700 133.900 226.200 134.200 ;
        RECT 220.900 133.800 221.300 133.900 ;
        RECT 217.400 133.300 219.300 133.600 ;
        RECT 215.100 133.100 216.900 133.300 ;
        RECT 212.600 132.800 213.500 133.100 ;
        RECT 213.100 131.100 213.500 132.800 ;
        RECT 214.200 131.100 214.600 133.100 ;
        RECT 215.000 133.000 217.000 133.100 ;
        RECT 215.000 131.100 215.400 133.000 ;
        RECT 216.600 131.100 217.000 133.000 ;
        RECT 217.400 131.100 217.800 133.300 ;
        RECT 218.900 133.200 219.300 133.300 ;
        RECT 223.800 132.800 224.100 133.900 ;
        RECT 225.400 133.800 226.200 133.900 ;
        RECT 227.000 133.600 227.400 135.300 ;
        RECT 228.700 135.200 229.100 135.300 ;
        RECT 230.300 135.200 230.600 135.800 ;
        RECT 231.300 135.900 231.600 136.500 ;
        RECT 231.900 136.500 232.300 136.600 ;
        RECT 234.200 136.500 234.600 136.600 ;
        RECT 231.900 136.200 234.600 136.500 ;
        RECT 231.300 135.700 233.700 135.900 ;
        RECT 235.800 135.700 236.200 139.900 ;
        RECT 237.000 136.800 237.400 137.200 ;
        RECT 237.000 136.200 237.300 136.800 ;
        RECT 237.700 136.200 238.100 139.900 ;
        RECT 240.600 136.400 241.000 139.900 ;
        RECT 236.600 135.900 237.300 136.200 ;
        RECT 237.600 135.900 238.100 136.200 ;
        RECT 240.500 135.900 241.000 136.400 ;
        RECT 242.200 136.200 242.600 139.900 ;
        RECT 241.300 135.900 242.600 136.200 ;
        RECT 236.600 135.800 237.000 135.900 ;
        RECT 231.300 135.600 236.200 135.700 ;
        RECT 233.300 135.500 236.200 135.600 ;
        RECT 233.400 135.400 236.200 135.500 ;
        RECT 237.600 135.200 237.900 135.900 ;
        RECT 227.900 134.900 228.300 135.000 ;
        RECT 227.900 134.600 229.800 134.900 ;
        RECT 230.200 134.800 230.600 135.200 ;
        RECT 232.600 135.100 233.000 135.200 ;
        RECT 232.600 134.800 235.100 135.100 ;
        RECT 237.400 134.800 237.900 135.200 ;
        RECT 229.400 134.500 229.800 134.600 ;
        RECT 230.300 134.200 230.600 134.800 ;
        RECT 233.400 134.700 233.800 134.800 ;
        RECT 234.700 134.700 235.100 134.800 ;
        RECT 233.900 134.200 234.300 134.300 ;
        RECT 237.600 134.200 237.900 134.800 ;
        RECT 238.200 134.400 238.600 135.200 ;
        RECT 240.500 134.200 240.800 135.900 ;
        RECT 241.300 134.900 241.600 135.900 ;
        RECT 243.800 135.600 244.200 139.900 ;
        RECT 245.400 135.600 245.800 139.900 ;
        RECT 247.000 135.600 247.400 139.900 ;
        RECT 248.600 135.600 249.000 139.900 ;
        RECT 243.000 135.200 244.200 135.600 ;
        RECT 244.700 135.200 245.800 135.600 ;
        RECT 246.300 135.200 247.400 135.600 ;
        RECT 248.100 135.200 249.000 135.600 ;
        RECT 241.100 134.500 241.600 134.900 ;
        RECT 230.300 133.900 235.800 134.200 ;
        RECT 230.500 133.800 230.900 133.900 ;
        RECT 222.900 132.700 223.300 132.800 ;
        RECT 219.800 132.100 220.200 132.500 ;
        RECT 221.900 132.400 223.300 132.700 ;
        RECT 223.800 132.400 224.200 132.800 ;
        RECT 221.900 132.100 222.200 132.400 ;
        RECT 224.600 132.100 225.000 132.500 ;
        RECT 219.500 131.800 220.200 132.100 ;
        RECT 219.500 131.100 220.100 131.800 ;
        RECT 221.800 131.100 222.200 132.100 ;
        RECT 224.000 131.800 225.000 132.100 ;
        RECT 224.000 131.100 224.400 131.800 ;
        RECT 226.200 131.100 226.600 133.500 ;
        RECT 227.000 133.300 228.900 133.600 ;
        RECT 227.000 131.100 227.400 133.300 ;
        RECT 228.500 133.200 228.900 133.300 ;
        RECT 233.400 132.800 233.700 133.900 ;
        RECT 235.000 133.800 235.800 133.900 ;
        RECT 236.600 133.800 237.900 134.200 ;
        RECT 239.000 134.100 239.400 134.200 ;
        RECT 240.500 134.100 241.000 134.200 ;
        RECT 238.600 133.800 241.000 134.100 ;
        RECT 232.500 132.700 232.900 132.800 ;
        RECT 229.400 132.100 229.800 132.500 ;
        RECT 231.500 132.400 232.900 132.700 ;
        RECT 233.400 132.400 233.800 132.800 ;
        RECT 231.500 132.100 231.800 132.400 ;
        RECT 234.200 132.100 234.600 132.500 ;
        RECT 229.100 131.800 229.800 132.100 ;
        RECT 229.100 131.100 229.700 131.800 ;
        RECT 231.400 131.100 231.800 132.100 ;
        RECT 233.600 131.800 234.600 132.100 ;
        RECT 233.600 131.100 234.000 131.800 ;
        RECT 235.800 131.100 236.200 133.500 ;
        RECT 236.700 133.100 237.000 133.800 ;
        RECT 238.600 133.600 239.000 133.800 ;
        RECT 237.500 133.100 239.300 133.300 ;
        RECT 240.500 133.100 240.800 133.800 ;
        RECT 241.300 133.700 241.600 134.500 ;
        RECT 242.100 134.800 242.600 135.200 ;
        RECT 242.100 134.400 242.500 134.800 ;
        RECT 243.000 133.800 243.400 135.200 ;
        RECT 244.700 134.500 245.100 135.200 ;
        RECT 246.300 134.500 246.700 135.200 ;
        RECT 248.100 134.500 248.500 135.200 ;
        RECT 243.800 134.100 245.100 134.500 ;
        RECT 245.500 134.100 246.700 134.500 ;
        RECT 247.200 134.100 248.500 134.500 ;
        RECT 248.900 134.100 249.800 134.500 ;
        RECT 244.700 133.800 245.100 134.100 ;
        RECT 246.300 133.800 246.700 134.100 ;
        RECT 248.100 133.800 248.500 134.100 ;
        RECT 249.400 133.800 249.800 134.100 ;
        RECT 241.300 133.400 242.600 133.700 ;
        RECT 243.000 133.400 244.200 133.800 ;
        RECT 244.700 133.400 245.800 133.800 ;
        RECT 246.300 133.400 247.400 133.800 ;
        RECT 248.100 133.400 249.000 133.800 ;
        RECT 236.600 131.100 237.000 133.100 ;
        RECT 237.400 133.000 239.400 133.100 ;
        RECT 237.400 131.100 237.800 133.000 ;
        RECT 239.000 131.100 239.400 133.000 ;
        RECT 240.500 132.800 241.000 133.100 ;
        RECT 240.600 131.100 241.000 132.800 ;
        RECT 242.200 131.100 242.600 133.400 ;
        RECT 243.800 131.100 244.200 133.400 ;
        RECT 245.400 131.100 245.800 133.400 ;
        RECT 247.000 131.100 247.400 133.400 ;
        RECT 248.600 131.100 249.000 133.400 ;
        RECT 0.600 127.500 1.000 129.900 ;
        RECT 2.800 129.200 3.200 129.900 ;
        RECT 2.200 128.900 3.200 129.200 ;
        RECT 5.000 128.900 5.400 129.900 ;
        RECT 7.100 129.200 7.700 129.900 ;
        RECT 7.000 128.900 7.700 129.200 ;
        RECT 2.200 128.500 2.600 128.900 ;
        RECT 5.000 128.600 5.300 128.900 ;
        RECT 3.000 128.200 3.400 128.600 ;
        RECT 3.900 128.300 5.300 128.600 ;
        RECT 7.000 128.500 7.400 128.900 ;
        RECT 3.900 128.200 4.300 128.300 ;
        RECT 1.000 127.100 1.800 127.200 ;
        RECT 3.100 127.100 3.400 128.200 ;
        RECT 7.900 127.700 8.300 127.800 ;
        RECT 9.400 127.700 9.800 129.900 ;
        RECT 10.500 128.200 10.900 129.900 ;
        RECT 10.500 127.900 11.400 128.200 ;
        RECT 12.600 127.900 13.000 129.900 ;
        RECT 13.400 128.000 13.800 129.900 ;
        RECT 15.000 128.000 15.400 129.900 ;
        RECT 13.400 127.900 15.400 128.000 ;
        RECT 15.800 128.000 16.200 129.900 ;
        RECT 17.400 128.000 17.800 129.900 ;
        RECT 15.800 127.900 17.800 128.000 ;
        RECT 18.200 127.900 18.600 129.900 ;
        RECT 7.900 127.400 9.800 127.700 ;
        RECT 5.900 127.100 6.300 127.200 ;
        RECT 1.000 126.800 6.500 127.100 ;
        RECT 2.500 126.700 2.900 126.800 ;
        RECT 1.700 126.200 2.100 126.300 ;
        RECT 1.700 126.100 4.200 126.200 ;
        RECT 5.400 126.100 5.800 126.200 ;
        RECT 1.700 125.900 5.800 126.100 ;
        RECT 3.800 125.800 5.800 125.900 ;
        RECT 0.600 125.500 3.400 125.600 ;
        RECT 0.600 125.400 3.500 125.500 ;
        RECT 0.600 125.300 5.500 125.400 ;
        RECT 0.600 121.100 1.000 125.300 ;
        RECT 3.100 125.100 5.500 125.300 ;
        RECT 2.200 124.500 4.900 124.800 ;
        RECT 2.200 124.400 2.600 124.500 ;
        RECT 4.500 124.400 4.900 124.500 ;
        RECT 5.200 124.500 5.500 125.100 ;
        RECT 6.200 125.200 6.500 126.800 ;
        RECT 7.000 126.400 7.400 126.500 ;
        RECT 7.000 126.100 8.900 126.400 ;
        RECT 8.500 126.000 8.900 126.100 ;
        RECT 7.700 125.700 8.100 125.800 ;
        RECT 9.400 125.700 9.800 127.400 ;
        RECT 7.700 125.400 9.800 125.700 ;
        RECT 6.200 124.900 7.400 125.200 ;
        RECT 5.900 124.500 6.300 124.600 ;
        RECT 5.200 124.200 6.300 124.500 ;
        RECT 7.100 124.400 7.400 124.900 ;
        RECT 7.100 124.000 7.800 124.400 ;
        RECT 3.900 123.700 4.300 123.800 ;
        RECT 5.300 123.700 5.700 123.800 ;
        RECT 2.200 123.100 2.600 123.500 ;
        RECT 3.900 123.400 5.700 123.700 ;
        RECT 5.000 123.100 5.300 123.400 ;
        RECT 7.000 123.100 7.400 123.500 ;
        RECT 2.200 122.800 3.200 123.100 ;
        RECT 2.800 121.100 3.200 122.800 ;
        RECT 5.000 121.100 5.400 123.100 ;
        RECT 7.100 121.100 7.700 123.100 ;
        RECT 9.400 121.100 9.800 125.400 ;
        RECT 10.200 124.400 10.600 125.200 ;
        RECT 11.000 125.100 11.400 127.900 ;
        RECT 11.800 126.800 12.200 127.600 ;
        RECT 12.700 127.200 13.000 127.900 ;
        RECT 13.500 127.700 15.300 127.900 ;
        RECT 15.900 127.700 17.700 127.900 ;
        RECT 14.600 127.200 15.000 127.400 ;
        RECT 16.200 127.200 16.600 127.400 ;
        RECT 18.200 127.200 18.500 127.900 ;
        RECT 19.000 127.500 19.400 129.900 ;
        RECT 21.200 129.200 21.600 129.900 ;
        RECT 20.600 128.900 21.600 129.200 ;
        RECT 23.400 128.900 23.800 129.900 ;
        RECT 25.500 129.200 26.100 129.900 ;
        RECT 25.400 128.900 26.100 129.200 ;
        RECT 20.600 128.500 21.000 128.900 ;
        RECT 23.400 128.600 23.700 128.900 ;
        RECT 21.400 128.200 21.800 128.600 ;
        RECT 22.300 128.300 23.700 128.600 ;
        RECT 25.400 128.500 25.800 128.900 ;
        RECT 22.300 128.200 22.700 128.300 ;
        RECT 21.500 127.200 21.800 128.200 ;
        RECT 26.300 127.700 26.700 127.800 ;
        RECT 27.800 127.700 28.200 129.900 ;
        RECT 30.500 128.000 30.900 129.500 ;
        RECT 32.600 128.500 33.000 129.500 ;
        RECT 26.300 127.400 28.200 127.700 ;
        RECT 12.600 126.800 13.900 127.200 ;
        RECT 14.600 126.900 15.400 127.200 ;
        RECT 15.000 126.800 15.400 126.900 ;
        RECT 15.800 126.900 16.600 127.200 ;
        RECT 15.800 126.800 16.200 126.900 ;
        RECT 17.300 126.800 18.600 127.200 ;
        RECT 19.400 127.100 20.200 127.200 ;
        RECT 21.400 127.100 21.800 127.200 ;
        RECT 24.300 127.100 24.700 127.200 ;
        RECT 19.400 126.800 24.900 127.100 ;
        RECT 12.600 125.100 13.000 125.200 ;
        RECT 13.600 125.100 13.900 126.800 ;
        RECT 14.200 125.800 14.600 126.600 ;
        RECT 16.600 125.800 17.000 126.600 ;
        RECT 17.300 125.100 17.600 126.800 ;
        RECT 20.900 126.700 21.300 126.800 ;
        RECT 20.100 126.200 20.500 126.300 ;
        RECT 20.100 125.900 22.600 126.200 ;
        RECT 22.200 125.800 22.600 125.900 ;
        RECT 19.000 125.500 21.800 125.600 ;
        RECT 19.000 125.400 21.900 125.500 ;
        RECT 19.000 125.300 23.900 125.400 ;
        RECT 18.200 125.100 18.600 125.200 ;
        RECT 11.000 124.800 13.300 125.100 ;
        RECT 13.600 124.800 14.100 125.100 ;
        RECT 11.000 121.100 11.400 124.800 ;
        RECT 13.000 124.200 13.300 124.800 ;
        RECT 13.000 123.800 13.400 124.200 ;
        RECT 13.700 121.100 14.100 124.800 ;
        RECT 17.100 124.800 17.600 125.100 ;
        RECT 17.900 124.800 18.600 125.100 ;
        RECT 17.100 121.100 17.500 124.800 ;
        RECT 17.900 124.200 18.200 124.800 ;
        RECT 17.800 123.800 18.200 124.200 ;
        RECT 19.000 121.100 19.400 125.300 ;
        RECT 21.500 125.100 23.900 125.300 ;
        RECT 20.600 124.500 23.300 124.800 ;
        RECT 20.600 124.400 21.000 124.500 ;
        RECT 22.900 124.400 23.300 124.500 ;
        RECT 23.600 124.500 23.900 125.100 ;
        RECT 24.600 125.200 24.900 126.800 ;
        RECT 25.400 126.400 25.800 126.500 ;
        RECT 25.400 126.100 27.300 126.400 ;
        RECT 26.900 126.000 27.300 126.100 ;
        RECT 26.100 125.700 26.500 125.800 ;
        RECT 27.800 125.700 28.200 127.400 ;
        RECT 30.100 127.700 30.900 128.000 ;
        RECT 30.100 127.500 30.500 127.700 ;
        RECT 30.100 127.200 30.400 127.500 ;
        RECT 32.700 127.400 33.000 128.500 ;
        RECT 29.400 126.800 30.400 127.200 ;
        RECT 30.900 127.100 33.000 127.400 ;
        RECT 33.400 128.500 33.800 129.500 ;
        RECT 33.400 127.400 33.700 128.500 ;
        RECT 35.500 128.000 35.900 129.500 ;
        RECT 38.200 128.500 38.600 129.500 ;
        RECT 35.500 127.700 36.300 128.000 ;
        RECT 35.900 127.500 36.300 127.700 ;
        RECT 33.400 127.100 35.500 127.400 ;
        RECT 30.900 126.900 31.400 127.100 ;
        RECT 30.100 126.200 30.400 126.800 ;
        RECT 30.700 126.500 31.400 126.900 ;
        RECT 35.000 126.900 35.500 127.100 ;
        RECT 36.000 127.200 36.300 127.500 ;
        RECT 38.200 127.400 38.500 128.500 ;
        RECT 40.300 128.000 40.700 129.500 ;
        RECT 43.800 128.900 44.200 129.900 ;
        RECT 43.800 128.200 44.100 128.900 ;
        RECT 40.300 127.700 41.100 128.000 ;
        RECT 40.700 127.500 41.100 127.700 ;
        RECT 36.000 127.100 37.000 127.200 ;
        RECT 37.400 127.100 37.800 127.200 ;
        RECT 38.200 127.100 40.300 127.400 ;
        RECT 28.600 126.100 29.000 126.200 ;
        RECT 29.400 126.100 29.800 126.200 ;
        RECT 28.600 125.800 29.800 126.100 ;
        RECT 26.100 125.400 28.200 125.700 ;
        RECT 29.400 125.400 29.800 125.800 ;
        RECT 30.100 125.800 30.600 126.200 ;
        RECT 24.600 124.900 25.800 125.200 ;
        RECT 24.300 124.500 24.700 124.600 ;
        RECT 23.600 124.200 24.700 124.500 ;
        RECT 25.500 124.400 25.800 124.900 ;
        RECT 25.500 124.000 26.200 124.400 ;
        RECT 22.300 123.700 22.700 123.800 ;
        RECT 23.700 123.700 24.100 123.800 ;
        RECT 20.600 123.100 21.000 123.500 ;
        RECT 22.300 123.400 24.100 123.700 ;
        RECT 23.400 123.100 23.700 123.400 ;
        RECT 25.400 123.100 25.800 123.500 ;
        RECT 20.600 122.800 21.600 123.100 ;
        RECT 21.200 121.100 21.600 122.800 ;
        RECT 23.400 121.100 23.800 123.100 ;
        RECT 25.500 121.100 26.100 123.100 ;
        RECT 27.800 121.100 28.200 125.400 ;
        RECT 30.100 124.900 30.400 125.800 ;
        RECT 31.100 125.500 31.400 126.500 ;
        RECT 31.800 125.800 32.200 126.600 ;
        RECT 32.600 125.800 33.000 126.600 ;
        RECT 33.400 125.800 33.800 126.600 ;
        RECT 34.200 125.800 34.600 126.600 ;
        RECT 35.000 126.500 35.700 126.900 ;
        RECT 36.000 126.800 37.800 127.100 ;
        RECT 39.800 126.900 40.300 127.100 ;
        RECT 40.800 127.200 41.100 127.500 ;
        RECT 43.800 127.800 44.200 128.200 ;
        RECT 44.600 127.800 45.000 128.600 ;
        RECT 45.500 128.200 45.900 128.600 ;
        RECT 45.400 127.800 45.800 128.200 ;
        RECT 46.200 127.900 46.600 129.900 ;
        RECT 48.600 129.100 49.000 129.200 ;
        RECT 50.200 129.100 50.600 129.900 ;
        RECT 48.600 128.800 50.600 129.100 ;
        RECT 52.300 129.200 52.900 129.900 ;
        RECT 52.300 128.900 53.000 129.200 ;
        RECT 54.600 128.900 55.000 129.900 ;
        RECT 56.800 129.200 57.200 129.900 ;
        RECT 56.800 128.900 57.800 129.200 ;
        RECT 43.800 127.200 44.100 127.800 ;
        RECT 40.800 127.100 41.800 127.200 ;
        RECT 43.000 127.100 43.400 127.200 ;
        RECT 35.000 125.500 35.300 126.500 ;
        RECT 31.100 125.200 33.000 125.500 ;
        RECT 30.100 124.600 30.900 124.900 ;
        RECT 30.500 121.100 30.900 124.600 ;
        RECT 32.700 123.500 33.000 125.200 ;
        RECT 32.600 121.500 33.000 123.500 ;
        RECT 33.400 125.200 35.300 125.500 ;
        RECT 33.400 123.500 33.700 125.200 ;
        RECT 36.000 124.900 36.300 126.800 ;
        RECT 36.600 125.400 37.000 126.200 ;
        RECT 38.200 125.800 38.600 126.600 ;
        RECT 39.000 125.800 39.400 126.600 ;
        RECT 39.800 126.500 40.500 126.900 ;
        RECT 40.800 126.800 43.400 127.100 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 39.800 125.500 40.100 126.500 ;
        RECT 35.500 124.600 36.300 124.900 ;
        RECT 38.200 125.200 40.100 125.500 ;
        RECT 33.400 121.500 33.800 123.500 ;
        RECT 35.500 121.100 35.900 124.600 ;
        RECT 38.200 123.500 38.500 125.200 ;
        RECT 40.800 124.900 41.100 126.800 ;
        RECT 41.400 126.100 41.800 126.200 ;
        RECT 42.200 126.100 42.600 126.200 ;
        RECT 41.400 125.800 42.600 126.100 ;
        RECT 41.400 125.400 41.800 125.800 ;
        RECT 43.000 125.400 43.400 126.200 ;
        RECT 43.800 125.100 44.100 126.800 ;
        RECT 46.300 126.200 46.600 127.900 ;
        RECT 50.200 127.700 50.600 128.800 ;
        RECT 52.600 128.500 53.000 128.900 ;
        RECT 54.700 128.600 55.000 128.900 ;
        RECT 54.700 128.300 56.100 128.600 ;
        RECT 55.700 128.200 56.100 128.300 ;
        RECT 56.600 128.200 57.000 128.600 ;
        RECT 57.400 128.500 57.800 128.900 ;
        RECT 51.700 127.700 52.100 127.800 ;
        RECT 50.200 127.400 52.100 127.700 ;
        RECT 47.000 126.400 47.400 127.200 ;
        RECT 45.400 126.100 45.800 126.200 ;
        RECT 46.200 126.100 46.600 126.200 ;
        RECT 47.800 126.100 48.200 126.200 ;
        RECT 49.400 126.100 49.800 126.200 ;
        RECT 45.400 125.800 46.600 126.100 ;
        RECT 47.400 125.800 49.800 126.100 ;
        RECT 45.500 125.100 45.800 125.800 ;
        RECT 47.400 125.600 47.800 125.800 ;
        RECT 50.200 125.700 50.600 127.400 ;
        RECT 53.700 127.100 54.100 127.200 ;
        RECT 56.600 127.100 56.900 128.200 ;
        RECT 59.000 127.500 59.400 129.900 ;
        RECT 61.100 128.200 61.500 129.900 ;
        RECT 60.600 127.900 61.500 128.200 ;
        RECT 62.200 127.900 62.600 129.900 ;
        RECT 63.000 128.000 63.400 129.900 ;
        RECT 64.600 128.000 65.000 129.900 ;
        RECT 63.000 127.900 65.000 128.000 ;
        RECT 58.200 127.100 59.000 127.200 ;
        RECT 53.500 126.800 59.000 127.100 ;
        RECT 59.800 126.800 60.200 127.600 ;
        RECT 52.600 126.400 53.000 126.500 ;
        RECT 51.100 126.100 53.000 126.400 ;
        RECT 51.100 126.000 51.500 126.100 ;
        RECT 51.900 125.700 52.300 125.800 ;
        RECT 50.200 125.400 52.300 125.700 ;
        RECT 40.300 124.600 41.100 124.900 ;
        RECT 43.300 124.700 44.200 125.100 ;
        RECT 38.200 121.500 38.600 123.500 ;
        RECT 40.300 121.100 40.700 124.600 ;
        RECT 43.300 121.100 43.700 124.700 ;
        RECT 45.400 121.100 45.800 125.100 ;
        RECT 46.200 124.800 48.200 125.100 ;
        RECT 46.200 121.100 46.600 124.800 ;
        RECT 47.800 121.100 48.200 124.800 ;
        RECT 50.200 121.100 50.600 125.400 ;
        RECT 53.500 125.200 53.800 126.800 ;
        RECT 57.100 126.700 57.500 126.800 ;
        RECT 57.900 126.200 58.300 126.300 ;
        RECT 55.800 125.900 58.300 126.200 ;
        RECT 60.600 126.100 61.000 127.900 ;
        RECT 62.300 127.200 62.600 127.900 ;
        RECT 63.100 127.700 64.900 127.900 ;
        RECT 65.400 127.600 65.800 129.900 ;
        RECT 67.000 128.200 67.400 129.900 ;
        RECT 67.000 127.900 67.500 128.200 ;
        RECT 64.200 127.200 64.600 127.400 ;
        RECT 65.400 127.300 66.700 127.600 ;
        RECT 62.200 126.800 63.500 127.200 ;
        RECT 64.200 126.900 65.000 127.200 ;
        RECT 64.600 126.800 65.000 126.900 ;
        RECT 55.800 125.800 56.200 125.900 ;
        RECT 60.600 125.800 62.500 126.100 ;
        RECT 56.600 125.500 59.400 125.600 ;
        RECT 56.500 125.400 59.400 125.500 ;
        RECT 52.600 124.900 53.800 125.200 ;
        RECT 54.500 125.300 59.400 125.400 ;
        RECT 54.500 125.100 56.900 125.300 ;
        RECT 52.600 124.400 52.900 124.900 ;
        RECT 52.200 124.000 52.900 124.400 ;
        RECT 53.700 124.500 54.100 124.600 ;
        RECT 54.500 124.500 54.800 125.100 ;
        RECT 53.700 124.200 54.800 124.500 ;
        RECT 55.100 124.500 57.800 124.800 ;
        RECT 55.100 124.400 55.500 124.500 ;
        RECT 57.400 124.400 57.800 124.500 ;
        RECT 54.300 123.700 54.700 123.800 ;
        RECT 55.700 123.700 56.100 123.800 ;
        RECT 52.600 123.100 53.000 123.500 ;
        RECT 54.300 123.400 56.100 123.700 ;
        RECT 54.700 123.100 55.000 123.400 ;
        RECT 57.400 123.100 57.800 123.500 ;
        RECT 52.300 121.100 52.900 123.100 ;
        RECT 54.600 121.100 55.000 123.100 ;
        RECT 56.800 122.800 57.800 123.100 ;
        RECT 56.800 121.100 57.200 122.800 ;
        RECT 59.000 121.100 59.400 125.300 ;
        RECT 60.600 121.100 61.000 125.800 ;
        RECT 62.200 125.200 62.500 125.800 ;
        RECT 61.400 124.400 61.800 125.200 ;
        RECT 62.200 125.100 62.600 125.200 ;
        RECT 63.200 125.100 63.500 126.800 ;
        RECT 63.800 125.800 64.200 126.600 ;
        RECT 65.500 126.200 65.900 126.600 ;
        RECT 65.400 125.800 65.900 126.200 ;
        RECT 66.400 126.500 66.700 127.300 ;
        RECT 67.200 127.200 67.500 127.900 ;
        RECT 69.400 127.600 69.800 129.900 ;
        RECT 71.000 127.600 71.400 129.900 ;
        RECT 72.600 127.600 73.000 129.900 ;
        RECT 74.200 127.600 74.600 129.900 ;
        RECT 77.700 128.200 78.100 129.500 ;
        RECT 79.800 128.500 80.200 129.500 ;
        RECT 77.700 128.000 78.600 128.200 ;
        RECT 77.300 127.800 78.600 128.000 ;
        RECT 77.300 127.700 78.100 127.800 ;
        RECT 69.400 127.200 70.300 127.600 ;
        RECT 71.000 127.200 72.100 127.600 ;
        RECT 72.600 127.200 73.700 127.600 ;
        RECT 74.200 127.200 75.400 127.600 ;
        RECT 77.300 127.500 77.700 127.700 ;
        RECT 77.300 127.200 77.600 127.500 ;
        RECT 79.900 127.400 80.200 128.500 ;
        RECT 82.100 127.900 82.900 129.900 ;
        RECT 84.900 128.200 85.300 129.900 ;
        RECT 67.000 127.100 67.500 127.200 ;
        RECT 67.800 127.100 68.200 127.200 ;
        RECT 67.000 126.800 68.200 127.100 ;
        RECT 68.600 126.900 69.000 127.200 ;
        RECT 69.900 126.900 70.300 127.200 ;
        RECT 71.700 126.900 72.100 127.200 ;
        RECT 73.300 126.900 73.700 127.200 ;
        RECT 66.400 126.100 66.900 126.500 ;
        RECT 66.400 125.100 66.700 126.100 ;
        RECT 67.200 125.100 67.500 126.800 ;
        RECT 68.600 126.500 69.500 126.900 ;
        RECT 69.900 126.500 71.200 126.900 ;
        RECT 71.700 126.500 72.900 126.900 ;
        RECT 73.300 126.500 74.600 126.900 ;
        RECT 69.900 125.800 70.300 126.500 ;
        RECT 71.700 125.800 72.100 126.500 ;
        RECT 73.300 125.800 73.700 126.500 ;
        RECT 75.000 125.800 75.400 127.200 ;
        RECT 76.600 126.800 77.600 127.200 ;
        RECT 78.100 127.100 80.200 127.400 ;
        RECT 78.100 126.900 78.600 127.100 ;
        RECT 62.200 124.800 62.900 125.100 ;
        RECT 63.200 124.800 63.700 125.100 ;
        RECT 62.600 124.200 62.900 124.800 ;
        RECT 62.600 123.800 63.000 124.200 ;
        RECT 63.300 121.100 63.700 124.800 ;
        RECT 65.400 124.800 66.700 125.100 ;
        RECT 65.400 121.100 65.800 124.800 ;
        RECT 67.000 124.600 67.500 125.100 ;
        RECT 69.400 125.400 70.300 125.800 ;
        RECT 71.000 125.400 72.100 125.800 ;
        RECT 72.600 125.400 73.700 125.800 ;
        RECT 74.200 125.400 75.400 125.800 ;
        RECT 76.600 125.400 77.000 126.200 ;
        RECT 67.000 121.100 67.400 124.600 ;
        RECT 69.400 121.100 69.800 125.400 ;
        RECT 71.000 121.100 71.400 125.400 ;
        RECT 72.600 121.100 73.000 125.400 ;
        RECT 74.200 121.100 74.600 125.400 ;
        RECT 77.300 124.900 77.600 126.800 ;
        RECT 77.900 126.500 78.600 126.900 ;
        RECT 78.300 125.500 78.600 126.500 ;
        RECT 79.000 125.800 79.400 126.600 ;
        RECT 79.800 125.800 80.200 126.600 ;
        RECT 81.400 126.400 81.800 127.200 ;
        RECT 82.300 126.200 82.600 127.900 ;
        RECT 84.600 127.800 85.800 128.200 ;
        RECT 84.600 127.200 84.900 127.800 ;
        RECT 83.000 126.800 83.400 127.200 ;
        RECT 84.600 126.800 85.000 127.200 ;
        RECT 83.000 126.600 83.300 126.800 ;
        RECT 82.900 126.200 83.300 126.600 ;
        RECT 80.600 126.100 81.000 126.200 ;
        RECT 80.600 125.800 81.400 126.100 ;
        RECT 82.200 125.800 82.600 126.200 ;
        RECT 81.000 125.600 81.400 125.800 ;
        RECT 82.300 125.700 82.600 125.800 ;
        RECT 78.300 125.200 80.200 125.500 ;
        RECT 82.300 125.400 83.300 125.700 ;
        RECT 83.800 125.400 84.200 126.200 ;
        RECT 77.300 124.600 78.100 124.900 ;
        RECT 77.700 121.100 78.100 124.600 ;
        RECT 79.900 123.500 80.200 125.200 ;
        RECT 83.000 125.200 83.300 125.400 ;
        RECT 79.800 121.500 80.200 123.500 ;
        RECT 80.600 124.800 82.600 125.100 ;
        RECT 80.600 121.100 81.000 124.800 ;
        RECT 82.200 121.400 82.600 124.800 ;
        RECT 83.000 121.700 83.400 125.200 ;
        RECT 83.800 121.400 84.200 125.100 ;
        RECT 84.600 124.400 85.000 125.200 ;
        RECT 82.200 121.100 84.200 121.400 ;
        RECT 85.400 121.100 85.800 127.800 ;
        RECT 87.000 127.600 87.400 129.900 ;
        RECT 88.600 128.200 89.000 129.900 ;
        RECT 88.600 127.900 89.100 128.200 ;
        RECT 92.100 128.000 92.500 129.500 ;
        RECT 94.200 128.500 94.600 129.500 ;
        RECT 86.200 126.800 86.600 127.600 ;
        RECT 87.000 127.300 88.300 127.600 ;
        RECT 87.100 126.200 87.500 126.600 ;
        RECT 87.000 125.800 87.500 126.200 ;
        RECT 88.000 126.500 88.300 127.300 ;
        RECT 88.800 127.200 89.100 127.900 ;
        RECT 91.700 127.700 92.500 128.000 ;
        RECT 91.700 127.500 92.100 127.700 ;
        RECT 91.700 127.200 92.000 127.500 ;
        RECT 94.300 127.400 94.600 128.500 ;
        RECT 88.600 126.800 89.100 127.200 ;
        RECT 89.400 127.100 89.800 127.200 ;
        RECT 91.000 127.100 92.000 127.200 ;
        RECT 89.400 126.800 92.000 127.100 ;
        RECT 92.500 127.100 94.600 127.400 ;
        RECT 95.000 128.500 95.400 129.500 ;
        RECT 95.000 127.400 95.300 128.500 ;
        RECT 97.100 128.000 97.500 129.500 ;
        RECT 102.700 129.200 103.500 129.900 ;
        RECT 102.200 128.800 103.500 129.200 ;
        RECT 97.100 127.700 97.900 128.000 ;
        RECT 102.700 127.900 103.500 128.800 ;
        RECT 107.300 128.000 107.700 129.500 ;
        RECT 109.400 128.500 109.800 129.500 ;
        RECT 97.500 127.500 97.900 127.700 ;
        RECT 95.000 127.100 97.100 127.400 ;
        RECT 92.500 126.900 93.000 127.100 ;
        RECT 88.000 126.100 88.500 126.500 ;
        RECT 88.000 125.100 88.300 126.100 ;
        RECT 88.800 125.100 89.100 126.800 ;
        RECT 90.200 126.100 90.600 126.200 ;
        RECT 91.000 126.100 91.400 126.200 ;
        RECT 90.200 125.800 91.400 126.100 ;
        RECT 91.000 125.400 91.400 125.800 ;
        RECT 87.000 124.800 88.300 125.100 ;
        RECT 87.000 121.100 87.400 124.800 ;
        RECT 88.600 124.600 89.100 125.100 ;
        RECT 91.700 124.900 92.000 126.800 ;
        RECT 92.300 126.500 93.000 126.900 ;
        RECT 96.600 126.900 97.100 127.100 ;
        RECT 97.600 127.200 97.900 127.500 ;
        RECT 97.600 127.100 98.600 127.200 ;
        RECT 100.600 127.100 101.000 127.200 ;
        RECT 92.700 125.500 93.000 126.500 ;
        RECT 93.400 125.800 93.800 126.600 ;
        RECT 94.200 125.800 94.600 126.600 ;
        RECT 95.000 125.800 95.400 126.600 ;
        RECT 95.800 125.800 96.200 126.600 ;
        RECT 96.600 126.500 97.300 126.900 ;
        RECT 97.600 126.800 101.000 127.100 ;
        RECT 102.200 126.800 102.600 127.200 ;
        RECT 96.600 125.500 96.900 126.500 ;
        RECT 92.700 125.200 94.600 125.500 ;
        RECT 91.700 124.600 92.500 124.900 ;
        RECT 88.600 121.100 89.000 124.600 ;
        RECT 92.100 121.100 92.500 124.600 ;
        RECT 94.300 123.500 94.600 125.200 ;
        RECT 94.200 121.500 94.600 123.500 ;
        RECT 95.000 125.200 96.900 125.500 ;
        RECT 95.000 123.500 95.300 125.200 ;
        RECT 97.600 124.900 97.900 126.800 ;
        RECT 102.300 126.600 102.600 126.800 ;
        RECT 102.300 126.200 102.700 126.600 ;
        RECT 103.000 126.200 103.300 127.900 ;
        RECT 106.900 127.700 107.700 128.000 ;
        RECT 106.900 127.500 107.300 127.700 ;
        RECT 106.900 127.200 107.200 127.500 ;
        RECT 109.500 127.400 109.800 128.500 ;
        RECT 112.100 128.000 112.500 129.500 ;
        RECT 114.200 128.500 114.600 129.500 ;
        RECT 103.800 126.400 104.200 127.200 ;
        RECT 106.200 127.100 107.200 127.200 ;
        RECT 104.600 126.800 107.200 127.100 ;
        RECT 107.700 127.100 109.800 127.400 ;
        RECT 111.700 127.700 112.500 128.000 ;
        RECT 111.700 127.500 112.100 127.700 ;
        RECT 111.700 127.200 112.000 127.500 ;
        RECT 114.300 127.400 114.600 128.500 ;
        RECT 115.000 128.000 115.400 129.900 ;
        RECT 116.600 128.000 117.000 129.900 ;
        RECT 115.000 127.900 117.000 128.000 ;
        RECT 117.400 127.900 117.800 129.900 ;
        RECT 118.500 128.200 118.900 129.900 ;
        RECT 118.500 127.900 119.400 128.200 ;
        RECT 115.100 127.700 116.900 127.900 ;
        RECT 110.200 127.100 110.600 127.200 ;
        RECT 111.000 127.100 112.000 127.200 ;
        RECT 107.700 126.900 108.200 127.100 ;
        RECT 104.600 126.200 104.900 126.800 ;
        RECT 98.200 125.400 98.600 126.200 ;
        RECT 101.400 125.400 101.800 126.200 ;
        RECT 103.000 125.800 103.400 126.200 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 104.200 125.800 105.000 126.100 ;
        RECT 105.400 126.100 105.800 126.200 ;
        RECT 106.200 126.100 106.600 126.200 ;
        RECT 105.400 125.800 106.600 126.100 ;
        RECT 103.000 125.700 103.300 125.800 ;
        RECT 102.300 125.400 103.300 125.700 ;
        RECT 104.200 125.600 104.600 125.800 ;
        RECT 106.200 125.400 106.600 125.800 ;
        RECT 102.300 125.100 102.600 125.400 ;
        RECT 97.100 124.600 97.900 124.900 ;
        RECT 95.000 121.500 95.400 123.500 ;
        RECT 97.100 121.100 97.500 124.600 ;
        RECT 101.400 121.400 101.800 125.100 ;
        RECT 102.200 121.700 102.600 125.100 ;
        RECT 103.000 124.800 105.000 125.100 ;
        RECT 103.000 121.400 103.400 124.800 ;
        RECT 101.400 121.100 103.400 121.400 ;
        RECT 104.600 121.100 105.000 124.800 ;
        RECT 106.900 124.900 107.200 126.800 ;
        RECT 107.500 126.500 108.200 126.900 ;
        RECT 110.200 126.800 112.000 127.100 ;
        RECT 112.500 127.100 114.600 127.400 ;
        RECT 115.400 127.200 115.800 127.400 ;
        RECT 117.400 127.200 117.700 127.900 ;
        RECT 112.500 126.900 113.000 127.100 ;
        RECT 107.900 125.500 108.200 126.500 ;
        RECT 108.600 125.800 109.000 126.600 ;
        RECT 109.400 125.800 109.800 126.600 ;
        RECT 107.900 125.200 109.800 125.500 ;
        RECT 111.000 125.400 111.400 126.200 ;
        RECT 106.900 124.600 107.700 124.900 ;
        RECT 107.300 121.100 107.700 124.600 ;
        RECT 109.500 123.500 109.800 125.200 ;
        RECT 111.700 124.900 112.000 126.800 ;
        RECT 112.300 126.500 113.000 126.900 ;
        RECT 115.000 126.900 115.800 127.200 ;
        RECT 116.500 127.100 117.800 127.200 ;
        RECT 118.200 127.100 118.600 127.200 ;
        RECT 115.000 126.800 115.400 126.900 ;
        RECT 116.500 126.800 118.600 127.100 ;
        RECT 112.700 125.500 113.000 126.500 ;
        RECT 113.400 125.800 113.800 126.600 ;
        RECT 114.200 125.800 114.600 126.600 ;
        RECT 115.000 126.100 115.400 126.200 ;
        RECT 115.800 126.100 116.200 126.600 ;
        RECT 115.000 125.800 116.200 126.100 ;
        RECT 112.700 125.200 114.600 125.500 ;
        RECT 111.700 124.600 112.500 124.900 ;
        RECT 109.400 121.500 109.800 123.500 ;
        RECT 112.100 121.100 112.500 124.600 ;
        RECT 114.300 123.500 114.600 125.200 ;
        RECT 116.500 125.100 116.800 126.800 ;
        RECT 119.000 126.100 119.400 127.900 ;
        RECT 119.800 126.800 120.200 127.600 ;
        RECT 120.600 127.500 121.000 129.900 ;
        RECT 122.800 129.200 123.200 129.900 ;
        RECT 122.200 128.900 123.200 129.200 ;
        RECT 125.000 128.900 125.400 129.900 ;
        RECT 127.100 129.200 127.700 129.900 ;
        RECT 127.000 128.900 127.700 129.200 ;
        RECT 122.200 128.500 122.600 128.900 ;
        RECT 125.000 128.600 125.300 128.900 ;
        RECT 123.000 127.800 123.400 128.600 ;
        RECT 123.900 128.300 125.300 128.600 ;
        RECT 127.000 128.500 127.400 128.900 ;
        RECT 123.900 128.200 124.300 128.300 ;
        RECT 121.000 127.100 121.800 127.200 ;
        RECT 123.100 127.100 123.400 127.800 ;
        RECT 127.900 127.700 128.300 127.800 ;
        RECT 129.400 127.700 129.800 129.900 ;
        RECT 127.900 127.400 129.800 127.700 ;
        RECT 125.900 127.100 126.300 127.200 ;
        RECT 121.000 126.800 126.500 127.100 ;
        RECT 122.500 126.700 122.900 126.800 ;
        RECT 117.400 125.800 119.400 126.100 ;
        RECT 121.700 126.200 122.100 126.300 ;
        RECT 121.700 125.900 124.200 126.200 ;
        RECT 123.800 125.800 124.200 125.900 ;
        RECT 117.400 125.200 117.700 125.800 ;
        RECT 117.400 125.100 117.800 125.200 ;
        RECT 114.200 121.500 114.600 123.500 ;
        RECT 116.300 124.800 116.800 125.100 ;
        RECT 117.100 124.800 117.800 125.100 ;
        RECT 116.300 121.100 116.700 124.800 ;
        RECT 117.100 124.200 117.400 124.800 ;
        RECT 118.200 124.400 118.600 125.200 ;
        RECT 117.000 123.800 117.400 124.200 ;
        RECT 119.000 121.100 119.400 125.800 ;
        RECT 120.600 125.500 123.400 125.600 ;
        RECT 120.600 125.400 123.500 125.500 ;
        RECT 120.600 125.300 125.500 125.400 ;
        RECT 120.600 121.100 121.000 125.300 ;
        RECT 123.100 125.100 125.500 125.300 ;
        RECT 122.200 124.500 124.900 124.800 ;
        RECT 122.200 124.400 122.600 124.500 ;
        RECT 124.500 124.400 124.900 124.500 ;
        RECT 125.200 124.500 125.500 125.100 ;
        RECT 126.200 125.200 126.500 126.800 ;
        RECT 127.000 126.400 127.400 126.500 ;
        RECT 127.000 126.100 128.900 126.400 ;
        RECT 128.500 126.000 128.900 126.100 ;
        RECT 127.700 125.700 128.100 125.800 ;
        RECT 129.400 125.700 129.800 127.400 ;
        RECT 127.700 125.400 129.800 125.700 ;
        RECT 126.200 124.900 127.400 125.200 ;
        RECT 125.900 124.500 126.300 124.600 ;
        RECT 125.200 124.200 126.300 124.500 ;
        RECT 127.100 124.400 127.400 124.900 ;
        RECT 127.100 124.000 127.800 124.400 ;
        RECT 123.900 123.700 124.300 123.800 ;
        RECT 125.300 123.700 125.700 123.800 ;
        RECT 122.200 123.100 122.600 123.500 ;
        RECT 123.900 123.400 125.700 123.700 ;
        RECT 125.000 123.100 125.300 123.400 ;
        RECT 127.000 123.100 127.400 123.500 ;
        RECT 122.200 122.800 123.200 123.100 ;
        RECT 122.800 121.100 123.200 122.800 ;
        RECT 125.000 121.100 125.400 123.100 ;
        RECT 127.100 121.100 127.700 123.100 ;
        RECT 129.400 121.100 129.800 125.400 ;
        RECT 130.200 127.700 130.600 129.900 ;
        RECT 132.300 129.200 132.900 129.900 ;
        RECT 132.300 128.900 133.000 129.200 ;
        RECT 134.600 128.900 135.000 129.900 ;
        RECT 136.800 129.200 137.200 129.900 ;
        RECT 136.800 128.900 137.800 129.200 ;
        RECT 132.600 128.500 133.000 128.900 ;
        RECT 134.700 128.600 135.000 128.900 ;
        RECT 134.700 128.300 136.100 128.600 ;
        RECT 135.700 128.200 136.100 128.300 ;
        RECT 136.600 128.200 137.000 128.600 ;
        RECT 137.400 128.500 137.800 128.900 ;
        RECT 131.700 127.700 132.100 127.800 ;
        RECT 130.200 127.400 132.100 127.700 ;
        RECT 130.200 125.700 130.600 127.400 ;
        RECT 133.700 127.100 134.600 127.200 ;
        RECT 136.600 127.100 136.900 128.200 ;
        RECT 139.000 127.500 139.400 129.900 ;
        RECT 141.100 128.200 141.500 129.900 ;
        RECT 140.600 127.900 141.500 128.200 ;
        RECT 142.200 127.900 142.600 129.900 ;
        RECT 143.000 128.000 143.400 129.900 ;
        RECT 144.600 128.000 145.000 129.900 ;
        RECT 143.000 127.900 145.000 128.000 ;
        RECT 145.400 128.000 145.800 129.900 ;
        RECT 147.000 128.000 147.400 129.900 ;
        RECT 145.400 127.900 147.400 128.000 ;
        RECT 147.800 127.900 148.200 129.900 ;
        RECT 138.200 127.100 139.000 127.200 ;
        RECT 133.500 126.800 139.000 127.100 ;
        RECT 139.800 126.800 140.200 127.600 ;
        RECT 132.600 126.400 133.000 126.500 ;
        RECT 131.100 126.100 133.000 126.400 ;
        RECT 131.100 126.000 131.500 126.100 ;
        RECT 131.900 125.700 132.300 125.800 ;
        RECT 130.200 125.400 132.300 125.700 ;
        RECT 130.200 121.100 130.600 125.400 ;
        RECT 133.500 125.200 133.800 126.800 ;
        RECT 137.100 126.700 137.500 126.800 ;
        RECT 136.600 126.200 137.000 126.300 ;
        RECT 137.900 126.200 138.300 126.300 ;
        RECT 135.800 125.900 138.300 126.200 ;
        RECT 140.600 126.100 141.000 127.900 ;
        RECT 142.300 127.200 142.600 127.900 ;
        RECT 143.100 127.700 144.900 127.900 ;
        RECT 145.500 127.700 147.300 127.900 ;
        RECT 144.200 127.200 144.600 127.400 ;
        RECT 145.800 127.200 146.200 127.400 ;
        RECT 147.800 127.200 148.100 127.900 ;
        RECT 150.200 127.700 150.600 129.900 ;
        RECT 152.300 129.200 152.900 129.900 ;
        RECT 152.300 128.900 153.000 129.200 ;
        RECT 154.600 128.900 155.000 129.900 ;
        RECT 156.800 129.200 157.200 129.900 ;
        RECT 156.800 128.900 157.800 129.200 ;
        RECT 152.600 128.500 153.000 128.900 ;
        RECT 154.700 128.600 155.000 128.900 ;
        RECT 154.700 128.300 156.100 128.600 ;
        RECT 155.700 128.200 156.100 128.300 ;
        RECT 156.600 128.200 157.000 128.600 ;
        RECT 157.400 128.500 157.800 128.900 ;
        RECT 151.700 127.700 152.100 127.800 ;
        RECT 150.200 127.400 152.100 127.700 ;
        RECT 142.200 126.800 143.500 127.200 ;
        RECT 144.200 127.100 145.000 127.200 ;
        RECT 145.400 127.100 146.200 127.200 ;
        RECT 144.200 126.900 146.200 127.100 ;
        RECT 144.600 126.800 145.800 126.900 ;
        RECT 146.900 126.800 148.200 127.200 ;
        RECT 135.800 125.800 136.200 125.900 ;
        RECT 140.600 125.800 142.500 126.100 ;
        RECT 136.600 125.500 139.400 125.600 ;
        RECT 136.500 125.400 139.400 125.500 ;
        RECT 132.600 124.900 133.800 125.200 ;
        RECT 134.500 125.300 139.400 125.400 ;
        RECT 134.500 125.100 136.900 125.300 ;
        RECT 132.600 124.400 132.900 124.900 ;
        RECT 132.200 124.000 132.900 124.400 ;
        RECT 133.700 124.500 134.100 124.600 ;
        RECT 134.500 124.500 134.800 125.100 ;
        RECT 133.700 124.200 134.800 124.500 ;
        RECT 135.100 124.500 137.800 124.800 ;
        RECT 135.100 124.400 135.500 124.500 ;
        RECT 137.400 124.400 137.800 124.500 ;
        RECT 134.300 123.700 134.700 123.800 ;
        RECT 135.700 123.700 136.100 123.800 ;
        RECT 132.600 123.100 133.000 123.500 ;
        RECT 134.300 123.400 136.100 123.700 ;
        RECT 134.700 123.100 135.000 123.400 ;
        RECT 137.400 123.100 137.800 123.500 ;
        RECT 132.300 121.100 132.900 123.100 ;
        RECT 134.600 121.100 135.000 123.100 ;
        RECT 136.800 122.800 137.800 123.100 ;
        RECT 136.800 121.100 137.200 122.800 ;
        RECT 139.000 121.100 139.400 125.300 ;
        RECT 140.600 121.100 141.000 125.800 ;
        RECT 142.200 125.200 142.500 125.800 ;
        RECT 141.400 124.400 141.800 125.200 ;
        RECT 142.200 125.100 142.600 125.200 ;
        RECT 143.200 125.100 143.500 126.800 ;
        RECT 143.800 125.800 144.200 126.600 ;
        RECT 146.200 125.800 146.600 126.600 ;
        RECT 146.900 125.100 147.200 126.800 ;
        RECT 150.200 125.700 150.600 127.400 ;
        RECT 153.700 127.100 154.600 127.200 ;
        RECT 156.600 127.100 156.900 128.200 ;
        RECT 159.000 127.500 159.400 129.900 ;
        RECT 161.100 128.200 161.500 129.900 ;
        RECT 160.600 127.900 161.500 128.200 ;
        RECT 162.200 127.900 162.600 129.900 ;
        RECT 163.000 128.000 163.400 129.900 ;
        RECT 164.600 128.000 165.000 129.900 ;
        RECT 163.000 127.900 165.000 128.000 ;
        RECT 165.400 128.500 165.800 129.500 ;
        RECT 158.200 127.100 159.000 127.200 ;
        RECT 153.500 126.800 159.000 127.100 ;
        RECT 159.800 126.800 160.200 127.600 ;
        RECT 152.600 126.400 153.000 126.500 ;
        RECT 151.100 126.100 153.000 126.400 ;
        RECT 151.100 126.000 151.500 126.100 ;
        RECT 151.900 125.700 152.300 125.800 ;
        RECT 150.200 125.400 152.300 125.700 ;
        RECT 147.800 125.100 148.200 125.200 ;
        RECT 142.200 124.800 142.900 125.100 ;
        RECT 143.200 124.800 143.700 125.100 ;
        RECT 142.600 124.200 142.900 124.800 ;
        RECT 142.600 123.800 143.000 124.200 ;
        RECT 143.300 121.100 143.700 124.800 ;
        RECT 146.700 124.800 147.200 125.100 ;
        RECT 147.500 124.800 148.200 125.100 ;
        RECT 146.700 121.100 147.100 124.800 ;
        RECT 147.500 124.200 147.800 124.800 ;
        RECT 147.400 123.800 147.800 124.200 ;
        RECT 150.200 121.100 150.600 125.400 ;
        RECT 153.500 125.200 153.800 126.800 ;
        RECT 157.100 126.700 157.500 126.800 ;
        RECT 156.600 126.200 157.000 126.300 ;
        RECT 157.900 126.200 158.300 126.300 ;
        RECT 155.800 125.900 158.300 126.200 ;
        RECT 160.600 126.100 161.000 127.900 ;
        RECT 162.300 127.200 162.600 127.900 ;
        RECT 163.100 127.700 164.900 127.900 ;
        RECT 165.400 127.400 165.700 128.500 ;
        RECT 167.500 128.000 167.900 129.500 ;
        RECT 170.200 128.000 170.600 129.900 ;
        RECT 171.800 128.000 172.200 129.900 ;
        RECT 167.500 127.700 168.300 128.000 ;
        RECT 170.200 127.900 172.200 128.000 ;
        RECT 172.600 127.900 173.000 129.900 ;
        RECT 173.700 128.200 174.100 129.900 ;
        RECT 173.700 127.900 174.600 128.200 ;
        RECT 170.300 127.700 172.100 127.900 ;
        RECT 167.900 127.500 168.300 127.700 ;
        RECT 164.200 127.200 164.600 127.400 ;
        RECT 161.400 127.100 161.800 127.200 ;
        RECT 162.200 127.100 163.500 127.200 ;
        RECT 161.400 126.800 163.500 127.100 ;
        RECT 164.200 126.900 165.000 127.200 ;
        RECT 165.400 127.100 167.500 127.400 ;
        RECT 164.600 126.800 165.000 126.900 ;
        RECT 167.000 126.900 167.500 127.100 ;
        RECT 168.000 127.200 168.300 127.500 ;
        RECT 170.600 127.200 171.000 127.400 ;
        RECT 172.600 127.200 172.900 127.900 ;
        RECT 155.800 125.800 156.200 125.900 ;
        RECT 160.600 125.800 162.500 126.100 ;
        RECT 156.600 125.500 159.400 125.600 ;
        RECT 156.500 125.400 159.400 125.500 ;
        RECT 152.600 124.900 153.800 125.200 ;
        RECT 154.500 125.300 159.400 125.400 ;
        RECT 154.500 125.100 156.900 125.300 ;
        RECT 152.600 124.400 152.900 124.900 ;
        RECT 152.200 124.000 152.900 124.400 ;
        RECT 153.700 124.500 154.100 124.600 ;
        RECT 154.500 124.500 154.800 125.100 ;
        RECT 153.700 124.200 154.800 124.500 ;
        RECT 155.100 124.500 157.800 124.800 ;
        RECT 155.100 124.400 155.500 124.500 ;
        RECT 157.400 124.400 157.800 124.500 ;
        RECT 154.300 123.700 154.700 123.800 ;
        RECT 155.700 123.700 156.100 123.800 ;
        RECT 152.600 123.100 153.000 123.500 ;
        RECT 154.300 123.400 156.100 123.700 ;
        RECT 154.700 123.100 155.000 123.400 ;
        RECT 157.400 123.100 157.800 123.500 ;
        RECT 152.300 121.100 152.900 123.100 ;
        RECT 154.600 121.100 155.000 123.100 ;
        RECT 156.800 122.800 157.800 123.100 ;
        RECT 156.800 121.100 157.200 122.800 ;
        RECT 159.000 121.100 159.400 125.300 ;
        RECT 160.600 121.100 161.000 125.800 ;
        RECT 162.200 125.200 162.500 125.800 ;
        RECT 161.400 124.400 161.800 125.200 ;
        RECT 162.200 125.100 162.600 125.200 ;
        RECT 163.200 125.100 163.500 126.800 ;
        RECT 163.800 125.800 164.200 126.600 ;
        RECT 165.400 125.800 165.800 126.600 ;
        RECT 166.200 125.800 166.600 126.600 ;
        RECT 167.000 126.500 167.700 126.900 ;
        RECT 168.000 126.800 169.000 127.200 ;
        RECT 170.200 126.900 171.000 127.200 ;
        RECT 170.200 126.800 170.600 126.900 ;
        RECT 171.700 126.800 173.000 127.200 ;
        RECT 167.000 125.500 167.300 126.500 ;
        RECT 165.400 125.200 167.300 125.500 ;
        RECT 162.200 124.800 162.900 125.100 ;
        RECT 163.200 124.800 163.700 125.100 ;
        RECT 162.600 124.200 162.900 124.800 ;
        RECT 162.600 123.800 163.000 124.200 ;
        RECT 163.300 121.100 163.700 124.800 ;
        RECT 165.400 123.500 165.700 125.200 ;
        RECT 168.000 124.900 168.300 126.800 ;
        RECT 168.600 125.400 169.000 126.200 ;
        RECT 171.000 125.800 171.400 126.600 ;
        RECT 171.700 125.100 172.000 126.800 ;
        RECT 174.200 126.100 174.600 127.900 ;
        RECT 175.000 126.800 175.400 127.600 ;
        RECT 175.800 127.500 176.200 129.900 ;
        RECT 178.000 129.200 178.400 129.900 ;
        RECT 177.400 128.900 178.400 129.200 ;
        RECT 180.200 128.900 180.600 129.900 ;
        RECT 182.300 129.200 182.900 129.900 ;
        RECT 182.200 128.900 182.900 129.200 ;
        RECT 177.400 128.500 177.800 128.900 ;
        RECT 180.200 128.600 180.500 128.900 ;
        RECT 178.200 127.800 178.600 128.600 ;
        RECT 179.100 128.300 180.500 128.600 ;
        RECT 182.200 128.500 182.600 128.900 ;
        RECT 179.100 128.200 179.500 128.300 ;
        RECT 176.200 127.100 177.000 127.200 ;
        RECT 178.300 127.100 178.600 127.800 ;
        RECT 183.100 127.700 183.500 127.800 ;
        RECT 184.600 127.700 185.000 129.900 ;
        RECT 183.100 127.400 185.000 127.700 ;
        RECT 181.100 127.100 181.500 127.200 ;
        RECT 176.200 126.800 181.700 127.100 ;
        RECT 177.700 126.700 178.100 126.800 ;
        RECT 172.600 125.800 174.600 126.100 ;
        RECT 176.900 126.200 177.300 126.300 ;
        RECT 178.200 126.200 178.600 126.300 ;
        RECT 181.400 126.200 181.700 126.800 ;
        RECT 182.200 126.400 182.600 126.500 ;
        RECT 176.900 125.900 179.400 126.200 ;
        RECT 179.000 125.800 179.400 125.900 ;
        RECT 181.400 125.800 181.800 126.200 ;
        RECT 182.200 126.100 184.100 126.400 ;
        RECT 183.700 126.000 184.100 126.100 ;
        RECT 172.600 125.200 172.900 125.800 ;
        RECT 172.600 125.100 173.000 125.200 ;
        RECT 167.500 124.600 168.300 124.900 ;
        RECT 171.500 124.800 172.000 125.100 ;
        RECT 172.300 124.800 173.000 125.100 ;
        RECT 165.400 121.500 165.800 123.500 ;
        RECT 167.500 122.200 167.900 124.600 ;
        RECT 167.000 121.800 167.900 122.200 ;
        RECT 167.500 121.100 167.900 121.800 ;
        RECT 171.500 121.100 171.900 124.800 ;
        RECT 172.300 124.200 172.600 124.800 ;
        RECT 173.400 124.400 173.800 125.200 ;
        RECT 172.200 123.800 172.600 124.200 ;
        RECT 174.200 121.100 174.600 125.800 ;
        RECT 175.800 125.500 178.600 125.600 ;
        RECT 175.800 125.400 178.700 125.500 ;
        RECT 175.800 125.300 180.700 125.400 ;
        RECT 175.800 121.100 176.200 125.300 ;
        RECT 178.300 125.100 180.700 125.300 ;
        RECT 177.400 124.500 180.100 124.800 ;
        RECT 177.400 124.400 177.800 124.500 ;
        RECT 179.700 124.400 180.100 124.500 ;
        RECT 180.400 124.500 180.700 125.100 ;
        RECT 181.400 125.200 181.700 125.800 ;
        RECT 182.900 125.700 183.300 125.800 ;
        RECT 184.600 125.700 185.000 127.400 ;
        RECT 185.400 128.500 185.800 129.500 ;
        RECT 185.400 127.400 185.700 128.500 ;
        RECT 187.500 128.000 187.900 129.500 ;
        RECT 191.500 129.200 192.300 129.900 ;
        RECT 191.000 128.800 192.300 129.200 ;
        RECT 187.500 127.700 188.300 128.000 ;
        RECT 191.500 127.900 192.300 128.800 ;
        RECT 196.100 128.000 196.500 129.500 ;
        RECT 198.200 128.500 198.600 129.500 ;
        RECT 187.900 127.500 188.300 127.700 ;
        RECT 185.400 127.100 187.500 127.400 ;
        RECT 187.000 126.900 187.500 127.100 ;
        RECT 188.000 127.200 188.300 127.500 ;
        RECT 188.000 127.100 189.000 127.200 ;
        RECT 185.400 125.800 185.800 126.600 ;
        RECT 186.200 125.800 186.600 126.600 ;
        RECT 187.000 126.500 187.700 126.900 ;
        RECT 188.000 126.800 189.700 127.100 ;
        RECT 191.000 126.800 191.400 127.200 ;
        RECT 182.900 125.400 185.000 125.700 ;
        RECT 187.000 125.500 187.300 126.500 ;
        RECT 181.400 124.900 182.600 125.200 ;
        RECT 181.100 124.500 181.500 124.600 ;
        RECT 180.400 124.200 181.500 124.500 ;
        RECT 182.300 124.400 182.600 124.900 ;
        RECT 182.300 124.000 183.000 124.400 ;
        RECT 179.100 123.700 179.500 123.800 ;
        RECT 180.500 123.700 180.900 123.800 ;
        RECT 177.400 123.100 177.800 123.500 ;
        RECT 179.100 123.400 180.900 123.700 ;
        RECT 180.200 123.100 180.500 123.400 ;
        RECT 182.200 123.100 182.600 123.500 ;
        RECT 177.400 122.800 178.400 123.100 ;
        RECT 178.000 121.100 178.400 122.800 ;
        RECT 180.200 121.100 180.600 123.100 ;
        RECT 182.300 121.100 182.900 123.100 ;
        RECT 184.600 121.100 185.000 125.400 ;
        RECT 185.400 125.200 187.300 125.500 ;
        RECT 185.400 123.500 185.700 125.200 ;
        RECT 188.000 124.900 188.300 126.800 ;
        RECT 189.400 126.200 189.700 126.800 ;
        RECT 191.100 126.600 191.400 126.800 ;
        RECT 191.100 126.200 191.500 126.600 ;
        RECT 191.800 126.200 192.100 127.900 ;
        RECT 195.700 127.700 196.500 128.000 ;
        RECT 195.700 127.500 196.100 127.700 ;
        RECT 195.700 127.200 196.000 127.500 ;
        RECT 198.300 127.400 198.600 128.500 ;
        RECT 192.600 126.400 193.000 127.200 ;
        RECT 195.000 127.100 196.000 127.200 ;
        RECT 193.400 126.800 196.000 127.100 ;
        RECT 196.500 127.100 198.600 127.400 ;
        RECT 200.600 127.700 201.000 129.900 ;
        RECT 202.700 129.200 203.300 129.900 ;
        RECT 202.700 128.900 203.400 129.200 ;
        RECT 205.000 128.900 205.400 129.900 ;
        RECT 207.200 129.200 207.600 129.900 ;
        RECT 207.200 128.900 208.200 129.200 ;
        RECT 203.000 128.500 203.400 128.900 ;
        RECT 205.100 128.600 205.400 128.900 ;
        RECT 205.100 128.300 206.500 128.600 ;
        RECT 206.100 128.200 206.500 128.300 ;
        RECT 207.000 127.800 207.400 128.600 ;
        RECT 207.800 128.500 208.200 128.900 ;
        RECT 202.100 127.700 202.500 127.800 ;
        RECT 200.600 127.400 202.500 127.700 ;
        RECT 196.500 126.900 197.000 127.100 ;
        RECT 193.400 126.200 193.700 126.800 ;
        RECT 188.600 125.400 189.000 126.200 ;
        RECT 189.400 125.800 189.800 126.200 ;
        RECT 190.200 125.400 190.600 126.200 ;
        RECT 191.800 125.800 192.200 126.200 ;
        RECT 193.400 126.100 193.800 126.200 ;
        RECT 193.000 125.800 193.800 126.100 ;
        RECT 191.800 125.700 192.100 125.800 ;
        RECT 191.100 125.400 192.100 125.700 ;
        RECT 193.000 125.600 193.400 125.800 ;
        RECT 195.000 125.400 195.400 126.200 ;
        RECT 191.100 125.100 191.400 125.400 ;
        RECT 187.500 124.600 188.300 124.900 ;
        RECT 185.400 121.500 185.800 123.500 ;
        RECT 187.500 121.100 187.900 124.600 ;
        RECT 190.200 121.400 190.600 125.100 ;
        RECT 191.000 121.700 191.400 125.100 ;
        RECT 191.800 124.800 193.800 125.100 ;
        RECT 191.800 121.400 192.200 124.800 ;
        RECT 190.200 121.100 192.200 121.400 ;
        RECT 193.400 121.100 193.800 124.800 ;
        RECT 195.700 124.900 196.000 126.800 ;
        RECT 196.300 126.500 197.000 126.900 ;
        RECT 196.700 125.500 197.000 126.500 ;
        RECT 197.400 125.800 197.800 126.600 ;
        RECT 198.200 125.800 198.600 126.600 ;
        RECT 200.600 125.700 201.000 127.400 ;
        RECT 204.100 127.100 204.500 127.200 ;
        RECT 207.000 127.100 207.300 127.800 ;
        RECT 209.400 127.500 209.800 129.900 ;
        RECT 211.500 128.200 211.900 129.900 ;
        RECT 211.000 127.900 211.900 128.200 ;
        RECT 212.600 127.900 213.000 129.900 ;
        RECT 213.400 128.000 213.800 129.900 ;
        RECT 215.000 128.000 215.400 129.900 ;
        RECT 213.400 127.900 215.400 128.000 ;
        RECT 215.800 128.500 216.200 129.500 ;
        RECT 208.600 127.100 209.400 127.200 ;
        RECT 203.900 126.800 209.400 127.100 ;
        RECT 210.200 126.800 210.600 127.600 ;
        RECT 203.000 126.400 203.400 126.500 ;
        RECT 201.500 126.100 203.400 126.400 ;
        RECT 201.500 126.000 201.900 126.100 ;
        RECT 202.300 125.700 202.700 125.800 ;
        RECT 196.700 125.200 198.600 125.500 ;
        RECT 195.700 124.600 196.500 124.900 ;
        RECT 196.100 121.100 196.500 124.600 ;
        RECT 198.300 123.500 198.600 125.200 ;
        RECT 198.200 121.500 198.600 123.500 ;
        RECT 200.600 125.400 202.700 125.700 ;
        RECT 200.600 121.100 201.000 125.400 ;
        RECT 203.900 125.200 204.200 126.800 ;
        RECT 207.500 126.700 207.900 126.800 ;
        RECT 207.000 126.200 207.400 126.300 ;
        RECT 208.300 126.200 208.700 126.300 ;
        RECT 206.200 125.900 208.700 126.200 ;
        RECT 211.000 126.100 211.400 127.900 ;
        RECT 212.700 127.200 213.000 127.900 ;
        RECT 213.500 127.700 215.300 127.900 ;
        RECT 215.800 127.400 216.100 128.500 ;
        RECT 217.900 128.200 218.300 129.500 ;
        RECT 217.400 128.000 218.300 128.200 ;
        RECT 220.900 128.200 221.300 129.900 ;
        RECT 217.400 127.800 218.700 128.000 ;
        RECT 220.900 127.900 221.800 128.200 ;
        RECT 223.000 127.900 223.400 129.900 ;
        RECT 223.800 128.000 224.200 129.900 ;
        RECT 225.400 128.000 225.800 129.900 ;
        RECT 223.800 127.900 225.800 128.000 ;
        RECT 217.900 127.700 218.700 127.800 ;
        RECT 218.300 127.500 218.700 127.700 ;
        RECT 214.600 127.200 215.000 127.400 ;
        RECT 211.800 127.100 212.200 127.200 ;
        RECT 212.600 127.100 213.900 127.200 ;
        RECT 211.800 126.800 213.900 127.100 ;
        RECT 214.600 126.900 215.400 127.200 ;
        RECT 215.800 127.100 217.900 127.400 ;
        RECT 215.000 126.800 215.400 126.900 ;
        RECT 217.400 126.900 217.900 127.100 ;
        RECT 218.400 127.200 218.700 127.500 ;
        RECT 206.200 125.800 206.600 125.900 ;
        RECT 211.000 125.800 212.900 126.100 ;
        RECT 207.000 125.500 209.800 125.600 ;
        RECT 206.900 125.400 209.800 125.500 ;
        RECT 203.000 124.900 204.200 125.200 ;
        RECT 204.900 125.300 209.800 125.400 ;
        RECT 204.900 125.100 207.300 125.300 ;
        RECT 203.000 124.400 203.300 124.900 ;
        RECT 202.600 124.200 203.300 124.400 ;
        RECT 204.100 124.500 204.500 124.600 ;
        RECT 204.900 124.500 205.200 125.100 ;
        RECT 204.100 124.200 205.200 124.500 ;
        RECT 205.500 124.500 208.200 124.800 ;
        RECT 205.500 124.400 205.900 124.500 ;
        RECT 207.800 124.400 208.200 124.500 ;
        RECT 202.200 124.000 203.300 124.200 ;
        RECT 202.200 123.800 202.900 124.000 ;
        RECT 204.700 123.700 205.100 123.800 ;
        RECT 206.100 123.700 206.500 123.800 ;
        RECT 203.000 123.100 203.400 123.500 ;
        RECT 204.700 123.400 206.500 123.700 ;
        RECT 205.100 123.100 205.400 123.400 ;
        RECT 207.800 123.100 208.200 123.500 ;
        RECT 202.700 121.100 203.300 123.100 ;
        RECT 205.000 121.100 205.400 123.100 ;
        RECT 207.200 122.800 208.200 123.100 ;
        RECT 207.200 121.100 207.600 122.800 ;
        RECT 209.400 121.100 209.800 125.300 ;
        RECT 211.000 121.100 211.400 125.800 ;
        RECT 212.600 125.200 212.900 125.800 ;
        RECT 211.800 124.400 212.200 125.200 ;
        RECT 212.600 125.100 213.000 125.200 ;
        RECT 213.600 125.100 213.900 126.800 ;
        RECT 214.200 125.800 214.600 126.600 ;
        RECT 215.800 125.800 216.200 126.600 ;
        RECT 216.600 125.800 217.000 126.600 ;
        RECT 217.400 126.500 218.100 126.900 ;
        RECT 218.400 126.800 219.400 127.200 ;
        RECT 217.400 125.500 217.700 126.500 ;
        RECT 215.800 125.200 217.700 125.500 ;
        RECT 212.600 124.800 213.300 125.100 ;
        RECT 213.600 124.800 214.100 125.100 ;
        RECT 213.000 124.200 213.300 124.800 ;
        RECT 213.000 123.800 213.400 124.200 ;
        RECT 213.700 121.100 214.100 124.800 ;
        RECT 215.800 123.500 216.100 125.200 ;
        RECT 218.400 124.900 218.700 126.800 ;
        RECT 219.000 125.400 219.400 126.200 ;
        RECT 217.900 124.600 218.700 124.900 ;
        RECT 215.800 121.500 216.200 123.500 ;
        RECT 217.900 121.100 218.300 124.600 ;
        RECT 220.600 124.400 221.000 125.200 ;
        RECT 221.400 125.100 221.800 127.900 ;
        RECT 222.200 126.800 222.600 127.600 ;
        RECT 223.100 127.200 223.400 127.900 ;
        RECT 223.900 127.700 225.700 127.900 ;
        RECT 226.200 127.700 226.600 129.900 ;
        RECT 228.300 129.200 228.900 129.900 ;
        RECT 228.300 128.900 229.000 129.200 ;
        RECT 230.600 128.900 231.000 129.900 ;
        RECT 232.800 129.200 233.200 129.900 ;
        RECT 232.800 128.900 233.800 129.200 ;
        RECT 228.600 128.500 229.000 128.900 ;
        RECT 230.700 128.600 231.000 128.900 ;
        RECT 230.700 128.300 232.100 128.600 ;
        RECT 231.700 128.200 232.100 128.300 ;
        RECT 232.600 128.200 233.000 128.600 ;
        RECT 233.400 128.500 233.800 128.900 ;
        RECT 227.700 127.700 228.100 127.800 ;
        RECT 226.200 127.400 228.100 127.700 ;
        RECT 225.000 127.200 225.400 127.400 ;
        RECT 223.000 126.800 224.300 127.200 ;
        RECT 225.000 126.900 225.800 127.200 ;
        RECT 225.400 126.800 225.800 126.900 ;
        RECT 224.000 125.200 224.300 126.800 ;
        RECT 224.600 125.800 225.000 126.600 ;
        RECT 226.200 125.700 226.600 127.400 ;
        RECT 229.700 127.100 230.100 127.200 ;
        RECT 232.600 127.100 232.900 128.200 ;
        RECT 235.000 127.500 235.400 129.900 ;
        RECT 237.100 129.200 237.500 129.900 ;
        RECT 236.600 128.800 237.500 129.200 ;
        RECT 237.100 128.200 237.500 128.800 ;
        RECT 236.600 127.900 237.500 128.200 ;
        RECT 239.800 127.900 240.200 129.900 ;
        RECT 240.500 128.200 240.900 128.600 ;
        RECT 234.200 127.100 235.000 127.200 ;
        RECT 229.500 126.800 235.000 127.100 ;
        RECT 235.800 126.800 236.200 127.600 ;
        RECT 228.600 126.400 229.000 126.500 ;
        RECT 227.100 126.100 229.000 126.400 ;
        RECT 227.100 126.000 227.500 126.100 ;
        RECT 227.900 125.700 228.300 125.800 ;
        RECT 226.200 125.400 228.300 125.700 ;
        RECT 223.000 125.100 223.400 125.200 ;
        RECT 221.400 124.800 223.700 125.100 ;
        RECT 224.000 124.800 225.000 125.200 ;
        RECT 221.400 121.100 221.800 124.800 ;
        RECT 223.400 124.200 223.700 124.800 ;
        RECT 223.400 123.800 223.800 124.200 ;
        RECT 224.100 121.100 224.500 124.800 ;
        RECT 226.200 121.100 226.600 125.400 ;
        RECT 229.500 125.200 229.800 126.800 ;
        RECT 233.100 126.700 233.500 126.800 ;
        RECT 233.900 126.200 234.300 126.300 ;
        RECT 231.800 125.900 234.300 126.200 ;
        RECT 231.800 125.800 232.200 125.900 ;
        RECT 232.600 125.500 235.400 125.600 ;
        RECT 232.500 125.400 235.400 125.500 ;
        RECT 228.600 124.900 229.800 125.200 ;
        RECT 230.500 125.300 235.400 125.400 ;
        RECT 230.500 125.100 232.900 125.300 ;
        RECT 228.600 124.400 228.900 124.900 ;
        RECT 228.200 124.000 228.900 124.400 ;
        RECT 229.700 124.500 230.100 124.600 ;
        RECT 230.500 124.500 230.800 125.100 ;
        RECT 229.700 124.200 230.800 124.500 ;
        RECT 231.100 124.500 233.800 124.800 ;
        RECT 231.100 124.400 231.500 124.500 ;
        RECT 233.400 124.400 233.800 124.500 ;
        RECT 230.300 123.700 230.700 123.800 ;
        RECT 231.700 123.700 232.100 123.800 ;
        RECT 228.600 123.100 229.000 123.500 ;
        RECT 230.300 123.400 232.100 123.700 ;
        RECT 230.700 123.100 231.000 123.400 ;
        RECT 233.400 123.100 233.800 123.500 ;
        RECT 228.300 121.100 228.900 123.100 ;
        RECT 230.600 121.100 231.000 123.100 ;
        RECT 232.800 122.800 233.800 123.100 ;
        RECT 232.800 121.100 233.200 122.800 ;
        RECT 235.000 121.100 235.400 125.300 ;
        RECT 236.600 121.100 237.000 127.900 ;
        RECT 239.000 126.400 239.400 127.200 ;
        RECT 238.200 126.100 238.600 126.200 ;
        RECT 239.800 126.100 240.100 127.900 ;
        RECT 240.600 127.800 241.000 128.200 ;
        RECT 241.400 127.700 241.800 129.900 ;
        RECT 243.500 129.200 244.100 129.900 ;
        RECT 243.500 128.900 244.200 129.200 ;
        RECT 245.800 128.900 246.200 129.900 ;
        RECT 248.000 129.200 248.400 129.900 ;
        RECT 248.000 128.900 249.000 129.200 ;
        RECT 243.800 128.500 244.200 128.900 ;
        RECT 245.900 128.600 246.200 128.900 ;
        RECT 245.900 128.300 247.300 128.600 ;
        RECT 246.900 128.200 247.300 128.300 ;
        RECT 247.800 128.200 248.200 128.600 ;
        RECT 248.600 128.500 249.000 128.900 ;
        RECT 242.900 127.700 243.300 127.800 ;
        RECT 241.400 127.400 243.300 127.700 ;
        RECT 240.600 126.800 241.000 127.200 ;
        RECT 240.600 126.200 240.900 126.800 ;
        RECT 240.600 126.100 241.000 126.200 ;
        RECT 238.200 125.800 239.000 126.100 ;
        RECT 239.800 125.800 241.000 126.100 ;
        RECT 238.600 125.600 239.000 125.800 ;
        RECT 237.400 124.400 237.800 125.200 ;
        RECT 240.600 125.100 240.900 125.800 ;
        RECT 241.400 125.700 241.800 127.400 ;
        RECT 244.900 127.100 245.800 127.200 ;
        RECT 247.800 127.100 248.100 128.200 ;
        RECT 250.200 127.500 250.600 129.900 ;
        RECT 249.400 127.100 250.200 127.200 ;
        RECT 244.700 126.800 250.200 127.100 ;
        RECT 243.800 126.400 244.200 126.500 ;
        RECT 242.300 126.100 244.200 126.400 ;
        RECT 242.300 126.000 242.700 126.100 ;
        RECT 243.100 125.700 243.500 125.800 ;
        RECT 241.400 125.400 243.500 125.700 ;
        RECT 238.200 124.800 240.200 125.100 ;
        RECT 238.200 121.100 238.600 124.800 ;
        RECT 239.800 121.100 240.200 124.800 ;
        RECT 240.600 121.100 241.000 125.100 ;
        RECT 241.400 121.100 241.800 125.400 ;
        RECT 244.700 125.200 245.000 126.800 ;
        RECT 248.300 126.700 248.700 126.800 ;
        RECT 249.100 126.200 249.500 126.300 ;
        RECT 245.400 126.100 245.800 126.200 ;
        RECT 247.000 126.100 249.500 126.200 ;
        RECT 245.400 125.900 249.500 126.100 ;
        RECT 245.400 125.800 247.400 125.900 ;
        RECT 247.800 125.500 250.600 125.600 ;
        RECT 247.700 125.400 250.600 125.500 ;
        RECT 243.800 124.900 245.000 125.200 ;
        RECT 245.700 125.300 250.600 125.400 ;
        RECT 245.700 125.100 248.100 125.300 ;
        RECT 243.800 124.400 244.100 124.900 ;
        RECT 243.400 124.000 244.100 124.400 ;
        RECT 244.900 124.500 245.300 124.600 ;
        RECT 245.700 124.500 246.000 125.100 ;
        RECT 244.900 124.200 246.000 124.500 ;
        RECT 246.300 124.500 249.000 124.800 ;
        RECT 246.300 124.400 246.700 124.500 ;
        RECT 248.600 124.400 249.000 124.500 ;
        RECT 245.500 123.700 245.900 123.800 ;
        RECT 246.900 123.700 247.300 123.800 ;
        RECT 243.800 123.100 244.200 123.500 ;
        RECT 245.500 123.400 247.300 123.700 ;
        RECT 245.900 123.100 246.200 123.400 ;
        RECT 248.600 123.100 249.000 123.500 ;
        RECT 243.500 121.100 244.100 123.100 ;
        RECT 245.800 121.100 246.200 123.100 ;
        RECT 248.000 122.800 249.000 123.100 ;
        RECT 248.000 121.100 248.400 122.800 ;
        RECT 250.200 121.100 250.600 125.300 ;
        RECT 1.400 115.600 1.800 119.900 ;
        RECT 3.000 115.600 3.400 119.900 ;
        RECT 4.600 115.600 5.000 119.900 ;
        RECT 6.200 115.600 6.600 119.900 ;
        RECT 0.600 115.200 1.800 115.600 ;
        RECT 2.300 115.200 3.400 115.600 ;
        RECT 3.900 115.200 5.000 115.600 ;
        RECT 5.700 115.200 6.600 115.600 ;
        RECT 0.600 113.800 1.000 115.200 ;
        RECT 2.300 114.500 2.700 115.200 ;
        RECT 3.900 114.500 4.300 115.200 ;
        RECT 5.700 114.500 6.100 115.200 ;
        RECT 8.600 115.100 9.000 119.900 ;
        RECT 10.600 116.800 11.000 117.200 ;
        RECT 9.400 115.800 9.800 116.600 ;
        RECT 10.600 116.200 10.900 116.800 ;
        RECT 11.300 116.200 11.700 119.900 ;
        RECT 10.200 115.900 10.900 116.200 ;
        RECT 11.200 115.900 11.700 116.200 ;
        RECT 10.200 115.800 10.600 115.900 ;
        RECT 10.200 115.100 10.500 115.800 ;
        RECT 11.200 115.200 11.500 115.900 ;
        RECT 13.400 115.700 13.800 119.900 ;
        RECT 15.600 118.200 16.000 119.900 ;
        RECT 15.000 117.900 16.000 118.200 ;
        RECT 17.800 117.900 18.200 119.900 ;
        RECT 19.900 117.900 20.500 119.900 ;
        RECT 15.000 117.500 15.400 117.900 ;
        RECT 17.800 117.600 18.100 117.900 ;
        RECT 16.700 117.300 18.500 117.600 ;
        RECT 19.800 117.500 20.200 117.900 ;
        RECT 16.700 117.200 17.100 117.300 ;
        RECT 18.100 117.200 18.500 117.300 ;
        RECT 15.000 116.500 15.400 116.600 ;
        RECT 17.300 116.500 17.700 116.600 ;
        RECT 15.000 116.200 17.700 116.500 ;
        RECT 18.000 116.500 19.100 116.800 ;
        RECT 18.000 115.900 18.300 116.500 ;
        RECT 18.700 116.400 19.100 116.500 ;
        RECT 19.900 116.600 20.600 117.000 ;
        RECT 19.900 116.100 20.200 116.600 ;
        RECT 15.900 115.700 18.300 115.900 ;
        RECT 13.400 115.600 18.300 115.700 ;
        RECT 19.000 115.800 20.200 116.100 ;
        RECT 13.400 115.500 16.300 115.600 ;
        RECT 13.400 115.400 16.200 115.500 ;
        RECT 8.600 114.800 10.500 115.100 ;
        RECT 11.000 114.800 11.500 115.200 ;
        RECT 1.400 114.100 2.700 114.500 ;
        RECT 3.100 114.100 4.300 114.500 ;
        RECT 4.800 114.100 6.100 114.500 ;
        RECT 6.500 114.100 7.400 114.500 ;
        RECT 2.300 113.800 2.700 114.100 ;
        RECT 3.900 113.800 4.300 114.100 ;
        RECT 5.700 113.800 6.100 114.100 ;
        RECT 7.000 113.800 7.400 114.100 ;
        RECT 0.600 113.400 1.800 113.800 ;
        RECT 2.300 113.400 3.400 113.800 ;
        RECT 3.900 113.400 5.000 113.800 ;
        RECT 5.700 113.400 6.600 113.800 ;
        RECT 7.800 113.400 8.200 114.200 ;
        RECT 1.400 111.100 1.800 113.400 ;
        RECT 3.000 111.100 3.400 113.400 ;
        RECT 4.600 111.100 5.000 113.400 ;
        RECT 6.200 111.100 6.600 113.400 ;
        RECT 8.600 113.100 9.000 114.800 ;
        RECT 11.200 114.200 11.500 114.800 ;
        RECT 11.800 115.100 12.200 115.200 ;
        RECT 12.600 115.100 13.000 115.200 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 11.800 114.800 13.000 115.100 ;
        RECT 14.500 114.800 17.000 115.100 ;
        RECT 11.800 114.400 12.200 114.800 ;
        RECT 14.500 114.700 14.900 114.800 ;
        RECT 15.800 114.700 16.200 114.800 ;
        RECT 15.300 114.200 15.700 114.300 ;
        RECT 19.000 114.200 19.300 115.800 ;
        RECT 22.200 115.600 22.600 119.900 ;
        RECT 20.500 115.300 22.600 115.600 ;
        RECT 23.000 117.500 23.400 119.500 ;
        RECT 25.100 119.200 25.500 119.900 ;
        RECT 25.100 118.800 25.800 119.200 ;
        RECT 23.000 115.800 23.300 117.500 ;
        RECT 25.100 116.400 25.500 118.800 ;
        RECT 25.100 116.100 25.900 116.400 ;
        RECT 23.000 115.500 24.900 115.800 ;
        RECT 20.500 115.200 20.900 115.300 ;
        RECT 21.300 114.900 21.700 115.000 ;
        RECT 19.800 114.600 21.700 114.900 ;
        RECT 19.800 114.500 20.200 114.600 ;
        RECT 10.200 113.800 11.500 114.200 ;
        RECT 12.600 114.100 13.000 114.200 ;
        RECT 12.200 113.800 13.000 114.100 ;
        RECT 13.800 113.900 19.300 114.200 ;
        RECT 13.800 113.800 14.600 113.900 ;
        RECT 10.300 113.100 10.600 113.800 ;
        RECT 12.200 113.600 12.600 113.800 ;
        RECT 11.100 113.100 12.900 113.300 ;
        RECT 8.600 112.800 9.500 113.100 ;
        RECT 9.100 111.100 9.500 112.800 ;
        RECT 10.200 111.100 10.600 113.100 ;
        RECT 11.000 113.000 13.000 113.100 ;
        RECT 11.000 111.100 11.400 113.000 ;
        RECT 12.600 111.100 13.000 113.000 ;
        RECT 13.400 111.100 13.800 113.500 ;
        RECT 15.900 112.800 16.200 113.900 ;
        RECT 17.400 113.800 17.800 113.900 ;
        RECT 18.700 113.800 19.100 113.900 ;
        RECT 22.200 113.600 22.600 115.300 ;
        RECT 23.000 114.400 23.400 115.200 ;
        RECT 23.800 114.400 24.200 115.200 ;
        RECT 24.600 114.500 24.900 115.500 ;
        RECT 24.600 114.100 25.300 114.500 ;
        RECT 25.600 114.200 25.900 116.100 ;
        RECT 27.800 116.100 28.200 116.200 ;
        RECT 28.600 116.100 29.000 119.900 ;
        RECT 27.800 115.800 29.000 116.100 ;
        RECT 29.400 115.800 29.800 116.600 ;
        RECT 31.500 116.200 31.900 119.900 ;
        RECT 32.200 116.800 32.600 117.200 ;
        RECT 32.300 116.200 32.600 116.800 ;
        RECT 31.500 115.900 32.000 116.200 ;
        RECT 32.300 115.900 33.000 116.200 ;
        RECT 26.200 115.100 26.600 115.600 ;
        RECT 26.200 114.800 28.100 115.100 ;
        RECT 27.800 114.200 28.100 114.800 ;
        RECT 24.600 113.900 25.100 114.100 ;
        RECT 20.700 113.300 22.600 113.600 ;
        RECT 20.700 113.200 21.100 113.300 ;
        RECT 15.000 112.100 15.400 112.500 ;
        RECT 15.800 112.400 16.200 112.800 ;
        RECT 16.700 112.700 17.100 112.800 ;
        RECT 16.700 112.400 18.100 112.700 ;
        RECT 17.800 112.100 18.100 112.400 ;
        RECT 19.800 112.100 20.200 112.500 ;
        RECT 15.000 111.800 16.000 112.100 ;
        RECT 15.600 111.100 16.000 111.800 ;
        RECT 17.800 111.100 18.200 112.100 ;
        RECT 19.800 111.800 20.500 112.100 ;
        RECT 19.900 111.100 20.500 111.800 ;
        RECT 22.200 111.100 22.600 113.300 ;
        RECT 23.000 113.600 25.100 113.900 ;
        RECT 25.600 113.800 26.600 114.200 ;
        RECT 23.000 112.500 23.300 113.600 ;
        RECT 25.600 113.500 25.900 113.800 ;
        RECT 25.500 113.300 25.900 113.500 ;
        RECT 27.800 113.400 28.200 114.200 ;
        RECT 25.100 113.000 25.900 113.300 ;
        RECT 28.600 113.100 29.000 115.800 ;
        RECT 29.400 115.100 29.800 115.200 ;
        RECT 31.000 115.100 31.400 115.200 ;
        RECT 29.400 114.800 31.400 115.100 ;
        RECT 31.000 114.400 31.400 114.800 ;
        RECT 31.700 114.200 32.000 115.900 ;
        RECT 32.600 115.800 33.000 115.900 ;
        RECT 33.400 115.700 33.800 119.900 ;
        RECT 35.600 118.200 36.000 119.900 ;
        RECT 35.000 117.900 36.000 118.200 ;
        RECT 37.800 117.900 38.200 119.900 ;
        RECT 39.900 117.900 40.500 119.900 ;
        RECT 35.000 117.500 35.400 117.900 ;
        RECT 37.800 117.600 38.100 117.900 ;
        RECT 36.700 117.300 38.500 117.600 ;
        RECT 39.800 117.500 40.200 117.900 ;
        RECT 36.700 117.200 37.100 117.300 ;
        RECT 38.100 117.200 38.500 117.300 ;
        RECT 35.000 116.500 35.400 116.600 ;
        RECT 37.300 116.500 37.700 116.600 ;
        RECT 35.000 116.200 37.700 116.500 ;
        RECT 38.000 116.500 39.100 116.800 ;
        RECT 38.000 115.900 38.300 116.500 ;
        RECT 38.700 116.400 39.100 116.500 ;
        RECT 39.900 116.600 40.600 117.000 ;
        RECT 39.900 116.100 40.200 116.600 ;
        RECT 35.900 115.700 38.300 115.900 ;
        RECT 33.400 115.600 38.300 115.700 ;
        RECT 39.000 115.800 40.200 116.100 ;
        RECT 33.400 115.500 36.300 115.600 ;
        RECT 33.400 115.400 36.200 115.500 ;
        RECT 36.600 115.100 37.000 115.200 ;
        RECT 37.400 115.100 37.800 115.200 ;
        RECT 34.500 114.800 37.800 115.100 ;
        RECT 34.500 114.700 34.900 114.800 ;
        RECT 35.300 114.200 35.700 114.300 ;
        RECT 39.000 114.200 39.300 115.800 ;
        RECT 42.200 115.600 42.600 119.900 ;
        RECT 43.400 116.800 43.800 117.200 ;
        RECT 43.400 116.200 43.700 116.800 ;
        RECT 44.100 116.200 44.500 119.900 ;
        RECT 43.000 115.900 43.700 116.200 ;
        RECT 44.000 115.900 44.500 116.200 ;
        RECT 43.000 115.800 43.400 115.900 ;
        RECT 40.500 115.300 42.600 115.600 ;
        RECT 40.500 115.200 40.900 115.300 ;
        RECT 41.300 114.900 41.700 115.000 ;
        RECT 39.800 114.600 41.700 114.900 ;
        RECT 39.800 114.500 40.200 114.600 ;
        RECT 30.200 114.100 30.600 114.200 ;
        RECT 30.200 113.800 31.000 114.100 ;
        RECT 31.700 113.800 33.000 114.200 ;
        RECT 33.800 113.900 39.400 114.200 ;
        RECT 33.800 113.800 34.600 113.900 ;
        RECT 30.600 113.600 31.000 113.800 ;
        RECT 30.300 113.100 32.100 113.300 ;
        RECT 32.600 113.100 32.900 113.800 ;
        RECT 23.000 111.500 23.400 112.500 ;
        RECT 25.100 111.500 25.500 113.000 ;
        RECT 28.600 112.800 29.500 113.100 ;
        RECT 29.100 111.100 29.500 112.800 ;
        RECT 30.200 113.000 32.200 113.100 ;
        RECT 30.200 111.100 30.600 113.000 ;
        RECT 31.800 111.100 32.200 113.000 ;
        RECT 32.600 111.100 33.000 113.100 ;
        RECT 33.400 111.100 33.800 113.500 ;
        RECT 35.900 112.800 36.200 113.900 ;
        RECT 38.700 113.800 39.400 113.900 ;
        RECT 42.200 113.600 42.600 115.300 ;
        RECT 43.000 115.100 43.400 115.200 ;
        RECT 44.000 115.100 44.300 115.900 ;
        RECT 47.800 115.600 48.200 119.900 ;
        RECT 49.900 117.900 50.500 119.900 ;
        RECT 52.200 117.900 52.600 119.900 ;
        RECT 54.400 118.200 54.800 119.900 ;
        RECT 54.400 117.900 55.400 118.200 ;
        RECT 50.200 117.500 50.600 117.900 ;
        RECT 52.300 117.600 52.600 117.900 ;
        RECT 51.900 117.300 53.700 117.600 ;
        RECT 55.000 117.500 55.400 117.900 ;
        RECT 51.900 117.200 52.300 117.300 ;
        RECT 53.300 117.200 53.700 117.300 ;
        RECT 49.800 116.600 50.500 117.000 ;
        RECT 50.200 116.100 50.500 116.600 ;
        RECT 51.300 116.500 52.400 116.800 ;
        RECT 51.300 116.400 51.700 116.500 ;
        RECT 50.200 115.800 51.400 116.100 ;
        RECT 47.800 115.300 49.900 115.600 ;
        RECT 43.000 114.800 44.300 115.100 ;
        RECT 44.000 114.200 44.300 114.800 ;
        RECT 44.600 114.400 45.000 115.200 ;
        RECT 43.000 113.800 44.300 114.200 ;
        RECT 45.400 114.100 45.800 114.200 ;
        RECT 46.200 114.100 46.600 114.200 ;
        RECT 45.000 113.800 46.600 114.100 ;
        RECT 40.700 113.300 42.600 113.600 ;
        RECT 40.700 113.200 41.100 113.300 ;
        RECT 35.000 112.100 35.400 112.500 ;
        RECT 35.800 112.400 36.200 112.800 ;
        RECT 36.700 112.700 37.100 112.800 ;
        RECT 36.700 112.400 38.100 112.700 ;
        RECT 37.800 112.100 38.100 112.400 ;
        RECT 39.800 112.100 40.200 112.500 ;
        RECT 35.000 111.800 36.000 112.100 ;
        RECT 35.600 111.100 36.000 111.800 ;
        RECT 37.800 111.100 38.200 112.100 ;
        RECT 39.800 111.800 40.500 112.100 ;
        RECT 39.900 111.100 40.500 111.800 ;
        RECT 42.200 111.100 42.600 113.300 ;
        RECT 43.100 113.100 43.400 113.800 ;
        RECT 45.000 113.600 45.400 113.800 ;
        RECT 47.800 113.600 48.200 115.300 ;
        RECT 49.500 115.200 49.900 115.300 ;
        RECT 48.700 114.900 49.100 115.000 ;
        RECT 48.700 114.600 50.600 114.900 ;
        RECT 50.200 114.500 50.600 114.600 ;
        RECT 51.100 114.200 51.400 115.800 ;
        RECT 52.100 115.900 52.400 116.500 ;
        RECT 52.700 116.500 53.100 116.600 ;
        RECT 55.000 116.500 55.400 116.600 ;
        RECT 52.700 116.200 55.400 116.500 ;
        RECT 52.100 115.700 54.500 115.900 ;
        RECT 56.600 115.700 57.000 119.900 ;
        RECT 58.700 116.200 59.100 119.900 ;
        RECT 59.400 116.800 59.800 117.200 ;
        RECT 59.500 116.200 59.800 116.800 ;
        RECT 58.200 115.800 59.200 116.200 ;
        RECT 59.500 115.900 60.200 116.200 ;
        RECT 52.100 115.600 57.000 115.700 ;
        RECT 54.100 115.500 57.000 115.600 ;
        RECT 54.200 115.400 57.000 115.500 ;
        RECT 53.400 115.100 53.800 115.200 ;
        RECT 53.400 114.800 55.900 115.100 ;
        RECT 55.500 114.700 55.900 114.800 ;
        RECT 58.200 114.400 58.600 115.200 ;
        RECT 54.700 114.200 55.100 114.300 ;
        RECT 58.900 114.200 59.200 115.800 ;
        RECT 59.800 115.800 60.200 115.900 ;
        RECT 60.600 115.800 61.000 116.600 ;
        RECT 59.800 115.100 60.100 115.800 ;
        RECT 61.400 115.100 61.800 119.900 ;
        RECT 64.900 116.400 65.300 119.900 ;
        RECT 67.000 117.500 67.400 119.500 ;
        RECT 64.500 116.100 65.300 116.400 ;
        RECT 64.500 115.800 65.000 116.100 ;
        RECT 67.100 115.800 67.400 117.500 ;
        RECT 63.800 115.100 64.200 115.600 ;
        RECT 59.800 114.800 61.800 115.100 ;
        RECT 51.100 113.900 56.600 114.200 ;
        RECT 51.300 113.800 51.700 113.900 ;
        RECT 54.200 113.800 54.600 113.900 ;
        RECT 55.800 113.800 56.600 113.900 ;
        RECT 57.400 114.100 57.800 114.200 ;
        RECT 57.400 113.800 58.200 114.100 ;
        RECT 58.900 113.800 60.200 114.200 ;
        RECT 47.800 113.300 49.700 113.600 ;
        RECT 43.900 113.100 45.700 113.300 ;
        RECT 43.000 111.100 43.400 113.100 ;
        RECT 43.800 113.000 45.800 113.100 ;
        RECT 43.800 111.100 44.200 113.000 ;
        RECT 45.400 111.100 45.800 113.000 ;
        RECT 47.800 111.100 48.200 113.300 ;
        RECT 49.300 113.200 49.700 113.300 ;
        RECT 54.200 112.800 54.500 113.800 ;
        RECT 57.800 113.600 58.200 113.800 ;
        RECT 53.300 112.700 53.700 112.800 ;
        RECT 50.200 112.100 50.600 112.500 ;
        RECT 52.300 112.400 53.700 112.700 ;
        RECT 54.200 112.400 54.600 112.800 ;
        RECT 52.300 112.100 52.600 112.400 ;
        RECT 55.000 112.100 55.400 112.500 ;
        RECT 49.900 111.800 50.600 112.100 ;
        RECT 49.900 111.100 50.500 111.800 ;
        RECT 52.200 111.100 52.600 112.100 ;
        RECT 54.400 111.800 55.400 112.100 ;
        RECT 54.400 111.100 54.800 111.800 ;
        RECT 56.600 111.100 57.000 113.500 ;
        RECT 57.500 113.100 59.300 113.300 ;
        RECT 59.800 113.100 60.100 113.800 ;
        RECT 61.400 113.100 61.800 114.800 ;
        RECT 63.000 114.800 64.200 115.100 ;
        RECT 62.200 114.100 62.600 114.200 ;
        RECT 63.000 114.100 63.300 114.800 ;
        RECT 64.500 114.200 64.800 115.800 ;
        RECT 65.500 115.500 67.400 115.800 ;
        RECT 67.800 117.500 68.200 119.500 ;
        RECT 69.900 119.200 70.300 119.900 ;
        RECT 69.900 118.800 70.600 119.200 ;
        RECT 67.800 115.800 68.100 117.500 ;
        RECT 69.900 116.400 70.300 118.800 ;
        RECT 69.900 116.100 70.700 116.400 ;
        RECT 67.800 115.500 69.700 115.800 ;
        RECT 65.500 114.500 65.800 115.500 ;
        RECT 62.200 113.800 63.300 114.100 ;
        RECT 63.800 113.800 64.800 114.200 ;
        RECT 65.100 114.100 65.800 114.500 ;
        RECT 66.200 114.400 66.600 115.200 ;
        RECT 67.000 114.400 67.400 115.200 ;
        RECT 67.800 114.400 68.200 115.200 ;
        RECT 68.600 114.400 69.000 115.200 ;
        RECT 69.400 114.500 69.700 115.500 ;
        RECT 62.200 113.400 62.600 113.800 ;
        RECT 64.500 113.500 64.800 113.800 ;
        RECT 65.300 113.900 65.800 114.100 ;
        RECT 69.400 114.100 70.100 114.500 ;
        RECT 70.400 114.200 70.700 116.100 ;
        RECT 71.000 114.800 71.400 115.600 ;
        RECT 69.400 113.900 69.900 114.100 ;
        RECT 65.300 113.600 67.400 113.900 ;
        RECT 57.400 113.000 59.400 113.100 ;
        RECT 57.400 111.100 57.800 113.000 ;
        RECT 59.000 111.100 59.400 113.000 ;
        RECT 59.800 111.100 60.200 113.100 ;
        RECT 60.900 112.800 61.800 113.100 ;
        RECT 64.500 113.300 64.900 113.500 ;
        RECT 64.500 113.000 65.300 113.300 ;
        RECT 60.900 111.100 61.300 112.800 ;
        RECT 64.900 111.500 65.300 113.000 ;
        RECT 67.100 112.500 67.400 113.600 ;
        RECT 67.000 111.500 67.400 112.500 ;
        RECT 67.800 113.600 69.900 113.900 ;
        RECT 70.400 113.800 71.400 114.200 ;
        RECT 67.800 112.500 68.100 113.600 ;
        RECT 70.400 113.500 70.700 113.800 ;
        RECT 70.300 113.300 70.700 113.500 ;
        RECT 72.600 113.400 73.000 114.200 ;
        RECT 69.900 113.000 70.700 113.300 ;
        RECT 73.400 113.100 73.800 119.900 ;
        RECT 76.900 119.200 77.300 119.900 ;
        RECT 76.900 118.800 77.800 119.200 ;
        RECT 74.200 115.800 74.600 116.600 ;
        RECT 76.900 116.400 77.300 118.800 ;
        RECT 79.000 117.500 79.400 119.500 ;
        RECT 76.500 116.100 77.300 116.400 ;
        RECT 75.000 115.100 75.400 115.200 ;
        RECT 75.800 115.100 76.200 115.600 ;
        RECT 75.000 114.800 76.200 115.100 ;
        RECT 76.500 114.200 76.800 116.100 ;
        RECT 79.100 115.800 79.400 117.500 ;
        RECT 81.100 116.200 81.500 119.900 ;
        RECT 81.800 116.800 82.200 117.200 ;
        RECT 81.900 116.200 82.200 116.800 ;
        RECT 81.100 115.900 81.600 116.200 ;
        RECT 81.900 115.900 82.600 116.200 ;
        RECT 77.500 115.500 79.400 115.800 ;
        RECT 77.500 114.500 77.800 115.500 ;
        RECT 75.800 113.800 76.800 114.200 ;
        RECT 77.100 114.100 77.800 114.500 ;
        RECT 78.200 114.400 78.600 115.200 ;
        RECT 79.000 114.400 79.400 115.200 ;
        RECT 80.600 114.400 81.000 115.200 ;
        RECT 81.300 114.200 81.600 115.900 ;
        RECT 82.200 115.800 82.600 115.900 ;
        RECT 83.000 115.800 83.400 116.600 ;
        RECT 82.200 115.100 82.500 115.800 ;
        RECT 83.800 115.100 84.200 119.900 ;
        RECT 85.400 115.700 85.800 119.900 ;
        RECT 87.600 118.200 88.000 119.900 ;
        RECT 87.000 117.900 88.000 118.200 ;
        RECT 89.800 117.900 90.200 119.900 ;
        RECT 91.900 117.900 92.500 119.900 ;
        RECT 87.000 117.500 87.400 117.900 ;
        RECT 89.800 117.600 90.100 117.900 ;
        RECT 88.700 117.300 90.500 117.600 ;
        RECT 91.800 117.500 92.200 117.900 ;
        RECT 88.700 117.200 89.100 117.300 ;
        RECT 90.100 117.200 90.500 117.300 ;
        RECT 87.000 116.500 87.400 116.600 ;
        RECT 89.300 116.500 89.700 116.600 ;
        RECT 87.000 116.200 89.700 116.500 ;
        RECT 90.000 116.500 91.100 116.800 ;
        RECT 90.000 115.900 90.300 116.500 ;
        RECT 90.700 116.400 91.100 116.500 ;
        RECT 91.900 116.600 92.600 117.000 ;
        RECT 91.900 116.100 92.200 116.600 ;
        RECT 87.900 115.700 90.300 115.900 ;
        RECT 85.400 115.600 90.300 115.700 ;
        RECT 91.000 115.800 92.200 116.100 ;
        RECT 85.400 115.500 88.300 115.600 ;
        RECT 85.400 115.400 88.200 115.500 ;
        RECT 91.000 115.200 91.300 115.800 ;
        RECT 94.200 115.600 94.600 119.900 ;
        RECT 92.500 115.300 94.600 115.600 ;
        RECT 92.500 115.200 92.900 115.300 ;
        RECT 88.600 115.100 89.000 115.200 ;
        RECT 82.200 114.800 84.200 115.100 ;
        RECT 76.500 113.500 76.800 113.800 ;
        RECT 77.300 113.900 77.800 114.100 ;
        RECT 79.800 114.100 80.200 114.200 ;
        RECT 77.300 113.600 79.400 113.900 ;
        RECT 79.800 113.800 80.600 114.100 ;
        RECT 81.300 113.800 82.600 114.200 ;
        RECT 80.200 113.600 80.600 113.800 ;
        RECT 76.500 113.300 76.900 113.500 ;
        RECT 67.800 111.500 68.200 112.500 ;
        RECT 69.900 111.500 70.300 113.000 ;
        RECT 73.400 112.800 74.300 113.100 ;
        RECT 76.500 113.000 77.300 113.300 ;
        RECT 73.900 112.200 74.300 112.800 ;
        RECT 73.900 111.800 74.600 112.200 ;
        RECT 73.900 111.100 74.300 111.800 ;
        RECT 76.900 111.500 77.300 113.000 ;
        RECT 79.100 112.500 79.400 113.600 ;
        RECT 79.900 113.100 81.700 113.300 ;
        RECT 82.200 113.100 82.500 113.800 ;
        RECT 83.800 113.100 84.200 114.800 ;
        RECT 86.500 114.800 89.000 115.100 ;
        RECT 91.000 114.800 91.400 115.200 ;
        RECT 93.300 114.900 93.700 115.000 ;
        RECT 86.500 114.700 86.900 114.800 ;
        RECT 87.300 114.200 87.700 114.300 ;
        RECT 91.000 114.200 91.300 114.800 ;
        RECT 91.800 114.600 93.700 114.900 ;
        RECT 91.800 114.500 92.200 114.600 ;
        RECT 84.600 113.400 85.000 114.200 ;
        RECT 85.800 113.900 91.300 114.200 ;
        RECT 85.800 113.800 86.600 113.900 ;
        RECT 79.000 111.500 79.400 112.500 ;
        RECT 79.800 113.000 81.800 113.100 ;
        RECT 79.800 111.100 80.200 113.000 ;
        RECT 81.400 111.100 81.800 113.000 ;
        RECT 82.200 111.100 82.600 113.100 ;
        RECT 83.300 112.800 84.200 113.100 ;
        RECT 83.300 111.100 83.700 112.800 ;
        RECT 85.400 111.100 85.800 113.500 ;
        RECT 87.900 113.200 88.200 113.900 ;
        RECT 90.700 113.800 91.100 113.900 ;
        RECT 94.200 113.600 94.600 115.300 ;
        RECT 92.700 113.300 94.600 113.600 ;
        RECT 95.000 113.400 95.400 114.200 ;
        RECT 92.700 113.200 93.100 113.300 ;
        RECT 87.000 112.100 87.400 112.500 ;
        RECT 87.800 112.400 88.200 113.200 ;
        RECT 88.700 112.700 89.100 112.800 ;
        RECT 88.700 112.400 90.100 112.700 ;
        RECT 89.800 112.100 90.100 112.400 ;
        RECT 91.800 112.100 92.200 112.500 ;
        RECT 87.000 111.800 88.000 112.100 ;
        RECT 87.600 111.100 88.000 111.800 ;
        RECT 89.800 111.100 90.200 112.100 ;
        RECT 91.800 111.800 92.500 112.100 ;
        RECT 91.900 111.100 92.500 111.800 ;
        RECT 94.200 111.100 94.600 113.300 ;
        RECT 95.800 113.100 96.200 119.900 ;
        RECT 96.600 116.100 97.000 116.600 ;
        RECT 97.400 116.100 97.800 116.200 ;
        RECT 96.600 115.800 97.800 116.100 ;
        RECT 98.200 115.100 98.600 119.900 ;
        RECT 101.800 116.800 102.200 117.200 ;
        RECT 99.000 115.800 99.400 116.600 ;
        RECT 101.800 116.200 102.100 116.800 ;
        RECT 102.500 116.200 102.900 119.900 ;
        RECT 101.400 115.900 102.100 116.200 ;
        RECT 102.400 115.900 102.900 116.200 ;
        RECT 101.400 115.800 101.800 115.900 ;
        RECT 101.400 115.100 101.700 115.800 ;
        RECT 98.200 114.800 101.700 115.100 ;
        RECT 96.600 114.100 97.000 114.200 ;
        RECT 97.400 114.100 97.800 114.200 ;
        RECT 96.600 113.800 97.800 114.100 ;
        RECT 97.400 113.400 97.800 113.800 ;
        RECT 98.200 113.100 98.600 114.800 ;
        RECT 102.400 114.200 102.700 115.900 ;
        RECT 103.000 114.400 103.400 115.200 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 103.800 114.800 105.000 115.100 ;
        RECT 105.400 115.100 105.800 119.900 ;
        RECT 107.400 116.800 107.800 117.200 ;
        RECT 106.200 115.800 106.600 116.600 ;
        RECT 107.400 116.200 107.700 116.800 ;
        RECT 108.100 116.200 108.500 119.900 ;
        RECT 107.000 115.900 107.700 116.200 ;
        RECT 108.000 115.900 108.500 116.200 ;
        RECT 107.000 115.800 107.400 115.900 ;
        RECT 107.000 115.100 107.300 115.800 ;
        RECT 108.000 115.200 108.300 115.900 ;
        RECT 110.200 115.600 110.600 119.900 ;
        RECT 112.300 117.900 112.900 119.900 ;
        RECT 114.600 117.900 115.000 119.900 ;
        RECT 116.800 118.200 117.200 119.900 ;
        RECT 116.800 117.900 117.800 118.200 ;
        RECT 112.600 117.500 113.000 117.900 ;
        RECT 114.700 117.600 115.000 117.900 ;
        RECT 114.300 117.300 116.100 117.600 ;
        RECT 117.400 117.500 117.800 117.900 ;
        RECT 114.300 117.200 114.700 117.300 ;
        RECT 115.700 117.200 116.100 117.300 ;
        RECT 112.200 116.600 112.900 117.000 ;
        RECT 112.600 116.100 112.900 116.600 ;
        RECT 113.700 116.500 114.800 116.800 ;
        RECT 113.700 116.400 114.100 116.500 ;
        RECT 112.600 115.800 113.800 116.100 ;
        RECT 110.200 115.300 112.300 115.600 ;
        RECT 105.400 114.800 107.300 115.100 ;
        RECT 107.800 114.800 108.300 115.200 ;
        RECT 101.400 113.800 102.700 114.200 ;
        RECT 103.800 114.200 104.100 114.800 ;
        RECT 103.800 114.100 104.200 114.200 ;
        RECT 103.400 113.800 104.200 114.100 ;
        RECT 100.600 113.100 101.000 113.200 ;
        RECT 101.500 113.100 101.800 113.800 ;
        RECT 103.400 113.600 103.800 113.800 ;
        RECT 104.600 113.400 105.000 114.200 ;
        RECT 102.300 113.100 104.100 113.300 ;
        RECT 105.400 113.100 105.800 114.800 ;
        RECT 108.000 114.200 108.300 114.800 ;
        RECT 108.600 114.400 109.000 115.200 ;
        RECT 107.000 113.800 108.300 114.200 ;
        RECT 109.400 114.100 109.800 114.200 ;
        RECT 109.000 113.800 109.800 114.100 ;
        RECT 107.100 113.100 107.400 113.800 ;
        RECT 109.000 113.600 109.400 113.800 ;
        RECT 110.200 113.600 110.600 115.300 ;
        RECT 111.900 115.200 112.300 115.300 ;
        RECT 111.100 114.900 111.500 115.000 ;
        RECT 111.100 114.600 113.000 114.900 ;
        RECT 112.600 114.500 113.000 114.600 ;
        RECT 113.500 114.200 113.800 115.800 ;
        RECT 114.500 115.900 114.800 116.500 ;
        RECT 115.100 116.500 115.500 116.600 ;
        RECT 117.400 116.500 117.800 116.600 ;
        RECT 115.100 116.200 117.800 116.500 ;
        RECT 114.500 115.700 116.900 115.900 ;
        RECT 119.000 115.700 119.400 119.900 ;
        RECT 114.500 115.600 119.400 115.700 ;
        RECT 116.500 115.500 119.400 115.600 ;
        RECT 116.600 115.400 119.400 115.500 ;
        RECT 119.800 115.600 120.200 119.900 ;
        RECT 121.900 117.900 122.500 119.900 ;
        RECT 124.200 117.900 124.600 119.900 ;
        RECT 126.400 118.200 126.800 119.900 ;
        RECT 126.400 117.900 127.400 118.200 ;
        RECT 122.200 117.500 122.600 117.900 ;
        RECT 124.300 117.600 124.600 117.900 ;
        RECT 123.900 117.300 125.700 117.600 ;
        RECT 127.000 117.500 127.400 117.900 ;
        RECT 123.900 117.200 124.300 117.300 ;
        RECT 125.300 117.200 125.700 117.300 ;
        RECT 121.800 116.600 122.500 117.000 ;
        RECT 122.200 116.100 122.500 116.600 ;
        RECT 123.300 116.500 124.400 116.800 ;
        RECT 123.300 116.400 123.700 116.500 ;
        RECT 122.200 115.800 123.400 116.100 ;
        RECT 119.800 115.300 121.900 115.600 ;
        RECT 114.200 115.100 114.600 115.200 ;
        RECT 115.800 115.100 116.200 115.200 ;
        RECT 114.200 114.800 118.300 115.100 ;
        RECT 117.900 114.700 118.300 114.800 ;
        RECT 117.100 114.200 117.500 114.300 ;
        RECT 113.500 113.900 119.000 114.200 ;
        RECT 113.700 113.800 114.100 113.900 ;
        RECT 110.200 113.300 112.100 113.600 ;
        RECT 107.900 113.100 109.700 113.300 ;
        RECT 95.800 112.800 96.700 113.100 ;
        RECT 98.200 112.800 99.100 113.100 ;
        RECT 100.600 112.800 101.800 113.100 ;
        RECT 96.300 112.200 96.700 112.800 ;
        RECT 96.300 111.800 97.000 112.200 ;
        RECT 96.300 111.100 96.700 111.800 ;
        RECT 98.700 111.100 99.100 112.800 ;
        RECT 101.400 111.100 101.800 112.800 ;
        RECT 102.200 113.000 104.200 113.100 ;
        RECT 102.200 111.100 102.600 113.000 ;
        RECT 103.800 111.100 104.200 113.000 ;
        RECT 105.400 112.800 106.300 113.100 ;
        RECT 105.900 111.100 106.300 112.800 ;
        RECT 107.000 111.100 107.400 113.100 ;
        RECT 107.800 113.000 109.800 113.100 ;
        RECT 107.800 111.100 108.200 113.000 ;
        RECT 109.400 111.100 109.800 113.000 ;
        RECT 110.200 111.100 110.600 113.300 ;
        RECT 111.700 113.200 112.100 113.300 ;
        RECT 116.600 112.800 116.900 113.900 ;
        RECT 118.200 113.800 119.000 113.900 ;
        RECT 119.800 113.600 120.200 115.300 ;
        RECT 121.500 115.200 121.900 115.300 ;
        RECT 120.700 114.900 121.100 115.000 ;
        RECT 120.700 114.600 122.600 114.900 ;
        RECT 122.200 114.500 122.600 114.600 ;
        RECT 123.100 114.200 123.400 115.800 ;
        RECT 124.100 115.900 124.400 116.500 ;
        RECT 124.700 116.500 125.100 116.600 ;
        RECT 127.000 116.500 127.400 116.600 ;
        RECT 124.700 116.200 127.400 116.500 ;
        RECT 124.100 115.700 126.500 115.900 ;
        RECT 128.600 115.700 129.000 119.900 ;
        RECT 124.100 115.600 129.000 115.700 ;
        RECT 126.100 115.500 129.000 115.600 ;
        RECT 126.200 115.400 129.000 115.500 ;
        RECT 130.200 115.600 130.600 119.900 ;
        RECT 131.800 115.600 132.200 119.900 ;
        RECT 133.400 115.600 133.800 119.900 ;
        RECT 135.000 115.600 135.400 119.900 ;
        RECT 136.600 117.500 137.000 119.500 ;
        RECT 136.600 115.800 136.900 117.500 ;
        RECT 138.700 116.400 139.100 119.900 ;
        RECT 138.700 116.100 139.500 116.400 ;
        RECT 130.200 115.200 131.100 115.600 ;
        RECT 131.800 115.200 132.900 115.600 ;
        RECT 133.400 115.200 134.500 115.600 ;
        RECT 135.000 115.200 136.200 115.600 ;
        RECT 136.600 115.500 138.500 115.800 ;
        RECT 125.400 115.100 125.800 115.200 ;
        RECT 125.400 114.800 127.900 115.100 ;
        RECT 127.500 114.700 127.900 114.800 ;
        RECT 130.700 114.500 131.100 115.200 ;
        RECT 132.500 114.500 132.900 115.200 ;
        RECT 134.100 114.500 134.500 115.200 ;
        RECT 126.700 114.200 127.100 114.300 ;
        RECT 123.000 114.100 128.600 114.200 ;
        RECT 129.400 114.100 130.300 114.500 ;
        RECT 130.700 114.100 132.000 114.500 ;
        RECT 132.500 114.100 133.700 114.500 ;
        RECT 134.100 114.100 135.400 114.500 ;
        RECT 123.000 113.900 129.800 114.100 ;
        RECT 123.000 113.800 123.700 113.900 ;
        RECT 115.700 112.700 116.100 112.800 ;
        RECT 112.600 112.100 113.000 112.500 ;
        RECT 114.700 112.400 116.100 112.700 ;
        RECT 116.600 112.400 117.000 112.800 ;
        RECT 114.700 112.100 115.000 112.400 ;
        RECT 117.400 112.100 117.800 112.500 ;
        RECT 112.300 111.800 113.000 112.100 ;
        RECT 112.300 111.100 112.900 111.800 ;
        RECT 114.600 111.100 115.000 112.100 ;
        RECT 116.800 111.800 117.800 112.100 ;
        RECT 116.800 111.100 117.200 111.800 ;
        RECT 119.000 111.100 119.400 113.500 ;
        RECT 119.800 113.300 121.700 113.600 ;
        RECT 119.800 111.100 120.200 113.300 ;
        RECT 121.300 113.200 121.700 113.300 ;
        RECT 126.200 112.800 126.500 113.900 ;
        RECT 127.800 113.800 129.800 113.900 ;
        RECT 130.700 113.800 131.100 114.100 ;
        RECT 132.500 113.800 132.900 114.100 ;
        RECT 134.100 113.800 134.500 114.100 ;
        RECT 135.800 113.800 136.200 115.200 ;
        RECT 136.600 114.400 137.000 115.200 ;
        RECT 137.400 114.400 137.800 115.200 ;
        RECT 138.200 114.500 138.500 115.500 ;
        RECT 138.200 114.100 138.900 114.500 ;
        RECT 139.200 114.200 139.500 116.100 ;
        RECT 139.800 115.100 140.200 115.600 ;
        RECT 142.200 115.100 142.600 119.900 ;
        RECT 144.200 116.800 144.600 117.200 ;
        RECT 143.000 115.800 143.400 116.600 ;
        RECT 144.200 116.200 144.500 116.800 ;
        RECT 144.900 116.200 145.300 119.900 ;
        RECT 143.800 115.900 144.500 116.200 ;
        RECT 144.800 115.900 145.300 116.200 ;
        RECT 143.800 115.800 144.200 115.900 ;
        RECT 143.800 115.100 144.100 115.800 ;
        RECT 139.800 114.800 141.700 115.100 ;
        RECT 141.400 114.200 141.700 114.800 ;
        RECT 142.200 114.800 144.100 115.100 ;
        RECT 139.200 114.100 140.200 114.200 ;
        RECT 140.600 114.100 141.000 114.200 ;
        RECT 138.200 113.900 138.700 114.100 ;
        RECT 125.300 112.700 125.700 112.800 ;
        RECT 122.200 112.100 122.600 112.500 ;
        RECT 124.300 112.400 125.700 112.700 ;
        RECT 126.200 112.400 126.600 112.800 ;
        RECT 124.300 112.100 124.600 112.400 ;
        RECT 127.000 112.100 127.400 112.500 ;
        RECT 121.900 111.800 122.600 112.100 ;
        RECT 121.900 111.100 122.500 111.800 ;
        RECT 124.200 111.100 124.600 112.100 ;
        RECT 126.400 111.800 127.400 112.100 ;
        RECT 126.400 111.100 126.800 111.800 ;
        RECT 128.600 111.100 129.000 113.500 ;
        RECT 130.200 113.400 131.100 113.800 ;
        RECT 131.800 113.400 132.900 113.800 ;
        RECT 133.400 113.400 134.500 113.800 ;
        RECT 135.000 113.400 136.200 113.800 ;
        RECT 136.600 113.600 138.700 113.900 ;
        RECT 139.200 113.800 141.000 114.100 ;
        RECT 130.200 111.100 130.600 113.400 ;
        RECT 131.800 111.100 132.200 113.400 ;
        RECT 133.400 111.100 133.800 113.400 ;
        RECT 135.000 111.100 135.400 113.400 ;
        RECT 136.600 112.500 136.900 113.600 ;
        RECT 139.200 113.500 139.500 113.800 ;
        RECT 139.100 113.300 139.500 113.500 ;
        RECT 141.400 113.400 141.800 114.200 ;
        RECT 138.700 113.000 139.500 113.300 ;
        RECT 142.200 113.100 142.600 114.800 ;
        RECT 144.800 114.200 145.100 115.900 ;
        RECT 148.600 115.600 149.000 119.900 ;
        RECT 150.700 117.900 151.300 119.900 ;
        RECT 153.000 117.900 153.400 119.900 ;
        RECT 155.200 118.200 155.600 119.900 ;
        RECT 155.200 117.900 156.200 118.200 ;
        RECT 151.000 117.500 151.400 117.900 ;
        RECT 153.100 117.600 153.400 117.900 ;
        RECT 152.700 117.300 154.500 117.600 ;
        RECT 155.800 117.500 156.200 117.900 ;
        RECT 152.700 117.200 153.100 117.300 ;
        RECT 154.100 117.200 154.500 117.300 ;
        RECT 150.600 116.600 151.300 117.000 ;
        RECT 151.000 116.100 151.300 116.600 ;
        RECT 152.100 116.500 153.200 116.800 ;
        RECT 152.100 116.400 152.500 116.500 ;
        RECT 151.000 115.800 152.200 116.100 ;
        RECT 148.600 115.300 150.700 115.600 ;
        RECT 145.400 115.100 145.800 115.200 ;
        RECT 146.200 115.100 146.600 115.200 ;
        RECT 145.400 114.800 146.600 115.100 ;
        RECT 145.400 114.400 145.800 114.800 ;
        RECT 143.800 113.800 145.100 114.200 ;
        RECT 146.200 114.100 146.600 114.200 ;
        RECT 147.000 114.100 147.400 114.200 ;
        RECT 145.800 113.800 147.400 114.100 ;
        RECT 143.900 113.100 144.200 113.800 ;
        RECT 145.800 113.600 146.200 113.800 ;
        RECT 148.600 113.600 149.000 115.300 ;
        RECT 150.300 115.200 150.700 115.300 ;
        RECT 151.900 115.200 152.200 115.800 ;
        RECT 152.900 115.900 153.200 116.500 ;
        RECT 153.500 116.500 153.900 116.600 ;
        RECT 155.800 116.500 156.200 116.600 ;
        RECT 153.500 116.200 156.200 116.500 ;
        RECT 152.900 115.700 155.300 115.900 ;
        RECT 157.400 115.700 157.800 119.900 ;
        RECT 158.600 116.800 159.000 117.200 ;
        RECT 158.600 116.200 158.900 116.800 ;
        RECT 159.300 116.200 159.700 119.900 ;
        RECT 158.200 115.900 158.900 116.200 ;
        RECT 159.200 115.900 159.700 116.200 ;
        RECT 158.200 115.800 158.600 115.900 ;
        RECT 152.900 115.600 157.800 115.700 ;
        RECT 154.900 115.500 157.800 115.600 ;
        RECT 155.000 115.400 157.800 115.500 ;
        RECT 149.500 114.900 149.900 115.000 ;
        RECT 149.500 114.600 151.400 114.900 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 154.200 115.100 154.600 115.200 ;
        RECT 154.200 114.800 156.700 115.100 ;
        RECT 151.000 114.500 151.400 114.600 ;
        RECT 151.900 114.200 152.200 114.800 ;
        RECT 155.000 114.700 155.400 114.800 ;
        RECT 156.300 114.700 156.700 114.800 ;
        RECT 155.500 114.200 155.900 114.300 ;
        RECT 159.200 114.200 159.500 115.900 ;
        RECT 161.400 115.700 161.800 119.900 ;
        RECT 163.600 118.200 164.000 119.900 ;
        RECT 163.000 117.900 164.000 118.200 ;
        RECT 165.800 117.900 166.200 119.900 ;
        RECT 167.900 117.900 168.500 119.900 ;
        RECT 163.000 117.500 163.400 117.900 ;
        RECT 165.800 117.600 166.100 117.900 ;
        RECT 164.700 117.300 166.500 117.600 ;
        RECT 167.800 117.500 168.200 117.900 ;
        RECT 164.700 117.200 165.100 117.300 ;
        RECT 166.100 117.200 166.500 117.300 ;
        RECT 163.000 116.500 163.400 116.600 ;
        RECT 165.300 116.500 165.700 116.600 ;
        RECT 163.000 116.200 165.700 116.500 ;
        RECT 166.000 116.500 167.100 116.800 ;
        RECT 166.000 115.900 166.300 116.500 ;
        RECT 166.700 116.400 167.100 116.500 ;
        RECT 167.900 116.600 168.600 117.000 ;
        RECT 167.900 116.100 168.200 116.600 ;
        RECT 163.900 115.700 166.300 115.900 ;
        RECT 161.400 115.600 166.300 115.700 ;
        RECT 167.000 115.800 168.200 116.100 ;
        RECT 161.400 115.500 164.300 115.600 ;
        RECT 161.400 115.400 164.200 115.500 ;
        RECT 159.800 114.400 160.200 115.200 ;
        RECT 164.600 115.100 165.000 115.200 ;
        RECT 162.500 114.800 165.000 115.100 ;
        RECT 162.500 114.700 162.900 114.800 ;
        RECT 163.300 114.200 163.700 114.300 ;
        RECT 167.000 114.200 167.300 115.800 ;
        RECT 170.200 115.600 170.600 119.900 ;
        RECT 172.300 117.200 172.700 119.900 ;
        RECT 171.800 116.800 172.700 117.200 ;
        RECT 173.000 116.800 173.400 117.200 ;
        RECT 172.300 116.200 172.700 116.800 ;
        RECT 173.100 116.200 173.400 116.800 ;
        RECT 172.300 115.900 172.800 116.200 ;
        RECT 173.100 115.900 173.800 116.200 ;
        RECT 168.500 115.300 170.600 115.600 ;
        RECT 168.500 115.200 168.900 115.300 ;
        RECT 169.300 114.900 169.700 115.000 ;
        RECT 167.800 114.600 169.700 114.900 ;
        RECT 167.800 114.500 168.200 114.600 ;
        RECT 151.900 113.900 157.400 114.200 ;
        RECT 152.100 113.800 152.500 113.900 ;
        RECT 148.600 113.300 150.500 113.600 ;
        RECT 144.700 113.100 146.500 113.300 ;
        RECT 136.600 111.500 137.000 112.500 ;
        RECT 138.700 111.500 139.100 113.000 ;
        RECT 142.200 112.800 143.100 113.100 ;
        RECT 142.700 111.100 143.100 112.800 ;
        RECT 143.800 111.100 144.200 113.100 ;
        RECT 144.600 113.000 146.600 113.100 ;
        RECT 144.600 111.100 145.000 113.000 ;
        RECT 146.200 111.100 146.600 113.000 ;
        RECT 148.600 111.100 149.000 113.300 ;
        RECT 150.100 113.200 150.500 113.300 ;
        RECT 155.000 112.800 155.300 113.900 ;
        RECT 156.600 113.800 157.400 113.900 ;
        RECT 158.200 113.800 159.500 114.200 ;
        RECT 160.600 114.100 161.000 114.200 ;
        RECT 160.200 113.800 161.000 114.100 ;
        RECT 161.800 113.900 167.300 114.200 ;
        RECT 161.800 113.800 162.600 113.900 ;
        RECT 154.100 112.700 154.500 112.800 ;
        RECT 151.000 112.100 151.400 112.500 ;
        RECT 153.100 112.400 154.500 112.700 ;
        RECT 155.000 112.400 155.400 112.800 ;
        RECT 153.100 112.100 153.400 112.400 ;
        RECT 155.800 112.100 156.200 112.500 ;
        RECT 150.700 111.800 151.400 112.100 ;
        RECT 150.700 111.100 151.300 111.800 ;
        RECT 153.000 111.100 153.400 112.100 ;
        RECT 155.200 111.800 156.200 112.100 ;
        RECT 155.200 111.100 155.600 111.800 ;
        RECT 157.400 111.100 157.800 113.500 ;
        RECT 158.300 113.100 158.600 113.800 ;
        RECT 160.200 113.600 160.600 113.800 ;
        RECT 159.100 113.100 160.900 113.300 ;
        RECT 158.200 111.100 158.600 113.100 ;
        RECT 159.000 113.000 161.000 113.100 ;
        RECT 159.000 111.100 159.400 113.000 ;
        RECT 160.600 111.100 161.000 113.000 ;
        RECT 161.400 111.100 161.800 113.500 ;
        RECT 163.900 112.800 164.200 113.900 ;
        RECT 166.700 113.800 167.100 113.900 ;
        RECT 170.200 113.600 170.600 115.300 ;
        RECT 171.800 114.400 172.200 115.200 ;
        RECT 172.500 114.200 172.800 115.900 ;
        RECT 173.400 115.800 173.800 115.900 ;
        RECT 174.200 115.800 174.600 116.600 ;
        RECT 173.400 115.100 173.700 115.800 ;
        RECT 175.000 115.100 175.400 119.900 ;
        RECT 176.600 117.500 177.000 119.500 ;
        RECT 178.700 119.200 179.100 119.900 ;
        RECT 178.200 118.800 179.100 119.200 ;
        RECT 176.600 115.800 176.900 117.500 ;
        RECT 178.700 116.400 179.100 118.800 ;
        RECT 182.200 116.400 182.600 119.900 ;
        RECT 178.700 116.100 179.500 116.400 ;
        RECT 176.600 115.500 178.500 115.800 ;
        RECT 173.400 114.800 175.400 115.100 ;
        RECT 171.000 114.100 171.400 114.200 ;
        RECT 171.000 113.800 171.800 114.100 ;
        RECT 172.500 113.800 173.800 114.200 ;
        RECT 171.400 113.600 171.800 113.800 ;
        RECT 168.700 113.300 170.600 113.600 ;
        RECT 168.700 113.200 169.100 113.300 ;
        RECT 163.000 112.100 163.400 112.500 ;
        RECT 163.800 112.400 164.200 112.800 ;
        RECT 164.700 112.700 165.100 112.800 ;
        RECT 164.700 112.400 166.100 112.700 ;
        RECT 165.800 112.100 166.100 112.400 ;
        RECT 167.800 112.100 168.200 112.500 ;
        RECT 163.000 111.800 164.000 112.100 ;
        RECT 163.600 111.100 164.000 111.800 ;
        RECT 165.800 111.100 166.200 112.100 ;
        RECT 167.800 111.800 168.500 112.100 ;
        RECT 167.900 111.100 168.500 111.800 ;
        RECT 170.200 111.100 170.600 113.300 ;
        RECT 171.100 113.100 172.900 113.300 ;
        RECT 173.400 113.100 173.700 113.800 ;
        RECT 175.000 113.100 175.400 114.800 ;
        RECT 176.600 114.400 177.000 115.200 ;
        RECT 177.400 114.400 177.800 115.200 ;
        RECT 178.200 114.500 178.500 115.500 ;
        RECT 175.800 113.400 176.200 114.200 ;
        RECT 178.200 114.100 178.900 114.500 ;
        RECT 179.200 114.200 179.500 116.100 ;
        RECT 182.100 115.900 182.600 116.400 ;
        RECT 183.800 116.200 184.200 119.900 ;
        RECT 182.900 115.900 184.200 116.200 ;
        RECT 179.800 115.100 180.200 115.600 ;
        RECT 181.400 115.100 181.800 115.200 ;
        RECT 179.800 114.800 181.800 115.100 ;
        RECT 182.100 114.200 182.400 115.900 ;
        RECT 182.900 114.900 183.200 115.900 ;
        RECT 182.700 114.500 183.200 114.900 ;
        RECT 178.200 113.900 178.700 114.100 ;
        RECT 176.600 113.600 178.700 113.900 ;
        RECT 179.200 113.800 180.200 114.200 ;
        RECT 182.100 113.800 182.600 114.200 ;
        RECT 171.000 113.000 173.000 113.100 ;
        RECT 171.000 111.100 171.400 113.000 ;
        RECT 172.600 111.100 173.000 113.000 ;
        RECT 173.400 111.100 173.800 113.100 ;
        RECT 174.500 112.800 175.400 113.100 ;
        RECT 174.500 111.100 174.900 112.800 ;
        RECT 176.600 112.500 176.900 113.600 ;
        RECT 179.200 113.500 179.500 113.800 ;
        RECT 179.100 113.300 179.500 113.500 ;
        RECT 178.700 113.000 179.500 113.300 ;
        RECT 182.100 113.100 182.400 113.800 ;
        RECT 182.900 113.700 183.200 114.500 ;
        RECT 183.700 114.800 184.200 115.200 ;
        RECT 183.700 114.400 184.100 114.800 ;
        RECT 182.900 113.400 184.200 113.700 ;
        RECT 184.600 113.400 185.000 114.200 ;
        RECT 176.600 111.500 177.000 112.500 ;
        RECT 178.700 111.500 179.100 113.000 ;
        RECT 182.100 112.800 182.600 113.100 ;
        RECT 182.200 111.100 182.600 112.800 ;
        RECT 183.800 111.100 184.200 113.400 ;
        RECT 185.400 113.100 185.800 119.900 ;
        RECT 186.200 115.800 186.600 116.600 ;
        RECT 187.000 115.800 187.400 116.600 ;
        RECT 187.800 116.100 188.200 119.900 ;
        RECT 189.800 116.800 190.200 117.200 ;
        RECT 189.800 116.200 190.100 116.800 ;
        RECT 190.500 116.200 190.900 119.900 ;
        RECT 189.400 116.100 190.100 116.200 ;
        RECT 187.800 115.900 190.100 116.100 ;
        RECT 190.400 115.900 190.900 116.200 ;
        RECT 193.900 116.200 194.300 119.900 ;
        RECT 194.600 116.800 195.000 117.200 ;
        RECT 194.700 116.200 195.000 116.800 ;
        RECT 193.900 115.900 194.400 116.200 ;
        RECT 194.700 115.900 195.400 116.200 ;
        RECT 187.800 115.800 189.800 115.900 ;
        RECT 187.800 113.100 188.200 115.800 ;
        RECT 190.400 114.200 190.700 115.900 ;
        RECT 191.000 114.400 191.400 115.200 ;
        RECT 193.400 114.400 193.800 115.200 ;
        RECT 194.100 114.200 194.400 115.900 ;
        RECT 195.000 115.800 195.400 115.900 ;
        RECT 195.800 115.800 196.200 116.600 ;
        RECT 195.000 115.100 195.300 115.800 ;
        RECT 196.600 115.100 197.000 119.900 ;
        RECT 195.000 114.800 197.000 115.100 ;
        RECT 188.600 113.400 189.000 114.200 ;
        RECT 189.400 113.800 190.700 114.200 ;
        RECT 191.800 114.100 192.200 114.200 ;
        RECT 192.600 114.100 193.000 114.200 ;
        RECT 191.400 113.800 193.400 114.100 ;
        RECT 194.100 113.800 195.400 114.200 ;
        RECT 189.500 113.100 189.800 113.800 ;
        RECT 191.400 113.600 191.800 113.800 ;
        RECT 193.000 113.600 193.400 113.800 ;
        RECT 190.300 113.100 192.100 113.300 ;
        RECT 192.700 113.100 194.500 113.300 ;
        RECT 195.000 113.100 195.300 113.800 ;
        RECT 196.600 113.100 197.000 114.800 ;
        RECT 199.800 115.600 200.200 119.900 ;
        RECT 201.900 117.900 202.500 119.900 ;
        RECT 204.200 117.900 204.600 119.900 ;
        RECT 206.400 118.200 206.800 119.900 ;
        RECT 206.400 117.900 207.400 118.200 ;
        RECT 202.200 117.500 202.600 117.900 ;
        RECT 204.300 117.600 204.600 117.900 ;
        RECT 203.900 117.300 205.700 117.600 ;
        RECT 207.000 117.500 207.400 117.900 ;
        RECT 203.900 117.200 204.300 117.300 ;
        RECT 205.300 117.200 205.700 117.300 ;
        RECT 201.800 116.600 202.500 117.000 ;
        RECT 202.200 116.100 202.500 116.600 ;
        RECT 203.300 116.500 204.400 116.800 ;
        RECT 203.300 116.400 203.700 116.500 ;
        RECT 202.200 115.800 203.400 116.100 ;
        RECT 199.800 115.300 201.900 115.600 ;
        RECT 197.400 114.100 197.800 114.200 ;
        RECT 199.800 114.100 200.200 115.300 ;
        RECT 201.500 115.200 201.900 115.300 ;
        RECT 200.700 114.900 201.100 115.000 ;
        RECT 200.700 114.600 202.600 114.900 ;
        RECT 202.200 114.500 202.600 114.600 ;
        RECT 197.400 113.800 200.200 114.100 ;
        RECT 203.100 114.200 203.400 115.800 ;
        RECT 204.100 115.900 204.400 116.500 ;
        RECT 204.700 116.500 205.100 116.600 ;
        RECT 207.000 116.500 207.400 116.600 ;
        RECT 204.700 116.200 207.400 116.500 ;
        RECT 204.100 115.700 206.500 115.900 ;
        RECT 208.600 115.700 209.000 119.900 ;
        RECT 204.100 115.600 209.000 115.700 ;
        RECT 206.100 115.500 209.000 115.600 ;
        RECT 206.200 115.400 209.000 115.500 ;
        RECT 209.400 115.700 209.800 119.900 ;
        RECT 211.600 118.200 212.000 119.900 ;
        RECT 211.000 117.900 212.000 118.200 ;
        RECT 213.800 117.900 214.200 119.900 ;
        RECT 215.900 117.900 216.500 119.900 ;
        RECT 211.000 117.500 211.400 117.900 ;
        RECT 213.800 117.600 214.100 117.900 ;
        RECT 212.700 117.300 214.500 117.600 ;
        RECT 215.800 117.500 216.200 117.900 ;
        RECT 212.700 117.200 213.100 117.300 ;
        RECT 214.100 117.200 214.500 117.300 ;
        RECT 211.000 116.500 211.400 116.600 ;
        RECT 213.300 116.500 213.700 116.600 ;
        RECT 211.000 116.200 213.700 116.500 ;
        RECT 214.000 116.500 215.100 116.800 ;
        RECT 214.000 115.900 214.300 116.500 ;
        RECT 214.700 116.400 215.100 116.500 ;
        RECT 215.900 116.600 216.600 117.000 ;
        RECT 215.900 116.100 216.200 116.600 ;
        RECT 211.900 115.700 214.300 115.900 ;
        RECT 209.400 115.600 214.300 115.700 ;
        RECT 215.000 115.800 216.200 116.100 ;
        RECT 209.400 115.500 212.300 115.600 ;
        RECT 209.400 115.400 212.200 115.500 ;
        RECT 203.800 115.100 204.200 115.200 ;
        RECT 205.400 115.100 205.800 115.200 ;
        RECT 212.600 115.100 213.000 115.200 ;
        RECT 203.800 114.800 207.900 115.100 ;
        RECT 207.500 114.700 207.900 114.800 ;
        RECT 210.500 114.800 213.000 115.100 ;
        RECT 210.500 114.700 210.900 114.800 ;
        RECT 206.700 114.200 207.100 114.300 ;
        RECT 211.300 114.200 211.700 114.300 ;
        RECT 215.000 114.200 215.300 115.800 ;
        RECT 218.200 115.600 218.600 119.900 ;
        RECT 220.300 116.200 220.700 119.900 ;
        RECT 221.000 116.800 221.400 117.200 ;
        RECT 221.100 116.200 221.400 116.800 ;
        RECT 223.000 116.400 223.400 119.900 ;
        RECT 219.800 115.800 220.800 116.200 ;
        RECT 221.100 115.900 221.800 116.200 ;
        RECT 221.400 115.800 221.800 115.900 ;
        RECT 222.900 115.900 223.400 116.400 ;
        RECT 224.600 116.200 225.000 119.900 ;
        RECT 223.700 115.900 225.000 116.200 ;
        RECT 225.400 117.500 225.800 119.500 ;
        RECT 216.500 115.300 218.600 115.600 ;
        RECT 216.500 115.200 216.900 115.300 ;
        RECT 217.300 114.900 217.700 115.000 ;
        RECT 215.800 114.600 217.700 114.900 ;
        RECT 215.800 114.500 216.200 114.600 ;
        RECT 203.100 113.900 208.600 114.200 ;
        RECT 203.300 113.800 203.700 113.900 ;
        RECT 206.200 113.800 206.600 113.900 ;
        RECT 207.800 113.800 208.600 113.900 ;
        RECT 209.800 113.900 215.400 114.200 ;
        RECT 209.800 113.800 210.600 113.900 ;
        RECT 197.400 113.400 197.800 113.800 ;
        RECT 199.800 113.600 200.200 113.800 ;
        RECT 185.400 112.800 186.300 113.100 ;
        RECT 185.900 112.200 186.300 112.800 ;
        RECT 187.300 112.800 188.200 113.100 ;
        RECT 185.900 111.800 186.600 112.200 ;
        RECT 185.900 111.100 186.300 111.800 ;
        RECT 187.300 111.100 187.700 112.800 ;
        RECT 189.400 111.100 189.800 113.100 ;
        RECT 190.200 113.000 192.200 113.100 ;
        RECT 190.200 111.100 190.600 113.000 ;
        RECT 191.800 111.100 192.200 113.000 ;
        RECT 192.600 113.000 194.600 113.100 ;
        RECT 192.600 111.100 193.000 113.000 ;
        RECT 194.200 111.100 194.600 113.000 ;
        RECT 195.000 111.100 195.400 113.100 ;
        RECT 196.100 112.800 197.000 113.100 ;
        RECT 199.800 113.300 201.700 113.600 ;
        RECT 196.100 111.100 196.500 112.800 ;
        RECT 199.800 111.100 200.200 113.300 ;
        RECT 201.300 113.200 201.700 113.300 ;
        RECT 206.200 112.800 206.500 113.800 ;
        RECT 205.300 112.700 205.700 112.800 ;
        RECT 202.200 112.100 202.600 112.500 ;
        RECT 204.300 112.400 205.700 112.700 ;
        RECT 206.200 112.400 206.600 112.800 ;
        RECT 204.300 112.100 204.600 112.400 ;
        RECT 207.000 112.100 207.400 112.500 ;
        RECT 201.900 111.800 202.600 112.100 ;
        RECT 201.900 111.100 202.500 111.800 ;
        RECT 204.200 111.100 204.600 112.100 ;
        RECT 206.400 111.800 207.400 112.100 ;
        RECT 206.400 111.100 206.800 111.800 ;
        RECT 208.600 111.100 209.000 113.500 ;
        RECT 209.400 111.100 209.800 113.500 ;
        RECT 211.900 112.800 212.200 113.900 ;
        RECT 214.700 113.800 215.400 113.900 ;
        RECT 218.200 113.600 218.600 115.300 ;
        RECT 219.800 114.400 220.200 115.200 ;
        RECT 220.500 114.200 220.800 115.800 ;
        RECT 222.200 114.800 222.600 115.200 ;
        RECT 219.000 114.100 219.400 114.200 ;
        RECT 219.000 113.800 219.800 114.100 ;
        RECT 220.500 113.800 221.800 114.200 ;
        RECT 222.200 114.100 222.500 114.800 ;
        RECT 222.900 114.200 223.200 115.900 ;
        RECT 223.700 114.900 224.000 115.900 ;
        RECT 225.400 115.800 225.700 117.500 ;
        RECT 227.500 116.400 227.900 119.900 ;
        RECT 230.200 117.500 230.600 119.500 ;
        RECT 227.500 116.100 228.300 116.400 ;
        RECT 225.400 115.500 227.300 115.800 ;
        RECT 223.500 114.500 224.000 114.900 ;
        RECT 222.900 114.100 223.400 114.200 ;
        RECT 222.200 113.800 223.400 114.100 ;
        RECT 219.400 113.600 219.800 113.800 ;
        RECT 216.700 113.300 218.600 113.600 ;
        RECT 216.700 113.200 217.100 113.300 ;
        RECT 211.000 112.100 211.400 112.500 ;
        RECT 211.800 112.400 212.200 112.800 ;
        RECT 212.700 112.700 213.100 112.800 ;
        RECT 212.700 112.400 214.100 112.700 ;
        RECT 213.800 112.100 214.100 112.400 ;
        RECT 215.800 112.100 216.200 112.500 ;
        RECT 211.000 111.800 212.000 112.100 ;
        RECT 211.600 111.100 212.000 111.800 ;
        RECT 213.800 111.100 214.200 112.100 ;
        RECT 215.800 111.800 216.500 112.100 ;
        RECT 215.900 111.100 216.500 111.800 ;
        RECT 218.200 111.100 218.600 113.300 ;
        RECT 219.100 113.100 220.900 113.300 ;
        RECT 221.400 113.100 221.700 113.800 ;
        RECT 222.900 113.100 223.200 113.800 ;
        RECT 223.700 113.700 224.000 114.500 ;
        RECT 224.500 114.800 225.000 115.200 ;
        RECT 224.500 114.400 224.900 114.800 ;
        RECT 225.400 114.400 225.800 115.200 ;
        RECT 226.200 114.400 226.600 115.200 ;
        RECT 227.000 114.500 227.300 115.500 ;
        RECT 227.000 114.100 227.700 114.500 ;
        RECT 228.000 114.200 228.300 116.100 ;
        RECT 230.200 115.800 230.500 117.500 ;
        RECT 232.300 116.400 232.700 119.900 ;
        RECT 232.300 116.100 233.100 116.400 ;
        RECT 228.600 114.800 229.000 115.600 ;
        RECT 230.200 115.500 232.100 115.800 ;
        RECT 230.200 114.400 230.600 115.200 ;
        RECT 231.000 114.400 231.400 115.200 ;
        RECT 231.800 114.500 232.100 115.500 ;
        RECT 227.000 113.900 227.500 114.100 ;
        RECT 223.700 113.400 225.000 113.700 ;
        RECT 219.000 113.000 221.000 113.100 ;
        RECT 219.000 111.100 219.400 113.000 ;
        RECT 220.600 111.100 221.000 113.000 ;
        RECT 221.400 111.100 221.800 113.100 ;
        RECT 222.900 112.800 223.400 113.100 ;
        RECT 223.000 111.100 223.400 112.800 ;
        RECT 224.600 111.100 225.000 113.400 ;
        RECT 225.400 113.600 227.500 113.900 ;
        RECT 228.000 113.800 229.000 114.200 ;
        RECT 231.800 114.100 232.500 114.500 ;
        RECT 232.800 114.200 233.100 116.100 ;
        RECT 235.000 116.200 235.400 119.900 ;
        RECT 236.600 116.400 237.000 119.900 ;
        RECT 235.000 115.900 236.300 116.200 ;
        RECT 236.600 115.900 237.100 116.400 ;
        RECT 233.400 114.800 233.800 115.600 ;
        RECT 235.000 114.800 235.500 115.200 ;
        RECT 235.100 114.400 235.500 114.800 ;
        RECT 236.000 114.900 236.300 115.900 ;
        RECT 236.000 114.500 236.500 114.900 ;
        RECT 231.800 113.900 232.300 114.100 ;
        RECT 225.400 112.500 225.700 113.600 ;
        RECT 228.000 113.500 228.300 113.800 ;
        RECT 227.900 113.300 228.300 113.500 ;
        RECT 227.500 113.000 228.300 113.300 ;
        RECT 230.200 113.600 232.300 113.900 ;
        RECT 232.800 113.800 233.800 114.200 ;
        RECT 225.400 111.500 225.800 112.500 ;
        RECT 227.500 112.200 227.900 113.000 ;
        RECT 227.000 111.800 227.900 112.200 ;
        RECT 227.500 111.500 227.900 111.800 ;
        RECT 230.200 112.500 230.500 113.600 ;
        RECT 232.800 113.500 233.100 113.800 ;
        RECT 236.000 113.700 236.300 114.500 ;
        RECT 236.800 114.200 237.100 115.900 ;
        RECT 236.600 113.800 237.100 114.200 ;
        RECT 232.700 113.300 233.100 113.500 ;
        RECT 232.300 113.200 233.100 113.300 ;
        RECT 231.800 113.000 233.100 113.200 ;
        RECT 235.000 113.400 236.300 113.700 ;
        RECT 231.800 112.800 232.700 113.000 ;
        RECT 230.200 111.500 230.600 112.500 ;
        RECT 232.300 111.500 232.700 112.800 ;
        RECT 235.000 111.100 235.400 113.400 ;
        RECT 236.800 113.100 237.100 113.800 ;
        RECT 238.200 113.400 238.600 114.200 ;
        RECT 236.600 112.800 237.100 113.100 ;
        RECT 239.000 113.100 239.400 119.900 ;
        RECT 239.800 115.800 240.200 116.600 ;
        RECT 240.600 115.700 241.000 119.900 ;
        RECT 242.800 118.200 243.200 119.900 ;
        RECT 242.200 117.900 243.200 118.200 ;
        RECT 245.000 117.900 245.400 119.900 ;
        RECT 247.100 117.900 247.700 119.900 ;
        RECT 242.200 117.500 242.600 117.900 ;
        RECT 245.000 117.600 245.300 117.900 ;
        RECT 243.900 117.300 245.700 117.600 ;
        RECT 247.000 117.500 247.400 117.900 ;
        RECT 243.900 117.200 244.300 117.300 ;
        RECT 245.300 117.200 245.700 117.300 ;
        RECT 242.200 116.500 242.600 116.600 ;
        RECT 244.500 116.500 244.900 116.600 ;
        RECT 242.200 116.200 244.900 116.500 ;
        RECT 245.200 116.500 246.300 116.800 ;
        RECT 245.200 115.900 245.500 116.500 ;
        RECT 245.900 116.400 246.300 116.500 ;
        RECT 247.100 116.600 247.800 117.000 ;
        RECT 247.100 116.100 247.400 116.600 ;
        RECT 243.100 115.700 245.500 115.900 ;
        RECT 240.600 115.600 245.500 115.700 ;
        RECT 246.200 115.800 247.400 116.100 ;
        RECT 240.600 115.500 243.500 115.600 ;
        RECT 240.600 115.400 243.400 115.500 ;
        RECT 243.800 115.100 244.200 115.200 ;
        RECT 241.700 114.800 244.200 115.100 ;
        RECT 241.700 114.700 242.100 114.800 ;
        RECT 243.000 114.700 243.400 114.800 ;
        RECT 242.500 114.200 242.900 114.300 ;
        RECT 246.200 114.200 246.500 115.800 ;
        RECT 249.400 115.600 249.800 119.900 ;
        RECT 247.700 115.300 249.800 115.600 ;
        RECT 247.700 115.200 248.100 115.300 ;
        RECT 248.500 114.900 248.900 115.000 ;
        RECT 247.000 114.600 248.900 114.900 ;
        RECT 247.000 114.500 247.400 114.600 ;
        RECT 241.000 113.900 246.500 114.200 ;
        RECT 241.000 113.800 241.800 113.900 ;
        RECT 239.000 112.800 239.900 113.100 ;
        RECT 236.600 111.100 237.000 112.800 ;
        RECT 239.500 111.100 239.900 112.800 ;
        RECT 240.600 111.100 241.000 113.500 ;
        RECT 243.100 112.800 243.400 113.900 ;
        RECT 245.900 113.800 246.300 113.900 ;
        RECT 249.400 113.600 249.800 115.300 ;
        RECT 247.900 113.300 249.800 113.600 ;
        RECT 247.900 113.200 248.300 113.300 ;
        RECT 242.200 112.100 242.600 112.500 ;
        RECT 243.000 112.400 243.400 112.800 ;
        RECT 243.900 112.700 244.300 112.800 ;
        RECT 243.900 112.400 245.300 112.700 ;
        RECT 245.000 112.100 245.300 112.400 ;
        RECT 247.000 112.100 247.400 112.500 ;
        RECT 242.200 111.800 243.200 112.100 ;
        RECT 242.800 111.100 243.200 111.800 ;
        RECT 245.000 111.100 245.400 112.100 ;
        RECT 247.000 111.800 247.700 112.100 ;
        RECT 247.100 111.100 247.700 111.800 ;
        RECT 249.400 111.100 249.800 113.300 ;
        RECT 0.600 107.500 1.000 109.900 ;
        RECT 2.800 109.200 3.200 109.900 ;
        RECT 2.200 108.900 3.200 109.200 ;
        RECT 5.000 108.900 5.400 109.900 ;
        RECT 7.100 109.200 7.700 109.900 ;
        RECT 7.000 108.900 7.700 109.200 ;
        RECT 2.200 108.500 2.600 108.900 ;
        RECT 5.000 108.600 5.300 108.900 ;
        RECT 3.000 108.200 3.400 108.600 ;
        RECT 3.900 108.300 5.300 108.600 ;
        RECT 7.000 108.500 7.400 108.900 ;
        RECT 3.900 108.200 4.300 108.300 ;
        RECT 1.000 107.100 1.800 107.200 ;
        RECT 3.100 107.100 3.400 108.200 ;
        RECT 7.900 107.700 8.300 107.800 ;
        RECT 9.400 107.700 9.800 109.900 ;
        RECT 11.000 108.200 11.400 109.900 ;
        RECT 7.900 107.400 9.800 107.700 ;
        RECT 5.900 107.100 6.300 107.200 ;
        RECT 9.400 107.100 9.800 107.400 ;
        RECT 10.900 107.900 11.400 108.200 ;
        RECT 10.900 107.200 11.200 107.900 ;
        RECT 12.600 107.600 13.000 109.900 ;
        RECT 11.700 107.300 13.000 107.600 ;
        RECT 13.400 107.700 13.800 109.900 ;
        RECT 15.500 109.200 16.100 109.900 ;
        RECT 15.500 108.900 16.200 109.200 ;
        RECT 17.800 108.900 18.200 109.900 ;
        RECT 20.000 109.200 20.400 109.900 ;
        RECT 20.000 108.900 21.000 109.200 ;
        RECT 15.800 108.500 16.200 108.900 ;
        RECT 17.900 108.600 18.200 108.900 ;
        RECT 17.900 108.300 19.300 108.600 ;
        RECT 18.900 108.200 19.300 108.300 ;
        RECT 19.800 108.200 20.200 108.600 ;
        RECT 20.600 108.500 21.000 108.900 ;
        RECT 14.900 107.700 15.300 107.800 ;
        RECT 13.400 107.400 15.300 107.700 ;
        RECT 10.200 107.100 10.600 107.200 ;
        RECT 1.000 106.800 6.500 107.100 ;
        RECT 2.500 106.700 2.900 106.800 ;
        RECT 1.700 106.200 2.100 106.300 ;
        RECT 3.000 106.200 3.400 106.300 ;
        RECT 1.700 105.900 4.200 106.200 ;
        RECT 3.800 105.800 4.200 105.900 ;
        RECT 0.600 105.500 3.400 105.600 ;
        RECT 0.600 105.400 3.500 105.500 ;
        RECT 0.600 105.300 5.500 105.400 ;
        RECT 0.600 101.100 1.000 105.300 ;
        RECT 3.100 105.100 5.500 105.300 ;
        RECT 2.200 104.500 4.900 104.800 ;
        RECT 2.200 104.400 2.600 104.500 ;
        RECT 4.500 104.400 4.900 104.500 ;
        RECT 5.200 104.500 5.500 105.100 ;
        RECT 6.200 105.200 6.500 106.800 ;
        RECT 9.400 106.800 10.600 107.100 ;
        RECT 10.900 106.800 11.400 107.200 ;
        RECT 7.000 106.400 7.400 106.500 ;
        RECT 7.000 106.100 8.900 106.400 ;
        RECT 8.500 106.000 8.900 106.100 ;
        RECT 7.700 105.700 8.100 105.800 ;
        RECT 9.400 105.700 9.800 106.800 ;
        RECT 7.700 105.400 9.800 105.700 ;
        RECT 6.200 104.900 7.400 105.200 ;
        RECT 5.900 104.500 6.300 104.600 ;
        RECT 5.200 104.200 6.300 104.500 ;
        RECT 7.100 104.400 7.400 104.900 ;
        RECT 7.100 104.000 7.800 104.400 ;
        RECT 3.900 103.700 4.300 103.800 ;
        RECT 5.300 103.700 5.700 103.800 ;
        RECT 2.200 103.100 2.600 103.500 ;
        RECT 3.900 103.400 5.700 103.700 ;
        RECT 5.000 103.100 5.300 103.400 ;
        RECT 7.000 103.100 7.400 103.500 ;
        RECT 2.200 102.800 3.200 103.100 ;
        RECT 2.800 101.100 3.200 102.800 ;
        RECT 5.000 101.100 5.400 103.100 ;
        RECT 7.100 101.100 7.700 103.100 ;
        RECT 9.400 101.100 9.800 105.400 ;
        RECT 10.900 105.100 11.200 106.800 ;
        RECT 11.700 106.500 12.000 107.300 ;
        RECT 11.500 106.100 12.000 106.500 ;
        RECT 11.700 105.100 12.000 106.100 ;
        RECT 12.500 106.200 12.900 106.600 ;
        RECT 12.500 105.800 13.000 106.200 ;
        RECT 13.400 105.700 13.800 107.400 ;
        RECT 16.900 107.100 17.300 107.200 ;
        RECT 18.200 107.100 18.600 107.200 ;
        RECT 19.800 107.100 20.100 108.200 ;
        RECT 22.200 107.500 22.600 109.900 ;
        RECT 24.300 108.200 24.700 109.900 ;
        RECT 23.800 107.900 24.700 108.200 ;
        RECT 25.400 107.900 25.800 109.900 ;
        RECT 26.200 108.000 26.600 109.900 ;
        RECT 27.800 108.000 28.200 109.900 ;
        RECT 26.200 107.900 28.200 108.000 ;
        RECT 21.400 107.100 22.200 107.200 ;
        RECT 16.700 106.800 22.200 107.100 ;
        RECT 23.000 106.800 23.400 107.600 ;
        RECT 15.800 106.400 16.200 106.500 ;
        RECT 14.300 106.100 16.200 106.400 ;
        RECT 14.300 106.000 14.700 106.100 ;
        RECT 15.100 105.700 15.500 105.800 ;
        RECT 13.400 105.400 15.500 105.700 ;
        RECT 10.900 104.600 11.400 105.100 ;
        RECT 11.700 104.800 13.000 105.100 ;
        RECT 11.000 101.100 11.400 104.600 ;
        RECT 12.600 101.100 13.000 104.800 ;
        RECT 13.400 101.100 13.800 105.400 ;
        RECT 16.700 105.200 17.000 106.800 ;
        RECT 20.300 106.700 20.700 106.800 ;
        RECT 19.800 106.200 20.200 106.300 ;
        RECT 21.100 106.200 21.500 106.300 ;
        RECT 19.000 105.900 21.500 106.200 ;
        RECT 23.000 106.200 23.300 106.800 ;
        RECT 19.000 105.800 19.400 105.900 ;
        RECT 23.000 105.800 23.400 106.200 ;
        RECT 23.800 106.100 24.200 107.900 ;
        RECT 25.500 107.200 25.800 107.900 ;
        RECT 26.300 107.700 28.100 107.900 ;
        RECT 28.600 107.700 29.000 109.900 ;
        RECT 30.700 109.200 31.300 109.900 ;
        RECT 30.700 108.900 31.400 109.200 ;
        RECT 33.000 108.900 33.400 109.900 ;
        RECT 35.200 109.200 35.600 109.900 ;
        RECT 35.200 108.900 36.200 109.200 ;
        RECT 31.000 108.500 31.400 108.900 ;
        RECT 33.100 108.600 33.400 108.900 ;
        RECT 33.100 108.300 34.500 108.600 ;
        RECT 34.100 108.200 34.500 108.300 ;
        RECT 35.000 108.200 35.400 108.600 ;
        RECT 35.800 108.500 36.200 108.900 ;
        RECT 30.100 107.700 30.500 107.800 ;
        RECT 28.600 107.400 30.500 107.700 ;
        RECT 27.400 107.200 27.800 107.400 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 25.400 107.100 26.700 107.200 ;
        RECT 24.600 106.800 26.700 107.100 ;
        RECT 27.400 106.900 28.200 107.200 ;
        RECT 27.800 106.800 28.200 106.900 ;
        RECT 23.800 105.800 25.700 106.100 ;
        RECT 19.800 105.500 22.600 105.600 ;
        RECT 19.700 105.400 22.600 105.500 ;
        RECT 15.800 104.900 17.000 105.200 ;
        RECT 17.700 105.300 22.600 105.400 ;
        RECT 17.700 105.100 20.100 105.300 ;
        RECT 15.800 104.400 16.100 104.900 ;
        RECT 15.400 104.000 16.100 104.400 ;
        RECT 16.900 104.500 17.300 104.600 ;
        RECT 17.700 104.500 18.000 105.100 ;
        RECT 16.900 104.200 18.000 104.500 ;
        RECT 18.300 104.500 21.000 104.800 ;
        RECT 18.300 104.400 18.700 104.500 ;
        RECT 20.600 104.400 21.000 104.500 ;
        RECT 17.500 103.700 17.900 103.800 ;
        RECT 18.900 103.700 19.300 103.800 ;
        RECT 15.800 103.100 16.200 103.500 ;
        RECT 17.500 103.400 19.300 103.700 ;
        RECT 17.900 103.100 18.200 103.400 ;
        RECT 20.600 103.100 21.000 103.500 ;
        RECT 15.500 101.100 16.100 103.100 ;
        RECT 17.800 101.100 18.200 103.100 ;
        RECT 20.000 102.800 21.000 103.100 ;
        RECT 20.000 101.100 20.400 102.800 ;
        RECT 22.200 101.100 22.600 105.300 ;
        RECT 23.800 101.100 24.200 105.800 ;
        RECT 25.400 105.200 25.700 105.800 ;
        RECT 24.600 104.400 25.000 105.200 ;
        RECT 25.400 105.100 25.800 105.200 ;
        RECT 26.400 105.100 26.700 106.800 ;
        RECT 27.000 105.800 27.400 106.600 ;
        RECT 28.600 105.700 29.000 107.400 ;
        RECT 32.100 107.100 32.500 107.200 ;
        RECT 34.200 107.100 34.600 107.200 ;
        RECT 35.000 107.100 35.300 108.200 ;
        RECT 37.400 107.500 37.800 109.900 ;
        RECT 39.000 107.600 39.400 109.900 ;
        RECT 40.600 107.600 41.000 109.900 ;
        RECT 42.200 107.600 42.600 109.900 ;
        RECT 43.800 107.600 44.200 109.900 ;
        RECT 45.700 109.200 46.100 109.900 ;
        RECT 45.400 108.800 46.100 109.200 ;
        RECT 45.700 108.200 46.100 108.800 ;
        RECT 49.400 108.500 49.800 109.500 ;
        RECT 45.700 107.900 46.600 108.200 ;
        RECT 38.200 107.200 39.400 107.600 ;
        RECT 39.900 107.200 41.000 107.600 ;
        RECT 41.500 107.200 42.600 107.600 ;
        RECT 43.300 107.200 44.200 107.600 ;
        RECT 36.600 107.100 37.400 107.200 ;
        RECT 31.900 106.800 37.400 107.100 ;
        RECT 31.000 106.400 31.400 106.500 ;
        RECT 29.500 106.100 31.400 106.400 ;
        RECT 29.500 106.000 29.900 106.100 ;
        RECT 30.300 105.700 30.700 105.800 ;
        RECT 28.600 105.400 30.700 105.700 ;
        RECT 25.400 104.800 26.100 105.100 ;
        RECT 26.400 104.800 26.900 105.100 ;
        RECT 25.800 104.200 26.100 104.800 ;
        RECT 25.800 103.800 26.200 104.200 ;
        RECT 26.500 101.100 26.900 104.800 ;
        RECT 28.600 101.100 29.000 105.400 ;
        RECT 31.900 105.200 32.200 106.800 ;
        RECT 35.500 106.700 35.900 106.800 ;
        RECT 36.300 106.200 36.700 106.300 ;
        RECT 32.600 106.100 33.000 106.200 ;
        RECT 34.200 106.100 36.700 106.200 ;
        RECT 32.600 105.900 36.700 106.100 ;
        RECT 32.600 105.800 34.600 105.900 ;
        RECT 38.200 105.800 38.600 107.200 ;
        RECT 39.900 106.900 40.300 107.200 ;
        RECT 41.500 106.900 41.900 107.200 ;
        RECT 43.300 106.900 43.700 107.200 ;
        RECT 39.000 106.500 40.300 106.900 ;
        RECT 40.700 106.500 41.900 106.900 ;
        RECT 42.400 106.500 43.700 106.900 ;
        RECT 39.900 105.800 40.300 106.500 ;
        RECT 41.500 105.800 41.900 106.500 ;
        RECT 43.300 105.800 43.700 106.500 ;
        RECT 35.000 105.500 37.800 105.600 ;
        RECT 34.900 105.400 37.800 105.500 ;
        RECT 38.200 105.400 39.400 105.800 ;
        RECT 39.900 105.400 41.000 105.800 ;
        RECT 41.500 105.400 42.600 105.800 ;
        RECT 43.300 105.400 44.200 105.800 ;
        RECT 31.000 104.900 32.200 105.200 ;
        RECT 32.900 105.300 37.800 105.400 ;
        RECT 32.900 105.100 35.300 105.300 ;
        RECT 31.000 104.400 31.300 104.900 ;
        RECT 30.600 104.000 31.300 104.400 ;
        RECT 32.100 104.500 32.500 104.600 ;
        RECT 32.900 104.500 33.200 105.100 ;
        RECT 32.100 104.200 33.200 104.500 ;
        RECT 33.500 104.500 36.200 104.800 ;
        RECT 33.500 104.400 33.900 104.500 ;
        RECT 35.800 104.400 36.200 104.500 ;
        RECT 32.700 103.700 33.100 103.800 ;
        RECT 34.100 103.700 34.500 103.800 ;
        RECT 31.000 103.100 31.400 103.500 ;
        RECT 32.700 103.400 34.500 103.700 ;
        RECT 33.100 103.100 33.400 103.400 ;
        RECT 35.800 103.100 36.200 103.500 ;
        RECT 30.700 101.100 31.300 103.100 ;
        RECT 33.000 101.100 33.400 103.100 ;
        RECT 35.200 102.800 36.200 103.100 ;
        RECT 35.200 101.100 35.600 102.800 ;
        RECT 37.400 101.100 37.800 105.300 ;
        RECT 39.000 101.100 39.400 105.400 ;
        RECT 40.600 101.100 41.000 105.400 ;
        RECT 42.200 101.100 42.600 105.400 ;
        RECT 43.800 101.100 44.200 105.400 ;
        RECT 45.400 104.400 45.800 105.200 ;
        RECT 46.200 101.100 46.600 107.900 ;
        RECT 47.000 107.100 47.400 107.600 ;
        RECT 49.400 107.400 49.700 108.500 ;
        RECT 51.500 108.000 51.900 109.500 ;
        RECT 51.500 107.700 52.300 108.000 ;
        RECT 51.900 107.500 52.300 107.700 ;
        RECT 47.800 107.100 48.200 107.200 ;
        RECT 49.400 107.100 51.500 107.400 ;
        RECT 47.000 106.800 48.200 107.100 ;
        RECT 51.000 106.900 51.500 107.100 ;
        RECT 52.000 107.200 52.300 107.500 ;
        RECT 54.200 107.700 54.600 109.900 ;
        RECT 56.300 109.200 56.900 109.900 ;
        RECT 56.300 108.900 57.000 109.200 ;
        RECT 58.600 108.900 59.000 109.900 ;
        RECT 60.800 109.200 61.200 109.900 ;
        RECT 60.800 108.900 61.800 109.200 ;
        RECT 56.600 108.500 57.000 108.900 ;
        RECT 58.700 108.600 59.000 108.900 ;
        RECT 58.700 108.300 60.100 108.600 ;
        RECT 59.700 108.200 60.100 108.300 ;
        RECT 60.600 108.200 61.000 108.600 ;
        RECT 61.400 108.500 61.800 108.900 ;
        RECT 55.700 107.700 56.100 107.800 ;
        RECT 54.200 107.400 56.200 107.700 ;
        RECT 49.400 105.800 49.800 106.600 ;
        RECT 50.200 105.800 50.600 106.600 ;
        RECT 51.000 106.500 51.700 106.900 ;
        RECT 52.000 106.800 53.000 107.200 ;
        RECT 51.000 105.500 51.300 106.500 ;
        RECT 49.400 105.200 51.300 105.500 ;
        RECT 49.400 103.500 49.700 105.200 ;
        RECT 52.000 104.900 52.300 106.800 ;
        RECT 52.600 106.100 53.000 106.200 ;
        RECT 54.200 106.100 54.600 107.400 ;
        RECT 55.800 106.800 56.200 107.400 ;
        RECT 57.700 107.100 58.100 107.200 ;
        RECT 59.000 107.100 59.400 107.200 ;
        RECT 60.600 107.100 60.900 108.200 ;
        RECT 63.000 107.500 63.400 109.900 ;
        RECT 64.100 108.200 64.500 109.900 ;
        RECT 64.100 107.900 65.000 108.200 ;
        RECT 66.200 107.900 66.600 109.900 ;
        RECT 67.000 108.000 67.400 109.900 ;
        RECT 68.600 108.000 69.000 109.900 ;
        RECT 67.000 107.900 69.000 108.000 ;
        RECT 69.400 108.000 69.800 109.900 ;
        RECT 71.000 108.000 71.400 109.900 ;
        RECT 69.400 107.900 71.400 108.000 ;
        RECT 71.800 107.900 72.200 109.900 ;
        RECT 72.900 108.200 73.300 109.900 ;
        RECT 72.900 107.900 73.800 108.200 ;
        RECT 62.200 107.100 63.000 107.200 ;
        RECT 57.500 106.800 63.000 107.100 ;
        RECT 56.600 106.400 57.000 106.500 ;
        RECT 52.600 105.800 54.600 106.100 ;
        RECT 55.100 106.100 57.000 106.400 ;
        RECT 55.100 106.000 55.500 106.100 ;
        RECT 52.600 105.400 53.000 105.800 ;
        RECT 54.200 105.700 54.600 105.800 ;
        RECT 55.900 105.700 56.300 105.800 ;
        RECT 54.200 105.400 56.300 105.700 ;
        RECT 51.500 104.600 52.300 104.900 ;
        RECT 49.400 101.500 49.800 103.500 ;
        RECT 51.500 102.200 51.900 104.600 ;
        RECT 51.000 101.800 51.900 102.200 ;
        RECT 51.500 101.100 51.900 101.800 ;
        RECT 54.200 101.100 54.600 105.400 ;
        RECT 57.500 105.200 57.800 106.800 ;
        RECT 61.100 106.700 61.500 106.800 ;
        RECT 60.600 106.200 61.000 106.300 ;
        RECT 61.900 106.200 62.300 106.300 ;
        RECT 59.800 105.900 62.300 106.200 ;
        RECT 59.800 105.800 60.200 105.900 ;
        RECT 60.600 105.500 63.400 105.600 ;
        RECT 60.500 105.400 63.400 105.500 ;
        RECT 56.600 104.900 57.800 105.200 ;
        RECT 58.500 105.300 63.400 105.400 ;
        RECT 58.500 105.100 60.900 105.300 ;
        RECT 56.600 104.400 56.900 104.900 ;
        RECT 56.200 104.000 56.900 104.400 ;
        RECT 57.700 104.500 58.100 104.600 ;
        RECT 58.500 104.500 58.800 105.100 ;
        RECT 57.700 104.200 58.800 104.500 ;
        RECT 59.100 104.500 61.800 104.800 ;
        RECT 59.100 104.400 59.500 104.500 ;
        RECT 61.400 104.400 61.800 104.500 ;
        RECT 58.300 103.700 58.700 103.800 ;
        RECT 59.700 103.700 60.100 103.800 ;
        RECT 56.600 103.100 57.000 103.500 ;
        RECT 58.300 103.400 60.100 103.700 ;
        RECT 58.700 103.100 59.000 103.400 ;
        RECT 61.400 103.100 61.800 103.500 ;
        RECT 56.300 101.100 56.900 103.100 ;
        RECT 58.600 101.100 59.000 103.100 ;
        RECT 60.800 102.800 61.800 103.100 ;
        RECT 60.800 101.100 61.200 102.800 ;
        RECT 63.000 101.100 63.400 105.300 ;
        RECT 63.800 104.400 64.200 105.200 ;
        RECT 64.600 105.100 65.000 107.900 ;
        RECT 65.400 106.800 65.800 107.600 ;
        RECT 66.300 107.200 66.600 107.900 ;
        RECT 67.100 107.700 68.900 107.900 ;
        RECT 69.500 107.700 71.300 107.900 ;
        RECT 68.200 107.200 68.600 107.400 ;
        RECT 69.800 107.200 70.200 107.400 ;
        RECT 71.800 107.200 72.100 107.900 ;
        RECT 66.200 106.800 67.500 107.200 ;
        RECT 68.200 107.100 69.000 107.200 ;
        RECT 69.400 107.100 70.200 107.200 ;
        RECT 68.200 106.900 70.200 107.100 ;
        RECT 70.900 107.100 72.200 107.200 ;
        RECT 72.600 107.100 73.000 107.200 ;
        RECT 68.600 106.800 69.800 106.900 ;
        RECT 70.900 106.800 73.000 107.100 ;
        RECT 66.200 105.100 66.600 105.200 ;
        RECT 67.200 105.100 67.500 106.800 ;
        RECT 67.800 105.800 68.200 106.600 ;
        RECT 70.200 105.800 70.600 106.600 ;
        RECT 70.900 105.100 71.200 106.800 ;
        RECT 73.400 106.100 73.800 107.900 ;
        RECT 75.000 107.700 75.400 109.900 ;
        RECT 77.100 109.200 77.700 109.900 ;
        RECT 77.100 108.900 77.800 109.200 ;
        RECT 79.400 108.900 79.800 109.900 ;
        RECT 81.600 109.200 82.000 109.900 ;
        RECT 81.600 108.900 82.600 109.200 ;
        RECT 77.400 108.500 77.800 108.900 ;
        RECT 79.500 108.600 79.800 108.900 ;
        RECT 79.500 108.300 80.900 108.600 ;
        RECT 80.500 108.200 80.900 108.300 ;
        RECT 81.400 107.800 81.800 108.600 ;
        RECT 82.200 108.500 82.600 108.900 ;
        RECT 76.500 107.700 76.900 107.800 ;
        RECT 74.200 107.100 74.600 107.600 ;
        RECT 75.000 107.400 76.900 107.700 ;
        RECT 75.000 107.100 75.400 107.400 ;
        RECT 78.500 107.100 78.900 107.200 ;
        RECT 81.400 107.100 81.700 107.800 ;
        RECT 83.800 107.500 84.200 109.900 ;
        RECT 84.600 107.500 85.000 109.900 ;
        RECT 86.800 109.200 87.200 109.900 ;
        RECT 86.200 108.900 87.200 109.200 ;
        RECT 89.000 108.900 89.400 109.900 ;
        RECT 91.100 109.200 91.700 109.900 ;
        RECT 91.000 108.900 91.700 109.200 ;
        RECT 86.200 108.500 86.600 108.900 ;
        RECT 89.000 108.600 89.300 108.900 ;
        RECT 87.000 108.200 87.400 108.600 ;
        RECT 87.900 108.300 89.300 108.600 ;
        RECT 91.000 108.500 91.400 108.900 ;
        RECT 87.900 108.200 88.300 108.300 ;
        RECT 83.000 107.100 83.800 107.200 ;
        RECT 85.000 107.100 85.800 107.200 ;
        RECT 87.100 107.100 87.400 108.200 ;
        RECT 91.900 107.700 92.300 107.800 ;
        RECT 93.400 107.700 93.800 109.900 ;
        RECT 94.200 108.000 94.600 109.900 ;
        RECT 95.800 108.000 96.200 109.900 ;
        RECT 94.200 107.900 96.200 108.000 ;
        RECT 96.600 107.900 97.000 109.900 ;
        RECT 97.700 108.200 98.100 109.900 ;
        RECT 100.600 109.100 101.000 109.200 ;
        RECT 101.700 109.100 102.100 109.900 ;
        RECT 100.600 108.800 102.100 109.100 ;
        RECT 101.700 108.200 102.100 108.800 ;
        RECT 104.100 108.200 104.500 109.900 ;
        RECT 107.500 109.200 107.900 109.900 ;
        RECT 108.900 109.200 109.300 109.900 ;
        RECT 107.500 108.800 108.200 109.200 ;
        RECT 108.600 108.800 109.300 109.200 ;
        RECT 107.500 108.200 107.900 108.800 ;
        RECT 97.700 107.900 98.600 108.200 ;
        RECT 101.700 107.900 102.600 108.200 ;
        RECT 104.100 107.900 105.000 108.200 ;
        RECT 94.300 107.700 96.100 107.900 ;
        RECT 91.900 107.400 93.800 107.700 ;
        RECT 89.900 107.100 90.300 107.200 ;
        RECT 74.200 106.800 75.400 107.100 ;
        RECT 71.800 105.800 73.800 106.100 ;
        RECT 71.800 105.200 72.100 105.800 ;
        RECT 71.800 105.100 72.200 105.200 ;
        RECT 64.600 104.800 66.900 105.100 ;
        RECT 67.200 104.800 67.700 105.100 ;
        RECT 64.600 101.100 65.000 104.800 ;
        RECT 66.600 104.200 66.900 104.800 ;
        RECT 66.600 103.800 67.000 104.200 ;
        RECT 67.300 101.100 67.700 104.800 ;
        RECT 70.700 104.800 71.200 105.100 ;
        RECT 71.500 104.800 72.200 105.100 ;
        RECT 70.700 101.100 71.100 104.800 ;
        RECT 71.500 104.200 71.800 104.800 ;
        RECT 72.600 104.400 73.000 105.200 ;
        RECT 71.400 103.800 71.800 104.200 ;
        RECT 73.400 101.100 73.800 105.800 ;
        RECT 75.000 105.700 75.400 106.800 ;
        RECT 78.300 106.800 90.500 107.100 ;
        RECT 77.400 106.400 77.800 106.500 ;
        RECT 75.900 106.100 77.800 106.400 ;
        RECT 75.900 106.000 76.300 106.100 ;
        RECT 76.700 105.700 77.100 105.800 ;
        RECT 75.000 105.400 77.100 105.700 ;
        RECT 75.000 101.100 75.400 105.400 ;
        RECT 78.300 105.200 78.600 106.800 ;
        RECT 81.900 106.700 82.300 106.800 ;
        RECT 86.500 106.700 86.900 106.800 ;
        RECT 82.700 106.200 83.100 106.300 ;
        RECT 79.800 106.100 80.200 106.200 ;
        RECT 80.600 106.100 83.100 106.200 ;
        RECT 79.800 105.900 83.100 106.100 ;
        RECT 85.700 106.200 86.100 106.300 ;
        RECT 87.000 106.200 87.400 106.300 ;
        RECT 85.700 105.900 88.200 106.200 ;
        RECT 79.800 105.800 81.000 105.900 ;
        RECT 87.800 105.800 88.200 105.900 ;
        RECT 81.400 105.500 84.200 105.600 ;
        RECT 81.300 105.400 84.200 105.500 ;
        RECT 77.400 104.900 78.600 105.200 ;
        RECT 79.300 105.300 84.200 105.400 ;
        RECT 79.300 105.100 81.700 105.300 ;
        RECT 77.400 104.400 77.700 104.900 ;
        RECT 77.000 104.000 77.700 104.400 ;
        RECT 78.500 104.500 78.900 104.600 ;
        RECT 79.300 104.500 79.600 105.100 ;
        RECT 78.500 104.200 79.600 104.500 ;
        RECT 79.900 104.500 82.600 104.800 ;
        RECT 79.900 104.400 80.300 104.500 ;
        RECT 82.200 104.400 82.600 104.500 ;
        RECT 79.100 103.700 79.500 103.800 ;
        RECT 80.500 103.700 80.900 103.800 ;
        RECT 77.400 103.100 77.800 103.500 ;
        RECT 79.100 103.400 80.900 103.700 ;
        RECT 79.500 103.100 79.800 103.400 ;
        RECT 82.200 103.100 82.600 103.500 ;
        RECT 77.100 101.100 77.700 103.100 ;
        RECT 79.400 101.100 79.800 103.100 ;
        RECT 81.600 102.800 82.600 103.100 ;
        RECT 81.600 101.100 82.000 102.800 ;
        RECT 83.800 101.100 84.200 105.300 ;
        RECT 84.600 105.500 87.400 105.600 ;
        RECT 84.600 105.400 87.500 105.500 ;
        RECT 84.600 105.300 89.500 105.400 ;
        RECT 84.600 101.100 85.000 105.300 ;
        RECT 87.100 105.100 89.500 105.300 ;
        RECT 86.200 104.500 88.900 104.800 ;
        RECT 86.200 104.400 86.600 104.500 ;
        RECT 88.500 104.400 88.900 104.500 ;
        RECT 89.200 104.500 89.500 105.100 ;
        RECT 90.200 105.200 90.500 106.800 ;
        RECT 91.000 106.400 91.400 106.500 ;
        RECT 91.000 106.100 92.900 106.400 ;
        RECT 92.500 106.000 92.900 106.100 ;
        RECT 91.700 105.700 92.100 105.800 ;
        RECT 93.400 105.700 93.800 107.400 ;
        RECT 94.600 107.200 95.000 107.400 ;
        RECT 96.600 107.200 96.900 107.900 ;
        RECT 94.200 106.900 95.000 107.200 ;
        RECT 94.200 106.800 94.600 106.900 ;
        RECT 95.700 106.800 97.000 107.200 ;
        RECT 95.000 105.800 95.400 106.600 ;
        RECT 91.700 105.400 93.800 105.700 ;
        RECT 90.200 104.900 91.400 105.200 ;
        RECT 89.900 104.500 90.300 104.600 ;
        RECT 89.200 104.200 90.300 104.500 ;
        RECT 91.100 104.400 91.400 104.900 ;
        RECT 91.100 104.000 91.800 104.400 ;
        RECT 87.900 103.700 88.300 103.800 ;
        RECT 89.300 103.700 89.700 103.800 ;
        RECT 86.200 103.100 86.600 103.500 ;
        RECT 87.900 103.400 89.700 103.700 ;
        RECT 89.000 103.100 89.300 103.400 ;
        RECT 91.000 103.100 91.400 103.500 ;
        RECT 86.200 102.800 87.200 103.100 ;
        RECT 86.800 101.100 87.200 102.800 ;
        RECT 89.000 101.100 89.400 103.100 ;
        RECT 91.100 101.100 91.700 103.100 ;
        RECT 93.400 101.100 93.800 105.400 ;
        RECT 95.700 105.100 96.000 106.800 ;
        RECT 96.600 105.100 97.000 105.200 ;
        RECT 95.500 104.800 96.000 105.100 ;
        RECT 96.300 104.800 97.000 105.100 ;
        RECT 95.500 102.200 95.900 104.800 ;
        RECT 96.300 104.200 96.600 104.800 ;
        RECT 97.400 104.400 97.800 105.200 ;
        RECT 96.200 103.800 96.600 104.200 ;
        RECT 95.000 101.800 95.900 102.200 ;
        RECT 95.500 101.100 95.900 101.800 ;
        RECT 98.200 101.100 98.600 107.900 ;
        RECT 99.000 107.100 99.400 107.600 ;
        RECT 99.800 107.100 100.200 107.200 ;
        RECT 99.000 106.800 100.200 107.100 ;
        RECT 99.000 105.100 99.400 105.200 ;
        RECT 101.400 105.100 101.800 105.200 ;
        RECT 99.000 104.800 101.800 105.100 ;
        RECT 101.400 104.400 101.800 104.800 ;
        RECT 102.200 101.100 102.600 107.900 ;
        RECT 103.000 107.100 103.400 107.600 ;
        RECT 103.800 107.100 104.200 107.200 ;
        RECT 103.000 106.800 104.200 107.100 ;
        RECT 104.600 106.100 105.000 107.900 ;
        RECT 107.000 107.900 107.900 108.200 ;
        RECT 108.900 108.200 109.300 108.800 ;
        RECT 112.300 108.200 112.700 109.900 ;
        RECT 108.900 107.900 109.800 108.200 ;
        RECT 105.400 106.800 105.800 107.600 ;
        RECT 106.200 106.800 106.600 107.600 ;
        RECT 104.600 105.800 105.700 106.100 ;
        RECT 103.800 104.400 104.200 105.200 ;
        RECT 104.600 101.100 105.000 105.800 ;
        RECT 105.400 105.200 105.700 105.800 ;
        RECT 105.400 104.800 105.800 105.200 ;
        RECT 107.000 101.100 107.400 107.900 ;
        RECT 107.800 105.100 108.200 105.200 ;
        RECT 108.600 105.100 109.000 105.200 ;
        RECT 107.800 104.800 109.000 105.100 ;
        RECT 107.800 104.400 108.200 104.800 ;
        RECT 108.600 104.400 109.000 104.800 ;
        RECT 109.400 101.100 109.800 107.900 ;
        RECT 111.800 107.900 112.700 108.200 ;
        RECT 110.200 106.800 110.600 107.600 ;
        RECT 111.000 106.800 111.400 107.600 ;
        RECT 111.000 105.100 111.400 105.200 ;
        RECT 111.800 105.100 112.200 107.900 ;
        RECT 114.200 107.600 114.600 109.900 ;
        RECT 115.800 107.600 116.200 109.900 ;
        RECT 117.400 107.600 117.800 109.900 ;
        RECT 119.000 107.600 119.400 109.900 ;
        RECT 121.900 108.200 122.300 109.900 ;
        RECT 124.300 108.200 124.700 109.900 ;
        RECT 121.400 107.900 122.300 108.200 ;
        RECT 123.800 107.900 124.700 108.200 ;
        RECT 125.400 107.900 125.800 109.900 ;
        RECT 126.200 108.000 126.600 109.900 ;
        RECT 127.800 108.000 128.200 109.900 ;
        RECT 129.900 108.200 130.300 109.900 ;
        RECT 131.300 109.200 131.700 109.900 ;
        RECT 134.700 109.200 135.100 109.900 ;
        RECT 131.000 108.800 131.700 109.200 ;
        RECT 134.200 108.800 135.100 109.200 ;
        RECT 126.200 107.900 128.200 108.000 ;
        RECT 129.400 107.900 130.300 108.200 ;
        RECT 131.300 108.200 131.700 108.800 ;
        RECT 134.700 108.200 135.100 108.800 ;
        RECT 131.300 107.900 132.200 108.200 ;
        RECT 114.200 107.200 115.100 107.600 ;
        RECT 115.800 107.200 116.900 107.600 ;
        RECT 117.400 107.200 118.500 107.600 ;
        RECT 119.000 107.200 120.200 107.600 ;
        RECT 114.700 106.900 115.100 107.200 ;
        RECT 116.500 106.900 116.900 107.200 ;
        RECT 118.100 106.900 118.500 107.200 ;
        RECT 114.700 106.500 116.000 106.900 ;
        RECT 116.500 106.500 117.700 106.900 ;
        RECT 118.100 106.500 119.400 106.900 ;
        RECT 114.700 105.800 115.100 106.500 ;
        RECT 116.500 105.800 116.900 106.500 ;
        RECT 118.100 105.800 118.500 106.500 ;
        RECT 119.800 105.800 120.200 107.200 ;
        RECT 120.600 106.800 121.000 107.600 ;
        RECT 114.200 105.400 115.100 105.800 ;
        RECT 115.800 105.400 116.900 105.800 ;
        RECT 117.400 105.400 118.500 105.800 ;
        RECT 119.000 105.400 120.200 105.800 ;
        RECT 111.000 104.800 112.200 105.100 ;
        RECT 111.800 101.100 112.200 104.800 ;
        RECT 112.600 104.400 113.000 105.200 ;
        RECT 114.200 101.100 114.600 105.400 ;
        RECT 115.800 101.100 116.200 105.400 ;
        RECT 117.400 101.100 117.800 105.400 ;
        RECT 119.000 101.100 119.400 105.400 ;
        RECT 121.400 101.100 121.800 107.900 ;
        RECT 122.200 107.100 122.600 107.200 ;
        RECT 123.000 107.100 123.400 107.600 ;
        RECT 122.200 106.800 123.400 107.100 ;
        RECT 123.800 106.100 124.200 107.900 ;
        RECT 125.500 107.200 125.800 107.900 ;
        RECT 126.300 107.700 128.100 107.900 ;
        RECT 127.400 107.200 127.800 107.400 ;
        RECT 125.400 106.800 126.700 107.200 ;
        RECT 127.400 106.900 128.200 107.200 ;
        RECT 127.800 106.800 128.200 106.900 ;
        RECT 128.600 106.800 129.000 107.600 ;
        RECT 123.800 105.800 125.700 106.100 ;
        RECT 122.200 105.100 122.600 105.200 ;
        RECT 123.000 105.100 123.400 105.200 ;
        RECT 122.200 104.800 123.400 105.100 ;
        RECT 122.200 104.400 122.600 104.800 ;
        RECT 123.800 101.100 124.200 105.800 ;
        RECT 125.400 105.200 125.700 105.800 ;
        RECT 124.600 104.400 125.000 105.200 ;
        RECT 125.400 105.100 125.800 105.200 ;
        RECT 126.400 105.100 126.700 106.800 ;
        RECT 127.000 105.800 127.400 106.600 ;
        RECT 125.400 104.800 126.100 105.100 ;
        RECT 126.400 104.800 126.900 105.100 ;
        RECT 125.800 104.200 126.100 104.800 ;
        RECT 125.800 103.800 126.200 104.200 ;
        RECT 126.500 101.100 126.900 104.800 ;
        RECT 129.400 101.100 129.800 107.900 ;
        RECT 130.200 104.400 130.600 105.200 ;
        RECT 131.000 104.400 131.400 105.200 ;
        RECT 131.800 101.100 132.200 107.900 ;
        RECT 134.200 107.900 135.100 108.200 ;
        RECT 132.600 107.100 133.000 107.600 ;
        RECT 133.400 107.100 133.800 107.600 ;
        RECT 132.600 106.800 133.800 107.100 ;
        RECT 132.600 104.100 133.000 104.200 ;
        RECT 134.200 104.100 134.600 107.900 ;
        RECT 135.800 107.700 136.200 109.900 ;
        RECT 137.900 109.200 138.500 109.900 ;
        RECT 137.900 108.900 138.600 109.200 ;
        RECT 140.200 108.900 140.600 109.900 ;
        RECT 142.400 109.200 142.800 109.900 ;
        RECT 142.400 108.900 143.400 109.200 ;
        RECT 138.200 108.500 138.600 108.900 ;
        RECT 140.300 108.600 140.600 108.900 ;
        RECT 140.300 108.300 141.700 108.600 ;
        RECT 141.300 108.200 141.700 108.300 ;
        RECT 142.200 107.800 142.600 108.600 ;
        RECT 143.000 108.500 143.400 108.900 ;
        RECT 137.300 107.700 137.700 107.800 ;
        RECT 135.800 107.400 137.700 107.700 ;
        RECT 135.800 105.700 136.200 107.400 ;
        RECT 139.300 107.100 139.700 107.200 ;
        RECT 142.200 107.100 142.500 107.800 ;
        RECT 144.600 107.500 145.000 109.900 ;
        RECT 146.200 107.600 146.600 109.900 ;
        RECT 147.800 107.600 148.200 109.900 ;
        RECT 149.400 107.600 149.800 109.900 ;
        RECT 151.000 107.600 151.400 109.900 ;
        RECT 155.500 108.200 155.900 109.900 ;
        RECT 155.000 107.900 155.900 108.200 ;
        RECT 156.600 108.500 157.000 109.500 ;
        RECT 146.200 107.200 147.100 107.600 ;
        RECT 147.800 107.200 148.900 107.600 ;
        RECT 149.400 107.200 150.500 107.600 ;
        RECT 151.000 107.200 152.200 107.600 ;
        RECT 143.800 107.100 144.600 107.200 ;
        RECT 145.400 107.100 145.800 107.200 ;
        RECT 139.100 106.900 145.800 107.100 ;
        RECT 146.700 106.900 147.100 107.200 ;
        RECT 148.500 106.900 148.900 107.200 ;
        RECT 150.100 106.900 150.500 107.200 ;
        RECT 139.100 106.800 146.300 106.900 ;
        RECT 138.200 106.400 138.600 106.500 ;
        RECT 136.700 106.100 138.600 106.400 ;
        RECT 136.700 106.000 137.100 106.100 ;
        RECT 137.500 105.700 137.900 105.800 ;
        RECT 135.800 105.400 137.900 105.700 ;
        RECT 135.000 104.400 135.400 105.200 ;
        RECT 132.600 103.800 134.600 104.100 ;
        RECT 134.200 101.100 134.600 103.800 ;
        RECT 135.800 101.100 136.200 105.400 ;
        RECT 139.100 105.200 139.400 106.800 ;
        RECT 142.700 106.700 143.100 106.800 ;
        RECT 145.400 106.500 146.300 106.800 ;
        RECT 146.700 106.500 148.000 106.900 ;
        RECT 148.500 106.500 149.700 106.900 ;
        RECT 150.100 106.500 151.400 106.900 ;
        RECT 142.200 106.200 142.600 106.300 ;
        RECT 143.500 106.200 143.900 106.300 ;
        RECT 141.400 105.900 143.900 106.200 ;
        RECT 141.400 105.800 141.800 105.900 ;
        RECT 146.700 105.800 147.100 106.500 ;
        RECT 148.500 105.800 148.900 106.500 ;
        RECT 150.100 105.800 150.500 106.500 ;
        RECT 151.800 105.800 152.200 107.200 ;
        RECT 153.400 107.100 153.800 107.200 ;
        RECT 154.200 107.100 154.600 107.600 ;
        RECT 153.400 106.800 154.600 107.100 ;
        RECT 154.200 106.100 154.600 106.200 ;
        RECT 155.000 106.100 155.400 107.900 ;
        RECT 156.600 107.400 156.900 108.500 ;
        RECT 158.700 108.000 159.100 109.500 ;
        RECT 158.700 107.700 159.500 108.000 ;
        RECT 162.700 107.900 163.500 109.900 ;
        RECT 165.700 108.200 166.100 109.900 ;
        RECT 165.700 107.900 166.600 108.200 ;
        RECT 167.800 108.000 168.200 109.900 ;
        RECT 169.400 108.000 169.800 109.900 ;
        RECT 167.800 107.900 169.800 108.000 ;
        RECT 170.200 107.900 170.600 109.900 ;
        RECT 171.100 108.200 171.500 108.600 ;
        RECT 159.100 107.500 159.500 107.700 ;
        RECT 156.600 107.100 158.700 107.400 ;
        RECT 158.200 106.900 158.700 107.100 ;
        RECT 159.200 107.200 159.500 107.500 ;
        RECT 159.200 107.100 160.200 107.200 ;
        RECT 162.200 107.100 162.600 107.200 ;
        RECT 154.200 105.800 155.400 106.100 ;
        RECT 156.600 105.800 157.000 106.600 ;
        RECT 157.400 105.800 157.800 106.600 ;
        RECT 158.200 106.500 158.900 106.900 ;
        RECT 159.200 106.800 162.600 107.100 ;
        RECT 142.200 105.500 145.000 105.600 ;
        RECT 142.100 105.400 145.000 105.500 ;
        RECT 138.200 104.900 139.400 105.200 ;
        RECT 140.100 105.300 145.000 105.400 ;
        RECT 140.100 105.100 142.500 105.300 ;
        RECT 138.200 104.400 138.500 104.900 ;
        RECT 137.800 104.000 138.500 104.400 ;
        RECT 139.300 104.500 139.700 104.600 ;
        RECT 140.100 104.500 140.400 105.100 ;
        RECT 139.300 104.200 140.400 104.500 ;
        RECT 140.700 104.500 143.400 104.800 ;
        RECT 140.700 104.400 141.100 104.500 ;
        RECT 143.000 104.400 143.400 104.500 ;
        RECT 139.900 103.700 140.300 103.800 ;
        RECT 141.300 103.700 141.700 103.800 ;
        RECT 138.200 103.100 138.600 103.500 ;
        RECT 139.900 103.400 141.700 103.700 ;
        RECT 140.300 103.100 140.600 103.400 ;
        RECT 143.000 103.100 143.400 103.500 ;
        RECT 137.900 101.100 138.500 103.100 ;
        RECT 140.200 101.100 140.600 103.100 ;
        RECT 142.400 102.800 143.400 103.100 ;
        RECT 142.400 101.100 142.800 102.800 ;
        RECT 144.600 101.100 145.000 105.300 ;
        RECT 146.200 105.400 147.100 105.800 ;
        RECT 147.800 105.400 148.900 105.800 ;
        RECT 149.400 105.400 150.500 105.800 ;
        RECT 151.000 105.400 152.200 105.800 ;
        RECT 146.200 101.100 146.600 105.400 ;
        RECT 147.800 101.100 148.200 105.400 ;
        RECT 149.400 101.100 149.800 105.400 ;
        RECT 151.000 101.100 151.400 105.400 ;
        RECT 155.000 101.100 155.400 105.800 ;
        RECT 158.200 105.500 158.500 106.500 ;
        RECT 156.600 105.200 158.500 105.500 ;
        RECT 155.800 104.400 156.200 105.200 ;
        RECT 156.600 103.500 156.900 105.200 ;
        RECT 159.200 104.900 159.500 106.800 ;
        RECT 162.300 106.600 162.600 106.800 ;
        RECT 162.300 106.200 162.700 106.600 ;
        RECT 163.000 106.200 163.300 107.900 ;
        RECT 163.800 106.400 164.200 107.200 ;
        RECT 159.800 105.400 160.200 106.200 ;
        RECT 161.400 105.400 161.800 106.200 ;
        RECT 163.000 105.800 163.400 106.200 ;
        RECT 164.600 106.100 165.000 106.200 ;
        RECT 164.200 105.800 165.000 106.100 ;
        RECT 166.200 106.100 166.600 107.900 ;
        RECT 167.900 107.700 169.700 107.900 ;
        RECT 167.000 106.800 167.400 107.600 ;
        RECT 168.200 107.200 168.600 107.400 ;
        RECT 170.200 107.200 170.500 107.900 ;
        RECT 171.000 107.800 171.400 108.200 ;
        RECT 171.800 107.900 172.200 109.900 ;
        RECT 175.500 108.200 175.900 109.900 ;
        RECT 167.800 106.900 168.600 107.200 ;
        RECT 169.300 107.100 170.600 107.200 ;
        RECT 171.000 107.100 171.400 107.200 ;
        RECT 167.800 106.800 168.200 106.900 ;
        RECT 169.300 106.800 171.400 107.100 ;
        RECT 167.800 106.100 168.100 106.800 ;
        RECT 166.200 105.800 168.100 106.100 ;
        RECT 168.600 105.800 169.000 106.600 ;
        RECT 163.000 105.700 163.300 105.800 ;
        RECT 162.300 105.400 163.300 105.700 ;
        RECT 164.200 105.600 164.600 105.800 ;
        RECT 162.300 105.100 162.600 105.400 ;
        RECT 158.700 104.600 159.500 104.900 ;
        RECT 156.600 101.500 157.000 103.500 ;
        RECT 158.700 101.100 159.100 104.600 ;
        RECT 161.400 101.400 161.800 105.100 ;
        RECT 162.200 101.700 162.600 105.100 ;
        RECT 163.000 104.800 165.000 105.100 ;
        RECT 163.000 101.400 163.400 104.800 ;
        RECT 161.400 101.100 163.400 101.400 ;
        RECT 164.600 101.100 165.000 104.800 ;
        RECT 165.400 104.400 165.800 105.200 ;
        RECT 166.200 101.100 166.600 105.800 ;
        RECT 169.300 105.100 169.600 106.800 ;
        RECT 171.000 106.100 171.400 106.200 ;
        RECT 171.900 106.100 172.200 107.900 ;
        RECT 175.000 107.900 175.900 108.200 ;
        RECT 172.600 106.400 173.000 107.200 ;
        RECT 173.400 106.100 173.800 106.200 ;
        RECT 175.000 106.100 175.400 107.900 ;
        RECT 171.000 105.800 172.200 106.100 ;
        RECT 173.000 105.800 175.400 106.100 ;
        RECT 170.200 105.100 170.600 105.200 ;
        RECT 171.100 105.100 171.400 105.800 ;
        RECT 173.000 105.600 173.400 105.800 ;
        RECT 169.100 104.800 169.600 105.100 ;
        RECT 169.900 104.800 170.600 105.100 ;
        RECT 169.100 101.100 169.500 104.800 ;
        RECT 169.900 104.200 170.200 104.800 ;
        RECT 169.800 103.800 170.200 104.200 ;
        RECT 171.000 101.100 171.400 105.100 ;
        RECT 171.800 104.800 173.800 105.100 ;
        RECT 171.800 101.100 172.200 104.800 ;
        RECT 173.400 101.100 173.800 104.800 ;
        RECT 175.000 101.100 175.400 105.800 ;
        RECT 176.600 107.700 177.000 109.900 ;
        RECT 178.700 109.200 179.300 109.900 ;
        RECT 178.700 108.900 179.400 109.200 ;
        RECT 181.000 108.900 181.400 109.900 ;
        RECT 183.200 109.200 183.600 109.900 ;
        RECT 183.200 108.900 184.200 109.200 ;
        RECT 179.000 108.500 179.400 108.900 ;
        RECT 181.100 108.600 181.400 108.900 ;
        RECT 181.100 108.300 182.500 108.600 ;
        RECT 182.100 108.200 182.500 108.300 ;
        RECT 183.000 108.200 183.400 108.600 ;
        RECT 183.800 108.500 184.200 108.900 ;
        RECT 178.100 107.700 178.500 107.800 ;
        RECT 176.600 107.400 178.500 107.700 ;
        RECT 176.600 105.700 177.000 107.400 ;
        RECT 180.100 107.100 180.500 107.200 ;
        RECT 182.200 107.100 182.600 107.200 ;
        RECT 183.000 107.100 183.300 108.200 ;
        RECT 185.400 107.500 185.800 109.900 ;
        RECT 186.200 107.900 186.600 109.900 ;
        RECT 187.000 108.000 187.400 109.900 ;
        RECT 188.600 108.000 189.000 109.900 ;
        RECT 187.000 107.900 189.000 108.000 ;
        RECT 186.300 107.200 186.600 107.900 ;
        RECT 187.100 107.700 188.900 107.900 ;
        RECT 189.400 107.700 189.800 109.900 ;
        RECT 191.500 109.200 192.100 109.900 ;
        RECT 191.500 108.900 192.200 109.200 ;
        RECT 193.800 108.900 194.200 109.900 ;
        RECT 196.000 109.200 196.400 109.900 ;
        RECT 196.000 108.900 197.000 109.200 ;
        RECT 191.800 108.500 192.200 108.900 ;
        RECT 193.900 108.600 194.200 108.900 ;
        RECT 193.900 108.300 195.300 108.600 ;
        RECT 194.900 108.200 195.300 108.300 ;
        RECT 195.800 108.200 196.200 108.600 ;
        RECT 196.600 108.500 197.000 108.900 ;
        RECT 190.900 107.700 191.300 107.800 ;
        RECT 189.400 107.400 191.300 107.700 ;
        RECT 188.200 107.200 188.600 107.400 ;
        RECT 184.600 107.100 185.400 107.200 ;
        RECT 179.900 106.800 185.400 107.100 ;
        RECT 186.200 106.800 187.500 107.200 ;
        RECT 188.200 106.900 189.000 107.200 ;
        RECT 188.600 106.800 189.000 106.900 ;
        RECT 179.000 106.400 179.400 106.500 ;
        RECT 177.500 106.100 179.400 106.400 ;
        RECT 177.500 106.000 177.900 106.100 ;
        RECT 178.300 105.700 178.700 105.800 ;
        RECT 176.600 105.400 178.700 105.700 ;
        RECT 175.800 104.100 176.200 105.200 ;
        RECT 176.600 104.100 177.000 105.400 ;
        RECT 178.200 104.800 178.600 105.400 ;
        RECT 179.900 105.200 180.200 106.800 ;
        RECT 183.500 106.700 183.900 106.800 ;
        RECT 184.300 106.200 184.700 106.300 ;
        RECT 181.400 106.100 181.800 106.200 ;
        RECT 182.200 106.100 184.700 106.200 ;
        RECT 181.400 105.900 184.700 106.100 ;
        RECT 181.400 105.800 182.600 105.900 ;
        RECT 183.000 105.500 185.800 105.600 ;
        RECT 182.900 105.400 185.800 105.500 ;
        RECT 179.000 104.900 180.200 105.200 ;
        RECT 180.900 105.300 185.800 105.400 ;
        RECT 180.900 105.100 183.300 105.300 ;
        RECT 179.000 104.400 179.300 104.900 ;
        RECT 175.800 103.800 177.000 104.100 ;
        RECT 178.600 104.000 179.300 104.400 ;
        RECT 180.100 104.500 180.500 104.600 ;
        RECT 180.900 104.500 181.200 105.100 ;
        RECT 180.100 104.200 181.200 104.500 ;
        RECT 181.500 104.500 184.200 104.800 ;
        RECT 181.500 104.400 181.900 104.500 ;
        RECT 183.800 104.400 184.200 104.500 ;
        RECT 176.600 101.100 177.000 103.800 ;
        RECT 180.700 103.700 181.100 103.800 ;
        RECT 182.100 103.700 182.500 103.800 ;
        RECT 179.000 103.100 179.400 103.500 ;
        RECT 180.700 103.400 182.500 103.700 ;
        RECT 181.100 103.100 181.400 103.400 ;
        RECT 183.800 103.100 184.200 103.500 ;
        RECT 178.700 101.100 179.300 103.100 ;
        RECT 181.000 101.100 181.400 103.100 ;
        RECT 183.200 102.800 184.200 103.100 ;
        RECT 183.200 101.100 183.600 102.800 ;
        RECT 185.400 101.100 185.800 105.300 ;
        RECT 186.200 105.100 186.600 105.200 ;
        RECT 187.200 105.100 187.500 106.800 ;
        RECT 187.800 105.800 188.200 106.600 ;
        RECT 189.400 105.700 189.800 107.400 ;
        RECT 192.900 107.100 193.300 107.200 ;
        RECT 195.800 107.100 196.100 108.200 ;
        RECT 198.200 107.500 198.600 109.900 ;
        RECT 200.300 107.900 201.100 109.900 ;
        RECT 206.500 108.000 206.900 109.500 ;
        RECT 208.600 108.500 209.000 109.500 ;
        RECT 197.400 107.100 198.200 107.200 ;
        RECT 192.700 106.800 198.200 107.100 ;
        RECT 199.800 106.800 200.200 107.200 ;
        RECT 191.800 106.400 192.200 106.500 ;
        RECT 190.300 106.100 192.200 106.400 ;
        RECT 190.300 106.000 190.700 106.100 ;
        RECT 191.100 105.700 191.500 105.800 ;
        RECT 189.400 105.400 191.500 105.700 ;
        RECT 186.200 104.800 186.900 105.100 ;
        RECT 187.200 104.800 187.700 105.100 ;
        RECT 186.600 104.200 186.900 104.800 ;
        RECT 186.600 103.800 187.000 104.200 ;
        RECT 187.300 102.200 187.700 104.800 ;
        RECT 187.300 101.800 188.200 102.200 ;
        RECT 187.300 101.100 187.700 101.800 ;
        RECT 189.400 101.100 189.800 105.400 ;
        RECT 192.700 105.200 193.000 106.800 ;
        RECT 196.300 106.700 196.700 106.800 ;
        RECT 199.900 106.600 200.200 106.800 ;
        RECT 197.100 106.200 197.500 106.300 ;
        RECT 199.900 106.200 200.300 106.600 ;
        RECT 200.600 106.200 200.900 107.900 ;
        RECT 206.100 107.700 206.900 108.000 ;
        RECT 206.100 107.500 206.500 107.700 ;
        RECT 206.100 107.200 206.400 107.500 ;
        RECT 208.700 107.400 209.000 108.500 ;
        RECT 209.400 108.000 209.800 109.900 ;
        RECT 211.000 108.000 211.400 109.900 ;
        RECT 209.400 107.900 211.400 108.000 ;
        RECT 211.800 107.900 212.200 109.900 ;
        RECT 209.500 107.700 211.300 107.900 ;
        RECT 201.400 106.400 201.800 107.200 ;
        RECT 202.200 107.100 202.600 107.200 ;
        RECT 205.400 107.100 206.400 107.200 ;
        RECT 202.200 106.800 206.400 107.100 ;
        RECT 206.900 107.100 209.000 107.400 ;
        RECT 209.800 107.200 210.200 107.400 ;
        RECT 211.800 107.200 212.100 107.900 ;
        RECT 212.600 107.500 213.000 109.900 ;
        RECT 214.800 109.200 215.200 109.900 ;
        RECT 214.200 108.900 215.200 109.200 ;
        RECT 217.000 108.900 217.400 109.900 ;
        RECT 219.100 109.200 219.700 109.900 ;
        RECT 219.000 108.900 219.700 109.200 ;
        RECT 214.200 108.500 214.600 108.900 ;
        RECT 217.000 108.600 217.300 108.900 ;
        RECT 215.000 107.800 215.400 108.600 ;
        RECT 215.900 108.300 217.300 108.600 ;
        RECT 219.000 108.500 219.400 108.900 ;
        RECT 215.900 108.200 216.300 108.300 ;
        RECT 206.900 106.900 207.400 107.100 ;
        RECT 194.200 106.100 194.600 106.200 ;
        RECT 195.000 106.100 197.500 106.200 ;
        RECT 194.200 105.900 197.500 106.100 ;
        RECT 194.200 105.800 195.400 105.900 ;
        RECT 195.800 105.500 198.600 105.600 ;
        RECT 195.700 105.400 198.600 105.500 ;
        RECT 199.000 105.400 199.400 106.200 ;
        RECT 200.600 105.800 201.000 106.200 ;
        RECT 202.200 106.100 202.600 106.200 ;
        RECT 203.000 106.100 203.400 106.200 ;
        RECT 201.800 105.800 203.400 106.100 ;
        RECT 200.600 105.700 200.900 105.800 ;
        RECT 199.900 105.400 200.900 105.700 ;
        RECT 201.800 105.600 202.200 105.800 ;
        RECT 205.400 105.400 205.800 106.200 ;
        RECT 191.800 104.900 193.000 105.200 ;
        RECT 193.700 105.300 198.600 105.400 ;
        RECT 193.700 105.100 196.100 105.300 ;
        RECT 191.800 104.400 192.100 104.900 ;
        RECT 191.400 104.000 192.100 104.400 ;
        RECT 192.900 104.500 193.300 104.600 ;
        RECT 193.700 104.500 194.000 105.100 ;
        RECT 192.900 104.200 194.000 104.500 ;
        RECT 194.300 104.500 197.000 104.800 ;
        RECT 194.300 104.400 194.700 104.500 ;
        RECT 196.600 104.400 197.000 104.500 ;
        RECT 193.500 103.700 193.900 103.800 ;
        RECT 194.900 103.700 195.300 103.800 ;
        RECT 191.800 103.100 192.200 103.500 ;
        RECT 193.500 103.400 195.300 103.700 ;
        RECT 193.900 103.100 194.200 103.400 ;
        RECT 196.600 103.100 197.000 103.500 ;
        RECT 191.500 101.100 192.100 103.100 ;
        RECT 193.800 101.100 194.200 103.100 ;
        RECT 196.000 102.800 197.000 103.100 ;
        RECT 196.000 101.100 196.400 102.800 ;
        RECT 198.200 101.100 198.600 105.300 ;
        RECT 199.900 105.100 200.200 105.400 ;
        RECT 199.000 101.400 199.400 105.100 ;
        RECT 199.800 101.700 200.200 105.100 ;
        RECT 200.600 104.800 202.600 105.100 ;
        RECT 200.600 101.400 201.000 104.800 ;
        RECT 199.000 101.100 201.000 101.400 ;
        RECT 202.200 101.100 202.600 104.800 ;
        RECT 206.100 104.900 206.400 106.800 ;
        RECT 206.700 106.500 207.400 106.900 ;
        RECT 209.400 106.900 210.200 107.200 ;
        RECT 209.400 106.800 209.800 106.900 ;
        RECT 210.900 106.800 212.200 107.200 ;
        RECT 213.000 107.100 213.800 107.200 ;
        RECT 215.100 107.100 215.400 107.800 ;
        RECT 219.900 107.700 220.300 107.800 ;
        RECT 221.400 107.700 221.800 109.900 ;
        RECT 222.500 109.200 222.900 109.900 ;
        RECT 222.200 108.800 222.900 109.200 ;
        RECT 222.500 108.200 222.900 108.800 ;
        RECT 224.600 108.500 225.000 109.500 ;
        RECT 222.500 107.900 223.400 108.200 ;
        RECT 219.900 107.400 221.800 107.700 ;
        RECT 217.900 107.100 218.300 107.200 ;
        RECT 213.000 106.800 218.500 107.100 ;
        RECT 207.100 105.500 207.400 106.500 ;
        RECT 207.800 105.800 208.200 106.600 ;
        RECT 208.600 105.800 209.000 106.600 ;
        RECT 210.200 105.800 210.600 106.600 ;
        RECT 207.100 105.200 209.000 105.500 ;
        RECT 206.100 104.600 206.900 104.900 ;
        RECT 206.500 101.100 206.900 104.600 ;
        RECT 208.700 103.500 209.000 105.200 ;
        RECT 210.900 105.100 211.200 106.800 ;
        RECT 214.500 106.700 214.900 106.800 ;
        RECT 213.700 106.200 214.100 106.300 ;
        RECT 215.000 106.200 215.400 106.300 ;
        RECT 213.700 105.900 216.200 106.200 ;
        RECT 215.800 105.800 216.200 105.900 ;
        RECT 212.600 105.500 215.400 105.600 ;
        RECT 212.600 105.400 215.500 105.500 ;
        RECT 212.600 105.300 217.500 105.400 ;
        RECT 211.800 105.100 212.200 105.200 ;
        RECT 208.600 101.500 209.000 103.500 ;
        RECT 210.700 104.800 211.200 105.100 ;
        RECT 211.500 104.800 212.200 105.100 ;
        RECT 210.700 101.100 211.100 104.800 ;
        RECT 211.500 104.200 211.800 104.800 ;
        RECT 211.400 103.800 211.800 104.200 ;
        RECT 212.600 101.100 213.000 105.300 ;
        RECT 215.100 105.100 217.500 105.300 ;
        RECT 214.200 104.500 216.900 104.800 ;
        RECT 214.200 104.400 214.600 104.500 ;
        RECT 216.500 104.400 216.900 104.500 ;
        RECT 217.200 104.500 217.500 105.100 ;
        RECT 218.200 105.200 218.500 106.800 ;
        RECT 219.000 106.400 219.400 106.500 ;
        RECT 219.000 106.100 220.900 106.400 ;
        RECT 220.500 106.000 220.900 106.100 ;
        RECT 219.700 105.700 220.100 105.800 ;
        RECT 221.400 105.700 221.800 107.400 ;
        RECT 219.700 105.400 221.800 105.700 ;
        RECT 218.200 104.900 219.400 105.200 ;
        RECT 217.900 104.500 218.300 104.600 ;
        RECT 217.200 104.200 218.300 104.500 ;
        RECT 219.100 104.400 219.400 104.900 ;
        RECT 219.100 104.200 219.800 104.400 ;
        RECT 219.100 104.000 220.200 104.200 ;
        RECT 219.500 103.800 220.200 104.000 ;
        RECT 215.900 103.700 216.300 103.800 ;
        RECT 217.300 103.700 217.700 103.800 ;
        RECT 214.200 103.100 214.600 103.500 ;
        RECT 215.900 103.400 217.700 103.700 ;
        RECT 217.000 103.100 217.300 103.400 ;
        RECT 219.000 103.100 219.400 103.500 ;
        RECT 214.200 102.800 215.200 103.100 ;
        RECT 214.800 101.100 215.200 102.800 ;
        RECT 217.000 101.100 217.400 103.100 ;
        RECT 219.100 101.100 219.700 103.100 ;
        RECT 221.400 101.100 221.800 105.400 ;
        RECT 222.200 104.400 222.600 105.200 ;
        RECT 223.000 101.100 223.400 107.900 ;
        RECT 223.800 106.800 224.200 107.600 ;
        RECT 224.600 107.400 224.900 108.500 ;
        RECT 226.700 108.000 227.100 109.500 ;
        RECT 226.700 107.700 227.500 108.000 ;
        RECT 227.100 107.500 227.500 107.700 ;
        RECT 224.600 107.100 226.700 107.400 ;
        RECT 226.200 106.900 226.700 107.100 ;
        RECT 227.200 107.200 227.500 107.500 ;
        RECT 229.400 107.600 229.800 109.900 ;
        RECT 232.600 107.600 233.000 109.900 ;
        RECT 234.200 107.600 234.600 109.900 ;
        RECT 235.800 107.600 236.200 109.900 ;
        RECT 237.400 107.600 237.800 109.900 ;
        RECT 240.300 108.200 240.700 109.900 ;
        RECT 239.800 107.900 240.700 108.200 ;
        RECT 241.400 107.900 241.800 109.900 ;
        RECT 242.200 108.000 242.600 109.900 ;
        RECT 243.800 108.000 244.200 109.900 ;
        RECT 242.200 107.900 244.200 108.000 ;
        RECT 229.400 107.300 230.500 107.600 ;
        RECT 223.800 106.200 224.100 106.800 ;
        RECT 223.800 105.800 224.200 106.200 ;
        RECT 224.600 105.800 225.000 106.600 ;
        RECT 225.400 105.800 225.800 106.600 ;
        RECT 226.200 106.500 226.900 106.900 ;
        RECT 227.200 106.800 228.200 107.200 ;
        RECT 226.200 105.500 226.500 106.500 ;
        RECT 224.600 105.200 226.500 105.500 ;
        RECT 227.200 105.200 227.500 106.800 ;
        RECT 227.800 105.400 228.200 106.200 ;
        RECT 229.400 105.800 229.800 106.600 ;
        RECT 230.200 105.800 230.500 107.300 ;
        RECT 232.600 107.200 233.500 107.600 ;
        RECT 234.200 107.200 235.300 107.600 ;
        RECT 235.800 107.200 236.900 107.600 ;
        RECT 237.400 107.200 238.600 107.600 ;
        RECT 231.800 106.900 232.200 107.200 ;
        RECT 233.100 106.900 233.500 107.200 ;
        RECT 234.900 106.900 235.300 107.200 ;
        RECT 236.500 106.900 236.900 107.200 ;
        RECT 231.800 106.500 232.700 106.900 ;
        RECT 233.100 106.500 234.400 106.900 ;
        RECT 234.900 106.500 236.100 106.900 ;
        RECT 236.500 106.500 237.800 106.900 ;
        RECT 233.100 105.800 233.500 106.500 ;
        RECT 234.900 105.800 235.300 106.500 ;
        RECT 236.500 105.800 236.900 106.500 ;
        RECT 238.200 105.800 238.600 107.200 ;
        RECT 239.000 106.800 239.400 107.600 ;
        RECT 239.000 106.200 239.300 106.800 ;
        RECT 239.000 105.800 239.400 106.200 ;
        RECT 239.800 106.100 240.200 107.900 ;
        RECT 241.500 107.200 241.800 107.900 ;
        RECT 242.300 107.700 244.100 107.900 ;
        RECT 245.400 107.600 245.800 109.900 ;
        RECT 247.000 107.600 247.400 109.900 ;
        RECT 248.600 107.600 249.000 109.900 ;
        RECT 250.200 107.600 250.600 109.900 ;
        RECT 243.400 107.200 243.800 107.400 ;
        RECT 245.400 107.200 246.300 107.600 ;
        RECT 247.000 107.200 248.100 107.600 ;
        RECT 248.600 107.200 249.700 107.600 ;
        RECT 250.200 107.200 251.400 107.600 ;
        RECT 241.400 106.800 242.700 107.200 ;
        RECT 243.400 106.900 244.200 107.200 ;
        RECT 243.800 106.800 244.200 106.900 ;
        RECT 245.900 106.900 246.300 107.200 ;
        RECT 247.700 106.900 248.100 107.200 ;
        RECT 249.300 106.900 249.700 107.200 ;
        RECT 239.800 105.800 241.700 106.100 ;
        RECT 230.200 105.400 230.800 105.800 ;
        RECT 232.600 105.400 233.500 105.800 ;
        RECT 234.200 105.400 235.300 105.800 ;
        RECT 235.800 105.400 236.900 105.800 ;
        RECT 237.400 105.400 238.600 105.800 ;
        RECT 224.600 103.500 224.900 105.200 ;
        RECT 227.000 104.900 227.500 105.200 ;
        RECT 230.200 105.100 230.500 105.400 ;
        RECT 226.700 104.600 227.500 104.900 ;
        RECT 229.400 104.800 230.500 105.100 ;
        RECT 224.600 101.500 225.000 103.500 ;
        RECT 226.700 101.100 227.100 104.600 ;
        RECT 229.400 101.100 229.800 104.800 ;
        RECT 232.600 101.100 233.000 105.400 ;
        RECT 234.200 101.100 234.600 105.400 ;
        RECT 235.800 101.100 236.200 105.400 ;
        RECT 237.400 101.100 237.800 105.400 ;
        RECT 239.800 101.100 240.200 105.800 ;
        RECT 241.400 105.200 241.700 105.800 ;
        RECT 240.600 104.400 241.000 105.200 ;
        RECT 241.400 105.100 241.800 105.200 ;
        RECT 242.400 105.100 242.700 106.800 ;
        RECT 243.000 105.800 243.400 106.600 ;
        RECT 245.900 106.500 247.200 106.900 ;
        RECT 247.700 106.500 248.900 106.900 ;
        RECT 249.300 106.500 250.600 106.900 ;
        RECT 245.900 105.800 246.300 106.500 ;
        RECT 247.700 105.800 248.100 106.500 ;
        RECT 249.300 105.800 249.700 106.500 ;
        RECT 251.000 105.800 251.400 107.200 ;
        RECT 245.400 105.400 246.300 105.800 ;
        RECT 247.000 105.400 248.100 105.800 ;
        RECT 248.600 105.400 249.700 105.800 ;
        RECT 250.200 105.400 251.400 105.800 ;
        RECT 241.400 104.800 242.100 105.100 ;
        RECT 242.400 104.800 242.900 105.100 ;
        RECT 241.800 104.200 242.100 104.800 ;
        RECT 241.800 103.800 242.200 104.200 ;
        RECT 242.500 101.100 242.900 104.800 ;
        RECT 245.400 101.100 245.800 105.400 ;
        RECT 247.000 101.100 247.400 105.400 ;
        RECT 248.600 101.100 249.000 105.400 ;
        RECT 250.200 101.100 250.600 105.400 ;
        RECT 1.700 99.200 2.100 99.900 ;
        RECT 1.700 98.800 2.600 99.200 ;
        RECT 1.000 96.800 1.400 97.200 ;
        RECT 1.000 96.200 1.300 96.800 ;
        RECT 1.700 96.200 2.100 98.800 ;
        RECT 0.600 95.900 1.300 96.200 ;
        RECT 1.600 95.900 2.100 96.200 ;
        RECT 0.600 95.800 1.000 95.900 ;
        RECT 1.600 94.200 1.900 95.900 ;
        RECT 3.800 95.700 4.200 99.900 ;
        RECT 6.000 98.200 6.400 99.900 ;
        RECT 5.400 97.900 6.400 98.200 ;
        RECT 8.200 97.900 8.600 99.900 ;
        RECT 10.300 97.900 10.900 99.900 ;
        RECT 5.400 97.500 5.800 97.900 ;
        RECT 8.200 97.600 8.500 97.900 ;
        RECT 7.100 97.300 8.900 97.600 ;
        RECT 10.200 97.500 10.600 97.900 ;
        RECT 7.100 97.200 7.500 97.300 ;
        RECT 8.500 97.200 8.900 97.300 ;
        RECT 5.400 96.500 5.800 96.600 ;
        RECT 7.700 96.500 8.100 96.600 ;
        RECT 5.400 96.200 8.100 96.500 ;
        RECT 8.400 96.500 9.500 96.800 ;
        RECT 8.400 95.900 8.700 96.500 ;
        RECT 9.100 96.400 9.500 96.500 ;
        RECT 10.300 96.600 11.000 97.000 ;
        RECT 10.300 96.100 10.600 96.600 ;
        RECT 6.300 95.700 8.700 95.900 ;
        RECT 3.800 95.600 8.700 95.700 ;
        RECT 9.400 95.800 10.600 96.100 ;
        RECT 3.800 95.500 6.700 95.600 ;
        RECT 3.800 95.400 6.600 95.500 ;
        RECT 2.200 94.400 2.600 95.200 ;
        RECT 7.000 95.100 7.400 95.200 ;
        RECT 4.900 94.800 7.400 95.100 ;
        RECT 4.900 94.700 5.300 94.800 ;
        RECT 5.700 94.200 6.100 94.300 ;
        RECT 9.400 94.200 9.700 95.800 ;
        RECT 12.600 95.600 13.000 99.900 ;
        RECT 15.300 96.400 15.700 99.900 ;
        RECT 17.400 97.500 17.800 99.500 ;
        RECT 14.900 96.100 15.700 96.400 ;
        RECT 10.900 95.300 13.000 95.600 ;
        RECT 10.900 95.200 11.300 95.300 ;
        RECT 11.700 94.900 12.100 95.000 ;
        RECT 10.200 94.600 12.100 94.900 ;
        RECT 10.200 94.500 10.600 94.600 ;
        RECT 0.600 93.800 1.900 94.200 ;
        RECT 3.000 94.100 3.400 94.200 ;
        RECT 2.600 93.800 3.400 94.100 ;
        RECT 4.200 93.900 9.700 94.200 ;
        RECT 4.200 93.800 5.000 93.900 ;
        RECT 0.700 93.100 1.000 93.800 ;
        RECT 2.600 93.600 3.000 93.800 ;
        RECT 1.500 93.100 3.300 93.300 ;
        RECT 0.600 91.100 1.000 93.100 ;
        RECT 1.400 93.000 3.400 93.100 ;
        RECT 1.400 91.100 1.800 93.000 ;
        RECT 3.000 91.100 3.400 93.000 ;
        RECT 3.800 91.100 4.200 93.500 ;
        RECT 6.300 93.200 6.600 93.900 ;
        RECT 9.100 93.800 9.500 93.900 ;
        RECT 12.600 93.600 13.000 95.300 ;
        RECT 13.400 95.100 13.800 95.200 ;
        RECT 14.200 95.100 14.600 95.600 ;
        RECT 13.400 94.800 14.600 95.100 ;
        RECT 14.900 94.200 15.200 96.100 ;
        RECT 17.500 95.800 17.800 97.500 ;
        RECT 15.900 95.500 17.800 95.800 ;
        RECT 15.900 94.500 16.200 95.500 ;
        RECT 14.200 93.800 15.200 94.200 ;
        RECT 15.500 94.100 16.200 94.500 ;
        RECT 16.600 94.400 17.000 95.200 ;
        RECT 17.400 94.400 17.800 95.200 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 19.000 95.100 19.400 99.900 ;
        RECT 21.000 96.800 21.400 97.200 ;
        RECT 19.800 95.800 20.200 96.600 ;
        RECT 21.000 96.200 21.300 96.800 ;
        RECT 21.700 96.200 22.100 99.900 ;
        RECT 20.600 95.900 21.300 96.200 ;
        RECT 21.600 95.900 22.100 96.200 ;
        RECT 20.600 95.800 21.000 95.900 ;
        RECT 20.600 95.100 20.900 95.800 ;
        RECT 19.000 94.800 20.900 95.100 ;
        RECT 11.100 93.300 13.000 93.600 ;
        RECT 11.100 93.200 11.500 93.300 ;
        RECT 5.400 92.100 5.800 92.500 ;
        RECT 6.200 92.400 6.600 93.200 ;
        RECT 7.100 92.700 7.500 92.800 ;
        RECT 7.100 92.400 8.500 92.700 ;
        RECT 8.200 92.100 8.500 92.400 ;
        RECT 10.200 92.100 10.600 92.500 ;
        RECT 5.400 91.800 6.400 92.100 ;
        RECT 6.000 91.100 6.400 91.800 ;
        RECT 8.200 91.100 8.600 92.100 ;
        RECT 10.200 91.800 10.900 92.100 ;
        RECT 10.300 91.100 10.900 91.800 ;
        RECT 12.600 91.100 13.000 93.300 ;
        RECT 14.900 93.500 15.200 93.800 ;
        RECT 15.700 93.900 16.200 94.100 ;
        RECT 18.200 94.200 18.500 94.800 ;
        RECT 15.700 93.600 17.800 93.900 ;
        RECT 14.900 93.300 15.300 93.500 ;
        RECT 14.900 93.200 15.700 93.300 ;
        RECT 14.900 93.000 16.200 93.200 ;
        RECT 15.300 92.800 16.200 93.000 ;
        RECT 15.300 91.500 15.700 92.800 ;
        RECT 17.500 92.500 17.800 93.600 ;
        RECT 18.200 93.400 18.600 94.200 ;
        RECT 19.000 93.100 19.400 94.800 ;
        RECT 21.600 94.200 21.900 95.900 ;
        RECT 22.200 94.400 22.600 95.200 ;
        RECT 24.600 95.100 25.000 99.900 ;
        RECT 26.600 96.800 27.000 97.200 ;
        RECT 25.400 95.800 25.800 96.600 ;
        RECT 26.600 96.200 26.900 96.800 ;
        RECT 27.300 96.200 27.700 99.900 ;
        RECT 26.200 95.900 26.900 96.200 ;
        RECT 27.200 95.900 27.700 96.200 ;
        RECT 30.700 96.200 31.100 99.900 ;
        RECT 31.400 96.800 31.800 97.200 ;
        RECT 31.500 96.200 31.800 96.800 ;
        RECT 30.700 95.900 31.200 96.200 ;
        RECT 31.500 95.900 32.200 96.200 ;
        RECT 26.200 95.800 26.600 95.900 ;
        RECT 26.200 95.100 26.500 95.800 ;
        RECT 24.600 94.800 26.500 95.100 ;
        RECT 19.800 94.100 20.200 94.200 ;
        RECT 20.600 94.100 21.900 94.200 ;
        RECT 23.000 94.100 23.400 94.200 ;
        RECT 19.800 93.800 21.900 94.100 ;
        RECT 22.600 93.800 23.400 94.100 ;
        RECT 20.700 93.100 21.000 93.800 ;
        RECT 22.600 93.600 23.000 93.800 ;
        RECT 23.800 93.400 24.200 94.200 ;
        RECT 21.500 93.100 23.300 93.300 ;
        RECT 24.600 93.100 25.000 94.800 ;
        RECT 27.200 94.200 27.500 95.900 ;
        RECT 27.800 94.400 28.200 95.200 ;
        RECT 30.200 94.400 30.600 95.200 ;
        RECT 30.900 94.200 31.200 95.900 ;
        RECT 31.800 95.800 32.200 95.900 ;
        RECT 32.600 95.700 33.000 99.900 ;
        RECT 34.800 98.200 35.200 99.900 ;
        RECT 34.200 97.900 35.200 98.200 ;
        RECT 37.000 97.900 37.400 99.900 ;
        RECT 39.100 97.900 39.700 99.900 ;
        RECT 34.200 97.500 34.600 97.900 ;
        RECT 37.000 97.600 37.300 97.900 ;
        RECT 35.900 97.300 37.700 97.600 ;
        RECT 39.000 97.500 39.400 97.900 ;
        RECT 35.900 97.200 36.300 97.300 ;
        RECT 37.300 97.200 37.700 97.300 ;
        RECT 34.200 96.500 34.600 96.600 ;
        RECT 36.500 96.500 36.900 96.600 ;
        RECT 34.200 96.200 36.900 96.500 ;
        RECT 37.200 96.500 38.300 96.800 ;
        RECT 37.200 95.900 37.500 96.500 ;
        RECT 37.900 96.400 38.300 96.500 ;
        RECT 39.100 96.600 39.800 97.000 ;
        RECT 39.100 96.100 39.400 96.600 ;
        RECT 35.100 95.700 37.500 95.900 ;
        RECT 32.600 95.600 37.500 95.700 ;
        RECT 38.200 95.800 39.400 96.100 ;
        RECT 32.600 95.500 35.500 95.600 ;
        RECT 32.600 95.400 35.400 95.500 ;
        RECT 35.800 95.100 36.200 95.200 ;
        RECT 33.700 94.800 36.200 95.100 ;
        RECT 33.700 94.700 34.100 94.800 ;
        RECT 35.000 94.700 35.400 94.800 ;
        RECT 34.500 94.200 34.900 94.300 ;
        RECT 38.200 94.200 38.500 95.800 ;
        RECT 41.400 95.600 41.800 99.900 ;
        RECT 42.600 96.800 43.000 97.200 ;
        RECT 42.600 96.200 42.900 96.800 ;
        RECT 43.300 96.200 43.700 99.900 ;
        RECT 42.200 95.900 42.900 96.200 ;
        RECT 43.200 95.900 43.700 96.200 ;
        RECT 45.400 97.500 45.800 99.500 ;
        RECT 47.500 99.200 47.900 99.900 ;
        RECT 47.500 98.800 48.200 99.200 ;
        RECT 42.200 95.800 42.600 95.900 ;
        RECT 39.700 95.300 41.800 95.600 ;
        RECT 39.700 95.200 40.100 95.300 ;
        RECT 40.500 94.900 40.900 95.000 ;
        RECT 39.000 94.600 40.900 94.900 ;
        RECT 39.000 94.500 39.400 94.600 ;
        RECT 26.200 93.800 27.500 94.200 ;
        RECT 28.600 94.100 29.000 94.200 ;
        RECT 29.400 94.100 29.800 94.200 ;
        RECT 28.200 93.800 30.200 94.100 ;
        RECT 30.900 93.800 32.200 94.200 ;
        RECT 33.000 93.900 38.500 94.200 ;
        RECT 33.000 93.800 33.800 93.900 ;
        RECT 26.300 93.100 26.600 93.800 ;
        RECT 28.200 93.600 28.600 93.800 ;
        RECT 29.800 93.600 30.200 93.800 ;
        RECT 27.100 93.100 28.900 93.300 ;
        RECT 29.500 93.100 31.300 93.300 ;
        RECT 31.800 93.100 32.100 93.800 ;
        RECT 19.000 92.800 19.900 93.100 ;
        RECT 17.400 91.500 17.800 92.500 ;
        RECT 19.500 91.100 19.900 92.800 ;
        RECT 20.600 91.100 21.000 93.100 ;
        RECT 21.400 93.000 23.400 93.100 ;
        RECT 21.400 91.100 21.800 93.000 ;
        RECT 23.000 91.100 23.400 93.000 ;
        RECT 24.600 92.800 25.500 93.100 ;
        RECT 25.100 91.100 25.500 92.800 ;
        RECT 26.200 91.100 26.600 93.100 ;
        RECT 27.000 93.000 29.000 93.100 ;
        RECT 27.000 91.100 27.400 93.000 ;
        RECT 28.600 91.100 29.000 93.000 ;
        RECT 29.400 93.000 31.400 93.100 ;
        RECT 29.400 91.100 29.800 93.000 ;
        RECT 31.000 91.100 31.400 93.000 ;
        RECT 31.800 91.100 32.200 93.100 ;
        RECT 32.600 91.100 33.000 93.500 ;
        RECT 35.100 93.200 35.400 93.900 ;
        RECT 37.900 93.800 38.500 93.900 ;
        RECT 34.200 92.100 34.600 92.500 ;
        RECT 35.000 92.400 35.400 93.200 ;
        RECT 38.200 93.200 38.500 93.800 ;
        RECT 41.400 93.600 41.800 95.300 ;
        RECT 43.200 94.200 43.500 95.900 ;
        RECT 45.400 95.800 45.700 97.500 ;
        RECT 47.500 96.400 47.900 98.800 ;
        RECT 47.500 96.100 48.300 96.400 ;
        RECT 45.400 95.500 47.300 95.800 ;
        RECT 43.800 94.400 44.200 95.200 ;
        RECT 45.400 94.400 45.800 95.200 ;
        RECT 46.200 94.400 46.600 95.200 ;
        RECT 47.000 94.500 47.300 95.500 ;
        RECT 42.200 93.800 43.500 94.200 ;
        RECT 44.600 94.100 45.000 94.200 ;
        RECT 44.200 93.800 45.000 94.100 ;
        RECT 47.000 94.100 47.700 94.500 ;
        RECT 48.000 94.200 48.300 96.100 ;
        RECT 51.800 95.700 52.200 99.900 ;
        RECT 54.000 98.200 54.400 99.900 ;
        RECT 53.400 97.900 54.400 98.200 ;
        RECT 56.200 97.900 56.600 99.900 ;
        RECT 58.300 97.900 58.900 99.900 ;
        RECT 53.400 97.500 53.800 97.900 ;
        RECT 56.200 97.600 56.500 97.900 ;
        RECT 55.100 97.300 56.900 97.600 ;
        RECT 58.200 97.500 58.600 97.900 ;
        RECT 55.100 97.200 55.500 97.300 ;
        RECT 56.500 97.200 56.900 97.300 ;
        RECT 53.400 96.500 53.800 96.600 ;
        RECT 55.700 96.500 56.100 96.600 ;
        RECT 53.400 96.200 56.100 96.500 ;
        RECT 56.400 96.500 57.500 96.800 ;
        RECT 56.400 95.900 56.700 96.500 ;
        RECT 57.100 96.400 57.500 96.500 ;
        RECT 58.300 96.600 59.000 97.000 ;
        RECT 58.300 96.100 58.600 96.600 ;
        RECT 54.300 95.700 56.700 95.900 ;
        RECT 51.800 95.600 56.700 95.700 ;
        RECT 57.400 95.800 58.600 96.100 ;
        RECT 48.600 95.100 49.000 95.600 ;
        RECT 51.800 95.500 54.700 95.600 ;
        RECT 51.800 95.400 54.600 95.500 ;
        RECT 51.000 95.100 51.400 95.200 ;
        RECT 55.000 95.100 55.400 95.200 ;
        RECT 48.600 94.800 51.400 95.100 ;
        RECT 52.900 94.800 55.400 95.100 ;
        RECT 52.900 94.700 53.300 94.800 ;
        RECT 53.700 94.200 54.100 94.300 ;
        RECT 57.400 94.200 57.700 95.800 ;
        RECT 60.600 95.600 61.000 99.900 ;
        RECT 58.900 95.300 61.000 95.600 ;
        RECT 61.400 97.500 61.800 99.500 ;
        RECT 61.400 95.800 61.700 97.500 ;
        RECT 63.500 96.400 63.900 99.900 ;
        RECT 63.500 96.100 64.300 96.400 ;
        RECT 61.400 95.500 63.300 95.800 ;
        RECT 58.900 95.200 59.300 95.300 ;
        RECT 59.700 94.900 60.100 95.000 ;
        RECT 58.200 94.600 60.100 94.900 ;
        RECT 58.200 94.500 58.600 94.600 ;
        RECT 47.000 93.900 47.500 94.100 ;
        RECT 39.900 93.300 41.800 93.600 ;
        RECT 39.900 93.200 40.300 93.300 ;
        RECT 38.200 92.800 38.600 93.200 ;
        RECT 35.900 92.700 36.300 92.800 ;
        RECT 35.900 92.400 37.300 92.700 ;
        RECT 37.000 92.100 37.300 92.400 ;
        RECT 39.000 92.100 39.400 92.500 ;
        RECT 34.200 91.800 35.200 92.100 ;
        RECT 34.800 91.100 35.200 91.800 ;
        RECT 37.000 91.100 37.400 92.100 ;
        RECT 39.000 91.800 39.700 92.100 ;
        RECT 39.100 91.100 39.700 91.800 ;
        RECT 41.400 91.100 41.800 93.300 ;
        RECT 42.300 93.100 42.600 93.800 ;
        RECT 44.200 93.600 44.600 93.800 ;
        RECT 45.400 93.600 47.500 93.900 ;
        RECT 48.000 93.800 49.000 94.200 ;
        RECT 52.200 93.900 57.700 94.200 ;
        RECT 52.200 93.800 53.000 93.900 ;
        RECT 43.100 93.100 44.900 93.300 ;
        RECT 42.200 91.100 42.600 93.100 ;
        RECT 43.000 93.000 45.000 93.100 ;
        RECT 43.000 91.100 43.400 93.000 ;
        RECT 44.600 91.100 45.000 93.000 ;
        RECT 45.400 92.500 45.700 93.600 ;
        RECT 48.000 93.500 48.300 93.800 ;
        RECT 47.900 93.300 48.300 93.500 ;
        RECT 47.500 93.000 48.300 93.300 ;
        RECT 45.400 91.500 45.800 92.500 ;
        RECT 47.500 91.500 47.900 93.000 ;
        RECT 51.800 91.100 52.200 93.500 ;
        RECT 54.300 92.800 54.600 93.900 ;
        RECT 57.100 93.800 57.500 93.900 ;
        RECT 60.600 93.600 61.000 95.300 ;
        RECT 61.400 94.400 61.800 95.200 ;
        RECT 62.200 94.400 62.600 95.200 ;
        RECT 63.000 94.500 63.300 95.500 ;
        RECT 63.000 94.100 63.700 94.500 ;
        RECT 64.000 94.200 64.300 96.100 ;
        RECT 64.600 94.800 65.000 95.600 ;
        RECT 67.000 95.100 67.400 99.900 ;
        RECT 69.000 96.800 69.400 97.200 ;
        RECT 67.800 95.800 68.200 96.600 ;
        RECT 69.000 96.200 69.300 96.800 ;
        RECT 69.700 96.200 70.100 99.900 ;
        RECT 68.600 95.900 69.300 96.200 ;
        RECT 69.600 95.900 70.100 96.200 ;
        RECT 73.100 96.200 73.500 99.900 ;
        RECT 73.800 96.800 74.200 97.200 ;
        RECT 73.900 96.200 74.200 96.800 ;
        RECT 73.100 95.900 73.600 96.200 ;
        RECT 73.900 95.900 74.600 96.200 ;
        RECT 68.600 95.800 69.000 95.900 ;
        RECT 68.600 95.100 68.900 95.800 ;
        RECT 67.000 94.800 68.900 95.100 ;
        RECT 63.000 93.900 63.500 94.100 ;
        RECT 59.100 93.300 61.000 93.600 ;
        RECT 59.100 93.200 59.500 93.300 ;
        RECT 53.400 92.100 53.800 92.500 ;
        RECT 54.200 92.400 54.600 92.800 ;
        RECT 55.100 92.700 55.500 92.800 ;
        RECT 55.100 92.400 56.500 92.700 ;
        RECT 56.200 92.100 56.500 92.400 ;
        RECT 58.200 92.100 58.600 92.500 ;
        RECT 53.400 91.800 54.400 92.100 ;
        RECT 54.000 91.100 54.400 91.800 ;
        RECT 56.200 91.100 56.600 92.100 ;
        RECT 58.200 91.800 58.900 92.100 ;
        RECT 58.300 91.100 58.900 91.800 ;
        RECT 60.600 91.100 61.000 93.300 ;
        RECT 61.400 93.600 63.500 93.900 ;
        RECT 64.000 93.800 65.000 94.200 ;
        RECT 65.400 94.100 65.800 94.200 ;
        RECT 66.200 94.100 66.600 94.200 ;
        RECT 65.400 93.800 66.600 94.100 ;
        RECT 61.400 92.500 61.700 93.600 ;
        RECT 64.000 93.500 64.300 93.800 ;
        RECT 63.900 93.300 64.300 93.500 ;
        RECT 66.200 93.400 66.600 93.800 ;
        RECT 63.500 93.000 64.300 93.300 ;
        RECT 67.000 93.100 67.400 94.800 ;
        RECT 69.600 94.200 69.900 95.900 ;
        RECT 73.300 95.200 73.600 95.900 ;
        RECT 74.200 95.800 74.600 95.900 ;
        RECT 75.000 95.700 75.400 99.900 ;
        RECT 77.200 98.200 77.600 99.900 ;
        RECT 76.600 97.900 77.600 98.200 ;
        RECT 79.400 97.900 79.800 99.900 ;
        RECT 81.500 97.900 82.100 99.900 ;
        RECT 76.600 97.500 77.000 97.900 ;
        RECT 79.400 97.600 79.700 97.900 ;
        RECT 78.300 97.300 80.100 97.600 ;
        RECT 81.400 97.500 81.800 97.900 ;
        RECT 78.300 97.200 78.700 97.300 ;
        RECT 79.700 97.200 80.100 97.300 ;
        RECT 76.600 96.500 77.000 96.600 ;
        RECT 78.900 96.500 79.300 96.600 ;
        RECT 76.600 96.200 79.300 96.500 ;
        RECT 79.600 96.500 80.700 96.800 ;
        RECT 79.600 95.900 79.900 96.500 ;
        RECT 80.300 96.400 80.700 96.500 ;
        RECT 81.500 96.600 82.200 97.000 ;
        RECT 81.500 96.100 81.800 96.600 ;
        RECT 77.500 95.700 79.900 95.900 ;
        RECT 75.000 95.600 79.900 95.700 ;
        RECT 80.600 95.800 81.800 96.100 ;
        RECT 75.000 95.500 77.900 95.600 ;
        RECT 75.000 95.400 77.800 95.500 ;
        RECT 70.200 94.400 70.600 95.200 ;
        RECT 71.000 95.100 71.400 95.200 ;
        RECT 72.600 95.100 73.000 95.200 ;
        RECT 71.000 94.800 73.000 95.100 ;
        RECT 72.600 94.400 73.000 94.800 ;
        RECT 73.300 94.800 73.800 95.200 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 76.100 94.800 78.600 95.100 ;
        RECT 73.300 94.200 73.600 94.800 ;
        RECT 76.100 94.700 76.500 94.800 ;
        RECT 77.400 94.700 77.800 94.800 ;
        RECT 76.900 94.200 77.300 94.300 ;
        RECT 80.600 94.200 80.900 95.800 ;
        RECT 83.800 95.600 84.200 99.900 ;
        RECT 82.100 95.300 84.200 95.600 ;
        RECT 84.600 95.700 85.000 99.900 ;
        RECT 86.800 98.200 87.200 99.900 ;
        RECT 86.200 97.900 87.200 98.200 ;
        RECT 89.000 97.900 89.400 99.900 ;
        RECT 91.100 97.900 91.700 99.900 ;
        RECT 86.200 97.500 86.600 97.900 ;
        RECT 89.000 97.600 89.300 97.900 ;
        RECT 87.900 97.300 89.700 97.600 ;
        RECT 91.000 97.500 91.400 97.900 ;
        RECT 87.900 97.200 88.300 97.300 ;
        RECT 89.300 97.200 89.700 97.300 ;
        RECT 86.200 96.500 86.600 96.600 ;
        RECT 88.500 96.500 88.900 96.600 ;
        RECT 86.200 96.200 88.900 96.500 ;
        RECT 89.200 96.500 90.300 96.800 ;
        RECT 89.200 95.900 89.500 96.500 ;
        RECT 89.900 96.400 90.300 96.500 ;
        RECT 91.100 96.600 91.800 97.000 ;
        RECT 91.100 96.100 91.400 96.600 ;
        RECT 87.100 95.700 89.500 95.900 ;
        RECT 84.600 95.600 89.500 95.700 ;
        RECT 90.200 95.800 91.400 96.100 ;
        RECT 84.600 95.500 87.500 95.600 ;
        RECT 84.600 95.400 87.400 95.500 ;
        RECT 82.100 95.200 82.500 95.300 ;
        RECT 82.900 94.900 83.300 95.000 ;
        RECT 81.400 94.600 83.300 94.900 ;
        RECT 81.400 94.500 81.800 94.600 ;
        RECT 68.600 93.800 69.900 94.200 ;
        RECT 71.000 94.100 71.400 94.200 ;
        RECT 70.600 93.800 71.400 94.100 ;
        RECT 71.800 94.100 72.200 94.200 ;
        RECT 71.800 93.800 72.600 94.100 ;
        RECT 73.300 93.800 74.600 94.200 ;
        RECT 75.400 93.900 80.900 94.200 ;
        RECT 75.400 93.800 76.200 93.900 ;
        RECT 68.700 93.100 69.000 93.800 ;
        RECT 70.600 93.600 71.000 93.800 ;
        RECT 72.200 93.600 72.600 93.800 ;
        RECT 69.500 93.100 71.300 93.300 ;
        RECT 71.900 93.100 73.700 93.300 ;
        RECT 74.200 93.100 74.500 93.800 ;
        RECT 61.400 91.500 61.800 92.500 ;
        RECT 63.500 92.200 63.900 93.000 ;
        RECT 67.000 92.800 67.900 93.100 ;
        RECT 63.500 91.800 64.200 92.200 ;
        RECT 63.500 91.500 63.900 91.800 ;
        RECT 67.500 91.100 67.900 92.800 ;
        RECT 68.600 91.100 69.000 93.100 ;
        RECT 69.400 93.000 71.400 93.100 ;
        RECT 69.400 91.100 69.800 93.000 ;
        RECT 71.000 91.100 71.400 93.000 ;
        RECT 71.800 93.000 73.800 93.100 ;
        RECT 71.800 91.100 72.200 93.000 ;
        RECT 73.400 91.100 73.800 93.000 ;
        RECT 74.200 91.100 74.600 93.100 ;
        RECT 75.000 91.100 75.400 93.500 ;
        RECT 77.500 92.800 77.800 93.900 ;
        RECT 80.300 93.800 80.700 93.900 ;
        RECT 83.800 93.600 84.200 95.300 ;
        RECT 87.800 95.100 88.200 95.200 ;
        RECT 89.400 95.100 89.800 95.200 ;
        RECT 85.700 94.800 89.800 95.100 ;
        RECT 85.700 94.700 86.100 94.800 ;
        RECT 86.500 94.200 86.900 94.300 ;
        RECT 90.200 94.200 90.500 95.800 ;
        RECT 93.400 95.600 93.800 99.900 ;
        RECT 94.200 95.800 94.600 96.600 ;
        RECT 91.700 95.300 93.800 95.600 ;
        RECT 91.700 95.200 92.100 95.300 ;
        RECT 92.500 94.900 92.900 95.000 ;
        RECT 91.000 94.600 92.900 94.900 ;
        RECT 91.000 94.500 91.400 94.600 ;
        RECT 85.000 93.900 90.500 94.200 ;
        RECT 85.000 93.800 85.800 93.900 ;
        RECT 82.300 93.300 84.200 93.600 ;
        RECT 82.300 93.200 82.700 93.300 ;
        RECT 76.600 92.100 77.000 92.500 ;
        RECT 77.400 92.400 77.800 92.800 ;
        RECT 78.300 92.700 78.700 92.800 ;
        RECT 78.300 92.400 79.700 92.700 ;
        RECT 79.400 92.100 79.700 92.400 ;
        RECT 81.400 92.100 81.800 92.500 ;
        RECT 76.600 91.800 77.600 92.100 ;
        RECT 77.200 91.100 77.600 91.800 ;
        RECT 79.400 91.100 79.800 92.100 ;
        RECT 81.400 91.800 82.100 92.100 ;
        RECT 81.500 91.100 82.100 91.800 ;
        RECT 83.800 91.100 84.200 93.300 ;
        RECT 84.600 91.100 85.000 93.500 ;
        RECT 87.100 92.800 87.400 93.900 ;
        RECT 87.800 93.800 88.200 93.900 ;
        RECT 89.900 93.800 90.300 93.900 ;
        RECT 93.400 93.600 93.800 95.300 ;
        RECT 91.900 93.300 93.800 93.600 ;
        RECT 91.900 93.200 92.300 93.300 ;
        RECT 86.200 92.100 86.600 92.500 ;
        RECT 87.000 92.400 87.400 92.800 ;
        RECT 87.900 92.700 88.300 92.800 ;
        RECT 87.900 92.400 89.300 92.700 ;
        RECT 89.000 92.100 89.300 92.400 ;
        RECT 91.000 92.100 91.400 92.500 ;
        RECT 86.200 91.800 87.200 92.100 ;
        RECT 86.800 91.100 87.200 91.800 ;
        RECT 89.000 91.100 89.400 92.100 ;
        RECT 91.000 91.800 91.700 92.100 ;
        RECT 91.100 91.100 91.700 91.800 ;
        RECT 93.400 91.100 93.800 93.300 ;
        RECT 95.000 93.100 95.400 99.900 ;
        RECT 96.600 95.800 97.000 96.600 ;
        RECT 97.400 96.100 97.800 99.900 ;
        RECT 101.000 96.800 101.400 97.200 ;
        RECT 101.000 96.200 101.300 96.800 ;
        RECT 101.700 96.200 102.100 99.900 ;
        RECT 100.600 96.100 101.300 96.200 ;
        RECT 97.400 95.900 101.300 96.100 ;
        RECT 97.400 95.800 101.000 95.900 ;
        RECT 101.600 95.800 102.600 96.200 ;
        RECT 95.800 94.100 96.200 94.200 ;
        RECT 96.600 94.100 97.000 94.200 ;
        RECT 95.800 93.800 97.000 94.100 ;
        RECT 95.800 93.400 96.200 93.800 ;
        RECT 97.400 93.100 97.800 95.800 ;
        RECT 101.600 94.200 101.900 95.800 ;
        RECT 103.800 95.700 104.200 99.900 ;
        RECT 106.000 98.200 106.400 99.900 ;
        RECT 105.400 97.900 106.400 98.200 ;
        RECT 108.200 97.900 108.600 99.900 ;
        RECT 110.300 97.900 110.900 99.900 ;
        RECT 105.400 97.500 105.800 97.900 ;
        RECT 108.200 97.600 108.500 97.900 ;
        RECT 107.100 97.300 108.900 97.600 ;
        RECT 110.200 97.500 110.600 97.900 ;
        RECT 107.100 97.200 107.500 97.300 ;
        RECT 108.500 97.200 108.900 97.300 ;
        RECT 105.400 96.500 105.800 96.600 ;
        RECT 107.700 96.500 108.100 96.600 ;
        RECT 105.400 96.200 108.100 96.500 ;
        RECT 108.400 96.500 109.500 96.800 ;
        RECT 108.400 95.900 108.700 96.500 ;
        RECT 109.100 96.400 109.500 96.500 ;
        RECT 110.300 96.600 111.000 97.000 ;
        RECT 110.300 96.100 110.600 96.600 ;
        RECT 106.300 95.700 108.700 95.900 ;
        RECT 103.800 95.600 108.700 95.700 ;
        RECT 109.400 95.800 110.600 96.100 ;
        RECT 103.800 95.500 106.700 95.600 ;
        RECT 103.800 95.400 106.600 95.500 ;
        RECT 102.200 95.100 102.600 95.200 ;
        RECT 103.000 95.100 103.400 95.200 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 102.200 94.800 103.400 95.100 ;
        RECT 104.900 94.800 107.400 95.100 ;
        RECT 102.200 94.400 102.600 94.800 ;
        RECT 104.900 94.700 105.300 94.800 ;
        RECT 106.200 94.700 106.600 94.800 ;
        RECT 105.700 94.200 106.100 94.300 ;
        RECT 109.400 94.200 109.700 95.800 ;
        RECT 112.600 95.600 113.000 99.900 ;
        RECT 110.900 95.300 113.000 95.600 ;
        RECT 110.900 95.200 111.300 95.300 ;
        RECT 111.700 94.900 112.100 95.000 ;
        RECT 110.200 94.600 112.100 94.900 ;
        RECT 110.200 94.500 110.600 94.600 ;
        RECT 98.200 94.100 98.600 94.200 ;
        RECT 99.800 94.100 100.200 94.200 ;
        RECT 98.200 93.800 100.200 94.100 ;
        RECT 100.600 93.800 101.900 94.200 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 102.600 93.800 103.400 94.100 ;
        RECT 104.200 93.900 109.700 94.200 ;
        RECT 104.200 93.800 105.000 93.900 ;
        RECT 98.200 93.400 98.600 93.800 ;
        RECT 100.700 93.100 101.000 93.800 ;
        RECT 102.600 93.600 103.000 93.800 ;
        RECT 101.500 93.100 103.300 93.300 ;
        RECT 94.500 92.800 95.400 93.100 ;
        RECT 96.900 92.800 97.800 93.100 ;
        RECT 94.500 92.200 94.900 92.800 ;
        RECT 94.500 91.800 95.400 92.200 ;
        RECT 94.500 91.100 94.900 91.800 ;
        RECT 96.900 91.100 97.300 92.800 ;
        RECT 100.600 91.100 101.000 93.100 ;
        RECT 101.400 93.000 103.400 93.100 ;
        RECT 101.400 91.100 101.800 93.000 ;
        RECT 103.000 91.100 103.400 93.000 ;
        RECT 103.800 91.100 104.200 93.500 ;
        RECT 106.300 93.200 106.600 93.900 ;
        RECT 109.100 93.800 109.500 93.900 ;
        RECT 112.600 93.600 113.000 95.300 ;
        RECT 114.200 95.100 114.600 99.900 ;
        RECT 115.000 95.800 115.400 96.600 ;
        RECT 115.800 95.100 116.200 95.200 ;
        RECT 114.200 94.800 116.200 95.100 ;
        RECT 111.100 93.300 113.000 93.600 ;
        RECT 113.400 93.400 113.800 94.200 ;
        RECT 111.100 93.200 111.500 93.300 ;
        RECT 105.400 92.100 105.800 92.500 ;
        RECT 106.200 92.400 106.600 93.200 ;
        RECT 107.100 92.700 107.500 92.800 ;
        RECT 107.100 92.400 108.500 92.700 ;
        RECT 108.200 92.100 108.500 92.400 ;
        RECT 110.200 92.100 110.600 92.500 ;
        RECT 105.400 91.800 106.400 92.100 ;
        RECT 106.000 91.100 106.400 91.800 ;
        RECT 108.200 91.100 108.600 92.100 ;
        RECT 110.200 91.800 110.900 92.100 ;
        RECT 110.300 91.100 110.900 91.800 ;
        RECT 112.600 91.100 113.000 93.300 ;
        RECT 114.200 93.100 114.600 94.800 ;
        RECT 115.000 94.100 115.400 94.200 ;
        RECT 115.800 94.100 116.200 94.200 ;
        RECT 115.000 93.800 116.200 94.100 ;
        RECT 115.800 93.400 116.200 93.800 ;
        RECT 116.600 93.100 117.000 99.900 ;
        RECT 117.400 95.800 117.800 96.600 ;
        RECT 120.100 96.400 120.500 99.900 ;
        RECT 122.200 97.500 122.600 99.500 ;
        RECT 119.700 96.100 120.500 96.400 ;
        RECT 119.000 94.800 119.400 95.600 ;
        RECT 119.700 94.200 120.000 96.100 ;
        RECT 122.300 95.800 122.600 97.500 ;
        RECT 120.700 95.500 122.600 95.800 ;
        RECT 123.000 95.900 123.400 99.900 ;
        RECT 124.600 97.900 125.000 99.900 ;
        RECT 120.700 94.500 121.000 95.500 ;
        RECT 123.000 95.200 123.300 95.900 ;
        RECT 124.600 95.800 124.900 97.900 ;
        RECT 123.700 95.500 124.900 95.800 ;
        RECT 127.000 95.600 127.400 99.900 ;
        RECT 128.600 95.600 129.000 99.900 ;
        RECT 130.200 95.600 130.600 99.900 ;
        RECT 131.800 95.600 132.200 99.900 ;
        RECT 119.000 93.800 120.000 94.200 ;
        RECT 120.300 94.100 121.000 94.500 ;
        RECT 121.400 94.400 121.800 95.200 ;
        RECT 122.200 94.400 122.600 95.200 ;
        RECT 123.000 94.800 123.400 95.200 ;
        RECT 119.700 93.500 120.000 93.800 ;
        RECT 120.500 93.900 121.000 94.100 ;
        RECT 120.500 93.600 122.600 93.900 ;
        RECT 119.700 93.300 120.100 93.500 ;
        RECT 114.200 92.800 115.100 93.100 ;
        RECT 116.600 92.800 117.500 93.100 ;
        RECT 119.700 93.000 120.500 93.300 ;
        RECT 114.700 91.100 115.100 92.800 ;
        RECT 117.100 92.200 117.500 92.800 ;
        RECT 116.600 91.800 117.500 92.200 ;
        RECT 117.100 91.100 117.500 91.800 ;
        RECT 120.100 92.200 120.500 93.000 ;
        RECT 122.300 92.500 122.600 93.600 ;
        RECT 123.000 93.100 123.300 94.800 ;
        RECT 123.700 93.800 124.000 95.500 ;
        RECT 127.000 95.200 127.900 95.600 ;
        RECT 128.600 95.200 129.700 95.600 ;
        RECT 130.200 95.200 131.300 95.600 ;
        RECT 131.800 95.200 133.000 95.600 ;
        RECT 124.600 94.800 125.000 95.200 ;
        RECT 124.600 94.400 124.900 94.800 ;
        RECT 124.400 94.000 125.000 94.400 ;
        RECT 125.400 93.800 125.800 94.600 ;
        RECT 127.500 94.500 127.900 95.200 ;
        RECT 129.300 94.500 129.700 95.200 ;
        RECT 130.900 94.500 131.300 95.200 ;
        RECT 127.500 94.100 128.800 94.500 ;
        RECT 129.300 94.100 130.500 94.500 ;
        RECT 130.900 94.100 132.200 94.500 ;
        RECT 127.500 93.800 127.900 94.100 ;
        RECT 129.300 93.800 129.700 94.100 ;
        RECT 130.900 93.800 131.300 94.100 ;
        RECT 132.600 93.800 133.000 95.200 ;
        RECT 123.600 93.700 124.000 93.800 ;
        RECT 123.600 93.500 125.100 93.700 ;
        RECT 123.600 93.400 125.700 93.500 ;
        RECT 124.800 93.200 125.700 93.400 ;
        RECT 125.400 93.100 125.700 93.200 ;
        RECT 127.000 93.400 127.900 93.800 ;
        RECT 128.600 93.400 129.700 93.800 ;
        RECT 130.200 93.400 131.300 93.800 ;
        RECT 131.800 93.400 133.000 93.800 ;
        RECT 133.400 93.400 133.800 94.200 ;
        RECT 123.000 92.600 123.700 93.100 ;
        RECT 120.100 91.800 121.000 92.200 ;
        RECT 120.100 91.500 120.500 91.800 ;
        RECT 122.200 91.500 122.600 92.500 ;
        RECT 123.300 92.200 123.700 92.600 ;
        RECT 123.000 91.800 123.700 92.200 ;
        RECT 123.300 91.100 123.700 91.800 ;
        RECT 125.400 91.100 125.800 93.100 ;
        RECT 127.000 91.100 127.400 93.400 ;
        RECT 128.600 91.100 129.000 93.400 ;
        RECT 130.200 91.100 130.600 93.400 ;
        RECT 131.800 91.100 132.200 93.400 ;
        RECT 134.200 93.100 134.600 99.900 ;
        RECT 135.000 95.800 135.400 96.600 ;
        RECT 136.600 96.400 137.000 99.900 ;
        RECT 136.500 95.900 137.000 96.400 ;
        RECT 138.200 96.200 138.600 99.900 ;
        RECT 139.800 96.400 140.200 99.900 ;
        RECT 137.300 95.900 138.600 96.200 ;
        RECT 139.700 95.900 140.200 96.400 ;
        RECT 141.400 96.200 141.800 99.900 ;
        RECT 143.000 96.400 143.400 99.900 ;
        RECT 140.500 95.900 141.800 96.200 ;
        RECT 142.900 95.900 143.400 96.400 ;
        RECT 144.600 96.200 145.000 99.900 ;
        RECT 143.700 95.900 145.000 96.200 ;
        RECT 145.400 96.200 145.800 99.900 ;
        RECT 147.000 96.400 147.400 99.900 ;
        RECT 149.400 96.400 149.800 99.900 ;
        RECT 145.400 95.900 146.700 96.200 ;
        RECT 147.000 95.900 147.500 96.400 ;
        RECT 135.000 95.200 135.300 95.800 ;
        RECT 135.000 94.800 135.400 95.200 ;
        RECT 136.500 94.200 136.800 95.900 ;
        RECT 137.300 94.900 137.600 95.900 ;
        RECT 137.100 94.500 137.600 94.900 ;
        RECT 136.500 93.800 137.000 94.200 ;
        RECT 136.500 93.100 136.800 93.800 ;
        RECT 137.300 93.700 137.600 94.500 ;
        RECT 139.700 94.200 140.000 95.900 ;
        RECT 140.500 94.900 140.800 95.900 ;
        RECT 140.300 94.500 140.800 94.900 ;
        RECT 139.700 93.800 140.200 94.200 ;
        RECT 137.300 93.400 138.600 93.700 ;
        RECT 134.200 92.800 135.100 93.100 ;
        RECT 136.500 92.800 137.000 93.100 ;
        RECT 134.700 91.100 135.100 92.800 ;
        RECT 136.600 91.100 137.000 92.800 ;
        RECT 138.200 91.100 138.600 93.400 ;
        RECT 139.700 93.200 140.000 93.800 ;
        RECT 140.500 93.700 140.800 94.500 ;
        RECT 142.900 94.200 143.200 95.900 ;
        RECT 143.700 94.900 144.000 95.900 ;
        RECT 143.500 94.500 144.000 94.900 ;
        RECT 142.900 93.800 143.400 94.200 ;
        RECT 140.500 93.400 141.800 93.700 ;
        RECT 139.700 92.800 140.200 93.200 ;
        RECT 139.800 91.100 140.200 92.800 ;
        RECT 141.400 91.100 141.800 93.400 ;
        RECT 142.900 93.100 143.200 93.800 ;
        RECT 143.700 93.700 144.000 94.500 ;
        RECT 146.400 94.900 146.700 95.900 ;
        RECT 146.400 94.500 146.900 94.900 ;
        RECT 146.400 93.700 146.700 94.500 ;
        RECT 147.200 94.200 147.500 95.900 ;
        RECT 149.300 95.900 149.800 96.400 ;
        RECT 151.000 96.200 151.400 99.900 ;
        RECT 155.300 99.200 155.700 99.900 ;
        RECT 155.000 98.800 155.700 99.200 ;
        RECT 155.300 96.400 155.700 98.800 ;
        RECT 157.400 97.500 157.800 99.500 ;
        RECT 150.100 95.900 151.400 96.200 ;
        RECT 154.900 96.100 155.700 96.400 ;
        RECT 149.300 94.200 149.600 95.900 ;
        RECT 150.100 94.900 150.400 95.900 ;
        RECT 149.900 94.500 150.400 94.900 ;
        RECT 153.400 95.100 153.800 95.200 ;
        RECT 154.200 95.100 154.600 95.600 ;
        RECT 153.400 94.800 154.600 95.100 ;
        RECT 147.000 93.800 147.500 94.200 ;
        RECT 148.600 94.100 149.000 94.200 ;
        RECT 149.300 94.100 149.800 94.200 ;
        RECT 148.600 93.800 149.800 94.100 ;
        RECT 143.700 93.400 145.000 93.700 ;
        RECT 142.900 92.800 143.400 93.100 ;
        RECT 143.000 91.100 143.400 92.800 ;
        RECT 144.600 91.100 145.000 93.400 ;
        RECT 145.400 93.400 146.700 93.700 ;
        RECT 145.400 91.100 145.800 93.400 ;
        RECT 147.200 93.100 147.500 93.800 ;
        RECT 147.000 92.800 147.500 93.100 ;
        RECT 149.300 93.100 149.600 93.800 ;
        RECT 150.100 93.700 150.400 94.500 ;
        RECT 154.900 94.200 155.200 96.100 ;
        RECT 157.500 95.800 157.800 97.500 ;
        RECT 158.500 96.300 158.900 99.900 ;
        RECT 158.500 95.900 159.400 96.300 ;
        RECT 155.900 95.500 157.800 95.800 ;
        RECT 155.900 94.500 156.200 95.500 ;
        RECT 154.200 93.800 155.200 94.200 ;
        RECT 155.500 94.100 156.200 94.500 ;
        RECT 156.600 94.400 157.000 95.200 ;
        RECT 157.400 94.400 157.800 95.200 ;
        RECT 158.200 94.800 158.600 95.600 ;
        RECT 150.100 93.400 151.400 93.700 ;
        RECT 149.300 92.800 149.800 93.100 ;
        RECT 147.000 91.100 147.400 92.800 ;
        RECT 149.400 91.100 149.800 92.800 ;
        RECT 151.000 91.100 151.400 93.400 ;
        RECT 154.900 93.500 155.200 93.800 ;
        RECT 155.700 93.900 156.200 94.100 ;
        RECT 159.000 94.200 159.300 95.900 ;
        RECT 160.600 95.600 161.000 99.900 ;
        RECT 162.700 97.900 163.300 99.900 ;
        RECT 165.000 97.900 165.400 99.900 ;
        RECT 167.200 98.200 167.600 99.900 ;
        RECT 167.200 97.900 168.200 98.200 ;
        RECT 163.000 97.500 163.400 97.900 ;
        RECT 165.100 97.600 165.400 97.900 ;
        RECT 164.700 97.300 166.500 97.600 ;
        RECT 167.800 97.500 168.200 97.900 ;
        RECT 164.700 97.200 165.100 97.300 ;
        RECT 166.100 97.200 166.500 97.300 ;
        RECT 162.600 96.600 163.300 97.000 ;
        RECT 163.000 96.100 163.300 96.600 ;
        RECT 164.100 96.500 165.200 96.800 ;
        RECT 164.100 96.400 164.500 96.500 ;
        RECT 163.000 95.800 164.200 96.100 ;
        RECT 160.600 95.300 162.700 95.600 ;
        RECT 155.700 93.600 157.800 93.900 ;
        RECT 154.900 93.300 155.300 93.500 ;
        RECT 154.900 93.000 155.700 93.300 ;
        RECT 155.300 91.500 155.700 93.000 ;
        RECT 157.500 92.500 157.800 93.600 ;
        RECT 157.400 91.500 157.800 92.500 ;
        RECT 159.000 93.800 159.400 94.200 ;
        RECT 159.000 92.200 159.300 93.800 ;
        RECT 160.600 93.600 161.000 95.300 ;
        RECT 162.300 95.200 162.700 95.300 ;
        RECT 161.500 94.900 161.900 95.000 ;
        RECT 161.500 94.600 163.400 94.900 ;
        RECT 163.000 94.500 163.400 94.600 ;
        RECT 163.900 94.200 164.200 95.800 ;
        RECT 164.900 95.900 165.200 96.500 ;
        RECT 165.500 96.500 165.900 96.600 ;
        RECT 167.800 96.500 168.200 96.600 ;
        RECT 165.500 96.200 168.200 96.500 ;
        RECT 164.900 95.700 167.300 95.900 ;
        RECT 169.400 95.700 169.800 99.900 ;
        RECT 164.900 95.600 169.800 95.700 ;
        RECT 166.900 95.500 169.800 95.600 ;
        RECT 167.000 95.400 169.800 95.500 ;
        RECT 170.200 95.700 170.600 99.900 ;
        RECT 172.400 98.200 172.800 99.900 ;
        RECT 171.800 97.900 172.800 98.200 ;
        RECT 174.600 97.900 175.000 99.900 ;
        RECT 176.700 97.900 177.300 99.900 ;
        RECT 171.800 97.500 172.200 97.900 ;
        RECT 174.600 97.600 174.900 97.900 ;
        RECT 173.500 97.300 175.300 97.600 ;
        RECT 176.600 97.500 177.000 97.900 ;
        RECT 173.500 97.200 173.900 97.300 ;
        RECT 174.900 97.200 175.300 97.300 ;
        RECT 171.800 96.500 172.200 96.600 ;
        RECT 174.100 96.500 174.500 96.600 ;
        RECT 171.800 96.200 174.500 96.500 ;
        RECT 174.800 96.500 175.900 96.800 ;
        RECT 174.800 95.900 175.100 96.500 ;
        RECT 175.500 96.400 175.900 96.500 ;
        RECT 176.700 96.600 177.400 97.000 ;
        RECT 176.700 96.100 177.000 96.600 ;
        RECT 172.700 95.700 175.100 95.900 ;
        RECT 170.200 95.600 175.100 95.700 ;
        RECT 175.800 95.800 177.000 96.100 ;
        RECT 170.200 95.500 173.100 95.600 ;
        RECT 170.200 95.400 173.000 95.500 ;
        RECT 175.800 95.200 176.100 95.800 ;
        RECT 179.000 95.600 179.400 99.900 ;
        RECT 177.300 95.300 179.400 95.600 ;
        RECT 177.300 95.200 177.700 95.300 ;
        RECT 164.600 95.100 165.000 95.200 ;
        RECT 166.200 95.100 166.600 95.200 ;
        RECT 173.400 95.100 173.800 95.200 ;
        RECT 164.600 94.800 168.700 95.100 ;
        RECT 168.300 94.700 168.700 94.800 ;
        RECT 171.300 94.800 173.800 95.100 ;
        RECT 175.800 94.800 176.200 95.200 ;
        RECT 178.100 94.900 178.500 95.000 ;
        RECT 171.300 94.700 171.700 94.800 ;
        RECT 167.500 94.200 167.900 94.300 ;
        RECT 172.100 94.200 172.500 94.300 ;
        RECT 175.800 94.200 176.100 94.800 ;
        RECT 176.600 94.600 178.500 94.900 ;
        RECT 176.600 94.500 177.000 94.600 ;
        RECT 163.900 94.100 169.400 94.200 ;
        RECT 170.600 94.100 176.100 94.200 ;
        RECT 163.900 93.900 176.100 94.100 ;
        RECT 164.100 93.800 164.500 93.900 ;
        RECT 160.600 93.300 162.500 93.600 ;
        RECT 159.800 93.100 160.200 93.200 ;
        RECT 160.600 93.100 161.000 93.300 ;
        RECT 162.100 93.200 162.500 93.300 ;
        RECT 159.800 92.800 161.000 93.100 ;
        RECT 167.000 92.800 167.300 93.900 ;
        RECT 168.600 93.800 171.400 93.900 ;
        RECT 159.800 92.400 160.200 92.800 ;
        RECT 159.000 91.100 159.400 92.200 ;
        RECT 160.600 91.100 161.000 92.800 ;
        RECT 166.100 92.700 166.500 92.800 ;
        RECT 163.000 92.100 163.400 92.500 ;
        RECT 165.100 92.400 166.500 92.700 ;
        RECT 167.000 92.400 167.400 92.800 ;
        RECT 165.100 92.100 165.400 92.400 ;
        RECT 167.800 92.100 168.200 92.500 ;
        RECT 162.700 91.800 163.400 92.100 ;
        RECT 162.700 91.100 163.300 91.800 ;
        RECT 165.000 91.100 165.400 92.100 ;
        RECT 167.200 91.800 168.200 92.100 ;
        RECT 167.200 91.100 167.600 91.800 ;
        RECT 169.400 91.100 169.800 93.500 ;
        RECT 170.200 91.100 170.600 93.500 ;
        RECT 172.700 92.800 173.000 93.900 ;
        RECT 175.500 93.800 175.900 93.900 ;
        RECT 179.000 93.600 179.400 95.300 ;
        RECT 177.500 93.300 179.400 93.600 ;
        RECT 177.500 93.200 177.900 93.300 ;
        RECT 171.800 92.100 172.200 92.500 ;
        RECT 172.600 92.400 173.000 92.800 ;
        RECT 173.500 92.700 173.900 92.800 ;
        RECT 173.500 92.400 174.900 92.700 ;
        RECT 174.600 92.100 174.900 92.400 ;
        RECT 176.600 92.100 177.000 92.500 ;
        RECT 171.800 91.800 172.800 92.100 ;
        RECT 172.400 91.100 172.800 91.800 ;
        RECT 174.600 91.100 175.000 92.100 ;
        RECT 176.600 91.800 177.300 92.100 ;
        RECT 176.700 91.100 177.300 91.800 ;
        RECT 179.000 91.100 179.400 93.300 ;
        RECT 179.800 95.600 180.200 99.900 ;
        RECT 181.900 97.900 182.500 99.900 ;
        RECT 184.200 97.900 184.600 99.900 ;
        RECT 186.400 98.200 186.800 99.900 ;
        RECT 186.400 97.900 187.400 98.200 ;
        RECT 182.200 97.500 182.600 97.900 ;
        RECT 184.300 97.600 184.600 97.900 ;
        RECT 183.900 97.300 185.700 97.600 ;
        RECT 187.000 97.500 187.400 97.900 ;
        RECT 183.900 97.200 184.300 97.300 ;
        RECT 185.300 97.200 185.700 97.300 ;
        RECT 181.800 96.600 182.500 97.000 ;
        RECT 182.200 96.100 182.500 96.600 ;
        RECT 183.300 96.500 184.400 96.800 ;
        RECT 183.300 96.400 183.700 96.500 ;
        RECT 182.200 95.800 183.400 96.100 ;
        RECT 179.800 95.300 181.900 95.600 ;
        RECT 179.800 93.600 180.200 95.300 ;
        RECT 181.500 95.200 181.900 95.300 ;
        RECT 183.100 95.200 183.400 95.800 ;
        RECT 184.100 95.900 184.400 96.500 ;
        RECT 184.700 96.500 185.100 96.600 ;
        RECT 187.000 96.500 187.400 96.600 ;
        RECT 184.700 96.200 187.400 96.500 ;
        RECT 184.100 95.700 186.500 95.900 ;
        RECT 188.600 95.700 189.000 99.900 ;
        RECT 184.100 95.600 189.000 95.700 ;
        RECT 186.100 95.500 189.000 95.600 ;
        RECT 186.200 95.400 189.000 95.500 ;
        RECT 180.700 94.900 181.100 95.000 ;
        RECT 180.700 94.600 182.600 94.900 ;
        RECT 183.000 94.800 183.400 95.200 ;
        RECT 185.400 95.100 185.800 95.200 ;
        RECT 190.200 95.100 190.600 99.900 ;
        RECT 192.200 96.800 192.600 97.200 ;
        RECT 191.000 95.800 191.400 96.600 ;
        RECT 192.200 96.200 192.500 96.800 ;
        RECT 192.900 96.200 193.300 99.900 ;
        RECT 191.800 95.900 192.500 96.200 ;
        RECT 192.800 95.900 193.300 96.200 ;
        RECT 191.800 95.800 192.200 95.900 ;
        RECT 191.800 95.100 192.100 95.800 ;
        RECT 185.400 94.800 187.900 95.100 ;
        RECT 182.200 94.500 182.600 94.600 ;
        RECT 183.100 94.200 183.400 94.800 ;
        RECT 186.200 94.700 186.600 94.800 ;
        RECT 187.500 94.700 187.900 94.800 ;
        RECT 190.200 94.800 192.100 95.100 ;
        RECT 186.700 94.200 187.100 94.300 ;
        RECT 183.100 93.900 188.600 94.200 ;
        RECT 183.300 93.800 183.700 93.900 ;
        RECT 179.800 93.300 181.700 93.600 ;
        RECT 179.800 91.100 180.200 93.300 ;
        RECT 181.300 93.200 181.700 93.300 ;
        RECT 186.200 92.800 186.500 93.900 ;
        RECT 187.800 93.800 188.600 93.900 ;
        RECT 185.300 92.700 185.700 92.800 ;
        RECT 182.200 92.100 182.600 92.500 ;
        RECT 184.300 92.400 185.700 92.700 ;
        RECT 186.200 92.400 186.600 92.800 ;
        RECT 184.300 92.100 184.600 92.400 ;
        RECT 187.000 92.100 187.400 92.500 ;
        RECT 181.900 91.800 182.600 92.100 ;
        RECT 181.900 91.100 182.500 91.800 ;
        RECT 184.200 91.100 184.600 92.100 ;
        RECT 186.400 91.800 187.400 92.100 ;
        RECT 186.400 91.100 186.800 91.800 ;
        RECT 188.600 91.100 189.000 93.500 ;
        RECT 189.400 93.400 189.800 94.200 ;
        RECT 190.200 93.100 190.600 94.800 ;
        RECT 192.800 94.200 193.100 95.900 ;
        RECT 195.000 95.600 195.400 99.900 ;
        RECT 197.100 97.900 197.700 99.900 ;
        RECT 199.400 97.900 199.800 99.900 ;
        RECT 201.600 98.200 202.000 99.900 ;
        RECT 201.600 97.900 202.600 98.200 ;
        RECT 197.400 97.500 197.800 97.900 ;
        RECT 199.500 97.600 199.800 97.900 ;
        RECT 199.100 97.300 200.900 97.600 ;
        RECT 202.200 97.500 202.600 97.900 ;
        RECT 199.100 97.200 199.500 97.300 ;
        RECT 200.500 97.200 200.900 97.300 ;
        RECT 197.000 96.600 197.700 97.000 ;
        RECT 197.400 96.100 197.700 96.600 ;
        RECT 198.500 96.500 199.600 96.800 ;
        RECT 198.500 96.400 198.900 96.500 ;
        RECT 197.400 95.800 198.600 96.100 ;
        RECT 195.000 95.300 197.100 95.600 ;
        RECT 193.400 94.400 193.800 95.200 ;
        RECT 191.000 94.100 191.400 94.200 ;
        RECT 191.800 94.100 193.100 94.200 ;
        RECT 194.200 94.100 194.600 94.200 ;
        RECT 191.000 93.800 193.100 94.100 ;
        RECT 193.800 93.800 194.600 94.100 ;
        RECT 191.900 93.100 192.200 93.800 ;
        RECT 193.800 93.600 194.200 93.800 ;
        RECT 195.000 93.600 195.400 95.300 ;
        RECT 196.700 95.200 197.100 95.300 ;
        RECT 198.300 95.200 198.600 95.800 ;
        RECT 199.300 95.900 199.600 96.500 ;
        RECT 199.900 96.500 200.300 96.600 ;
        RECT 202.200 96.500 202.600 96.600 ;
        RECT 199.900 96.200 202.600 96.500 ;
        RECT 199.300 95.700 201.700 95.900 ;
        RECT 203.800 95.700 204.200 99.900 ;
        RECT 206.600 96.800 207.000 97.200 ;
        RECT 206.600 96.200 206.900 96.800 ;
        RECT 207.300 96.200 207.700 99.900 ;
        RECT 206.200 95.900 206.900 96.200 ;
        RECT 207.200 95.900 207.700 96.200 ;
        RECT 209.400 97.500 209.800 99.500 ;
        RECT 211.500 99.200 211.900 99.900 ;
        RECT 211.000 98.800 211.900 99.200 ;
        RECT 206.200 95.800 206.600 95.900 ;
        RECT 199.300 95.600 204.200 95.700 ;
        RECT 201.300 95.500 204.200 95.600 ;
        RECT 201.400 95.400 204.200 95.500 ;
        RECT 195.900 94.900 196.300 95.000 ;
        RECT 195.900 94.600 197.800 94.900 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 200.600 95.100 201.000 95.200 ;
        RECT 204.600 95.100 205.000 95.200 ;
        RECT 207.200 95.100 207.500 95.900 ;
        RECT 209.400 95.800 209.700 97.500 ;
        RECT 211.500 96.400 211.900 98.800 ;
        RECT 211.500 96.100 212.300 96.400 ;
        RECT 209.400 95.500 211.300 95.800 ;
        RECT 200.600 94.800 203.100 95.100 ;
        RECT 204.600 94.800 207.500 95.100 ;
        RECT 197.400 94.500 197.800 94.600 ;
        RECT 198.300 94.200 198.600 94.800 ;
        RECT 201.400 94.700 201.800 94.800 ;
        RECT 202.700 94.700 203.100 94.800 ;
        RECT 201.900 94.200 202.300 94.300 ;
        RECT 207.200 94.200 207.500 94.800 ;
        RECT 207.800 94.400 208.200 95.200 ;
        RECT 209.400 94.400 209.800 95.200 ;
        RECT 210.200 94.400 210.600 95.200 ;
        RECT 211.000 94.500 211.300 95.500 ;
        RECT 198.300 93.900 203.800 94.200 ;
        RECT 198.500 93.800 198.900 93.900 ;
        RECT 195.000 93.300 196.900 93.600 ;
        RECT 192.700 93.100 194.500 93.300 ;
        RECT 190.200 92.800 191.100 93.100 ;
        RECT 190.700 91.100 191.100 92.800 ;
        RECT 191.800 91.100 192.200 93.100 ;
        RECT 192.600 93.000 194.600 93.100 ;
        RECT 192.600 91.100 193.000 93.000 ;
        RECT 194.200 91.100 194.600 93.000 ;
        RECT 195.000 91.100 195.400 93.300 ;
        RECT 196.500 93.200 196.900 93.300 ;
        RECT 201.400 92.800 201.700 93.900 ;
        RECT 203.000 93.800 203.800 93.900 ;
        RECT 206.200 93.800 207.500 94.200 ;
        RECT 208.600 94.100 209.000 94.200 ;
        RECT 208.200 93.800 209.000 94.100 ;
        RECT 211.000 94.100 211.700 94.500 ;
        RECT 212.000 94.200 212.300 96.100 ;
        RECT 214.200 95.800 214.600 96.600 ;
        RECT 212.600 94.800 213.000 95.600 ;
        RECT 211.000 93.900 211.500 94.100 ;
        RECT 200.500 92.700 200.900 92.800 ;
        RECT 197.400 92.100 197.800 92.500 ;
        RECT 199.500 92.400 200.900 92.700 ;
        RECT 201.400 92.400 201.800 92.800 ;
        RECT 199.500 92.100 199.800 92.400 ;
        RECT 202.200 92.100 202.600 92.500 ;
        RECT 197.100 91.800 197.800 92.100 ;
        RECT 197.100 91.100 197.700 91.800 ;
        RECT 199.400 91.100 199.800 92.100 ;
        RECT 201.600 91.800 202.600 92.100 ;
        RECT 201.600 91.100 202.000 91.800 ;
        RECT 203.800 91.100 204.200 93.500 ;
        RECT 206.300 93.100 206.600 93.800 ;
        RECT 208.200 93.600 208.600 93.800 ;
        RECT 209.400 93.600 211.500 93.900 ;
        RECT 212.000 93.800 213.000 94.200 ;
        RECT 207.100 93.100 208.900 93.300 ;
        RECT 206.200 91.100 206.600 93.100 ;
        RECT 207.000 93.000 209.000 93.100 ;
        RECT 207.000 91.100 207.400 93.000 ;
        RECT 208.600 91.100 209.000 93.000 ;
        RECT 209.400 92.500 209.700 93.600 ;
        RECT 212.000 93.500 212.300 93.800 ;
        RECT 211.900 93.300 212.300 93.500 ;
        RECT 211.500 93.000 212.300 93.300 ;
        RECT 215.000 93.100 215.400 99.900 ;
        RECT 216.600 95.600 217.000 99.900 ;
        RECT 218.700 97.900 219.300 99.900 ;
        RECT 221.000 97.900 221.400 99.900 ;
        RECT 223.200 98.200 223.600 99.900 ;
        RECT 223.200 97.900 224.200 98.200 ;
        RECT 219.000 97.500 219.400 97.900 ;
        RECT 221.100 97.600 221.400 97.900 ;
        RECT 220.700 97.300 222.500 97.600 ;
        RECT 223.800 97.500 224.200 97.900 ;
        RECT 220.700 97.200 221.100 97.300 ;
        RECT 222.100 97.200 222.500 97.300 ;
        RECT 218.600 96.600 219.300 97.000 ;
        RECT 219.000 96.100 219.300 96.600 ;
        RECT 220.100 96.500 221.200 96.800 ;
        RECT 220.100 96.400 220.500 96.500 ;
        RECT 219.000 95.800 220.200 96.100 ;
        RECT 216.600 95.300 218.700 95.600 ;
        RECT 215.800 93.400 216.200 94.200 ;
        RECT 216.600 93.600 217.000 95.300 ;
        RECT 218.300 95.200 218.700 95.300 ;
        RECT 219.900 95.200 220.200 95.800 ;
        RECT 220.900 95.900 221.200 96.500 ;
        RECT 221.500 96.500 221.900 96.600 ;
        RECT 223.800 96.500 224.200 96.600 ;
        RECT 221.500 96.200 224.200 96.500 ;
        RECT 220.900 95.700 223.300 95.900 ;
        RECT 225.400 95.700 225.800 99.900 ;
        RECT 226.600 96.800 227.000 97.200 ;
        RECT 226.600 96.200 226.900 96.800 ;
        RECT 227.300 96.200 227.700 99.900 ;
        RECT 226.200 95.900 226.900 96.200 ;
        RECT 227.200 95.900 227.700 96.200 ;
        RECT 230.700 96.200 231.100 99.900 ;
        RECT 231.400 96.800 231.800 97.200 ;
        RECT 231.500 96.200 231.800 96.800 ;
        RECT 230.700 95.900 231.200 96.200 ;
        RECT 231.500 95.900 232.200 96.200 ;
        RECT 226.200 95.800 226.600 95.900 ;
        RECT 220.900 95.600 225.800 95.700 ;
        RECT 222.900 95.500 225.800 95.600 ;
        RECT 223.000 95.400 225.800 95.500 ;
        RECT 217.500 94.900 217.900 95.000 ;
        RECT 217.500 94.600 219.400 94.900 ;
        RECT 219.800 94.800 220.200 95.200 ;
        RECT 222.200 95.100 222.600 95.200 ;
        RECT 222.200 94.800 224.700 95.100 ;
        RECT 219.000 94.500 219.400 94.600 ;
        RECT 219.900 94.200 220.200 94.800 ;
        RECT 223.000 94.700 223.400 94.800 ;
        RECT 224.300 94.700 224.700 94.800 ;
        RECT 226.200 94.800 226.600 95.200 ;
        RECT 223.500 94.200 223.900 94.300 ;
        RECT 226.200 94.200 226.500 94.800 ;
        RECT 227.200 94.200 227.500 95.900 ;
        RECT 227.800 95.100 228.200 95.200 ;
        RECT 228.600 95.100 229.000 95.200 ;
        RECT 227.800 94.800 229.000 95.100 ;
        RECT 227.800 94.400 228.200 94.800 ;
        RECT 230.200 94.400 230.600 95.200 ;
        RECT 230.900 94.200 231.200 95.900 ;
        RECT 231.800 95.800 232.200 95.900 ;
        RECT 232.600 95.800 233.000 96.600 ;
        RECT 231.800 95.100 232.100 95.800 ;
        RECT 233.400 95.100 233.800 99.900 ;
        RECT 235.000 95.700 235.400 99.900 ;
        RECT 237.200 98.200 237.600 99.900 ;
        RECT 236.600 97.900 237.600 98.200 ;
        RECT 239.400 97.900 239.800 99.900 ;
        RECT 241.500 97.900 242.100 99.900 ;
        RECT 236.600 97.500 237.000 97.900 ;
        RECT 239.400 97.600 239.700 97.900 ;
        RECT 238.300 97.300 240.100 97.600 ;
        RECT 241.400 97.500 241.800 97.900 ;
        RECT 238.300 97.200 238.700 97.300 ;
        RECT 239.700 97.200 240.100 97.300 ;
        RECT 236.600 96.500 237.000 96.600 ;
        RECT 238.900 96.500 239.300 96.600 ;
        RECT 236.600 96.200 239.300 96.500 ;
        RECT 239.600 96.500 240.700 96.800 ;
        RECT 239.600 95.900 239.900 96.500 ;
        RECT 240.300 96.400 240.700 96.500 ;
        RECT 241.500 96.600 242.200 97.000 ;
        RECT 241.500 96.100 241.800 96.600 ;
        RECT 237.500 95.700 239.900 95.900 ;
        RECT 235.000 95.600 239.900 95.700 ;
        RECT 240.600 95.800 241.800 96.100 ;
        RECT 235.000 95.500 237.900 95.600 ;
        RECT 235.000 95.400 237.800 95.500 ;
        RECT 238.200 95.100 238.600 95.200 ;
        RECT 231.800 94.800 233.800 95.100 ;
        RECT 219.900 93.900 225.400 94.200 ;
        RECT 220.100 93.800 220.500 93.900 ;
        RECT 209.400 91.500 209.800 92.500 ;
        RECT 211.500 91.500 211.900 93.000 ;
        RECT 214.500 92.800 215.400 93.100 ;
        RECT 216.600 93.300 218.500 93.600 ;
        RECT 214.500 91.100 214.900 92.800 ;
        RECT 216.600 91.100 217.000 93.300 ;
        RECT 218.100 93.200 218.500 93.300 ;
        RECT 223.000 92.800 223.300 93.900 ;
        RECT 224.600 93.800 225.400 93.900 ;
        RECT 226.200 93.800 227.500 94.200 ;
        RECT 228.600 94.100 229.000 94.200 ;
        RECT 229.400 94.100 229.800 94.200 ;
        RECT 228.200 93.800 230.200 94.100 ;
        RECT 230.900 93.800 232.200 94.200 ;
        RECT 222.100 92.700 222.500 92.800 ;
        RECT 219.000 92.100 219.400 92.500 ;
        RECT 221.100 92.400 222.500 92.700 ;
        RECT 223.000 92.400 223.400 92.800 ;
        RECT 221.100 92.100 221.400 92.400 ;
        RECT 223.800 92.100 224.200 92.500 ;
        RECT 218.700 91.800 219.400 92.100 ;
        RECT 218.700 91.100 219.300 91.800 ;
        RECT 221.000 91.100 221.400 92.100 ;
        RECT 223.200 91.800 224.200 92.100 ;
        RECT 223.200 91.100 223.600 91.800 ;
        RECT 225.400 91.100 225.800 93.500 ;
        RECT 226.300 93.100 226.600 93.800 ;
        RECT 228.200 93.600 228.600 93.800 ;
        RECT 229.800 93.600 230.200 93.800 ;
        RECT 227.100 93.100 228.900 93.300 ;
        RECT 229.500 93.100 231.300 93.300 ;
        RECT 231.800 93.100 232.100 93.800 ;
        RECT 233.400 93.100 233.800 94.800 ;
        RECT 236.100 94.800 238.600 95.100 ;
        RECT 236.100 94.700 236.500 94.800 ;
        RECT 237.400 94.700 237.800 94.800 ;
        RECT 236.900 94.200 237.300 94.300 ;
        RECT 240.600 94.200 240.900 95.800 ;
        RECT 243.800 95.600 244.200 99.900 ;
        RECT 244.600 95.800 245.000 96.600 ;
        RECT 242.100 95.300 244.200 95.600 ;
        RECT 242.100 95.200 242.500 95.300 ;
        RECT 242.900 94.900 243.300 95.000 ;
        RECT 241.400 94.600 243.300 94.900 ;
        RECT 241.400 94.500 241.800 94.600 ;
        RECT 234.200 93.400 234.600 94.200 ;
        RECT 235.400 93.900 240.900 94.200 ;
        RECT 235.400 93.800 236.200 93.900 ;
        RECT 226.200 91.100 226.600 93.100 ;
        RECT 227.000 93.000 229.000 93.100 ;
        RECT 227.000 91.100 227.400 93.000 ;
        RECT 228.600 91.100 229.000 93.000 ;
        RECT 229.400 93.000 231.400 93.100 ;
        RECT 229.400 91.100 229.800 93.000 ;
        RECT 231.000 91.100 231.400 93.000 ;
        RECT 231.800 91.100 232.200 93.100 ;
        RECT 232.900 92.800 233.800 93.100 ;
        RECT 232.900 91.100 233.300 92.800 ;
        RECT 235.000 91.100 235.400 93.500 ;
        RECT 237.500 92.800 237.800 93.900 ;
        RECT 240.300 93.800 240.700 93.900 ;
        RECT 243.800 93.600 244.200 95.300 ;
        RECT 242.300 93.300 244.200 93.600 ;
        RECT 242.300 93.200 242.700 93.300 ;
        RECT 236.600 92.100 237.000 92.500 ;
        RECT 237.400 92.400 237.800 92.800 ;
        RECT 238.300 92.700 238.700 92.800 ;
        RECT 238.300 92.400 239.700 92.700 ;
        RECT 239.400 92.100 239.700 92.400 ;
        RECT 241.400 92.100 241.800 92.500 ;
        RECT 236.600 91.800 237.600 92.100 ;
        RECT 237.200 91.100 237.600 91.800 ;
        RECT 239.400 91.100 239.800 92.100 ;
        RECT 241.400 91.800 242.100 92.100 ;
        RECT 241.500 91.100 242.100 91.800 ;
        RECT 243.800 91.100 244.200 93.300 ;
        RECT 245.400 93.100 245.800 99.900 ;
        RECT 247.000 97.500 247.400 99.500 ;
        RECT 249.100 99.200 249.500 99.900 ;
        RECT 248.600 98.800 249.500 99.200 ;
        RECT 247.000 95.800 247.300 97.500 ;
        RECT 249.100 96.400 249.500 98.800 ;
        RECT 249.100 96.100 249.900 96.400 ;
        RECT 247.000 95.500 248.900 95.800 ;
        RECT 247.000 94.400 247.400 95.200 ;
        RECT 247.800 94.400 248.200 95.200 ;
        RECT 248.600 94.500 248.900 95.500 ;
        RECT 246.200 93.400 246.600 94.200 ;
        RECT 248.600 94.100 249.300 94.500 ;
        RECT 249.600 94.200 249.900 96.100 ;
        RECT 250.200 95.100 250.600 95.600 ;
        RECT 251.000 95.100 251.400 95.200 ;
        RECT 250.200 94.800 251.400 95.100 ;
        RECT 248.600 93.900 249.100 94.100 ;
        RECT 247.000 93.600 249.100 93.900 ;
        RECT 249.600 93.800 250.600 94.200 ;
        RECT 244.900 92.800 245.800 93.100 ;
        RECT 244.900 92.200 245.300 92.800 ;
        RECT 244.600 91.800 245.300 92.200 ;
        RECT 244.900 91.100 245.300 91.800 ;
        RECT 247.000 92.500 247.300 93.600 ;
        RECT 249.600 93.500 249.900 93.800 ;
        RECT 249.500 93.300 249.900 93.500 ;
        RECT 249.100 93.000 249.900 93.300 ;
        RECT 247.000 91.500 247.400 92.500 ;
        RECT 249.100 91.500 249.500 93.000 ;
        RECT 1.400 87.600 1.800 89.900 ;
        RECT 3.000 87.600 3.400 89.900 ;
        RECT 4.600 87.600 5.000 89.900 ;
        RECT 6.200 87.600 6.600 89.900 ;
        RECT 8.100 89.200 8.500 89.900 ;
        RECT 7.800 88.800 8.500 89.200 ;
        RECT 8.100 88.200 8.500 88.800 ;
        RECT 8.100 87.900 9.000 88.200 ;
        RECT 1.400 87.200 2.300 87.600 ;
        RECT 3.000 87.200 4.100 87.600 ;
        RECT 4.600 87.200 5.700 87.600 ;
        RECT 6.200 87.200 7.400 87.600 ;
        RECT 1.900 86.900 2.300 87.200 ;
        RECT 3.700 86.900 4.100 87.200 ;
        RECT 5.300 86.900 5.700 87.200 ;
        RECT 1.900 86.500 3.200 86.900 ;
        RECT 3.700 86.500 4.900 86.900 ;
        RECT 5.300 86.500 6.600 86.900 ;
        RECT 1.900 85.800 2.300 86.500 ;
        RECT 3.700 85.800 4.100 86.500 ;
        RECT 5.300 85.800 5.700 86.500 ;
        RECT 7.000 85.800 7.400 87.200 ;
        RECT 1.400 85.400 2.300 85.800 ;
        RECT 3.000 85.400 4.100 85.800 ;
        RECT 4.600 85.400 5.700 85.800 ;
        RECT 6.200 85.400 7.400 85.800 ;
        RECT 1.400 81.100 1.800 85.400 ;
        RECT 3.000 81.100 3.400 85.400 ;
        RECT 4.600 81.100 5.000 85.400 ;
        RECT 6.200 81.100 6.600 85.400 ;
        RECT 7.800 84.400 8.200 85.200 ;
        RECT 8.600 81.100 9.000 87.900 ;
        RECT 9.400 86.800 9.800 87.600 ;
        RECT 10.200 87.500 10.600 89.900 ;
        RECT 12.400 89.200 12.800 89.900 ;
        RECT 11.800 88.900 12.800 89.200 ;
        RECT 14.600 88.900 15.000 89.900 ;
        RECT 16.700 89.200 17.300 89.900 ;
        RECT 16.600 88.900 17.300 89.200 ;
        RECT 11.800 88.500 12.200 88.900 ;
        RECT 14.600 88.600 14.900 88.900 ;
        RECT 12.600 88.200 13.000 88.600 ;
        RECT 13.500 88.300 14.900 88.600 ;
        RECT 16.600 88.500 17.000 88.900 ;
        RECT 13.500 88.200 13.900 88.300 ;
        RECT 10.600 87.100 11.400 87.200 ;
        RECT 12.700 87.100 13.000 88.200 ;
        RECT 17.500 87.700 17.900 87.800 ;
        RECT 19.000 87.700 19.400 89.900 ;
        RECT 17.500 87.400 19.400 87.700 ;
        RECT 15.500 87.100 15.900 87.200 ;
        RECT 10.600 86.800 16.100 87.100 ;
        RECT 12.100 86.700 12.500 86.800 ;
        RECT 11.300 86.200 11.700 86.300 ;
        RECT 11.300 86.100 13.800 86.200 ;
        RECT 14.200 86.100 14.600 86.200 ;
        RECT 11.300 85.900 14.600 86.100 ;
        RECT 13.400 85.800 14.600 85.900 ;
        RECT 15.000 86.100 15.400 86.200 ;
        RECT 15.800 86.100 16.100 86.800 ;
        RECT 16.600 86.400 17.000 86.500 ;
        RECT 16.600 86.100 18.500 86.400 ;
        RECT 15.000 85.800 16.100 86.100 ;
        RECT 18.100 86.000 18.500 86.100 ;
        RECT 10.200 85.500 13.000 85.600 ;
        RECT 10.200 85.400 13.100 85.500 ;
        RECT 10.200 85.300 15.100 85.400 ;
        RECT 10.200 81.100 10.600 85.300 ;
        RECT 12.700 85.100 15.100 85.300 ;
        RECT 11.800 84.500 14.500 84.800 ;
        RECT 11.800 84.400 12.200 84.500 ;
        RECT 14.100 84.400 14.500 84.500 ;
        RECT 14.800 84.500 15.100 85.100 ;
        RECT 15.800 85.200 16.100 85.800 ;
        RECT 17.300 85.700 17.700 85.800 ;
        RECT 19.000 85.700 19.400 87.400 ;
        RECT 17.300 85.400 19.400 85.700 ;
        RECT 15.800 84.900 17.000 85.200 ;
        RECT 15.500 84.500 15.900 84.600 ;
        RECT 14.800 84.200 15.900 84.500 ;
        RECT 16.700 84.400 17.000 84.900 ;
        RECT 16.700 84.000 17.400 84.400 ;
        RECT 13.500 83.700 13.900 83.800 ;
        RECT 14.900 83.700 15.300 83.800 ;
        RECT 11.800 83.100 12.200 83.500 ;
        RECT 13.500 83.400 15.300 83.700 ;
        RECT 14.600 83.100 14.900 83.400 ;
        RECT 16.600 83.100 17.000 83.500 ;
        RECT 11.800 82.800 12.800 83.100 ;
        RECT 12.400 81.100 12.800 82.800 ;
        RECT 14.600 81.100 15.000 83.100 ;
        RECT 16.700 81.100 17.300 83.100 ;
        RECT 19.000 81.100 19.400 85.400 ;
        RECT 19.800 87.700 20.200 89.900 ;
        RECT 21.900 89.200 22.500 89.900 ;
        RECT 21.900 88.900 22.600 89.200 ;
        RECT 24.200 88.900 24.600 89.900 ;
        RECT 26.400 89.200 26.800 89.900 ;
        RECT 26.400 88.900 27.400 89.200 ;
        RECT 22.200 88.500 22.600 88.900 ;
        RECT 24.300 88.600 24.600 88.900 ;
        RECT 24.300 88.300 25.700 88.600 ;
        RECT 25.300 88.200 25.700 88.300 ;
        RECT 26.200 88.200 26.600 88.600 ;
        RECT 27.000 88.500 27.400 88.900 ;
        RECT 21.300 87.700 21.700 87.800 ;
        RECT 19.800 87.400 21.700 87.700 ;
        RECT 19.800 85.700 20.200 87.400 ;
        RECT 23.300 87.100 23.700 87.200 ;
        RECT 26.200 87.100 26.500 88.200 ;
        RECT 28.600 87.500 29.000 89.900 ;
        RECT 31.300 88.000 31.700 89.500 ;
        RECT 33.400 88.500 33.800 89.500 ;
        RECT 34.500 89.200 34.900 89.900 ;
        RECT 34.200 88.800 34.900 89.200 ;
        RECT 30.900 87.700 31.700 88.000 ;
        RECT 30.900 87.500 31.300 87.700 ;
        RECT 30.900 87.200 31.200 87.500 ;
        RECT 33.500 87.400 33.800 88.500 ;
        RECT 34.500 88.200 34.900 88.800 ;
        RECT 36.600 88.500 37.000 89.500 ;
        RECT 34.500 87.900 35.400 88.200 ;
        RECT 27.800 87.100 28.600 87.200 ;
        RECT 23.100 86.800 28.600 87.100 ;
        RECT 30.200 86.800 31.200 87.200 ;
        RECT 31.700 87.100 33.800 87.400 ;
        RECT 31.700 86.900 32.200 87.100 ;
        RECT 22.200 86.400 22.600 86.500 ;
        RECT 20.700 86.100 22.600 86.400 ;
        RECT 23.100 86.200 23.400 86.800 ;
        RECT 26.700 86.700 27.100 86.800 ;
        RECT 26.200 86.200 26.600 86.300 ;
        RECT 27.500 86.200 27.900 86.300 ;
        RECT 20.700 86.000 21.100 86.100 ;
        RECT 23.000 85.800 23.400 86.200 ;
        RECT 25.400 85.900 27.900 86.200 ;
        RECT 25.400 85.800 25.800 85.900 ;
        RECT 21.500 85.700 21.900 85.800 ;
        RECT 19.800 85.400 21.900 85.700 ;
        RECT 19.800 81.100 20.200 85.400 ;
        RECT 23.100 85.200 23.400 85.800 ;
        RECT 26.200 85.500 29.000 85.600 ;
        RECT 26.100 85.400 29.000 85.500 ;
        RECT 30.200 85.400 30.600 86.200 ;
        RECT 22.200 84.900 23.400 85.200 ;
        RECT 24.100 85.300 29.000 85.400 ;
        RECT 24.100 85.100 26.500 85.300 ;
        RECT 22.200 84.400 22.500 84.900 ;
        RECT 21.800 84.000 22.500 84.400 ;
        RECT 23.300 84.500 23.700 84.600 ;
        RECT 24.100 84.500 24.400 85.100 ;
        RECT 23.300 84.200 24.400 84.500 ;
        RECT 24.700 84.500 27.400 84.800 ;
        RECT 24.700 84.400 25.100 84.500 ;
        RECT 27.000 84.400 27.400 84.500 ;
        RECT 23.900 83.700 24.300 83.800 ;
        RECT 25.300 83.700 25.700 83.800 ;
        RECT 22.200 83.100 22.600 83.500 ;
        RECT 23.900 83.400 25.700 83.700 ;
        RECT 24.300 83.100 24.600 83.400 ;
        RECT 27.000 83.100 27.400 83.500 ;
        RECT 21.900 81.100 22.500 83.100 ;
        RECT 24.200 81.100 24.600 83.100 ;
        RECT 26.400 82.800 27.400 83.100 ;
        RECT 26.400 81.100 26.800 82.800 ;
        RECT 28.600 81.100 29.000 85.300 ;
        RECT 30.900 84.900 31.200 86.800 ;
        RECT 31.500 86.500 32.200 86.900 ;
        RECT 31.900 85.500 32.200 86.500 ;
        RECT 32.600 85.800 33.000 86.600 ;
        RECT 33.400 85.800 33.800 86.600 ;
        RECT 31.900 85.200 33.800 85.500 ;
        RECT 30.900 84.600 31.700 84.900 ;
        RECT 31.300 82.200 31.700 84.600 ;
        RECT 33.500 83.500 33.800 85.200 ;
        RECT 34.200 84.400 34.600 85.200 ;
        RECT 31.300 81.800 32.200 82.200 ;
        RECT 31.300 81.100 31.700 81.800 ;
        RECT 33.400 81.500 33.800 83.500 ;
        RECT 35.000 81.100 35.400 87.900 ;
        RECT 35.800 86.800 36.200 87.600 ;
        RECT 36.600 87.400 36.900 88.500 ;
        RECT 38.700 88.000 39.100 89.500 ;
        RECT 42.700 89.200 43.100 89.900 ;
        RECT 42.200 88.800 43.100 89.200 ;
        RECT 42.700 88.200 43.100 88.800 ;
        RECT 38.700 87.700 39.500 88.000 ;
        RECT 39.100 87.500 39.500 87.700 ;
        RECT 42.200 87.900 43.100 88.200 ;
        RECT 36.600 87.100 38.700 87.400 ;
        RECT 38.200 86.900 38.700 87.100 ;
        RECT 39.200 87.200 39.500 87.500 ;
        RECT 39.200 87.100 40.200 87.200 ;
        RECT 40.600 87.100 41.000 87.200 ;
        RECT 36.600 85.800 37.000 86.600 ;
        RECT 37.400 85.800 37.800 86.600 ;
        RECT 38.200 86.500 38.900 86.900 ;
        RECT 39.200 86.800 41.000 87.100 ;
        RECT 41.400 86.800 41.800 87.600 ;
        RECT 38.200 85.500 38.500 86.500 ;
        RECT 36.600 85.200 38.500 85.500 ;
        RECT 36.600 83.500 36.900 85.200 ;
        RECT 39.200 84.900 39.500 86.800 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 41.400 86.100 41.700 86.800 ;
        RECT 39.800 85.800 41.700 86.100 ;
        RECT 39.800 85.400 40.200 85.800 ;
        RECT 38.700 84.600 39.500 84.900 ;
        RECT 36.600 81.500 37.000 83.500 ;
        RECT 38.700 81.100 39.100 84.600 ;
        RECT 42.200 81.100 42.600 87.900 ;
        RECT 45.400 87.700 45.800 89.900 ;
        RECT 47.500 89.200 48.100 89.900 ;
        RECT 47.500 88.900 48.200 89.200 ;
        RECT 49.800 88.900 50.200 89.900 ;
        RECT 52.000 89.200 52.400 89.900 ;
        RECT 52.000 88.900 53.000 89.200 ;
        RECT 47.800 88.500 48.200 88.900 ;
        RECT 49.900 88.600 50.200 88.900 ;
        RECT 49.900 88.300 51.300 88.600 ;
        RECT 50.900 88.200 51.300 88.300 ;
        RECT 51.800 88.200 52.200 88.600 ;
        RECT 52.600 88.500 53.000 88.900 ;
        RECT 46.900 87.700 47.300 87.800 ;
        RECT 45.400 87.400 47.300 87.700 ;
        RECT 45.400 85.700 45.800 87.400 ;
        RECT 48.900 87.100 49.300 87.200 ;
        RECT 51.800 87.100 52.100 88.200 ;
        RECT 54.200 87.500 54.600 89.900 ;
        RECT 55.000 88.000 55.400 89.900 ;
        RECT 56.600 88.000 57.000 89.900 ;
        RECT 55.000 87.900 57.000 88.000 ;
        RECT 57.400 87.900 57.800 89.900 ;
        RECT 58.500 88.200 58.900 89.900 ;
        RECT 58.500 87.900 59.400 88.200 ;
        RECT 62.500 88.000 62.900 89.500 ;
        RECT 64.600 88.500 65.000 89.500 ;
        RECT 55.100 87.700 56.900 87.900 ;
        RECT 55.400 87.200 55.800 87.400 ;
        RECT 57.400 87.200 57.700 87.900 ;
        RECT 53.400 87.100 54.200 87.200 ;
        RECT 48.700 86.800 54.200 87.100 ;
        RECT 55.000 86.900 55.800 87.200 ;
        RECT 55.000 86.800 55.400 86.900 ;
        RECT 56.500 86.800 57.800 87.200 ;
        RECT 47.800 86.400 48.200 86.500 ;
        RECT 46.300 86.100 48.200 86.400 ;
        RECT 46.300 86.000 46.700 86.100 ;
        RECT 47.100 85.700 47.500 85.800 ;
        RECT 45.400 85.400 47.500 85.700 ;
        RECT 43.000 85.100 43.400 85.200 ;
        RECT 43.800 85.100 44.200 85.200 ;
        RECT 43.000 84.800 44.200 85.100 ;
        RECT 43.000 84.400 43.400 84.800 ;
        RECT 45.400 81.100 45.800 85.400 ;
        RECT 48.700 85.200 49.000 86.800 ;
        RECT 52.300 86.700 52.700 86.800 ;
        RECT 53.100 86.200 53.500 86.300 ;
        RECT 49.400 86.100 49.800 86.200 ;
        RECT 51.000 86.100 53.500 86.200 ;
        RECT 49.400 85.900 53.500 86.100 ;
        RECT 49.400 85.800 51.400 85.900 ;
        RECT 55.800 85.800 56.200 86.600 ;
        RECT 51.800 85.500 54.600 85.600 ;
        RECT 51.700 85.400 54.600 85.500 ;
        RECT 47.800 84.900 49.000 85.200 ;
        RECT 49.700 85.300 54.600 85.400 ;
        RECT 49.700 85.100 52.100 85.300 ;
        RECT 47.800 84.400 48.100 84.900 ;
        RECT 47.400 84.000 48.100 84.400 ;
        RECT 48.900 84.500 49.300 84.600 ;
        RECT 49.700 84.500 50.000 85.100 ;
        RECT 48.900 84.200 50.000 84.500 ;
        RECT 50.300 84.500 53.000 84.800 ;
        RECT 50.300 84.400 50.700 84.500 ;
        RECT 52.600 84.400 53.000 84.500 ;
        RECT 49.500 83.700 49.900 83.800 ;
        RECT 50.900 83.700 51.300 83.800 ;
        RECT 47.800 83.100 48.200 83.500 ;
        RECT 49.500 83.400 51.300 83.700 ;
        RECT 49.900 83.100 50.200 83.400 ;
        RECT 52.600 83.100 53.000 83.500 ;
        RECT 47.500 81.100 48.100 83.100 ;
        RECT 49.800 81.100 50.200 83.100 ;
        RECT 52.000 82.800 53.000 83.100 ;
        RECT 52.000 81.100 52.400 82.800 ;
        RECT 54.200 81.100 54.600 85.300 ;
        RECT 56.500 85.100 56.800 86.800 ;
        RECT 59.000 86.100 59.400 87.900 ;
        RECT 62.100 87.700 62.900 88.000 ;
        RECT 59.800 87.100 60.200 87.600 ;
        RECT 62.100 87.500 62.500 87.700 ;
        RECT 62.100 87.200 62.400 87.500 ;
        RECT 64.700 87.400 65.000 88.500 ;
        RECT 60.600 87.100 61.000 87.200 ;
        RECT 59.800 86.800 61.000 87.100 ;
        RECT 61.400 86.800 62.400 87.200 ;
        RECT 62.900 87.100 65.000 87.400 ;
        RECT 65.400 87.700 65.800 89.900 ;
        RECT 67.500 89.200 68.100 89.900 ;
        RECT 67.500 88.900 68.200 89.200 ;
        RECT 69.800 88.900 70.200 89.900 ;
        RECT 72.000 89.200 72.400 89.900 ;
        RECT 72.000 88.900 73.000 89.200 ;
        RECT 67.800 88.500 68.200 88.900 ;
        RECT 69.900 88.600 70.200 88.900 ;
        RECT 69.900 88.300 71.300 88.600 ;
        RECT 70.900 88.200 71.300 88.300 ;
        RECT 71.800 88.200 72.200 88.600 ;
        RECT 72.600 88.500 73.000 88.900 ;
        RECT 66.900 87.700 67.300 87.800 ;
        RECT 65.400 87.400 67.300 87.700 ;
        RECT 62.900 86.900 63.400 87.100 ;
        RECT 57.400 85.800 59.400 86.100 ;
        RECT 57.400 85.200 57.700 85.800 ;
        RECT 57.400 85.100 57.800 85.200 ;
        RECT 56.300 84.800 56.800 85.100 ;
        RECT 57.100 84.800 57.800 85.100 ;
        RECT 56.300 81.100 56.700 84.800 ;
        RECT 57.100 84.200 57.400 84.800 ;
        RECT 58.200 84.400 58.600 85.200 ;
        RECT 57.000 83.800 57.400 84.200 ;
        RECT 59.000 81.100 59.400 85.800 ;
        RECT 61.400 85.400 61.800 86.200 ;
        RECT 62.100 84.900 62.400 86.800 ;
        RECT 62.700 86.500 63.400 86.900 ;
        RECT 63.100 85.500 63.400 86.500 ;
        RECT 63.800 85.800 64.200 86.600 ;
        RECT 64.600 85.800 65.000 86.600 ;
        RECT 65.400 85.700 65.800 87.400 ;
        RECT 68.900 87.100 69.300 87.200 ;
        RECT 71.800 87.100 72.100 88.200 ;
        RECT 74.200 87.500 74.600 89.900 ;
        RECT 75.800 87.600 76.200 89.900 ;
        RECT 77.400 87.600 77.800 89.900 ;
        RECT 79.000 87.600 79.400 89.900 ;
        RECT 80.600 87.600 81.000 89.900 ;
        RECT 82.500 89.200 82.900 89.900 ;
        RECT 84.900 89.200 85.300 89.900 ;
        RECT 82.500 88.800 83.400 89.200 ;
        RECT 84.600 88.800 85.300 89.200 ;
        RECT 82.500 88.200 82.900 88.800 ;
        RECT 84.900 88.200 85.300 88.800 ;
        RECT 87.300 88.200 87.700 89.900 ;
        RECT 90.700 89.200 91.100 89.900 ;
        RECT 90.200 88.800 91.100 89.200 ;
        RECT 90.700 88.200 91.100 88.800 ;
        RECT 82.500 87.900 83.400 88.200 ;
        RECT 84.900 87.900 85.800 88.200 ;
        RECT 87.300 87.900 88.200 88.200 ;
        RECT 75.000 87.200 76.200 87.600 ;
        RECT 76.700 87.200 77.800 87.600 ;
        RECT 78.300 87.200 79.400 87.600 ;
        RECT 80.100 87.200 81.000 87.600 ;
        RECT 73.400 87.100 74.200 87.200 ;
        RECT 68.700 86.800 74.200 87.100 ;
        RECT 67.800 86.400 68.200 86.500 ;
        RECT 66.300 86.100 68.200 86.400 ;
        RECT 66.300 86.000 66.700 86.100 ;
        RECT 67.100 85.700 67.500 85.800 ;
        RECT 63.100 85.200 65.000 85.500 ;
        RECT 62.100 84.600 62.900 84.900 ;
        RECT 62.500 82.200 62.900 84.600 ;
        RECT 64.700 83.500 65.000 85.200 ;
        RECT 62.500 81.800 63.400 82.200 ;
        RECT 62.500 81.100 62.900 81.800 ;
        RECT 64.600 81.500 65.000 83.500 ;
        RECT 65.400 85.400 67.500 85.700 ;
        RECT 65.400 81.100 65.800 85.400 ;
        RECT 68.700 85.200 69.000 86.800 ;
        RECT 72.300 86.700 72.700 86.800 ;
        RECT 73.100 86.200 73.500 86.300 ;
        RECT 70.200 86.100 70.600 86.200 ;
        RECT 71.000 86.100 73.500 86.200 ;
        RECT 70.200 85.900 73.500 86.100 ;
        RECT 70.200 85.800 71.400 85.900 ;
        RECT 75.000 85.800 75.400 87.200 ;
        RECT 76.700 86.900 77.100 87.200 ;
        RECT 78.300 86.900 78.700 87.200 ;
        RECT 80.100 86.900 80.500 87.200 ;
        RECT 81.400 86.900 81.800 87.200 ;
        RECT 75.800 86.500 77.100 86.900 ;
        RECT 77.500 86.500 78.700 86.900 ;
        RECT 79.200 86.500 80.500 86.900 ;
        RECT 80.900 86.500 81.800 86.900 ;
        RECT 76.700 85.800 77.100 86.500 ;
        RECT 78.300 85.800 78.700 86.500 ;
        RECT 80.100 85.800 80.500 86.500 ;
        RECT 71.800 85.500 74.600 85.600 ;
        RECT 71.700 85.400 74.600 85.500 ;
        RECT 75.000 85.400 76.200 85.800 ;
        RECT 76.700 85.400 77.800 85.800 ;
        RECT 78.300 85.400 79.400 85.800 ;
        RECT 80.100 85.400 81.000 85.800 ;
        RECT 67.800 84.900 69.000 85.200 ;
        RECT 69.700 85.300 74.600 85.400 ;
        RECT 69.700 85.100 72.100 85.300 ;
        RECT 67.800 84.400 68.100 84.900 ;
        RECT 67.400 84.200 68.100 84.400 ;
        RECT 68.900 84.500 69.300 84.600 ;
        RECT 69.700 84.500 70.000 85.100 ;
        RECT 68.900 84.200 70.000 84.500 ;
        RECT 70.300 84.500 73.000 84.800 ;
        RECT 70.300 84.400 70.700 84.500 ;
        RECT 72.600 84.400 73.000 84.500 ;
        RECT 67.000 84.000 68.100 84.200 ;
        RECT 67.000 83.800 67.700 84.000 ;
        RECT 69.500 83.700 69.900 83.800 ;
        RECT 70.900 83.700 71.300 83.800 ;
        RECT 67.800 83.100 68.200 83.500 ;
        RECT 69.500 83.400 71.300 83.700 ;
        RECT 69.900 83.100 70.200 83.400 ;
        RECT 72.600 83.100 73.000 83.500 ;
        RECT 67.500 81.100 68.100 83.100 ;
        RECT 69.800 81.100 70.200 83.100 ;
        RECT 72.000 82.800 73.000 83.100 ;
        RECT 72.000 81.100 72.400 82.800 ;
        RECT 74.200 81.100 74.600 85.300 ;
        RECT 75.800 81.100 76.200 85.400 ;
        RECT 77.400 81.100 77.800 85.400 ;
        RECT 79.000 81.100 79.400 85.400 ;
        RECT 80.600 81.100 81.000 85.400 ;
        RECT 82.200 84.400 82.600 85.200 ;
        RECT 83.000 81.100 83.400 87.900 ;
        RECT 83.800 87.100 84.200 87.600 ;
        RECT 84.600 87.100 85.000 87.200 ;
        RECT 83.800 86.800 85.000 87.100 ;
        RECT 84.600 84.400 85.000 85.200 ;
        RECT 85.400 81.100 85.800 87.900 ;
        RECT 86.200 86.800 86.600 87.600 ;
        RECT 87.800 86.100 88.200 87.900 ;
        RECT 90.200 87.900 91.100 88.200 ;
        RECT 92.100 88.200 92.500 89.900 ;
        RECT 95.500 89.200 95.900 89.900 ;
        RECT 96.900 89.200 97.300 89.900 ;
        RECT 95.500 88.800 96.200 89.200 ;
        RECT 96.600 88.800 97.300 89.200 ;
        RECT 95.500 88.200 95.900 88.800 ;
        RECT 92.100 87.900 93.000 88.200 ;
        RECT 88.600 87.100 89.000 87.600 ;
        RECT 89.400 87.100 89.800 87.600 ;
        RECT 88.600 86.800 89.800 87.100 ;
        RECT 87.800 85.800 88.900 86.100 ;
        RECT 87.000 84.400 87.400 85.200 ;
        RECT 87.800 81.100 88.200 85.800 ;
        RECT 88.600 85.200 88.900 85.800 ;
        RECT 88.600 84.800 89.000 85.200 ;
        RECT 90.200 81.100 90.600 87.900 ;
        RECT 91.800 86.100 92.200 86.200 ;
        RECT 91.000 85.800 92.200 86.100 ;
        RECT 91.000 85.200 91.300 85.800 ;
        RECT 91.000 83.800 91.400 85.200 ;
        RECT 91.800 84.400 92.200 85.200 ;
        RECT 92.600 81.100 93.000 87.900 ;
        RECT 95.000 87.900 95.900 88.200 ;
        RECT 96.900 88.200 97.300 88.800 ;
        RECT 101.900 89.200 102.300 89.900 ;
        RECT 104.300 89.200 104.700 89.900 ;
        RECT 101.900 88.800 102.600 89.200 ;
        RECT 104.300 88.800 105.000 89.200 ;
        RECT 101.900 88.200 102.300 88.800 ;
        RECT 104.300 88.200 104.700 88.800 ;
        RECT 96.900 87.900 97.800 88.200 ;
        RECT 93.400 87.100 93.800 87.600 ;
        RECT 94.200 87.100 94.600 87.600 ;
        RECT 93.400 86.800 94.600 87.100 ;
        RECT 95.000 81.100 95.400 87.900 ;
        RECT 95.800 84.400 96.200 85.200 ;
        RECT 96.600 84.400 97.000 85.200 ;
        RECT 97.400 81.100 97.800 87.900 ;
        RECT 101.400 87.900 102.300 88.200 ;
        RECT 103.800 87.900 104.700 88.200 ;
        RECT 98.200 87.100 98.600 87.600 ;
        RECT 100.600 87.100 101.000 87.600 ;
        RECT 98.200 86.800 101.000 87.100 ;
        RECT 101.400 81.100 101.800 87.900 ;
        RECT 103.000 86.800 103.400 87.600 ;
        RECT 102.200 84.400 102.600 85.200 ;
        RECT 103.800 81.100 104.200 87.900 ;
        RECT 105.400 87.500 105.800 89.900 ;
        RECT 107.600 89.200 108.000 89.900 ;
        RECT 107.000 88.900 108.000 89.200 ;
        RECT 109.800 88.900 110.200 89.900 ;
        RECT 111.900 89.200 112.500 89.900 ;
        RECT 111.800 88.900 112.500 89.200 ;
        RECT 107.000 88.500 107.400 88.900 ;
        RECT 109.800 88.600 110.100 88.900 ;
        RECT 107.800 87.800 108.200 88.600 ;
        RECT 108.700 88.300 110.100 88.600 ;
        RECT 111.800 88.500 112.200 88.900 ;
        RECT 108.700 88.200 109.100 88.300 ;
        RECT 105.800 87.100 106.600 87.200 ;
        RECT 107.900 87.100 108.200 87.800 ;
        RECT 112.700 87.700 113.100 87.800 ;
        RECT 114.200 87.700 114.600 89.900 ;
        RECT 115.000 88.000 115.400 89.900 ;
        RECT 116.600 88.000 117.000 89.900 ;
        RECT 115.000 87.900 117.000 88.000 ;
        RECT 117.400 87.900 117.800 89.900 ;
        RECT 118.500 88.200 118.900 89.900 ;
        RECT 120.600 88.500 121.000 89.500 ;
        RECT 118.500 87.900 119.400 88.200 ;
        RECT 115.100 87.700 116.900 87.900 ;
        RECT 112.700 87.400 114.600 87.700 ;
        RECT 110.700 87.100 111.100 87.200 ;
        RECT 105.800 86.800 111.300 87.100 ;
        RECT 107.300 86.700 107.700 86.800 ;
        RECT 106.500 86.200 106.900 86.300 ;
        RECT 106.500 86.100 109.000 86.200 ;
        RECT 110.200 86.100 110.600 86.200 ;
        RECT 106.500 85.900 110.600 86.100 ;
        RECT 108.600 85.800 110.600 85.900 ;
        RECT 105.400 85.500 108.200 85.600 ;
        RECT 105.400 85.400 108.300 85.500 ;
        RECT 105.400 85.300 110.300 85.400 ;
        RECT 104.600 84.400 105.000 85.200 ;
        RECT 105.400 81.100 105.800 85.300 ;
        RECT 107.900 85.100 110.300 85.300 ;
        RECT 107.000 84.500 109.700 84.800 ;
        RECT 107.000 84.400 107.400 84.500 ;
        RECT 109.300 84.400 109.700 84.500 ;
        RECT 110.000 84.500 110.300 85.100 ;
        RECT 111.000 85.200 111.300 86.800 ;
        RECT 111.800 86.400 112.200 86.500 ;
        RECT 111.800 86.100 113.700 86.400 ;
        RECT 113.300 86.000 113.700 86.100 ;
        RECT 112.500 85.700 112.900 85.800 ;
        RECT 114.200 85.700 114.600 87.400 ;
        RECT 115.400 87.200 115.800 87.400 ;
        RECT 117.400 87.200 117.700 87.900 ;
        RECT 115.000 86.900 115.800 87.200 ;
        RECT 115.000 86.800 115.400 86.900 ;
        RECT 116.500 86.800 117.800 87.200 ;
        RECT 115.800 85.800 116.200 86.600 ;
        RECT 116.500 86.200 116.800 86.800 ;
        RECT 116.500 85.800 117.000 86.200 ;
        RECT 119.000 86.100 119.400 87.900 ;
        RECT 119.800 86.800 120.200 87.600 ;
        RECT 120.600 87.400 120.900 88.500 ;
        RECT 122.700 88.000 123.100 89.500 ;
        RECT 125.400 88.000 125.800 89.900 ;
        RECT 127.000 88.000 127.400 89.900 ;
        RECT 122.700 87.700 123.500 88.000 ;
        RECT 125.400 87.900 127.400 88.000 ;
        RECT 127.800 87.900 128.200 89.900 ;
        RECT 128.900 88.200 129.300 89.900 ;
        RECT 128.900 87.900 129.800 88.200 ;
        RECT 125.500 87.700 127.300 87.900 ;
        RECT 123.100 87.500 123.500 87.700 ;
        RECT 120.600 87.100 122.700 87.400 ;
        RECT 122.200 86.900 122.700 87.100 ;
        RECT 123.200 87.200 123.500 87.500 ;
        RECT 125.800 87.200 126.200 87.400 ;
        RECT 127.800 87.200 128.100 87.900 ;
        RECT 117.400 85.800 119.400 86.100 ;
        RECT 120.600 85.800 121.000 86.600 ;
        RECT 121.400 85.800 121.800 86.600 ;
        RECT 122.200 86.500 122.900 86.900 ;
        RECT 123.200 86.800 124.200 87.200 ;
        RECT 125.400 86.900 126.200 87.200 ;
        RECT 125.400 86.800 125.800 86.900 ;
        RECT 126.900 86.800 128.200 87.200 ;
        RECT 112.500 85.400 114.600 85.700 ;
        RECT 111.000 84.900 112.200 85.200 ;
        RECT 110.700 84.500 111.100 84.600 ;
        RECT 110.000 84.200 111.100 84.500 ;
        RECT 111.900 84.400 112.200 84.900 ;
        RECT 111.900 84.000 112.600 84.400 ;
        RECT 108.700 83.700 109.100 83.800 ;
        RECT 110.100 83.700 110.500 83.800 ;
        RECT 107.000 83.100 107.400 83.500 ;
        RECT 108.700 83.400 110.500 83.700 ;
        RECT 109.800 83.100 110.100 83.400 ;
        RECT 111.800 83.100 112.200 83.500 ;
        RECT 107.000 82.800 108.000 83.100 ;
        RECT 107.600 81.100 108.000 82.800 ;
        RECT 109.800 81.100 110.200 83.100 ;
        RECT 111.900 81.100 112.500 83.100 ;
        RECT 114.200 81.100 114.600 85.400 ;
        RECT 116.500 85.100 116.800 85.800 ;
        RECT 117.400 85.200 117.700 85.800 ;
        RECT 117.400 85.100 117.800 85.200 ;
        RECT 116.300 84.800 116.800 85.100 ;
        RECT 117.100 84.800 117.800 85.100 ;
        RECT 116.300 81.100 116.700 84.800 ;
        RECT 117.100 84.200 117.400 84.800 ;
        RECT 118.200 84.400 118.600 85.200 ;
        RECT 117.000 83.800 117.400 84.200 ;
        RECT 119.000 81.100 119.400 85.800 ;
        RECT 122.200 85.500 122.500 86.500 ;
        RECT 120.600 85.200 122.500 85.500 ;
        RECT 120.600 83.500 120.900 85.200 ;
        RECT 123.200 84.900 123.500 86.800 ;
        RECT 123.800 86.100 124.200 86.200 ;
        RECT 124.600 86.100 125.000 86.200 ;
        RECT 123.800 85.800 125.000 86.100 ;
        RECT 126.200 85.800 126.600 86.600 ;
        RECT 126.900 86.200 127.200 86.800 ;
        RECT 126.900 85.800 127.400 86.200 ;
        RECT 129.400 86.100 129.800 87.900 ;
        RECT 131.000 87.700 131.400 89.900 ;
        RECT 133.100 89.200 133.700 89.900 ;
        RECT 133.100 88.900 133.800 89.200 ;
        RECT 135.400 88.900 135.800 89.900 ;
        RECT 137.600 89.200 138.000 89.900 ;
        RECT 137.600 88.900 138.600 89.200 ;
        RECT 133.400 88.500 133.800 88.900 ;
        RECT 135.500 88.600 135.800 88.900 ;
        RECT 135.500 88.300 136.900 88.600 ;
        RECT 136.500 88.200 136.900 88.300 ;
        RECT 137.400 88.200 137.800 88.600 ;
        RECT 138.200 88.500 138.600 88.900 ;
        RECT 132.500 87.700 132.900 87.800 ;
        RECT 130.200 86.800 130.600 87.600 ;
        RECT 131.000 87.400 132.900 87.700 ;
        RECT 127.800 85.800 129.800 86.100 ;
        RECT 123.800 85.400 124.200 85.800 ;
        RECT 126.900 85.100 127.200 85.800 ;
        RECT 127.800 85.200 128.100 85.800 ;
        RECT 127.800 85.100 128.200 85.200 ;
        RECT 122.700 84.600 123.500 84.900 ;
        RECT 126.700 84.800 127.200 85.100 ;
        RECT 127.500 84.800 128.200 85.100 ;
        RECT 120.600 81.500 121.000 83.500 ;
        RECT 122.700 82.200 123.100 84.600 ;
        RECT 122.200 81.800 123.100 82.200 ;
        RECT 122.700 81.100 123.100 81.800 ;
        RECT 126.700 81.100 127.100 84.800 ;
        RECT 127.500 84.200 127.800 84.800 ;
        RECT 128.600 84.400 129.000 85.200 ;
        RECT 127.400 83.800 127.800 84.200 ;
        RECT 129.400 81.100 129.800 85.800 ;
        RECT 131.000 85.700 131.400 87.400 ;
        RECT 134.500 87.100 134.900 87.200 ;
        RECT 137.400 87.100 137.700 88.200 ;
        RECT 139.800 87.500 140.200 89.900 ;
        RECT 140.600 87.700 141.000 89.900 ;
        RECT 142.700 89.200 143.300 89.900 ;
        RECT 142.700 88.900 143.400 89.200 ;
        RECT 145.000 88.900 145.400 89.900 ;
        RECT 147.200 89.200 147.600 89.900 ;
        RECT 147.200 88.900 148.200 89.200 ;
        RECT 143.000 88.500 143.400 88.900 ;
        RECT 145.100 88.600 145.400 88.900 ;
        RECT 145.100 88.300 146.500 88.600 ;
        RECT 146.100 88.200 146.500 88.300 ;
        RECT 147.000 88.200 147.400 88.600 ;
        RECT 147.800 88.500 148.200 88.900 ;
        RECT 142.100 87.700 142.500 87.800 ;
        RECT 140.600 87.400 142.500 87.700 ;
        RECT 139.000 87.100 139.800 87.200 ;
        RECT 134.300 86.800 139.800 87.100 ;
        RECT 133.400 86.400 133.800 86.500 ;
        RECT 131.900 86.100 133.800 86.400 ;
        RECT 134.300 86.200 134.600 86.800 ;
        RECT 137.900 86.700 138.300 86.800 ;
        RECT 138.700 86.200 139.100 86.300 ;
        RECT 131.900 86.000 132.300 86.100 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 135.000 86.100 135.400 86.200 ;
        RECT 136.600 86.100 139.100 86.200 ;
        RECT 135.000 85.900 139.100 86.100 ;
        RECT 135.000 85.800 137.000 85.900 ;
        RECT 132.700 85.700 133.100 85.800 ;
        RECT 131.000 85.400 133.100 85.700 ;
        RECT 131.000 81.100 131.400 85.400 ;
        RECT 134.300 85.200 134.600 85.800 ;
        RECT 140.600 85.700 141.000 87.400 ;
        RECT 144.100 87.100 144.500 87.200 ;
        RECT 147.000 87.100 147.300 88.200 ;
        RECT 149.400 87.500 149.800 89.900 ;
        RECT 153.100 88.200 153.500 89.900 ;
        RECT 152.600 87.900 153.500 88.200 ;
        RECT 154.200 87.900 154.600 89.900 ;
        RECT 155.000 88.000 155.400 89.900 ;
        RECT 156.600 88.000 157.000 89.900 ;
        RECT 155.000 87.900 157.000 88.000 ;
        RECT 159.000 87.900 159.400 89.900 ;
        RECT 159.700 88.200 160.100 88.600 ;
        RECT 148.600 87.100 149.400 87.200 ;
        RECT 143.900 86.800 149.400 87.100 ;
        RECT 151.000 87.100 151.400 87.200 ;
        RECT 151.800 87.100 152.200 87.600 ;
        RECT 151.000 86.800 152.200 87.100 ;
        RECT 143.000 86.400 143.400 86.500 ;
        RECT 141.500 86.100 143.400 86.400 ;
        RECT 141.500 86.000 141.900 86.100 ;
        RECT 142.300 85.700 142.700 85.800 ;
        RECT 137.400 85.500 140.200 85.600 ;
        RECT 137.300 85.400 140.200 85.500 ;
        RECT 133.400 84.900 134.600 85.200 ;
        RECT 135.300 85.300 140.200 85.400 ;
        RECT 135.300 85.100 137.700 85.300 ;
        RECT 133.400 84.400 133.700 84.900 ;
        RECT 133.000 84.000 133.700 84.400 ;
        RECT 134.500 84.500 134.900 84.600 ;
        RECT 135.300 84.500 135.600 85.100 ;
        RECT 134.500 84.200 135.600 84.500 ;
        RECT 135.900 84.500 138.600 84.800 ;
        RECT 135.900 84.400 136.300 84.500 ;
        RECT 138.200 84.400 138.600 84.500 ;
        RECT 135.100 83.700 135.500 83.800 ;
        RECT 136.500 83.700 136.900 83.800 ;
        RECT 133.400 83.100 133.800 83.500 ;
        RECT 135.100 83.400 136.900 83.700 ;
        RECT 135.500 83.100 135.800 83.400 ;
        RECT 138.200 83.100 138.600 83.500 ;
        RECT 133.100 81.100 133.700 83.100 ;
        RECT 135.400 81.100 135.800 83.100 ;
        RECT 137.600 82.800 138.600 83.100 ;
        RECT 137.600 81.100 138.000 82.800 ;
        RECT 139.800 81.100 140.200 85.300 ;
        RECT 140.600 85.400 142.700 85.700 ;
        RECT 140.600 81.100 141.000 85.400 ;
        RECT 143.900 85.200 144.200 86.800 ;
        RECT 147.500 86.700 147.900 86.800 ;
        RECT 147.000 86.200 147.400 86.300 ;
        RECT 148.300 86.200 148.700 86.300 ;
        RECT 146.200 85.900 148.700 86.200 ;
        RECT 152.600 86.100 153.000 87.900 ;
        RECT 154.300 87.200 154.600 87.900 ;
        RECT 155.100 87.700 156.900 87.900 ;
        RECT 156.200 87.200 156.600 87.400 ;
        RECT 153.400 87.100 153.800 87.200 ;
        RECT 154.200 87.100 155.500 87.200 ;
        RECT 153.400 86.800 155.500 87.100 ;
        RECT 156.200 87.100 157.000 87.200 ;
        RECT 156.200 86.900 157.700 87.100 ;
        RECT 156.600 86.800 157.700 86.900 ;
        RECT 146.200 85.800 146.600 85.900 ;
        RECT 152.600 85.800 154.500 86.100 ;
        RECT 147.000 85.500 149.800 85.600 ;
        RECT 146.900 85.400 149.800 85.500 ;
        RECT 143.000 84.900 144.200 85.200 ;
        RECT 144.900 85.300 149.800 85.400 ;
        RECT 144.900 85.100 147.300 85.300 ;
        RECT 143.000 84.400 143.300 84.900 ;
        RECT 142.600 84.000 143.300 84.400 ;
        RECT 144.100 84.500 144.500 84.600 ;
        RECT 144.900 84.500 145.200 85.100 ;
        RECT 144.100 84.200 145.200 84.500 ;
        RECT 145.500 84.500 148.200 84.800 ;
        RECT 145.500 84.400 145.900 84.500 ;
        RECT 147.800 84.400 148.200 84.500 ;
        RECT 144.700 83.700 145.100 83.800 ;
        RECT 146.100 83.700 146.500 83.800 ;
        RECT 143.000 83.100 143.400 83.500 ;
        RECT 144.700 83.400 146.500 83.700 ;
        RECT 145.100 83.100 145.400 83.400 ;
        RECT 147.800 83.100 148.200 83.500 ;
        RECT 142.700 81.100 143.300 83.100 ;
        RECT 145.000 81.100 145.400 83.100 ;
        RECT 147.200 82.800 148.200 83.100 ;
        RECT 147.200 81.100 147.600 82.800 ;
        RECT 149.400 81.100 149.800 85.300 ;
        RECT 152.600 81.100 153.000 85.800 ;
        RECT 154.200 85.200 154.500 85.800 ;
        RECT 153.400 84.400 153.800 85.200 ;
        RECT 154.200 85.100 154.600 85.200 ;
        RECT 155.200 85.100 155.500 86.800 ;
        RECT 155.800 85.800 156.200 86.600 ;
        RECT 157.400 86.200 157.700 86.800 ;
        RECT 158.200 86.400 158.600 87.200 ;
        RECT 157.400 86.100 157.800 86.200 ;
        RECT 159.000 86.100 159.300 87.900 ;
        RECT 159.800 87.800 160.200 88.200 ;
        RECT 162.500 88.000 162.900 89.500 ;
        RECT 164.600 88.500 165.000 89.500 ;
        RECT 166.200 88.900 166.600 89.900 ;
        RECT 162.100 87.700 162.900 88.000 ;
        RECT 162.100 87.500 162.500 87.700 ;
        RECT 162.100 87.200 162.400 87.500 ;
        RECT 164.700 87.400 165.000 88.500 ;
        RECT 165.400 87.800 165.800 88.600 ;
        RECT 166.300 88.100 166.600 88.900 ;
        RECT 167.900 88.200 168.300 88.600 ;
        RECT 167.800 88.100 168.200 88.200 ;
        RECT 166.200 87.800 168.200 88.100 ;
        RECT 168.600 87.900 169.000 89.900 ;
        RECT 161.400 86.800 162.400 87.200 ;
        RECT 162.900 87.100 165.000 87.400 ;
        RECT 166.300 87.200 166.600 87.800 ;
        RECT 162.900 86.900 163.400 87.100 ;
        RECT 159.800 86.100 160.200 86.200 ;
        RECT 157.400 85.800 158.200 86.100 ;
        RECT 159.000 85.800 160.200 86.100 ;
        RECT 160.600 86.100 161.000 86.200 ;
        RECT 161.400 86.100 161.800 86.200 ;
        RECT 160.600 85.800 161.800 86.100 ;
        RECT 157.800 85.600 158.200 85.800 ;
        RECT 159.800 85.100 160.100 85.800 ;
        RECT 161.400 85.400 161.800 85.800 ;
        RECT 154.200 84.800 154.900 85.100 ;
        RECT 155.200 84.800 155.700 85.100 ;
        RECT 154.600 84.200 154.900 84.800 ;
        RECT 154.600 83.800 155.000 84.200 ;
        RECT 155.300 81.100 155.700 84.800 ;
        RECT 157.400 84.800 159.400 85.100 ;
        RECT 157.400 81.100 157.800 84.800 ;
        RECT 159.000 81.100 159.400 84.800 ;
        RECT 159.800 81.100 160.200 85.100 ;
        RECT 162.100 84.900 162.400 86.800 ;
        RECT 162.700 86.500 163.400 86.900 ;
        RECT 166.200 86.800 166.600 87.200 ;
        RECT 167.800 87.100 168.200 87.200 ;
        RECT 168.700 87.100 169.000 87.900 ;
        RECT 171.000 87.700 171.400 89.900 ;
        RECT 173.100 89.200 173.700 89.900 ;
        RECT 173.100 88.900 173.800 89.200 ;
        RECT 175.400 88.900 175.800 89.900 ;
        RECT 177.600 89.200 178.000 89.900 ;
        RECT 177.600 88.900 178.600 89.200 ;
        RECT 173.400 88.500 173.800 88.900 ;
        RECT 175.500 88.600 175.800 88.900 ;
        RECT 175.500 88.300 176.900 88.600 ;
        RECT 176.500 88.200 176.900 88.300 ;
        RECT 177.400 88.200 177.800 88.600 ;
        RECT 178.200 88.500 178.600 88.900 ;
        RECT 172.500 87.700 172.900 87.800 ;
        RECT 171.000 87.400 172.900 87.700 ;
        RECT 167.800 86.800 169.000 87.100 ;
        RECT 163.100 85.500 163.400 86.500 ;
        RECT 163.800 85.800 164.200 86.600 ;
        RECT 164.600 85.800 165.000 86.600 ;
        RECT 163.100 85.200 165.000 85.500 ;
        RECT 162.100 84.600 162.900 84.900 ;
        RECT 162.500 82.200 162.900 84.600 ;
        RECT 164.700 83.500 165.000 85.200 ;
        RECT 166.300 85.100 166.600 86.800 ;
        RECT 167.000 85.400 167.400 86.200 ;
        RECT 167.800 86.100 168.200 86.200 ;
        RECT 168.700 86.100 169.000 86.800 ;
        RECT 169.400 86.400 169.800 87.200 ;
        RECT 170.200 86.100 170.600 86.200 ;
        RECT 167.800 85.800 169.000 86.100 ;
        RECT 169.800 85.800 170.600 86.100 ;
        RECT 167.900 85.100 168.200 85.800 ;
        RECT 169.800 85.600 170.200 85.800 ;
        RECT 171.000 85.700 171.400 87.400 ;
        RECT 174.500 87.100 174.900 87.200 ;
        RECT 175.800 87.100 176.200 87.200 ;
        RECT 177.400 87.100 177.700 88.200 ;
        RECT 179.800 87.500 180.200 89.900 ;
        RECT 182.500 88.000 182.900 89.500 ;
        RECT 184.600 88.500 185.000 89.500 ;
        RECT 182.100 87.700 182.900 88.000 ;
        RECT 182.100 87.500 182.500 87.700 ;
        RECT 182.100 87.200 182.400 87.500 ;
        RECT 184.700 87.400 185.000 88.500 ;
        RECT 179.000 87.100 179.800 87.200 ;
        RECT 174.300 86.800 179.800 87.100 ;
        RECT 181.400 86.800 182.400 87.200 ;
        RECT 182.900 87.100 185.000 87.400 ;
        RECT 185.400 88.500 185.800 89.500 ;
        RECT 185.400 87.400 185.700 88.500 ;
        RECT 187.500 88.000 187.900 89.500 ;
        RECT 190.200 88.500 190.600 89.500 ;
        RECT 187.500 87.700 188.300 88.000 ;
        RECT 187.900 87.500 188.300 87.700 ;
        RECT 185.400 87.100 187.500 87.400 ;
        RECT 182.900 86.900 183.400 87.100 ;
        RECT 173.400 86.400 173.800 86.500 ;
        RECT 171.900 86.100 173.800 86.400 ;
        RECT 171.900 86.000 172.300 86.100 ;
        RECT 172.700 85.700 173.100 85.800 ;
        RECT 171.000 85.400 173.100 85.700 ;
        RECT 166.200 84.700 167.100 85.100 ;
        RECT 162.500 81.800 163.400 82.200 ;
        RECT 162.500 81.100 162.900 81.800 ;
        RECT 164.600 81.500 165.000 83.500 ;
        RECT 166.700 81.100 167.100 84.700 ;
        RECT 167.800 81.100 168.200 85.100 ;
        RECT 168.600 84.800 170.600 85.100 ;
        RECT 168.600 81.100 169.000 84.800 ;
        RECT 170.200 81.100 170.600 84.800 ;
        RECT 171.000 81.100 171.400 85.400 ;
        RECT 174.300 85.200 174.600 86.800 ;
        RECT 177.900 86.700 178.300 86.800 ;
        RECT 178.700 86.200 179.100 86.300 ;
        RECT 182.100 86.200 182.400 86.800 ;
        RECT 182.700 86.500 183.400 86.900 ;
        RECT 187.000 86.900 187.500 87.100 ;
        RECT 188.000 87.200 188.300 87.500 ;
        RECT 190.200 87.400 190.500 88.500 ;
        RECT 192.300 88.000 192.700 89.500 ;
        RECT 196.300 89.200 196.700 89.900 ;
        RECT 195.800 88.800 196.700 89.200 ;
        RECT 196.300 88.200 196.700 88.800 ;
        RECT 198.700 88.200 199.100 89.900 ;
        RECT 192.300 87.700 193.100 88.000 ;
        RECT 192.700 87.500 193.100 87.700 ;
        RECT 195.800 87.900 196.700 88.200 ;
        RECT 198.200 87.900 199.100 88.200 ;
        RECT 199.800 87.900 200.200 89.900 ;
        RECT 200.600 88.000 201.000 89.900 ;
        RECT 202.200 88.000 202.600 89.900 ;
        RECT 200.600 87.900 202.600 88.000 ;
        RECT 176.600 85.900 179.100 86.200 ;
        RECT 180.600 86.100 181.000 86.200 ;
        RECT 181.400 86.100 181.800 86.200 ;
        RECT 176.600 85.800 177.000 85.900 ;
        RECT 180.600 85.800 181.800 86.100 ;
        RECT 177.400 85.500 180.200 85.600 ;
        RECT 177.300 85.400 180.200 85.500 ;
        RECT 181.400 85.400 181.800 85.800 ;
        RECT 182.100 85.800 182.600 86.200 ;
        RECT 173.400 84.900 174.600 85.200 ;
        RECT 175.300 85.300 180.200 85.400 ;
        RECT 175.300 85.100 177.700 85.300 ;
        RECT 173.400 84.400 173.700 84.900 ;
        RECT 173.000 84.000 173.700 84.400 ;
        RECT 174.500 84.500 174.900 84.600 ;
        RECT 175.300 84.500 175.600 85.100 ;
        RECT 174.500 84.200 175.600 84.500 ;
        RECT 175.900 84.500 178.600 84.800 ;
        RECT 175.900 84.400 176.300 84.500 ;
        RECT 178.200 84.400 178.600 84.500 ;
        RECT 175.100 83.700 175.500 83.800 ;
        RECT 176.500 83.700 176.900 83.800 ;
        RECT 173.400 83.100 173.800 83.500 ;
        RECT 175.100 83.400 176.900 83.700 ;
        RECT 175.500 83.100 175.800 83.400 ;
        RECT 178.200 83.100 178.600 83.500 ;
        RECT 173.100 81.100 173.700 83.100 ;
        RECT 175.400 81.100 175.800 83.100 ;
        RECT 177.600 82.800 178.600 83.100 ;
        RECT 177.600 81.100 178.000 82.800 ;
        RECT 179.800 81.100 180.200 85.300 ;
        RECT 182.100 84.900 182.400 85.800 ;
        RECT 183.100 85.500 183.400 86.500 ;
        RECT 183.800 85.800 184.200 86.600 ;
        RECT 184.600 85.800 185.000 86.600 ;
        RECT 185.400 85.800 185.800 86.600 ;
        RECT 186.200 85.800 186.600 86.600 ;
        RECT 187.000 86.500 187.700 86.900 ;
        RECT 188.000 86.800 189.000 87.200 ;
        RECT 190.200 87.100 192.300 87.400 ;
        RECT 191.800 86.900 192.300 87.100 ;
        RECT 192.800 87.200 193.100 87.500 ;
        RECT 187.000 85.500 187.300 86.500 ;
        RECT 183.100 85.200 185.000 85.500 ;
        RECT 182.100 84.600 182.900 84.900 ;
        RECT 182.500 81.100 182.900 84.600 ;
        RECT 184.700 83.500 185.000 85.200 ;
        RECT 184.600 81.500 185.000 83.500 ;
        RECT 185.400 85.200 187.300 85.500 ;
        RECT 185.400 83.500 185.700 85.200 ;
        RECT 188.000 84.900 188.300 86.800 ;
        RECT 188.600 85.400 189.000 86.200 ;
        RECT 190.200 85.800 190.600 86.600 ;
        RECT 191.000 85.800 191.400 86.600 ;
        RECT 191.800 86.500 192.500 86.900 ;
        RECT 192.800 86.800 193.800 87.200 ;
        RECT 195.000 86.800 195.400 87.600 ;
        RECT 191.800 85.500 192.100 86.500 ;
        RECT 187.500 84.600 188.300 84.900 ;
        RECT 190.200 85.200 192.100 85.500 ;
        RECT 185.400 81.500 185.800 83.500 ;
        RECT 187.500 82.200 187.900 84.600 ;
        RECT 190.200 83.500 190.500 85.200 ;
        RECT 192.800 84.900 193.100 86.800 ;
        RECT 193.400 86.100 193.800 86.200 ;
        RECT 195.000 86.100 195.300 86.800 ;
        RECT 193.400 85.800 195.300 86.100 ;
        RECT 193.400 85.400 193.800 85.800 ;
        RECT 192.300 84.600 193.100 84.900 ;
        RECT 187.500 81.800 188.200 82.200 ;
        RECT 187.500 81.100 187.900 81.800 ;
        RECT 190.200 81.500 190.600 83.500 ;
        RECT 192.300 82.200 192.700 84.600 ;
        RECT 192.300 81.800 193.000 82.200 ;
        RECT 192.300 81.100 192.700 81.800 ;
        RECT 195.800 81.100 196.200 87.900 ;
        RECT 197.400 86.800 197.800 87.600 ;
        RECT 198.200 86.100 198.600 87.900 ;
        RECT 199.900 87.200 200.200 87.900 ;
        RECT 200.700 87.700 202.500 87.900 ;
        RECT 204.600 87.700 205.000 89.900 ;
        RECT 206.700 89.200 207.300 89.900 ;
        RECT 206.700 88.900 207.400 89.200 ;
        RECT 209.000 88.900 209.400 89.900 ;
        RECT 211.200 89.200 211.600 89.900 ;
        RECT 211.200 88.900 212.200 89.200 ;
        RECT 207.000 88.500 207.400 88.900 ;
        RECT 209.100 88.600 209.400 88.900 ;
        RECT 209.100 88.300 210.500 88.600 ;
        RECT 210.100 88.200 210.500 88.300 ;
        RECT 211.000 88.200 211.400 88.600 ;
        RECT 211.800 88.500 212.200 88.900 ;
        RECT 206.100 87.700 206.500 87.800 ;
        RECT 204.600 87.400 206.500 87.700 ;
        RECT 201.800 87.200 202.200 87.400 ;
        RECT 199.800 86.800 201.100 87.200 ;
        RECT 201.800 86.900 202.600 87.200 ;
        RECT 202.200 86.800 202.600 86.900 ;
        RECT 198.200 85.800 200.100 86.100 ;
        RECT 196.600 84.400 197.000 85.200 ;
        RECT 198.200 81.100 198.600 85.800 ;
        RECT 199.800 85.200 200.100 85.800 ;
        RECT 200.800 85.200 201.100 86.800 ;
        RECT 201.400 86.100 201.800 86.600 ;
        RECT 203.000 86.100 203.400 86.200 ;
        RECT 201.400 85.800 203.400 86.100 ;
        RECT 204.600 85.700 205.000 87.400 ;
        RECT 208.100 87.100 208.500 87.200 ;
        RECT 211.000 87.100 211.300 88.200 ;
        RECT 213.400 87.500 213.800 89.900 ;
        RECT 216.100 88.000 216.500 89.500 ;
        RECT 218.200 88.500 218.600 89.500 ;
        RECT 215.700 87.700 216.500 88.000 ;
        RECT 215.700 87.500 216.100 87.700 ;
        RECT 215.700 87.200 216.000 87.500 ;
        RECT 218.300 87.400 218.600 88.500 ;
        RECT 220.300 89.200 220.700 89.900 ;
        RECT 220.300 88.800 221.000 89.200 ;
        RECT 220.300 88.200 220.700 88.800 ;
        RECT 219.800 87.900 220.700 88.200 ;
        RECT 221.400 88.500 221.800 89.500 ;
        RECT 212.600 87.100 213.400 87.200 ;
        RECT 215.000 87.100 216.000 87.200 ;
        RECT 207.900 86.800 213.400 87.100 ;
        RECT 214.200 86.800 216.000 87.100 ;
        RECT 216.500 87.100 218.600 87.400 ;
        RECT 216.500 86.900 217.000 87.100 ;
        RECT 207.000 86.400 207.400 86.500 ;
        RECT 205.500 86.100 207.400 86.400 ;
        RECT 205.500 86.000 205.900 86.100 ;
        RECT 206.300 85.700 206.700 85.800 ;
        RECT 204.600 85.400 206.700 85.700 ;
        RECT 199.000 84.400 199.400 85.200 ;
        RECT 199.800 85.100 200.200 85.200 ;
        RECT 199.800 84.800 200.500 85.100 ;
        RECT 200.800 84.800 201.800 85.200 ;
        RECT 200.200 84.200 200.500 84.800 ;
        RECT 200.200 83.800 200.600 84.200 ;
        RECT 200.900 81.100 201.300 84.800 ;
        RECT 204.600 81.100 205.000 85.400 ;
        RECT 207.900 85.200 208.200 86.800 ;
        RECT 211.500 86.700 211.900 86.800 ;
        RECT 212.300 86.200 212.700 86.300 ;
        RECT 210.200 85.900 212.700 86.200 ;
        RECT 214.200 86.200 214.500 86.800 ;
        RECT 210.200 85.800 210.600 85.900 ;
        RECT 214.200 85.800 214.600 86.200 ;
        RECT 211.000 85.500 213.800 85.600 ;
        RECT 210.900 85.400 213.800 85.500 ;
        RECT 215.000 85.400 215.400 86.200 ;
        RECT 207.000 84.900 208.200 85.200 ;
        RECT 208.900 85.300 213.800 85.400 ;
        RECT 208.900 85.100 211.300 85.300 ;
        RECT 207.000 84.400 207.300 84.900 ;
        RECT 206.600 84.000 207.300 84.400 ;
        RECT 208.100 84.500 208.500 84.600 ;
        RECT 208.900 84.500 209.200 85.100 ;
        RECT 208.100 84.200 209.200 84.500 ;
        RECT 209.500 84.500 212.200 84.800 ;
        RECT 209.500 84.400 209.900 84.500 ;
        RECT 211.800 84.400 212.200 84.500 ;
        RECT 208.700 83.700 209.100 83.800 ;
        RECT 210.100 83.700 210.500 83.800 ;
        RECT 207.000 83.100 207.400 83.500 ;
        RECT 208.700 83.400 210.500 83.700 ;
        RECT 209.100 83.100 209.400 83.400 ;
        RECT 211.800 83.100 212.200 83.500 ;
        RECT 206.700 81.100 207.300 83.100 ;
        RECT 209.000 81.100 209.400 83.100 ;
        RECT 211.200 82.800 212.200 83.100 ;
        RECT 211.200 81.100 211.600 82.800 ;
        RECT 213.400 81.100 213.800 85.300 ;
        RECT 215.700 84.900 216.000 86.800 ;
        RECT 216.300 86.500 217.000 86.900 ;
        RECT 219.000 86.800 219.400 87.600 ;
        RECT 216.700 85.500 217.000 86.500 ;
        RECT 217.400 85.800 217.800 86.600 ;
        RECT 218.200 85.800 218.600 86.600 ;
        RECT 216.700 85.200 218.600 85.500 ;
        RECT 215.700 84.600 216.500 84.900 ;
        RECT 216.100 81.100 216.500 84.600 ;
        RECT 218.300 83.500 218.600 85.200 ;
        RECT 218.200 81.500 218.600 83.500 ;
        RECT 219.800 81.100 220.200 87.900 ;
        RECT 221.400 87.400 221.700 88.500 ;
        RECT 223.500 88.000 223.900 89.500 ;
        RECT 227.500 88.200 227.900 89.900 ;
        RECT 223.500 87.700 224.300 88.000 ;
        RECT 223.900 87.500 224.300 87.700 ;
        RECT 227.000 87.900 227.900 88.200 ;
        RECT 228.600 87.900 229.000 89.900 ;
        RECT 229.400 88.000 229.800 89.900 ;
        RECT 231.000 88.000 231.400 89.900 ;
        RECT 229.400 87.900 231.400 88.000 ;
        RECT 221.400 87.100 223.500 87.400 ;
        RECT 223.000 86.900 223.500 87.100 ;
        RECT 224.000 87.200 224.300 87.500 ;
        RECT 221.400 85.800 221.800 86.600 ;
        RECT 222.200 85.800 222.600 86.600 ;
        RECT 223.000 86.500 223.700 86.900 ;
        RECT 224.000 86.800 225.000 87.200 ;
        RECT 226.200 87.100 226.600 87.600 ;
        RECT 225.400 86.800 226.600 87.100 ;
        RECT 223.000 85.500 223.300 86.500 ;
        RECT 221.400 85.200 223.300 85.500 ;
        RECT 220.600 84.400 221.000 85.200 ;
        RECT 221.400 83.500 221.700 85.200 ;
        RECT 224.000 84.900 224.300 86.800 ;
        RECT 224.600 86.100 225.000 86.200 ;
        RECT 225.400 86.100 225.700 86.800 ;
        RECT 224.600 85.800 225.700 86.100 ;
        RECT 227.000 86.100 227.400 87.900 ;
        RECT 228.700 87.200 229.000 87.900 ;
        RECT 229.500 87.700 231.300 87.900 ;
        RECT 231.800 87.500 232.200 89.900 ;
        RECT 234.000 89.200 234.400 89.900 ;
        RECT 233.400 88.900 234.400 89.200 ;
        RECT 236.200 88.900 236.600 89.900 ;
        RECT 238.300 89.200 238.900 89.900 ;
        RECT 238.200 88.900 238.900 89.200 ;
        RECT 233.400 88.500 233.800 88.900 ;
        RECT 236.200 88.600 236.500 88.900 ;
        RECT 234.200 88.200 234.600 88.600 ;
        RECT 235.100 88.300 236.500 88.600 ;
        RECT 238.200 88.500 238.600 88.900 ;
        RECT 235.100 88.200 235.500 88.300 ;
        RECT 230.600 87.200 231.000 87.400 ;
        RECT 228.600 86.800 229.900 87.200 ;
        RECT 230.600 86.900 231.400 87.200 ;
        RECT 231.000 86.800 231.400 86.900 ;
        RECT 232.200 87.100 233.000 87.200 ;
        RECT 234.300 87.100 234.600 88.200 ;
        RECT 239.100 87.700 239.500 87.800 ;
        RECT 240.600 87.700 241.000 89.900 ;
        RECT 241.400 88.000 241.800 89.900 ;
        RECT 243.000 88.000 243.400 89.900 ;
        RECT 241.400 87.900 243.400 88.000 ;
        RECT 243.800 87.900 244.200 89.900 ;
        RECT 241.500 87.700 243.300 87.900 ;
        RECT 239.100 87.400 241.000 87.700 ;
        RECT 237.100 87.100 237.500 87.200 ;
        RECT 232.200 86.800 237.700 87.100 ;
        RECT 227.000 85.800 228.900 86.100 ;
        RECT 224.600 85.400 225.000 85.800 ;
        RECT 223.500 84.600 224.300 84.900 ;
        RECT 221.400 81.500 221.800 83.500 ;
        RECT 223.500 82.200 223.900 84.600 ;
        RECT 223.500 81.800 224.200 82.200 ;
        RECT 223.500 81.100 223.900 81.800 ;
        RECT 227.000 81.100 227.400 85.800 ;
        RECT 228.600 85.200 228.900 85.800 ;
        RECT 229.600 85.200 229.900 86.800 ;
        RECT 233.700 86.700 234.100 86.800 ;
        RECT 230.200 85.800 230.600 86.600 ;
        RECT 232.900 86.200 233.300 86.300 ;
        RECT 234.200 86.200 234.600 86.300 ;
        RECT 232.900 85.900 235.400 86.200 ;
        RECT 235.000 85.800 235.400 85.900 ;
        RECT 231.800 85.500 234.600 85.600 ;
        RECT 231.800 85.400 234.700 85.500 ;
        RECT 231.800 85.300 236.700 85.400 ;
        RECT 227.800 84.400 228.200 85.200 ;
        RECT 228.600 85.100 229.000 85.200 ;
        RECT 228.600 84.800 229.300 85.100 ;
        RECT 229.600 84.800 230.600 85.200 ;
        RECT 229.000 84.200 229.300 84.800 ;
        RECT 229.000 83.800 229.400 84.200 ;
        RECT 229.700 81.100 230.100 84.800 ;
        RECT 231.800 81.100 232.200 85.300 ;
        RECT 234.300 85.100 236.700 85.300 ;
        RECT 233.400 84.500 236.100 84.800 ;
        RECT 233.400 84.400 233.800 84.500 ;
        RECT 235.700 84.400 236.100 84.500 ;
        RECT 236.400 84.500 236.700 85.100 ;
        RECT 237.400 85.200 237.700 86.800 ;
        RECT 238.200 86.400 238.600 86.500 ;
        RECT 238.200 86.100 240.100 86.400 ;
        RECT 239.700 86.000 240.100 86.100 ;
        RECT 238.900 85.700 239.300 85.800 ;
        RECT 240.600 85.700 241.000 87.400 ;
        RECT 241.800 87.200 242.200 87.400 ;
        RECT 243.800 87.200 244.100 87.900 ;
        RECT 245.400 87.600 245.800 89.900 ;
        RECT 247.000 87.600 247.400 89.900 ;
        RECT 248.600 87.600 249.000 89.900 ;
        RECT 250.200 87.600 250.600 89.900 ;
        RECT 244.600 87.200 245.800 87.600 ;
        RECT 246.300 87.200 247.400 87.600 ;
        RECT 247.900 87.200 249.000 87.600 ;
        RECT 249.700 87.200 250.600 87.600 ;
        RECT 241.400 86.900 242.200 87.200 ;
        RECT 241.400 86.800 241.800 86.900 ;
        RECT 242.900 86.800 244.200 87.200 ;
        RECT 242.200 85.800 242.600 86.600 ;
        RECT 242.900 86.100 243.200 86.800 ;
        RECT 243.800 86.100 244.200 86.200 ;
        RECT 242.900 85.800 244.200 86.100 ;
        RECT 244.600 85.800 245.000 87.200 ;
        RECT 246.300 86.900 246.700 87.200 ;
        RECT 247.900 86.900 248.300 87.200 ;
        RECT 249.700 86.900 250.100 87.200 ;
        RECT 251.000 86.900 251.400 87.200 ;
        RECT 245.400 86.500 246.700 86.900 ;
        RECT 247.100 86.500 248.300 86.900 ;
        RECT 248.800 86.500 250.100 86.900 ;
        RECT 250.500 86.500 251.400 86.900 ;
        RECT 246.300 85.800 246.700 86.500 ;
        RECT 247.900 85.800 248.300 86.500 ;
        RECT 249.700 85.800 250.100 86.500 ;
        RECT 238.900 85.400 241.000 85.700 ;
        RECT 237.400 84.900 238.600 85.200 ;
        RECT 237.100 84.500 237.500 84.600 ;
        RECT 236.400 84.200 237.500 84.500 ;
        RECT 238.300 84.400 238.600 84.900 ;
        RECT 238.300 84.000 239.000 84.400 ;
        RECT 235.100 83.700 235.500 83.800 ;
        RECT 236.500 83.700 236.900 83.800 ;
        RECT 233.400 83.100 233.800 83.500 ;
        RECT 235.100 83.400 236.900 83.700 ;
        RECT 236.200 83.100 236.500 83.400 ;
        RECT 238.200 83.100 238.600 83.500 ;
        RECT 233.400 82.800 234.400 83.100 ;
        RECT 234.000 81.100 234.400 82.800 ;
        RECT 236.200 81.100 236.600 83.100 ;
        RECT 238.300 81.100 238.900 83.100 ;
        RECT 240.600 81.100 241.000 85.400 ;
        RECT 242.900 85.100 243.200 85.800 ;
        RECT 244.600 85.400 245.800 85.800 ;
        RECT 246.300 85.400 247.400 85.800 ;
        RECT 247.900 85.400 249.000 85.800 ;
        RECT 249.700 85.400 250.600 85.800 ;
        RECT 243.800 85.100 244.200 85.200 ;
        RECT 242.700 84.800 243.200 85.100 ;
        RECT 243.500 84.800 244.200 85.100 ;
        RECT 242.700 81.100 243.100 84.800 ;
        RECT 243.500 84.200 243.800 84.800 ;
        RECT 243.400 83.800 243.800 84.200 ;
        RECT 245.400 81.100 245.800 85.400 ;
        RECT 247.000 81.100 247.400 85.400 ;
        RECT 248.600 81.100 249.000 85.400 ;
        RECT 250.200 81.100 250.600 85.400 ;
        RECT 0.600 75.700 1.000 79.900 ;
        RECT 2.800 78.200 3.200 79.900 ;
        RECT 2.200 77.900 3.200 78.200 ;
        RECT 5.000 77.900 5.400 79.900 ;
        RECT 7.100 77.900 7.700 79.900 ;
        RECT 2.200 77.500 2.600 77.900 ;
        RECT 5.000 77.600 5.300 77.900 ;
        RECT 3.900 77.300 5.700 77.600 ;
        RECT 7.000 77.500 7.400 77.900 ;
        RECT 3.900 77.200 4.300 77.300 ;
        RECT 5.300 77.200 5.700 77.300 ;
        RECT 2.200 76.500 2.600 76.600 ;
        RECT 4.500 76.500 4.900 76.600 ;
        RECT 2.200 76.200 4.900 76.500 ;
        RECT 5.200 76.500 6.300 76.800 ;
        RECT 5.200 75.900 5.500 76.500 ;
        RECT 5.900 76.400 6.300 76.500 ;
        RECT 7.100 76.600 7.800 77.000 ;
        RECT 7.100 76.100 7.400 76.600 ;
        RECT 3.100 75.700 5.500 75.900 ;
        RECT 0.600 75.600 5.500 75.700 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 0.600 75.500 3.500 75.600 ;
        RECT 0.600 75.400 3.400 75.500 ;
        RECT 6.200 75.200 6.500 75.800 ;
        RECT 9.400 75.600 9.800 79.900 ;
        RECT 11.800 76.200 12.200 79.900 ;
        RECT 11.100 75.900 12.200 76.200 ;
        RECT 12.600 76.200 13.000 79.900 ;
        RECT 14.200 76.200 14.600 79.900 ;
        RECT 12.600 75.900 14.600 76.200 ;
        RECT 15.000 75.900 15.400 79.900 ;
        RECT 16.100 76.300 16.500 79.900 ;
        RECT 16.100 75.900 17.000 76.300 ;
        RECT 19.500 76.200 19.900 79.900 ;
        RECT 20.200 76.800 20.600 77.200 ;
        RECT 20.300 76.200 20.600 76.800 ;
        RECT 19.500 75.900 20.000 76.200 ;
        RECT 20.300 75.900 21.000 76.200 ;
        RECT 11.100 75.600 11.400 75.900 ;
        RECT 7.700 75.300 9.800 75.600 ;
        RECT 7.700 75.200 8.100 75.300 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 1.700 74.800 4.200 75.100 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 8.500 74.900 8.900 75.000 ;
        RECT 1.700 74.700 2.100 74.800 ;
        RECT 3.000 74.700 3.400 74.800 ;
        RECT 2.500 74.200 2.900 74.300 ;
        RECT 6.200 74.200 6.500 74.800 ;
        RECT 7.000 74.600 8.900 74.900 ;
        RECT 7.000 74.500 7.400 74.600 ;
        RECT 1.000 73.900 6.500 74.200 ;
        RECT 1.000 73.800 1.800 73.900 ;
        RECT 0.600 71.100 1.000 73.500 ;
        RECT 3.100 72.800 3.400 73.900 ;
        RECT 5.900 73.800 6.300 73.900 ;
        RECT 9.400 73.600 9.800 75.300 ;
        RECT 10.800 75.200 11.400 75.600 ;
        RECT 13.000 75.200 13.400 75.400 ;
        RECT 15.000 75.200 15.300 75.900 ;
        RECT 7.900 73.300 9.800 73.600 ;
        RECT 11.100 73.700 11.400 75.200 ;
        RECT 11.800 74.400 12.200 75.200 ;
        RECT 12.600 74.900 13.400 75.200 ;
        RECT 14.200 74.900 15.400 75.200 ;
        RECT 12.600 74.800 13.000 74.900 ;
        RECT 13.400 73.800 13.800 74.600 ;
        RECT 11.100 73.400 12.200 73.700 ;
        RECT 7.900 73.200 8.300 73.300 ;
        RECT 2.200 72.100 2.600 72.500 ;
        RECT 3.000 72.400 3.400 72.800 ;
        RECT 3.900 72.700 4.300 72.800 ;
        RECT 3.900 72.400 5.300 72.700 ;
        RECT 5.000 72.100 5.300 72.400 ;
        RECT 7.000 72.100 7.400 72.500 ;
        RECT 2.200 71.800 3.200 72.100 ;
        RECT 2.800 71.100 3.200 71.800 ;
        RECT 5.000 71.100 5.400 72.100 ;
        RECT 7.000 71.800 7.700 72.100 ;
        RECT 7.100 71.100 7.700 71.800 ;
        RECT 9.400 71.100 9.800 73.300 ;
        RECT 11.800 71.100 12.200 73.400 ;
        RECT 14.200 73.100 14.500 74.900 ;
        RECT 15.000 74.800 15.400 74.900 ;
        RECT 15.800 74.800 16.200 75.600 ;
        RECT 16.600 74.200 16.900 75.900 ;
        RECT 19.700 75.200 20.000 75.900 ;
        RECT 20.600 75.800 21.000 75.900 ;
        RECT 21.400 75.800 21.800 76.600 ;
        RECT 19.000 74.400 19.400 75.200 ;
        RECT 19.700 74.800 20.200 75.200 ;
        RECT 20.600 75.100 20.900 75.800 ;
        RECT 22.200 75.100 22.600 79.900 ;
        RECT 23.800 76.200 24.200 79.900 ;
        RECT 25.400 76.200 25.800 79.900 ;
        RECT 23.800 75.900 25.800 76.200 ;
        RECT 26.200 75.900 26.600 79.900 ;
        RECT 27.300 76.300 27.700 79.900 ;
        RECT 27.300 75.900 28.200 76.300 ;
        RECT 30.700 76.200 31.100 79.900 ;
        RECT 31.400 76.800 31.800 77.200 ;
        RECT 31.500 76.200 31.800 76.800 ;
        RECT 30.700 75.900 31.200 76.200 ;
        RECT 31.500 75.900 32.200 76.200 ;
        RECT 24.200 75.200 24.600 75.400 ;
        RECT 26.200 75.200 26.500 75.900 ;
        RECT 20.600 74.800 22.600 75.100 ;
        RECT 23.800 74.900 24.600 75.200 ;
        RECT 25.400 74.900 26.600 75.200 ;
        RECT 23.800 74.800 24.200 74.900 ;
        RECT 19.700 74.200 20.000 74.800 ;
        RECT 16.600 73.800 17.000 74.200 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 18.200 73.800 19.000 74.100 ;
        RECT 19.700 73.800 21.000 74.200 ;
        RECT 15.000 73.100 15.400 73.200 ;
        RECT 16.600 73.100 16.900 73.800 ;
        RECT 18.600 73.600 19.000 73.800 ;
        RECT 14.200 71.100 14.600 73.100 ;
        RECT 15.000 72.800 16.900 73.100 ;
        RECT 14.900 72.400 15.300 72.800 ;
        RECT 16.600 72.100 16.900 72.800 ;
        RECT 17.400 72.400 17.800 73.200 ;
        RECT 18.300 73.100 20.100 73.300 ;
        RECT 20.600 73.100 20.900 73.800 ;
        RECT 22.200 73.100 22.600 74.800 ;
        RECT 23.000 73.400 23.400 74.200 ;
        RECT 24.600 73.800 25.000 74.600 ;
        RECT 18.200 73.000 20.200 73.100 ;
        RECT 16.600 71.100 17.000 72.100 ;
        RECT 18.200 71.100 18.600 73.000 ;
        RECT 19.800 71.100 20.200 73.000 ;
        RECT 20.600 71.100 21.000 73.100 ;
        RECT 21.700 72.800 22.600 73.100 ;
        RECT 25.400 73.100 25.700 74.900 ;
        RECT 26.200 74.800 26.600 74.900 ;
        RECT 27.000 74.800 27.400 75.600 ;
        RECT 27.800 74.200 28.100 75.900 ;
        RECT 30.200 74.400 30.600 75.200 ;
        RECT 30.900 74.200 31.200 75.900 ;
        RECT 31.800 75.800 32.200 75.900 ;
        RECT 32.600 75.800 33.000 76.600 ;
        RECT 31.800 75.100 32.100 75.800 ;
        RECT 33.400 75.100 33.800 79.900 ;
        RECT 35.000 75.700 35.400 79.900 ;
        RECT 37.200 78.200 37.600 79.900 ;
        RECT 36.600 77.900 37.600 78.200 ;
        RECT 39.400 77.900 39.800 79.900 ;
        RECT 41.500 77.900 42.100 79.900 ;
        RECT 36.600 77.500 37.000 77.900 ;
        RECT 39.400 77.600 39.700 77.900 ;
        RECT 38.300 77.300 40.100 77.600 ;
        RECT 41.400 77.500 41.800 77.900 ;
        RECT 38.300 77.200 38.700 77.300 ;
        RECT 39.700 77.200 40.100 77.300 ;
        RECT 36.600 76.500 37.000 76.600 ;
        RECT 38.900 76.500 39.300 76.600 ;
        RECT 36.600 76.200 39.300 76.500 ;
        RECT 39.600 76.500 40.700 76.800 ;
        RECT 39.600 75.900 39.900 76.500 ;
        RECT 40.300 76.400 40.700 76.500 ;
        RECT 41.500 76.600 42.200 77.000 ;
        RECT 41.500 76.100 41.800 76.600 ;
        RECT 37.500 75.700 39.900 75.900 ;
        RECT 35.000 75.600 39.900 75.700 ;
        RECT 40.600 75.800 41.800 76.100 ;
        RECT 35.000 75.500 37.900 75.600 ;
        RECT 35.000 75.400 37.800 75.500 ;
        RECT 38.200 75.100 38.600 75.200 ;
        RECT 31.800 74.800 33.800 75.100 ;
        RECT 27.800 73.800 28.200 74.200 ;
        RECT 29.400 74.100 29.800 74.200 ;
        RECT 30.900 74.100 32.200 74.200 ;
        RECT 32.600 74.100 33.000 74.200 ;
        RECT 29.400 73.800 30.200 74.100 ;
        RECT 30.900 73.800 33.000 74.100 ;
        RECT 26.200 73.100 26.600 73.200 ;
        RECT 27.800 73.100 28.100 73.800 ;
        RECT 29.800 73.600 30.200 73.800 ;
        RECT 21.700 71.100 22.100 72.800 ;
        RECT 25.400 71.100 25.800 73.100 ;
        RECT 26.200 72.800 28.100 73.100 ;
        RECT 26.100 72.400 26.500 72.800 ;
        RECT 27.800 72.100 28.100 72.800 ;
        RECT 28.600 72.400 29.000 73.200 ;
        RECT 29.500 73.100 31.300 73.300 ;
        RECT 31.800 73.100 32.100 73.800 ;
        RECT 33.400 73.100 33.800 74.800 ;
        RECT 36.100 74.800 38.600 75.100 ;
        RECT 36.100 74.700 36.500 74.800 ;
        RECT 37.400 74.700 37.800 74.800 ;
        RECT 36.900 74.200 37.300 74.300 ;
        RECT 40.600 74.200 40.900 75.800 ;
        RECT 43.800 75.600 44.200 79.900 ;
        RECT 42.100 75.300 44.200 75.600 ;
        RECT 44.600 77.500 45.000 79.500 ;
        RECT 44.600 75.800 44.900 77.500 ;
        RECT 46.700 76.400 47.100 79.900 ;
        RECT 46.700 76.100 47.500 76.400 ;
        RECT 52.300 76.300 52.700 79.900 ;
        RECT 44.600 75.500 46.500 75.800 ;
        RECT 42.100 75.200 42.500 75.300 ;
        RECT 42.900 74.900 43.300 75.000 ;
        RECT 41.400 74.600 43.300 74.900 ;
        RECT 41.400 74.500 41.800 74.600 ;
        RECT 34.200 73.400 34.600 74.200 ;
        RECT 35.400 73.900 40.900 74.200 ;
        RECT 35.400 73.800 36.200 73.900 ;
        RECT 29.400 73.000 31.400 73.100 ;
        RECT 27.800 71.100 28.200 72.100 ;
        RECT 29.400 71.100 29.800 73.000 ;
        RECT 31.000 71.100 31.400 73.000 ;
        RECT 31.800 71.100 32.200 73.100 ;
        RECT 32.900 72.800 33.800 73.100 ;
        RECT 32.900 71.100 33.300 72.800 ;
        RECT 35.000 71.100 35.400 73.500 ;
        RECT 37.500 72.800 37.800 73.900 ;
        RECT 40.300 73.800 40.700 73.900 ;
        RECT 43.800 73.600 44.200 75.300 ;
        RECT 44.600 74.400 45.000 75.200 ;
        RECT 45.400 74.400 45.800 75.200 ;
        RECT 46.200 74.500 46.500 75.500 ;
        RECT 46.200 74.100 46.900 74.500 ;
        RECT 47.200 74.200 47.500 76.100 ;
        RECT 51.800 75.900 52.700 76.300 ;
        RECT 53.400 75.900 53.800 79.900 ;
        RECT 54.200 76.200 54.600 79.900 ;
        RECT 55.800 76.200 56.200 79.900 ;
        RECT 54.200 75.900 56.200 76.200 ;
        RECT 47.800 75.100 48.200 75.600 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 47.800 74.800 49.800 75.100 ;
        RECT 51.900 74.200 52.200 75.900 ;
        RECT 52.600 74.800 53.000 75.600 ;
        RECT 53.500 75.200 53.800 75.900 ;
        RECT 56.600 75.600 57.000 79.900 ;
        RECT 58.700 77.900 59.300 79.900 ;
        RECT 61.000 77.900 61.400 79.900 ;
        RECT 63.200 78.200 63.600 79.900 ;
        RECT 63.200 77.900 64.200 78.200 ;
        RECT 59.000 77.500 59.400 77.900 ;
        RECT 61.100 77.600 61.400 77.900 ;
        RECT 60.700 77.300 62.500 77.600 ;
        RECT 63.800 77.500 64.200 77.900 ;
        RECT 60.700 77.200 61.100 77.300 ;
        RECT 62.100 77.200 62.500 77.300 ;
        RECT 58.200 77.000 58.900 77.200 ;
        RECT 58.200 76.800 59.300 77.000 ;
        RECT 58.600 76.600 59.300 76.800 ;
        RECT 59.000 76.100 59.300 76.600 ;
        RECT 60.100 76.500 61.200 76.800 ;
        RECT 60.100 76.400 60.500 76.500 ;
        RECT 59.000 75.800 60.200 76.100 ;
        RECT 55.400 75.200 55.800 75.400 ;
        RECT 56.600 75.300 58.700 75.600 ;
        RECT 53.400 74.900 54.600 75.200 ;
        RECT 55.400 74.900 56.200 75.200 ;
        RECT 53.400 74.800 53.800 74.900 ;
        RECT 54.200 74.800 54.600 74.900 ;
        RECT 55.800 74.800 56.200 74.900 ;
        RECT 46.200 73.900 46.700 74.100 ;
        RECT 42.300 73.300 44.200 73.600 ;
        RECT 42.300 73.200 42.700 73.300 ;
        RECT 36.600 72.100 37.000 72.500 ;
        RECT 37.400 72.400 37.800 72.800 ;
        RECT 38.300 72.700 38.700 72.800 ;
        RECT 38.300 72.400 39.700 72.700 ;
        RECT 39.400 72.100 39.700 72.400 ;
        RECT 41.400 72.100 41.800 72.500 ;
        RECT 36.600 71.800 37.600 72.100 ;
        RECT 37.200 71.100 37.600 71.800 ;
        RECT 39.400 71.100 39.800 72.100 ;
        RECT 41.400 71.800 42.100 72.100 ;
        RECT 41.500 71.100 42.100 71.800 ;
        RECT 43.800 71.100 44.200 73.300 ;
        RECT 44.600 73.600 46.700 73.900 ;
        RECT 47.200 73.800 48.200 74.200 ;
        RECT 51.800 73.800 52.200 74.200 ;
        RECT 44.600 72.500 44.900 73.600 ;
        RECT 47.200 73.500 47.500 73.800 ;
        RECT 47.100 73.300 47.500 73.500 ;
        RECT 46.700 73.000 47.500 73.300 ;
        RECT 49.400 73.100 49.800 73.200 ;
        RECT 51.000 73.100 51.400 73.200 ;
        RECT 51.900 73.100 52.200 73.800 ;
        RECT 53.400 73.100 53.800 73.200 ;
        RECT 54.300 73.100 54.600 74.800 ;
        RECT 55.000 73.800 55.400 74.600 ;
        RECT 44.600 71.500 45.000 72.500 ;
        RECT 46.700 71.500 47.100 73.000 ;
        RECT 49.400 72.800 51.400 73.100 ;
        RECT 51.800 72.800 53.800 73.100 ;
        RECT 51.000 72.400 51.400 72.800 ;
        RECT 51.900 72.100 52.200 72.800 ;
        RECT 53.500 72.400 53.900 72.800 ;
        RECT 51.800 71.100 52.200 72.100 ;
        RECT 54.200 71.100 54.600 73.100 ;
        RECT 56.600 73.600 57.000 75.300 ;
        RECT 58.300 75.200 58.700 75.300 ;
        RECT 57.500 74.900 57.900 75.000 ;
        RECT 57.500 74.600 59.400 74.900 ;
        RECT 59.000 74.500 59.400 74.600 ;
        RECT 59.900 74.200 60.200 75.800 ;
        RECT 60.900 75.900 61.200 76.500 ;
        RECT 61.500 76.500 61.900 76.600 ;
        RECT 63.800 76.500 64.200 76.600 ;
        RECT 61.500 76.200 64.200 76.500 ;
        RECT 60.900 75.700 63.300 75.900 ;
        RECT 65.400 75.700 65.800 79.900 ;
        RECT 67.000 76.400 67.400 79.900 ;
        RECT 60.900 75.600 65.800 75.700 ;
        RECT 62.900 75.500 65.800 75.600 ;
        RECT 63.000 75.400 65.800 75.500 ;
        RECT 66.900 75.900 67.400 76.400 ;
        RECT 68.600 76.200 69.000 79.900 ;
        RECT 67.700 75.900 69.000 76.200 ;
        RECT 69.400 76.200 69.800 79.900 ;
        RECT 71.000 76.400 71.400 79.900 ;
        RECT 69.400 75.900 70.700 76.200 ;
        RECT 71.000 75.900 71.500 76.400 ;
        RECT 73.900 76.200 74.300 79.900 ;
        RECT 74.600 76.800 75.000 77.200 ;
        RECT 74.700 76.200 75.000 76.800 ;
        RECT 73.900 75.900 74.400 76.200 ;
        RECT 74.700 75.900 75.400 76.200 ;
        RECT 62.200 75.100 62.600 75.200 ;
        RECT 62.200 74.800 64.700 75.100 ;
        RECT 64.300 74.700 64.700 74.800 ;
        RECT 63.500 74.200 63.900 74.300 ;
        RECT 66.900 74.200 67.200 75.900 ;
        RECT 67.700 74.900 68.000 75.900 ;
        RECT 67.500 74.500 68.000 74.900 ;
        RECT 59.900 73.900 65.400 74.200 ;
        RECT 60.100 73.800 60.500 73.900 ;
        RECT 56.600 73.300 58.500 73.600 ;
        RECT 56.600 71.100 57.000 73.300 ;
        RECT 58.100 73.200 58.500 73.300 ;
        RECT 63.000 72.800 63.300 73.900 ;
        RECT 64.600 73.800 65.400 73.900 ;
        RECT 66.900 73.800 67.400 74.200 ;
        RECT 62.100 72.700 62.500 72.800 ;
        RECT 59.000 72.100 59.400 72.500 ;
        RECT 61.100 72.400 62.500 72.700 ;
        RECT 63.000 72.400 63.400 72.800 ;
        RECT 61.100 72.100 61.400 72.400 ;
        RECT 63.800 72.100 64.200 72.500 ;
        RECT 58.700 71.800 59.400 72.100 ;
        RECT 58.700 71.100 59.300 71.800 ;
        RECT 61.000 71.100 61.400 72.100 ;
        RECT 63.200 71.800 64.200 72.100 ;
        RECT 63.200 71.100 63.600 71.800 ;
        RECT 65.400 71.100 65.800 73.500 ;
        RECT 66.900 73.100 67.200 73.800 ;
        RECT 67.700 73.700 68.000 74.500 ;
        RECT 68.500 75.100 69.000 75.200 ;
        RECT 69.400 75.100 69.900 75.200 ;
        RECT 68.500 74.800 69.900 75.100 ;
        RECT 68.500 74.400 68.900 74.800 ;
        RECT 69.500 74.400 69.900 74.800 ;
        RECT 70.400 74.900 70.700 75.900 ;
        RECT 70.400 74.500 70.900 74.900 ;
        RECT 70.400 73.700 70.700 74.500 ;
        RECT 71.200 74.200 71.500 75.900 ;
        RECT 74.100 75.200 74.400 75.900 ;
        RECT 75.000 75.800 75.400 75.900 ;
        RECT 75.800 75.800 76.200 76.600 ;
        RECT 73.400 74.400 73.800 75.200 ;
        RECT 74.100 74.800 74.600 75.200 ;
        RECT 75.000 75.100 75.300 75.800 ;
        RECT 76.600 75.100 77.000 79.900 ;
        RECT 78.200 75.700 78.600 79.900 ;
        RECT 80.400 78.200 80.800 79.900 ;
        RECT 79.800 77.900 80.800 78.200 ;
        RECT 82.600 77.900 83.000 79.900 ;
        RECT 84.700 77.900 85.300 79.900 ;
        RECT 79.800 77.500 80.200 77.900 ;
        RECT 82.600 77.600 82.900 77.900 ;
        RECT 81.500 77.300 83.300 77.600 ;
        RECT 84.600 77.500 85.000 77.900 ;
        RECT 81.500 77.200 81.900 77.300 ;
        RECT 82.900 77.200 83.300 77.300 ;
        RECT 79.800 76.500 80.200 76.600 ;
        RECT 82.100 76.500 82.500 76.600 ;
        RECT 79.800 76.200 82.500 76.500 ;
        RECT 82.800 76.500 83.900 76.800 ;
        RECT 82.800 75.900 83.100 76.500 ;
        RECT 83.500 76.400 83.900 76.500 ;
        RECT 84.700 76.600 85.400 77.000 ;
        RECT 84.700 76.100 85.000 76.600 ;
        RECT 80.700 75.700 83.100 75.900 ;
        RECT 78.200 75.600 83.100 75.700 ;
        RECT 83.800 75.800 85.000 76.100 ;
        RECT 78.200 75.500 81.100 75.600 ;
        RECT 78.200 75.400 81.000 75.500 ;
        RECT 81.400 75.100 81.800 75.200 ;
        RECT 75.000 74.800 77.000 75.100 ;
        RECT 74.100 74.200 74.400 74.800 ;
        RECT 71.000 74.100 71.500 74.200 ;
        RECT 72.600 74.100 73.000 74.200 ;
        RECT 71.000 73.800 73.400 74.100 ;
        RECT 74.100 73.800 75.400 74.200 ;
        RECT 67.700 73.400 69.000 73.700 ;
        RECT 66.900 72.800 67.400 73.100 ;
        RECT 67.000 71.100 67.400 72.800 ;
        RECT 68.600 71.100 69.000 73.400 ;
        RECT 69.400 73.400 70.700 73.700 ;
        RECT 69.400 71.100 69.800 73.400 ;
        RECT 71.200 73.100 71.500 73.800 ;
        RECT 73.000 73.600 73.400 73.800 ;
        RECT 72.700 73.100 74.500 73.300 ;
        RECT 75.000 73.100 75.300 73.800 ;
        RECT 76.600 73.100 77.000 74.800 ;
        RECT 79.300 74.800 81.800 75.100 ;
        RECT 79.300 74.700 79.700 74.800 ;
        RECT 80.100 74.200 80.500 74.300 ;
        RECT 83.800 74.200 84.100 75.800 ;
        RECT 87.000 75.600 87.400 79.900 ;
        RECT 87.800 76.200 88.200 79.900 ;
        RECT 89.400 79.600 91.400 79.900 ;
        RECT 89.400 76.200 89.800 79.600 ;
        RECT 87.800 75.900 89.800 76.200 ;
        RECT 90.200 75.900 90.600 79.300 ;
        RECT 91.000 75.900 91.400 79.600 ;
        RECT 90.200 75.600 90.500 75.900 ;
        RECT 85.300 75.300 87.400 75.600 ;
        RECT 85.300 75.200 85.700 75.300 ;
        RECT 86.100 74.900 86.500 75.000 ;
        RECT 84.600 74.600 86.500 74.900 ;
        RECT 84.600 74.500 85.000 74.600 ;
        RECT 77.400 73.400 77.800 74.200 ;
        RECT 78.600 73.900 84.100 74.200 ;
        RECT 78.600 73.800 79.400 73.900 ;
        RECT 80.600 73.800 81.000 73.900 ;
        RECT 83.500 73.800 83.900 73.900 ;
        RECT 71.000 72.800 71.500 73.100 ;
        RECT 72.600 73.000 74.600 73.100 ;
        RECT 71.000 71.100 71.400 72.800 ;
        RECT 72.600 71.100 73.000 73.000 ;
        RECT 74.200 71.100 74.600 73.000 ;
        RECT 75.000 71.100 75.400 73.100 ;
        RECT 76.100 72.800 77.000 73.100 ;
        RECT 76.100 71.100 76.500 72.800 ;
        RECT 78.200 71.100 78.600 73.500 ;
        RECT 80.700 72.800 81.000 73.800 ;
        RECT 87.000 73.600 87.400 75.300 ;
        RECT 88.200 75.200 88.600 75.400 ;
        RECT 89.500 75.300 90.500 75.600 ;
        RECT 89.500 75.200 89.800 75.300 ;
        RECT 87.800 74.900 88.600 75.200 ;
        RECT 87.800 74.800 88.200 74.900 ;
        RECT 89.400 74.800 89.800 75.200 ;
        RECT 91.000 74.800 91.400 75.600 ;
        RECT 88.600 73.800 89.000 74.600 ;
        RECT 85.500 73.300 87.400 73.600 ;
        RECT 85.500 73.200 85.900 73.300 ;
        RECT 79.800 72.100 80.200 72.500 ;
        RECT 80.600 72.400 81.000 72.800 ;
        RECT 81.500 72.700 81.900 72.800 ;
        RECT 81.500 72.400 82.900 72.700 ;
        RECT 82.600 72.100 82.900 72.400 ;
        RECT 84.600 72.100 85.000 72.500 ;
        RECT 79.800 71.800 80.800 72.100 ;
        RECT 80.400 71.100 80.800 71.800 ;
        RECT 82.600 71.100 83.000 72.100 ;
        RECT 84.600 71.800 85.300 72.100 ;
        RECT 84.700 71.100 85.300 71.800 ;
        RECT 87.000 71.100 87.400 73.300 ;
        RECT 89.500 73.100 89.800 74.800 ;
        RECT 90.100 74.400 90.500 74.800 ;
        RECT 90.200 74.200 90.500 74.400 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 91.800 73.400 92.200 74.200 ;
        RECT 92.600 73.100 93.000 79.900 ;
        RECT 93.400 75.800 93.800 76.600 ;
        RECT 94.200 75.800 94.600 76.600 ;
        RECT 95.000 73.100 95.400 79.900 ;
        RECT 97.400 75.100 97.800 79.900 ;
        RECT 101.000 76.800 101.400 77.200 ;
        RECT 98.200 75.800 98.600 76.600 ;
        RECT 101.000 76.200 101.300 76.800 ;
        RECT 101.700 76.200 102.100 79.900 ;
        RECT 104.600 77.900 105.000 79.900 ;
        RECT 100.600 75.900 101.300 76.200 ;
        RECT 101.600 75.900 102.100 76.200 ;
        RECT 100.600 75.800 101.000 75.900 ;
        RECT 100.600 75.100 100.900 75.800 ;
        RECT 97.400 74.800 100.900 75.100 ;
        RECT 95.800 73.400 96.200 74.200 ;
        RECT 96.600 73.400 97.000 74.200 ;
        RECT 89.300 71.100 90.100 73.100 ;
        RECT 92.600 72.800 93.500 73.100 ;
        RECT 93.100 72.200 93.500 72.800 ;
        RECT 92.600 71.800 93.500 72.200 ;
        RECT 93.100 71.100 93.500 71.800 ;
        RECT 94.500 72.800 95.400 73.100 ;
        RECT 97.400 73.100 97.800 74.800 ;
        RECT 101.600 74.200 101.900 75.900 ;
        RECT 104.700 75.800 105.000 77.900 ;
        RECT 106.200 75.900 106.600 79.900 ;
        RECT 104.700 75.500 105.900 75.800 ;
        RECT 102.200 74.400 102.600 75.200 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 100.600 73.800 101.900 74.200 ;
        RECT 103.000 74.100 103.400 74.200 ;
        RECT 102.600 73.800 103.400 74.100 ;
        RECT 103.800 73.800 104.200 74.600 ;
        RECT 104.700 74.400 105.000 74.800 ;
        RECT 104.700 74.100 105.200 74.400 ;
        RECT 104.800 74.000 105.200 74.100 ;
        RECT 105.600 73.800 105.900 75.500 ;
        RECT 106.300 75.200 106.600 75.900 ;
        RECT 106.200 74.800 106.600 75.200 ;
        RECT 100.700 73.100 101.000 73.800 ;
        RECT 102.600 73.600 103.000 73.800 ;
        RECT 105.600 73.700 106.000 73.800 ;
        RECT 104.500 73.500 106.000 73.700 ;
        RECT 103.900 73.400 106.000 73.500 ;
        RECT 101.500 73.100 103.300 73.300 ;
        RECT 103.900 73.200 104.800 73.400 ;
        RECT 103.900 73.100 104.200 73.200 ;
        RECT 106.300 73.100 106.600 74.800 ;
        RECT 107.000 73.400 107.400 74.200 ;
        RECT 97.400 72.800 98.300 73.100 ;
        RECT 94.500 71.100 94.900 72.800 ;
        RECT 97.900 71.100 98.300 72.800 ;
        RECT 100.600 71.100 101.000 73.100 ;
        RECT 101.400 73.000 103.400 73.100 ;
        RECT 101.400 71.100 101.800 73.000 ;
        RECT 103.000 71.100 103.400 73.000 ;
        RECT 103.800 71.100 104.200 73.100 ;
        RECT 105.900 72.600 106.600 73.100 ;
        RECT 107.800 73.100 108.200 79.900 ;
        RECT 108.600 75.800 109.000 76.600 ;
        RECT 109.700 76.300 110.100 79.900 ;
        RECT 112.100 76.300 112.500 79.900 ;
        RECT 116.100 76.400 116.500 79.900 ;
        RECT 118.200 77.500 118.600 79.500 ;
        RECT 109.700 75.900 110.600 76.300 ;
        RECT 112.100 75.900 113.000 76.300 ;
        RECT 109.400 74.800 109.800 75.600 ;
        RECT 110.200 74.200 110.500 75.900 ;
        RECT 112.600 75.800 113.000 75.900 ;
        RECT 115.700 76.100 116.500 76.400 ;
        RECT 111.000 75.100 111.400 75.200 ;
        RECT 111.800 75.100 112.200 75.600 ;
        RECT 111.000 74.800 112.200 75.100 ;
        RECT 112.600 74.200 112.900 75.800 ;
        RECT 115.000 74.800 115.400 75.600 ;
        RECT 115.700 74.200 116.000 76.100 ;
        RECT 118.300 75.800 118.600 77.500 ;
        RECT 116.700 75.500 118.600 75.800 ;
        RECT 116.700 74.500 117.000 75.500 ;
        RECT 108.600 74.100 109.000 74.200 ;
        RECT 110.200 74.100 110.600 74.200 ;
        RECT 108.600 73.800 110.600 74.100 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 115.000 73.800 116.000 74.200 ;
        RECT 116.300 74.100 117.000 74.500 ;
        RECT 117.400 74.400 117.800 75.200 ;
        RECT 118.200 74.400 118.600 75.200 ;
        RECT 119.800 75.100 120.200 79.900 ;
        RECT 120.600 75.800 121.000 76.600 ;
        RECT 121.700 76.300 122.100 79.900 ;
        RECT 125.700 76.400 126.100 79.900 ;
        RECT 128.600 79.600 130.600 79.900 ;
        RECT 127.800 77.500 128.200 79.500 ;
        RECT 121.700 75.900 122.600 76.300 ;
        RECT 125.300 76.100 126.100 76.400 ;
        RECT 121.400 75.100 121.800 75.600 ;
        RECT 119.800 74.800 121.800 75.100 ;
        RECT 122.200 75.100 122.500 75.900 ;
        RECT 123.000 75.100 123.400 75.200 ;
        RECT 122.200 74.800 123.400 75.100 ;
        RECT 123.800 75.100 124.200 75.200 ;
        RECT 124.600 75.100 125.000 75.600 ;
        RECT 123.800 74.800 125.000 75.100 ;
        RECT 107.800 72.800 108.700 73.100 ;
        RECT 105.900 72.200 106.300 72.600 ;
        RECT 108.300 72.200 108.700 72.800 ;
        RECT 105.900 71.800 106.600 72.200 ;
        RECT 108.300 71.800 109.000 72.200 ;
        RECT 110.200 72.100 110.500 73.800 ;
        RECT 111.000 73.100 111.400 73.200 ;
        RECT 111.800 73.100 112.200 73.200 ;
        RECT 111.000 72.800 112.200 73.100 ;
        RECT 111.000 72.400 111.400 72.800 ;
        RECT 112.600 72.100 112.900 73.800 ;
        RECT 115.700 73.500 116.000 73.800 ;
        RECT 116.500 73.900 117.000 74.100 ;
        RECT 116.500 73.600 118.600 73.900 ;
        RECT 115.700 73.300 116.100 73.500 ;
        RECT 113.400 72.400 113.800 73.200 ;
        RECT 115.700 73.000 116.500 73.300 ;
        RECT 116.100 72.200 116.500 73.000 ;
        RECT 118.300 72.500 118.600 73.600 ;
        RECT 119.000 73.400 119.400 74.200 ;
        RECT 119.800 73.100 120.200 74.800 ;
        RECT 122.200 74.200 122.500 74.800 ;
        RECT 125.300 74.200 125.600 76.100 ;
        RECT 127.900 75.800 128.200 77.500 ;
        RECT 128.600 75.900 129.000 79.600 ;
        RECT 129.400 75.900 129.800 79.300 ;
        RECT 130.200 76.200 130.600 79.600 ;
        RECT 131.800 76.200 132.200 79.900 ;
        RECT 130.200 75.900 132.200 76.200 ;
        RECT 132.600 77.500 133.000 79.500 ;
        RECT 126.300 75.500 128.200 75.800 ;
        RECT 129.500 75.600 129.800 75.900 ;
        RECT 132.600 75.800 132.900 77.500 ;
        RECT 134.700 76.400 135.100 79.900 ;
        RECT 138.200 77.900 138.600 79.900 ;
        RECT 134.700 76.100 135.500 76.400 ;
        RECT 126.300 74.500 126.600 75.500 ;
        RECT 122.200 73.800 122.600 74.200 ;
        RECT 124.600 73.800 125.600 74.200 ;
        RECT 125.900 74.100 126.600 74.500 ;
        RECT 127.000 74.400 127.400 75.200 ;
        RECT 127.800 74.400 128.200 75.200 ;
        RECT 128.600 74.800 129.000 75.600 ;
        RECT 129.500 75.300 130.500 75.600 ;
        RECT 132.600 75.500 134.500 75.800 ;
        RECT 130.200 75.200 130.500 75.300 ;
        RECT 131.400 75.200 131.800 75.400 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 131.400 74.900 132.200 75.200 ;
        RECT 131.800 74.800 132.200 74.900 ;
        RECT 129.500 74.400 129.900 74.800 ;
        RECT 129.500 74.200 129.800 74.400 ;
        RECT 119.800 72.800 120.700 73.100 ;
        RECT 105.900 71.100 106.300 71.800 ;
        RECT 108.300 71.100 108.700 71.800 ;
        RECT 110.200 71.100 110.600 72.100 ;
        RECT 112.600 71.100 113.000 72.100 ;
        RECT 115.800 71.800 116.500 72.200 ;
        RECT 116.100 71.500 116.500 71.800 ;
        RECT 118.200 71.500 118.600 72.500 ;
        RECT 120.300 71.100 120.700 72.800 ;
        RECT 122.200 72.100 122.500 73.800 ;
        RECT 125.300 73.500 125.600 73.800 ;
        RECT 126.100 73.900 126.600 74.100 ;
        RECT 126.100 73.600 128.200 73.900 ;
        RECT 129.400 73.800 129.800 74.200 ;
        RECT 125.300 73.300 125.700 73.500 ;
        RECT 123.000 72.400 123.400 73.200 ;
        RECT 125.300 73.000 126.100 73.300 ;
        RECT 122.200 71.100 122.600 72.100 ;
        RECT 125.700 71.500 126.100 73.000 ;
        RECT 127.900 72.500 128.200 73.600 ;
        RECT 130.200 73.100 130.500 74.800 ;
        RECT 131.000 73.800 131.400 74.600 ;
        RECT 131.800 74.200 132.100 74.800 ;
        RECT 132.600 74.400 133.000 75.200 ;
        RECT 133.400 74.400 133.800 75.200 ;
        RECT 134.200 74.500 134.500 75.500 ;
        RECT 135.200 75.200 135.500 76.100 ;
        RECT 138.300 75.800 138.600 77.900 ;
        RECT 139.800 75.900 140.200 79.900 ;
        RECT 135.000 74.800 135.500 75.200 ;
        RECT 135.800 75.100 136.200 75.600 ;
        RECT 138.300 75.500 139.500 75.800 ;
        RECT 136.600 75.100 137.000 75.200 ;
        RECT 135.800 74.800 137.000 75.100 ;
        RECT 138.200 74.800 138.600 75.200 ;
        RECT 131.800 73.800 132.200 74.200 ;
        RECT 134.200 74.100 134.900 74.500 ;
        RECT 135.200 74.200 135.500 74.800 ;
        RECT 134.200 73.900 134.700 74.100 ;
        RECT 132.600 73.600 134.700 73.900 ;
        RECT 135.200 73.800 136.200 74.200 ;
        RECT 137.400 73.800 137.800 74.600 ;
        RECT 138.300 74.400 138.600 74.800 ;
        RECT 138.300 74.100 138.800 74.400 ;
        RECT 138.400 74.000 138.800 74.100 ;
        RECT 139.200 73.800 139.500 75.500 ;
        RECT 139.900 75.200 140.200 75.900 ;
        RECT 139.800 74.800 140.200 75.200 ;
        RECT 127.800 71.500 128.200 72.500 ;
        RECT 129.900 72.200 130.700 73.100 ;
        RECT 129.400 71.800 130.700 72.200 ;
        RECT 129.900 71.100 130.700 71.800 ;
        RECT 132.600 72.500 132.900 73.600 ;
        RECT 135.200 73.500 135.500 73.800 ;
        RECT 139.200 73.700 139.600 73.800 ;
        RECT 138.100 73.500 139.600 73.700 ;
        RECT 135.100 73.300 135.500 73.500 ;
        RECT 134.700 73.000 135.500 73.300 ;
        RECT 137.500 73.400 139.600 73.500 ;
        RECT 137.500 73.200 138.400 73.400 ;
        RECT 137.500 73.100 137.800 73.200 ;
        RECT 139.900 73.100 140.200 74.800 ;
        RECT 140.600 73.400 141.000 74.200 ;
        RECT 132.600 71.500 133.000 72.500 ;
        RECT 134.700 71.500 135.100 73.000 ;
        RECT 137.400 71.100 137.800 73.100 ;
        RECT 139.500 72.600 140.200 73.100 ;
        RECT 141.400 73.100 141.800 79.900 ;
        RECT 142.200 75.800 142.600 76.600 ;
        RECT 143.000 76.200 143.400 79.900 ;
        RECT 144.600 76.400 145.000 79.900 ;
        RECT 143.000 75.900 144.300 76.200 ;
        RECT 144.600 75.900 145.100 76.400 ;
        RECT 144.000 74.900 144.300 75.900 ;
        RECT 144.000 74.500 144.500 74.900 ;
        RECT 144.000 73.700 144.300 74.500 ;
        RECT 144.800 74.200 145.100 75.900 ;
        RECT 147.800 75.600 148.200 79.900 ;
        RECT 149.900 77.900 150.500 79.900 ;
        RECT 152.200 77.900 152.600 79.900 ;
        RECT 154.400 78.200 154.800 79.900 ;
        RECT 154.400 77.900 155.400 78.200 ;
        RECT 150.200 77.500 150.600 77.900 ;
        RECT 152.300 77.600 152.600 77.900 ;
        RECT 151.900 77.300 153.700 77.600 ;
        RECT 155.000 77.500 155.400 77.900 ;
        RECT 151.900 77.200 152.300 77.300 ;
        RECT 153.300 77.200 153.700 77.300 ;
        RECT 149.800 76.600 150.500 77.000 ;
        RECT 150.200 76.100 150.500 76.600 ;
        RECT 151.300 76.500 152.400 76.800 ;
        RECT 151.300 76.400 151.700 76.500 ;
        RECT 150.200 75.800 151.400 76.100 ;
        RECT 147.800 75.300 149.900 75.600 ;
        RECT 144.600 74.100 145.100 74.200 ;
        RECT 147.000 74.100 147.400 74.200 ;
        RECT 144.600 73.800 147.400 74.100 ;
        RECT 143.000 73.400 144.300 73.700 ;
        RECT 141.400 72.800 142.300 73.100 ;
        RECT 139.500 71.100 139.900 72.600 ;
        RECT 141.900 72.200 142.300 72.800 ;
        RECT 141.400 71.800 142.300 72.200 ;
        RECT 141.900 71.100 142.300 71.800 ;
        RECT 143.000 71.100 143.400 73.400 ;
        RECT 144.800 73.100 145.100 73.800 ;
        RECT 144.600 72.800 145.100 73.100 ;
        RECT 147.800 73.600 148.200 75.300 ;
        RECT 149.500 75.200 149.900 75.300 ;
        RECT 151.100 75.100 151.400 75.800 ;
        RECT 152.100 75.900 152.400 76.500 ;
        RECT 152.700 76.500 153.100 76.600 ;
        RECT 155.000 76.500 155.400 76.600 ;
        RECT 152.700 76.200 155.400 76.500 ;
        RECT 152.100 75.700 154.500 75.900 ;
        RECT 156.600 75.700 157.000 79.900 ;
        RECT 157.400 75.800 157.800 77.200 ;
        RECT 152.100 75.600 157.000 75.700 ;
        RECT 154.100 75.500 157.000 75.600 ;
        RECT 154.200 75.400 157.000 75.500 ;
        RECT 151.800 75.100 152.200 75.200 ;
        RECT 148.700 74.900 149.100 75.000 ;
        RECT 148.700 74.600 150.600 74.900 ;
        RECT 151.000 74.800 152.200 75.100 ;
        RECT 153.400 75.100 153.800 75.200 ;
        RECT 158.200 75.100 158.600 79.900 ;
        RECT 159.800 76.200 160.200 79.900 ;
        RECT 161.400 76.200 161.800 79.900 ;
        RECT 159.800 75.900 161.800 76.200 ;
        RECT 162.200 75.900 162.600 79.900 ;
        RECT 163.800 76.400 164.200 79.900 ;
        RECT 163.700 75.900 164.200 76.400 ;
        RECT 165.400 76.200 165.800 79.900 ;
        RECT 164.500 75.900 165.800 76.200 ;
        RECT 167.500 76.200 167.900 79.900 ;
        RECT 168.200 76.800 168.600 77.200 ;
        RECT 168.300 76.200 168.600 76.800 ;
        RECT 167.500 75.900 168.000 76.200 ;
        RECT 168.300 75.900 169.000 76.200 ;
        RECT 160.200 75.200 160.600 75.400 ;
        RECT 162.200 75.200 162.500 75.900 ;
        RECT 159.800 75.100 160.600 75.200 ;
        RECT 153.400 74.800 155.900 75.100 ;
        RECT 150.200 74.500 150.600 74.600 ;
        RECT 151.100 74.200 151.400 74.800 ;
        RECT 154.200 74.700 154.600 74.800 ;
        RECT 155.500 74.700 155.900 74.800 ;
        RECT 158.200 74.900 160.600 75.100 ;
        RECT 161.400 74.900 162.600 75.200 ;
        RECT 158.200 74.800 160.200 74.900 ;
        RECT 161.400 74.800 161.800 74.900 ;
        RECT 162.200 74.800 162.600 74.900 ;
        RECT 154.700 74.200 155.100 74.300 ;
        RECT 151.100 74.100 156.600 74.200 ;
        RECT 157.400 74.100 157.800 74.200 ;
        RECT 151.100 73.900 157.800 74.100 ;
        RECT 151.300 73.800 151.700 73.900 ;
        RECT 147.800 73.300 149.700 73.600 ;
        RECT 144.600 71.100 145.000 72.800 ;
        RECT 147.800 71.100 148.200 73.300 ;
        RECT 149.300 73.200 149.700 73.300 ;
        RECT 154.200 72.800 154.500 73.900 ;
        RECT 155.800 73.800 157.800 73.900 ;
        RECT 153.300 72.700 153.700 72.800 ;
        RECT 150.200 72.100 150.600 72.500 ;
        RECT 152.300 72.400 153.700 72.700 ;
        RECT 154.200 72.400 154.600 72.800 ;
        RECT 152.300 72.100 152.600 72.400 ;
        RECT 155.000 72.100 155.400 72.500 ;
        RECT 149.900 71.800 150.600 72.100 ;
        RECT 149.900 71.100 150.500 71.800 ;
        RECT 152.200 71.100 152.600 72.100 ;
        RECT 154.400 71.800 155.400 72.100 ;
        RECT 154.400 71.100 154.800 71.800 ;
        RECT 156.600 71.100 157.000 73.500 ;
        RECT 158.200 73.100 158.600 74.800 ;
        RECT 160.600 73.800 161.000 74.600 ;
        RECT 157.700 72.800 158.600 73.100 ;
        RECT 161.400 73.100 161.700 74.800 ;
        RECT 163.700 74.200 164.000 75.900 ;
        RECT 164.500 74.900 164.800 75.900 ;
        RECT 167.700 75.200 168.000 75.900 ;
        RECT 168.600 75.800 169.000 75.900 ;
        RECT 169.400 75.800 169.800 76.600 ;
        RECT 164.300 74.500 164.800 74.900 ;
        RECT 166.200 75.100 166.600 75.200 ;
        RECT 167.000 75.100 167.400 75.200 ;
        RECT 166.200 74.800 167.400 75.100 ;
        RECT 163.700 73.800 164.200 74.200 ;
        RECT 157.700 71.100 158.100 72.800 ;
        RECT 161.400 71.100 161.800 73.100 ;
        RECT 162.200 72.800 162.600 73.200 ;
        RECT 163.700 73.100 164.000 73.800 ;
        RECT 164.500 73.700 164.800 74.500 ;
        RECT 167.000 74.400 167.400 74.800 ;
        RECT 167.700 74.800 168.200 75.200 ;
        RECT 168.600 75.100 168.900 75.800 ;
        RECT 170.200 75.100 170.600 79.900 ;
        RECT 171.800 75.700 172.200 79.900 ;
        RECT 174.000 78.200 174.400 79.900 ;
        RECT 173.400 77.900 174.400 78.200 ;
        RECT 176.200 77.900 176.600 79.900 ;
        RECT 178.300 77.900 178.900 79.900 ;
        RECT 173.400 77.500 173.800 77.900 ;
        RECT 176.200 77.600 176.500 77.900 ;
        RECT 175.100 77.300 176.900 77.600 ;
        RECT 178.200 77.500 178.600 77.900 ;
        RECT 175.100 77.200 175.500 77.300 ;
        RECT 176.500 77.200 176.900 77.300 ;
        RECT 173.400 76.500 173.800 76.600 ;
        RECT 175.700 76.500 176.100 76.600 ;
        RECT 173.400 76.200 176.100 76.500 ;
        RECT 176.400 76.500 177.500 76.800 ;
        RECT 176.400 75.900 176.700 76.500 ;
        RECT 177.100 76.400 177.500 76.500 ;
        RECT 178.300 76.600 179.000 77.000 ;
        RECT 178.300 76.100 178.600 76.600 ;
        RECT 174.300 75.700 176.700 75.900 ;
        RECT 171.800 75.600 176.700 75.700 ;
        RECT 177.400 75.800 178.600 76.100 ;
        RECT 171.800 75.500 174.700 75.600 ;
        RECT 171.800 75.400 174.600 75.500 ;
        RECT 175.000 75.100 175.400 75.200 ;
        RECT 168.600 74.800 170.600 75.100 ;
        RECT 167.700 74.200 168.000 74.800 ;
        RECT 166.200 74.100 166.600 74.200 ;
        RECT 166.200 73.800 167.000 74.100 ;
        RECT 167.700 73.800 169.000 74.200 ;
        RECT 164.500 73.400 165.800 73.700 ;
        RECT 166.600 73.600 167.000 73.800 ;
        RECT 163.700 72.800 164.200 73.100 ;
        RECT 162.100 72.400 162.500 72.800 ;
        RECT 163.800 71.100 164.200 72.800 ;
        RECT 165.400 71.100 165.800 73.400 ;
        RECT 166.300 73.100 168.100 73.300 ;
        RECT 168.600 73.100 168.900 73.800 ;
        RECT 170.200 73.100 170.600 74.800 ;
        RECT 172.900 74.800 175.400 75.100 ;
        RECT 172.900 74.700 173.300 74.800 ;
        RECT 174.200 74.700 174.600 74.800 ;
        RECT 173.700 74.200 174.100 74.300 ;
        RECT 177.400 74.200 177.700 75.800 ;
        RECT 180.600 75.600 181.000 79.900 ;
        RECT 181.800 76.800 182.200 77.200 ;
        RECT 181.800 76.200 182.100 76.800 ;
        RECT 182.500 76.200 182.900 79.900 ;
        RECT 181.400 75.900 182.100 76.200 ;
        RECT 182.400 75.900 182.900 76.200 ;
        RECT 184.600 77.500 185.000 79.500 ;
        RECT 181.400 75.800 181.800 75.900 ;
        RECT 178.900 75.300 181.000 75.600 ;
        RECT 178.900 75.200 179.300 75.300 ;
        RECT 179.700 74.900 180.100 75.000 ;
        RECT 178.200 74.600 180.100 74.900 ;
        RECT 178.200 74.500 178.600 74.600 ;
        RECT 171.000 73.400 171.400 74.200 ;
        RECT 172.200 73.900 177.700 74.200 ;
        RECT 172.200 73.800 173.000 73.900 ;
        RECT 166.200 73.000 168.200 73.100 ;
        RECT 166.200 71.100 166.600 73.000 ;
        RECT 167.800 71.100 168.200 73.000 ;
        RECT 168.600 71.100 169.000 73.100 ;
        RECT 169.700 72.800 170.600 73.100 ;
        RECT 169.700 71.100 170.100 72.800 ;
        RECT 171.800 71.100 172.200 73.500 ;
        RECT 174.300 72.800 174.600 73.900 ;
        RECT 177.100 73.800 177.500 73.900 ;
        RECT 180.600 73.600 181.000 75.300 ;
        RECT 182.400 74.200 182.700 75.900 ;
        RECT 184.600 75.800 184.900 77.500 ;
        RECT 186.700 76.400 187.100 79.900 ;
        RECT 189.400 77.500 189.800 79.500 ;
        RECT 186.700 76.100 187.500 76.400 ;
        RECT 184.600 75.500 186.500 75.800 ;
        RECT 183.000 74.400 183.400 75.200 ;
        RECT 184.600 74.400 185.000 75.200 ;
        RECT 185.400 74.400 185.800 75.200 ;
        RECT 186.200 74.500 186.500 75.500 ;
        RECT 181.400 73.800 182.700 74.200 ;
        RECT 183.800 74.100 184.200 74.200 ;
        RECT 183.400 73.800 184.200 74.100 ;
        RECT 186.200 74.100 186.900 74.500 ;
        RECT 187.200 74.200 187.500 76.100 ;
        RECT 189.400 75.800 189.700 77.500 ;
        RECT 191.500 76.400 191.900 79.900 ;
        RECT 195.500 77.200 195.900 79.900 ;
        RECT 195.000 76.800 195.900 77.200 ;
        RECT 196.200 76.800 196.600 77.200 ;
        RECT 191.500 76.100 192.300 76.400 ;
        RECT 187.800 75.100 188.200 75.600 ;
        RECT 189.400 75.500 191.300 75.800 ;
        RECT 188.600 75.100 189.000 75.200 ;
        RECT 187.800 74.800 189.000 75.100 ;
        RECT 189.400 74.400 189.800 75.200 ;
        RECT 190.200 74.400 190.600 75.200 ;
        RECT 191.000 74.500 191.300 75.500 ;
        RECT 186.200 73.900 186.700 74.100 ;
        RECT 179.100 73.300 181.000 73.600 ;
        RECT 179.100 73.200 179.500 73.300 ;
        RECT 173.400 72.100 173.800 72.500 ;
        RECT 174.200 72.400 174.600 72.800 ;
        RECT 175.100 72.700 175.500 72.800 ;
        RECT 175.100 72.400 176.500 72.700 ;
        RECT 176.200 72.100 176.500 72.400 ;
        RECT 178.200 72.100 178.600 72.500 ;
        RECT 173.400 71.800 174.400 72.100 ;
        RECT 174.000 71.100 174.400 71.800 ;
        RECT 176.200 71.100 176.600 72.100 ;
        RECT 178.200 71.800 178.900 72.100 ;
        RECT 178.300 71.100 178.900 71.800 ;
        RECT 180.600 71.100 181.000 73.300 ;
        RECT 181.500 73.200 181.800 73.800 ;
        RECT 183.400 73.600 183.800 73.800 ;
        RECT 184.600 73.600 186.700 73.900 ;
        RECT 187.200 73.800 188.200 74.200 ;
        RECT 191.000 74.100 191.700 74.500 ;
        RECT 192.000 74.200 192.300 76.100 ;
        RECT 195.500 76.200 195.900 76.800 ;
        RECT 196.300 76.200 196.600 76.800 ;
        RECT 195.500 75.900 196.000 76.200 ;
        RECT 196.300 75.900 197.000 76.200 ;
        RECT 192.600 74.800 193.000 75.600 ;
        RECT 194.200 75.100 194.600 75.200 ;
        RECT 195.000 75.100 195.400 75.200 ;
        RECT 194.200 74.800 195.400 75.100 ;
        RECT 195.000 74.400 195.400 74.800 ;
        RECT 195.700 74.200 196.000 75.900 ;
        RECT 196.600 75.800 197.000 75.900 ;
        RECT 197.400 75.800 197.800 76.600 ;
        RECT 196.600 75.100 196.900 75.800 ;
        RECT 198.200 75.100 198.600 79.900 ;
        RECT 196.600 74.800 198.600 75.100 ;
        RECT 191.000 73.900 191.500 74.100 ;
        RECT 181.400 71.100 181.800 73.200 ;
        RECT 182.300 73.100 184.100 73.300 ;
        RECT 182.200 73.000 184.200 73.100 ;
        RECT 182.200 71.100 182.600 73.000 ;
        RECT 183.800 71.100 184.200 73.000 ;
        RECT 184.600 72.500 184.900 73.600 ;
        RECT 187.200 73.500 187.500 73.800 ;
        RECT 187.100 73.300 187.500 73.500 ;
        RECT 186.700 73.000 187.500 73.300 ;
        RECT 189.400 73.600 191.500 73.900 ;
        RECT 192.000 73.800 193.000 74.200 ;
        RECT 193.400 74.100 193.800 74.200 ;
        RECT 194.200 74.100 194.600 74.200 ;
        RECT 193.400 73.800 195.000 74.100 ;
        RECT 195.700 73.800 197.000 74.200 ;
        RECT 184.600 71.500 185.000 72.500 ;
        RECT 186.700 71.500 187.100 73.000 ;
        RECT 189.400 72.500 189.700 73.600 ;
        RECT 192.000 73.500 192.300 73.800 ;
        RECT 194.600 73.600 195.000 73.800 ;
        RECT 191.900 73.300 192.300 73.500 ;
        RECT 191.500 73.000 192.300 73.300 ;
        RECT 194.300 73.100 196.100 73.300 ;
        RECT 196.600 73.100 196.900 73.800 ;
        RECT 198.200 73.100 198.600 74.800 ;
        RECT 199.000 73.400 199.400 74.200 ;
        RECT 199.800 73.400 200.200 74.200 ;
        RECT 194.200 73.000 196.200 73.100 ;
        RECT 189.400 71.500 189.800 72.500 ;
        RECT 191.500 72.200 191.900 73.000 ;
        RECT 191.000 71.800 191.900 72.200 ;
        RECT 191.500 71.500 191.900 71.800 ;
        RECT 194.200 71.100 194.600 73.000 ;
        RECT 195.800 71.100 196.200 73.000 ;
        RECT 196.600 71.100 197.000 73.100 ;
        RECT 197.700 72.800 198.600 73.100 ;
        RECT 200.600 73.100 201.000 79.900 ;
        RECT 203.800 79.600 205.800 79.900 ;
        RECT 201.400 75.800 201.800 76.600 ;
        RECT 203.800 75.900 204.200 79.600 ;
        RECT 204.600 75.800 205.000 79.300 ;
        RECT 205.400 76.200 205.800 79.600 ;
        RECT 207.000 76.200 207.400 79.900 ;
        RECT 205.400 75.900 207.400 76.200 ;
        RECT 207.800 77.500 208.200 79.500 ;
        RECT 204.700 75.600 205.000 75.800 ;
        RECT 207.800 75.800 208.100 77.500 ;
        RECT 209.900 76.400 210.300 79.900 ;
        RECT 209.900 76.100 210.700 76.400 ;
        RECT 203.800 74.800 204.200 75.600 ;
        RECT 204.700 75.300 205.700 75.600 ;
        RECT 207.800 75.500 209.700 75.800 ;
        RECT 205.400 75.200 205.700 75.300 ;
        RECT 206.600 75.200 207.000 75.400 ;
        RECT 205.400 74.800 205.800 75.200 ;
        RECT 206.600 74.900 207.400 75.200 ;
        RECT 207.000 74.800 207.400 74.900 ;
        RECT 204.700 74.400 205.100 74.800 ;
        RECT 204.700 74.200 205.000 74.400 ;
        RECT 202.200 74.100 202.600 74.200 ;
        RECT 204.600 74.100 205.000 74.200 ;
        RECT 202.200 73.800 205.000 74.100 ;
        RECT 205.400 73.100 205.700 74.800 ;
        RECT 206.200 73.800 206.600 74.600 ;
        RECT 207.800 74.400 208.200 75.200 ;
        RECT 208.600 74.400 209.000 75.200 ;
        RECT 209.400 74.500 209.700 75.500 ;
        RECT 209.400 74.100 210.100 74.500 ;
        RECT 210.400 74.200 210.700 76.100 ;
        RECT 211.000 75.100 211.400 75.600 ;
        RECT 211.800 75.100 212.200 75.200 ;
        RECT 211.000 74.800 212.200 75.100 ;
        RECT 209.400 73.900 209.900 74.100 ;
        RECT 207.800 73.600 209.900 73.900 ;
        RECT 210.400 73.800 211.400 74.200 ;
        RECT 200.600 72.800 201.500 73.100 ;
        RECT 197.700 71.100 198.100 72.800 ;
        RECT 201.100 71.100 201.500 72.800 ;
        RECT 205.100 71.100 205.900 73.100 ;
        RECT 207.800 72.500 208.100 73.600 ;
        RECT 210.400 73.500 210.700 73.800 ;
        RECT 210.300 73.300 210.700 73.500 ;
        RECT 212.600 73.400 213.000 74.200 ;
        RECT 209.900 73.000 210.700 73.300 ;
        RECT 213.400 73.100 213.800 79.900 ;
        RECT 214.200 75.800 214.600 76.600 ;
        RECT 215.000 76.100 215.400 76.200 ;
        RECT 215.800 76.100 216.200 79.900 ;
        RECT 215.000 75.800 216.200 76.100 ;
        RECT 215.000 73.400 215.400 74.200 ;
        RECT 215.800 73.100 216.200 75.800 ;
        RECT 216.600 75.800 217.000 76.600 ;
        RECT 218.700 76.200 219.100 79.900 ;
        RECT 219.400 76.800 219.800 77.200 ;
        RECT 219.500 76.200 219.800 76.800 ;
        RECT 222.500 76.400 222.900 79.900 ;
        RECT 224.600 77.500 225.000 79.500 ;
        RECT 218.700 75.900 219.200 76.200 ;
        RECT 219.500 75.900 220.200 76.200 ;
        RECT 216.600 75.100 216.900 75.800 ;
        RECT 218.200 75.100 218.600 75.200 ;
        RECT 216.600 74.800 218.600 75.100 ;
        RECT 218.200 74.400 218.600 74.800 ;
        RECT 218.900 74.200 219.200 75.900 ;
        RECT 219.800 75.800 220.200 75.900 ;
        RECT 222.100 76.100 222.900 76.400 ;
        RECT 219.800 75.100 220.200 75.200 ;
        RECT 221.400 75.100 221.800 75.600 ;
        RECT 219.800 74.800 221.800 75.100 ;
        RECT 222.100 74.200 222.400 76.100 ;
        RECT 224.700 75.800 225.000 77.500 ;
        RECT 223.100 75.500 225.000 75.800 ;
        RECT 225.400 75.600 225.800 79.900 ;
        RECT 227.500 77.900 228.100 79.900 ;
        RECT 229.800 77.900 230.200 79.900 ;
        RECT 232.000 78.200 232.400 79.900 ;
        RECT 232.000 77.900 233.000 78.200 ;
        RECT 227.800 77.500 228.200 77.900 ;
        RECT 229.900 77.600 230.200 77.900 ;
        RECT 229.500 77.300 231.300 77.600 ;
        RECT 232.600 77.500 233.000 77.900 ;
        RECT 229.500 77.200 229.900 77.300 ;
        RECT 230.900 77.200 231.300 77.300 ;
        RECT 227.400 76.600 228.100 77.000 ;
        RECT 227.800 76.100 228.100 76.600 ;
        RECT 228.900 76.500 230.000 76.800 ;
        RECT 228.900 76.400 229.300 76.500 ;
        RECT 227.800 75.800 229.000 76.100 ;
        RECT 223.100 74.500 223.400 75.500 ;
        RECT 225.400 75.300 227.500 75.600 ;
        RECT 217.400 74.100 217.800 74.200 ;
        RECT 217.400 73.800 218.200 74.100 ;
        RECT 218.900 73.800 220.200 74.200 ;
        RECT 220.600 74.100 221.000 74.200 ;
        RECT 221.400 74.100 222.400 74.200 ;
        RECT 222.700 74.100 223.400 74.500 ;
        RECT 223.800 74.400 224.200 75.200 ;
        RECT 224.600 74.400 225.000 75.200 ;
        RECT 220.600 73.800 222.400 74.100 ;
        RECT 217.800 73.600 218.200 73.800 ;
        RECT 217.500 73.100 219.300 73.300 ;
        RECT 219.800 73.100 220.100 73.800 ;
        RECT 222.100 73.500 222.400 73.800 ;
        RECT 222.900 73.900 223.400 74.100 ;
        RECT 222.900 73.600 225.000 73.900 ;
        RECT 222.100 73.300 222.500 73.500 ;
        RECT 207.800 71.500 208.200 72.500 ;
        RECT 209.900 72.200 210.300 73.000 ;
        RECT 213.400 72.800 214.300 73.100 ;
        RECT 215.800 72.800 216.700 73.100 ;
        RECT 213.900 72.200 214.300 72.800 ;
        RECT 209.400 71.800 210.300 72.200 ;
        RECT 213.400 71.800 214.300 72.200 ;
        RECT 209.900 71.500 210.300 71.800 ;
        RECT 213.900 71.100 214.300 71.800 ;
        RECT 216.300 71.100 216.700 72.800 ;
        RECT 217.400 73.000 219.400 73.100 ;
        RECT 217.400 71.100 217.800 73.000 ;
        RECT 219.000 71.100 219.400 73.000 ;
        RECT 219.800 71.100 220.200 73.100 ;
        RECT 222.100 73.000 222.900 73.300 ;
        RECT 222.500 71.500 222.900 73.000 ;
        RECT 224.700 72.500 225.000 73.600 ;
        RECT 224.600 71.500 225.000 72.500 ;
        RECT 225.400 73.600 225.800 75.300 ;
        RECT 227.100 75.200 227.500 75.300 ;
        RECT 226.300 74.900 226.700 75.000 ;
        RECT 226.300 74.600 228.200 74.900 ;
        RECT 227.800 74.500 228.200 74.600 ;
        RECT 228.700 74.200 229.000 75.800 ;
        RECT 229.700 75.900 230.000 76.500 ;
        RECT 230.300 76.500 230.700 76.600 ;
        RECT 232.600 76.500 233.000 76.600 ;
        RECT 230.300 76.200 233.000 76.500 ;
        RECT 229.700 75.700 232.100 75.900 ;
        RECT 234.200 75.700 234.600 79.900 ;
        RECT 229.700 75.600 234.600 75.700 ;
        RECT 231.700 75.500 234.600 75.600 ;
        RECT 231.800 75.400 234.600 75.500 ;
        RECT 235.800 75.600 236.200 79.900 ;
        RECT 237.400 75.600 237.800 79.900 ;
        RECT 239.000 75.600 239.400 79.900 ;
        RECT 240.600 75.600 241.000 79.900 ;
        RECT 243.500 76.300 243.900 79.900 ;
        RECT 243.000 75.900 243.900 76.300 ;
        RECT 244.600 75.900 245.000 79.900 ;
        RECT 245.400 76.200 245.800 79.900 ;
        RECT 247.000 76.200 247.400 79.900 ;
        RECT 248.200 76.800 248.600 77.200 ;
        RECT 248.200 76.200 248.500 76.800 ;
        RECT 248.900 76.200 249.300 79.900 ;
        RECT 245.400 75.900 247.400 76.200 ;
        RECT 247.800 75.900 248.500 76.200 ;
        RECT 248.800 75.900 249.300 76.200 ;
        RECT 235.800 75.200 236.700 75.600 ;
        RECT 237.400 75.200 238.500 75.600 ;
        RECT 239.000 75.200 240.100 75.600 ;
        RECT 240.600 75.200 241.800 75.600 ;
        RECT 229.400 75.100 229.800 75.200 ;
        RECT 231.000 75.100 231.400 75.200 ;
        RECT 229.400 74.800 233.500 75.100 ;
        RECT 233.100 74.700 233.500 74.800 ;
        RECT 236.300 74.500 236.700 75.200 ;
        RECT 238.100 74.500 238.500 75.200 ;
        RECT 239.700 74.500 240.100 75.200 ;
        RECT 232.300 74.200 232.700 74.300 ;
        RECT 228.700 73.900 234.200 74.200 ;
        RECT 228.900 73.800 229.300 73.900 ;
        RECT 225.400 73.300 227.300 73.600 ;
        RECT 225.400 71.100 225.800 73.300 ;
        RECT 226.900 73.200 227.300 73.300 ;
        RECT 231.800 73.200 232.100 73.900 ;
        RECT 233.400 73.800 234.200 73.900 ;
        RECT 235.000 74.100 235.900 74.500 ;
        RECT 236.300 74.100 237.600 74.500 ;
        RECT 238.100 74.100 239.300 74.500 ;
        RECT 239.700 74.100 241.000 74.500 ;
        RECT 235.000 73.800 235.400 74.100 ;
        RECT 236.300 73.800 236.700 74.100 ;
        RECT 238.100 73.800 238.500 74.100 ;
        RECT 239.700 73.800 240.100 74.100 ;
        RECT 241.400 73.800 241.800 75.200 ;
        RECT 243.100 74.200 243.400 75.900 ;
        RECT 243.800 74.800 244.200 75.600 ;
        RECT 244.700 75.200 245.000 75.900 ;
        RECT 247.800 75.800 248.200 75.900 ;
        RECT 246.600 75.200 247.000 75.400 ;
        RECT 244.600 74.900 245.800 75.200 ;
        RECT 246.600 74.900 247.400 75.200 ;
        RECT 244.600 74.800 245.000 74.900 ;
        RECT 243.000 73.800 243.400 74.200 ;
        RECT 230.900 72.700 231.300 72.800 ;
        RECT 227.800 72.100 228.200 72.500 ;
        RECT 229.900 72.400 231.300 72.700 ;
        RECT 231.800 72.400 232.200 73.200 ;
        RECT 229.900 72.100 230.200 72.400 ;
        RECT 232.600 72.100 233.000 72.500 ;
        RECT 227.500 71.800 228.200 72.100 ;
        RECT 227.500 71.100 228.100 71.800 ;
        RECT 229.800 71.100 230.200 72.100 ;
        RECT 232.000 71.800 233.000 72.100 ;
        RECT 232.000 71.100 232.400 71.800 ;
        RECT 234.200 71.100 234.600 73.500 ;
        RECT 235.800 73.400 236.700 73.800 ;
        RECT 237.400 73.400 238.500 73.800 ;
        RECT 239.000 73.400 240.100 73.800 ;
        RECT 240.600 73.400 241.800 73.800 ;
        RECT 235.800 71.100 236.200 73.400 ;
        RECT 237.400 71.100 237.800 73.400 ;
        RECT 239.000 71.100 239.400 73.400 ;
        RECT 240.600 71.100 241.000 73.400 ;
        RECT 242.200 72.400 242.600 73.200 ;
        RECT 243.100 73.100 243.400 73.800 ;
        RECT 244.600 73.100 245.000 73.200 ;
        RECT 245.500 73.100 245.800 74.900 ;
        RECT 247.000 74.800 247.400 74.900 ;
        RECT 246.200 73.800 246.600 74.600 ;
        RECT 248.800 74.200 249.100 75.900 ;
        RECT 249.400 75.100 249.800 75.200 ;
        RECT 251.800 75.100 252.200 75.200 ;
        RECT 249.400 74.800 252.200 75.100 ;
        RECT 249.400 74.400 249.800 74.800 ;
        RECT 247.800 73.800 249.100 74.200 ;
        RECT 250.200 74.100 250.600 74.200 ;
        RECT 249.800 73.800 250.600 74.100 ;
        RECT 247.900 73.100 248.200 73.800 ;
        RECT 249.800 73.600 250.200 73.800 ;
        RECT 248.700 73.100 250.500 73.300 ;
        RECT 243.000 72.800 245.000 73.100 ;
        RECT 243.100 72.100 243.400 72.800 ;
        RECT 244.700 72.400 245.100 72.800 ;
        RECT 243.000 71.100 243.400 72.100 ;
        RECT 245.400 71.100 245.800 73.100 ;
        RECT 247.800 71.100 248.200 73.100 ;
        RECT 248.600 73.000 250.600 73.100 ;
        RECT 248.600 71.100 249.000 73.000 ;
        RECT 250.200 71.100 250.600 73.000 ;
        RECT 1.900 68.200 2.300 69.900 ;
        RECT 1.400 67.900 2.300 68.200 ;
        RECT 3.000 67.900 3.400 69.900 ;
        RECT 3.800 68.000 4.200 69.900 ;
        RECT 5.400 68.000 5.800 69.900 ;
        RECT 8.100 68.000 8.500 69.500 ;
        RECT 10.200 68.500 10.600 69.500 ;
        RECT 3.800 67.900 5.800 68.000 ;
        RECT 0.600 66.800 1.000 67.600 ;
        RECT 1.400 66.100 1.800 67.900 ;
        RECT 3.100 67.200 3.400 67.900 ;
        RECT 3.900 67.700 5.700 67.900 ;
        RECT 7.700 67.700 8.500 68.000 ;
        RECT 7.700 67.500 8.100 67.700 ;
        RECT 5.000 67.200 5.400 67.400 ;
        RECT 7.700 67.200 8.000 67.500 ;
        RECT 10.300 67.400 10.600 68.500 ;
        RECT 11.000 67.500 11.400 69.900 ;
        RECT 13.200 69.200 13.600 69.900 ;
        RECT 12.600 68.900 13.600 69.200 ;
        RECT 15.400 68.900 15.800 69.900 ;
        RECT 17.500 69.200 18.100 69.900 ;
        RECT 17.400 68.900 18.100 69.200 ;
        RECT 12.600 68.500 13.000 68.900 ;
        RECT 15.400 68.600 15.700 68.900 ;
        RECT 13.400 68.200 13.800 68.600 ;
        RECT 14.300 68.300 15.700 68.600 ;
        RECT 17.400 68.500 17.800 68.900 ;
        RECT 14.300 68.200 14.700 68.300 ;
        RECT 3.000 66.800 4.300 67.200 ;
        RECT 5.000 66.900 5.800 67.200 ;
        RECT 5.400 66.800 5.800 66.900 ;
        RECT 7.000 66.800 8.000 67.200 ;
        RECT 8.500 67.100 10.600 67.400 ;
        RECT 11.400 67.100 12.200 67.200 ;
        RECT 13.500 67.100 13.800 68.200 ;
        RECT 18.300 67.700 18.700 67.800 ;
        RECT 19.800 67.700 20.200 69.900 ;
        RECT 18.300 67.400 20.200 67.700 ;
        RECT 20.600 67.500 21.000 69.900 ;
        RECT 22.800 69.200 23.200 69.900 ;
        RECT 22.200 68.900 23.200 69.200 ;
        RECT 25.000 68.900 25.400 69.900 ;
        RECT 27.100 69.200 27.700 69.900 ;
        RECT 27.000 68.900 27.700 69.200 ;
        RECT 22.200 68.500 22.600 68.900 ;
        RECT 25.000 68.600 25.300 68.900 ;
        RECT 23.000 68.200 23.400 68.600 ;
        RECT 23.900 68.300 25.300 68.600 ;
        RECT 27.000 68.500 27.400 68.900 ;
        RECT 23.900 68.200 24.300 68.300 ;
        RECT 15.000 67.100 15.400 67.200 ;
        RECT 16.300 67.100 16.700 67.200 ;
        RECT 8.500 66.900 9.000 67.100 ;
        RECT 1.400 65.800 3.300 66.100 ;
        RECT 1.400 61.100 1.800 65.800 ;
        RECT 3.000 65.200 3.300 65.800 ;
        RECT 2.200 64.400 2.600 65.200 ;
        RECT 3.000 65.100 3.400 65.200 ;
        RECT 4.000 65.100 4.300 66.800 ;
        RECT 4.600 65.800 5.000 66.600 ;
        RECT 7.700 66.200 8.000 66.800 ;
        RECT 8.300 66.500 9.000 66.900 ;
        RECT 11.400 66.800 16.900 67.100 ;
        RECT 12.900 66.700 13.300 66.800 ;
        RECT 6.200 66.100 6.600 66.200 ;
        RECT 7.000 66.100 7.400 66.200 ;
        RECT 6.200 65.800 7.400 66.100 ;
        RECT 7.000 65.400 7.400 65.800 ;
        RECT 7.700 65.800 8.200 66.200 ;
        RECT 3.000 64.800 3.700 65.100 ;
        RECT 4.000 64.800 4.500 65.100 ;
        RECT 3.400 64.200 3.700 64.800 ;
        RECT 3.400 63.800 3.800 64.200 ;
        RECT 4.100 61.100 4.500 64.800 ;
        RECT 7.700 64.900 8.000 65.800 ;
        RECT 8.700 65.500 9.000 66.500 ;
        RECT 9.400 65.800 9.800 66.600 ;
        RECT 10.200 65.800 10.600 66.600 ;
        RECT 12.100 66.200 12.500 66.300 ;
        RECT 12.100 65.900 14.600 66.200 ;
        RECT 14.200 65.800 14.600 65.900 ;
        RECT 11.000 65.500 13.800 65.600 ;
        RECT 8.700 65.200 10.600 65.500 ;
        RECT 7.700 64.600 8.500 64.900 ;
        RECT 8.100 61.100 8.500 64.600 ;
        RECT 10.300 63.500 10.600 65.200 ;
        RECT 10.200 61.500 10.600 63.500 ;
        RECT 11.000 65.400 13.900 65.500 ;
        RECT 11.000 65.300 15.900 65.400 ;
        RECT 11.000 61.100 11.400 65.300 ;
        RECT 13.500 65.100 15.900 65.300 ;
        RECT 12.600 64.500 15.300 64.800 ;
        RECT 12.600 64.400 13.000 64.500 ;
        RECT 14.900 64.400 15.300 64.500 ;
        RECT 15.600 64.500 15.900 65.100 ;
        RECT 16.600 65.200 16.900 66.800 ;
        RECT 17.400 66.400 17.800 66.500 ;
        RECT 17.400 66.100 19.300 66.400 ;
        RECT 18.900 66.000 19.300 66.100 ;
        RECT 18.100 65.700 18.500 65.800 ;
        RECT 19.800 65.700 20.200 67.400 ;
        RECT 21.000 67.100 21.800 67.200 ;
        RECT 23.100 67.100 23.400 68.200 ;
        RECT 27.900 67.700 28.300 67.800 ;
        RECT 29.400 67.700 29.800 69.900 ;
        RECT 27.900 67.400 29.800 67.700 ;
        RECT 25.900 67.100 26.300 67.200 ;
        RECT 21.000 66.800 26.500 67.100 ;
        RECT 22.500 66.700 22.900 66.800 ;
        RECT 21.700 66.200 22.100 66.300 ;
        RECT 26.200 66.200 26.500 66.800 ;
        RECT 27.000 66.400 27.400 66.500 ;
        RECT 21.700 66.100 24.200 66.200 ;
        RECT 25.400 66.100 25.800 66.200 ;
        RECT 21.700 65.900 25.800 66.100 ;
        RECT 23.800 65.800 25.800 65.900 ;
        RECT 26.200 65.800 26.600 66.200 ;
        RECT 27.000 66.100 28.900 66.400 ;
        RECT 28.500 66.000 28.900 66.100 ;
        RECT 18.100 65.400 20.200 65.700 ;
        RECT 16.600 64.900 17.800 65.200 ;
        RECT 16.300 64.500 16.700 64.600 ;
        RECT 15.600 64.200 16.700 64.500 ;
        RECT 17.500 64.400 17.800 64.900 ;
        RECT 17.500 64.000 18.200 64.400 ;
        RECT 14.300 63.700 14.700 63.800 ;
        RECT 15.700 63.700 16.100 63.800 ;
        RECT 12.600 63.100 13.000 63.500 ;
        RECT 14.300 63.400 16.100 63.700 ;
        RECT 15.400 63.100 15.700 63.400 ;
        RECT 17.400 63.100 17.800 63.500 ;
        RECT 12.600 62.800 13.600 63.100 ;
        RECT 13.200 61.100 13.600 62.800 ;
        RECT 15.400 61.100 15.800 63.100 ;
        RECT 17.500 61.100 18.100 63.100 ;
        RECT 19.800 61.100 20.200 65.400 ;
        RECT 20.600 65.500 23.400 65.600 ;
        RECT 20.600 65.400 23.500 65.500 ;
        RECT 20.600 65.300 25.500 65.400 ;
        RECT 20.600 61.100 21.000 65.300 ;
        RECT 23.100 65.100 25.500 65.300 ;
        RECT 22.200 64.500 24.900 64.800 ;
        RECT 22.200 64.400 22.600 64.500 ;
        RECT 24.500 64.400 24.900 64.500 ;
        RECT 25.200 64.500 25.500 65.100 ;
        RECT 26.200 65.200 26.500 65.800 ;
        RECT 27.700 65.700 28.100 65.800 ;
        RECT 29.400 65.700 29.800 67.400 ;
        RECT 30.200 68.500 30.600 69.500 ;
        RECT 30.200 67.400 30.500 68.500 ;
        RECT 32.300 68.000 32.700 69.500 ;
        RECT 35.000 68.500 35.400 69.500 ;
        RECT 32.300 67.700 33.100 68.000 ;
        RECT 32.700 67.500 33.100 67.700 ;
        RECT 30.200 67.100 32.300 67.400 ;
        RECT 31.800 66.900 32.300 67.100 ;
        RECT 32.800 67.200 33.100 67.500 ;
        RECT 35.000 67.400 35.300 68.500 ;
        RECT 37.100 68.000 37.500 69.500 ;
        RECT 41.700 68.000 42.100 69.500 ;
        RECT 43.800 68.500 44.200 69.500 ;
        RECT 37.100 67.700 37.900 68.000 ;
        RECT 37.500 67.500 37.900 67.700 ;
        RECT 30.200 65.800 30.600 66.600 ;
        RECT 31.000 65.800 31.400 66.600 ;
        RECT 31.800 66.500 32.500 66.900 ;
        RECT 32.800 66.800 33.800 67.200 ;
        RECT 35.000 67.100 37.100 67.400 ;
        RECT 36.600 66.900 37.100 67.100 ;
        RECT 37.600 67.200 37.900 67.500 ;
        RECT 41.300 67.700 42.100 68.000 ;
        RECT 41.300 67.500 41.700 67.700 ;
        RECT 41.300 67.200 41.600 67.500 ;
        RECT 43.900 67.400 44.200 68.500 ;
        RECT 46.500 68.000 46.900 69.500 ;
        RECT 48.600 68.500 49.000 69.500 ;
        RECT 37.600 67.100 38.600 67.200 ;
        RECT 39.800 67.100 40.200 67.200 ;
        RECT 27.700 65.400 29.800 65.700 ;
        RECT 31.800 65.500 32.100 66.500 ;
        RECT 26.200 64.900 27.400 65.200 ;
        RECT 25.900 64.500 26.300 64.600 ;
        RECT 25.200 64.200 26.300 64.500 ;
        RECT 27.100 64.400 27.400 64.900 ;
        RECT 27.100 64.000 27.800 64.400 ;
        RECT 23.900 63.700 24.300 63.800 ;
        RECT 25.300 63.700 25.700 63.800 ;
        RECT 22.200 63.100 22.600 63.500 ;
        RECT 23.900 63.400 25.700 63.700 ;
        RECT 25.000 63.100 25.300 63.400 ;
        RECT 27.000 63.100 27.400 63.500 ;
        RECT 22.200 62.800 23.200 63.100 ;
        RECT 22.800 61.100 23.200 62.800 ;
        RECT 25.000 61.100 25.400 63.100 ;
        RECT 27.100 61.100 27.700 63.100 ;
        RECT 29.400 61.100 29.800 65.400 ;
        RECT 30.200 65.200 32.100 65.500 ;
        RECT 30.200 63.500 30.500 65.200 ;
        RECT 32.800 64.900 33.100 66.800 ;
        RECT 33.400 66.100 33.800 66.200 ;
        RECT 34.200 66.100 34.600 66.200 ;
        RECT 33.400 65.800 34.600 66.100 ;
        RECT 35.000 65.800 35.400 66.600 ;
        RECT 35.800 65.800 36.200 66.600 ;
        RECT 36.600 66.500 37.300 66.900 ;
        RECT 37.600 66.800 40.200 67.100 ;
        RECT 40.600 66.800 41.600 67.200 ;
        RECT 42.100 67.100 44.200 67.400 ;
        RECT 46.100 67.700 46.900 68.000 ;
        RECT 46.100 67.500 46.500 67.700 ;
        RECT 46.100 67.200 46.400 67.500 ;
        RECT 48.700 67.400 49.000 68.500 ;
        RECT 52.300 67.900 53.100 69.900 ;
        RECT 56.500 67.900 57.300 69.900 ;
        RECT 60.300 68.200 60.700 69.900 ;
        RECT 59.800 67.900 60.700 68.200 ;
        RECT 61.400 68.000 61.800 69.900 ;
        RECT 63.000 68.000 63.400 69.900 ;
        RECT 61.400 67.900 63.400 68.000 ;
        RECT 63.800 67.900 64.200 69.900 ;
        RECT 65.900 67.900 66.700 69.900 ;
        RECT 69.900 68.200 70.300 69.900 ;
        RECT 69.400 67.900 70.300 68.200 ;
        RECT 72.900 68.000 73.300 69.500 ;
        RECT 75.000 68.500 75.400 69.500 ;
        RECT 42.100 66.900 42.600 67.100 ;
        RECT 33.400 65.400 33.800 65.800 ;
        RECT 36.600 65.500 36.900 66.500 ;
        RECT 32.300 64.600 33.100 64.900 ;
        RECT 35.000 65.200 36.900 65.500 ;
        RECT 30.200 61.500 30.600 63.500 ;
        RECT 32.300 61.100 32.700 64.600 ;
        RECT 35.000 63.500 35.300 65.200 ;
        RECT 37.600 64.900 37.900 66.800 ;
        RECT 41.300 66.200 41.600 66.800 ;
        RECT 41.900 66.500 42.600 66.900 ;
        RECT 45.400 66.800 46.400 67.200 ;
        RECT 46.900 67.100 49.000 67.400 ;
        RECT 46.900 66.900 47.400 67.100 ;
        RECT 38.200 65.400 38.600 66.200 ;
        RECT 40.600 65.400 41.000 66.200 ;
        RECT 41.300 65.800 41.800 66.200 ;
        RECT 37.100 64.600 37.900 64.900 ;
        RECT 41.300 64.900 41.600 65.800 ;
        RECT 42.300 65.500 42.600 66.500 ;
        RECT 43.000 65.800 43.400 66.600 ;
        RECT 43.800 66.100 44.200 66.600 ;
        RECT 46.100 66.200 46.400 66.800 ;
        RECT 46.700 66.500 47.400 66.900 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 51.900 66.600 52.200 66.800 ;
        RECT 44.600 66.100 45.000 66.200 ;
        RECT 43.800 65.800 45.000 66.100 ;
        RECT 42.300 65.200 44.200 65.500 ;
        RECT 45.400 65.400 45.800 66.200 ;
        RECT 46.100 65.800 46.600 66.200 ;
        RECT 41.300 64.600 42.100 64.900 ;
        RECT 35.000 61.500 35.400 63.500 ;
        RECT 37.100 61.100 37.500 64.600 ;
        RECT 41.700 61.100 42.100 64.600 ;
        RECT 43.900 63.500 44.200 65.200 ;
        RECT 46.100 64.900 46.400 65.800 ;
        RECT 47.100 65.500 47.400 66.500 ;
        RECT 47.800 65.800 48.200 66.600 ;
        RECT 48.600 66.100 49.000 66.600 ;
        RECT 51.900 66.200 52.300 66.600 ;
        RECT 52.600 66.200 52.900 67.900 ;
        RECT 53.400 66.400 53.800 67.200 ;
        RECT 55.800 66.400 56.200 67.200 ;
        RECT 56.700 66.200 57.000 67.900 ;
        RECT 57.400 66.800 57.800 67.200 ;
        RECT 59.000 66.800 59.400 67.600 ;
        RECT 59.800 67.100 60.200 67.900 ;
        RECT 61.500 67.700 63.300 67.900 ;
        RECT 61.800 67.200 62.200 67.400 ;
        RECT 63.800 67.200 64.100 67.900 ;
        RECT 66.200 67.800 66.600 67.900 ;
        RECT 61.400 67.100 62.200 67.200 ;
        RECT 59.800 66.900 62.200 67.100 ;
        RECT 59.800 66.800 61.800 66.900 ;
        RECT 62.900 66.800 64.200 67.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 57.400 66.600 57.700 66.800 ;
        RECT 57.300 66.200 57.700 66.600 ;
        RECT 50.200 66.100 50.600 66.200 ;
        RECT 48.600 65.800 50.600 66.100 ;
        RECT 47.100 65.200 49.000 65.500 ;
        RECT 51.000 65.400 51.400 66.200 ;
        RECT 52.600 65.800 53.000 66.200 ;
        RECT 54.200 66.100 54.600 66.200 ;
        RECT 53.800 65.800 54.600 66.100 ;
        RECT 55.000 66.100 55.400 66.200 ;
        RECT 55.000 65.800 55.800 66.100 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 52.600 65.700 52.900 65.800 ;
        RECT 51.900 65.400 52.900 65.700 ;
        RECT 53.800 65.600 54.200 65.800 ;
        RECT 55.400 65.600 55.800 65.800 ;
        RECT 56.700 65.700 57.000 65.800 ;
        RECT 56.700 65.400 57.700 65.700 ;
        RECT 58.200 65.400 58.600 66.200 ;
        RECT 46.100 64.600 46.900 64.900 ;
        RECT 43.800 61.500 44.200 63.500 ;
        RECT 46.500 61.100 46.900 64.600 ;
        RECT 48.700 63.500 49.000 65.200 ;
        RECT 51.900 65.100 52.200 65.400 ;
        RECT 57.400 65.100 57.700 65.400 ;
        RECT 48.600 61.500 49.000 63.500 ;
        RECT 51.000 61.400 51.400 65.100 ;
        RECT 51.800 61.700 52.200 65.100 ;
        RECT 52.600 64.800 54.600 65.100 ;
        RECT 52.600 61.400 53.000 64.800 ;
        RECT 51.000 61.100 53.000 61.400 ;
        RECT 54.200 61.100 54.600 64.800 ;
        RECT 55.000 64.800 57.000 65.100 ;
        RECT 55.000 61.100 55.400 64.800 ;
        RECT 56.600 61.400 57.000 64.800 ;
        RECT 57.400 61.700 57.800 65.100 ;
        RECT 58.200 61.400 58.600 65.100 ;
        RECT 56.600 61.100 58.600 61.400 ;
        RECT 59.800 61.100 60.200 66.800 ;
        RECT 62.200 65.800 62.600 66.600 ;
        RECT 60.600 64.400 61.000 65.200 ;
        RECT 62.900 65.100 63.200 66.800 ;
        RECT 65.500 66.600 65.800 66.800 ;
        RECT 65.500 66.200 65.900 66.600 ;
        RECT 66.200 66.200 66.500 67.800 ;
        RECT 67.000 66.400 67.400 67.200 ;
        RECT 68.600 66.800 69.000 67.600 ;
        RECT 63.800 66.100 64.200 66.200 ;
        RECT 64.600 66.100 65.000 66.200 ;
        RECT 63.800 65.800 65.000 66.100 ;
        RECT 64.600 65.400 65.000 65.800 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 67.800 66.100 68.200 66.200 ;
        RECT 69.400 66.100 69.800 67.900 ;
        RECT 72.500 67.700 73.300 68.000 ;
        RECT 72.500 67.500 72.900 67.700 ;
        RECT 72.500 67.200 72.800 67.500 ;
        RECT 75.100 67.400 75.400 68.500 ;
        RECT 77.300 68.200 78.100 69.900 ;
        RECT 77.300 67.900 78.600 68.200 ;
        RECT 79.800 67.900 80.200 69.900 ;
        RECT 80.600 68.000 81.000 69.900 ;
        RECT 82.200 68.000 82.600 69.900 ;
        RECT 84.300 68.200 84.700 69.900 ;
        RECT 80.600 67.900 82.600 68.000 ;
        RECT 83.800 67.900 84.700 68.200 ;
        RECT 85.400 67.900 85.800 69.900 ;
        RECT 87.500 68.400 87.900 69.900 ;
        RECT 87.500 67.900 88.200 68.400 ;
        RECT 90.100 67.900 90.900 69.900 ;
        RECT 93.900 69.100 94.300 69.900 ;
        RECT 93.900 68.800 96.100 69.100 ;
        RECT 93.900 68.200 94.300 68.800 ;
        RECT 93.400 67.900 94.300 68.200 ;
        RECT 95.800 68.200 96.100 68.800 ;
        RECT 71.800 66.800 72.800 67.200 ;
        RECT 73.300 67.100 75.400 67.400 ;
        RECT 77.500 67.800 78.600 67.900 ;
        RECT 73.300 66.900 73.800 67.100 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 67.400 65.800 68.200 66.100 ;
        RECT 68.600 65.800 69.800 66.100 ;
        RECT 66.200 65.700 66.500 65.800 ;
        RECT 65.500 65.400 66.500 65.700 ;
        RECT 67.400 65.600 67.800 65.800 ;
        RECT 63.800 65.100 64.200 65.200 ;
        RECT 65.500 65.100 65.800 65.400 ;
        RECT 68.600 65.200 68.900 65.800 ;
        RECT 62.700 64.800 63.200 65.100 ;
        RECT 63.500 64.800 64.200 65.100 ;
        RECT 62.700 62.200 63.100 64.800 ;
        RECT 63.500 64.200 63.800 64.800 ;
        RECT 63.400 63.800 63.800 64.200 ;
        RECT 62.200 61.800 63.100 62.200 ;
        RECT 62.700 61.100 63.100 61.800 ;
        RECT 64.600 61.400 65.000 65.100 ;
        RECT 65.400 61.700 65.800 65.100 ;
        RECT 66.200 64.800 68.200 65.100 ;
        RECT 68.600 64.800 69.000 65.200 ;
        RECT 66.200 61.400 66.600 64.800 ;
        RECT 64.600 61.100 66.600 61.400 ;
        RECT 67.800 61.100 68.200 64.800 ;
        RECT 69.400 61.100 69.800 65.800 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 70.200 65.200 70.500 65.800 ;
        RECT 71.800 65.400 72.200 66.200 ;
        RECT 70.200 64.400 70.600 65.200 ;
        RECT 72.500 64.900 72.800 66.800 ;
        RECT 73.100 66.500 73.800 66.900 ;
        RECT 73.500 65.500 73.800 66.500 ;
        RECT 74.200 65.800 74.600 66.600 ;
        RECT 75.000 65.800 75.400 66.600 ;
        RECT 76.600 66.400 77.000 67.200 ;
        RECT 77.500 66.200 77.800 67.800 ;
        RECT 79.900 67.200 80.200 67.900 ;
        RECT 80.700 67.700 82.500 67.900 ;
        RECT 81.800 67.200 82.200 67.400 ;
        RECT 78.200 66.800 78.600 67.200 ;
        RECT 79.800 66.800 81.100 67.200 ;
        RECT 81.800 66.900 82.600 67.200 ;
        RECT 78.200 66.600 78.500 66.800 ;
        RECT 78.100 66.200 78.500 66.600 ;
        RECT 80.800 66.200 81.100 66.800 ;
        RECT 82.200 66.800 82.600 66.900 ;
        RECT 83.000 66.800 83.400 67.600 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 75.800 65.800 76.600 66.100 ;
        RECT 77.400 65.800 77.800 66.200 ;
        RECT 76.200 65.600 76.600 65.800 ;
        RECT 77.500 65.700 77.800 65.800 ;
        RECT 73.500 65.200 75.400 65.500 ;
        RECT 77.500 65.400 78.500 65.700 ;
        RECT 79.000 65.400 79.400 66.200 ;
        RECT 80.600 65.800 81.100 66.200 ;
        RECT 81.400 65.800 81.800 66.600 ;
        RECT 82.200 66.100 82.500 66.800 ;
        RECT 83.800 66.100 84.200 67.900 ;
        RECT 85.500 67.800 85.800 67.900 ;
        RECT 85.500 67.600 86.400 67.800 ;
        RECT 85.500 67.500 87.600 67.600 ;
        RECT 86.100 67.300 87.600 67.500 ;
        RECT 87.200 67.200 87.600 67.300 ;
        RECT 85.400 66.400 85.800 67.200 ;
        RECT 86.400 66.900 86.800 67.000 ;
        RECT 86.300 66.600 86.800 66.900 ;
        RECT 86.300 66.200 86.600 66.600 ;
        RECT 82.200 65.800 84.200 66.100 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 72.500 64.600 73.300 64.900 ;
        RECT 72.900 62.200 73.300 64.600 ;
        RECT 75.100 63.500 75.400 65.200 ;
        RECT 78.200 65.100 78.500 65.400 ;
        RECT 79.800 65.100 80.200 65.200 ;
        RECT 80.800 65.100 81.100 65.800 ;
        RECT 72.600 61.800 73.300 62.200 ;
        RECT 72.900 61.100 73.300 61.800 ;
        RECT 75.000 61.500 75.400 63.500 ;
        RECT 75.800 64.800 77.800 65.100 ;
        RECT 75.800 61.100 76.200 64.800 ;
        RECT 77.400 61.400 77.800 64.800 ;
        RECT 78.200 61.700 78.600 65.100 ;
        RECT 79.000 61.400 79.400 65.100 ;
        RECT 79.800 64.800 80.500 65.100 ;
        RECT 80.800 64.800 81.300 65.100 ;
        RECT 80.200 64.200 80.500 64.800 ;
        RECT 80.200 63.800 80.600 64.200 ;
        RECT 77.400 61.100 79.400 61.400 ;
        RECT 80.900 61.100 81.300 64.800 ;
        RECT 83.800 61.100 84.200 65.800 ;
        RECT 87.200 65.500 87.500 67.200 ;
        RECT 87.900 66.200 88.200 67.900 ;
        RECT 89.400 66.400 89.800 67.200 ;
        RECT 90.300 66.200 90.600 67.900 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 92.600 66.800 93.000 67.600 ;
        RECT 91.000 66.600 91.300 66.800 ;
        RECT 90.900 66.200 91.300 66.600 ;
        RECT 87.800 65.800 88.200 66.200 ;
        RECT 88.600 66.100 89.000 66.200 ;
        RECT 88.600 65.800 89.400 66.100 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 86.300 65.200 87.500 65.500 ;
        RECT 84.600 64.400 85.000 65.200 ;
        RECT 86.300 63.100 86.600 65.200 ;
        RECT 87.900 65.100 88.200 65.800 ;
        RECT 89.000 65.600 89.400 65.800 ;
        RECT 90.300 65.700 90.600 65.800 ;
        RECT 90.300 65.400 91.300 65.700 ;
        RECT 91.800 65.400 92.200 66.200 ;
        RECT 91.000 65.100 91.300 65.400 ;
        RECT 86.200 61.100 86.600 63.100 ;
        RECT 87.800 61.100 88.200 65.100 ;
        RECT 88.600 64.800 90.600 65.100 ;
        RECT 88.600 61.100 89.000 64.800 ;
        RECT 90.200 61.400 90.600 64.800 ;
        RECT 91.000 61.700 91.400 65.100 ;
        RECT 91.800 61.400 92.200 65.100 ;
        RECT 90.200 61.100 92.200 61.400 ;
        RECT 93.400 61.100 93.800 67.900 ;
        RECT 95.800 67.800 96.200 68.200 ;
        RECT 96.600 67.700 97.000 69.900 ;
        RECT 98.700 69.200 99.300 69.900 ;
        RECT 98.700 68.900 99.400 69.200 ;
        RECT 101.000 68.900 101.400 69.900 ;
        RECT 103.200 69.200 103.600 69.900 ;
        RECT 103.200 68.900 104.200 69.200 ;
        RECT 99.000 68.500 99.400 68.900 ;
        RECT 101.100 68.600 101.400 68.900 ;
        RECT 101.100 68.300 102.500 68.600 ;
        RECT 102.100 68.200 102.500 68.300 ;
        RECT 103.000 68.200 103.400 68.600 ;
        RECT 103.800 68.500 104.200 68.900 ;
        RECT 98.100 67.700 98.500 67.800 ;
        RECT 96.600 67.400 98.500 67.700 ;
        RECT 96.600 65.700 97.000 67.400 ;
        RECT 100.100 67.100 100.500 67.200 ;
        RECT 103.000 67.100 103.300 68.200 ;
        RECT 105.400 67.500 105.800 69.900 ;
        RECT 106.200 67.800 106.600 68.600 ;
        RECT 104.600 67.100 105.400 67.200 ;
        RECT 99.900 66.800 105.400 67.100 ;
        RECT 99.000 66.400 99.400 66.500 ;
        RECT 97.500 66.100 99.400 66.400 ;
        RECT 97.500 66.000 97.900 66.100 ;
        RECT 98.300 65.700 98.700 65.800 ;
        RECT 96.600 65.400 98.700 65.700 ;
        RECT 94.200 64.400 94.600 65.200 ;
        RECT 96.600 61.100 97.000 65.400 ;
        RECT 99.900 65.200 100.200 66.800 ;
        RECT 103.500 66.700 103.900 66.800 ;
        RECT 104.300 66.200 104.700 66.300 ;
        RECT 100.600 66.100 101.000 66.200 ;
        RECT 102.200 66.100 104.700 66.200 ;
        RECT 100.600 65.900 104.700 66.100 ;
        RECT 100.600 65.800 102.600 65.900 ;
        RECT 103.000 65.500 105.800 65.600 ;
        RECT 102.900 65.400 105.800 65.500 ;
        RECT 99.000 64.900 100.200 65.200 ;
        RECT 100.900 65.300 105.800 65.400 ;
        RECT 100.900 65.100 103.300 65.300 ;
        RECT 99.000 64.400 99.300 64.900 ;
        RECT 98.600 64.000 99.300 64.400 ;
        RECT 100.100 64.500 100.500 64.600 ;
        RECT 100.900 64.500 101.200 65.100 ;
        RECT 100.100 64.200 101.200 64.500 ;
        RECT 101.500 64.500 104.200 64.800 ;
        RECT 101.500 64.400 101.900 64.500 ;
        RECT 103.800 64.400 104.200 64.500 ;
        RECT 100.700 63.700 101.100 63.800 ;
        RECT 102.100 63.700 102.500 63.800 ;
        RECT 99.000 63.100 99.400 63.500 ;
        RECT 100.700 63.400 102.500 63.700 ;
        RECT 101.100 63.100 101.400 63.400 ;
        RECT 103.800 63.100 104.200 63.500 ;
        RECT 98.700 61.100 99.300 63.100 ;
        RECT 101.000 61.100 101.400 63.100 ;
        RECT 103.200 62.800 104.200 63.100 ;
        RECT 103.200 61.100 103.600 62.800 ;
        RECT 105.400 61.100 105.800 65.300 ;
        RECT 107.000 61.100 107.400 69.900 ;
        RECT 109.100 69.200 109.500 69.900 ;
        RECT 111.500 69.200 111.900 69.900 ;
        RECT 109.100 68.800 109.800 69.200 ;
        RECT 111.000 68.800 111.900 69.200 ;
        RECT 109.100 68.200 109.500 68.800 ;
        RECT 111.500 68.200 111.900 68.800 ;
        RECT 108.600 67.900 109.500 68.200 ;
        RECT 111.000 67.900 111.900 68.200 ;
        RECT 112.900 68.200 113.300 69.900 ;
        RECT 116.300 68.200 117.100 69.900 ;
        RECT 112.900 67.900 113.800 68.200 ;
        RECT 107.800 66.800 108.200 67.600 ;
        RECT 108.600 61.100 109.000 67.900 ;
        RECT 109.400 67.100 109.800 67.200 ;
        RECT 110.200 67.100 110.600 67.600 ;
        RECT 109.400 66.800 110.600 67.100 ;
        RECT 109.400 64.400 109.800 65.200 ;
        RECT 111.000 61.100 111.400 67.900 ;
        RECT 112.600 66.100 113.000 66.200 ;
        RECT 113.400 66.100 113.800 67.900 ;
        RECT 115.800 67.900 117.100 68.200 ;
        RECT 115.800 67.800 116.900 67.900 ;
        RECT 114.200 66.800 114.600 67.600 ;
        RECT 115.800 66.800 116.200 67.200 ;
        RECT 115.900 66.600 116.200 66.800 ;
        RECT 115.900 66.200 116.300 66.600 ;
        RECT 116.600 66.200 116.900 67.800 ;
        RECT 119.000 67.700 119.400 69.900 ;
        RECT 121.100 69.200 121.700 69.900 ;
        RECT 121.100 68.900 121.800 69.200 ;
        RECT 123.400 68.900 123.800 69.900 ;
        RECT 125.600 69.200 126.000 69.900 ;
        RECT 125.600 68.900 126.600 69.200 ;
        RECT 121.400 68.500 121.800 68.900 ;
        RECT 123.500 68.600 123.800 68.900 ;
        RECT 123.500 68.300 124.900 68.600 ;
        RECT 124.500 68.200 124.900 68.300 ;
        RECT 125.400 68.200 125.800 68.600 ;
        RECT 126.200 68.500 126.600 68.900 ;
        RECT 120.500 67.700 120.900 67.800 ;
        RECT 119.000 67.400 120.900 67.700 ;
        RECT 117.400 66.400 117.800 67.200 ;
        RECT 112.600 65.800 113.800 66.100 ;
        RECT 111.800 64.400 112.200 65.200 ;
        RECT 112.600 64.400 113.000 65.200 ;
        RECT 113.400 61.100 113.800 65.800 ;
        RECT 115.000 65.400 115.400 66.200 ;
        RECT 116.600 65.800 117.000 66.200 ;
        RECT 118.200 66.100 118.600 66.200 ;
        RECT 117.800 65.800 118.600 66.100 ;
        RECT 116.600 65.700 116.900 65.800 ;
        RECT 115.900 65.400 116.900 65.700 ;
        RECT 117.800 65.600 118.200 65.800 ;
        RECT 119.000 65.700 119.400 67.400 ;
        RECT 122.500 67.100 122.900 67.200 ;
        RECT 125.400 67.100 125.700 68.200 ;
        RECT 127.800 67.500 128.200 69.900 ;
        RECT 129.900 68.200 130.300 69.900 ;
        RECT 129.400 67.900 130.300 68.200 ;
        RECT 131.000 67.900 131.400 69.900 ;
        RECT 131.800 68.000 132.200 69.900 ;
        RECT 133.400 68.000 133.800 69.900 ;
        RECT 131.800 67.900 133.800 68.000 ;
        RECT 135.800 67.900 136.200 69.900 ;
        RECT 138.200 68.900 138.600 69.900 ;
        RECT 136.500 68.200 136.900 68.600 ;
        RECT 136.600 68.100 137.000 68.200 ;
        RECT 138.200 68.100 138.500 68.900 ;
        RECT 127.000 67.100 127.800 67.200 ;
        RECT 122.300 66.800 127.800 67.100 ;
        RECT 128.600 66.800 129.000 67.600 ;
        RECT 121.400 66.400 121.800 66.500 ;
        RECT 119.900 66.100 121.800 66.400 ;
        RECT 122.300 66.200 122.600 66.800 ;
        RECT 125.900 66.700 126.300 66.800 ;
        RECT 125.400 66.200 125.800 66.300 ;
        RECT 126.700 66.200 127.100 66.300 ;
        RECT 119.900 66.000 120.300 66.100 ;
        RECT 122.200 65.800 122.600 66.200 ;
        RECT 124.600 65.900 127.100 66.200 ;
        RECT 129.400 66.100 129.800 67.900 ;
        RECT 131.100 67.200 131.400 67.900 ;
        RECT 131.900 67.700 133.700 67.900 ;
        RECT 133.000 67.200 133.400 67.400 ;
        RECT 131.000 66.800 132.300 67.200 ;
        RECT 133.000 66.900 133.800 67.200 ;
        RECT 124.600 65.800 125.000 65.900 ;
        RECT 129.400 65.800 131.300 66.100 ;
        RECT 120.700 65.700 121.100 65.800 ;
        RECT 119.000 65.400 121.100 65.700 ;
        RECT 115.900 65.100 116.200 65.400 ;
        RECT 115.000 61.400 115.400 65.100 ;
        RECT 115.800 61.700 116.200 65.100 ;
        RECT 116.600 64.800 118.600 65.100 ;
        RECT 116.600 61.400 117.000 64.800 ;
        RECT 115.000 61.100 117.000 61.400 ;
        RECT 118.200 61.100 118.600 64.800 ;
        RECT 119.000 61.100 119.400 65.400 ;
        RECT 122.300 65.200 122.600 65.800 ;
        RECT 125.400 65.500 128.200 65.600 ;
        RECT 125.300 65.400 128.200 65.500 ;
        RECT 121.400 64.900 122.600 65.200 ;
        RECT 123.300 65.300 128.200 65.400 ;
        RECT 123.300 65.100 125.700 65.300 ;
        RECT 121.400 64.400 121.700 64.900 ;
        RECT 121.000 64.000 121.700 64.400 ;
        RECT 122.500 64.500 122.900 64.600 ;
        RECT 123.300 64.500 123.600 65.100 ;
        RECT 122.500 64.200 123.600 64.500 ;
        RECT 123.900 64.500 126.600 64.800 ;
        RECT 123.900 64.400 124.300 64.500 ;
        RECT 126.200 64.400 126.600 64.500 ;
        RECT 123.100 63.700 123.500 63.800 ;
        RECT 124.500 63.700 124.900 63.800 ;
        RECT 121.400 63.100 121.800 63.500 ;
        RECT 123.100 63.400 124.900 63.700 ;
        RECT 123.500 63.100 123.800 63.400 ;
        RECT 126.200 63.100 126.600 63.500 ;
        RECT 121.100 61.100 121.700 63.100 ;
        RECT 123.400 61.100 123.800 63.100 ;
        RECT 125.600 62.800 126.600 63.100 ;
        RECT 125.600 61.100 126.000 62.800 ;
        RECT 127.800 61.100 128.200 65.300 ;
        RECT 129.400 61.100 129.800 65.800 ;
        RECT 131.000 65.200 131.300 65.800 ;
        RECT 130.200 64.400 130.600 65.200 ;
        RECT 131.000 65.100 131.400 65.200 ;
        RECT 132.000 65.100 132.300 66.800 ;
        RECT 133.400 66.800 133.800 66.900 ;
        RECT 132.600 65.800 133.000 66.600 ;
        RECT 133.400 66.100 133.700 66.800 ;
        RECT 135.000 66.400 135.400 67.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 135.800 66.100 136.100 67.900 ;
        RECT 136.600 67.800 138.500 68.100 ;
        RECT 139.000 67.800 139.400 68.600 ;
        RECT 138.200 67.200 138.500 67.800 ;
        RECT 139.800 67.500 140.200 69.900 ;
        RECT 142.000 69.200 142.400 69.900 ;
        RECT 141.400 68.900 142.400 69.200 ;
        RECT 144.200 68.900 144.600 69.900 ;
        RECT 146.300 69.200 146.900 69.900 ;
        RECT 146.200 68.900 146.900 69.200 ;
        RECT 141.400 68.500 141.800 68.900 ;
        RECT 144.200 68.600 144.500 68.900 ;
        RECT 142.200 68.200 142.600 68.600 ;
        RECT 143.100 68.300 144.500 68.600 ;
        RECT 146.200 68.500 146.600 68.900 ;
        RECT 143.100 68.200 143.500 68.300 ;
        RECT 138.200 66.800 138.600 67.200 ;
        RECT 140.200 67.100 141.000 67.200 ;
        RECT 142.300 67.100 142.600 68.200 ;
        RECT 147.100 67.700 147.500 67.800 ;
        RECT 148.600 67.700 149.000 69.900 ;
        RECT 147.100 67.400 149.000 67.700 ;
        RECT 151.000 67.500 151.400 69.900 ;
        RECT 153.200 69.200 153.600 69.900 ;
        RECT 152.600 68.900 153.600 69.200 ;
        RECT 155.400 68.900 155.800 69.900 ;
        RECT 157.500 69.200 158.100 69.900 ;
        RECT 157.400 68.900 158.100 69.200 ;
        RECT 152.600 68.500 153.000 68.900 ;
        RECT 155.400 68.600 155.700 68.900 ;
        RECT 153.400 68.200 153.800 68.600 ;
        RECT 154.300 68.300 155.700 68.600 ;
        RECT 157.400 68.500 157.800 68.900 ;
        RECT 154.300 68.200 154.700 68.300 ;
        RECT 145.100 67.100 145.500 67.200 ;
        RECT 140.200 66.800 145.700 67.100 ;
        RECT 136.600 66.100 137.000 66.200 ;
        RECT 133.400 65.800 135.000 66.100 ;
        RECT 135.800 65.800 137.000 66.100 ;
        RECT 134.600 65.600 135.000 65.800 ;
        RECT 136.600 65.100 136.900 65.800 ;
        RECT 137.400 65.400 137.800 66.200 ;
        RECT 138.200 65.100 138.500 66.800 ;
        RECT 141.700 66.700 142.100 66.800 ;
        RECT 140.900 66.200 141.300 66.300 ;
        RECT 142.200 66.200 142.600 66.300 ;
        RECT 140.900 65.900 143.400 66.200 ;
        RECT 143.000 65.800 143.400 65.900 ;
        RECT 144.600 66.100 145.000 66.200 ;
        RECT 145.400 66.100 145.700 66.800 ;
        RECT 146.200 66.400 146.600 66.500 ;
        RECT 146.200 66.100 148.100 66.400 ;
        RECT 144.600 65.800 145.700 66.100 ;
        RECT 147.700 66.000 148.100 66.100 ;
        RECT 139.800 65.500 142.600 65.600 ;
        RECT 139.800 65.400 142.700 65.500 ;
        RECT 139.800 65.300 144.700 65.400 ;
        RECT 131.000 64.800 131.700 65.100 ;
        RECT 132.000 64.800 132.500 65.100 ;
        RECT 131.400 64.200 131.700 64.800 ;
        RECT 131.400 63.800 131.800 64.200 ;
        RECT 132.100 61.100 132.500 64.800 ;
        RECT 134.200 64.800 136.200 65.100 ;
        RECT 134.200 61.100 134.600 64.800 ;
        RECT 135.800 61.100 136.200 64.800 ;
        RECT 136.600 61.100 137.000 65.100 ;
        RECT 137.700 64.700 138.600 65.100 ;
        RECT 137.700 61.100 138.100 64.700 ;
        RECT 139.800 61.100 140.200 65.300 ;
        RECT 142.300 65.100 144.700 65.300 ;
        RECT 141.400 64.500 144.100 64.800 ;
        RECT 141.400 64.400 141.800 64.500 ;
        RECT 143.700 64.400 144.100 64.500 ;
        RECT 144.400 64.500 144.700 65.100 ;
        RECT 145.400 65.200 145.700 65.800 ;
        RECT 146.900 65.700 147.300 65.800 ;
        RECT 148.600 65.700 149.000 67.400 ;
        RECT 151.400 67.100 152.200 67.200 ;
        RECT 153.500 67.100 153.800 68.200 ;
        RECT 158.300 67.700 158.700 67.800 ;
        RECT 159.800 67.700 160.200 69.900 ;
        RECT 161.900 68.200 162.300 69.900 ;
        RECT 158.300 67.400 160.200 67.700 ;
        RECT 161.400 67.900 162.300 68.200 ;
        RECT 163.000 67.900 163.400 69.900 ;
        RECT 163.800 68.000 164.200 69.900 ;
        RECT 165.400 68.000 165.800 69.900 ;
        RECT 163.800 67.900 165.800 68.000 ;
        RECT 167.500 67.900 168.300 69.900 ;
        RECT 170.200 68.500 170.600 69.500 ;
        RECT 156.300 67.100 156.700 67.200 ;
        RECT 159.800 67.100 160.200 67.400 ;
        RECT 160.600 67.100 161.000 67.600 ;
        RECT 151.400 66.800 156.900 67.100 ;
        RECT 152.900 66.700 153.300 66.800 ;
        RECT 152.100 66.200 152.500 66.300 ;
        RECT 152.100 66.100 154.600 66.200 ;
        RECT 155.800 66.100 156.200 66.200 ;
        RECT 152.100 65.900 156.200 66.100 ;
        RECT 154.200 65.800 156.200 65.900 ;
        RECT 146.900 65.400 149.000 65.700 ;
        RECT 145.400 64.900 146.600 65.200 ;
        RECT 145.100 64.500 145.500 64.600 ;
        RECT 144.400 64.200 145.500 64.500 ;
        RECT 146.300 64.400 146.600 64.900 ;
        RECT 146.300 64.000 147.000 64.400 ;
        RECT 143.100 63.700 143.500 63.800 ;
        RECT 144.500 63.700 144.900 63.800 ;
        RECT 141.400 63.100 141.800 63.500 ;
        RECT 143.100 63.400 144.900 63.700 ;
        RECT 144.200 63.100 144.500 63.400 ;
        RECT 146.200 63.100 146.600 63.500 ;
        RECT 141.400 62.800 142.400 63.100 ;
        RECT 142.000 61.100 142.400 62.800 ;
        RECT 144.200 61.100 144.600 63.100 ;
        RECT 146.300 61.100 146.900 63.100 ;
        RECT 148.600 61.100 149.000 65.400 ;
        RECT 151.000 65.500 153.800 65.600 ;
        RECT 151.000 65.400 153.900 65.500 ;
        RECT 151.000 65.300 155.900 65.400 ;
        RECT 151.000 61.100 151.400 65.300 ;
        RECT 153.500 65.100 155.900 65.300 ;
        RECT 152.600 64.500 155.300 64.800 ;
        RECT 152.600 64.400 153.000 64.500 ;
        RECT 154.900 64.400 155.300 64.500 ;
        RECT 155.600 64.500 155.900 65.100 ;
        RECT 156.600 65.200 156.900 66.800 ;
        RECT 159.800 66.800 161.000 67.100 ;
        RECT 157.400 66.400 157.800 66.500 ;
        RECT 157.400 66.100 159.300 66.400 ;
        RECT 158.900 66.000 159.300 66.100 ;
        RECT 158.100 65.700 158.500 65.800 ;
        RECT 159.800 65.700 160.200 66.800 ;
        RECT 158.100 65.400 160.200 65.700 ;
        RECT 156.600 64.900 157.800 65.200 ;
        RECT 156.300 64.500 156.700 64.600 ;
        RECT 155.600 64.200 156.700 64.500 ;
        RECT 157.500 64.400 157.800 64.900 ;
        RECT 157.500 64.000 158.200 64.400 ;
        RECT 154.300 63.700 154.700 63.800 ;
        RECT 155.700 63.700 156.100 63.800 ;
        RECT 152.600 63.100 153.000 63.500 ;
        RECT 154.300 63.400 156.100 63.700 ;
        RECT 155.400 63.100 155.700 63.400 ;
        RECT 157.400 63.100 157.800 63.500 ;
        RECT 152.600 62.800 153.600 63.100 ;
        RECT 153.200 61.100 153.600 62.800 ;
        RECT 155.400 61.100 155.800 63.100 ;
        RECT 157.500 61.100 158.100 63.100 ;
        RECT 159.800 61.100 160.200 65.400 ;
        RECT 161.400 66.100 161.800 67.900 ;
        RECT 163.100 67.200 163.400 67.900 ;
        RECT 163.900 67.700 165.700 67.900 ;
        RECT 165.000 67.200 165.400 67.400 ;
        RECT 163.000 66.800 164.300 67.200 ;
        RECT 165.000 67.100 165.800 67.200 ;
        RECT 166.200 67.100 166.600 67.200 ;
        RECT 165.000 66.900 166.600 67.100 ;
        RECT 165.400 66.800 166.600 66.900 ;
        RECT 167.000 66.800 167.400 67.200 ;
        RECT 161.400 65.800 163.300 66.100 ;
        RECT 161.400 61.100 161.800 65.800 ;
        RECT 163.000 65.200 163.300 65.800 ;
        RECT 162.200 64.400 162.600 65.200 ;
        RECT 163.000 65.100 163.400 65.200 ;
        RECT 164.000 65.100 164.300 66.800 ;
        RECT 167.100 66.600 167.400 66.800 ;
        RECT 164.600 65.800 165.000 66.600 ;
        RECT 167.100 66.200 167.500 66.600 ;
        RECT 167.800 66.200 168.100 67.900 ;
        RECT 170.200 67.400 170.500 68.500 ;
        RECT 172.300 68.200 172.700 69.500 ;
        RECT 171.800 68.000 172.700 68.200 ;
        RECT 171.800 67.800 173.100 68.000 ;
        RECT 172.300 67.700 173.100 67.800 ;
        RECT 172.700 67.500 173.100 67.700 ;
        RECT 175.000 67.500 175.400 69.900 ;
        RECT 177.200 69.200 177.600 69.900 ;
        RECT 176.600 68.900 177.600 69.200 ;
        RECT 179.400 68.900 179.800 69.900 ;
        RECT 181.500 69.200 182.100 69.900 ;
        RECT 181.400 68.900 182.100 69.200 ;
        RECT 176.600 68.500 177.000 68.900 ;
        RECT 179.400 68.600 179.700 68.900 ;
        RECT 177.400 67.800 177.800 68.600 ;
        RECT 178.300 68.300 179.700 68.600 ;
        RECT 181.400 68.500 181.800 68.900 ;
        RECT 178.300 68.200 178.700 68.300 ;
        RECT 168.600 66.400 169.000 67.200 ;
        RECT 170.200 67.100 172.300 67.400 ;
        RECT 171.800 66.900 172.300 67.100 ;
        RECT 172.800 67.200 173.100 67.500 ;
        RECT 165.400 66.100 165.800 66.200 ;
        RECT 166.200 66.100 166.600 66.200 ;
        RECT 165.400 65.800 166.600 66.100 ;
        RECT 166.200 65.400 166.600 65.800 ;
        RECT 167.800 65.800 168.200 66.200 ;
        RECT 169.400 66.100 169.800 66.200 ;
        RECT 169.000 65.800 169.800 66.100 ;
        RECT 170.200 65.800 170.600 66.600 ;
        RECT 171.000 65.800 171.400 66.600 ;
        RECT 171.800 66.500 172.500 66.900 ;
        RECT 172.800 66.800 173.800 67.200 ;
        RECT 175.400 67.100 176.200 67.200 ;
        RECT 177.500 67.100 177.800 67.800 ;
        RECT 182.300 67.700 182.700 67.800 ;
        RECT 183.800 67.700 184.200 69.900 ;
        RECT 184.900 69.200 185.300 69.900 ;
        RECT 184.600 68.800 185.300 69.200 ;
        RECT 184.900 68.200 185.300 68.800 ;
        RECT 188.900 68.200 189.300 69.500 ;
        RECT 191.000 68.500 191.400 69.500 ;
        RECT 184.900 67.900 185.800 68.200 ;
        RECT 188.900 68.000 189.800 68.200 ;
        RECT 182.300 67.400 184.200 67.700 ;
        RECT 180.300 67.100 180.700 67.200 ;
        RECT 175.400 66.800 180.900 67.100 ;
        RECT 167.800 65.700 168.100 65.800 ;
        RECT 167.100 65.400 168.100 65.700 ;
        RECT 169.000 65.600 169.400 65.800 ;
        RECT 171.800 65.500 172.100 66.500 ;
        RECT 167.100 65.100 167.400 65.400 ;
        RECT 170.200 65.200 172.100 65.500 ;
        RECT 163.000 64.800 163.700 65.100 ;
        RECT 164.000 64.800 164.500 65.100 ;
        RECT 163.400 64.200 163.700 64.800 ;
        RECT 163.400 63.800 163.800 64.200 ;
        RECT 164.100 61.100 164.500 64.800 ;
        RECT 166.200 61.400 166.600 65.100 ;
        RECT 167.000 61.700 167.400 65.100 ;
        RECT 167.800 64.800 169.800 65.100 ;
        RECT 167.800 61.400 168.200 64.800 ;
        RECT 166.200 61.100 168.200 61.400 ;
        RECT 169.400 61.100 169.800 64.800 ;
        RECT 170.200 63.500 170.500 65.200 ;
        RECT 172.800 64.900 173.100 66.800 ;
        RECT 176.900 66.700 177.300 66.800 ;
        RECT 176.100 66.200 176.500 66.300 ;
        RECT 173.400 65.400 173.800 66.200 ;
        RECT 176.100 66.100 178.600 66.200 ;
        RECT 179.000 66.100 179.400 66.200 ;
        RECT 176.100 65.900 179.400 66.100 ;
        RECT 178.200 65.800 179.400 65.900 ;
        RECT 175.000 65.500 177.800 65.600 ;
        RECT 175.000 65.400 177.900 65.500 ;
        RECT 172.300 64.600 173.100 64.900 ;
        RECT 175.000 65.300 179.900 65.400 ;
        RECT 170.200 61.500 170.600 63.500 ;
        RECT 172.300 61.100 172.700 64.600 ;
        RECT 175.000 61.100 175.400 65.300 ;
        RECT 177.500 65.100 179.900 65.300 ;
        RECT 176.600 64.500 179.300 64.800 ;
        RECT 176.600 64.400 177.000 64.500 ;
        RECT 178.900 64.400 179.300 64.500 ;
        RECT 179.600 64.500 179.900 65.100 ;
        RECT 180.600 65.200 180.900 66.800 ;
        RECT 181.400 66.400 181.800 66.500 ;
        RECT 181.400 66.100 183.300 66.400 ;
        RECT 182.900 66.000 183.300 66.100 ;
        RECT 182.100 65.700 182.500 65.800 ;
        RECT 183.800 65.700 184.200 67.400 ;
        RECT 182.100 65.400 184.200 65.700 ;
        RECT 180.600 64.900 181.800 65.200 ;
        RECT 180.300 64.500 180.700 64.600 ;
        RECT 179.600 64.200 180.700 64.500 ;
        RECT 181.500 64.400 181.800 64.900 ;
        RECT 181.500 64.000 182.200 64.400 ;
        RECT 178.300 63.700 178.700 63.800 ;
        RECT 179.700 63.700 180.100 63.800 ;
        RECT 176.600 63.100 177.000 63.500 ;
        RECT 178.300 63.400 180.100 63.700 ;
        RECT 179.400 63.100 179.700 63.400 ;
        RECT 181.400 63.100 181.800 63.500 ;
        RECT 176.600 62.800 177.600 63.100 ;
        RECT 177.200 61.100 177.600 62.800 ;
        RECT 179.400 61.100 179.800 63.100 ;
        RECT 181.500 61.100 182.100 63.100 ;
        RECT 183.800 61.100 184.200 65.400 ;
        RECT 184.600 64.400 185.000 65.200 ;
        RECT 185.400 61.100 185.800 67.900 ;
        RECT 188.500 67.800 189.800 68.000 ;
        RECT 188.500 67.700 189.300 67.800 ;
        RECT 186.200 66.800 186.600 67.600 ;
        RECT 188.500 67.500 188.900 67.700 ;
        RECT 188.500 67.200 188.800 67.500 ;
        RECT 191.100 67.400 191.400 68.500 ;
        RECT 193.100 67.900 193.900 69.900 ;
        RECT 197.700 69.200 198.100 69.500 ;
        RECT 197.400 68.800 198.100 69.200 ;
        RECT 197.700 68.000 198.100 68.800 ;
        RECT 199.800 68.500 200.200 69.500 ;
        RECT 187.800 66.800 188.800 67.200 ;
        RECT 189.300 67.100 191.400 67.400 ;
        RECT 189.300 66.900 189.800 67.100 ;
        RECT 187.800 65.400 188.200 66.200 ;
        RECT 188.500 64.900 188.800 66.800 ;
        RECT 189.100 66.500 189.800 66.900 ;
        RECT 192.600 66.800 193.000 67.200 ;
        RECT 192.700 66.600 193.000 66.800 ;
        RECT 189.500 65.500 189.800 66.500 ;
        RECT 190.200 65.800 190.600 66.600 ;
        RECT 191.000 65.800 191.400 66.600 ;
        RECT 192.700 66.200 193.100 66.600 ;
        RECT 193.400 66.200 193.700 67.900 ;
        RECT 197.300 67.700 198.100 68.000 ;
        RECT 197.300 67.500 197.700 67.700 ;
        RECT 197.300 67.200 197.600 67.500 ;
        RECT 199.900 67.400 200.200 68.500 ;
        RECT 203.500 68.200 204.300 69.900 ;
        RECT 207.000 68.200 207.400 69.900 ;
        RECT 203.000 67.900 204.300 68.200 ;
        RECT 206.900 67.900 207.400 68.200 ;
        RECT 203.000 67.800 204.100 67.900 ;
        RECT 194.200 66.400 194.600 67.200 ;
        RECT 196.600 66.800 197.600 67.200 ;
        RECT 198.100 67.100 200.200 67.400 ;
        RECT 202.200 67.100 202.600 67.200 ;
        RECT 203.000 67.100 203.400 67.200 ;
        RECT 198.100 66.900 198.600 67.100 ;
        RECT 189.500 65.200 191.400 65.500 ;
        RECT 191.800 65.400 192.200 66.200 ;
        RECT 193.400 65.800 193.800 66.200 ;
        RECT 195.000 66.100 195.400 66.200 ;
        RECT 194.600 65.800 195.400 66.100 ;
        RECT 195.800 66.100 196.200 66.200 ;
        RECT 196.600 66.100 197.000 66.200 ;
        RECT 195.800 65.800 197.000 66.100 ;
        RECT 193.400 65.700 193.700 65.800 ;
        RECT 192.700 65.400 193.700 65.700 ;
        RECT 194.600 65.600 195.000 65.800 ;
        RECT 196.600 65.400 197.000 65.800 ;
        RECT 188.500 64.600 189.300 64.900 ;
        RECT 188.900 61.100 189.300 64.600 ;
        RECT 191.100 63.500 191.400 65.200 ;
        RECT 192.700 65.100 193.000 65.400 ;
        RECT 191.000 61.500 191.400 63.500 ;
        RECT 191.800 61.400 192.200 65.100 ;
        RECT 192.600 61.700 193.000 65.100 ;
        RECT 193.400 64.800 195.400 65.100 ;
        RECT 193.400 61.400 193.800 64.800 ;
        RECT 191.800 61.100 193.800 61.400 ;
        RECT 195.000 61.100 195.400 64.800 ;
        RECT 197.300 64.900 197.600 66.800 ;
        RECT 197.900 66.500 198.600 66.900 ;
        RECT 202.200 66.800 203.400 67.100 ;
        RECT 203.100 66.600 203.400 66.800 ;
        RECT 198.300 65.500 198.600 66.500 ;
        RECT 199.000 65.800 199.400 66.600 ;
        RECT 199.800 65.800 200.200 66.600 ;
        RECT 203.100 66.200 203.500 66.600 ;
        RECT 203.800 66.200 204.100 67.800 ;
        RECT 206.900 67.200 207.200 67.900 ;
        RECT 208.600 67.600 209.000 69.900 ;
        RECT 207.700 67.300 209.000 67.600 ;
        RECT 209.400 67.600 209.800 69.900 ;
        RECT 211.000 68.200 211.400 69.900 ;
        RECT 211.000 67.900 211.500 68.200 ;
        RECT 212.600 68.000 213.000 69.900 ;
        RECT 214.200 68.000 214.600 69.900 ;
        RECT 212.600 67.900 214.600 68.000 ;
        RECT 215.000 67.900 215.400 69.900 ;
        RECT 209.400 67.300 210.700 67.600 ;
        RECT 204.600 66.400 205.000 67.200 ;
        RECT 205.400 67.100 205.800 67.200 ;
        RECT 206.900 67.100 207.400 67.200 ;
        RECT 205.400 66.800 207.400 67.100 ;
        RECT 200.600 66.100 201.000 66.200 ;
        RECT 202.200 66.100 202.600 66.200 ;
        RECT 200.600 65.800 202.600 66.100 ;
        RECT 198.300 65.200 200.200 65.500 ;
        RECT 202.200 65.400 202.600 65.800 ;
        RECT 203.800 65.800 204.200 66.200 ;
        RECT 205.400 66.100 205.800 66.200 ;
        RECT 205.000 65.800 205.800 66.100 ;
        RECT 203.800 65.700 204.100 65.800 ;
        RECT 203.100 65.400 204.100 65.700 ;
        RECT 205.000 65.600 205.400 65.800 ;
        RECT 197.300 64.600 198.100 64.900 ;
        RECT 197.700 61.100 198.100 64.600 ;
        RECT 199.900 63.500 200.200 65.200 ;
        RECT 203.100 65.100 203.400 65.400 ;
        RECT 206.900 65.100 207.200 66.800 ;
        RECT 207.700 66.500 208.000 67.300 ;
        RECT 207.500 66.100 208.000 66.500 ;
        RECT 207.700 65.100 208.000 66.100 ;
        RECT 208.500 66.200 208.900 66.600 ;
        RECT 209.500 66.200 209.900 66.600 ;
        RECT 208.500 66.100 209.000 66.200 ;
        RECT 209.400 66.100 209.900 66.200 ;
        RECT 208.500 65.800 209.900 66.100 ;
        RECT 210.400 66.500 210.700 67.300 ;
        RECT 211.200 67.200 211.500 67.900 ;
        RECT 212.700 67.700 214.500 67.900 ;
        RECT 213.000 67.200 213.400 67.400 ;
        RECT 215.000 67.200 215.300 67.900 ;
        RECT 215.800 67.700 216.200 69.900 ;
        RECT 217.900 69.200 218.500 69.900 ;
        RECT 217.900 68.900 218.600 69.200 ;
        RECT 220.200 68.900 220.600 69.900 ;
        RECT 222.400 69.200 222.800 69.900 ;
        RECT 222.400 68.900 223.400 69.200 ;
        RECT 218.200 68.500 218.600 68.900 ;
        RECT 220.300 68.600 220.600 68.900 ;
        RECT 220.300 68.300 221.700 68.600 ;
        RECT 221.300 68.200 221.700 68.300 ;
        RECT 222.200 68.200 222.600 68.600 ;
        RECT 223.000 68.500 223.400 68.900 ;
        RECT 217.300 67.700 217.700 67.800 ;
        RECT 215.800 67.400 217.700 67.700 ;
        RECT 211.000 66.800 211.500 67.200 ;
        RECT 212.600 66.900 213.400 67.200 ;
        RECT 212.600 66.800 213.000 66.900 ;
        RECT 214.100 66.800 215.400 67.200 ;
        RECT 210.400 66.100 210.900 66.500 ;
        RECT 210.400 65.100 210.700 66.100 ;
        RECT 211.200 65.100 211.500 66.800 ;
        RECT 213.400 65.800 213.800 66.600 ;
        RECT 214.100 65.100 214.400 66.800 ;
        RECT 215.000 66.200 215.300 66.800 ;
        RECT 215.000 65.800 215.400 66.200 ;
        RECT 215.800 65.700 216.200 67.400 ;
        RECT 219.300 67.100 219.700 67.200 ;
        RECT 222.200 67.100 222.500 68.200 ;
        RECT 224.600 67.500 225.000 69.900 ;
        RECT 227.300 68.000 227.700 69.500 ;
        RECT 229.400 68.500 229.800 69.500 ;
        RECT 226.900 67.700 227.700 68.000 ;
        RECT 226.900 67.500 227.300 67.700 ;
        RECT 226.900 67.200 227.200 67.500 ;
        RECT 229.500 67.400 229.800 68.500 ;
        RECT 231.500 68.200 231.900 69.900 ;
        RECT 231.000 67.900 231.900 68.200 ;
        RECT 223.800 67.100 224.600 67.200 ;
        RECT 219.100 66.800 224.600 67.100 ;
        RECT 225.400 67.100 225.800 67.200 ;
        RECT 226.200 67.100 227.200 67.200 ;
        RECT 225.400 66.800 227.200 67.100 ;
        RECT 227.700 67.100 229.800 67.400 ;
        RECT 227.700 66.900 228.200 67.100 ;
        RECT 218.200 66.400 218.600 66.500 ;
        RECT 216.700 66.100 218.600 66.400 ;
        RECT 216.700 66.000 217.100 66.100 ;
        RECT 217.500 65.700 217.900 65.800 ;
        RECT 215.800 65.400 217.900 65.700 ;
        RECT 215.000 65.100 215.400 65.200 ;
        RECT 199.800 61.500 200.200 63.500 ;
        RECT 202.200 61.400 202.600 65.100 ;
        RECT 203.000 61.700 203.400 65.100 ;
        RECT 203.800 64.800 205.800 65.100 ;
        RECT 203.800 61.400 204.200 64.800 ;
        RECT 202.200 61.100 204.200 61.400 ;
        RECT 205.400 61.100 205.800 64.800 ;
        RECT 206.900 64.600 207.400 65.100 ;
        RECT 207.700 64.800 209.000 65.100 ;
        RECT 207.000 61.100 207.400 64.600 ;
        RECT 208.600 61.100 209.000 64.800 ;
        RECT 209.400 64.800 210.700 65.100 ;
        RECT 209.400 61.100 209.800 64.800 ;
        RECT 211.000 64.600 211.500 65.100 ;
        RECT 213.900 64.800 214.400 65.100 ;
        RECT 214.700 64.800 215.400 65.100 ;
        RECT 211.000 61.100 211.400 64.600 ;
        RECT 213.900 61.100 214.300 64.800 ;
        RECT 214.700 64.200 215.000 64.800 ;
        RECT 214.600 63.800 215.000 64.200 ;
        RECT 215.800 61.100 216.200 65.400 ;
        RECT 219.100 65.200 219.400 66.800 ;
        RECT 222.700 66.700 223.100 66.800 ;
        RECT 223.500 66.200 223.900 66.300 ;
        RECT 220.600 66.100 221.000 66.200 ;
        RECT 221.400 66.100 223.900 66.200 ;
        RECT 220.600 65.900 223.900 66.100 ;
        RECT 220.600 65.800 221.800 65.900 ;
        RECT 222.200 65.500 225.000 65.600 ;
        RECT 222.100 65.400 225.000 65.500 ;
        RECT 226.200 65.400 226.600 66.200 ;
        RECT 218.200 64.900 219.400 65.200 ;
        RECT 220.100 65.300 225.000 65.400 ;
        RECT 220.100 65.100 222.500 65.300 ;
        RECT 218.200 64.400 218.500 64.900 ;
        RECT 217.800 64.000 218.500 64.400 ;
        RECT 219.300 64.500 219.700 64.600 ;
        RECT 220.100 64.500 220.400 65.100 ;
        RECT 219.300 64.200 220.400 64.500 ;
        RECT 220.700 64.500 223.400 64.800 ;
        RECT 220.700 64.400 221.100 64.500 ;
        RECT 223.000 64.400 223.400 64.500 ;
        RECT 219.900 63.700 220.300 63.800 ;
        RECT 221.300 63.700 221.700 63.800 ;
        RECT 218.200 63.100 218.600 63.500 ;
        RECT 219.900 63.400 221.700 63.700 ;
        RECT 220.300 63.100 220.600 63.400 ;
        RECT 223.000 63.100 223.400 63.500 ;
        RECT 217.900 61.100 218.500 63.100 ;
        RECT 220.200 61.100 220.600 63.100 ;
        RECT 222.400 62.800 223.400 63.100 ;
        RECT 222.400 61.100 222.800 62.800 ;
        RECT 224.600 61.100 225.000 65.300 ;
        RECT 226.900 64.900 227.200 66.800 ;
        RECT 227.500 66.500 228.200 66.900 ;
        RECT 230.200 66.800 230.600 67.600 ;
        RECT 227.900 65.500 228.200 66.500 ;
        RECT 228.600 65.800 229.000 66.600 ;
        RECT 229.400 65.800 229.800 66.600 ;
        RECT 227.900 65.200 229.800 65.500 ;
        RECT 226.900 64.600 227.700 64.900 ;
        RECT 227.300 61.100 227.700 64.600 ;
        RECT 229.500 63.500 229.800 65.200 ;
        RECT 229.400 61.500 229.800 63.500 ;
        RECT 231.000 61.100 231.400 67.900 ;
        RECT 232.600 67.700 233.000 69.900 ;
        RECT 234.700 69.200 235.300 69.900 ;
        RECT 234.700 68.900 235.400 69.200 ;
        RECT 237.000 68.900 237.400 69.900 ;
        RECT 239.200 69.200 239.600 69.900 ;
        RECT 239.200 68.900 240.200 69.200 ;
        RECT 235.000 68.500 235.400 68.900 ;
        RECT 237.100 68.600 237.400 68.900 ;
        RECT 237.100 68.300 238.500 68.600 ;
        RECT 238.100 68.200 238.500 68.300 ;
        RECT 239.000 68.200 239.400 68.600 ;
        RECT 239.800 68.500 240.200 68.900 ;
        RECT 235.800 67.800 236.200 68.200 ;
        RECT 234.100 67.700 234.500 67.800 ;
        RECT 232.600 67.400 234.500 67.700 ;
        RECT 232.600 65.700 233.000 67.400 ;
        RECT 235.800 67.200 236.100 67.800 ;
        RECT 235.800 67.100 236.500 67.200 ;
        RECT 239.000 67.100 239.300 68.200 ;
        RECT 241.400 67.500 241.800 69.900 ;
        RECT 242.200 67.500 242.600 69.900 ;
        RECT 244.400 69.200 244.800 69.900 ;
        RECT 243.800 68.900 244.800 69.200 ;
        RECT 246.600 68.900 247.000 69.900 ;
        RECT 248.700 69.200 249.300 69.900 ;
        RECT 248.600 68.900 249.300 69.200 ;
        RECT 243.800 68.500 244.200 68.900 ;
        RECT 246.600 68.600 246.900 68.900 ;
        RECT 244.600 68.200 245.000 68.600 ;
        RECT 245.500 68.300 246.900 68.600 ;
        RECT 248.600 68.500 249.000 68.900 ;
        RECT 245.500 68.200 245.900 68.300 ;
        RECT 240.600 67.100 241.400 67.200 ;
        RECT 242.600 67.100 243.400 67.200 ;
        RECT 244.700 67.100 245.000 68.200 ;
        RECT 249.500 67.700 249.900 67.800 ;
        RECT 251.000 67.700 251.400 69.900 ;
        RECT 249.500 67.400 251.400 67.700 ;
        RECT 247.500 67.100 247.900 67.200 ;
        RECT 235.800 66.800 248.100 67.100 ;
        RECT 235.000 66.400 235.400 66.500 ;
        RECT 233.500 66.100 235.400 66.400 ;
        RECT 233.500 66.000 233.900 66.100 ;
        RECT 234.300 65.700 234.700 65.800 ;
        RECT 232.600 65.400 234.700 65.700 ;
        RECT 231.800 64.400 232.200 65.200 ;
        RECT 232.600 61.100 233.000 65.400 ;
        RECT 235.900 65.200 236.200 66.800 ;
        RECT 239.500 66.700 239.900 66.800 ;
        RECT 244.100 66.700 244.500 66.800 ;
        RECT 239.000 66.200 239.400 66.300 ;
        RECT 240.300 66.200 240.700 66.300 ;
        RECT 238.200 65.900 240.700 66.200 ;
        RECT 243.300 66.200 243.700 66.300 ;
        RECT 243.300 65.900 245.800 66.200 ;
        RECT 238.200 65.800 238.600 65.900 ;
        RECT 245.400 65.800 245.800 65.900 ;
        RECT 239.000 65.500 241.800 65.600 ;
        RECT 238.900 65.400 241.800 65.500 ;
        RECT 235.000 64.900 236.200 65.200 ;
        RECT 236.900 65.300 241.800 65.400 ;
        RECT 236.900 65.100 239.300 65.300 ;
        RECT 235.000 64.400 235.300 64.900 ;
        RECT 234.600 64.000 235.300 64.400 ;
        RECT 236.100 64.500 236.500 64.600 ;
        RECT 236.900 64.500 237.200 65.100 ;
        RECT 236.100 64.200 237.200 64.500 ;
        RECT 237.500 64.500 240.200 64.800 ;
        RECT 237.500 64.400 237.900 64.500 ;
        RECT 239.800 64.400 240.200 64.500 ;
        RECT 236.700 63.700 237.100 63.800 ;
        RECT 238.100 63.700 238.500 63.800 ;
        RECT 235.000 63.100 235.400 63.500 ;
        RECT 236.700 63.400 238.500 63.700 ;
        RECT 237.100 63.100 237.400 63.400 ;
        RECT 239.800 63.100 240.200 63.500 ;
        RECT 234.700 61.100 235.300 63.100 ;
        RECT 237.000 61.100 237.400 63.100 ;
        RECT 239.200 62.800 240.200 63.100 ;
        RECT 239.200 61.100 239.600 62.800 ;
        RECT 241.400 61.100 241.800 65.300 ;
        RECT 242.200 65.500 245.000 65.600 ;
        RECT 242.200 65.400 245.100 65.500 ;
        RECT 242.200 65.300 247.100 65.400 ;
        RECT 242.200 61.100 242.600 65.300 ;
        RECT 244.700 65.100 247.100 65.300 ;
        RECT 243.800 64.500 246.500 64.800 ;
        RECT 243.800 64.400 244.200 64.500 ;
        RECT 246.100 64.400 246.500 64.500 ;
        RECT 246.800 64.500 247.100 65.100 ;
        RECT 247.800 65.200 248.100 66.800 ;
        RECT 248.600 66.400 249.000 66.500 ;
        RECT 248.600 66.100 250.500 66.400 ;
        RECT 250.100 66.000 250.500 66.100 ;
        RECT 249.300 65.700 249.700 65.800 ;
        RECT 251.000 65.700 251.400 67.400 ;
        RECT 249.300 65.400 251.400 65.700 ;
        RECT 247.800 64.900 249.000 65.200 ;
        RECT 247.500 64.500 247.900 64.600 ;
        RECT 246.800 64.200 247.900 64.500 ;
        RECT 248.700 64.400 249.000 64.900 ;
        RECT 248.700 64.000 249.400 64.400 ;
        RECT 245.500 63.700 245.900 63.800 ;
        RECT 246.900 63.700 247.300 63.800 ;
        RECT 243.800 63.100 244.200 63.500 ;
        RECT 245.500 63.400 247.300 63.700 ;
        RECT 246.600 63.100 246.900 63.400 ;
        RECT 248.600 63.100 249.000 63.500 ;
        RECT 243.800 62.800 244.800 63.100 ;
        RECT 244.400 61.100 244.800 62.800 ;
        RECT 246.600 61.100 247.000 63.100 ;
        RECT 248.700 61.100 249.300 63.100 ;
        RECT 251.000 61.100 251.400 65.400 ;
        RECT 1.400 55.100 1.800 59.900 ;
        RECT 3.400 56.800 3.800 57.200 ;
        RECT 2.200 55.800 2.600 56.600 ;
        RECT 3.400 56.200 3.700 56.800 ;
        RECT 4.100 56.200 4.500 59.900 ;
        RECT 3.000 55.900 3.700 56.200 ;
        RECT 4.000 55.900 4.500 56.200 ;
        RECT 3.000 55.800 3.400 55.900 ;
        RECT 3.000 55.100 3.300 55.800 ;
        RECT 4.000 55.200 4.300 55.900 ;
        RECT 6.200 55.700 6.600 59.900 ;
        RECT 8.400 58.200 8.800 59.900 ;
        RECT 7.800 57.900 8.800 58.200 ;
        RECT 10.600 57.900 11.000 59.900 ;
        RECT 12.700 57.900 13.300 59.900 ;
        RECT 7.800 57.500 8.200 57.900 ;
        RECT 10.600 57.600 10.900 57.900 ;
        RECT 9.500 57.300 11.300 57.600 ;
        RECT 12.600 57.500 13.000 57.900 ;
        RECT 9.500 57.200 9.900 57.300 ;
        RECT 10.900 57.200 11.300 57.300 ;
        RECT 7.800 56.500 8.200 56.600 ;
        RECT 10.100 56.500 10.500 56.600 ;
        RECT 7.800 56.200 10.500 56.500 ;
        RECT 10.800 56.500 11.900 56.800 ;
        RECT 10.800 55.900 11.100 56.500 ;
        RECT 11.500 56.400 11.900 56.500 ;
        RECT 12.700 56.600 13.400 57.000 ;
        RECT 12.700 56.100 13.000 56.600 ;
        RECT 8.700 55.700 11.100 55.900 ;
        RECT 6.200 55.600 11.100 55.700 ;
        RECT 11.800 55.800 13.000 56.100 ;
        RECT 6.200 55.500 9.100 55.600 ;
        RECT 6.200 55.400 9.000 55.500 ;
        RECT 1.400 54.800 3.300 55.100 ;
        RECT 3.800 54.800 4.300 55.200 ;
        RECT 0.600 53.400 1.000 54.200 ;
        RECT 1.400 53.100 1.800 54.800 ;
        RECT 4.000 54.200 4.300 54.800 ;
        RECT 4.600 54.400 5.000 55.200 ;
        RECT 9.400 55.100 9.800 55.200 ;
        RECT 7.300 54.800 9.800 55.100 ;
        RECT 7.300 54.700 7.700 54.800 ;
        RECT 8.600 54.700 9.000 54.800 ;
        RECT 8.100 54.200 8.500 54.300 ;
        RECT 11.800 54.200 12.100 55.800 ;
        RECT 15.000 55.600 15.400 59.900 ;
        RECT 13.300 55.300 15.400 55.600 ;
        RECT 15.800 55.700 16.200 59.900 ;
        RECT 18.000 58.200 18.400 59.900 ;
        RECT 17.400 57.900 18.400 58.200 ;
        RECT 20.200 57.900 20.600 59.900 ;
        RECT 22.300 57.900 22.900 59.900 ;
        RECT 17.400 57.500 17.800 57.900 ;
        RECT 20.200 57.600 20.500 57.900 ;
        RECT 19.100 57.300 20.900 57.600 ;
        RECT 22.200 57.500 22.600 57.900 ;
        RECT 19.100 57.200 19.500 57.300 ;
        RECT 20.500 57.200 20.900 57.300 ;
        RECT 24.600 57.100 25.000 59.900 ;
        RECT 25.400 57.100 25.800 57.200 ;
        RECT 17.400 56.500 17.800 56.600 ;
        RECT 19.700 56.500 20.100 56.600 ;
        RECT 17.400 56.200 20.100 56.500 ;
        RECT 20.400 56.500 21.500 56.800 ;
        RECT 20.400 55.900 20.700 56.500 ;
        RECT 21.100 56.400 21.500 56.500 ;
        RECT 22.300 56.600 23.000 57.000 ;
        RECT 24.600 56.800 25.800 57.100 ;
        RECT 22.300 56.100 22.600 56.600 ;
        RECT 18.300 55.700 20.700 55.900 ;
        RECT 15.800 55.600 20.700 55.700 ;
        RECT 21.400 55.800 22.600 56.100 ;
        RECT 15.800 55.500 18.700 55.600 ;
        RECT 15.800 55.400 18.600 55.500 ;
        RECT 13.300 55.200 13.700 55.300 ;
        RECT 14.100 54.900 14.500 55.000 ;
        RECT 12.600 54.600 14.500 54.900 ;
        RECT 12.600 54.500 13.000 54.600 ;
        RECT 3.000 53.800 4.300 54.200 ;
        RECT 5.400 54.100 5.800 54.200 ;
        RECT 5.000 53.800 5.800 54.100 ;
        RECT 6.600 53.900 12.100 54.200 ;
        RECT 6.600 53.800 7.400 53.900 ;
        RECT 3.100 53.100 3.400 53.800 ;
        RECT 5.000 53.600 5.400 53.800 ;
        RECT 3.900 53.100 5.700 53.300 ;
        RECT 1.400 52.800 2.300 53.100 ;
        RECT 1.900 51.100 2.300 52.800 ;
        RECT 3.000 51.100 3.400 53.100 ;
        RECT 3.800 53.000 5.800 53.100 ;
        RECT 3.800 51.100 4.200 53.000 ;
        RECT 5.400 51.100 5.800 53.000 ;
        RECT 6.200 51.100 6.600 53.500 ;
        RECT 8.700 52.800 9.000 53.900 ;
        RECT 11.500 53.800 11.900 53.900 ;
        RECT 15.000 53.600 15.400 55.300 ;
        RECT 19.000 55.100 19.400 55.200 ;
        RECT 16.900 54.800 19.400 55.100 ;
        RECT 16.900 54.700 17.300 54.800 ;
        RECT 17.700 54.200 18.100 54.300 ;
        RECT 21.400 54.200 21.700 55.800 ;
        RECT 24.600 55.600 25.000 56.800 ;
        RECT 22.900 55.300 25.000 55.600 ;
        RECT 22.900 55.200 23.300 55.300 ;
        RECT 23.700 54.900 24.100 55.000 ;
        RECT 22.200 54.600 24.100 54.900 ;
        RECT 22.200 54.500 22.600 54.600 ;
        RECT 16.200 53.900 21.700 54.200 ;
        RECT 16.200 53.800 17.000 53.900 ;
        RECT 13.500 53.300 15.400 53.600 ;
        RECT 13.500 53.200 13.900 53.300 ;
        RECT 7.800 52.100 8.200 52.500 ;
        RECT 8.600 52.400 9.000 52.800 ;
        RECT 9.500 52.700 9.900 52.800 ;
        RECT 9.500 52.400 10.900 52.700 ;
        RECT 10.600 52.100 10.900 52.400 ;
        RECT 12.600 52.100 13.000 52.500 ;
        RECT 7.800 51.800 8.800 52.100 ;
        RECT 8.400 51.100 8.800 51.800 ;
        RECT 10.600 51.100 11.000 52.100 ;
        RECT 12.600 51.800 13.300 52.100 ;
        RECT 12.700 51.100 13.300 51.800 ;
        RECT 15.000 51.100 15.400 53.300 ;
        RECT 15.800 51.100 16.200 53.500 ;
        RECT 18.300 52.800 18.600 53.900 ;
        RECT 21.100 53.800 21.500 53.900 ;
        RECT 24.600 53.600 25.000 55.300 ;
        RECT 26.200 55.100 26.600 59.900 ;
        RECT 28.200 56.800 28.600 57.200 ;
        RECT 27.000 55.800 27.400 56.600 ;
        RECT 28.200 56.200 28.500 56.800 ;
        RECT 28.900 56.200 29.300 59.900 ;
        RECT 27.800 55.900 28.500 56.200 ;
        RECT 28.800 55.900 29.300 56.200 ;
        RECT 27.800 55.800 28.200 55.900 ;
        RECT 27.800 55.100 28.100 55.800 ;
        RECT 26.200 54.800 28.100 55.100 ;
        RECT 23.100 53.300 25.000 53.600 ;
        RECT 25.400 53.400 25.800 54.200 ;
        RECT 23.100 53.200 23.500 53.300 ;
        RECT 17.400 52.100 17.800 52.500 ;
        RECT 18.200 52.400 18.600 52.800 ;
        RECT 19.100 52.700 19.500 52.800 ;
        RECT 19.100 52.400 20.500 52.700 ;
        RECT 20.200 52.100 20.500 52.400 ;
        RECT 22.200 52.100 22.600 52.500 ;
        RECT 17.400 51.800 18.400 52.100 ;
        RECT 18.000 51.100 18.400 51.800 ;
        RECT 20.200 51.100 20.600 52.100 ;
        RECT 22.200 51.800 22.900 52.100 ;
        RECT 22.300 51.100 22.900 51.800 ;
        RECT 24.600 51.100 25.000 53.300 ;
        RECT 26.200 53.100 26.600 54.800 ;
        RECT 28.800 54.200 29.100 55.900 ;
        RECT 31.000 55.600 31.400 59.900 ;
        RECT 33.100 57.900 33.700 59.900 ;
        RECT 35.400 57.900 35.800 59.900 ;
        RECT 37.600 58.200 38.000 59.900 ;
        RECT 37.600 57.900 38.600 58.200 ;
        RECT 33.400 57.500 33.800 57.900 ;
        RECT 35.500 57.600 35.800 57.900 ;
        RECT 35.100 57.300 36.900 57.600 ;
        RECT 38.200 57.500 38.600 57.900 ;
        RECT 35.100 57.200 35.500 57.300 ;
        RECT 36.500 57.200 36.900 57.300 ;
        RECT 33.000 56.600 33.700 57.000 ;
        RECT 33.400 56.100 33.700 56.600 ;
        RECT 34.500 56.500 35.600 56.800 ;
        RECT 34.500 56.400 34.900 56.500 ;
        RECT 33.400 55.800 34.600 56.100 ;
        RECT 31.000 55.300 33.100 55.600 ;
        RECT 29.400 54.400 29.800 55.200 ;
        RECT 27.800 53.800 29.100 54.200 ;
        RECT 30.200 54.100 30.600 54.200 ;
        RECT 29.800 53.800 30.600 54.100 ;
        RECT 27.900 53.100 28.200 53.800 ;
        RECT 29.800 53.600 30.200 53.800 ;
        RECT 31.000 53.600 31.400 55.300 ;
        RECT 32.700 55.200 33.100 55.300 ;
        RECT 31.900 54.900 32.300 55.000 ;
        RECT 31.900 54.600 33.800 54.900 ;
        RECT 33.400 54.500 33.800 54.600 ;
        RECT 34.300 54.200 34.600 55.800 ;
        RECT 35.300 55.900 35.600 56.500 ;
        RECT 35.900 56.500 36.300 56.600 ;
        RECT 38.200 56.500 38.600 56.600 ;
        RECT 35.900 56.200 38.600 56.500 ;
        RECT 35.300 55.700 37.700 55.900 ;
        RECT 39.800 55.700 40.200 59.900 ;
        RECT 42.500 59.200 42.900 59.900 ;
        RECT 42.500 58.800 43.400 59.200 ;
        RECT 42.500 56.400 42.900 58.800 ;
        RECT 44.600 57.500 45.000 59.500 ;
        RECT 35.300 55.600 40.200 55.700 ;
        RECT 42.100 56.100 42.900 56.400 ;
        RECT 37.300 55.500 40.200 55.600 ;
        RECT 37.400 55.400 40.200 55.500 ;
        RECT 36.600 55.100 37.000 55.200 ;
        RECT 36.600 54.800 39.100 55.100 ;
        RECT 41.400 54.800 41.800 55.600 ;
        RECT 38.700 54.700 39.100 54.800 ;
        RECT 37.900 54.200 38.300 54.300 ;
        RECT 42.100 54.200 42.400 56.100 ;
        RECT 44.700 55.800 45.000 57.500 ;
        RECT 43.100 55.500 45.000 55.800 ;
        RECT 45.400 57.500 45.800 59.500 ;
        RECT 47.500 59.200 47.900 59.900 ;
        RECT 47.000 58.800 47.900 59.200 ;
        RECT 45.400 55.800 45.700 57.500 ;
        RECT 47.500 56.400 47.900 58.800 ;
        RECT 51.800 57.500 52.200 59.500 ;
        RECT 53.900 59.200 54.300 59.900 ;
        RECT 53.900 58.800 54.600 59.200 ;
        RECT 47.500 56.100 48.300 56.400 ;
        RECT 45.400 55.500 47.300 55.800 ;
        RECT 43.100 54.500 43.400 55.500 ;
        RECT 34.300 53.900 39.800 54.200 ;
        RECT 34.500 53.800 34.900 53.900 ;
        RECT 31.000 53.300 32.900 53.600 ;
        RECT 28.700 53.100 30.500 53.300 ;
        RECT 26.200 52.800 27.100 53.100 ;
        RECT 26.700 51.100 27.100 52.800 ;
        RECT 27.800 51.100 28.200 53.100 ;
        RECT 28.600 53.000 30.600 53.100 ;
        RECT 28.600 51.100 29.000 53.000 ;
        RECT 30.200 51.100 30.600 53.000 ;
        RECT 31.000 51.100 31.400 53.300 ;
        RECT 32.500 53.200 32.900 53.300 ;
        RECT 37.400 52.800 37.700 53.900 ;
        RECT 39.000 53.800 39.800 53.900 ;
        RECT 41.400 53.800 42.400 54.200 ;
        RECT 42.700 54.100 43.400 54.500 ;
        RECT 43.800 54.400 44.200 55.200 ;
        RECT 44.600 54.400 45.000 55.200 ;
        RECT 45.400 54.400 45.800 55.200 ;
        RECT 46.200 54.400 46.600 55.200 ;
        RECT 47.000 54.500 47.300 55.500 ;
        RECT 42.100 53.500 42.400 53.800 ;
        RECT 42.900 53.900 43.400 54.100 ;
        RECT 47.000 54.100 47.700 54.500 ;
        RECT 48.000 54.200 48.300 56.100 ;
        RECT 51.800 55.800 52.100 57.500 ;
        RECT 53.900 56.400 54.300 58.800 ;
        RECT 53.900 56.100 54.700 56.400 ;
        RECT 48.600 54.800 49.000 55.600 ;
        RECT 51.800 55.500 53.700 55.800 ;
        RECT 51.800 54.400 52.200 55.200 ;
        RECT 52.600 54.400 53.000 55.200 ;
        RECT 53.400 54.500 53.700 55.500 ;
        RECT 47.000 53.900 47.500 54.100 ;
        RECT 42.900 53.600 45.000 53.900 ;
        RECT 36.500 52.700 36.900 52.800 ;
        RECT 33.400 52.100 33.800 52.500 ;
        RECT 35.500 52.400 36.900 52.700 ;
        RECT 37.400 52.400 37.800 52.800 ;
        RECT 35.500 52.100 35.800 52.400 ;
        RECT 38.200 52.100 38.600 52.500 ;
        RECT 33.100 51.800 33.800 52.100 ;
        RECT 33.100 51.100 33.700 51.800 ;
        RECT 35.400 51.100 35.800 52.100 ;
        RECT 37.600 51.800 38.600 52.100 ;
        RECT 37.600 51.100 38.000 51.800 ;
        RECT 39.800 51.100 40.200 53.500 ;
        RECT 42.100 53.300 42.500 53.500 ;
        RECT 42.100 53.000 42.900 53.300 ;
        RECT 42.500 51.500 42.900 53.000 ;
        RECT 44.700 52.500 45.000 53.600 ;
        RECT 44.600 51.500 45.000 52.500 ;
        RECT 45.400 53.600 47.500 53.900 ;
        RECT 48.000 53.800 49.000 54.200 ;
        RECT 53.400 54.100 54.100 54.500 ;
        RECT 54.400 54.200 54.700 56.100 ;
        RECT 56.600 56.200 57.000 59.900 ;
        RECT 58.200 56.200 58.600 59.900 ;
        RECT 56.600 55.900 58.600 56.200 ;
        RECT 59.000 55.900 59.400 59.900 ;
        RECT 59.800 55.900 60.200 59.900 ;
        RECT 60.600 56.200 61.000 59.900 ;
        RECT 62.200 56.200 62.600 59.900 ;
        RECT 60.600 55.900 62.600 56.200 ;
        RECT 64.300 56.200 64.700 59.900 ;
        RECT 65.000 56.800 65.400 57.200 ;
        RECT 65.100 56.200 65.400 56.800 ;
        RECT 64.300 55.900 64.800 56.200 ;
        RECT 65.100 55.900 65.800 56.200 ;
        RECT 55.000 54.800 55.400 55.600 ;
        RECT 57.000 55.200 57.400 55.400 ;
        RECT 59.000 55.200 59.300 55.900 ;
        RECT 59.900 55.200 60.200 55.900 ;
        RECT 61.800 55.200 62.200 55.400 ;
        RECT 56.600 54.900 57.400 55.200 ;
        RECT 58.200 54.900 59.400 55.200 ;
        RECT 56.600 54.800 57.000 54.900 ;
        RECT 53.400 53.900 53.900 54.100 ;
        RECT 45.400 52.500 45.700 53.600 ;
        RECT 48.000 53.500 48.300 53.800 ;
        RECT 47.900 53.300 48.300 53.500 ;
        RECT 47.500 53.000 48.300 53.300 ;
        RECT 51.800 53.600 53.900 53.900 ;
        RECT 54.400 53.800 55.400 54.200 ;
        RECT 57.400 53.800 57.800 54.600 ;
        RECT 45.400 51.500 45.800 52.500 ;
        RECT 47.500 51.500 47.900 53.000 ;
        RECT 51.800 52.500 52.100 53.600 ;
        RECT 54.400 53.500 54.700 53.800 ;
        RECT 54.300 53.300 54.700 53.500 ;
        RECT 53.900 53.000 54.700 53.300 ;
        RECT 58.200 53.100 58.500 54.900 ;
        RECT 59.000 54.800 59.400 54.900 ;
        RECT 59.800 54.900 61.000 55.200 ;
        RECT 61.800 54.900 62.600 55.200 ;
        RECT 59.800 54.800 60.200 54.900 ;
        RECT 59.000 53.100 59.400 53.200 ;
        RECT 59.800 53.100 60.200 53.200 ;
        RECT 60.700 53.100 61.000 54.900 ;
        RECT 62.200 54.800 62.600 54.900 ;
        RECT 61.400 53.800 61.800 54.600 ;
        RECT 63.800 54.400 64.200 55.200 ;
        RECT 64.500 54.200 64.800 55.900 ;
        RECT 65.400 55.800 65.800 55.900 ;
        RECT 66.200 55.800 66.600 56.600 ;
        RECT 65.400 55.100 65.700 55.800 ;
        RECT 67.000 55.100 67.400 59.900 ;
        RECT 68.600 55.700 69.000 59.900 ;
        RECT 70.800 58.200 71.200 59.900 ;
        RECT 70.200 57.900 71.200 58.200 ;
        RECT 73.000 57.900 73.400 59.900 ;
        RECT 75.100 57.900 75.700 59.900 ;
        RECT 70.200 57.500 70.600 57.900 ;
        RECT 73.000 57.600 73.300 57.900 ;
        RECT 71.900 57.300 73.700 57.600 ;
        RECT 75.000 57.500 75.400 57.900 ;
        RECT 71.900 57.200 72.300 57.300 ;
        RECT 73.300 57.200 73.700 57.300 ;
        RECT 70.200 56.500 70.600 56.600 ;
        RECT 72.500 56.500 72.900 56.600 ;
        RECT 70.200 56.200 72.900 56.500 ;
        RECT 73.200 56.500 74.300 56.800 ;
        RECT 73.200 55.900 73.500 56.500 ;
        RECT 73.900 56.400 74.300 56.500 ;
        RECT 75.100 56.600 75.800 57.000 ;
        RECT 75.100 56.100 75.400 56.600 ;
        RECT 71.100 55.700 73.500 55.900 ;
        RECT 68.600 55.600 73.500 55.700 ;
        RECT 74.200 55.800 75.400 56.100 ;
        RECT 68.600 55.500 71.500 55.600 ;
        RECT 68.600 55.400 71.400 55.500 ;
        RECT 71.800 55.100 72.200 55.200 ;
        RECT 65.400 54.800 67.400 55.100 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 64.500 54.100 65.800 54.200 ;
        RECT 66.200 54.100 66.600 54.200 ;
        RECT 63.000 53.800 63.800 54.100 ;
        RECT 64.500 53.800 66.600 54.100 ;
        RECT 63.400 53.600 63.800 53.800 ;
        RECT 63.100 53.100 64.900 53.300 ;
        RECT 65.400 53.100 65.700 53.800 ;
        RECT 67.000 53.100 67.400 54.800 ;
        RECT 69.700 54.800 72.200 55.100 ;
        RECT 69.700 54.700 70.100 54.800 ;
        RECT 71.000 54.700 71.400 54.800 ;
        RECT 70.500 54.200 70.900 54.300 ;
        RECT 74.200 54.200 74.500 55.800 ;
        RECT 77.400 55.600 77.800 59.900 ;
        RECT 80.100 56.400 80.500 59.900 ;
        RECT 82.200 57.500 82.600 59.500 ;
        RECT 84.900 59.200 85.300 59.900 ;
        RECT 84.600 58.800 85.300 59.200 ;
        RECT 79.700 56.100 80.500 56.400 ;
        RECT 75.700 55.300 77.800 55.600 ;
        RECT 75.700 55.200 76.100 55.300 ;
        RECT 76.500 54.900 76.900 55.000 ;
        RECT 75.000 54.600 76.900 54.900 ;
        RECT 75.000 54.500 75.400 54.600 ;
        RECT 67.800 53.400 68.200 54.200 ;
        RECT 69.000 53.900 74.500 54.200 ;
        RECT 69.000 53.800 69.800 53.900 ;
        RECT 51.800 51.500 52.200 52.500 ;
        RECT 53.900 51.500 54.300 53.000 ;
        RECT 58.200 51.100 58.600 53.100 ;
        RECT 59.000 52.800 60.200 53.100 ;
        RECT 58.900 52.400 59.300 52.800 ;
        RECT 59.900 52.400 60.300 52.800 ;
        RECT 60.600 51.100 61.000 53.100 ;
        RECT 63.000 53.000 65.000 53.100 ;
        RECT 63.000 51.100 63.400 53.000 ;
        RECT 64.600 51.100 65.000 53.000 ;
        RECT 65.400 51.100 65.800 53.100 ;
        RECT 66.500 52.800 67.400 53.100 ;
        RECT 66.500 51.100 66.900 52.800 ;
        RECT 68.600 51.100 69.000 53.500 ;
        RECT 71.100 52.800 71.400 53.900 ;
        RECT 73.900 53.800 74.300 53.900 ;
        RECT 77.400 53.600 77.800 55.300 ;
        RECT 79.000 54.800 79.400 55.600 ;
        RECT 79.700 55.200 80.000 56.100 ;
        RECT 82.300 55.800 82.600 57.500 ;
        RECT 84.900 56.400 85.300 58.800 ;
        RECT 87.000 57.500 87.400 59.500 ;
        RECT 80.700 55.500 82.600 55.800 ;
        RECT 84.500 56.100 85.300 56.400 ;
        RECT 79.700 54.800 80.200 55.200 ;
        RECT 79.700 54.200 80.000 54.800 ;
        RECT 80.700 54.500 81.000 55.500 ;
        RECT 79.000 53.800 80.000 54.200 ;
        RECT 80.300 54.100 81.000 54.500 ;
        RECT 81.400 54.400 81.800 55.200 ;
        RECT 82.200 54.400 82.600 55.200 ;
        RECT 83.800 54.800 84.200 55.600 ;
        RECT 84.500 54.200 84.800 56.100 ;
        RECT 87.100 55.800 87.400 57.500 ;
        RECT 85.500 55.500 87.400 55.800 ;
        RECT 87.800 57.500 88.200 59.500 ;
        RECT 89.900 59.200 90.300 59.900 ;
        RECT 89.400 58.800 90.300 59.200 ;
        RECT 87.800 55.800 88.100 57.500 ;
        RECT 89.900 56.400 90.300 58.800 ;
        RECT 92.600 57.500 93.000 59.500 ;
        RECT 89.900 56.100 90.700 56.400 ;
        RECT 87.800 55.500 89.700 55.800 ;
        RECT 85.500 54.500 85.800 55.500 ;
        RECT 75.900 53.300 77.800 53.600 ;
        RECT 75.900 53.200 76.300 53.300 ;
        RECT 70.200 52.100 70.600 52.500 ;
        RECT 71.000 52.400 71.400 52.800 ;
        RECT 71.900 52.700 72.300 52.800 ;
        RECT 71.900 52.400 73.300 52.700 ;
        RECT 73.000 52.100 73.300 52.400 ;
        RECT 75.000 52.100 75.400 52.500 ;
        RECT 70.200 51.800 71.200 52.100 ;
        RECT 70.800 51.100 71.200 51.800 ;
        RECT 73.000 51.100 73.400 52.100 ;
        RECT 75.000 51.800 75.700 52.100 ;
        RECT 75.100 51.100 75.700 51.800 ;
        RECT 77.400 51.100 77.800 53.300 ;
        RECT 79.700 53.500 80.000 53.800 ;
        RECT 80.500 53.900 81.000 54.100 ;
        RECT 80.500 53.600 82.600 53.900 ;
        RECT 83.800 53.800 84.800 54.200 ;
        RECT 85.100 54.100 85.800 54.500 ;
        RECT 86.200 54.400 86.600 55.200 ;
        RECT 87.000 54.400 87.400 55.200 ;
        RECT 87.800 54.400 88.200 55.200 ;
        RECT 88.600 54.400 89.000 55.200 ;
        RECT 89.400 54.500 89.700 55.500 ;
        RECT 79.700 53.300 80.100 53.500 ;
        RECT 79.700 53.000 80.500 53.300 ;
        RECT 80.100 51.500 80.500 53.000 ;
        RECT 82.300 52.500 82.600 53.600 ;
        RECT 84.500 53.500 84.800 53.800 ;
        RECT 85.300 53.900 85.800 54.100 ;
        RECT 89.400 54.100 90.100 54.500 ;
        RECT 90.400 54.200 90.700 56.100 ;
        RECT 92.600 55.800 92.900 57.500 ;
        RECT 94.700 56.400 95.100 59.900 ;
        RECT 94.700 56.100 95.500 56.400 ;
        RECT 91.000 54.800 91.400 55.600 ;
        RECT 92.600 55.500 94.500 55.800 ;
        RECT 92.600 54.400 93.000 55.200 ;
        RECT 93.400 54.400 93.800 55.200 ;
        RECT 94.200 54.500 94.500 55.500 ;
        RECT 95.200 55.200 95.500 56.100 ;
        RECT 99.000 55.600 99.400 59.900 ;
        RECT 101.100 57.900 101.700 59.900 ;
        RECT 103.400 57.900 103.800 59.900 ;
        RECT 105.600 58.200 106.000 59.900 ;
        RECT 105.600 57.900 106.600 58.200 ;
        RECT 101.400 57.500 101.800 57.900 ;
        RECT 103.500 57.600 103.800 57.900 ;
        RECT 103.100 57.300 104.900 57.600 ;
        RECT 106.200 57.500 106.600 57.900 ;
        RECT 103.100 57.200 103.500 57.300 ;
        RECT 104.500 57.200 104.900 57.300 ;
        RECT 101.000 56.600 101.700 57.000 ;
        RECT 101.400 56.100 101.700 56.600 ;
        RECT 102.500 56.500 103.600 56.800 ;
        RECT 102.500 56.400 102.900 56.500 ;
        RECT 101.400 55.800 102.600 56.100 ;
        RECT 95.000 54.800 95.500 55.200 ;
        RECT 95.800 55.100 96.200 55.600 ;
        RECT 99.000 55.300 101.100 55.600 ;
        RECT 96.600 55.100 97.000 55.200 ;
        RECT 95.800 54.800 97.000 55.100 ;
        RECT 89.400 53.900 89.900 54.100 ;
        RECT 85.300 53.600 87.400 53.900 ;
        RECT 84.500 53.300 84.900 53.500 ;
        RECT 84.500 53.000 85.300 53.300 ;
        RECT 82.200 51.500 82.600 52.500 ;
        RECT 84.900 51.500 85.300 53.000 ;
        RECT 87.100 52.500 87.400 53.600 ;
        RECT 87.000 51.500 87.400 52.500 ;
        RECT 87.800 53.600 89.900 53.900 ;
        RECT 90.400 53.800 91.400 54.200 ;
        RECT 94.200 54.100 94.900 54.500 ;
        RECT 95.200 54.200 95.500 54.800 ;
        RECT 94.200 53.900 94.700 54.100 ;
        RECT 87.800 52.500 88.100 53.600 ;
        RECT 90.400 53.500 90.700 53.800 ;
        RECT 90.300 53.300 90.700 53.500 ;
        RECT 89.900 53.000 90.700 53.300 ;
        RECT 92.600 53.600 94.700 53.900 ;
        RECT 95.200 53.800 96.200 54.200 ;
        RECT 87.800 51.500 88.200 52.500 ;
        RECT 89.900 51.500 90.300 53.000 ;
        RECT 92.600 52.500 92.900 53.600 ;
        RECT 95.200 53.500 95.500 53.800 ;
        RECT 95.100 53.300 95.500 53.500 ;
        RECT 94.700 53.000 95.500 53.300 ;
        RECT 99.000 53.600 99.400 55.300 ;
        RECT 100.700 55.200 101.100 55.300 ;
        RECT 99.900 54.900 100.300 55.000 ;
        RECT 99.900 54.600 101.800 54.900 ;
        RECT 101.400 54.500 101.800 54.600 ;
        RECT 102.300 54.200 102.600 55.800 ;
        RECT 103.300 55.900 103.600 56.500 ;
        RECT 103.900 56.500 104.300 56.600 ;
        RECT 106.200 56.500 106.600 56.600 ;
        RECT 103.900 56.200 106.600 56.500 ;
        RECT 103.300 55.700 105.700 55.900 ;
        RECT 107.800 55.700 108.200 59.900 ;
        RECT 103.300 55.600 108.200 55.700 ;
        RECT 105.300 55.500 108.200 55.600 ;
        RECT 105.400 55.400 108.200 55.500 ;
        RECT 104.600 55.100 105.000 55.200 ;
        RECT 109.400 55.100 109.800 59.900 ;
        RECT 111.400 56.800 111.800 57.200 ;
        RECT 110.200 55.800 110.600 56.600 ;
        RECT 111.400 56.200 111.700 56.800 ;
        RECT 112.100 56.200 112.500 59.900 ;
        RECT 115.500 59.200 115.900 59.900 ;
        RECT 115.500 58.800 116.200 59.200 ;
        RECT 115.500 56.300 115.900 58.800 ;
        RECT 111.000 55.900 111.700 56.200 ;
        RECT 112.000 55.900 112.500 56.200 ;
        RECT 115.000 55.900 115.900 56.300 ;
        RECT 111.000 55.800 111.400 55.900 ;
        RECT 111.000 55.100 111.300 55.800 ;
        RECT 104.600 54.800 107.100 55.100 ;
        RECT 105.400 54.700 105.800 54.800 ;
        RECT 106.700 54.700 107.100 54.800 ;
        RECT 109.400 54.800 111.300 55.100 ;
        RECT 105.900 54.200 106.300 54.300 ;
        RECT 102.300 53.900 107.800 54.200 ;
        RECT 102.500 53.800 102.900 53.900 ;
        RECT 99.000 53.300 100.900 53.600 ;
        RECT 92.600 51.500 93.000 52.500 ;
        RECT 94.700 51.500 95.100 53.000 ;
        RECT 99.000 51.100 99.400 53.300 ;
        RECT 100.500 53.200 100.900 53.300 ;
        RECT 105.400 52.800 105.700 53.900 ;
        RECT 107.000 53.800 107.800 53.900 ;
        RECT 104.500 52.700 104.900 52.800 ;
        RECT 101.400 52.100 101.800 52.500 ;
        RECT 103.500 52.400 104.900 52.700 ;
        RECT 105.400 52.400 105.800 52.800 ;
        RECT 103.500 52.100 103.800 52.400 ;
        RECT 106.200 52.100 106.600 52.500 ;
        RECT 101.100 51.800 101.800 52.100 ;
        RECT 101.100 51.100 101.700 51.800 ;
        RECT 103.400 51.100 103.800 52.100 ;
        RECT 105.600 51.800 106.600 52.100 ;
        RECT 105.600 51.100 106.000 51.800 ;
        RECT 107.800 51.100 108.200 53.500 ;
        RECT 108.600 53.400 109.000 54.200 ;
        RECT 109.400 53.100 109.800 54.800 ;
        RECT 112.000 54.200 112.300 55.900 ;
        RECT 112.600 54.400 113.000 55.200 ;
        RECT 115.100 54.200 115.400 55.900 ;
        RECT 116.600 55.800 117.000 56.600 ;
        RECT 115.800 55.100 116.200 55.600 ;
        RECT 117.400 55.100 117.800 59.900 ;
        RECT 118.200 56.800 118.600 57.200 ;
        RECT 118.200 56.100 118.500 56.800 ;
        RECT 119.000 56.100 119.400 59.900 ;
        RECT 118.200 55.800 119.400 56.100 ;
        RECT 115.800 54.800 117.800 55.100 ;
        RECT 110.200 54.100 110.600 54.200 ;
        RECT 111.000 54.100 112.300 54.200 ;
        RECT 113.400 54.100 113.800 54.200 ;
        RECT 110.200 53.800 112.300 54.100 ;
        RECT 113.000 53.800 113.800 54.100 ;
        RECT 115.000 53.800 115.400 54.200 ;
        RECT 111.100 53.100 111.400 53.800 ;
        RECT 113.000 53.600 113.400 53.800 ;
        RECT 111.900 53.100 113.700 53.300 ;
        RECT 109.400 52.800 110.300 53.100 ;
        RECT 109.900 51.100 110.300 52.800 ;
        RECT 111.000 51.100 111.400 53.100 ;
        RECT 111.800 53.000 113.800 53.100 ;
        RECT 111.800 51.100 112.200 53.000 ;
        RECT 113.400 51.100 113.800 53.000 ;
        RECT 114.200 52.400 114.600 53.200 ;
        RECT 115.100 52.100 115.400 53.800 ;
        RECT 117.400 53.100 117.800 54.800 ;
        RECT 118.200 53.400 118.600 54.200 ;
        RECT 115.000 51.100 115.400 52.100 ;
        RECT 116.900 52.800 117.800 53.100 ;
        RECT 116.900 51.100 117.300 52.800 ;
        RECT 119.000 51.100 119.400 55.800 ;
        RECT 120.600 57.500 121.000 59.500 ;
        RECT 122.700 59.200 123.100 59.900 ;
        RECT 122.700 58.800 123.400 59.200 ;
        RECT 120.600 55.800 120.900 57.500 ;
        RECT 122.700 56.400 123.100 58.800 ;
        RECT 122.700 56.100 123.500 56.400 ;
        RECT 120.600 55.500 122.500 55.800 ;
        RECT 120.600 54.400 121.000 55.200 ;
        RECT 121.400 54.400 121.800 55.200 ;
        RECT 122.200 54.500 122.500 55.500 ;
        RECT 122.200 54.100 122.900 54.500 ;
        RECT 123.200 54.200 123.500 56.100 ;
        RECT 125.400 55.800 125.800 56.600 ;
        RECT 126.200 56.100 126.600 59.900 ;
        RECT 128.200 56.800 128.600 57.200 ;
        RECT 128.200 56.200 128.500 56.800 ;
        RECT 128.900 56.200 129.300 59.900 ;
        RECT 127.800 56.100 128.500 56.200 ;
        RECT 126.200 55.900 128.500 56.100 ;
        RECT 128.800 55.900 129.300 56.200 ;
        RECT 126.200 55.800 128.200 55.900 ;
        RECT 123.800 54.800 124.200 55.600 ;
        RECT 122.200 53.900 122.700 54.100 ;
        RECT 120.600 53.600 122.700 53.900 ;
        RECT 123.200 53.800 124.200 54.200 ;
        RECT 119.800 52.400 120.200 53.200 ;
        RECT 120.600 52.500 120.900 53.600 ;
        RECT 123.200 53.500 123.500 53.800 ;
        RECT 123.100 53.300 123.500 53.500 ;
        RECT 122.700 53.000 123.500 53.300 ;
        RECT 126.200 53.100 126.600 55.800 ;
        RECT 127.800 55.100 128.200 55.200 ;
        RECT 128.800 55.100 129.100 55.900 ;
        RECT 131.000 55.700 131.400 59.900 ;
        RECT 133.200 58.200 133.600 59.900 ;
        RECT 132.600 57.900 133.600 58.200 ;
        RECT 135.400 57.900 135.800 59.900 ;
        RECT 137.500 57.900 138.100 59.900 ;
        RECT 132.600 57.500 133.000 57.900 ;
        RECT 135.400 57.600 135.700 57.900 ;
        RECT 134.300 57.300 136.100 57.600 ;
        RECT 137.400 57.500 137.800 57.900 ;
        RECT 134.300 57.200 134.700 57.300 ;
        RECT 135.700 57.200 136.100 57.300 ;
        RECT 132.600 56.500 133.000 56.600 ;
        RECT 134.900 56.500 135.300 56.600 ;
        RECT 132.600 56.200 135.300 56.500 ;
        RECT 135.600 56.500 136.700 56.800 ;
        RECT 135.600 55.900 135.900 56.500 ;
        RECT 136.300 56.400 136.700 56.500 ;
        RECT 137.500 56.600 138.200 57.000 ;
        RECT 137.500 56.100 137.800 56.600 ;
        RECT 133.500 55.700 135.900 55.900 ;
        RECT 131.000 55.600 135.900 55.700 ;
        RECT 136.600 55.800 137.800 56.100 ;
        RECT 131.000 55.500 133.900 55.600 ;
        RECT 131.000 55.400 133.800 55.500 ;
        RECT 127.800 54.800 129.100 55.100 ;
        RECT 128.800 54.200 129.100 54.800 ;
        RECT 129.400 54.400 129.800 55.200 ;
        RECT 134.200 55.100 134.600 55.200 ;
        RECT 132.100 54.800 134.600 55.100 ;
        RECT 132.100 54.700 132.500 54.800 ;
        RECT 133.400 54.700 133.800 54.800 ;
        RECT 132.900 54.200 133.300 54.300 ;
        RECT 136.600 54.200 136.900 55.800 ;
        RECT 139.800 55.600 140.200 59.900 ;
        RECT 140.600 56.200 141.000 59.900 ;
        RECT 142.200 56.200 142.600 59.900 ;
        RECT 140.600 55.900 142.600 56.200 ;
        RECT 143.000 55.900 143.400 59.900 ;
        RECT 144.100 56.300 144.500 59.900 ;
        RECT 148.100 56.400 148.500 59.900 ;
        RECT 150.200 57.500 150.600 59.500 ;
        RECT 144.100 55.900 145.000 56.300 ;
        RECT 147.700 56.100 148.500 56.400 ;
        RECT 138.100 55.300 140.200 55.600 ;
        RECT 138.100 55.200 138.500 55.300 ;
        RECT 138.900 54.900 139.300 55.000 ;
        RECT 137.400 54.600 139.300 54.900 ;
        RECT 137.400 54.500 137.800 54.600 ;
        RECT 127.000 53.400 127.400 54.200 ;
        RECT 127.800 53.800 129.100 54.200 ;
        RECT 130.200 54.100 130.600 54.200 ;
        RECT 129.800 53.800 130.600 54.100 ;
        RECT 131.400 53.900 136.900 54.200 ;
        RECT 131.400 53.800 132.200 53.900 ;
        RECT 127.900 53.100 128.200 53.800 ;
        RECT 129.800 53.600 130.200 53.800 ;
        RECT 128.700 53.100 130.500 53.300 ;
        RECT 120.600 51.500 121.000 52.500 ;
        RECT 122.700 51.500 123.100 53.000 ;
        RECT 125.700 52.800 126.600 53.100 ;
        RECT 125.700 51.100 126.100 52.800 ;
        RECT 127.800 51.100 128.200 53.100 ;
        RECT 128.600 53.000 130.600 53.100 ;
        RECT 128.600 51.100 129.000 53.000 ;
        RECT 130.200 51.100 130.600 53.000 ;
        RECT 131.000 51.100 131.400 53.500 ;
        RECT 133.500 53.200 133.800 53.900 ;
        RECT 136.300 53.800 136.700 53.900 ;
        RECT 139.800 53.600 140.200 55.300 ;
        RECT 141.000 55.200 141.400 55.400 ;
        RECT 143.000 55.200 143.300 55.900 ;
        RECT 140.600 54.900 141.400 55.200 ;
        RECT 142.200 54.900 143.400 55.200 ;
        RECT 140.600 54.800 141.000 54.900 ;
        RECT 141.400 53.800 141.800 54.600 ;
        RECT 138.300 53.300 140.200 53.600 ;
        RECT 138.300 53.200 138.700 53.300 ;
        RECT 132.600 52.100 133.000 52.500 ;
        RECT 133.400 52.400 133.800 53.200 ;
        RECT 134.300 52.700 134.700 52.800 ;
        RECT 134.300 52.400 135.700 52.700 ;
        RECT 135.400 52.100 135.700 52.400 ;
        RECT 137.400 52.100 137.800 52.500 ;
        RECT 132.600 51.800 133.600 52.100 ;
        RECT 133.200 51.100 133.600 51.800 ;
        RECT 135.400 51.100 135.800 52.100 ;
        RECT 137.400 51.800 138.100 52.100 ;
        RECT 137.500 51.100 138.100 51.800 ;
        RECT 139.800 51.100 140.200 53.300 ;
        RECT 142.200 53.100 142.500 54.900 ;
        RECT 143.000 54.800 143.400 54.900 ;
        RECT 143.800 54.800 144.200 55.600 ;
        RECT 144.600 54.200 144.900 55.900 ;
        RECT 146.200 55.100 146.600 55.200 ;
        RECT 147.000 55.100 147.400 55.600 ;
        RECT 146.200 54.800 147.400 55.100 ;
        RECT 147.700 54.200 148.000 56.100 ;
        RECT 150.300 55.800 150.600 57.500 ;
        RECT 153.900 56.200 154.300 59.900 ;
        RECT 154.600 56.800 155.000 57.200 ;
        RECT 154.700 56.200 155.000 56.800 ;
        RECT 153.900 55.900 154.400 56.200 ;
        RECT 154.700 55.900 155.400 56.200 ;
        RECT 148.700 55.500 150.600 55.800 ;
        RECT 148.700 54.500 149.000 55.500 ;
        RECT 144.600 53.800 145.000 54.200 ;
        RECT 146.200 54.100 146.600 54.200 ;
        RECT 147.000 54.100 148.000 54.200 ;
        RECT 148.300 54.100 149.000 54.500 ;
        RECT 149.400 54.400 149.800 55.200 ;
        RECT 150.200 54.400 150.600 55.200 ;
        RECT 153.400 54.400 153.800 55.200 ;
        RECT 154.100 54.200 154.400 55.900 ;
        RECT 155.000 55.800 155.400 55.900 ;
        RECT 155.800 55.800 156.200 56.600 ;
        RECT 155.000 55.100 155.300 55.800 ;
        RECT 156.600 55.100 157.000 59.900 ;
        RECT 158.200 55.700 158.600 59.900 ;
        RECT 160.400 58.200 160.800 59.900 ;
        RECT 159.800 57.900 160.800 58.200 ;
        RECT 162.600 57.900 163.000 59.900 ;
        RECT 164.700 57.900 165.300 59.900 ;
        RECT 159.800 57.500 160.200 57.900 ;
        RECT 162.600 57.600 162.900 57.900 ;
        RECT 161.500 57.300 163.300 57.600 ;
        RECT 164.600 57.500 165.000 57.900 ;
        RECT 161.500 57.200 161.900 57.300 ;
        RECT 162.900 57.200 163.300 57.300 ;
        RECT 159.800 56.500 160.200 56.600 ;
        RECT 162.100 56.500 162.500 56.600 ;
        RECT 159.800 56.200 162.500 56.500 ;
        RECT 162.800 56.500 163.900 56.800 ;
        RECT 162.800 55.900 163.100 56.500 ;
        RECT 163.500 56.400 163.900 56.500 ;
        RECT 164.700 56.600 165.400 57.000 ;
        RECT 164.700 56.100 165.000 56.600 ;
        RECT 160.700 55.700 163.100 55.900 ;
        RECT 158.200 55.600 163.100 55.700 ;
        RECT 163.800 55.800 165.000 56.100 ;
        RECT 158.200 55.500 161.100 55.600 ;
        RECT 158.200 55.400 161.000 55.500 ;
        RECT 161.400 55.100 161.800 55.200 ;
        RECT 155.000 54.800 157.000 55.100 ;
        RECT 146.200 53.800 148.000 54.100 ;
        RECT 143.000 53.100 143.400 53.200 ;
        RECT 144.600 53.100 144.900 53.800 ;
        RECT 147.700 53.500 148.000 53.800 ;
        RECT 148.500 53.900 149.000 54.100 ;
        RECT 152.600 54.100 153.000 54.200 ;
        RECT 148.500 53.600 150.600 53.900 ;
        RECT 152.600 53.800 153.400 54.100 ;
        RECT 154.100 53.800 155.400 54.200 ;
        RECT 153.000 53.600 153.400 53.800 ;
        RECT 147.700 53.300 148.100 53.500 ;
        RECT 142.200 51.100 142.600 53.100 ;
        RECT 143.000 52.800 144.900 53.100 ;
        RECT 142.900 52.400 143.300 52.800 ;
        RECT 144.600 52.100 144.900 52.800 ;
        RECT 145.400 52.400 145.800 53.200 ;
        RECT 147.700 53.000 148.500 53.300 ;
        RECT 144.600 51.100 145.000 52.100 ;
        RECT 148.100 51.500 148.500 53.000 ;
        RECT 150.300 52.500 150.600 53.600 ;
        RECT 152.700 53.100 154.500 53.300 ;
        RECT 155.000 53.100 155.300 53.800 ;
        RECT 156.600 53.100 157.000 54.800 ;
        RECT 159.300 54.800 161.800 55.100 ;
        RECT 159.300 54.700 159.700 54.800 ;
        RECT 160.600 54.700 161.000 54.800 ;
        RECT 160.100 54.200 160.500 54.300 ;
        RECT 163.800 54.200 164.100 55.800 ;
        RECT 167.000 55.600 167.400 59.900 ;
        RECT 165.300 55.300 167.400 55.600 ;
        RECT 165.300 55.200 165.700 55.300 ;
        RECT 166.100 54.900 166.500 55.000 ;
        RECT 164.600 54.600 166.500 54.900 ;
        RECT 164.600 54.500 165.000 54.600 ;
        RECT 157.400 53.400 157.800 54.200 ;
        RECT 158.600 53.900 164.100 54.200 ;
        RECT 158.600 53.800 159.400 53.900 ;
        RECT 150.200 51.500 150.600 52.500 ;
        RECT 152.600 53.000 154.600 53.100 ;
        RECT 152.600 51.100 153.000 53.000 ;
        RECT 154.200 51.100 154.600 53.000 ;
        RECT 155.000 51.100 155.400 53.100 ;
        RECT 156.100 52.800 157.000 53.100 ;
        RECT 156.100 51.100 156.500 52.800 ;
        RECT 158.200 51.100 158.600 53.500 ;
        RECT 160.700 52.800 161.000 53.900 ;
        RECT 163.500 53.800 163.900 53.900 ;
        RECT 167.000 53.600 167.400 55.300 ;
        RECT 165.500 53.300 167.400 53.600 ;
        RECT 165.500 53.200 165.900 53.300 ;
        RECT 159.800 52.100 160.200 52.500 ;
        RECT 160.600 52.400 161.000 52.800 ;
        RECT 161.500 52.700 161.900 52.800 ;
        RECT 161.500 52.400 162.900 52.700 ;
        RECT 162.600 52.100 162.900 52.400 ;
        RECT 164.600 52.100 165.000 52.500 ;
        RECT 159.800 51.800 160.800 52.100 ;
        RECT 160.400 51.100 160.800 51.800 ;
        RECT 162.600 51.100 163.000 52.100 ;
        RECT 164.600 51.800 165.300 52.100 ;
        RECT 164.700 51.100 165.300 51.800 ;
        RECT 167.000 51.100 167.400 53.300 ;
        RECT 167.800 55.600 168.200 59.900 ;
        RECT 169.900 57.900 170.500 59.900 ;
        RECT 172.200 57.900 172.600 59.900 ;
        RECT 174.400 58.200 174.800 59.900 ;
        RECT 174.400 57.900 175.400 58.200 ;
        RECT 170.200 57.500 170.600 57.900 ;
        RECT 172.300 57.600 172.600 57.900 ;
        RECT 171.900 57.300 173.700 57.600 ;
        RECT 175.000 57.500 175.400 57.900 ;
        RECT 171.900 57.200 172.300 57.300 ;
        RECT 173.300 57.200 173.700 57.300 ;
        RECT 169.800 56.600 170.500 57.000 ;
        RECT 170.200 56.100 170.500 56.600 ;
        RECT 171.300 56.500 172.400 56.800 ;
        RECT 171.300 56.400 171.700 56.500 ;
        RECT 170.200 55.800 171.400 56.100 ;
        RECT 167.800 55.300 169.900 55.600 ;
        RECT 167.800 53.600 168.200 55.300 ;
        RECT 169.500 55.200 169.900 55.300 ;
        RECT 168.700 54.900 169.100 55.000 ;
        RECT 168.700 54.600 170.600 54.900 ;
        RECT 170.200 54.500 170.600 54.600 ;
        RECT 171.100 54.200 171.400 55.800 ;
        RECT 172.100 55.900 172.400 56.500 ;
        RECT 172.700 56.500 173.100 56.600 ;
        RECT 175.000 56.500 175.400 56.600 ;
        RECT 172.700 56.200 175.400 56.500 ;
        RECT 172.100 55.700 174.500 55.900 ;
        RECT 176.600 55.700 177.000 59.900 ;
        RECT 172.100 55.600 177.000 55.700 ;
        RECT 174.100 55.500 177.000 55.600 ;
        RECT 174.200 55.400 177.000 55.500 ;
        RECT 177.400 55.700 177.800 59.900 ;
        RECT 179.600 58.200 180.000 59.900 ;
        RECT 179.000 57.900 180.000 58.200 ;
        RECT 181.800 57.900 182.200 59.900 ;
        RECT 183.900 57.900 184.500 59.900 ;
        RECT 179.000 57.500 179.400 57.900 ;
        RECT 181.800 57.600 182.100 57.900 ;
        RECT 180.700 57.300 182.500 57.600 ;
        RECT 183.800 57.500 184.200 57.900 ;
        RECT 180.700 57.200 181.100 57.300 ;
        RECT 182.100 57.200 182.500 57.300 ;
        RECT 179.000 56.500 179.400 56.600 ;
        RECT 181.300 56.500 181.700 56.600 ;
        RECT 179.000 56.200 181.700 56.500 ;
        RECT 182.000 56.500 183.100 56.800 ;
        RECT 182.000 55.900 182.300 56.500 ;
        RECT 182.700 56.400 183.100 56.500 ;
        RECT 183.900 56.600 184.600 57.000 ;
        RECT 183.900 56.100 184.200 56.600 ;
        RECT 179.900 55.700 182.300 55.900 ;
        RECT 177.400 55.600 182.300 55.700 ;
        RECT 183.000 55.800 184.200 56.100 ;
        RECT 177.400 55.500 180.300 55.600 ;
        RECT 177.400 55.400 180.200 55.500 ;
        RECT 173.400 55.100 173.800 55.200 ;
        RECT 180.600 55.100 181.000 55.200 ;
        RECT 182.200 55.100 182.600 55.200 ;
        RECT 173.400 54.800 175.900 55.100 ;
        RECT 175.500 54.700 175.900 54.800 ;
        RECT 178.500 54.800 182.600 55.100 ;
        RECT 178.500 54.700 178.900 54.800 ;
        RECT 174.700 54.200 175.100 54.300 ;
        RECT 179.300 54.200 179.700 54.300 ;
        RECT 183.000 54.200 183.300 55.800 ;
        RECT 186.200 55.600 186.600 59.900 ;
        RECT 187.000 55.900 187.400 59.900 ;
        RECT 187.800 56.200 188.200 59.900 ;
        RECT 189.400 56.200 189.800 59.900 ;
        RECT 187.800 55.900 189.800 56.200 ;
        RECT 190.500 56.300 190.900 59.900 ;
        RECT 194.500 59.200 194.900 59.900 ;
        RECT 194.500 58.800 195.400 59.200 ;
        RECT 194.500 56.400 194.900 58.800 ;
        RECT 196.600 57.500 197.000 59.500 ;
        RECT 190.500 55.900 191.400 56.300 ;
        RECT 194.100 56.100 194.900 56.400 ;
        RECT 184.500 55.300 186.600 55.600 ;
        RECT 184.500 55.200 184.900 55.300 ;
        RECT 185.300 54.900 185.700 55.000 ;
        RECT 183.800 54.600 185.700 54.900 ;
        RECT 183.800 54.500 184.200 54.600 ;
        RECT 171.100 53.900 176.600 54.200 ;
        RECT 171.300 53.800 171.700 53.900 ;
        RECT 174.200 53.800 174.600 53.900 ;
        RECT 175.800 53.800 176.600 53.900 ;
        RECT 177.800 53.900 183.300 54.200 ;
        RECT 177.800 53.800 178.600 53.900 ;
        RECT 167.800 53.300 169.700 53.600 ;
        RECT 167.800 51.100 168.200 53.300 ;
        RECT 169.300 53.200 169.700 53.300 ;
        RECT 174.200 52.800 174.500 53.800 ;
        RECT 173.300 52.700 173.700 52.800 ;
        RECT 170.200 52.100 170.600 52.500 ;
        RECT 172.300 52.400 173.700 52.700 ;
        RECT 174.200 52.400 174.600 52.800 ;
        RECT 172.300 52.100 172.600 52.400 ;
        RECT 175.000 52.100 175.400 52.500 ;
        RECT 169.900 51.800 170.600 52.100 ;
        RECT 169.900 51.100 170.500 51.800 ;
        RECT 172.200 51.100 172.600 52.100 ;
        RECT 174.400 51.800 175.400 52.100 ;
        RECT 174.400 51.100 174.800 51.800 ;
        RECT 176.600 51.100 177.000 53.500 ;
        RECT 177.400 51.100 177.800 53.500 ;
        RECT 179.900 52.800 180.200 53.900 ;
        RECT 180.600 53.800 181.000 53.900 ;
        RECT 182.700 53.800 183.100 53.900 ;
        RECT 186.200 53.600 186.600 55.300 ;
        RECT 187.100 55.200 187.400 55.900 ;
        RECT 189.000 55.200 189.400 55.400 ;
        RECT 187.000 54.900 188.200 55.200 ;
        RECT 189.000 54.900 189.800 55.200 ;
        RECT 187.000 54.800 187.400 54.900 ;
        RECT 184.700 53.300 186.600 53.600 ;
        RECT 184.700 53.200 185.100 53.300 ;
        RECT 179.000 52.100 179.400 52.500 ;
        RECT 179.800 52.400 180.200 52.800 ;
        RECT 180.700 52.700 181.100 52.800 ;
        RECT 180.700 52.400 182.100 52.700 ;
        RECT 181.800 52.100 182.100 52.400 ;
        RECT 183.800 52.100 184.200 52.500 ;
        RECT 179.000 51.800 180.000 52.100 ;
        RECT 179.600 51.100 180.000 51.800 ;
        RECT 181.800 51.100 182.200 52.100 ;
        RECT 183.800 51.800 184.500 52.100 ;
        RECT 183.900 51.100 184.500 51.800 ;
        RECT 186.200 51.100 186.600 53.300 ;
        RECT 187.000 52.800 187.400 53.200 ;
        RECT 187.900 53.100 188.200 54.900 ;
        RECT 189.400 54.800 189.800 54.900 ;
        RECT 190.200 54.800 190.600 55.600 ;
        RECT 188.600 54.100 189.000 54.600 ;
        RECT 190.200 54.100 190.500 54.800 ;
        RECT 188.600 53.800 190.500 54.100 ;
        RECT 191.000 54.200 191.300 55.900 ;
        RECT 191.800 55.100 192.200 55.200 ;
        RECT 193.400 55.100 193.800 55.600 ;
        RECT 191.800 54.800 193.800 55.100 ;
        RECT 194.100 54.200 194.400 56.100 ;
        RECT 196.700 55.800 197.000 57.500 ;
        RECT 198.700 56.300 199.100 59.900 ;
        RECT 198.200 55.900 199.100 56.300 ;
        RECT 199.800 55.900 200.200 59.900 ;
        RECT 200.600 56.200 201.000 59.900 ;
        RECT 202.200 56.200 202.600 59.900 ;
        RECT 200.600 55.900 202.600 56.200 ;
        RECT 204.600 56.200 205.000 59.900 ;
        RECT 206.200 56.400 206.600 59.900 ;
        RECT 204.600 55.900 205.900 56.200 ;
        RECT 206.200 55.900 206.700 56.400 ;
        RECT 195.100 55.500 197.000 55.800 ;
        RECT 195.100 54.500 195.400 55.500 ;
        RECT 191.000 53.800 191.400 54.200 ;
        RECT 193.400 53.800 194.400 54.200 ;
        RECT 194.700 54.100 195.400 54.500 ;
        RECT 195.800 54.400 196.200 55.200 ;
        RECT 196.600 54.400 197.000 55.200 ;
        RECT 198.300 54.200 198.600 55.900 ;
        RECT 199.000 54.800 199.400 55.600 ;
        RECT 199.900 55.200 200.200 55.900 ;
        RECT 201.800 55.200 202.200 55.400 ;
        RECT 199.800 54.900 201.000 55.200 ;
        RECT 201.800 55.100 202.600 55.200 ;
        RECT 203.000 55.100 203.400 55.200 ;
        RECT 201.800 54.900 203.400 55.100 ;
        RECT 199.800 54.800 200.200 54.900 ;
        RECT 187.100 52.400 187.500 52.800 ;
        RECT 187.800 51.100 188.200 53.100 ;
        RECT 191.000 52.100 191.300 53.800 ;
        RECT 194.100 53.500 194.400 53.800 ;
        RECT 194.900 53.900 195.400 54.100 ;
        RECT 194.900 53.600 197.000 53.900 ;
        RECT 198.200 53.800 198.600 54.200 ;
        RECT 194.100 53.300 194.500 53.500 ;
        RECT 191.800 52.400 192.200 53.200 ;
        RECT 194.100 53.000 194.900 53.300 ;
        RECT 191.000 51.100 191.400 52.100 ;
        RECT 194.500 51.500 194.900 53.000 ;
        RECT 196.700 52.500 197.000 53.600 ;
        RECT 196.600 51.500 197.000 52.500 ;
        RECT 197.400 52.400 197.800 53.200 ;
        RECT 198.300 53.100 198.600 53.800 ;
        RECT 199.800 53.100 200.200 53.200 ;
        RECT 200.700 53.100 201.000 54.900 ;
        RECT 202.200 54.800 203.400 54.900 ;
        RECT 205.600 54.900 205.900 55.900 ;
        RECT 201.400 53.800 201.800 54.600 ;
        RECT 205.600 54.500 206.100 54.900 ;
        RECT 205.600 53.700 205.900 54.500 ;
        RECT 206.400 54.200 206.700 55.900 ;
        RECT 208.600 55.600 209.000 59.900 ;
        RECT 210.200 55.600 210.600 59.900 ;
        RECT 211.800 55.600 212.200 59.900 ;
        RECT 213.400 55.600 213.800 59.900 ;
        RECT 215.000 55.600 215.400 59.900 ;
        RECT 217.100 57.900 217.700 59.900 ;
        RECT 219.400 57.900 219.800 59.900 ;
        RECT 221.600 58.200 222.000 59.900 ;
        RECT 221.600 57.900 222.600 58.200 ;
        RECT 217.400 57.500 217.800 57.900 ;
        RECT 219.500 57.600 219.800 57.900 ;
        RECT 219.100 57.300 220.900 57.600 ;
        RECT 222.200 57.500 222.600 57.900 ;
        RECT 219.100 57.200 219.500 57.300 ;
        RECT 220.500 57.200 220.900 57.300 ;
        RECT 217.000 56.600 217.700 57.000 ;
        RECT 217.400 56.100 217.700 56.600 ;
        RECT 218.500 56.500 219.600 56.800 ;
        RECT 218.500 56.400 218.900 56.500 ;
        RECT 217.400 55.800 218.600 56.100 ;
        RECT 208.600 55.200 209.500 55.600 ;
        RECT 210.200 55.200 211.300 55.600 ;
        RECT 211.800 55.200 212.900 55.600 ;
        RECT 213.400 55.200 214.600 55.600 ;
        RECT 209.100 54.500 209.500 55.200 ;
        RECT 210.900 54.500 211.300 55.200 ;
        RECT 212.500 54.500 212.900 55.200 ;
        RECT 206.200 53.800 206.700 54.200 ;
        RECT 207.800 54.100 208.700 54.500 ;
        RECT 209.100 54.100 210.400 54.500 ;
        RECT 210.900 54.100 212.100 54.500 ;
        RECT 212.500 54.100 213.800 54.500 ;
        RECT 207.800 53.800 208.200 54.100 ;
        RECT 209.100 53.800 209.500 54.100 ;
        RECT 210.900 53.800 211.300 54.100 ;
        RECT 212.500 53.800 212.900 54.100 ;
        RECT 214.200 53.800 214.600 55.200 ;
        RECT 198.200 52.800 200.200 53.100 ;
        RECT 198.300 52.100 198.600 52.800 ;
        RECT 199.900 52.400 200.300 52.800 ;
        RECT 198.200 51.100 198.600 52.100 ;
        RECT 200.600 51.100 201.000 53.100 ;
        RECT 204.600 53.400 205.900 53.700 ;
        RECT 204.600 51.100 205.000 53.400 ;
        RECT 206.400 53.100 206.700 53.800 ;
        RECT 206.200 52.800 206.700 53.100 ;
        RECT 208.600 53.400 209.500 53.800 ;
        RECT 210.200 53.400 211.300 53.800 ;
        RECT 211.800 53.400 212.900 53.800 ;
        RECT 213.400 53.400 214.600 53.800 ;
        RECT 215.000 55.300 217.100 55.600 ;
        RECT 215.000 53.600 215.400 55.300 ;
        RECT 216.700 55.200 217.100 55.300 ;
        RECT 218.300 55.200 218.600 55.800 ;
        RECT 219.300 55.900 219.600 56.500 ;
        RECT 219.900 56.500 220.300 56.600 ;
        RECT 222.200 56.500 222.600 56.600 ;
        RECT 219.900 56.200 222.600 56.500 ;
        RECT 219.300 55.700 221.700 55.900 ;
        RECT 223.800 55.700 224.200 59.900 ;
        RECT 224.600 55.900 225.000 59.900 ;
        RECT 225.400 56.200 225.800 59.900 ;
        RECT 227.000 56.200 227.400 59.900 ;
        RECT 225.400 55.900 227.400 56.200 ;
        RECT 219.300 55.600 224.200 55.700 ;
        RECT 221.300 55.500 224.200 55.600 ;
        RECT 221.400 55.400 224.200 55.500 ;
        RECT 224.700 55.200 225.000 55.900 ;
        RECT 227.800 55.600 228.200 59.900 ;
        RECT 229.900 57.900 230.500 59.900 ;
        RECT 232.200 57.900 232.600 59.900 ;
        RECT 234.400 58.200 234.800 59.900 ;
        RECT 234.400 57.900 235.400 58.200 ;
        RECT 230.200 57.500 230.600 57.900 ;
        RECT 232.300 57.600 232.600 57.900 ;
        RECT 231.900 57.300 233.700 57.600 ;
        RECT 235.000 57.500 235.400 57.900 ;
        RECT 231.900 57.200 232.300 57.300 ;
        RECT 233.300 57.200 233.700 57.300 ;
        RECT 229.800 56.600 230.500 57.000 ;
        RECT 230.200 56.100 230.500 56.600 ;
        RECT 231.300 56.500 232.400 56.800 ;
        RECT 231.300 56.400 231.700 56.500 ;
        RECT 230.200 55.800 231.400 56.100 ;
        RECT 226.600 55.200 227.000 55.400 ;
        RECT 227.800 55.300 229.900 55.600 ;
        RECT 215.900 54.900 216.300 55.000 ;
        RECT 215.900 54.600 217.800 54.900 ;
        RECT 218.200 54.800 218.600 55.200 ;
        RECT 220.600 55.100 221.000 55.200 ;
        RECT 220.600 54.800 223.100 55.100 ;
        RECT 224.600 54.900 225.800 55.200 ;
        RECT 226.600 54.900 227.400 55.200 ;
        RECT 224.600 54.800 225.000 54.900 ;
        RECT 217.400 54.500 217.800 54.600 ;
        RECT 218.300 54.200 218.600 54.800 ;
        RECT 221.400 54.700 221.800 54.800 ;
        RECT 222.700 54.700 223.100 54.800 ;
        RECT 221.900 54.200 222.300 54.300 ;
        RECT 218.300 53.900 223.800 54.200 ;
        RECT 218.500 53.800 218.900 53.900 ;
        RECT 206.200 51.100 206.600 52.800 ;
        RECT 208.600 51.100 209.000 53.400 ;
        RECT 210.200 51.100 210.600 53.400 ;
        RECT 211.800 51.100 212.200 53.400 ;
        RECT 213.400 51.100 213.800 53.400 ;
        RECT 215.000 53.300 216.900 53.600 ;
        RECT 215.000 51.100 215.400 53.300 ;
        RECT 216.500 53.200 216.900 53.300 ;
        RECT 221.400 52.800 221.700 53.900 ;
        RECT 223.000 53.800 223.800 53.900 ;
        RECT 224.600 54.100 225.000 54.200 ;
        RECT 225.500 54.100 225.800 54.900 ;
        RECT 227.000 54.800 227.400 54.900 ;
        RECT 224.600 53.800 225.800 54.100 ;
        RECT 226.200 53.800 226.600 54.600 ;
        RECT 220.500 52.700 220.900 52.800 ;
        RECT 217.400 52.100 217.800 52.500 ;
        RECT 219.500 52.400 220.900 52.700 ;
        RECT 221.400 52.400 221.800 52.800 ;
        RECT 219.500 52.100 219.800 52.400 ;
        RECT 222.200 52.100 222.600 52.500 ;
        RECT 217.100 51.800 217.800 52.100 ;
        RECT 217.100 51.100 217.700 51.800 ;
        RECT 219.400 51.100 219.800 52.100 ;
        RECT 221.600 51.800 222.600 52.100 ;
        RECT 221.600 51.100 222.000 51.800 ;
        RECT 223.800 51.100 224.200 53.500 ;
        RECT 224.600 52.800 225.000 53.200 ;
        RECT 225.500 53.100 225.800 53.800 ;
        RECT 224.700 52.400 225.100 52.800 ;
        RECT 225.400 51.100 225.800 53.100 ;
        RECT 227.800 53.600 228.200 55.300 ;
        RECT 229.500 55.200 229.900 55.300 ;
        RECT 231.100 55.200 231.400 55.800 ;
        RECT 232.100 55.900 232.400 56.500 ;
        RECT 232.700 56.500 233.100 56.600 ;
        RECT 235.000 56.500 235.400 56.600 ;
        RECT 232.700 56.200 235.400 56.500 ;
        RECT 232.100 55.700 234.500 55.900 ;
        RECT 236.600 55.700 237.000 59.900 ;
        RECT 237.800 56.800 238.200 57.200 ;
        RECT 237.800 56.200 238.100 56.800 ;
        RECT 238.500 56.200 238.900 59.900 ;
        RECT 237.400 55.900 238.100 56.200 ;
        RECT 238.400 55.900 238.900 56.200 ;
        RECT 237.400 55.800 237.800 55.900 ;
        RECT 232.100 55.600 237.000 55.700 ;
        RECT 234.100 55.500 237.000 55.600 ;
        RECT 234.200 55.400 237.000 55.500 ;
        RECT 238.400 55.200 238.700 55.900 ;
        RECT 240.600 55.600 241.000 59.900 ;
        RECT 242.700 57.900 243.300 59.900 ;
        RECT 245.000 57.900 245.400 59.900 ;
        RECT 247.200 58.200 247.600 59.900 ;
        RECT 247.200 57.900 248.200 58.200 ;
        RECT 243.000 57.500 243.400 57.900 ;
        RECT 245.100 57.600 245.400 57.900 ;
        RECT 244.700 57.300 246.500 57.600 ;
        RECT 247.800 57.500 248.200 57.900 ;
        RECT 244.700 57.200 245.100 57.300 ;
        RECT 246.100 57.200 246.500 57.300 ;
        RECT 242.600 56.600 243.300 57.000 ;
        RECT 243.000 56.100 243.300 56.600 ;
        RECT 244.100 56.500 245.200 56.800 ;
        RECT 244.100 56.400 244.500 56.500 ;
        RECT 243.000 55.800 244.200 56.100 ;
        RECT 240.600 55.300 242.700 55.600 ;
        RECT 228.700 54.900 229.100 55.000 ;
        RECT 228.700 54.600 230.600 54.900 ;
        RECT 231.000 54.800 231.400 55.200 ;
        RECT 233.400 55.100 233.800 55.200 ;
        RECT 233.400 54.800 235.900 55.100 ;
        RECT 238.200 54.800 238.700 55.200 ;
        RECT 230.200 54.500 230.600 54.600 ;
        RECT 231.100 54.200 231.400 54.800 ;
        RECT 234.200 54.700 234.600 54.800 ;
        RECT 235.500 54.700 235.900 54.800 ;
        RECT 234.700 54.200 235.100 54.300 ;
        RECT 238.400 54.200 238.700 54.800 ;
        RECT 239.000 54.400 239.400 55.200 ;
        RECT 231.100 53.900 236.600 54.200 ;
        RECT 231.300 53.800 231.700 53.900 ;
        RECT 227.800 53.300 229.700 53.600 ;
        RECT 227.800 51.100 228.200 53.300 ;
        RECT 229.300 53.200 229.700 53.300 ;
        RECT 234.200 52.800 234.500 53.900 ;
        RECT 235.800 53.800 236.600 53.900 ;
        RECT 237.400 53.800 238.700 54.200 ;
        RECT 239.800 54.100 240.200 54.200 ;
        RECT 239.400 53.800 240.200 54.100 ;
        RECT 233.300 52.700 233.700 52.800 ;
        RECT 230.200 52.100 230.600 52.500 ;
        RECT 232.300 52.400 233.700 52.700 ;
        RECT 234.200 52.400 234.600 52.800 ;
        RECT 232.300 52.100 232.600 52.400 ;
        RECT 235.000 52.100 235.400 52.500 ;
        RECT 229.900 51.800 230.600 52.100 ;
        RECT 229.900 51.100 230.500 51.800 ;
        RECT 232.200 51.100 232.600 52.100 ;
        RECT 234.400 51.800 235.400 52.100 ;
        RECT 234.400 51.100 234.800 51.800 ;
        RECT 236.600 51.100 237.000 53.500 ;
        RECT 237.500 53.100 237.800 53.800 ;
        RECT 239.400 53.600 239.800 53.800 ;
        RECT 240.600 53.600 241.000 55.300 ;
        RECT 242.300 55.200 242.700 55.300 ;
        RECT 241.500 54.900 241.900 55.000 ;
        RECT 241.500 54.600 243.400 54.900 ;
        RECT 243.000 54.500 243.400 54.600 ;
        RECT 243.900 54.200 244.200 55.800 ;
        RECT 244.900 55.900 245.200 56.500 ;
        RECT 245.500 56.500 245.900 56.600 ;
        RECT 247.800 56.500 248.200 56.600 ;
        RECT 245.500 56.200 248.200 56.500 ;
        RECT 244.900 55.700 247.300 55.900 ;
        RECT 249.400 55.700 249.800 59.900 ;
        RECT 244.900 55.600 249.800 55.700 ;
        RECT 246.900 55.500 249.800 55.600 ;
        RECT 247.000 55.400 249.800 55.500 ;
        RECT 246.200 55.100 246.600 55.200 ;
        RECT 246.200 54.800 248.700 55.100 ;
        RECT 247.000 54.700 247.400 54.800 ;
        RECT 248.300 54.700 248.700 54.800 ;
        RECT 247.500 54.200 247.900 54.300 ;
        RECT 243.900 53.900 249.400 54.200 ;
        RECT 244.100 53.800 244.500 53.900 ;
        RECT 246.200 53.800 246.600 53.900 ;
        RECT 240.600 53.300 242.500 53.600 ;
        RECT 238.300 53.100 240.100 53.300 ;
        RECT 237.400 51.100 237.800 53.100 ;
        RECT 238.200 53.000 240.200 53.100 ;
        RECT 238.200 51.100 238.600 53.000 ;
        RECT 239.800 51.100 240.200 53.000 ;
        RECT 240.600 51.100 241.000 53.300 ;
        RECT 242.100 53.200 242.500 53.300 ;
        RECT 247.000 52.800 247.300 53.900 ;
        RECT 248.600 53.800 249.400 53.900 ;
        RECT 246.100 52.700 246.500 52.800 ;
        RECT 243.000 52.100 243.400 52.500 ;
        RECT 245.100 52.400 246.500 52.700 ;
        RECT 247.000 52.400 247.400 52.800 ;
        RECT 245.100 52.100 245.400 52.400 ;
        RECT 247.800 52.100 248.200 52.500 ;
        RECT 242.700 51.800 243.400 52.100 ;
        RECT 242.700 51.100 243.300 51.800 ;
        RECT 245.000 51.100 245.400 52.100 ;
        RECT 247.200 51.800 248.200 52.100 ;
        RECT 247.200 51.100 247.600 51.800 ;
        RECT 249.400 51.100 249.800 53.500 ;
        RECT 2.200 47.600 2.600 49.900 ;
        RECT 3.800 47.600 4.200 49.900 ;
        RECT 5.400 47.600 5.800 49.900 ;
        RECT 7.000 47.600 7.400 49.900 ;
        RECT 8.600 47.600 9.000 49.900 ;
        RECT 11.500 48.200 11.900 49.900 ;
        RECT 11.000 47.900 11.900 48.200 ;
        RECT 12.600 47.900 13.000 49.900 ;
        RECT 13.400 48.000 13.800 49.900 ;
        RECT 15.000 48.000 15.400 49.900 ;
        RECT 13.400 47.900 15.400 48.000 ;
        RECT 1.500 47.300 2.600 47.600 ;
        RECT 1.500 45.800 1.800 47.300 ;
        RECT 3.000 47.200 4.200 47.600 ;
        RECT 4.700 47.200 5.800 47.600 ;
        RECT 6.300 47.200 7.400 47.600 ;
        RECT 8.100 47.200 9.000 47.600 ;
        RECT 2.200 45.800 2.600 46.600 ;
        RECT 3.000 45.800 3.400 47.200 ;
        RECT 4.700 46.900 5.100 47.200 ;
        RECT 6.300 46.900 6.700 47.200 ;
        RECT 8.100 46.900 8.500 47.200 ;
        RECT 9.400 46.900 9.800 47.200 ;
        RECT 3.800 46.500 5.100 46.900 ;
        RECT 5.500 46.500 6.700 46.900 ;
        RECT 7.200 46.500 8.500 46.900 ;
        RECT 8.900 46.500 9.800 46.900 ;
        RECT 10.200 46.800 10.600 47.600 ;
        RECT 4.700 45.800 5.100 46.500 ;
        RECT 6.300 45.800 6.700 46.500 ;
        RECT 8.100 45.800 8.500 46.500 ;
        RECT 11.000 46.100 11.400 47.900 ;
        RECT 12.700 47.200 13.000 47.900 ;
        RECT 13.500 47.700 15.300 47.900 ;
        RECT 15.800 47.500 16.200 49.900 ;
        RECT 18.000 49.200 18.400 49.900 ;
        RECT 17.400 48.900 18.400 49.200 ;
        RECT 20.200 48.900 20.600 49.900 ;
        RECT 22.300 49.200 22.900 49.900 ;
        RECT 22.200 48.900 22.900 49.200 ;
        RECT 17.400 48.500 17.800 48.900 ;
        RECT 20.200 48.600 20.500 48.900 ;
        RECT 18.200 48.200 18.600 48.600 ;
        RECT 19.100 48.300 20.500 48.600 ;
        RECT 22.200 48.500 22.600 48.900 ;
        RECT 19.100 48.200 19.500 48.300 ;
        RECT 14.600 47.200 15.000 47.400 ;
        RECT 12.600 46.800 13.900 47.200 ;
        RECT 14.600 46.900 15.400 47.200 ;
        RECT 15.000 46.800 15.400 46.900 ;
        RECT 16.200 47.100 17.000 47.200 ;
        RECT 18.300 47.100 18.600 48.200 ;
        RECT 23.100 47.700 23.500 47.800 ;
        RECT 24.600 47.700 25.000 49.900 ;
        RECT 27.300 49.200 27.700 49.500 ;
        RECT 27.300 48.800 28.200 49.200 ;
        RECT 27.300 48.000 27.700 48.800 ;
        RECT 29.400 48.500 29.800 49.500 ;
        RECT 23.100 47.400 25.000 47.700 ;
        RECT 21.100 47.100 21.500 47.200 ;
        RECT 16.200 46.800 21.700 47.100 ;
        RECT 11.000 45.800 12.900 46.100 ;
        RECT 1.200 45.400 1.800 45.800 ;
        RECT 3.000 45.400 4.200 45.800 ;
        RECT 4.700 45.400 5.800 45.800 ;
        RECT 6.300 45.400 7.400 45.800 ;
        RECT 8.100 45.400 9.000 45.800 ;
        RECT 1.500 45.100 1.800 45.400 ;
        RECT 1.500 44.800 2.600 45.100 ;
        RECT 2.200 41.100 2.600 44.800 ;
        RECT 3.800 41.100 4.200 45.400 ;
        RECT 5.400 41.100 5.800 45.400 ;
        RECT 7.000 41.100 7.400 45.400 ;
        RECT 8.600 41.100 9.000 45.400 ;
        RECT 11.000 41.100 11.400 45.800 ;
        RECT 12.600 45.200 12.900 45.800 ;
        RECT 13.600 45.200 13.900 46.800 ;
        RECT 17.700 46.700 18.100 46.800 ;
        RECT 14.200 45.800 14.600 46.600 ;
        RECT 16.900 46.200 17.300 46.300 ;
        RECT 18.200 46.200 18.600 46.300 ;
        RECT 16.900 45.900 19.400 46.200 ;
        RECT 19.000 45.800 19.400 45.900 ;
        RECT 15.800 45.500 18.600 45.600 ;
        RECT 15.800 45.400 18.700 45.500 ;
        RECT 15.800 45.300 20.700 45.400 ;
        RECT 11.800 44.400 12.200 45.200 ;
        RECT 12.600 45.100 13.000 45.200 ;
        RECT 12.600 44.800 13.300 45.100 ;
        RECT 13.600 44.800 14.600 45.200 ;
        RECT 13.000 44.200 13.300 44.800 ;
        RECT 13.000 43.800 13.400 44.200 ;
        RECT 13.700 41.100 14.100 44.800 ;
        RECT 15.800 41.100 16.200 45.300 ;
        RECT 18.300 45.100 20.700 45.300 ;
        RECT 17.400 44.500 20.100 44.800 ;
        RECT 17.400 44.400 17.800 44.500 ;
        RECT 19.700 44.400 20.100 44.500 ;
        RECT 20.400 44.500 20.700 45.100 ;
        RECT 21.400 45.200 21.700 46.800 ;
        RECT 22.200 46.400 22.600 46.500 ;
        RECT 22.200 46.100 24.100 46.400 ;
        RECT 23.700 46.000 24.100 46.100 ;
        RECT 22.900 45.700 23.300 45.800 ;
        RECT 24.600 45.700 25.000 47.400 ;
        RECT 26.900 47.700 27.700 48.000 ;
        RECT 26.900 47.500 27.300 47.700 ;
        RECT 26.900 47.200 27.200 47.500 ;
        RECT 29.500 47.400 29.800 48.500 ;
        RECT 31.500 48.200 31.900 49.900 ;
        RECT 31.000 47.900 31.900 48.200 ;
        RECT 32.600 47.900 33.000 49.900 ;
        RECT 33.400 48.000 33.800 49.900 ;
        RECT 35.000 48.000 35.400 49.900 ;
        RECT 33.400 47.900 35.400 48.000 ;
        RECT 26.200 46.800 27.200 47.200 ;
        RECT 27.700 47.100 29.800 47.400 ;
        RECT 27.700 46.900 28.200 47.100 ;
        RECT 25.400 46.100 25.800 46.200 ;
        RECT 26.200 46.100 26.600 46.200 ;
        RECT 25.400 45.800 26.600 46.100 ;
        RECT 22.900 45.400 25.000 45.700 ;
        RECT 26.200 45.400 26.600 45.800 ;
        RECT 21.400 44.900 22.600 45.200 ;
        RECT 21.100 44.500 21.500 44.600 ;
        RECT 20.400 44.200 21.500 44.500 ;
        RECT 22.300 44.400 22.600 44.900 ;
        RECT 22.300 44.000 23.000 44.400 ;
        RECT 19.100 43.700 19.500 43.800 ;
        RECT 20.500 43.700 20.900 43.800 ;
        RECT 17.400 43.100 17.800 43.500 ;
        RECT 19.100 43.400 20.900 43.700 ;
        RECT 20.200 43.100 20.500 43.400 ;
        RECT 22.200 43.100 22.600 43.500 ;
        RECT 17.400 42.800 18.400 43.100 ;
        RECT 18.000 41.100 18.400 42.800 ;
        RECT 20.200 41.100 20.600 43.100 ;
        RECT 22.300 41.100 22.900 43.100 ;
        RECT 24.600 41.100 25.000 45.400 ;
        RECT 26.900 44.900 27.200 46.800 ;
        RECT 27.500 46.500 28.200 46.900 ;
        RECT 30.200 46.800 30.600 47.600 ;
        RECT 27.900 45.500 28.200 46.500 ;
        RECT 28.600 45.800 29.000 46.600 ;
        RECT 29.400 45.800 29.800 46.600 ;
        RECT 31.000 46.100 31.400 47.900 ;
        RECT 32.700 47.200 33.000 47.900 ;
        RECT 33.500 47.700 35.300 47.900 ;
        RECT 35.800 47.700 36.200 49.900 ;
        RECT 37.900 49.200 38.500 49.900 ;
        RECT 37.900 48.900 38.600 49.200 ;
        RECT 40.200 48.900 40.600 49.900 ;
        RECT 42.400 49.200 42.800 49.900 ;
        RECT 42.400 48.900 43.400 49.200 ;
        RECT 38.200 48.500 38.600 48.900 ;
        RECT 40.300 48.600 40.600 48.900 ;
        RECT 40.300 48.300 41.700 48.600 ;
        RECT 41.300 48.200 41.700 48.300 ;
        RECT 42.200 48.200 42.600 48.600 ;
        RECT 43.000 48.500 43.400 48.900 ;
        RECT 37.300 47.700 37.700 47.800 ;
        RECT 35.800 47.400 37.700 47.700 ;
        RECT 34.600 47.200 35.000 47.400 ;
        RECT 32.600 46.800 33.900 47.200 ;
        RECT 34.600 46.900 35.400 47.200 ;
        RECT 35.000 46.800 35.400 46.900 ;
        RECT 31.000 45.800 32.900 46.100 ;
        RECT 27.900 45.200 29.800 45.500 ;
        RECT 26.900 44.600 27.700 44.900 ;
        RECT 27.300 41.100 27.700 44.600 ;
        RECT 29.500 43.500 29.800 45.200 ;
        RECT 29.400 41.500 29.800 43.500 ;
        RECT 31.000 41.100 31.400 45.800 ;
        RECT 32.600 45.200 32.900 45.800 ;
        RECT 31.800 44.400 32.200 45.200 ;
        RECT 32.600 45.100 33.000 45.200 ;
        RECT 33.600 45.100 33.900 46.800 ;
        RECT 34.200 45.800 34.600 46.600 ;
        RECT 35.800 45.700 36.200 47.400 ;
        RECT 39.300 47.100 39.700 47.200 ;
        RECT 42.200 47.100 42.500 48.200 ;
        RECT 44.600 47.500 45.000 49.900 ;
        RECT 45.700 49.200 46.100 49.900 ;
        RECT 50.700 49.200 51.100 49.900 ;
        RECT 45.700 48.800 46.600 49.200 ;
        RECT 50.700 48.800 51.400 49.200 ;
        RECT 45.700 48.200 46.100 48.800 ;
        RECT 50.700 48.200 51.100 48.800 ;
        RECT 45.700 47.900 46.600 48.200 ;
        RECT 43.800 47.100 44.600 47.200 ;
        RECT 45.400 47.100 45.800 47.200 ;
        RECT 39.100 46.800 45.800 47.100 ;
        RECT 38.200 46.400 38.600 46.500 ;
        RECT 36.700 46.100 38.600 46.400 ;
        RECT 39.100 46.200 39.400 46.800 ;
        RECT 42.700 46.700 43.100 46.800 ;
        RECT 42.200 46.200 42.600 46.300 ;
        RECT 43.500 46.200 43.900 46.300 ;
        RECT 36.700 46.000 37.100 46.100 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 41.400 45.900 43.900 46.200 ;
        RECT 41.400 45.800 41.800 45.900 ;
        RECT 37.500 45.700 37.900 45.800 ;
        RECT 35.800 45.400 37.900 45.700 ;
        RECT 32.600 44.800 33.300 45.100 ;
        RECT 33.600 44.800 34.100 45.100 ;
        RECT 33.000 44.200 33.300 44.800 ;
        RECT 33.000 43.800 33.400 44.200 ;
        RECT 33.700 41.100 34.100 44.800 ;
        RECT 35.800 41.100 36.200 45.400 ;
        RECT 39.100 45.200 39.400 45.800 ;
        RECT 42.200 45.500 45.000 45.600 ;
        RECT 42.100 45.400 45.000 45.500 ;
        RECT 38.200 44.900 39.400 45.200 ;
        RECT 40.100 45.300 45.000 45.400 ;
        RECT 40.100 45.100 42.500 45.300 ;
        RECT 38.200 44.400 38.500 44.900 ;
        RECT 37.800 44.000 38.500 44.400 ;
        RECT 39.300 44.500 39.700 44.600 ;
        RECT 40.100 44.500 40.400 45.100 ;
        RECT 39.300 44.200 40.400 44.500 ;
        RECT 40.700 44.500 43.400 44.800 ;
        RECT 40.700 44.400 41.100 44.500 ;
        RECT 43.000 44.400 43.400 44.500 ;
        RECT 39.900 43.700 40.300 43.800 ;
        RECT 41.300 43.700 41.700 43.800 ;
        RECT 38.200 43.100 38.600 43.500 ;
        RECT 39.900 43.400 41.700 43.700 ;
        RECT 40.300 43.100 40.600 43.400 ;
        RECT 43.000 43.100 43.400 43.500 ;
        RECT 37.900 41.100 38.500 43.100 ;
        RECT 40.200 41.100 40.600 43.100 ;
        RECT 42.400 42.800 43.400 43.100 ;
        RECT 42.400 41.100 42.800 42.800 ;
        RECT 44.600 41.100 45.000 45.300 ;
        RECT 45.400 43.800 45.800 45.200 ;
        RECT 46.200 41.100 46.600 47.900 ;
        RECT 50.200 47.900 51.100 48.200 ;
        RECT 50.200 41.100 50.600 47.900 ;
        RECT 51.800 47.700 52.200 49.900 ;
        RECT 53.900 49.200 54.500 49.900 ;
        RECT 53.900 48.900 54.600 49.200 ;
        RECT 56.200 48.900 56.600 49.900 ;
        RECT 58.400 49.200 58.800 49.900 ;
        RECT 58.400 48.900 59.400 49.200 ;
        RECT 54.200 48.500 54.600 48.900 ;
        RECT 56.300 48.600 56.600 48.900 ;
        RECT 56.300 48.300 57.700 48.600 ;
        RECT 57.300 48.200 57.700 48.300 ;
        RECT 58.200 48.200 58.600 48.600 ;
        RECT 59.000 48.500 59.400 48.900 ;
        RECT 53.300 47.700 53.700 47.800 ;
        RECT 51.800 47.400 53.700 47.700 ;
        RECT 51.800 45.700 52.200 47.400 ;
        RECT 55.300 47.100 55.700 47.200 ;
        RECT 58.200 47.100 58.500 48.200 ;
        RECT 60.600 47.500 61.000 49.900 ;
        RECT 61.400 47.500 61.800 49.900 ;
        RECT 63.600 49.200 64.000 49.900 ;
        RECT 63.000 48.900 64.000 49.200 ;
        RECT 65.800 48.900 66.200 49.900 ;
        RECT 67.900 49.200 68.500 49.900 ;
        RECT 67.800 48.900 68.500 49.200 ;
        RECT 63.000 48.500 63.400 48.900 ;
        RECT 65.800 48.600 66.100 48.900 ;
        RECT 63.800 48.200 64.200 48.600 ;
        RECT 64.700 48.300 66.100 48.600 ;
        RECT 67.800 48.500 68.200 48.900 ;
        RECT 64.700 48.200 65.100 48.300 ;
        RECT 59.800 47.100 60.600 47.200 ;
        RECT 55.100 46.800 60.600 47.100 ;
        RECT 61.800 47.100 62.600 47.200 ;
        RECT 63.900 47.100 64.200 48.200 ;
        RECT 68.700 47.700 69.100 47.800 ;
        RECT 70.200 47.700 70.600 49.900 ;
        RECT 71.000 48.000 71.400 49.900 ;
        RECT 72.600 48.000 73.000 49.900 ;
        RECT 71.000 47.900 73.000 48.000 ;
        RECT 73.400 47.900 73.800 49.900 ;
        RECT 74.500 48.200 74.900 49.900 ;
        RECT 74.500 47.900 75.400 48.200 ;
        RECT 71.100 47.700 72.900 47.900 ;
        RECT 68.700 47.400 70.600 47.700 ;
        RECT 66.700 47.100 67.100 47.200 ;
        RECT 61.800 46.800 67.300 47.100 ;
        RECT 54.200 46.400 54.600 46.500 ;
        RECT 52.700 46.100 54.600 46.400 ;
        RECT 52.700 46.000 53.100 46.100 ;
        RECT 53.500 45.700 53.900 45.800 ;
        RECT 51.800 45.400 53.900 45.700 ;
        RECT 51.000 44.100 51.400 45.200 ;
        RECT 51.800 44.100 52.200 45.400 ;
        RECT 55.100 45.200 55.400 46.800 ;
        RECT 58.700 46.700 59.100 46.800 ;
        RECT 63.300 46.700 63.700 46.800 ;
        RECT 58.200 46.200 58.600 46.300 ;
        RECT 59.500 46.200 59.900 46.300 ;
        RECT 57.400 45.900 59.900 46.200 ;
        RECT 62.500 46.200 62.900 46.300 ;
        RECT 62.500 45.900 65.000 46.200 ;
        RECT 57.400 45.800 57.800 45.900 ;
        RECT 64.600 45.800 65.000 45.900 ;
        RECT 58.200 45.500 61.000 45.600 ;
        RECT 58.100 45.400 61.000 45.500 ;
        RECT 54.200 44.900 55.400 45.200 ;
        RECT 56.100 45.300 61.000 45.400 ;
        RECT 56.100 45.100 58.500 45.300 ;
        RECT 54.200 44.400 54.500 44.900 ;
        RECT 51.000 43.800 52.200 44.100 ;
        RECT 53.800 44.000 54.500 44.400 ;
        RECT 55.300 44.500 55.700 44.600 ;
        RECT 56.100 44.500 56.400 45.100 ;
        RECT 55.300 44.200 56.400 44.500 ;
        RECT 56.700 44.500 59.400 44.800 ;
        RECT 56.700 44.400 57.100 44.500 ;
        RECT 59.000 44.400 59.400 44.500 ;
        RECT 51.800 41.100 52.200 43.800 ;
        RECT 55.900 43.700 56.300 43.800 ;
        RECT 57.300 43.700 57.700 43.800 ;
        RECT 54.200 43.100 54.600 43.500 ;
        RECT 55.900 43.400 57.700 43.700 ;
        RECT 56.300 43.100 56.600 43.400 ;
        RECT 59.000 43.100 59.400 43.500 ;
        RECT 53.900 41.100 54.500 43.100 ;
        RECT 56.200 41.100 56.600 43.100 ;
        RECT 58.400 42.800 59.400 43.100 ;
        RECT 58.400 41.100 58.800 42.800 ;
        RECT 60.600 41.100 61.000 45.300 ;
        RECT 61.400 45.500 64.200 45.600 ;
        RECT 61.400 45.400 64.300 45.500 ;
        RECT 61.400 45.300 66.300 45.400 ;
        RECT 61.400 41.100 61.800 45.300 ;
        RECT 63.900 45.100 66.300 45.300 ;
        RECT 63.000 44.500 65.700 44.800 ;
        RECT 63.000 44.400 63.400 44.500 ;
        RECT 65.300 44.400 65.700 44.500 ;
        RECT 66.000 44.500 66.300 45.100 ;
        RECT 67.000 45.200 67.300 46.800 ;
        RECT 67.800 46.400 68.200 46.500 ;
        RECT 67.800 46.100 69.700 46.400 ;
        RECT 69.300 46.000 69.700 46.100 ;
        RECT 68.500 45.700 68.900 45.800 ;
        RECT 70.200 45.700 70.600 47.400 ;
        RECT 71.400 47.200 71.800 47.400 ;
        RECT 73.400 47.200 73.700 47.900 ;
        RECT 71.000 46.900 71.800 47.200 ;
        RECT 71.000 46.800 71.400 46.900 ;
        RECT 72.500 46.800 73.800 47.200 ;
        RECT 71.800 45.800 72.200 46.600 ;
        RECT 68.500 45.400 70.600 45.700 ;
        RECT 67.000 44.900 68.200 45.200 ;
        RECT 66.700 44.500 67.100 44.600 ;
        RECT 66.000 44.200 67.100 44.500 ;
        RECT 67.900 44.400 68.200 44.900 ;
        RECT 67.900 44.000 68.600 44.400 ;
        RECT 64.700 43.700 65.100 43.800 ;
        RECT 66.100 43.700 66.500 43.800 ;
        RECT 63.000 43.100 63.400 43.500 ;
        RECT 64.700 43.400 66.500 43.700 ;
        RECT 65.800 43.100 66.100 43.400 ;
        RECT 67.800 43.100 68.200 43.500 ;
        RECT 63.000 42.800 64.000 43.100 ;
        RECT 63.600 41.100 64.000 42.800 ;
        RECT 65.800 41.100 66.200 43.100 ;
        RECT 67.900 41.100 68.500 43.100 ;
        RECT 70.200 41.100 70.600 45.400 ;
        RECT 72.500 45.100 72.800 46.800 ;
        RECT 75.000 46.100 75.400 47.900 ;
        RECT 75.800 46.800 76.200 47.600 ;
        RECT 76.600 47.500 77.000 49.900 ;
        RECT 78.800 49.200 79.200 49.900 ;
        RECT 78.200 48.900 79.200 49.200 ;
        RECT 81.000 48.900 81.400 49.900 ;
        RECT 83.100 49.200 83.700 49.900 ;
        RECT 83.000 48.900 83.700 49.200 ;
        RECT 78.200 48.500 78.600 48.900 ;
        RECT 81.000 48.600 81.300 48.900 ;
        RECT 79.000 48.200 79.400 48.600 ;
        RECT 79.900 48.300 81.300 48.600 ;
        RECT 83.000 48.500 83.400 48.900 ;
        RECT 79.900 48.200 80.300 48.300 ;
        RECT 77.000 47.100 77.800 47.200 ;
        RECT 79.100 47.100 79.400 48.200 ;
        RECT 83.900 47.700 84.300 47.800 ;
        RECT 85.400 47.700 85.800 49.900 ;
        RECT 87.500 48.200 87.900 49.900 ;
        RECT 83.900 47.400 85.800 47.700 ;
        RECT 87.000 47.900 87.900 48.200 ;
        RECT 88.600 47.900 89.000 49.900 ;
        RECT 89.400 48.000 89.800 49.900 ;
        RECT 91.000 48.000 91.400 49.900 ;
        RECT 89.400 47.900 91.400 48.000 ;
        RECT 81.900 47.100 82.300 47.200 ;
        RECT 85.400 47.100 85.800 47.400 ;
        RECT 86.200 47.100 86.600 47.600 ;
        RECT 77.000 46.800 82.500 47.100 ;
        RECT 78.500 46.700 78.900 46.800 ;
        RECT 73.400 45.800 75.400 46.100 ;
        RECT 77.700 46.200 78.100 46.300 ;
        RECT 77.700 45.900 80.200 46.200 ;
        RECT 79.800 45.800 80.200 45.900 ;
        RECT 73.400 45.200 73.700 45.800 ;
        RECT 73.400 45.100 73.800 45.200 ;
        RECT 72.300 44.800 72.800 45.100 ;
        RECT 73.100 44.800 73.800 45.100 ;
        RECT 72.300 41.100 72.700 44.800 ;
        RECT 73.100 44.200 73.400 44.800 ;
        RECT 74.200 44.400 74.600 45.200 ;
        RECT 73.000 43.800 73.400 44.200 ;
        RECT 75.000 41.100 75.400 45.800 ;
        RECT 76.600 45.500 79.400 45.600 ;
        RECT 76.600 45.400 79.500 45.500 ;
        RECT 76.600 45.300 81.500 45.400 ;
        RECT 76.600 41.100 77.000 45.300 ;
        RECT 79.100 45.100 81.500 45.300 ;
        RECT 78.200 44.500 80.900 44.800 ;
        RECT 78.200 44.400 78.600 44.500 ;
        RECT 80.500 44.400 80.900 44.500 ;
        RECT 81.200 44.500 81.500 45.100 ;
        RECT 82.200 45.200 82.500 46.800 ;
        RECT 85.400 46.800 86.600 47.100 ;
        RECT 83.000 46.400 83.400 46.500 ;
        RECT 83.000 46.100 84.900 46.400 ;
        RECT 84.500 46.000 84.900 46.100 ;
        RECT 83.700 45.700 84.100 45.800 ;
        RECT 85.400 45.700 85.800 46.800 ;
        RECT 83.700 45.400 85.800 45.700 ;
        RECT 82.200 44.900 83.400 45.200 ;
        RECT 81.900 44.500 82.300 44.600 ;
        RECT 81.200 44.200 82.300 44.500 ;
        RECT 83.100 44.400 83.400 44.900 ;
        RECT 83.100 44.000 83.800 44.400 ;
        RECT 79.900 43.700 80.300 43.800 ;
        RECT 81.300 43.700 81.700 43.800 ;
        RECT 78.200 43.100 78.600 43.500 ;
        RECT 79.900 43.400 81.700 43.700 ;
        RECT 81.000 43.100 81.300 43.400 ;
        RECT 83.000 43.100 83.400 43.500 ;
        RECT 78.200 42.800 79.200 43.100 ;
        RECT 78.800 41.100 79.200 42.800 ;
        RECT 81.000 41.100 81.400 43.100 ;
        RECT 83.100 41.100 83.700 43.100 ;
        RECT 85.400 41.100 85.800 45.400 ;
        RECT 87.000 46.100 87.400 47.900 ;
        RECT 88.700 47.200 89.000 47.900 ;
        RECT 89.500 47.700 91.300 47.900 ;
        RECT 91.800 47.700 92.200 49.900 ;
        RECT 93.900 49.200 94.500 49.900 ;
        RECT 93.900 48.900 94.600 49.200 ;
        RECT 96.200 48.900 96.600 49.900 ;
        RECT 98.400 49.200 98.800 49.900 ;
        RECT 98.400 48.900 99.400 49.200 ;
        RECT 94.200 48.500 94.600 48.900 ;
        RECT 96.300 48.600 96.600 48.900 ;
        RECT 96.300 48.300 97.700 48.600 ;
        RECT 97.300 48.200 97.700 48.300 ;
        RECT 98.200 48.200 98.600 48.600 ;
        RECT 99.000 48.500 99.400 48.900 ;
        RECT 93.300 47.700 93.700 47.800 ;
        RECT 91.800 47.400 93.700 47.700 ;
        RECT 90.600 47.200 91.000 47.400 ;
        RECT 87.800 47.100 88.200 47.200 ;
        RECT 88.600 47.100 89.900 47.200 ;
        RECT 87.800 46.800 89.900 47.100 ;
        RECT 90.600 46.900 91.400 47.200 ;
        RECT 91.000 46.800 91.400 46.900 ;
        RECT 87.000 45.800 88.900 46.100 ;
        RECT 87.000 41.100 87.400 45.800 ;
        RECT 88.600 45.200 88.900 45.800 ;
        RECT 87.800 44.400 88.200 45.200 ;
        RECT 88.600 45.100 89.000 45.200 ;
        RECT 89.600 45.100 89.900 46.800 ;
        RECT 90.200 45.800 90.600 46.600 ;
        RECT 91.800 45.700 92.200 47.400 ;
        RECT 95.300 47.100 95.700 47.200 ;
        RECT 98.200 47.100 98.500 48.200 ;
        RECT 100.600 47.500 101.000 49.900 ;
        RECT 104.300 48.200 104.700 49.900 ;
        RECT 103.800 47.900 104.700 48.200 ;
        RECT 105.400 47.900 105.800 49.900 ;
        RECT 106.200 48.000 106.600 49.900 ;
        RECT 107.800 48.000 108.200 49.900 ;
        RECT 109.400 48.200 109.800 49.900 ;
        RECT 106.200 47.900 108.200 48.000 ;
        RECT 109.300 47.900 109.800 48.200 ;
        RECT 99.800 47.100 100.600 47.200 ;
        RECT 95.100 46.800 100.600 47.100 ;
        RECT 101.400 47.100 101.800 47.200 ;
        RECT 103.000 47.100 103.400 47.600 ;
        RECT 101.400 46.800 103.400 47.100 ;
        RECT 94.200 46.400 94.600 46.500 ;
        RECT 92.700 46.100 94.600 46.400 ;
        RECT 92.700 46.000 93.100 46.100 ;
        RECT 93.500 45.700 93.900 45.800 ;
        RECT 91.800 45.400 93.900 45.700 ;
        RECT 88.600 44.800 89.300 45.100 ;
        RECT 89.600 44.800 90.100 45.100 ;
        RECT 89.000 44.200 89.300 44.800 ;
        RECT 89.000 43.800 89.400 44.200 ;
        RECT 89.700 41.100 90.100 44.800 ;
        RECT 91.800 41.100 92.200 45.400 ;
        RECT 95.100 45.200 95.400 46.800 ;
        RECT 98.700 46.700 99.100 46.800 ;
        RECT 98.200 46.200 98.600 46.300 ;
        RECT 99.500 46.200 99.900 46.300 ;
        RECT 97.400 45.900 99.900 46.200 ;
        RECT 103.800 46.100 104.200 47.900 ;
        RECT 105.500 47.200 105.800 47.900 ;
        RECT 106.300 47.700 108.100 47.900 ;
        RECT 107.400 47.200 107.800 47.400 ;
        RECT 109.300 47.200 109.600 47.900 ;
        RECT 111.000 47.600 111.400 49.900 ;
        RECT 112.600 47.600 113.000 49.900 ;
        RECT 114.200 47.600 114.600 49.900 ;
        RECT 115.800 47.600 116.200 49.900 ;
        RECT 117.400 47.600 117.800 49.900 ;
        RECT 119.000 48.000 119.400 49.900 ;
        RECT 120.600 48.000 121.000 49.900 ;
        RECT 119.000 47.900 121.000 48.000 ;
        RECT 121.400 47.900 121.800 49.900 ;
        RECT 122.500 48.200 122.900 49.900 ;
        RECT 122.500 47.900 123.400 48.200 ;
        RECT 119.100 47.700 120.900 47.900 ;
        RECT 110.100 47.300 111.400 47.600 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 105.400 47.100 106.700 47.200 ;
        RECT 104.600 46.800 106.700 47.100 ;
        RECT 107.400 46.900 108.200 47.200 ;
        RECT 107.800 46.800 108.200 46.900 ;
        RECT 109.300 46.800 109.800 47.200 ;
        RECT 97.400 45.800 97.800 45.900 ;
        RECT 103.800 45.800 105.700 46.100 ;
        RECT 98.200 45.500 101.000 45.600 ;
        RECT 98.100 45.400 101.000 45.500 ;
        RECT 94.200 44.900 95.400 45.200 ;
        RECT 96.100 45.300 101.000 45.400 ;
        RECT 96.100 45.100 98.500 45.300 ;
        RECT 94.200 44.400 94.500 44.900 ;
        RECT 93.800 44.000 94.500 44.400 ;
        RECT 95.300 44.500 95.700 44.600 ;
        RECT 96.100 44.500 96.400 45.100 ;
        RECT 95.300 44.200 96.400 44.500 ;
        RECT 96.700 44.500 99.400 44.800 ;
        RECT 96.700 44.400 97.100 44.500 ;
        RECT 99.000 44.400 99.400 44.500 ;
        RECT 95.900 43.700 96.300 43.800 ;
        RECT 97.300 43.700 97.700 43.800 ;
        RECT 94.200 43.100 94.600 43.500 ;
        RECT 95.900 43.400 97.700 43.700 ;
        RECT 96.300 43.100 96.600 43.400 ;
        RECT 99.000 43.100 99.400 43.500 ;
        RECT 93.900 41.100 94.500 43.100 ;
        RECT 96.200 41.100 96.600 43.100 ;
        RECT 98.400 42.800 99.400 43.100 ;
        RECT 98.400 41.100 98.800 42.800 ;
        RECT 100.600 41.100 101.000 45.300 ;
        RECT 103.800 41.100 104.200 45.800 ;
        RECT 105.400 45.200 105.700 45.800 ;
        RECT 104.600 44.400 105.000 45.200 ;
        RECT 105.400 45.100 105.800 45.200 ;
        RECT 106.400 45.100 106.700 46.800 ;
        RECT 107.000 45.800 107.400 46.600 ;
        RECT 109.300 45.100 109.600 46.800 ;
        RECT 110.100 46.500 110.400 47.300 ;
        RECT 111.800 47.200 113.000 47.600 ;
        RECT 113.500 47.200 114.600 47.600 ;
        RECT 115.100 47.200 116.200 47.600 ;
        RECT 116.900 47.200 117.800 47.600 ;
        RECT 119.400 47.200 119.800 47.400 ;
        RECT 121.400 47.200 121.700 47.900 ;
        RECT 109.900 46.100 110.400 46.500 ;
        RECT 110.100 45.100 110.400 46.100 ;
        RECT 110.900 46.200 111.300 46.600 ;
        RECT 110.900 45.800 111.400 46.200 ;
        RECT 111.800 45.800 112.200 47.200 ;
        RECT 113.500 46.900 113.900 47.200 ;
        RECT 115.100 46.900 115.500 47.200 ;
        RECT 116.900 46.900 117.300 47.200 ;
        RECT 118.200 46.900 118.600 47.200 ;
        RECT 112.600 46.500 113.900 46.900 ;
        RECT 114.300 46.500 115.500 46.900 ;
        RECT 116.000 46.500 117.300 46.900 ;
        RECT 117.700 46.500 118.600 46.900 ;
        RECT 119.000 46.900 119.800 47.200 ;
        RECT 120.500 47.100 121.800 47.200 ;
        RECT 122.200 47.100 122.600 47.200 ;
        RECT 119.000 46.800 119.400 46.900 ;
        RECT 120.500 46.800 122.600 47.100 ;
        RECT 113.500 45.800 113.900 46.500 ;
        RECT 115.100 45.800 115.500 46.500 ;
        RECT 116.900 45.800 117.300 46.500 ;
        RECT 119.800 45.800 120.200 46.600 ;
        RECT 111.800 45.400 113.000 45.800 ;
        RECT 113.500 45.400 114.600 45.800 ;
        RECT 115.100 45.400 116.200 45.800 ;
        RECT 116.900 45.400 117.800 45.800 ;
        RECT 105.400 44.800 106.100 45.100 ;
        RECT 106.400 44.800 106.900 45.100 ;
        RECT 105.800 44.200 106.100 44.800 ;
        RECT 105.800 43.800 106.200 44.200 ;
        RECT 106.500 41.100 106.900 44.800 ;
        RECT 109.300 44.600 109.800 45.100 ;
        RECT 110.100 44.800 111.400 45.100 ;
        RECT 109.400 41.100 109.800 44.600 ;
        RECT 111.000 41.100 111.400 44.800 ;
        RECT 112.600 41.100 113.000 45.400 ;
        RECT 114.200 41.100 114.600 45.400 ;
        RECT 115.800 41.100 116.200 45.400 ;
        RECT 117.400 41.100 117.800 45.400 ;
        RECT 120.500 45.100 120.800 46.800 ;
        RECT 123.000 46.100 123.400 47.900 ;
        RECT 124.600 47.700 125.000 49.900 ;
        RECT 126.700 49.200 127.300 49.900 ;
        RECT 126.700 48.900 127.400 49.200 ;
        RECT 129.000 48.900 129.400 49.900 ;
        RECT 131.200 49.200 131.600 49.900 ;
        RECT 131.200 48.900 132.200 49.200 ;
        RECT 127.000 48.500 127.400 48.900 ;
        RECT 129.100 48.600 129.400 48.900 ;
        RECT 129.100 48.300 130.500 48.600 ;
        RECT 130.100 48.200 130.500 48.300 ;
        RECT 131.000 48.200 131.400 48.600 ;
        RECT 131.800 48.500 132.200 48.900 ;
        RECT 126.100 47.700 126.500 47.800 ;
        RECT 123.800 46.800 124.200 47.600 ;
        RECT 124.600 47.400 126.500 47.700 ;
        RECT 121.400 45.800 123.400 46.100 ;
        RECT 121.400 45.200 121.700 45.800 ;
        RECT 121.400 45.100 121.800 45.200 ;
        RECT 120.300 44.800 120.800 45.100 ;
        RECT 121.100 44.800 121.800 45.100 ;
        RECT 120.300 41.100 120.700 44.800 ;
        RECT 121.100 44.200 121.400 44.800 ;
        RECT 122.200 44.400 122.600 45.200 ;
        RECT 121.000 43.800 121.400 44.200 ;
        RECT 123.000 41.100 123.400 45.800 ;
        RECT 124.600 45.700 125.000 47.400 ;
        RECT 128.100 47.100 128.500 47.200 ;
        RECT 131.000 47.100 131.300 48.200 ;
        RECT 133.400 47.500 133.800 49.900 ;
        RECT 134.200 47.600 134.600 49.900 ;
        RECT 135.800 48.200 136.200 49.900 ;
        RECT 138.700 48.200 139.100 49.900 ;
        RECT 135.800 47.900 136.300 48.200 ;
        RECT 134.200 47.300 135.500 47.600 ;
        RECT 132.600 47.100 133.400 47.200 ;
        RECT 127.900 46.800 133.400 47.100 ;
        RECT 127.000 46.400 127.400 46.500 ;
        RECT 125.500 46.100 127.400 46.400 ;
        RECT 127.900 46.200 128.200 46.800 ;
        RECT 131.500 46.700 131.900 46.800 ;
        RECT 132.300 46.200 132.700 46.300 ;
        RECT 134.300 46.200 134.700 46.600 ;
        RECT 125.500 46.000 125.900 46.100 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 130.200 45.900 132.700 46.200 ;
        RECT 130.200 45.800 130.600 45.900 ;
        RECT 134.200 45.800 134.700 46.200 ;
        RECT 135.200 46.500 135.500 47.300 ;
        RECT 136.000 47.200 136.300 47.900 ;
        RECT 135.800 46.800 136.300 47.200 ;
        RECT 135.200 46.100 135.700 46.500 ;
        RECT 126.300 45.700 126.700 45.800 ;
        RECT 124.600 45.400 126.700 45.700 ;
        RECT 123.800 44.100 124.200 44.200 ;
        RECT 124.600 44.100 125.000 45.400 ;
        RECT 127.900 45.200 128.200 45.800 ;
        RECT 131.000 45.500 133.800 45.600 ;
        RECT 130.900 45.400 133.800 45.500 ;
        RECT 127.000 44.900 128.200 45.200 ;
        RECT 128.900 45.300 133.800 45.400 ;
        RECT 128.900 45.100 131.300 45.300 ;
        RECT 127.000 44.400 127.300 44.900 ;
        RECT 123.800 43.800 125.000 44.100 ;
        RECT 126.600 44.000 127.300 44.400 ;
        RECT 128.100 44.500 128.500 44.600 ;
        RECT 128.900 44.500 129.200 45.100 ;
        RECT 128.100 44.200 129.200 44.500 ;
        RECT 129.500 44.500 132.200 44.800 ;
        RECT 129.500 44.400 129.900 44.500 ;
        RECT 131.800 44.400 132.200 44.500 ;
        RECT 124.600 41.100 125.000 43.800 ;
        RECT 128.700 43.700 129.100 43.800 ;
        RECT 130.100 43.700 130.500 43.800 ;
        RECT 127.000 43.100 127.400 43.500 ;
        RECT 128.700 43.400 130.500 43.700 ;
        RECT 129.100 43.100 129.400 43.400 ;
        RECT 131.800 43.100 132.200 43.500 ;
        RECT 126.700 41.100 127.300 43.100 ;
        RECT 129.000 41.100 129.400 43.100 ;
        RECT 131.200 42.800 132.200 43.100 ;
        RECT 131.200 41.100 131.600 42.800 ;
        RECT 133.400 41.100 133.800 45.300 ;
        RECT 135.200 45.100 135.500 46.100 ;
        RECT 136.000 45.100 136.300 46.800 ;
        RECT 134.200 44.800 135.500 45.100 ;
        RECT 134.200 41.100 134.600 44.800 ;
        RECT 135.800 44.600 136.300 45.100 ;
        RECT 138.200 47.900 139.100 48.200 ;
        RECT 135.800 41.100 136.200 44.600 ;
        RECT 138.200 41.100 138.600 47.900 ;
        RECT 139.800 47.500 140.200 49.900 ;
        RECT 142.000 49.200 142.400 49.900 ;
        RECT 141.400 48.900 142.400 49.200 ;
        RECT 144.200 48.900 144.600 49.900 ;
        RECT 146.300 49.200 146.900 49.900 ;
        RECT 146.200 48.900 146.900 49.200 ;
        RECT 148.600 49.100 149.000 49.900 ;
        RECT 152.900 49.200 153.300 49.500 ;
        RECT 149.400 49.100 149.800 49.200 ;
        RECT 141.400 48.500 141.800 48.900 ;
        RECT 144.200 48.600 144.500 48.900 ;
        RECT 142.200 48.200 142.600 48.600 ;
        RECT 143.100 48.300 144.500 48.600 ;
        RECT 146.200 48.500 146.600 48.900 ;
        RECT 148.600 48.800 149.800 49.100 ;
        RECT 152.600 48.800 153.300 49.200 ;
        RECT 143.100 48.200 143.500 48.300 ;
        RECT 139.000 47.100 139.400 47.200 ;
        RECT 140.200 47.100 141.000 47.200 ;
        RECT 142.300 47.100 142.600 48.200 ;
        RECT 147.100 47.700 147.500 47.800 ;
        RECT 148.600 47.700 149.000 48.800 ;
        RECT 152.900 48.000 153.300 48.800 ;
        RECT 155.000 48.500 155.400 49.500 ;
        RECT 147.100 47.400 149.000 47.700 ;
        RECT 145.100 47.100 145.500 47.200 ;
        RECT 139.000 46.800 145.700 47.100 ;
        RECT 141.700 46.700 142.100 46.800 ;
        RECT 140.900 46.200 141.300 46.300 ;
        RECT 142.200 46.200 142.600 46.300 ;
        RECT 140.900 45.900 143.400 46.200 ;
        RECT 143.000 45.800 143.400 45.900 ;
        RECT 144.600 46.100 145.000 46.200 ;
        RECT 145.400 46.100 145.700 46.800 ;
        RECT 146.200 46.400 146.600 46.500 ;
        RECT 146.200 46.100 148.100 46.400 ;
        RECT 144.600 45.800 145.700 46.100 ;
        RECT 147.700 46.000 148.100 46.100 ;
        RECT 139.800 45.500 142.600 45.600 ;
        RECT 139.800 45.400 142.700 45.500 ;
        RECT 139.800 45.300 144.700 45.400 ;
        RECT 139.800 41.100 140.200 45.300 ;
        RECT 142.300 45.100 144.700 45.300 ;
        RECT 141.400 44.500 144.100 44.800 ;
        RECT 141.400 44.400 141.800 44.500 ;
        RECT 143.700 44.400 144.100 44.500 ;
        RECT 144.400 44.500 144.700 45.100 ;
        RECT 145.400 45.200 145.700 45.800 ;
        RECT 146.900 45.700 147.300 45.800 ;
        RECT 148.600 45.700 149.000 47.400 ;
        RECT 152.500 47.700 153.300 48.000 ;
        RECT 152.500 47.500 152.900 47.700 ;
        RECT 152.500 47.200 152.800 47.500 ;
        RECT 155.100 47.400 155.400 48.500 ;
        RECT 157.100 48.200 157.500 49.900 ;
        RECT 156.600 47.900 157.500 48.200 ;
        RECT 158.200 47.900 158.600 49.900 ;
        RECT 159.000 48.000 159.400 49.900 ;
        RECT 160.600 48.000 161.000 49.900 ;
        RECT 162.200 48.200 162.600 49.900 ;
        RECT 159.000 47.900 161.000 48.000 ;
        RECT 162.100 47.900 162.600 48.200 ;
        RECT 151.800 46.800 152.800 47.200 ;
        RECT 153.300 47.100 155.400 47.400 ;
        RECT 153.300 46.900 153.800 47.100 ;
        RECT 146.900 45.400 149.000 45.700 ;
        RECT 151.800 45.400 152.200 46.200 ;
        RECT 145.400 44.900 146.600 45.200 ;
        RECT 145.100 44.500 145.500 44.600 ;
        RECT 144.400 44.200 145.500 44.500 ;
        RECT 146.300 44.400 146.600 44.900 ;
        RECT 146.300 44.000 147.000 44.400 ;
        RECT 143.100 43.700 143.500 43.800 ;
        RECT 144.500 43.700 144.900 43.800 ;
        RECT 141.400 43.100 141.800 43.500 ;
        RECT 143.100 43.400 144.900 43.700 ;
        RECT 144.200 43.100 144.500 43.400 ;
        RECT 146.200 43.100 146.600 43.500 ;
        RECT 141.400 42.800 142.400 43.100 ;
        RECT 142.000 41.100 142.400 42.800 ;
        RECT 144.200 41.100 144.600 43.100 ;
        RECT 146.300 41.100 146.900 43.100 ;
        RECT 148.600 41.100 149.000 45.400 ;
        RECT 152.500 44.900 152.800 46.800 ;
        RECT 153.100 46.500 153.800 46.900 ;
        RECT 155.800 46.800 156.200 47.600 ;
        RECT 153.500 45.500 153.800 46.500 ;
        RECT 154.200 45.800 154.600 46.600 ;
        RECT 155.000 45.800 155.400 46.600 ;
        RECT 156.600 46.100 157.000 47.900 ;
        RECT 158.300 47.200 158.600 47.900 ;
        RECT 159.100 47.700 160.900 47.900 ;
        RECT 160.200 47.200 160.600 47.400 ;
        RECT 162.100 47.200 162.400 47.900 ;
        RECT 163.800 47.600 164.200 49.900 ;
        RECT 165.400 48.200 165.800 49.900 ;
        RECT 162.900 47.300 164.200 47.600 ;
        RECT 165.300 47.900 165.800 48.200 ;
        RECT 158.200 46.800 159.500 47.200 ;
        RECT 160.200 46.900 161.000 47.200 ;
        RECT 160.600 46.800 161.000 46.900 ;
        RECT 162.100 46.800 162.600 47.200 ;
        RECT 156.600 45.800 158.500 46.100 ;
        RECT 153.500 45.200 155.400 45.500 ;
        RECT 152.500 44.600 153.300 44.900 ;
        RECT 152.900 41.100 153.300 44.600 ;
        RECT 155.100 43.500 155.400 45.200 ;
        RECT 155.000 41.500 155.400 43.500 ;
        RECT 156.600 41.100 157.000 45.800 ;
        RECT 158.200 45.200 158.500 45.800 ;
        RECT 157.400 44.400 157.800 45.200 ;
        RECT 158.200 45.100 158.600 45.200 ;
        RECT 159.200 45.100 159.500 46.800 ;
        RECT 159.800 45.800 160.200 46.600 ;
        RECT 162.100 45.100 162.400 46.800 ;
        RECT 162.900 46.500 163.200 47.300 ;
        RECT 162.700 46.100 163.200 46.500 ;
        RECT 162.900 45.100 163.200 46.100 ;
        RECT 165.300 47.200 165.600 47.900 ;
        RECT 167.000 47.600 167.400 49.900 ;
        RECT 168.600 48.200 169.000 49.900 ;
        RECT 166.100 47.300 167.400 47.600 ;
        RECT 168.500 47.900 169.000 48.200 ;
        RECT 165.300 46.800 165.800 47.200 ;
        RECT 165.300 45.100 165.600 46.800 ;
        RECT 166.100 46.500 166.400 47.300 ;
        RECT 165.900 46.100 166.400 46.500 ;
        RECT 166.100 45.100 166.400 46.100 ;
        RECT 168.500 47.200 168.800 47.900 ;
        RECT 170.200 47.600 170.600 49.900 ;
        RECT 169.300 47.300 170.600 47.600 ;
        RECT 171.000 47.600 171.400 49.900 ;
        RECT 172.600 48.200 173.000 49.900 ;
        RECT 172.600 47.900 173.100 48.200 ;
        RECT 171.000 47.300 172.300 47.600 ;
        RECT 168.500 46.800 169.000 47.200 ;
        RECT 168.500 45.100 168.800 46.800 ;
        RECT 169.300 46.500 169.600 47.300 ;
        RECT 169.100 46.100 169.600 46.500 ;
        RECT 169.300 45.100 169.600 46.100 ;
        RECT 172.000 46.500 172.300 47.300 ;
        RECT 172.800 47.200 173.100 47.900 ;
        RECT 174.200 47.600 174.600 49.900 ;
        RECT 175.800 48.200 176.200 49.900 ;
        RECT 178.200 48.200 178.600 49.900 ;
        RECT 175.800 47.900 176.300 48.200 ;
        RECT 174.200 47.300 175.500 47.600 ;
        RECT 172.600 46.800 173.100 47.200 ;
        RECT 172.000 46.100 172.500 46.500 ;
        RECT 172.000 45.100 172.300 46.100 ;
        RECT 172.800 45.100 173.100 46.800 ;
        RECT 175.200 46.500 175.500 47.300 ;
        RECT 176.000 47.200 176.300 47.900 ;
        RECT 175.800 46.800 176.300 47.200 ;
        RECT 175.200 46.100 175.700 46.500 ;
        RECT 175.200 45.100 175.500 46.100 ;
        RECT 176.000 45.100 176.300 46.800 ;
        RECT 158.200 44.800 158.900 45.100 ;
        RECT 159.200 44.800 159.700 45.100 ;
        RECT 158.600 44.200 158.900 44.800 ;
        RECT 158.600 43.800 159.000 44.200 ;
        RECT 159.300 41.100 159.700 44.800 ;
        RECT 162.100 44.600 162.600 45.100 ;
        RECT 162.900 44.800 164.200 45.100 ;
        RECT 162.200 41.100 162.600 44.600 ;
        RECT 163.800 41.100 164.200 44.800 ;
        RECT 165.300 44.600 165.800 45.100 ;
        RECT 166.100 44.800 167.400 45.100 ;
        RECT 165.400 41.100 165.800 44.600 ;
        RECT 167.000 41.100 167.400 44.800 ;
        RECT 168.500 44.600 169.000 45.100 ;
        RECT 169.300 44.800 170.600 45.100 ;
        RECT 168.600 41.100 169.000 44.600 ;
        RECT 170.200 41.100 170.600 44.800 ;
        RECT 171.000 44.800 172.300 45.100 ;
        RECT 171.000 41.100 171.400 44.800 ;
        RECT 172.600 44.600 173.100 45.100 ;
        RECT 174.200 44.800 175.500 45.100 ;
        RECT 172.600 41.100 173.000 44.600 ;
        RECT 174.200 41.100 174.600 44.800 ;
        RECT 175.800 44.600 176.300 45.100 ;
        RECT 178.100 47.900 178.600 48.200 ;
        RECT 178.100 47.200 178.400 47.900 ;
        RECT 179.800 47.600 180.200 49.900 ;
        RECT 178.900 47.300 180.200 47.600 ;
        RECT 181.400 47.600 181.800 49.900 ;
        RECT 183.000 47.600 183.400 49.900 ;
        RECT 184.600 47.600 185.000 49.900 ;
        RECT 186.200 47.600 186.600 49.900 ;
        RECT 187.800 48.500 188.200 49.500 ;
        RECT 189.900 49.200 190.300 49.500 ;
        RECT 189.900 48.800 190.600 49.200 ;
        RECT 178.100 46.800 178.600 47.200 ;
        RECT 178.100 45.100 178.400 46.800 ;
        RECT 178.900 46.500 179.200 47.300 ;
        RECT 181.400 47.200 182.300 47.600 ;
        RECT 183.000 47.200 184.100 47.600 ;
        RECT 184.600 47.200 185.700 47.600 ;
        RECT 186.200 47.200 187.400 47.600 ;
        RECT 180.600 46.900 181.000 47.200 ;
        RECT 181.900 46.900 182.300 47.200 ;
        RECT 183.700 46.900 184.100 47.200 ;
        RECT 185.300 46.900 185.700 47.200 ;
        RECT 180.600 46.500 181.500 46.900 ;
        RECT 181.900 46.500 183.200 46.900 ;
        RECT 183.700 46.500 184.900 46.900 ;
        RECT 185.300 46.500 186.600 46.900 ;
        RECT 178.700 46.100 179.200 46.500 ;
        RECT 178.900 45.100 179.200 46.100 ;
        RECT 181.900 45.800 182.300 46.500 ;
        RECT 183.700 45.800 184.100 46.500 ;
        RECT 185.300 45.800 185.700 46.500 ;
        RECT 187.000 45.800 187.400 47.200 ;
        RECT 187.800 47.400 188.100 48.500 ;
        RECT 189.900 48.000 190.300 48.800 ;
        RECT 189.900 47.700 190.700 48.000 ;
        RECT 190.300 47.500 190.700 47.700 ;
        RECT 187.800 47.100 189.900 47.400 ;
        RECT 189.400 46.900 189.900 47.100 ;
        RECT 190.400 47.200 190.700 47.500 ;
        RECT 192.600 47.700 193.000 49.900 ;
        RECT 194.700 49.200 195.300 49.900 ;
        RECT 194.700 48.900 195.400 49.200 ;
        RECT 197.000 48.900 197.400 49.900 ;
        RECT 199.200 49.200 199.600 49.900 ;
        RECT 199.200 48.900 200.200 49.200 ;
        RECT 195.000 48.500 195.400 48.900 ;
        RECT 197.100 48.600 197.400 48.900 ;
        RECT 197.100 48.300 198.500 48.600 ;
        RECT 198.100 48.200 198.500 48.300 ;
        RECT 199.000 48.200 199.400 48.600 ;
        RECT 199.800 48.500 200.200 48.900 ;
        RECT 194.100 47.700 194.500 47.800 ;
        RECT 192.600 47.400 194.500 47.700 ;
        RECT 187.800 45.800 188.200 46.600 ;
        RECT 188.600 45.800 189.000 46.600 ;
        RECT 189.400 46.500 190.100 46.900 ;
        RECT 190.400 46.800 191.400 47.200 ;
        RECT 181.400 45.400 182.300 45.800 ;
        RECT 183.000 45.400 184.100 45.800 ;
        RECT 184.600 45.400 185.700 45.800 ;
        RECT 186.200 45.400 187.400 45.800 ;
        RECT 189.400 45.500 189.700 46.500 ;
        RECT 178.100 44.600 178.600 45.100 ;
        RECT 178.900 44.800 180.200 45.100 ;
        RECT 175.800 41.100 176.200 44.600 ;
        RECT 178.200 41.100 178.600 44.600 ;
        RECT 179.800 41.100 180.200 44.800 ;
        RECT 181.400 41.100 181.800 45.400 ;
        RECT 183.000 41.100 183.400 45.400 ;
        RECT 184.600 41.100 185.000 45.400 ;
        RECT 186.200 41.100 186.600 45.400 ;
        RECT 187.800 45.200 189.700 45.500 ;
        RECT 187.800 43.500 188.100 45.200 ;
        RECT 190.400 44.900 190.700 46.800 ;
        RECT 191.000 45.400 191.400 46.200 ;
        RECT 192.600 45.700 193.000 47.400 ;
        RECT 196.100 47.100 196.500 47.200 ;
        RECT 199.000 47.100 199.300 48.200 ;
        RECT 201.400 47.500 201.800 49.900 ;
        RECT 205.700 49.200 206.100 49.500 ;
        RECT 205.400 48.800 206.100 49.200 ;
        RECT 205.700 48.000 206.100 48.800 ;
        RECT 207.800 48.500 208.200 49.500 ;
        RECT 205.300 47.700 206.100 48.000 ;
        RECT 205.300 47.500 205.700 47.700 ;
        RECT 205.300 47.200 205.600 47.500 ;
        RECT 207.900 47.400 208.200 48.500 ;
        RECT 200.600 47.100 201.400 47.200 ;
        RECT 203.000 47.100 203.400 47.200 ;
        RECT 195.900 46.800 203.400 47.100 ;
        RECT 204.600 46.800 205.600 47.200 ;
        RECT 206.100 47.100 208.200 47.400 ;
        RECT 208.600 47.700 209.000 49.900 ;
        RECT 210.700 49.200 211.300 49.900 ;
        RECT 210.700 48.900 211.400 49.200 ;
        RECT 213.000 48.900 213.400 49.900 ;
        RECT 215.200 49.200 215.600 49.900 ;
        RECT 215.200 48.900 216.200 49.200 ;
        RECT 211.000 48.500 211.400 48.900 ;
        RECT 213.100 48.600 213.400 48.900 ;
        RECT 213.100 48.300 214.500 48.600 ;
        RECT 214.100 48.200 214.500 48.300 ;
        RECT 215.000 48.200 215.400 48.600 ;
        RECT 215.800 48.500 216.200 48.900 ;
        RECT 210.100 47.700 210.500 47.800 ;
        RECT 208.600 47.400 210.500 47.700 ;
        RECT 206.100 46.900 206.600 47.100 ;
        RECT 195.000 46.400 195.400 46.500 ;
        RECT 193.500 46.100 195.400 46.400 ;
        RECT 195.900 46.200 196.200 46.800 ;
        RECT 199.500 46.700 199.900 46.800 ;
        RECT 199.000 46.200 199.400 46.300 ;
        RECT 200.300 46.200 200.700 46.300 ;
        RECT 193.500 46.000 193.900 46.100 ;
        RECT 195.800 45.800 196.200 46.200 ;
        RECT 198.200 45.900 200.700 46.200 ;
        RECT 198.200 45.800 198.600 45.900 ;
        RECT 194.300 45.700 194.700 45.800 ;
        RECT 192.600 45.400 194.700 45.700 ;
        RECT 189.900 44.600 190.700 44.900 ;
        RECT 187.800 41.500 188.200 43.500 ;
        RECT 189.900 41.100 190.300 44.600 ;
        RECT 192.600 41.100 193.000 45.400 ;
        RECT 195.900 45.200 196.200 45.800 ;
        RECT 199.000 45.500 201.800 45.600 ;
        RECT 198.900 45.400 201.800 45.500 ;
        RECT 204.600 45.400 205.000 46.200 ;
        RECT 195.000 44.900 196.200 45.200 ;
        RECT 196.900 45.300 201.800 45.400 ;
        RECT 196.900 45.100 199.300 45.300 ;
        RECT 195.000 44.400 195.300 44.900 ;
        RECT 194.600 44.000 195.300 44.400 ;
        RECT 196.100 44.500 196.500 44.600 ;
        RECT 196.900 44.500 197.200 45.100 ;
        RECT 196.100 44.200 197.200 44.500 ;
        RECT 197.500 44.500 200.200 44.800 ;
        RECT 197.500 44.400 197.900 44.500 ;
        RECT 199.800 44.400 200.200 44.500 ;
        RECT 196.700 43.700 197.100 43.800 ;
        RECT 198.100 43.700 198.500 43.800 ;
        RECT 195.000 43.100 195.400 43.500 ;
        RECT 196.700 43.400 198.500 43.700 ;
        RECT 197.100 43.100 197.400 43.400 ;
        RECT 199.800 43.100 200.200 43.500 ;
        RECT 194.700 41.100 195.300 43.100 ;
        RECT 197.000 41.100 197.400 43.100 ;
        RECT 199.200 42.800 200.200 43.100 ;
        RECT 199.200 41.100 199.600 42.800 ;
        RECT 201.400 41.100 201.800 45.300 ;
        RECT 205.300 44.900 205.600 46.800 ;
        RECT 205.900 46.500 206.600 46.900 ;
        RECT 206.300 45.500 206.600 46.500 ;
        RECT 207.000 45.800 207.400 46.600 ;
        RECT 207.800 45.800 208.200 46.600 ;
        RECT 208.600 45.700 209.000 47.400 ;
        RECT 212.100 47.100 212.500 47.200 ;
        RECT 215.000 47.100 215.300 48.200 ;
        RECT 217.400 47.500 217.800 49.900 ;
        RECT 219.500 48.200 219.900 49.900 ;
        RECT 219.000 47.900 219.900 48.200 ;
        RECT 220.600 47.900 221.000 49.900 ;
        RECT 221.400 48.000 221.800 49.900 ;
        RECT 223.000 48.000 223.400 49.900 ;
        RECT 224.600 48.800 225.000 49.900 ;
        RECT 221.400 47.900 223.400 48.000 ;
        RECT 216.600 47.100 217.400 47.200 ;
        RECT 211.900 46.800 217.400 47.100 ;
        RECT 218.200 46.800 218.600 47.600 ;
        RECT 211.000 46.400 211.400 46.500 ;
        RECT 209.500 46.100 211.400 46.400 ;
        RECT 211.900 46.200 212.200 46.800 ;
        RECT 215.500 46.700 215.900 46.800 ;
        RECT 215.000 46.200 215.400 46.300 ;
        RECT 216.300 46.200 216.700 46.300 ;
        RECT 209.500 46.000 209.900 46.100 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 214.200 45.900 216.700 46.200 ;
        RECT 219.000 46.100 219.400 47.900 ;
        RECT 220.700 47.200 221.000 47.900 ;
        RECT 221.500 47.700 223.300 47.900 ;
        RECT 223.800 47.800 224.200 48.600 ;
        RECT 222.600 47.200 223.000 47.400 ;
        RECT 224.700 47.200 225.000 48.800 ;
        RECT 219.800 47.100 220.200 47.200 ;
        RECT 220.600 47.100 221.900 47.200 ;
        RECT 219.800 46.800 221.900 47.100 ;
        RECT 222.600 46.900 223.400 47.200 ;
        RECT 223.000 46.800 223.400 46.900 ;
        RECT 224.600 46.800 225.000 47.200 ;
        RECT 226.200 48.500 226.600 49.500 ;
        RECT 228.300 49.200 228.700 49.500 ;
        RECT 227.800 48.800 228.700 49.200 ;
        RECT 226.200 47.400 226.500 48.500 ;
        RECT 228.300 48.000 228.700 48.800 ;
        RECT 232.900 48.000 233.300 49.500 ;
        RECT 235.000 48.500 235.400 49.500 ;
        RECT 228.300 47.700 229.100 48.000 ;
        RECT 228.700 47.500 229.100 47.700 ;
        RECT 226.200 47.100 228.300 47.400 ;
        RECT 214.200 45.800 214.600 45.900 ;
        RECT 219.000 45.800 220.900 46.100 ;
        RECT 210.300 45.700 210.700 45.800 ;
        RECT 206.300 45.200 208.200 45.500 ;
        RECT 205.300 44.600 206.100 44.900 ;
        RECT 205.700 41.100 206.100 44.600 ;
        RECT 207.900 43.500 208.200 45.200 ;
        RECT 207.800 41.500 208.200 43.500 ;
        RECT 208.600 45.400 210.700 45.700 ;
        RECT 208.600 41.100 209.000 45.400 ;
        RECT 211.900 45.200 212.200 45.800 ;
        RECT 215.000 45.500 217.800 45.600 ;
        RECT 214.900 45.400 217.800 45.500 ;
        RECT 211.000 44.900 212.200 45.200 ;
        RECT 212.900 45.300 217.800 45.400 ;
        RECT 212.900 45.100 215.300 45.300 ;
        RECT 211.000 44.400 211.300 44.900 ;
        RECT 210.600 44.000 211.300 44.400 ;
        RECT 212.100 44.500 212.500 44.600 ;
        RECT 212.900 44.500 213.200 45.100 ;
        RECT 212.100 44.200 213.200 44.500 ;
        RECT 213.500 44.500 216.200 44.800 ;
        RECT 213.500 44.400 213.900 44.500 ;
        RECT 215.800 44.400 216.200 44.500 ;
        RECT 212.700 43.700 213.100 43.800 ;
        RECT 214.100 43.700 214.500 43.800 ;
        RECT 211.000 43.100 211.400 43.500 ;
        RECT 212.700 43.400 214.500 43.700 ;
        RECT 213.100 43.100 213.400 43.400 ;
        RECT 215.800 43.100 216.200 43.500 ;
        RECT 210.700 41.100 211.300 43.100 ;
        RECT 213.000 41.100 213.400 43.100 ;
        RECT 215.200 42.800 216.200 43.100 ;
        RECT 215.200 41.100 215.600 42.800 ;
        RECT 217.400 41.100 217.800 45.300 ;
        RECT 219.000 41.100 219.400 45.800 ;
        RECT 220.600 45.200 220.900 45.800 ;
        RECT 219.800 44.400 220.200 45.200 ;
        RECT 220.600 45.100 221.000 45.200 ;
        RECT 221.600 45.100 221.900 46.800 ;
        RECT 222.200 45.800 222.600 46.600 ;
        RECT 224.700 45.100 225.000 46.800 ;
        RECT 227.800 46.900 228.300 47.100 ;
        RECT 228.800 47.200 229.100 47.500 ;
        RECT 232.500 47.700 233.300 48.000 ;
        RECT 232.500 47.500 232.900 47.700 ;
        RECT 232.500 47.200 232.800 47.500 ;
        RECT 235.100 47.400 235.400 48.500 ;
        RECT 235.800 48.000 236.200 49.900 ;
        RECT 237.400 48.000 237.800 49.900 ;
        RECT 235.800 47.900 237.800 48.000 ;
        RECT 238.200 47.900 238.600 49.900 ;
        RECT 239.300 48.200 239.700 49.900 ;
        RECT 239.300 47.900 240.200 48.200 ;
        RECT 235.900 47.700 237.700 47.900 ;
        RECT 225.400 45.400 225.800 46.200 ;
        RECT 226.200 45.800 226.600 46.600 ;
        RECT 227.000 45.800 227.400 46.600 ;
        RECT 227.800 46.500 228.500 46.900 ;
        RECT 228.800 46.800 229.800 47.200 ;
        RECT 231.800 47.100 232.800 47.200 ;
        RECT 230.200 46.800 232.800 47.100 ;
        RECT 233.300 47.100 235.400 47.400 ;
        RECT 236.200 47.200 236.600 47.400 ;
        RECT 238.200 47.200 238.500 47.900 ;
        RECT 233.300 46.900 233.800 47.100 ;
        RECT 227.800 45.500 228.100 46.500 ;
        RECT 226.200 45.200 228.100 45.500 ;
        RECT 220.600 44.800 221.300 45.100 ;
        RECT 221.600 44.800 222.100 45.100 ;
        RECT 221.000 44.200 221.300 44.800 ;
        RECT 221.000 43.800 221.400 44.200 ;
        RECT 221.700 41.100 222.100 44.800 ;
        RECT 224.600 44.700 225.500 45.100 ;
        RECT 225.100 41.100 225.500 44.700 ;
        RECT 226.200 43.500 226.500 45.200 ;
        RECT 228.800 44.900 229.100 46.800 ;
        RECT 229.400 46.100 229.800 46.200 ;
        RECT 230.200 46.100 230.500 46.800 ;
        RECT 229.400 45.800 230.500 46.100 ;
        RECT 231.000 46.100 231.400 46.200 ;
        RECT 231.800 46.100 232.200 46.200 ;
        RECT 231.000 45.800 232.200 46.100 ;
        RECT 229.400 45.400 229.800 45.800 ;
        RECT 231.800 45.400 232.200 45.800 ;
        RECT 228.300 44.600 229.100 44.900 ;
        RECT 232.500 44.900 232.800 46.800 ;
        RECT 233.100 46.500 233.800 46.900 ;
        RECT 235.800 46.900 236.600 47.200 ;
        RECT 237.300 47.100 238.600 47.200 ;
        RECT 239.000 47.100 239.400 47.200 ;
        RECT 235.800 46.800 236.200 46.900 ;
        RECT 237.300 46.800 239.400 47.100 ;
        RECT 233.500 45.500 233.800 46.500 ;
        RECT 234.200 45.800 234.600 46.600 ;
        RECT 235.000 45.800 235.400 46.600 ;
        RECT 236.600 45.800 237.000 46.600 ;
        RECT 233.500 45.200 235.400 45.500 ;
        RECT 232.500 44.600 233.300 44.900 ;
        RECT 226.200 41.500 226.600 43.500 ;
        RECT 228.300 41.100 228.700 44.600 ;
        RECT 232.900 41.100 233.300 44.600 ;
        RECT 235.100 43.500 235.400 45.200 ;
        RECT 237.300 45.100 237.600 46.800 ;
        RECT 239.800 46.100 240.200 47.900 ;
        RECT 240.600 46.800 241.000 47.600 ;
        RECT 241.400 47.500 241.800 49.900 ;
        RECT 243.600 49.200 244.000 49.900 ;
        RECT 243.000 48.900 244.000 49.200 ;
        RECT 245.800 48.900 246.200 49.900 ;
        RECT 247.900 49.200 248.500 49.900 ;
        RECT 247.800 48.900 248.500 49.200 ;
        RECT 243.000 48.500 243.400 48.900 ;
        RECT 245.800 48.600 246.100 48.900 ;
        RECT 243.800 48.200 244.200 48.600 ;
        RECT 244.700 48.300 246.100 48.600 ;
        RECT 247.800 48.500 248.200 48.900 ;
        RECT 244.700 48.200 245.100 48.300 ;
        RECT 241.800 47.100 242.600 47.200 ;
        RECT 243.900 47.100 244.200 48.200 ;
        RECT 248.700 47.700 249.100 47.800 ;
        RECT 250.200 47.700 250.600 49.900 ;
        RECT 248.700 47.400 250.600 47.700 ;
        RECT 246.700 47.100 247.100 47.200 ;
        RECT 241.800 46.800 247.300 47.100 ;
        RECT 243.300 46.700 243.700 46.800 ;
        RECT 238.200 45.800 240.200 46.100 ;
        RECT 242.500 46.200 242.900 46.300 ;
        RECT 243.800 46.200 244.200 46.300 ;
        RECT 242.500 45.900 245.000 46.200 ;
        RECT 244.600 45.800 245.000 45.900 ;
        RECT 238.200 45.200 238.500 45.800 ;
        RECT 238.200 45.100 238.600 45.200 ;
        RECT 235.000 41.500 235.400 43.500 ;
        RECT 237.100 44.800 237.600 45.100 ;
        RECT 237.900 44.800 238.600 45.100 ;
        RECT 237.100 41.100 237.500 44.800 ;
        RECT 237.900 44.200 238.200 44.800 ;
        RECT 239.000 44.400 239.400 45.200 ;
        RECT 237.800 43.800 238.200 44.200 ;
        RECT 239.800 41.100 240.200 45.800 ;
        RECT 241.400 45.500 244.200 45.600 ;
        RECT 241.400 45.400 244.300 45.500 ;
        RECT 241.400 45.300 246.300 45.400 ;
        RECT 241.400 41.100 241.800 45.300 ;
        RECT 243.900 45.100 246.300 45.300 ;
        RECT 243.000 44.500 245.700 44.800 ;
        RECT 243.000 44.400 243.400 44.500 ;
        RECT 245.300 44.400 245.700 44.500 ;
        RECT 246.000 44.500 246.300 45.100 ;
        RECT 247.000 45.200 247.300 46.800 ;
        RECT 247.800 46.400 248.200 46.500 ;
        RECT 247.800 46.100 249.700 46.400 ;
        RECT 249.300 46.000 249.700 46.100 ;
        RECT 248.500 45.700 248.900 45.800 ;
        RECT 250.200 45.700 250.600 47.400 ;
        RECT 248.500 45.400 250.600 45.700 ;
        RECT 247.000 44.900 248.200 45.200 ;
        RECT 246.700 44.500 247.100 44.600 ;
        RECT 246.000 44.200 247.100 44.500 ;
        RECT 247.900 44.400 248.200 44.900 ;
        RECT 247.900 44.000 248.600 44.400 ;
        RECT 244.700 43.700 245.100 43.800 ;
        RECT 246.100 43.700 246.500 43.800 ;
        RECT 243.000 43.100 243.400 43.500 ;
        RECT 244.700 43.400 246.500 43.700 ;
        RECT 245.800 43.100 246.100 43.400 ;
        RECT 247.800 43.100 248.200 43.500 ;
        RECT 243.000 42.800 244.000 43.100 ;
        RECT 243.600 41.100 244.000 42.800 ;
        RECT 245.800 41.100 246.200 43.100 ;
        RECT 247.900 41.100 248.500 43.100 ;
        RECT 250.200 41.100 250.600 45.400 ;
        RECT 0.600 35.700 1.000 39.900 ;
        RECT 2.800 38.200 3.200 39.900 ;
        RECT 2.200 37.900 3.200 38.200 ;
        RECT 5.000 37.900 5.400 39.900 ;
        RECT 7.100 37.900 7.700 39.900 ;
        RECT 2.200 37.500 2.600 37.900 ;
        RECT 5.000 37.600 5.300 37.900 ;
        RECT 3.900 37.300 5.700 37.600 ;
        RECT 7.000 37.500 7.400 37.900 ;
        RECT 3.900 37.200 4.300 37.300 ;
        RECT 5.300 37.200 5.700 37.300 ;
        RECT 2.200 36.500 2.600 36.600 ;
        RECT 4.500 36.500 4.900 36.600 ;
        RECT 2.200 36.200 4.900 36.500 ;
        RECT 5.200 36.500 6.300 36.800 ;
        RECT 5.200 35.900 5.500 36.500 ;
        RECT 5.900 36.400 6.300 36.500 ;
        RECT 7.100 36.600 7.800 37.000 ;
        RECT 7.100 36.100 7.400 36.600 ;
        RECT 3.100 35.700 5.500 35.900 ;
        RECT 0.600 35.600 5.500 35.700 ;
        RECT 6.200 35.800 7.400 36.100 ;
        RECT 0.600 35.500 3.500 35.600 ;
        RECT 0.600 35.400 3.400 35.500 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 1.700 34.800 4.200 35.100 ;
        RECT 1.700 34.700 2.100 34.800 ;
        RECT 3.000 34.700 3.400 34.800 ;
        RECT 2.500 34.200 2.900 34.300 ;
        RECT 6.200 34.200 6.500 35.800 ;
        RECT 9.400 35.600 9.800 39.900 ;
        RECT 12.100 39.200 12.500 39.900 ;
        RECT 12.100 38.800 13.000 39.200 ;
        RECT 12.100 36.400 12.500 38.800 ;
        RECT 14.200 37.500 14.600 39.500 ;
        RECT 11.700 36.100 12.500 36.400 ;
        RECT 7.700 35.300 9.800 35.600 ;
        RECT 7.700 35.200 8.100 35.300 ;
        RECT 9.400 35.100 9.800 35.300 ;
        RECT 11.000 35.100 11.400 35.600 ;
        RECT 8.500 34.900 8.900 35.000 ;
        RECT 7.000 34.600 8.900 34.900 ;
        RECT 9.400 34.800 11.400 35.100 ;
        RECT 7.000 34.500 7.400 34.600 ;
        RECT 1.000 33.900 6.500 34.200 ;
        RECT 1.000 33.800 1.800 33.900 ;
        RECT 0.600 31.100 1.000 33.500 ;
        RECT 3.100 32.800 3.400 33.900 ;
        RECT 3.800 33.800 4.200 33.900 ;
        RECT 5.900 33.800 6.300 33.900 ;
        RECT 9.400 33.600 9.800 34.800 ;
        RECT 11.700 34.200 12.000 36.100 ;
        RECT 14.300 35.800 14.600 37.500 ;
        RECT 16.300 36.200 16.700 39.900 ;
        RECT 17.000 36.800 17.400 37.200 ;
        RECT 17.100 36.200 17.400 36.800 ;
        RECT 16.300 35.900 16.800 36.200 ;
        RECT 17.100 35.900 17.800 36.200 ;
        RECT 12.700 35.500 14.600 35.800 ;
        RECT 12.700 34.500 13.000 35.500 ;
        RECT 11.000 33.800 12.000 34.200 ;
        RECT 12.300 34.100 13.000 34.500 ;
        RECT 13.400 34.400 13.800 35.200 ;
        RECT 14.200 34.400 14.600 35.200 ;
        RECT 15.800 34.400 16.200 35.200 ;
        RECT 16.500 34.200 16.800 35.900 ;
        RECT 17.400 35.800 17.800 35.900 ;
        RECT 18.200 35.800 18.600 36.600 ;
        RECT 17.400 35.100 17.700 35.800 ;
        RECT 19.000 35.100 19.400 39.900 ;
        RECT 20.600 35.700 21.000 39.900 ;
        RECT 22.800 38.200 23.200 39.900 ;
        RECT 22.200 37.900 23.200 38.200 ;
        RECT 25.000 37.900 25.400 39.900 ;
        RECT 27.100 37.900 27.700 39.900 ;
        RECT 22.200 37.500 22.600 37.900 ;
        RECT 25.000 37.600 25.300 37.900 ;
        RECT 23.900 37.300 25.700 37.600 ;
        RECT 27.000 37.500 27.400 37.900 ;
        RECT 23.900 37.200 24.300 37.300 ;
        RECT 25.300 37.200 25.700 37.300 ;
        RECT 22.200 36.500 22.600 36.600 ;
        RECT 24.500 36.500 24.900 36.600 ;
        RECT 22.200 36.200 24.900 36.500 ;
        RECT 25.200 36.500 26.300 36.800 ;
        RECT 25.200 35.900 25.500 36.500 ;
        RECT 25.900 36.400 26.300 36.500 ;
        RECT 27.100 36.600 27.800 37.000 ;
        RECT 27.100 36.100 27.400 36.600 ;
        RECT 23.100 35.700 25.500 35.900 ;
        RECT 20.600 35.600 25.500 35.700 ;
        RECT 26.200 35.800 27.400 36.100 ;
        RECT 20.600 35.500 23.500 35.600 ;
        RECT 20.600 35.400 23.400 35.500 ;
        RECT 23.800 35.100 24.200 35.200 ;
        RECT 17.400 34.800 19.400 35.100 ;
        RECT 7.800 33.300 9.800 33.600 ;
        RECT 7.800 33.200 8.300 33.300 ;
        RECT 7.800 32.800 8.200 33.200 ;
        RECT 2.200 32.100 2.600 32.500 ;
        RECT 3.000 32.400 3.400 32.800 ;
        RECT 3.900 32.700 4.300 32.800 ;
        RECT 3.900 32.400 5.300 32.700 ;
        RECT 5.000 32.100 5.300 32.400 ;
        RECT 7.000 32.100 7.400 32.500 ;
        RECT 2.200 31.800 3.200 32.100 ;
        RECT 2.800 31.100 3.200 31.800 ;
        RECT 5.000 31.100 5.400 32.100 ;
        RECT 7.000 31.800 7.700 32.100 ;
        RECT 7.100 31.100 7.700 31.800 ;
        RECT 9.400 31.100 9.800 33.300 ;
        RECT 11.700 33.500 12.000 33.800 ;
        RECT 12.500 33.900 13.000 34.100 ;
        RECT 15.000 34.100 15.400 34.200 ;
        RECT 16.500 34.100 17.800 34.200 ;
        RECT 18.200 34.100 18.600 34.200 ;
        RECT 12.500 33.600 14.600 33.900 ;
        RECT 15.000 33.800 15.800 34.100 ;
        RECT 16.500 33.800 18.600 34.100 ;
        RECT 15.400 33.600 15.800 33.800 ;
        RECT 11.700 33.300 12.100 33.500 ;
        RECT 11.700 33.000 12.500 33.300 ;
        RECT 12.100 31.500 12.500 33.000 ;
        RECT 14.300 32.500 14.600 33.600 ;
        RECT 15.100 33.100 16.900 33.300 ;
        RECT 17.400 33.100 17.700 33.800 ;
        RECT 19.000 33.100 19.400 34.800 ;
        RECT 21.700 34.800 24.200 35.100 ;
        RECT 21.700 34.700 22.100 34.800 ;
        RECT 23.000 34.700 23.400 34.800 ;
        RECT 22.500 34.200 22.900 34.300 ;
        RECT 26.200 34.200 26.500 35.800 ;
        RECT 29.400 35.600 29.800 39.900 ;
        RECT 27.700 35.300 29.800 35.600 ;
        RECT 30.200 37.500 30.600 39.500 ;
        RECT 32.300 39.200 32.700 39.900 ;
        RECT 36.900 39.200 37.300 39.900 ;
        RECT 32.300 38.800 33.000 39.200 ;
        RECT 36.900 38.800 37.800 39.200 ;
        RECT 30.200 35.800 30.500 37.500 ;
        RECT 32.300 36.400 32.700 38.800 ;
        RECT 36.900 36.400 37.300 38.800 ;
        RECT 39.000 37.500 39.400 39.500 ;
        RECT 32.300 36.100 33.100 36.400 ;
        RECT 30.200 35.500 32.100 35.800 ;
        RECT 27.700 35.200 28.100 35.300 ;
        RECT 28.500 34.900 28.900 35.000 ;
        RECT 27.000 34.600 28.900 34.900 ;
        RECT 27.000 34.500 27.400 34.600 ;
        RECT 19.800 33.400 20.200 34.200 ;
        RECT 21.000 33.900 26.500 34.200 ;
        RECT 21.000 33.800 21.800 33.900 ;
        RECT 14.200 31.500 14.600 32.500 ;
        RECT 15.000 33.000 17.000 33.100 ;
        RECT 15.000 31.100 15.400 33.000 ;
        RECT 16.600 31.100 17.000 33.000 ;
        RECT 17.400 31.100 17.800 33.100 ;
        RECT 18.500 32.800 19.400 33.100 ;
        RECT 18.500 31.100 18.900 32.800 ;
        RECT 20.600 31.100 21.000 33.500 ;
        RECT 23.100 32.800 23.400 33.900 ;
        RECT 25.900 33.800 26.300 33.900 ;
        RECT 29.400 33.600 29.800 35.300 ;
        RECT 30.200 34.400 30.600 35.200 ;
        RECT 31.000 34.400 31.400 35.200 ;
        RECT 31.800 34.500 32.100 35.500 ;
        RECT 31.800 34.100 32.500 34.500 ;
        RECT 32.800 34.200 33.100 36.100 ;
        RECT 36.500 36.100 37.300 36.400 ;
        RECT 33.400 34.800 33.800 35.600 ;
        RECT 35.800 34.800 36.200 35.600 ;
        RECT 36.500 34.200 36.800 36.100 ;
        RECT 39.100 35.800 39.400 37.500 ;
        RECT 37.500 35.500 39.400 35.800 ;
        RECT 37.500 34.500 37.800 35.500 ;
        RECT 31.800 33.900 32.300 34.100 ;
        RECT 27.900 33.300 29.800 33.600 ;
        RECT 27.900 33.200 28.300 33.300 ;
        RECT 22.200 32.100 22.600 32.500 ;
        RECT 23.000 32.400 23.400 32.800 ;
        RECT 23.900 32.700 24.300 32.800 ;
        RECT 23.900 32.400 25.300 32.700 ;
        RECT 25.000 32.100 25.300 32.400 ;
        RECT 27.000 32.100 27.400 32.500 ;
        RECT 22.200 31.800 23.200 32.100 ;
        RECT 22.800 31.100 23.200 31.800 ;
        RECT 25.000 31.100 25.400 32.100 ;
        RECT 27.000 31.800 27.700 32.100 ;
        RECT 27.100 31.100 27.700 31.800 ;
        RECT 29.400 31.100 29.800 33.300 ;
        RECT 30.200 33.600 32.300 33.900 ;
        RECT 32.800 33.800 33.800 34.200 ;
        RECT 35.800 33.800 36.800 34.200 ;
        RECT 37.100 34.100 37.800 34.500 ;
        RECT 38.200 34.400 38.600 35.200 ;
        RECT 39.000 34.400 39.400 35.200 ;
        RECT 40.600 35.100 41.000 39.900 ;
        RECT 42.600 36.800 43.000 37.200 ;
        RECT 41.400 35.800 41.800 36.600 ;
        RECT 42.600 36.200 42.900 36.800 ;
        RECT 43.300 36.200 43.700 39.900 ;
        RECT 46.200 36.400 46.600 39.900 ;
        RECT 42.200 35.900 42.900 36.200 ;
        RECT 43.200 35.900 43.700 36.200 ;
        RECT 46.100 35.900 46.600 36.400 ;
        RECT 47.800 36.200 48.200 39.900 ;
        RECT 46.900 35.900 48.200 36.200 ;
        RECT 42.200 35.800 42.600 35.900 ;
        RECT 42.200 35.100 42.500 35.800 ;
        RECT 40.600 34.800 42.500 35.100 ;
        RECT 30.200 32.500 30.500 33.600 ;
        RECT 32.800 33.500 33.100 33.800 ;
        RECT 32.700 33.300 33.100 33.500 ;
        RECT 32.300 33.000 33.100 33.300 ;
        RECT 36.500 33.500 36.800 33.800 ;
        RECT 37.300 33.900 37.800 34.100 ;
        RECT 37.300 33.600 39.400 33.900 ;
        RECT 36.500 33.300 36.900 33.500 ;
        RECT 36.500 33.000 37.300 33.300 ;
        RECT 30.200 31.500 30.600 32.500 ;
        RECT 32.300 31.500 32.700 33.000 ;
        RECT 36.900 31.500 37.300 33.000 ;
        RECT 39.100 32.500 39.400 33.600 ;
        RECT 39.800 33.400 40.200 34.200 ;
        RECT 40.600 33.100 41.000 34.800 ;
        RECT 43.200 34.200 43.500 35.900 ;
        RECT 43.800 34.400 44.200 35.200 ;
        RECT 46.100 34.200 46.400 35.900 ;
        RECT 46.900 34.900 47.200 35.900 ;
        RECT 46.700 34.500 47.200 34.900 ;
        RECT 42.200 33.800 43.500 34.200 ;
        RECT 44.600 34.100 45.000 34.200 ;
        RECT 46.100 34.100 46.600 34.200 ;
        RECT 44.200 33.800 46.600 34.100 ;
        RECT 42.300 33.100 42.600 33.800 ;
        RECT 44.200 33.600 44.600 33.800 ;
        RECT 43.100 33.100 44.900 33.300 ;
        RECT 46.100 33.100 46.400 33.800 ;
        RECT 46.900 33.700 47.200 34.500 ;
        RECT 47.700 34.800 48.200 35.200 ;
        RECT 51.000 35.100 51.400 39.900 ;
        RECT 53.000 36.800 53.400 37.200 ;
        RECT 51.800 35.800 52.200 36.600 ;
        RECT 53.000 36.200 53.300 36.800 ;
        RECT 53.700 36.200 54.100 39.900 ;
        RECT 52.600 35.900 53.300 36.200 ;
        RECT 53.600 35.900 54.100 36.200 ;
        RECT 55.800 37.500 56.200 39.500 ;
        RECT 57.900 39.200 58.300 39.900 ;
        RECT 57.900 38.800 58.600 39.200 ;
        RECT 52.600 35.800 53.000 35.900 ;
        RECT 52.600 35.100 52.900 35.800 ;
        RECT 51.000 34.800 52.900 35.100 ;
        RECT 47.700 34.400 48.100 34.800 ;
        RECT 46.900 33.400 48.200 33.700 ;
        RECT 50.200 33.400 50.600 34.200 ;
        RECT 40.600 32.800 41.500 33.100 ;
        RECT 39.000 31.500 39.400 32.500 ;
        RECT 41.100 31.100 41.500 32.800 ;
        RECT 42.200 31.100 42.600 33.100 ;
        RECT 43.000 33.000 45.000 33.100 ;
        RECT 43.000 31.100 43.400 33.000 ;
        RECT 44.600 31.100 45.000 33.000 ;
        RECT 46.100 32.800 46.600 33.100 ;
        RECT 46.200 31.100 46.600 32.800 ;
        RECT 47.800 31.100 48.200 33.400 ;
        RECT 51.000 33.100 51.400 34.800 ;
        RECT 53.600 34.200 53.900 35.900 ;
        RECT 55.800 35.800 56.100 37.500 ;
        RECT 57.900 36.400 58.300 38.800 ;
        RECT 62.500 36.400 62.900 39.900 ;
        RECT 64.600 37.500 65.000 39.500 ;
        RECT 67.300 39.200 67.700 39.900 ;
        RECT 67.000 38.800 67.700 39.200 ;
        RECT 57.900 36.100 58.700 36.400 ;
        RECT 55.800 35.500 57.700 35.800 ;
        RECT 54.200 35.100 54.600 35.200 ;
        RECT 55.000 35.100 55.400 35.200 ;
        RECT 54.200 34.800 55.400 35.100 ;
        RECT 54.200 34.400 54.600 34.800 ;
        RECT 55.800 34.400 56.200 35.200 ;
        RECT 56.600 34.400 57.000 35.200 ;
        RECT 57.400 34.500 57.700 35.500 ;
        RECT 52.600 33.800 53.900 34.200 ;
        RECT 55.000 34.100 55.400 34.200 ;
        RECT 54.600 33.800 55.400 34.100 ;
        RECT 57.400 34.100 58.100 34.500 ;
        RECT 58.400 34.200 58.700 36.100 ;
        RECT 62.100 36.100 62.900 36.400 ;
        RECT 59.000 35.100 59.400 35.600 ;
        RECT 59.000 34.800 60.100 35.100 ;
        RECT 61.400 34.800 61.800 35.600 ;
        RECT 57.400 33.900 57.900 34.100 ;
        RECT 52.700 33.200 53.000 33.800 ;
        RECT 54.600 33.600 55.000 33.800 ;
        RECT 55.800 33.600 57.900 33.900 ;
        RECT 58.400 33.800 59.400 34.200 ;
        RECT 59.800 34.100 60.100 34.800 ;
        RECT 62.100 34.200 62.400 36.100 ;
        RECT 64.700 35.800 65.000 37.500 ;
        RECT 67.300 36.400 67.700 38.800 ;
        RECT 69.400 37.500 69.800 39.500 ;
        RECT 63.100 35.500 65.000 35.800 ;
        RECT 66.900 36.100 67.700 36.400 ;
        RECT 63.100 34.500 63.400 35.500 ;
        RECT 61.400 34.100 62.400 34.200 ;
        RECT 62.700 34.100 63.400 34.500 ;
        RECT 63.800 34.400 64.200 35.200 ;
        RECT 64.600 34.400 65.000 35.200 ;
        RECT 66.200 34.800 66.600 35.600 ;
        RECT 66.900 34.200 67.200 36.100 ;
        RECT 69.500 35.800 69.800 37.500 ;
        RECT 71.000 36.400 71.400 39.900 ;
        RECT 67.900 35.500 69.800 35.800 ;
        RECT 70.900 35.900 71.400 36.400 ;
        RECT 72.600 36.200 73.000 39.900 ;
        RECT 71.700 35.900 73.000 36.200 ;
        RECT 67.900 34.500 68.200 35.500 ;
        RECT 59.800 33.800 62.400 34.100 ;
        RECT 51.000 32.800 51.900 33.100 ;
        RECT 51.500 31.100 51.900 32.800 ;
        RECT 52.600 31.100 53.000 33.200 ;
        RECT 53.500 33.100 55.300 33.300 ;
        RECT 53.400 33.000 55.400 33.100 ;
        RECT 53.400 31.100 53.800 33.000 ;
        RECT 55.000 31.100 55.400 33.000 ;
        RECT 55.800 32.500 56.100 33.600 ;
        RECT 58.400 33.500 58.700 33.800 ;
        RECT 58.300 33.300 58.700 33.500 ;
        RECT 57.900 33.000 58.700 33.300 ;
        RECT 62.100 33.500 62.400 33.800 ;
        RECT 62.900 33.900 63.400 34.100 ;
        RECT 62.900 33.600 65.000 33.900 ;
        RECT 66.200 33.800 67.200 34.200 ;
        RECT 67.500 34.100 68.200 34.500 ;
        RECT 68.600 34.400 69.000 35.200 ;
        RECT 69.400 34.400 69.800 35.200 ;
        RECT 62.100 33.300 62.500 33.500 ;
        RECT 62.100 33.000 62.900 33.300 ;
        RECT 55.800 31.500 56.200 32.500 ;
        RECT 57.900 31.500 58.300 33.000 ;
        RECT 62.500 31.500 62.900 33.000 ;
        RECT 64.700 32.500 65.000 33.600 ;
        RECT 66.900 33.500 67.200 33.800 ;
        RECT 67.700 33.900 68.200 34.100 ;
        RECT 70.900 34.200 71.200 35.900 ;
        RECT 71.700 34.900 72.000 35.900 ;
        RECT 73.400 35.700 73.800 39.900 ;
        RECT 75.600 38.200 76.000 39.900 ;
        RECT 75.000 37.900 76.000 38.200 ;
        RECT 77.800 37.900 78.200 39.900 ;
        RECT 79.900 37.900 80.500 39.900 ;
        RECT 75.000 37.500 75.400 37.900 ;
        RECT 77.800 37.600 78.100 37.900 ;
        RECT 76.700 37.300 78.500 37.600 ;
        RECT 79.800 37.500 80.200 37.900 ;
        RECT 76.700 37.200 77.100 37.300 ;
        RECT 78.100 37.200 78.500 37.300 ;
        RECT 75.000 36.500 75.400 36.600 ;
        RECT 77.300 36.500 77.700 36.600 ;
        RECT 75.000 36.200 77.700 36.500 ;
        RECT 78.000 36.500 79.100 36.800 ;
        RECT 78.000 35.900 78.300 36.500 ;
        RECT 78.700 36.400 79.100 36.500 ;
        RECT 79.900 36.600 80.600 37.000 ;
        RECT 79.900 36.100 80.200 36.600 ;
        RECT 75.900 35.700 78.300 35.900 ;
        RECT 73.400 35.600 78.300 35.700 ;
        RECT 79.000 35.800 80.200 36.100 ;
        RECT 73.400 35.500 76.300 35.600 ;
        RECT 73.400 35.400 76.200 35.500 ;
        RECT 71.500 34.500 72.000 34.900 ;
        RECT 67.700 33.600 69.800 33.900 ;
        RECT 66.900 33.300 67.300 33.500 ;
        RECT 66.900 33.000 67.700 33.300 ;
        RECT 64.600 31.500 65.000 32.500 ;
        RECT 67.300 31.500 67.700 33.000 ;
        RECT 69.500 32.500 69.800 33.600 ;
        RECT 70.900 33.800 71.400 34.200 ;
        RECT 70.900 33.100 71.200 33.800 ;
        RECT 71.700 33.700 72.000 34.500 ;
        RECT 72.500 34.800 73.000 35.200 ;
        RECT 76.600 35.100 77.000 35.200 ;
        RECT 74.500 34.800 77.000 35.100 ;
        RECT 72.500 34.400 72.900 34.800 ;
        RECT 74.500 34.700 74.900 34.800 ;
        RECT 75.300 34.200 75.700 34.300 ;
        RECT 79.000 34.200 79.300 35.800 ;
        RECT 82.200 35.600 82.600 39.900 ;
        RECT 80.500 35.300 82.600 35.600 ;
        RECT 80.500 35.200 80.900 35.300 ;
        RECT 81.300 34.900 81.700 35.000 ;
        RECT 79.800 34.600 81.700 34.900 ;
        RECT 79.800 34.500 80.200 34.600 ;
        RECT 73.800 33.900 79.300 34.200 ;
        RECT 73.800 33.800 74.600 33.900 ;
        RECT 71.700 33.400 73.000 33.700 ;
        RECT 70.900 32.800 71.400 33.100 ;
        RECT 69.400 31.500 69.800 32.500 ;
        RECT 71.000 31.100 71.400 32.800 ;
        RECT 72.600 31.100 73.000 33.400 ;
        RECT 73.400 31.100 73.800 33.500 ;
        RECT 75.900 32.800 76.200 33.900 ;
        RECT 77.400 33.800 77.800 33.900 ;
        RECT 78.700 33.800 79.100 33.900 ;
        RECT 82.200 33.600 82.600 35.300 ;
        RECT 80.700 33.300 82.600 33.600 ;
        RECT 83.000 33.400 83.400 34.200 ;
        RECT 80.700 33.200 81.100 33.300 ;
        RECT 75.000 32.100 75.400 32.500 ;
        RECT 75.800 32.400 76.200 32.800 ;
        RECT 76.700 32.700 77.100 32.800 ;
        RECT 76.700 32.400 78.100 32.700 ;
        RECT 77.800 32.100 78.100 32.400 ;
        RECT 79.800 32.100 80.200 32.500 ;
        RECT 75.000 31.800 76.000 32.100 ;
        RECT 75.600 31.100 76.000 31.800 ;
        RECT 77.800 31.100 78.200 32.100 ;
        RECT 79.800 31.800 80.500 32.100 ;
        RECT 79.900 31.100 80.500 31.800 ;
        RECT 82.200 31.100 82.600 33.300 ;
        RECT 83.800 33.100 84.200 39.900 ;
        RECT 84.600 35.800 85.000 36.600 ;
        RECT 85.400 36.200 85.800 39.900 ;
        RECT 87.000 36.200 87.400 39.900 ;
        RECT 85.400 35.900 87.400 36.200 ;
        RECT 87.800 35.900 88.200 39.900 ;
        RECT 89.900 36.300 90.300 39.900 ;
        RECT 92.900 39.200 93.300 39.900 ;
        RECT 92.900 38.800 93.800 39.200 ;
        RECT 92.900 36.400 93.300 38.800 ;
        RECT 95.000 37.500 95.400 39.500 ;
        RECT 89.400 35.900 90.300 36.300 ;
        RECT 92.500 36.100 93.300 36.400 ;
        RECT 85.800 35.200 86.200 35.400 ;
        RECT 87.800 35.200 88.100 35.900 ;
        RECT 85.400 34.900 86.200 35.200 ;
        RECT 87.000 34.900 88.200 35.200 ;
        RECT 85.400 34.800 85.800 34.900 ;
        RECT 86.200 33.800 86.600 34.600 ;
        RECT 87.000 34.200 87.300 34.900 ;
        RECT 87.800 34.800 88.200 34.900 ;
        RECT 89.500 34.200 89.800 35.900 ;
        RECT 90.200 34.800 90.600 35.600 ;
        RECT 91.800 34.800 92.200 35.600 ;
        RECT 92.500 34.200 92.800 36.100 ;
        RECT 95.100 35.800 95.400 37.500 ;
        RECT 96.600 36.400 97.000 39.900 ;
        RECT 93.500 35.500 95.400 35.800 ;
        RECT 96.500 35.900 97.000 36.400 ;
        RECT 98.200 36.200 98.600 39.900 ;
        RECT 102.500 39.200 102.900 39.900 ;
        RECT 102.200 38.800 102.900 39.200 ;
        RECT 102.500 36.400 102.900 38.800 ;
        RECT 104.600 37.500 105.000 39.500 ;
        RECT 97.300 35.900 98.600 36.200 ;
        RECT 102.100 36.100 102.900 36.400 ;
        RECT 93.500 34.500 93.800 35.500 ;
        RECT 87.000 33.800 87.400 34.200 ;
        RECT 89.400 34.100 89.800 34.200 ;
        RECT 87.800 33.800 89.800 34.100 ;
        RECT 91.800 33.800 92.800 34.200 ;
        RECT 93.100 34.100 93.800 34.500 ;
        RECT 94.200 34.400 94.600 35.200 ;
        RECT 95.000 34.400 95.400 35.200 ;
        RECT 87.000 33.100 87.300 33.800 ;
        RECT 87.800 33.200 88.100 33.800 ;
        RECT 83.800 32.800 84.700 33.100 ;
        RECT 84.300 32.200 84.700 32.800 ;
        RECT 84.300 31.800 85.000 32.200 ;
        RECT 84.300 31.100 84.700 31.800 ;
        RECT 87.000 31.100 87.400 33.100 ;
        RECT 87.800 32.800 88.200 33.200 ;
        RECT 87.700 32.400 88.100 32.800 ;
        RECT 88.600 32.400 89.000 33.200 ;
        RECT 89.500 32.100 89.800 33.800 ;
        RECT 92.500 33.500 92.800 33.800 ;
        RECT 93.300 33.900 93.800 34.100 ;
        RECT 96.500 34.200 96.800 35.900 ;
        RECT 97.300 34.900 97.600 35.900 ;
        RECT 97.100 34.500 97.600 34.900 ;
        RECT 93.300 33.600 95.400 33.900 ;
        RECT 92.500 33.300 92.900 33.500 ;
        RECT 92.500 33.000 93.300 33.300 ;
        RECT 89.400 31.100 89.800 32.100 ;
        RECT 92.900 31.500 93.300 33.000 ;
        RECT 95.100 32.500 95.400 33.600 ;
        RECT 96.500 33.800 97.000 34.200 ;
        RECT 96.500 33.200 96.800 33.800 ;
        RECT 97.300 33.700 97.600 34.500 ;
        RECT 98.100 34.800 98.600 35.200 ;
        RECT 101.400 34.800 101.800 35.600 ;
        RECT 98.100 34.400 98.500 34.800 ;
        RECT 102.100 34.200 102.400 36.100 ;
        RECT 104.700 35.800 105.000 37.500 ;
        RECT 106.700 36.200 107.100 39.900 ;
        RECT 107.400 36.800 107.800 37.200 ;
        RECT 107.500 36.200 107.800 36.800 ;
        RECT 106.700 35.900 107.200 36.200 ;
        RECT 107.500 35.900 108.200 36.200 ;
        RECT 103.100 35.500 105.000 35.800 ;
        RECT 103.100 34.500 103.400 35.500 ;
        RECT 101.400 33.800 102.400 34.200 ;
        RECT 102.700 34.100 103.400 34.500 ;
        RECT 103.800 34.400 104.200 35.200 ;
        RECT 104.600 34.400 105.000 35.200 ;
        RECT 106.200 34.400 106.600 35.200 ;
        RECT 106.900 34.200 107.200 35.900 ;
        RECT 107.800 35.800 108.200 35.900 ;
        RECT 108.600 35.800 109.000 36.600 ;
        RECT 107.800 35.100 108.100 35.800 ;
        RECT 109.400 35.100 109.800 39.900 ;
        RECT 111.000 35.700 111.400 39.900 ;
        RECT 113.200 38.200 113.600 39.900 ;
        RECT 112.600 37.900 113.600 38.200 ;
        RECT 115.400 37.900 115.800 39.900 ;
        RECT 117.500 37.900 118.100 39.900 ;
        RECT 112.600 37.500 113.000 37.900 ;
        RECT 115.400 37.600 115.700 37.900 ;
        RECT 114.300 37.300 116.100 37.600 ;
        RECT 117.400 37.500 117.800 37.900 ;
        RECT 114.300 37.200 114.700 37.300 ;
        RECT 115.700 37.200 116.100 37.300 ;
        RECT 117.900 37.000 118.600 37.200 ;
        RECT 117.500 36.800 118.600 37.000 ;
        RECT 112.600 36.500 113.000 36.600 ;
        RECT 114.900 36.500 115.300 36.600 ;
        RECT 112.600 36.200 115.300 36.500 ;
        RECT 115.600 36.500 116.700 36.800 ;
        RECT 115.600 35.900 115.900 36.500 ;
        RECT 116.300 36.400 116.700 36.500 ;
        RECT 117.500 36.600 118.200 36.800 ;
        RECT 117.500 36.100 117.800 36.600 ;
        RECT 113.500 35.700 115.900 35.900 ;
        RECT 111.000 35.600 115.900 35.700 ;
        RECT 116.600 35.800 117.800 36.100 ;
        RECT 111.000 35.500 113.900 35.600 ;
        RECT 111.000 35.400 113.800 35.500 ;
        RECT 114.200 35.100 114.600 35.200 ;
        RECT 107.800 34.800 109.800 35.100 ;
        RECT 97.300 33.400 98.600 33.700 ;
        RECT 96.500 32.800 97.000 33.200 ;
        RECT 95.000 31.500 95.400 32.500 ;
        RECT 96.600 31.100 97.000 32.800 ;
        RECT 98.200 31.100 98.600 33.400 ;
        RECT 102.100 33.500 102.400 33.800 ;
        RECT 102.900 33.900 103.400 34.100 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 102.900 33.600 105.000 33.900 ;
        RECT 105.400 33.800 106.200 34.100 ;
        RECT 106.900 33.800 108.200 34.200 ;
        RECT 105.800 33.600 106.200 33.800 ;
        RECT 102.100 33.300 102.500 33.500 ;
        RECT 102.100 33.000 102.900 33.300 ;
        RECT 102.500 31.500 102.900 33.000 ;
        RECT 104.700 32.500 105.000 33.600 ;
        RECT 105.500 33.100 107.300 33.300 ;
        RECT 107.800 33.100 108.100 33.800 ;
        RECT 109.400 33.100 109.800 34.800 ;
        RECT 112.100 34.800 114.600 35.100 ;
        RECT 115.800 35.100 116.200 35.200 ;
        RECT 116.600 35.100 116.900 35.800 ;
        RECT 119.800 35.600 120.200 39.900 ;
        RECT 118.100 35.300 120.200 35.600 ;
        RECT 120.600 37.500 121.000 39.500 ;
        RECT 122.700 39.200 123.100 39.900 ;
        RECT 122.200 38.800 123.100 39.200 ;
        RECT 120.600 35.800 120.900 37.500 ;
        RECT 122.700 36.400 123.100 38.800 ;
        RECT 127.300 36.400 127.700 39.900 ;
        RECT 129.400 37.500 129.800 39.500 ;
        RECT 122.700 36.100 123.500 36.400 ;
        RECT 120.600 35.500 122.500 35.800 ;
        RECT 118.100 35.200 118.500 35.300 ;
        RECT 115.800 34.800 116.900 35.100 ;
        RECT 118.900 34.900 119.300 35.000 ;
        RECT 112.100 34.700 112.500 34.800 ;
        RECT 113.400 34.700 113.800 34.800 ;
        RECT 112.900 34.200 113.300 34.300 ;
        RECT 116.600 34.200 116.900 34.800 ;
        RECT 117.400 34.600 119.300 34.900 ;
        RECT 117.400 34.500 117.800 34.600 ;
        RECT 110.200 33.400 110.600 34.200 ;
        RECT 111.400 33.900 116.900 34.200 ;
        RECT 111.400 33.800 112.200 33.900 ;
        RECT 104.600 31.500 105.000 32.500 ;
        RECT 105.400 33.000 107.400 33.100 ;
        RECT 105.400 31.100 105.800 33.000 ;
        RECT 107.000 31.100 107.400 33.000 ;
        RECT 107.800 31.100 108.200 33.100 ;
        RECT 108.900 32.800 109.800 33.100 ;
        RECT 108.900 31.100 109.300 32.800 ;
        RECT 111.000 31.100 111.400 33.500 ;
        RECT 113.500 32.800 113.800 33.900 ;
        RECT 116.300 33.800 116.700 33.900 ;
        RECT 119.800 33.600 120.200 35.300 ;
        RECT 120.600 34.400 121.000 35.200 ;
        RECT 121.400 34.400 121.800 35.200 ;
        RECT 122.200 34.500 122.500 35.500 ;
        RECT 122.200 34.100 122.900 34.500 ;
        RECT 123.200 34.200 123.500 36.100 ;
        RECT 126.900 36.100 127.700 36.400 ;
        RECT 123.800 34.800 124.200 35.600 ;
        RECT 126.200 34.800 126.600 35.600 ;
        RECT 126.900 34.200 127.200 36.100 ;
        RECT 129.500 35.800 129.800 37.500 ;
        RECT 127.900 35.500 129.800 35.800 ;
        RECT 130.200 35.600 130.600 39.900 ;
        RECT 132.300 37.900 132.900 39.900 ;
        RECT 134.600 37.900 135.000 39.900 ;
        RECT 136.800 38.200 137.200 39.900 ;
        RECT 136.800 37.900 137.800 38.200 ;
        RECT 132.600 37.500 133.000 37.900 ;
        RECT 134.700 37.600 135.000 37.900 ;
        RECT 134.300 37.300 136.100 37.600 ;
        RECT 137.400 37.500 137.800 37.900 ;
        RECT 134.300 37.200 134.700 37.300 ;
        RECT 135.700 37.200 136.100 37.300 ;
        RECT 132.200 36.600 132.900 37.000 ;
        RECT 132.600 36.100 132.900 36.600 ;
        RECT 133.700 36.500 134.800 36.800 ;
        RECT 133.700 36.400 134.100 36.500 ;
        RECT 132.600 35.800 133.800 36.100 ;
        RECT 127.900 34.500 128.200 35.500 ;
        RECT 130.200 35.300 132.300 35.600 ;
        RECT 122.200 33.900 122.700 34.100 ;
        RECT 118.300 33.300 120.200 33.600 ;
        RECT 118.300 33.200 118.700 33.300 ;
        RECT 112.600 32.100 113.000 32.500 ;
        RECT 113.400 32.400 113.800 32.800 ;
        RECT 114.300 32.700 114.700 32.800 ;
        RECT 114.300 32.400 115.700 32.700 ;
        RECT 115.400 32.100 115.700 32.400 ;
        RECT 117.400 32.100 117.800 32.500 ;
        RECT 112.600 31.800 113.600 32.100 ;
        RECT 113.200 31.100 113.600 31.800 ;
        RECT 115.400 31.100 115.800 32.100 ;
        RECT 117.400 31.800 118.100 32.100 ;
        RECT 117.500 31.100 118.100 31.800 ;
        RECT 119.800 31.100 120.200 33.300 ;
        RECT 120.600 33.600 122.700 33.900 ;
        RECT 123.200 33.800 124.200 34.200 ;
        RECT 126.200 33.800 127.200 34.200 ;
        RECT 127.500 34.100 128.200 34.500 ;
        RECT 128.600 34.400 129.000 35.200 ;
        RECT 129.400 34.400 129.800 35.200 ;
        RECT 120.600 32.500 120.900 33.600 ;
        RECT 123.200 33.500 123.500 33.800 ;
        RECT 123.100 33.300 123.500 33.500 ;
        RECT 122.700 33.000 123.500 33.300 ;
        RECT 126.900 33.500 127.200 33.800 ;
        RECT 127.700 33.900 128.200 34.100 ;
        RECT 127.700 33.600 129.800 33.900 ;
        RECT 126.900 33.300 127.300 33.500 ;
        RECT 126.900 33.000 127.700 33.300 ;
        RECT 120.600 31.500 121.000 32.500 ;
        RECT 122.700 31.500 123.100 33.000 ;
        RECT 127.300 32.200 127.700 33.000 ;
        RECT 129.500 32.500 129.800 33.600 ;
        RECT 127.000 31.800 127.700 32.200 ;
        RECT 127.300 31.500 127.700 31.800 ;
        RECT 129.400 31.500 129.800 32.500 ;
        RECT 130.200 33.600 130.600 35.300 ;
        RECT 131.900 35.200 132.300 35.300 ;
        RECT 131.100 34.900 131.500 35.000 ;
        RECT 131.100 34.600 133.000 34.900 ;
        RECT 132.600 34.500 133.000 34.600 ;
        RECT 133.500 34.200 133.800 35.800 ;
        RECT 134.500 35.900 134.800 36.500 ;
        RECT 135.100 36.500 135.500 36.600 ;
        RECT 137.400 36.500 137.800 36.600 ;
        RECT 135.100 36.200 137.800 36.500 ;
        RECT 134.500 35.700 136.900 35.900 ;
        RECT 139.000 35.700 139.400 39.900 ;
        RECT 134.500 35.600 139.400 35.700 ;
        RECT 136.500 35.500 139.400 35.600 ;
        RECT 136.600 35.400 139.400 35.500 ;
        RECT 135.800 35.100 136.200 35.200 ;
        RECT 135.800 34.800 138.300 35.100 ;
        RECT 136.600 34.700 137.000 34.800 ;
        RECT 137.900 34.700 138.300 34.800 ;
        RECT 137.100 34.200 137.500 34.300 ;
        RECT 133.500 33.900 139.000 34.200 ;
        RECT 133.700 33.800 134.100 33.900 ;
        RECT 130.200 33.300 132.100 33.600 ;
        RECT 130.200 31.100 130.600 33.300 ;
        RECT 131.700 33.200 132.100 33.300 ;
        RECT 136.600 33.200 136.900 33.900 ;
        RECT 138.200 33.800 139.000 33.900 ;
        RECT 135.700 32.700 136.100 32.800 ;
        RECT 132.600 32.100 133.000 32.500 ;
        RECT 134.700 32.400 136.100 32.700 ;
        RECT 136.600 32.400 137.000 33.200 ;
        RECT 134.700 32.100 135.000 32.400 ;
        RECT 137.400 32.100 137.800 32.500 ;
        RECT 132.300 31.800 133.000 32.100 ;
        RECT 132.300 31.100 132.900 31.800 ;
        RECT 134.600 31.100 135.000 32.100 ;
        RECT 136.800 31.800 137.800 32.100 ;
        RECT 136.800 31.100 137.200 31.800 ;
        RECT 139.000 31.100 139.400 33.500 ;
        RECT 139.800 33.400 140.200 34.200 ;
        RECT 140.600 33.100 141.000 39.900 ;
        RECT 141.400 35.800 141.800 36.600 ;
        RECT 140.600 32.800 141.500 33.100 ;
        RECT 141.100 32.200 141.500 32.800 ;
        RECT 140.600 31.800 141.500 32.200 ;
        RECT 141.100 31.100 141.500 31.800 ;
        RECT 143.000 31.100 143.400 39.900 ;
        RECT 146.500 39.200 146.900 39.900 ;
        RECT 146.200 38.800 146.900 39.200 ;
        RECT 146.500 36.400 146.900 38.800 ;
        RECT 148.600 37.500 149.000 39.500 ;
        RECT 146.100 36.100 146.900 36.400 ;
        RECT 145.400 34.800 145.800 35.600 ;
        RECT 146.100 34.200 146.400 36.100 ;
        RECT 148.700 35.800 149.000 37.500 ;
        RECT 147.100 35.500 149.000 35.800 ;
        RECT 151.000 35.600 151.400 39.900 ;
        RECT 153.100 37.900 153.700 39.900 ;
        RECT 155.400 37.900 155.800 39.900 ;
        RECT 157.600 38.200 158.000 39.900 ;
        RECT 157.600 37.900 158.600 38.200 ;
        RECT 153.400 37.500 153.800 37.900 ;
        RECT 155.500 37.600 155.800 37.900 ;
        RECT 155.100 37.300 156.900 37.600 ;
        RECT 158.200 37.500 158.600 37.900 ;
        RECT 155.100 37.200 155.500 37.300 ;
        RECT 156.500 37.200 156.900 37.300 ;
        RECT 153.000 36.600 153.700 37.000 ;
        RECT 153.400 36.100 153.700 36.600 ;
        RECT 154.500 36.500 155.600 36.800 ;
        RECT 154.500 36.400 154.900 36.500 ;
        RECT 153.400 35.800 154.600 36.100 ;
        RECT 147.100 34.500 147.400 35.500 ;
        RECT 151.000 35.300 153.100 35.600 ;
        RECT 145.400 33.800 146.400 34.200 ;
        RECT 146.700 34.100 147.400 34.500 ;
        RECT 147.800 34.400 148.200 35.200 ;
        RECT 148.600 34.400 149.000 35.200 ;
        RECT 146.100 33.500 146.400 33.800 ;
        RECT 146.900 33.900 147.400 34.100 ;
        RECT 146.900 33.600 149.000 33.900 ;
        RECT 146.100 33.300 146.500 33.500 ;
        RECT 146.100 33.000 146.900 33.300 ;
        RECT 146.500 31.500 146.900 33.000 ;
        RECT 148.700 32.500 149.000 33.600 ;
        RECT 148.600 31.500 149.000 32.500 ;
        RECT 151.000 33.600 151.400 35.300 ;
        RECT 152.700 35.200 153.100 35.300 ;
        RECT 151.900 34.900 152.300 35.000 ;
        RECT 151.900 34.600 153.800 34.900 ;
        RECT 153.400 34.500 153.800 34.600 ;
        RECT 154.300 34.200 154.600 35.800 ;
        RECT 155.300 35.900 155.600 36.500 ;
        RECT 155.900 36.500 156.300 36.600 ;
        RECT 158.200 36.500 158.600 36.600 ;
        RECT 155.900 36.200 158.600 36.500 ;
        RECT 155.300 35.700 157.700 35.900 ;
        RECT 159.800 35.700 160.200 39.900 ;
        RECT 161.400 36.400 161.800 39.900 ;
        RECT 155.300 35.600 160.200 35.700 ;
        RECT 157.300 35.500 160.200 35.600 ;
        RECT 157.400 35.400 160.200 35.500 ;
        RECT 161.300 35.900 161.800 36.400 ;
        RECT 163.000 36.200 163.400 39.900 ;
        RECT 162.100 35.900 163.400 36.200 ;
        RECT 163.800 36.200 164.200 39.900 ;
        RECT 165.400 36.400 165.800 39.900 ;
        RECT 163.800 35.900 165.100 36.200 ;
        RECT 165.400 35.900 165.900 36.400 ;
        RECT 156.600 35.100 157.000 35.200 ;
        RECT 156.600 34.800 159.100 35.100 ;
        RECT 157.400 34.700 157.800 34.800 ;
        RECT 158.700 34.700 159.100 34.800 ;
        RECT 157.900 34.200 158.300 34.300 ;
        RECT 161.300 34.200 161.600 35.900 ;
        RECT 162.100 34.900 162.400 35.900 ;
        RECT 161.900 34.500 162.400 34.900 ;
        RECT 154.300 33.900 159.800 34.200 ;
        RECT 154.500 33.800 154.900 33.900 ;
        RECT 156.600 33.800 157.000 33.900 ;
        RECT 151.000 33.300 152.900 33.600 ;
        RECT 151.000 31.100 151.400 33.300 ;
        RECT 152.500 33.200 152.900 33.300 ;
        RECT 157.400 33.200 157.700 33.900 ;
        RECT 159.000 33.800 159.800 33.900 ;
        RECT 161.300 33.800 161.800 34.200 ;
        RECT 156.500 32.700 156.900 32.800 ;
        RECT 153.400 32.100 153.800 32.500 ;
        RECT 155.500 32.400 156.900 32.700 ;
        RECT 157.400 32.400 157.800 33.200 ;
        RECT 155.500 32.100 155.800 32.400 ;
        RECT 158.200 32.100 158.600 32.500 ;
        RECT 153.100 31.800 153.800 32.100 ;
        RECT 153.100 31.100 153.700 31.800 ;
        RECT 155.400 31.100 155.800 32.100 ;
        RECT 157.600 31.800 158.600 32.100 ;
        RECT 157.600 31.100 158.000 31.800 ;
        RECT 159.800 31.100 160.200 33.500 ;
        RECT 161.300 33.100 161.600 33.800 ;
        RECT 162.100 33.700 162.400 34.500 ;
        RECT 164.800 34.900 165.100 35.900 ;
        RECT 164.800 34.500 165.300 34.900 ;
        RECT 164.800 33.700 165.100 34.500 ;
        RECT 165.600 34.200 165.900 35.900 ;
        RECT 167.000 35.800 167.400 36.600 ;
        RECT 165.400 34.100 165.900 34.200 ;
        RECT 167.000 34.100 167.400 34.200 ;
        RECT 165.400 33.800 167.400 34.100 ;
        RECT 162.100 33.400 163.400 33.700 ;
        RECT 161.300 32.800 161.800 33.100 ;
        RECT 161.400 31.100 161.800 32.800 ;
        RECT 163.000 31.100 163.400 33.400 ;
        RECT 163.800 33.400 165.100 33.700 ;
        RECT 163.800 31.100 164.200 33.400 ;
        RECT 165.600 33.100 165.900 33.800 ;
        RECT 167.800 33.100 168.200 39.900 ;
        RECT 169.400 37.500 169.800 39.500 ;
        RECT 171.500 39.200 171.900 39.900 ;
        RECT 171.000 38.800 171.900 39.200 ;
        RECT 169.400 35.800 169.700 37.500 ;
        RECT 171.500 36.400 171.900 38.800 ;
        RECT 171.500 36.100 172.300 36.400 ;
        RECT 169.400 35.500 171.300 35.800 ;
        RECT 168.600 34.800 169.000 35.200 ;
        RECT 168.600 34.200 168.900 34.800 ;
        RECT 169.400 34.400 169.800 35.200 ;
        RECT 170.200 34.400 170.600 35.200 ;
        RECT 171.000 34.500 171.300 35.500 ;
        RECT 168.600 33.400 169.000 34.200 ;
        RECT 171.000 34.100 171.700 34.500 ;
        RECT 172.000 34.200 172.300 36.100 ;
        RECT 174.200 36.200 174.600 39.900 ;
        RECT 175.800 36.400 176.200 39.900 ;
        RECT 177.400 37.500 177.800 39.500 ;
        RECT 179.500 39.200 179.900 39.900 ;
        RECT 179.500 38.800 180.200 39.200 ;
        RECT 174.200 35.900 175.500 36.200 ;
        RECT 175.800 35.900 176.300 36.400 ;
        RECT 172.600 35.100 173.000 35.600 ;
        RECT 173.400 35.100 173.800 35.200 ;
        RECT 172.600 34.800 173.800 35.100 ;
        RECT 175.200 34.900 175.500 35.900 ;
        RECT 175.200 34.500 175.700 34.900 ;
        RECT 171.000 33.900 171.500 34.100 ;
        RECT 169.400 33.600 171.500 33.900 ;
        RECT 172.000 33.800 173.000 34.200 ;
        RECT 165.400 32.800 165.900 33.100 ;
        RECT 167.300 32.800 168.200 33.100 ;
        RECT 165.400 31.100 165.800 32.800 ;
        RECT 167.300 32.200 167.700 32.800 ;
        RECT 169.400 32.500 169.700 33.600 ;
        RECT 172.000 33.500 172.300 33.800 ;
        RECT 175.200 33.700 175.500 34.500 ;
        RECT 176.000 34.200 176.300 35.900 ;
        RECT 177.400 35.800 177.700 37.500 ;
        RECT 179.500 36.400 179.900 38.800 ;
        RECT 179.500 36.100 180.300 36.400 ;
        RECT 177.400 35.500 179.300 35.800 ;
        RECT 177.400 34.400 177.800 35.200 ;
        RECT 178.200 34.400 178.600 35.200 ;
        RECT 179.000 34.500 179.300 35.500 ;
        RECT 175.800 33.800 176.300 34.200 ;
        RECT 179.000 34.100 179.700 34.500 ;
        RECT 180.000 34.200 180.300 36.100 ;
        RECT 180.600 35.100 181.000 35.600 ;
        RECT 183.000 35.100 183.400 39.900 ;
        RECT 185.000 36.800 185.400 37.200 ;
        RECT 183.800 35.800 184.200 36.600 ;
        RECT 185.000 36.200 185.300 36.800 ;
        RECT 185.700 36.200 186.100 39.900 ;
        RECT 184.600 35.900 185.300 36.200 ;
        RECT 184.600 35.800 185.000 35.900 ;
        RECT 185.600 35.800 186.600 36.200 ;
        RECT 184.600 35.100 184.900 35.800 ;
        RECT 180.600 34.800 181.700 35.100 ;
        RECT 179.000 33.900 179.500 34.100 ;
        RECT 171.900 33.300 172.300 33.500 ;
        RECT 171.500 33.000 172.300 33.300 ;
        RECT 174.200 33.400 175.500 33.700 ;
        RECT 167.300 31.800 168.200 32.200 ;
        RECT 167.300 31.100 167.700 31.800 ;
        RECT 169.400 31.500 169.800 32.500 ;
        RECT 171.500 31.500 171.900 33.000 ;
        RECT 174.200 31.100 174.600 33.400 ;
        RECT 176.000 33.100 176.300 33.800 ;
        RECT 175.800 32.800 176.300 33.100 ;
        RECT 177.400 33.600 179.500 33.900 ;
        RECT 180.000 33.800 181.000 34.200 ;
        RECT 181.400 34.100 181.700 34.800 ;
        RECT 183.000 34.800 184.900 35.100 ;
        RECT 182.200 34.100 182.600 34.200 ;
        RECT 181.400 33.800 182.600 34.100 ;
        RECT 175.800 31.100 176.200 32.800 ;
        RECT 177.400 32.500 177.700 33.600 ;
        RECT 180.000 33.500 180.300 33.800 ;
        RECT 179.900 33.300 180.300 33.500 ;
        RECT 182.200 33.400 182.600 33.800 ;
        RECT 179.500 33.000 180.300 33.300 ;
        RECT 183.000 33.100 183.400 34.800 ;
        RECT 185.600 34.200 185.900 35.800 ;
        RECT 187.800 35.600 188.200 39.900 ;
        RECT 189.900 37.900 190.500 39.900 ;
        RECT 192.200 37.900 192.600 39.900 ;
        RECT 194.400 38.200 194.800 39.900 ;
        RECT 194.400 37.900 195.400 38.200 ;
        RECT 190.200 37.500 190.600 37.900 ;
        RECT 192.300 37.600 192.600 37.900 ;
        RECT 191.900 37.300 193.700 37.600 ;
        RECT 195.000 37.500 195.400 37.900 ;
        RECT 191.900 37.200 192.300 37.300 ;
        RECT 193.300 37.200 193.700 37.300 ;
        RECT 189.800 36.600 190.500 37.000 ;
        RECT 190.200 36.100 190.500 36.600 ;
        RECT 191.300 36.500 192.400 36.800 ;
        RECT 191.300 36.400 191.700 36.500 ;
        RECT 190.200 35.800 191.400 36.100 ;
        RECT 187.800 35.300 189.900 35.600 ;
        RECT 186.200 34.400 186.600 35.200 ;
        RECT 184.600 33.800 185.900 34.200 ;
        RECT 187.000 34.100 187.400 34.200 ;
        RECT 186.600 33.800 187.400 34.100 ;
        RECT 184.700 33.100 185.000 33.800 ;
        RECT 186.600 33.600 187.000 33.800 ;
        RECT 187.800 33.600 188.200 35.300 ;
        RECT 189.500 35.200 189.900 35.300 ;
        RECT 191.100 35.100 191.400 35.800 ;
        RECT 192.100 35.900 192.400 36.500 ;
        RECT 192.700 36.500 193.100 36.600 ;
        RECT 195.000 36.500 195.400 36.600 ;
        RECT 192.700 36.200 195.400 36.500 ;
        RECT 192.100 35.700 194.500 35.900 ;
        RECT 196.600 35.700 197.000 39.900 ;
        RECT 192.100 35.600 197.000 35.700 ;
        RECT 194.100 35.500 197.000 35.600 ;
        RECT 197.400 37.500 197.800 39.500 ;
        RECT 199.500 39.200 199.900 39.900 ;
        RECT 199.000 38.800 199.900 39.200 ;
        RECT 197.400 35.800 197.700 37.500 ;
        RECT 199.500 36.400 199.900 38.800 ;
        RECT 199.500 36.100 200.300 36.400 ;
        RECT 197.400 35.500 199.300 35.800 ;
        RECT 194.200 35.400 197.000 35.500 ;
        RECT 191.800 35.100 192.200 35.200 ;
        RECT 188.700 34.900 189.100 35.000 ;
        RECT 188.700 34.600 190.600 34.900 ;
        RECT 191.000 34.800 192.200 35.100 ;
        RECT 193.400 35.100 193.800 35.200 ;
        RECT 193.400 34.800 195.900 35.100 ;
        RECT 190.200 34.500 190.600 34.600 ;
        RECT 191.100 34.200 191.400 34.800 ;
        RECT 195.500 34.700 195.900 34.800 ;
        RECT 197.400 34.400 197.800 35.200 ;
        RECT 198.200 34.400 198.600 35.200 ;
        RECT 199.000 34.500 199.300 35.500 ;
        RECT 194.700 34.200 195.100 34.300 ;
        RECT 191.100 33.900 196.600 34.200 ;
        RECT 199.000 34.100 199.700 34.500 ;
        RECT 200.000 34.200 200.300 36.100 ;
        RECT 203.800 35.600 204.200 39.900 ;
        RECT 205.900 37.900 206.500 39.900 ;
        RECT 208.200 37.900 208.600 39.900 ;
        RECT 210.400 38.200 210.800 39.900 ;
        RECT 210.400 37.900 211.400 38.200 ;
        RECT 206.200 37.500 206.600 37.900 ;
        RECT 208.300 37.600 208.600 37.900 ;
        RECT 207.900 37.300 209.700 37.600 ;
        RECT 211.000 37.500 211.400 37.900 ;
        RECT 207.900 37.200 208.300 37.300 ;
        RECT 209.300 37.200 209.700 37.300 ;
        RECT 205.800 36.600 206.500 37.000 ;
        RECT 206.200 36.100 206.500 36.600 ;
        RECT 207.300 36.500 208.400 36.800 ;
        RECT 207.300 36.400 207.700 36.500 ;
        RECT 206.200 35.800 207.400 36.100 ;
        RECT 200.600 34.800 201.000 35.600 ;
        RECT 203.800 35.300 205.900 35.600 ;
        RECT 199.000 33.900 199.500 34.100 ;
        RECT 191.300 33.800 191.700 33.900 ;
        RECT 187.800 33.300 189.700 33.600 ;
        RECT 185.500 33.100 187.300 33.300 ;
        RECT 177.400 31.500 177.800 32.500 ;
        RECT 179.500 31.500 179.900 33.000 ;
        RECT 183.000 32.800 183.900 33.100 ;
        RECT 183.500 31.100 183.900 32.800 ;
        RECT 184.600 31.100 185.000 33.100 ;
        RECT 185.400 33.000 187.400 33.100 ;
        RECT 185.400 31.100 185.800 33.000 ;
        RECT 187.000 31.100 187.400 33.000 ;
        RECT 187.800 31.100 188.200 33.300 ;
        RECT 189.300 33.200 189.700 33.300 ;
        RECT 194.200 32.800 194.500 33.900 ;
        RECT 195.800 33.800 196.600 33.900 ;
        RECT 197.400 33.600 199.500 33.900 ;
        RECT 200.000 33.800 201.000 34.200 ;
        RECT 193.300 32.700 193.700 32.800 ;
        RECT 190.200 32.100 190.600 32.500 ;
        RECT 192.300 32.400 193.700 32.700 ;
        RECT 194.200 32.400 194.600 32.800 ;
        RECT 192.300 32.100 192.600 32.400 ;
        RECT 195.000 32.100 195.400 32.500 ;
        RECT 189.900 31.800 190.600 32.100 ;
        RECT 189.900 31.100 190.500 31.800 ;
        RECT 192.200 31.100 192.600 32.100 ;
        RECT 194.400 31.800 195.400 32.100 ;
        RECT 194.400 31.100 194.800 31.800 ;
        RECT 196.600 31.100 197.000 33.500 ;
        RECT 197.400 32.500 197.700 33.600 ;
        RECT 200.000 33.500 200.300 33.800 ;
        RECT 199.900 33.300 200.300 33.500 ;
        RECT 199.500 33.000 200.300 33.300 ;
        RECT 203.800 33.600 204.200 35.300 ;
        RECT 205.500 35.200 205.900 35.300 ;
        RECT 207.100 35.200 207.400 35.800 ;
        RECT 208.100 35.900 208.400 36.500 ;
        RECT 208.700 36.500 209.100 36.600 ;
        RECT 211.000 36.500 211.400 36.600 ;
        RECT 208.700 36.200 211.400 36.500 ;
        RECT 208.100 35.700 210.500 35.900 ;
        RECT 212.600 35.700 213.000 39.900 ;
        RECT 213.400 35.800 213.800 36.600 ;
        RECT 208.100 35.600 213.000 35.700 ;
        RECT 210.100 35.500 213.000 35.600 ;
        RECT 210.200 35.400 213.000 35.500 ;
        RECT 204.700 34.900 205.100 35.000 ;
        RECT 204.700 34.600 206.600 34.900 ;
        RECT 207.000 34.800 207.400 35.200 ;
        RECT 208.600 35.100 209.000 35.200 ;
        RECT 209.400 35.100 209.800 35.200 ;
        RECT 208.600 34.800 211.900 35.100 ;
        RECT 206.200 34.500 206.600 34.600 ;
        RECT 207.100 34.200 207.400 34.800 ;
        RECT 211.500 34.700 211.900 34.800 ;
        RECT 210.700 34.200 211.100 34.300 ;
        RECT 207.100 33.900 212.600 34.200 ;
        RECT 207.300 33.800 207.700 33.900 ;
        RECT 203.800 33.300 205.700 33.600 ;
        RECT 197.400 31.500 197.800 32.500 ;
        RECT 199.500 31.500 199.900 33.000 ;
        RECT 203.000 32.100 203.400 32.200 ;
        RECT 203.800 32.100 204.200 33.300 ;
        RECT 205.300 33.200 205.700 33.300 ;
        RECT 210.200 32.800 210.500 33.900 ;
        RECT 211.800 33.800 212.600 33.900 ;
        RECT 209.300 32.700 209.700 32.800 ;
        RECT 206.200 32.100 206.600 32.500 ;
        RECT 208.300 32.400 209.700 32.700 ;
        RECT 210.200 32.400 210.600 32.800 ;
        RECT 208.300 32.100 208.600 32.400 ;
        RECT 211.000 32.100 211.400 32.500 ;
        RECT 203.000 31.800 204.200 32.100 ;
        RECT 203.800 31.100 204.200 31.800 ;
        RECT 205.900 31.800 206.600 32.100 ;
        RECT 205.900 31.100 206.500 31.800 ;
        RECT 208.200 31.100 208.600 32.100 ;
        RECT 210.400 31.800 211.400 32.100 ;
        RECT 210.400 31.100 210.800 31.800 ;
        RECT 212.600 31.100 213.000 33.500 ;
        RECT 214.200 33.100 214.600 39.900 ;
        RECT 215.800 37.500 216.200 39.500 ;
        RECT 215.800 35.800 216.100 37.500 ;
        RECT 217.900 36.400 218.300 39.900 ;
        RECT 217.900 36.100 218.700 36.400 ;
        RECT 215.800 35.500 217.700 35.800 ;
        RECT 215.800 34.400 216.200 35.200 ;
        RECT 216.600 34.400 217.000 35.200 ;
        RECT 217.400 34.500 217.700 35.500 ;
        RECT 215.000 33.400 215.400 34.200 ;
        RECT 217.400 34.100 218.100 34.500 ;
        RECT 218.400 34.200 218.700 36.100 ;
        RECT 221.900 36.200 222.300 39.900 ;
        RECT 222.600 36.800 223.000 37.200 ;
        RECT 222.700 36.200 223.000 36.800 ;
        RECT 221.900 35.900 222.400 36.200 ;
        RECT 222.700 35.900 223.400 36.200 ;
        RECT 219.000 35.100 219.400 35.600 ;
        RECT 219.800 35.100 220.200 35.200 ;
        RECT 219.000 34.800 220.200 35.100 ;
        RECT 221.400 34.400 221.800 35.200 ;
        RECT 222.100 34.200 222.400 35.900 ;
        RECT 223.000 35.800 223.400 35.900 ;
        RECT 223.800 35.800 224.200 36.600 ;
        RECT 223.000 35.100 223.300 35.800 ;
        RECT 224.600 35.100 225.000 39.900 ;
        RECT 228.100 36.400 228.500 39.900 ;
        RECT 230.200 37.500 230.600 39.500 ;
        RECT 227.700 36.100 228.500 36.400 ;
        RECT 227.000 35.100 227.400 35.600 ;
        RECT 223.000 34.800 225.000 35.100 ;
        RECT 217.400 33.900 217.900 34.100 ;
        RECT 215.800 33.600 217.900 33.900 ;
        RECT 218.400 33.800 219.400 34.200 ;
        RECT 220.600 34.100 221.000 34.200 ;
        RECT 220.600 33.800 221.400 34.100 ;
        RECT 222.100 33.800 223.400 34.200 ;
        RECT 213.700 32.800 214.600 33.100 ;
        RECT 213.700 32.200 214.100 32.800 ;
        RECT 215.800 32.500 216.100 33.600 ;
        RECT 218.400 33.500 218.700 33.800 ;
        RECT 221.000 33.600 221.400 33.800 ;
        RECT 218.300 33.300 218.700 33.500 ;
        RECT 217.900 33.000 218.700 33.300 ;
        RECT 220.700 33.100 222.500 33.300 ;
        RECT 223.000 33.100 223.300 33.800 ;
        RECT 224.600 33.100 225.000 34.800 ;
        RECT 226.200 34.800 227.400 35.100 ;
        RECT 226.200 34.200 226.500 34.800 ;
        RECT 227.700 34.200 228.000 36.100 ;
        RECT 230.300 35.800 230.600 37.500 ;
        RECT 232.300 36.300 232.700 39.900 ;
        RECT 231.800 35.900 232.700 36.300 ;
        RECT 233.400 35.900 233.800 39.900 ;
        RECT 234.200 36.200 234.600 39.900 ;
        RECT 235.800 36.200 236.200 39.900 ;
        RECT 234.200 35.900 236.200 36.200 ;
        RECT 237.900 36.200 238.300 39.900 ;
        RECT 238.600 36.800 239.000 37.200 ;
        RECT 238.700 36.200 239.000 36.800 ;
        RECT 237.900 35.900 238.400 36.200 ;
        RECT 238.700 35.900 239.400 36.200 ;
        RECT 228.700 35.500 230.600 35.800 ;
        RECT 228.700 34.500 229.000 35.500 ;
        RECT 225.400 34.100 225.800 34.200 ;
        RECT 226.200 34.100 226.600 34.200 ;
        RECT 225.400 33.800 226.600 34.100 ;
        RECT 227.000 33.800 228.000 34.200 ;
        RECT 228.300 34.100 229.000 34.500 ;
        RECT 229.400 34.400 229.800 35.200 ;
        RECT 230.200 34.400 230.600 35.200 ;
        RECT 231.900 34.200 232.200 35.900 ;
        RECT 232.600 34.800 233.000 35.600 ;
        RECT 233.500 35.200 233.800 35.900 ;
        RECT 235.400 35.200 235.800 35.400 ;
        RECT 233.400 34.900 234.600 35.200 ;
        RECT 235.400 34.900 236.200 35.200 ;
        RECT 233.400 34.800 233.800 34.900 ;
        RECT 225.400 33.400 225.800 33.800 ;
        RECT 227.700 33.500 228.000 33.800 ;
        RECT 228.500 33.900 229.000 34.100 ;
        RECT 228.500 33.600 230.600 33.900 ;
        RECT 231.800 33.800 232.200 34.200 ;
        RECT 220.600 33.000 222.600 33.100 ;
        RECT 213.700 31.800 214.600 32.200 ;
        RECT 213.700 31.100 214.100 31.800 ;
        RECT 215.800 31.500 216.200 32.500 ;
        RECT 217.900 31.500 218.300 33.000 ;
        RECT 220.600 31.100 221.000 33.000 ;
        RECT 222.200 31.100 222.600 33.000 ;
        RECT 223.000 31.100 223.400 33.100 ;
        RECT 224.100 32.800 225.000 33.100 ;
        RECT 227.700 33.300 228.100 33.500 ;
        RECT 227.700 33.000 228.500 33.300 ;
        RECT 224.100 31.100 224.500 32.800 ;
        RECT 228.100 31.500 228.500 33.000 ;
        RECT 230.300 32.500 230.600 33.600 ;
        RECT 230.200 31.500 230.600 32.500 ;
        RECT 231.000 32.400 231.400 33.200 ;
        RECT 231.900 33.100 232.200 33.800 ;
        RECT 233.400 33.100 233.800 33.200 ;
        RECT 234.300 33.100 234.600 34.900 ;
        RECT 235.800 34.800 236.200 34.900 ;
        RECT 235.000 33.800 235.400 34.600 ;
        RECT 235.800 34.100 236.100 34.800 ;
        RECT 237.400 34.400 237.800 35.200 ;
        RECT 238.100 34.200 238.400 35.900 ;
        RECT 239.000 35.800 239.400 35.900 ;
        RECT 239.800 35.800 240.200 36.600 ;
        RECT 239.000 35.100 239.300 35.800 ;
        RECT 240.600 35.100 241.000 39.900 ;
        RECT 242.200 35.700 242.600 39.900 ;
        RECT 244.400 38.200 244.800 39.900 ;
        RECT 243.800 37.900 244.800 38.200 ;
        RECT 246.600 37.900 247.000 39.900 ;
        RECT 248.700 37.900 249.300 39.900 ;
        RECT 243.800 37.500 244.200 37.900 ;
        RECT 246.600 37.600 246.900 37.900 ;
        RECT 245.500 37.300 247.300 37.600 ;
        RECT 248.600 37.500 249.000 37.900 ;
        RECT 245.500 37.200 245.900 37.300 ;
        RECT 246.900 37.200 247.300 37.300 ;
        RECT 243.800 36.500 244.200 36.600 ;
        RECT 246.100 36.500 246.500 36.600 ;
        RECT 243.800 36.200 246.500 36.500 ;
        RECT 246.800 36.500 247.900 36.800 ;
        RECT 246.800 35.900 247.100 36.500 ;
        RECT 247.500 36.400 247.900 36.500 ;
        RECT 248.700 36.600 249.400 37.000 ;
        RECT 248.700 36.100 249.000 36.600 ;
        RECT 244.700 35.700 247.100 35.900 ;
        RECT 242.200 35.600 247.100 35.700 ;
        RECT 247.800 35.800 249.000 36.100 ;
        RECT 242.200 35.500 245.100 35.600 ;
        RECT 242.200 35.400 245.000 35.500 ;
        RECT 245.400 35.100 245.800 35.200 ;
        RECT 239.000 34.800 241.000 35.100 ;
        RECT 236.600 34.100 237.000 34.200 ;
        RECT 238.100 34.100 239.400 34.200 ;
        RECT 239.800 34.100 240.200 34.200 ;
        RECT 235.800 33.800 237.400 34.100 ;
        RECT 238.100 33.800 240.200 34.100 ;
        RECT 237.000 33.600 237.400 33.800 ;
        RECT 236.700 33.100 238.500 33.300 ;
        RECT 239.000 33.100 239.300 33.800 ;
        RECT 240.600 33.100 241.000 34.800 ;
        RECT 243.300 34.800 245.800 35.100 ;
        RECT 243.300 34.700 243.700 34.800 ;
        RECT 244.600 34.700 245.000 34.800 ;
        RECT 244.100 34.200 244.500 34.300 ;
        RECT 247.800 34.200 248.100 35.800 ;
        RECT 251.000 35.600 251.400 39.900 ;
        RECT 249.300 35.300 251.400 35.600 ;
        RECT 249.300 35.200 249.700 35.300 ;
        RECT 250.100 34.900 250.500 35.000 ;
        RECT 248.600 34.600 250.500 34.900 ;
        RECT 248.600 34.500 249.000 34.600 ;
        RECT 241.400 33.400 241.800 34.200 ;
        RECT 242.600 33.900 248.100 34.200 ;
        RECT 242.600 33.800 243.400 33.900 ;
        RECT 231.800 32.800 233.800 33.100 ;
        RECT 231.900 32.100 232.200 32.800 ;
        RECT 233.500 32.400 233.900 32.800 ;
        RECT 231.800 31.100 232.200 32.100 ;
        RECT 234.200 31.100 234.600 33.100 ;
        RECT 236.600 33.000 238.600 33.100 ;
        RECT 236.600 31.100 237.000 33.000 ;
        RECT 238.200 31.100 238.600 33.000 ;
        RECT 239.000 31.100 239.400 33.100 ;
        RECT 240.100 32.800 241.000 33.100 ;
        RECT 240.100 31.100 240.500 32.800 ;
        RECT 242.200 31.100 242.600 33.500 ;
        RECT 244.700 32.800 245.000 33.900 ;
        RECT 247.500 33.800 247.900 33.900 ;
        RECT 251.000 33.600 251.400 35.300 ;
        RECT 249.500 33.300 251.400 33.600 ;
        RECT 249.500 33.200 249.900 33.300 ;
        RECT 243.800 32.100 244.200 32.500 ;
        RECT 244.600 32.400 245.000 32.800 ;
        RECT 245.500 32.700 245.900 32.800 ;
        RECT 245.500 32.400 246.900 32.700 ;
        RECT 246.600 32.100 246.900 32.400 ;
        RECT 248.600 32.100 249.000 32.500 ;
        RECT 243.800 31.800 244.800 32.100 ;
        RECT 244.400 31.100 244.800 31.800 ;
        RECT 246.600 31.100 247.000 32.100 ;
        RECT 248.600 31.800 249.300 32.100 ;
        RECT 248.700 31.100 249.300 31.800 ;
        RECT 251.000 31.100 251.400 33.300 ;
        RECT 1.900 28.200 2.300 29.900 ;
        RECT 1.400 27.900 2.300 28.200 ;
        RECT 3.000 27.900 3.400 29.900 ;
        RECT 3.800 28.000 4.200 29.900 ;
        RECT 5.400 28.000 5.800 29.900 ;
        RECT 7.500 28.200 7.900 29.900 ;
        RECT 3.800 27.900 5.800 28.000 ;
        RECT 7.000 27.900 7.900 28.200 ;
        RECT 8.600 27.900 9.000 29.900 ;
        RECT 9.400 28.000 9.800 29.900 ;
        RECT 11.000 28.000 11.400 29.900 ;
        RECT 9.400 27.900 11.400 28.000 ;
        RECT 0.600 26.800 1.000 27.600 ;
        RECT 1.400 26.100 1.800 27.900 ;
        RECT 3.100 27.200 3.400 27.900 ;
        RECT 3.900 27.700 5.700 27.900 ;
        RECT 5.000 27.200 5.400 27.400 ;
        RECT 3.000 26.800 4.300 27.200 ;
        RECT 5.000 26.900 5.800 27.200 ;
        RECT 5.400 26.800 5.800 26.900 ;
        RECT 6.200 26.800 6.600 27.600 ;
        RECT 1.400 25.800 3.300 26.100 ;
        RECT 1.400 21.100 1.800 25.800 ;
        RECT 3.000 25.200 3.300 25.800 ;
        RECT 2.200 24.400 2.600 25.200 ;
        RECT 3.000 25.100 3.400 25.200 ;
        RECT 4.000 25.100 4.300 26.800 ;
        RECT 4.600 25.800 5.000 26.600 ;
        RECT 7.000 26.100 7.400 27.900 ;
        RECT 8.700 27.200 9.000 27.900 ;
        RECT 9.500 27.700 11.300 27.900 ;
        RECT 11.800 27.500 12.200 29.900 ;
        RECT 14.000 29.200 14.400 29.900 ;
        RECT 13.400 28.900 14.400 29.200 ;
        RECT 16.200 28.900 16.600 29.900 ;
        RECT 18.300 29.200 18.900 29.900 ;
        RECT 18.200 28.900 18.900 29.200 ;
        RECT 13.400 28.500 13.800 28.900 ;
        RECT 16.200 28.600 16.500 28.900 ;
        RECT 14.200 28.200 14.600 28.600 ;
        RECT 15.100 28.300 16.500 28.600 ;
        RECT 18.200 28.500 18.600 28.900 ;
        RECT 15.100 28.200 15.500 28.300 ;
        RECT 10.600 27.200 11.000 27.400 ;
        RECT 8.600 26.800 9.900 27.200 ;
        RECT 10.600 26.900 11.400 27.200 ;
        RECT 11.000 26.800 11.400 26.900 ;
        RECT 12.200 27.100 13.000 27.200 ;
        RECT 14.300 27.100 14.600 28.200 ;
        RECT 19.100 27.700 19.500 27.800 ;
        RECT 20.600 27.700 21.000 29.900 ;
        RECT 19.100 27.400 21.000 27.700 ;
        RECT 21.400 27.500 21.800 29.900 ;
        RECT 23.600 29.200 24.000 29.900 ;
        RECT 23.000 28.900 24.000 29.200 ;
        RECT 25.800 28.900 26.200 29.900 ;
        RECT 27.900 29.200 28.500 29.900 ;
        RECT 27.800 28.900 28.500 29.200 ;
        RECT 23.000 28.500 23.400 28.900 ;
        RECT 25.800 28.600 26.100 28.900 ;
        RECT 23.800 28.200 24.200 28.600 ;
        RECT 24.700 28.300 26.100 28.600 ;
        RECT 27.800 28.500 28.200 28.900 ;
        RECT 24.700 28.200 25.100 28.300 ;
        RECT 16.600 27.100 17.500 27.200 ;
        RECT 12.200 26.800 17.700 27.100 ;
        RECT 7.000 25.800 8.900 26.100 ;
        RECT 3.000 24.800 3.700 25.100 ;
        RECT 4.000 24.800 4.500 25.100 ;
        RECT 3.400 24.200 3.700 24.800 ;
        RECT 3.400 23.800 3.800 24.200 ;
        RECT 4.100 21.100 4.500 24.800 ;
        RECT 7.000 21.100 7.400 25.800 ;
        RECT 8.600 25.200 8.900 25.800 ;
        RECT 9.600 25.200 9.900 26.800 ;
        RECT 13.700 26.700 14.100 26.800 ;
        RECT 10.200 25.800 10.600 26.600 ;
        RECT 12.900 26.200 13.300 26.300 ;
        RECT 14.200 26.200 14.600 26.300 ;
        RECT 17.400 26.200 17.700 26.800 ;
        RECT 18.200 26.400 18.600 26.500 ;
        RECT 12.900 25.900 15.400 26.200 ;
        RECT 15.000 25.800 15.400 25.900 ;
        RECT 17.400 25.800 17.800 26.200 ;
        RECT 18.200 26.100 20.100 26.400 ;
        RECT 19.700 26.000 20.100 26.100 ;
        RECT 11.800 25.500 14.600 25.600 ;
        RECT 11.800 25.400 14.700 25.500 ;
        RECT 11.800 25.300 16.700 25.400 ;
        RECT 7.800 24.400 8.200 25.200 ;
        RECT 8.600 25.100 9.000 25.200 ;
        RECT 8.600 24.800 9.300 25.100 ;
        RECT 9.600 24.800 10.600 25.200 ;
        RECT 9.000 24.200 9.300 24.800 ;
        RECT 9.000 23.800 9.400 24.200 ;
        RECT 9.700 21.100 10.100 24.800 ;
        RECT 11.800 21.100 12.200 25.300 ;
        RECT 14.300 25.100 16.700 25.300 ;
        RECT 13.400 24.500 16.100 24.800 ;
        RECT 13.400 24.400 13.800 24.500 ;
        RECT 15.700 24.400 16.100 24.500 ;
        RECT 16.400 24.500 16.700 25.100 ;
        RECT 17.400 25.200 17.700 25.800 ;
        RECT 18.900 25.700 19.300 25.800 ;
        RECT 20.600 25.700 21.000 27.400 ;
        RECT 21.800 27.100 22.600 27.200 ;
        RECT 23.900 27.100 24.200 28.200 ;
        RECT 28.700 27.700 29.100 27.800 ;
        RECT 30.200 27.700 30.600 29.900 ;
        RECT 28.700 27.400 30.600 27.700 ;
        RECT 26.700 27.100 27.100 27.200 ;
        RECT 21.800 26.800 27.300 27.100 ;
        RECT 23.300 26.700 23.700 26.800 ;
        RECT 22.500 26.200 22.900 26.300 ;
        RECT 22.500 25.900 25.000 26.200 ;
        RECT 24.600 25.800 25.000 25.900 ;
        RECT 26.200 26.100 26.600 26.200 ;
        RECT 27.000 26.100 27.300 26.800 ;
        RECT 27.800 26.400 28.200 26.500 ;
        RECT 27.800 26.100 29.700 26.400 ;
        RECT 26.200 25.800 27.300 26.100 ;
        RECT 29.300 26.000 29.700 26.100 ;
        RECT 18.900 25.400 21.000 25.700 ;
        RECT 17.400 24.900 18.600 25.200 ;
        RECT 17.100 24.500 17.500 24.600 ;
        RECT 16.400 24.200 17.500 24.500 ;
        RECT 18.300 24.400 18.600 24.900 ;
        RECT 18.300 24.000 19.000 24.400 ;
        RECT 15.100 23.700 15.500 23.800 ;
        RECT 16.500 23.700 16.900 23.800 ;
        RECT 13.400 23.100 13.800 23.500 ;
        RECT 15.100 23.400 16.900 23.700 ;
        RECT 16.200 23.100 16.500 23.400 ;
        RECT 18.200 23.100 18.600 23.500 ;
        RECT 13.400 22.800 14.400 23.100 ;
        RECT 14.000 21.100 14.400 22.800 ;
        RECT 16.200 21.100 16.600 23.100 ;
        RECT 18.300 21.100 18.900 23.100 ;
        RECT 20.600 21.100 21.000 25.400 ;
        RECT 21.400 25.500 24.200 25.600 ;
        RECT 21.400 25.400 24.300 25.500 ;
        RECT 21.400 25.300 26.300 25.400 ;
        RECT 21.400 21.100 21.800 25.300 ;
        RECT 23.900 25.100 26.300 25.300 ;
        RECT 23.000 24.500 25.700 24.800 ;
        RECT 23.000 24.400 23.400 24.500 ;
        RECT 25.300 24.400 25.700 24.500 ;
        RECT 26.000 24.500 26.300 25.100 ;
        RECT 27.000 25.200 27.300 25.800 ;
        RECT 28.500 25.700 28.900 25.800 ;
        RECT 30.200 25.700 30.600 27.400 ;
        RECT 28.500 25.400 30.600 25.700 ;
        RECT 27.000 24.900 28.200 25.200 ;
        RECT 26.700 24.500 27.100 24.600 ;
        RECT 26.000 24.200 27.100 24.500 ;
        RECT 27.900 24.400 28.200 24.900 ;
        RECT 27.900 24.000 28.600 24.400 ;
        RECT 24.700 23.700 25.100 23.800 ;
        RECT 26.100 23.700 26.500 23.800 ;
        RECT 23.000 23.100 23.400 23.500 ;
        RECT 24.700 23.400 26.500 23.700 ;
        RECT 25.800 23.100 26.100 23.400 ;
        RECT 27.800 23.100 28.200 23.500 ;
        RECT 23.000 22.800 24.000 23.100 ;
        RECT 23.600 21.100 24.000 22.800 ;
        RECT 25.800 21.100 26.200 23.100 ;
        RECT 27.900 21.100 28.500 23.100 ;
        RECT 30.200 21.100 30.600 25.400 ;
        RECT 31.000 27.700 31.400 29.900 ;
        RECT 33.100 29.200 33.700 29.900 ;
        RECT 33.100 28.900 33.800 29.200 ;
        RECT 35.400 28.900 35.800 29.900 ;
        RECT 37.600 29.200 38.000 29.900 ;
        RECT 37.600 28.900 38.600 29.200 ;
        RECT 33.400 28.500 33.800 28.900 ;
        RECT 35.500 28.600 35.800 28.900 ;
        RECT 35.500 28.300 36.900 28.600 ;
        RECT 36.500 28.200 36.900 28.300 ;
        RECT 37.400 27.800 37.800 28.600 ;
        RECT 38.200 28.500 38.600 28.900 ;
        RECT 32.500 27.700 32.900 27.800 ;
        RECT 31.000 27.400 32.900 27.700 ;
        RECT 31.000 25.700 31.400 27.400 ;
        RECT 34.500 27.100 34.900 27.200 ;
        RECT 37.400 27.100 37.700 27.800 ;
        RECT 39.800 27.500 40.200 29.900 ;
        RECT 40.600 27.700 41.000 29.900 ;
        RECT 42.700 29.200 43.300 29.900 ;
        RECT 42.700 28.900 43.400 29.200 ;
        RECT 45.000 28.900 45.400 29.900 ;
        RECT 47.200 29.200 47.600 29.900 ;
        RECT 47.200 28.900 48.200 29.200 ;
        RECT 43.000 28.500 43.400 28.900 ;
        RECT 45.100 28.600 45.400 28.900 ;
        RECT 45.100 28.300 46.500 28.600 ;
        RECT 46.100 28.200 46.500 28.300 ;
        RECT 47.000 28.200 47.400 28.600 ;
        RECT 47.800 28.500 48.200 28.900 ;
        RECT 42.100 27.700 42.500 27.800 ;
        RECT 40.600 27.400 42.500 27.700 ;
        RECT 39.000 27.100 39.800 27.200 ;
        RECT 34.300 26.800 39.800 27.100 ;
        RECT 33.400 26.400 33.800 26.500 ;
        RECT 31.900 26.100 33.800 26.400 ;
        RECT 31.900 26.000 32.300 26.100 ;
        RECT 32.700 25.700 33.100 25.800 ;
        RECT 31.000 25.400 33.100 25.700 ;
        RECT 31.000 21.100 31.400 25.400 ;
        RECT 34.300 25.200 34.600 26.800 ;
        RECT 37.900 26.700 38.300 26.800 ;
        RECT 37.400 26.200 37.800 26.300 ;
        RECT 38.700 26.200 39.100 26.300 ;
        RECT 36.600 25.900 39.100 26.200 ;
        RECT 36.600 25.800 37.000 25.900 ;
        RECT 40.600 25.700 41.000 27.400 ;
        RECT 44.100 27.100 44.500 27.200 ;
        RECT 47.000 27.100 47.300 28.200 ;
        RECT 49.400 27.500 49.800 29.900 ;
        RECT 51.800 28.500 52.200 29.500 ;
        RECT 53.900 29.200 54.300 29.500 ;
        RECT 53.900 28.800 54.600 29.200 ;
        RECT 51.800 27.400 52.100 28.500 ;
        RECT 53.900 28.000 54.300 28.800 ;
        RECT 56.600 28.000 57.000 29.900 ;
        RECT 58.200 28.000 58.600 29.900 ;
        RECT 53.900 27.700 54.700 28.000 ;
        RECT 56.600 27.900 58.600 28.000 ;
        RECT 59.000 27.900 59.400 29.900 ;
        RECT 60.100 28.200 60.500 29.900 ;
        RECT 60.100 27.900 61.000 28.200 ;
        RECT 56.700 27.700 58.500 27.900 ;
        RECT 54.300 27.500 54.700 27.700 ;
        RECT 48.600 27.100 49.400 27.200 ;
        RECT 51.800 27.100 53.900 27.400 ;
        RECT 43.900 26.800 49.400 27.100 ;
        RECT 53.400 26.900 53.900 27.100 ;
        RECT 54.400 27.200 54.700 27.500 ;
        RECT 57.000 27.200 57.400 27.400 ;
        RECT 59.000 27.200 59.300 27.900 ;
        RECT 43.000 26.400 43.400 26.500 ;
        RECT 41.500 26.100 43.400 26.400 ;
        RECT 41.500 26.000 41.900 26.100 ;
        RECT 42.300 25.700 42.700 25.800 ;
        RECT 37.400 25.500 40.200 25.600 ;
        RECT 37.300 25.400 40.200 25.500 ;
        RECT 33.400 24.900 34.600 25.200 ;
        RECT 35.300 25.300 40.200 25.400 ;
        RECT 35.300 25.100 37.700 25.300 ;
        RECT 33.400 24.400 33.700 24.900 ;
        RECT 33.000 24.000 33.700 24.400 ;
        RECT 34.500 24.500 34.900 24.600 ;
        RECT 35.300 24.500 35.600 25.100 ;
        RECT 34.500 24.200 35.600 24.500 ;
        RECT 35.900 24.500 38.600 24.800 ;
        RECT 35.900 24.400 36.300 24.500 ;
        RECT 38.200 24.400 38.600 24.500 ;
        RECT 35.100 23.700 35.500 23.800 ;
        RECT 36.500 23.700 36.900 23.800 ;
        RECT 33.400 23.100 33.800 23.500 ;
        RECT 35.100 23.400 36.900 23.700 ;
        RECT 35.500 23.100 35.800 23.400 ;
        RECT 38.200 23.100 38.600 23.500 ;
        RECT 33.100 21.100 33.700 23.100 ;
        RECT 35.400 21.100 35.800 23.100 ;
        RECT 37.600 22.800 38.600 23.100 ;
        RECT 37.600 21.100 38.000 22.800 ;
        RECT 39.800 21.100 40.200 25.300 ;
        RECT 40.600 25.400 42.700 25.700 ;
        RECT 40.600 21.100 41.000 25.400 ;
        RECT 43.900 25.200 44.200 26.800 ;
        RECT 47.500 26.700 47.900 26.800 ;
        RECT 47.000 26.200 47.400 26.300 ;
        RECT 48.300 26.200 48.700 26.300 ;
        RECT 46.200 25.900 48.700 26.200 ;
        RECT 46.200 25.800 46.600 25.900 ;
        RECT 51.800 25.800 52.200 26.600 ;
        RECT 52.600 25.800 53.000 26.600 ;
        RECT 53.400 26.500 54.100 26.900 ;
        RECT 54.400 26.800 55.400 27.200 ;
        RECT 56.600 26.900 57.400 27.200 ;
        RECT 56.600 26.800 57.000 26.900 ;
        RECT 58.100 26.800 59.400 27.200 ;
        RECT 47.000 25.500 49.800 25.600 ;
        RECT 53.400 25.500 53.700 26.500 ;
        RECT 46.900 25.400 49.800 25.500 ;
        RECT 43.000 24.900 44.200 25.200 ;
        RECT 44.900 25.300 49.800 25.400 ;
        RECT 44.900 25.100 47.300 25.300 ;
        RECT 43.000 24.400 43.300 24.900 ;
        RECT 42.600 24.000 43.300 24.400 ;
        RECT 44.100 24.500 44.500 24.600 ;
        RECT 44.900 24.500 45.200 25.100 ;
        RECT 44.100 24.200 45.200 24.500 ;
        RECT 45.500 24.500 48.200 24.800 ;
        RECT 45.500 24.400 45.900 24.500 ;
        RECT 47.800 24.400 48.200 24.500 ;
        RECT 44.700 23.700 45.100 23.800 ;
        RECT 46.100 23.700 46.500 23.800 ;
        RECT 43.000 23.100 43.400 23.500 ;
        RECT 44.700 23.400 46.500 23.700 ;
        RECT 45.100 23.100 45.400 23.400 ;
        RECT 47.800 23.100 48.200 23.500 ;
        RECT 42.700 21.100 43.300 23.100 ;
        RECT 45.000 21.100 45.400 23.100 ;
        RECT 47.200 22.800 48.200 23.100 ;
        RECT 47.200 21.100 47.600 22.800 ;
        RECT 49.400 21.100 49.800 25.300 ;
        RECT 51.800 25.200 53.700 25.500 ;
        RECT 51.800 23.500 52.100 25.200 ;
        RECT 54.400 24.900 54.700 26.800 ;
        RECT 55.000 25.400 55.400 26.200 ;
        RECT 57.400 25.800 57.800 26.600 ;
        RECT 58.100 25.100 58.400 26.800 ;
        RECT 60.600 26.100 61.000 27.900 ;
        RECT 61.400 26.800 61.800 27.600 ;
        RECT 62.200 27.500 62.600 29.900 ;
        RECT 64.400 29.200 64.800 29.900 ;
        RECT 63.800 28.900 64.800 29.200 ;
        RECT 66.600 28.900 67.000 29.900 ;
        RECT 68.700 29.200 69.300 29.900 ;
        RECT 68.600 28.900 69.300 29.200 ;
        RECT 63.800 28.500 64.200 28.900 ;
        RECT 66.600 28.600 66.900 28.900 ;
        RECT 64.600 28.200 65.000 28.600 ;
        RECT 65.500 28.300 66.900 28.600 ;
        RECT 68.600 28.500 69.000 28.900 ;
        RECT 65.500 28.200 65.900 28.300 ;
        RECT 62.600 27.100 63.400 27.200 ;
        RECT 64.700 27.100 65.000 28.200 ;
        RECT 69.500 27.700 69.900 27.800 ;
        RECT 71.000 27.700 71.400 29.900 ;
        RECT 73.700 29.200 74.100 29.500 ;
        RECT 73.400 28.800 74.100 29.200 ;
        RECT 73.700 28.000 74.100 28.800 ;
        RECT 75.800 28.500 76.200 29.500 ;
        RECT 69.500 27.400 71.400 27.700 ;
        RECT 66.200 27.100 66.600 27.200 ;
        RECT 67.500 27.100 67.900 27.200 ;
        RECT 62.600 26.800 68.100 27.100 ;
        RECT 64.100 26.700 64.500 26.800 ;
        RECT 59.000 25.800 61.000 26.100 ;
        RECT 63.300 26.200 63.700 26.300 ;
        RECT 63.300 25.900 65.800 26.200 ;
        RECT 65.400 25.800 65.800 25.900 ;
        RECT 59.000 25.200 59.300 25.800 ;
        RECT 59.000 25.100 59.400 25.200 ;
        RECT 53.900 24.600 54.700 24.900 ;
        RECT 57.900 24.800 58.400 25.100 ;
        RECT 58.700 24.800 59.400 25.100 ;
        RECT 51.800 21.500 52.200 23.500 ;
        RECT 53.900 21.100 54.300 24.600 ;
        RECT 57.900 21.100 58.300 24.800 ;
        RECT 58.700 24.200 59.000 24.800 ;
        RECT 59.800 24.400 60.200 25.200 ;
        RECT 58.600 23.800 59.000 24.200 ;
        RECT 60.600 21.100 61.000 25.800 ;
        RECT 62.200 25.500 65.000 25.600 ;
        RECT 62.200 25.400 65.100 25.500 ;
        RECT 62.200 25.300 67.100 25.400 ;
        RECT 62.200 21.100 62.600 25.300 ;
        RECT 64.700 25.100 67.100 25.300 ;
        RECT 63.800 24.500 66.500 24.800 ;
        RECT 63.800 24.400 64.200 24.500 ;
        RECT 66.100 24.400 66.500 24.500 ;
        RECT 66.800 24.500 67.100 25.100 ;
        RECT 67.800 25.200 68.100 26.800 ;
        RECT 68.600 26.400 69.000 26.500 ;
        RECT 68.600 26.100 70.500 26.400 ;
        RECT 70.100 26.000 70.500 26.100 ;
        RECT 69.300 25.700 69.700 25.800 ;
        RECT 71.000 25.700 71.400 27.400 ;
        RECT 73.300 27.700 74.100 28.000 ;
        RECT 73.300 27.500 73.700 27.700 ;
        RECT 73.300 27.200 73.600 27.500 ;
        RECT 75.900 27.400 76.200 28.500 ;
        RECT 77.900 28.200 78.300 29.900 ;
        RECT 77.400 27.900 78.300 28.200 ;
        RECT 79.000 27.900 79.400 29.900 ;
        RECT 79.800 28.000 80.200 29.900 ;
        RECT 81.400 28.000 81.800 29.900 ;
        RECT 79.800 27.900 81.800 28.000 ;
        RECT 82.200 28.000 82.600 29.900 ;
        RECT 83.800 28.000 84.200 29.900 ;
        RECT 82.200 27.900 84.200 28.000 ;
        RECT 84.600 27.900 85.000 29.900 ;
        RECT 72.600 26.800 73.600 27.200 ;
        RECT 74.100 27.100 76.200 27.400 ;
        RECT 74.100 26.900 74.600 27.100 ;
        RECT 69.300 25.400 71.400 25.700 ;
        RECT 72.600 25.400 73.000 26.200 ;
        RECT 67.800 24.900 69.000 25.200 ;
        RECT 67.500 24.500 67.900 24.600 ;
        RECT 66.800 24.200 67.900 24.500 ;
        RECT 68.700 24.400 69.000 24.900 ;
        RECT 68.700 24.000 69.400 24.400 ;
        RECT 65.500 23.700 65.900 23.800 ;
        RECT 66.900 23.700 67.300 23.800 ;
        RECT 63.800 23.100 64.200 23.500 ;
        RECT 65.500 23.400 67.300 23.700 ;
        RECT 66.600 23.100 66.900 23.400 ;
        RECT 68.600 23.100 69.000 23.500 ;
        RECT 63.800 22.800 64.800 23.100 ;
        RECT 64.400 21.100 64.800 22.800 ;
        RECT 66.600 21.100 67.000 23.100 ;
        RECT 68.700 21.100 69.300 23.100 ;
        RECT 71.000 21.100 71.400 25.400 ;
        RECT 73.300 24.900 73.600 26.800 ;
        RECT 73.900 26.500 74.600 26.900 ;
        RECT 76.600 26.800 77.000 27.600 ;
        RECT 74.300 25.500 74.600 26.500 ;
        RECT 75.000 25.800 75.400 26.600 ;
        RECT 75.800 25.800 76.200 26.600 ;
        RECT 77.400 26.100 77.800 27.900 ;
        RECT 79.100 27.200 79.400 27.900 ;
        RECT 79.900 27.700 81.700 27.900 ;
        RECT 82.300 27.700 84.100 27.900 ;
        RECT 81.000 27.200 81.400 27.400 ;
        RECT 82.600 27.200 83.000 27.400 ;
        RECT 84.600 27.200 84.900 27.900 ;
        RECT 85.400 27.700 85.800 29.900 ;
        RECT 87.500 29.200 88.100 29.900 ;
        RECT 87.500 28.900 88.200 29.200 ;
        RECT 89.800 28.900 90.200 29.900 ;
        RECT 92.000 29.200 92.400 29.900 ;
        RECT 92.000 28.900 93.000 29.200 ;
        RECT 87.800 28.500 88.200 28.900 ;
        RECT 89.900 28.600 90.200 28.900 ;
        RECT 89.900 28.300 91.300 28.600 ;
        RECT 90.900 28.200 91.300 28.300 ;
        RECT 91.800 28.200 92.200 28.600 ;
        RECT 92.600 28.500 93.000 28.900 ;
        RECT 86.900 27.700 87.300 27.800 ;
        RECT 85.400 27.400 87.300 27.700 ;
        RECT 78.200 27.100 78.600 27.200 ;
        RECT 79.000 27.100 80.300 27.200 ;
        RECT 78.200 26.800 80.300 27.100 ;
        RECT 81.000 27.100 81.800 27.200 ;
        RECT 82.200 27.100 83.000 27.200 ;
        RECT 81.000 26.900 83.000 27.100 ;
        RECT 81.400 26.800 82.600 26.900 ;
        RECT 83.700 26.800 85.000 27.200 ;
        RECT 77.400 25.800 79.300 26.100 ;
        RECT 74.300 25.200 76.200 25.500 ;
        RECT 73.300 24.600 74.100 24.900 ;
        RECT 73.700 21.100 74.100 24.600 ;
        RECT 75.900 23.500 76.200 25.200 ;
        RECT 75.800 21.500 76.200 23.500 ;
        RECT 77.400 21.100 77.800 25.800 ;
        RECT 79.000 25.200 79.300 25.800 ;
        RECT 78.200 24.400 78.600 25.200 ;
        RECT 79.000 25.100 79.400 25.200 ;
        RECT 80.000 25.100 80.300 26.800 ;
        RECT 80.600 25.800 81.000 26.600 ;
        RECT 83.000 25.800 83.400 26.600 ;
        RECT 83.700 26.200 84.000 26.800 ;
        RECT 83.700 25.800 84.200 26.200 ;
        RECT 83.700 25.100 84.000 25.800 ;
        RECT 85.400 25.700 85.800 27.400 ;
        RECT 88.900 27.100 89.300 27.200 ;
        RECT 91.800 27.100 92.100 28.200 ;
        RECT 94.200 27.500 94.600 29.900 ;
        RECT 96.600 27.700 97.000 29.900 ;
        RECT 98.700 29.200 99.300 29.900 ;
        RECT 98.700 28.900 99.400 29.200 ;
        RECT 101.000 28.900 101.400 29.900 ;
        RECT 103.200 29.200 103.600 29.900 ;
        RECT 103.200 28.900 104.200 29.200 ;
        RECT 99.000 28.500 99.400 28.900 ;
        RECT 101.100 28.600 101.400 28.900 ;
        RECT 101.100 28.300 102.500 28.600 ;
        RECT 102.100 28.200 102.500 28.300 ;
        RECT 103.000 28.200 103.400 28.600 ;
        RECT 103.800 28.500 104.200 28.900 ;
        RECT 98.100 27.700 98.500 27.800 ;
        RECT 96.600 27.400 98.500 27.700 ;
        RECT 93.400 27.100 94.200 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 88.700 26.800 96.200 27.100 ;
        RECT 87.800 26.400 88.200 26.500 ;
        RECT 86.300 26.100 88.200 26.400 ;
        RECT 86.300 26.000 86.700 26.100 ;
        RECT 87.100 25.700 87.500 25.800 ;
        RECT 85.400 25.400 87.500 25.700 ;
        RECT 84.600 25.100 85.000 25.200 ;
        RECT 79.000 24.800 79.700 25.100 ;
        RECT 80.000 24.800 80.500 25.100 ;
        RECT 79.400 24.200 79.700 24.800 ;
        RECT 79.400 23.800 79.800 24.200 ;
        RECT 80.100 21.100 80.500 24.800 ;
        RECT 83.500 24.800 84.000 25.100 ;
        RECT 84.300 24.800 85.000 25.100 ;
        RECT 83.500 21.100 83.900 24.800 ;
        RECT 84.300 24.200 84.600 24.800 ;
        RECT 84.200 23.800 84.600 24.200 ;
        RECT 85.400 21.100 85.800 25.400 ;
        RECT 88.700 25.200 89.000 26.800 ;
        RECT 92.300 26.700 92.700 26.800 ;
        RECT 93.100 26.200 93.500 26.300 ;
        RECT 90.200 26.100 90.600 26.200 ;
        RECT 91.000 26.100 93.500 26.200 ;
        RECT 90.200 25.900 93.500 26.100 ;
        RECT 90.200 25.800 91.400 25.900 ;
        RECT 96.600 25.700 97.000 27.400 ;
        RECT 100.100 27.100 100.500 27.200 ;
        RECT 103.000 27.100 103.300 28.200 ;
        RECT 105.400 27.500 105.800 29.900 ;
        RECT 107.500 28.200 107.900 29.900 ;
        RECT 107.000 27.900 107.900 28.200 ;
        RECT 108.600 27.900 109.000 29.900 ;
        RECT 109.400 28.000 109.800 29.900 ;
        RECT 111.000 28.000 111.400 29.900 ;
        RECT 109.400 27.900 111.400 28.000 ;
        RECT 111.800 28.000 112.200 29.900 ;
        RECT 113.400 28.000 113.800 29.900 ;
        RECT 111.800 27.900 113.800 28.000 ;
        RECT 104.600 27.100 105.400 27.200 ;
        RECT 99.900 26.800 105.400 27.100 ;
        RECT 106.200 26.800 106.600 27.600 ;
        RECT 99.000 26.400 99.400 26.500 ;
        RECT 97.500 26.100 99.400 26.400 ;
        RECT 99.900 26.200 100.200 26.800 ;
        RECT 103.500 26.700 103.900 26.800 ;
        RECT 103.000 26.200 103.400 26.300 ;
        RECT 104.300 26.200 104.700 26.300 ;
        RECT 97.500 26.000 97.900 26.100 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 102.200 25.900 104.700 26.200 ;
        RECT 107.000 26.100 107.400 27.900 ;
        RECT 108.700 27.200 109.000 27.900 ;
        RECT 109.500 27.700 111.300 27.900 ;
        RECT 111.900 27.700 113.700 27.900 ;
        RECT 114.200 27.800 114.600 29.900 ;
        RECT 115.300 28.200 115.700 29.900 ;
        RECT 115.300 27.900 116.200 28.200 ;
        RECT 110.600 27.200 111.000 27.400 ;
        RECT 112.200 27.200 112.600 27.400 ;
        RECT 114.200 27.200 114.500 27.800 ;
        RECT 107.800 27.100 108.200 27.200 ;
        RECT 108.600 27.100 109.900 27.200 ;
        RECT 107.800 26.800 109.900 27.100 ;
        RECT 110.600 26.900 111.400 27.200 ;
        RECT 111.000 26.800 111.400 26.900 ;
        RECT 111.800 26.900 112.600 27.200 ;
        RECT 111.800 26.800 112.200 26.900 ;
        RECT 113.300 26.800 114.600 27.200 ;
        RECT 102.200 25.800 102.600 25.900 ;
        RECT 107.000 25.800 108.900 26.100 ;
        RECT 98.300 25.700 98.700 25.800 ;
        RECT 91.800 25.500 94.600 25.600 ;
        RECT 91.700 25.400 94.600 25.500 ;
        RECT 87.800 24.900 89.000 25.200 ;
        RECT 89.700 25.300 94.600 25.400 ;
        RECT 89.700 25.100 92.100 25.300 ;
        RECT 87.800 24.400 88.100 24.900 ;
        RECT 87.400 24.000 88.100 24.400 ;
        RECT 88.900 24.500 89.300 24.600 ;
        RECT 89.700 24.500 90.000 25.100 ;
        RECT 88.900 24.200 90.000 24.500 ;
        RECT 90.300 24.500 93.000 24.800 ;
        RECT 90.300 24.400 90.700 24.500 ;
        RECT 92.600 24.400 93.000 24.500 ;
        RECT 89.500 23.700 89.900 23.800 ;
        RECT 90.900 23.700 91.300 23.800 ;
        RECT 87.800 23.100 88.200 23.500 ;
        RECT 89.500 23.400 91.300 23.700 ;
        RECT 89.900 23.100 90.200 23.400 ;
        RECT 92.600 23.100 93.000 23.500 ;
        RECT 87.500 21.100 88.100 23.100 ;
        RECT 89.800 21.100 90.200 23.100 ;
        RECT 92.000 22.800 93.000 23.100 ;
        RECT 92.000 21.100 92.400 22.800 ;
        RECT 94.200 21.100 94.600 25.300 ;
        RECT 96.600 25.400 98.700 25.700 ;
        RECT 96.600 21.100 97.000 25.400 ;
        RECT 99.900 25.200 100.200 25.800 ;
        RECT 103.000 25.500 105.800 25.600 ;
        RECT 102.900 25.400 105.800 25.500 ;
        RECT 99.000 24.900 100.200 25.200 ;
        RECT 100.900 25.300 105.800 25.400 ;
        RECT 100.900 25.100 103.300 25.300 ;
        RECT 99.000 24.400 99.300 24.900 ;
        RECT 98.600 24.000 99.300 24.400 ;
        RECT 100.100 24.500 100.500 24.600 ;
        RECT 100.900 24.500 101.200 25.100 ;
        RECT 100.100 24.200 101.200 24.500 ;
        RECT 101.500 24.500 104.200 24.800 ;
        RECT 101.500 24.400 101.900 24.500 ;
        RECT 103.800 24.400 104.200 24.500 ;
        RECT 100.700 23.700 101.100 23.800 ;
        RECT 102.100 23.700 102.500 23.800 ;
        RECT 99.000 23.100 99.400 23.500 ;
        RECT 100.700 23.400 102.500 23.700 ;
        RECT 101.100 23.100 101.400 23.400 ;
        RECT 103.800 23.100 104.200 23.500 ;
        RECT 98.700 21.100 99.300 23.100 ;
        RECT 101.000 21.100 101.400 23.100 ;
        RECT 103.200 22.800 104.200 23.100 ;
        RECT 103.200 21.100 103.600 22.800 ;
        RECT 105.400 21.100 105.800 25.300 ;
        RECT 107.000 21.100 107.400 25.800 ;
        RECT 108.600 25.200 108.900 25.800 ;
        RECT 107.800 24.400 108.200 25.200 ;
        RECT 108.600 25.100 109.000 25.200 ;
        RECT 109.600 25.100 109.900 26.800 ;
        RECT 110.200 25.800 110.600 26.600 ;
        RECT 111.000 26.100 111.400 26.200 ;
        RECT 112.600 26.100 113.000 26.600 ;
        RECT 111.000 25.800 113.000 26.100 ;
        RECT 113.300 25.100 113.600 26.800 ;
        RECT 115.800 26.100 116.200 27.900 ;
        RECT 116.600 26.800 117.000 27.600 ;
        RECT 117.400 27.500 117.800 29.900 ;
        RECT 119.600 29.200 120.000 29.900 ;
        RECT 119.000 28.900 120.000 29.200 ;
        RECT 121.800 28.900 122.200 29.900 ;
        RECT 123.900 29.200 124.500 29.900 ;
        RECT 123.800 28.900 124.500 29.200 ;
        RECT 119.000 28.500 119.400 28.900 ;
        RECT 121.800 28.600 122.100 28.900 ;
        RECT 119.800 28.200 120.200 28.600 ;
        RECT 120.700 28.300 122.100 28.600 ;
        RECT 123.800 28.500 124.200 28.900 ;
        RECT 120.700 28.200 121.100 28.300 ;
        RECT 117.800 27.100 118.600 27.200 ;
        RECT 119.900 27.100 120.200 28.200 ;
        RECT 124.700 27.700 125.100 27.800 ;
        RECT 126.200 27.700 126.600 29.900 ;
        RECT 127.000 28.000 127.400 29.900 ;
        RECT 128.600 28.000 129.000 29.900 ;
        RECT 127.000 27.900 129.000 28.000 ;
        RECT 129.400 27.900 129.800 29.900 ;
        RECT 130.500 28.200 130.900 29.900 ;
        RECT 130.500 27.900 131.400 28.200 ;
        RECT 127.100 27.700 128.900 27.900 ;
        RECT 124.700 27.400 126.600 27.700 ;
        RECT 122.700 27.100 123.100 27.200 ;
        RECT 117.800 26.800 123.300 27.100 ;
        RECT 119.300 26.700 119.700 26.800 ;
        RECT 114.200 25.800 116.200 26.100 ;
        RECT 118.500 26.200 118.900 26.300 ;
        RECT 119.800 26.200 120.200 26.300 ;
        RECT 118.500 25.900 121.000 26.200 ;
        RECT 120.600 25.800 121.000 25.900 ;
        RECT 122.200 26.100 122.600 26.200 ;
        RECT 123.000 26.100 123.300 26.800 ;
        RECT 123.800 26.400 124.200 26.500 ;
        RECT 123.800 26.100 125.700 26.400 ;
        RECT 122.200 25.800 123.300 26.100 ;
        RECT 125.300 26.000 125.700 26.100 ;
        RECT 114.200 25.200 114.500 25.800 ;
        RECT 114.200 25.100 114.600 25.200 ;
        RECT 108.600 24.800 109.300 25.100 ;
        RECT 109.600 24.800 110.100 25.100 ;
        RECT 109.000 24.200 109.300 24.800 ;
        RECT 109.000 23.800 109.400 24.200 ;
        RECT 109.700 21.100 110.100 24.800 ;
        RECT 113.100 24.800 113.600 25.100 ;
        RECT 113.900 24.800 114.600 25.100 ;
        RECT 113.100 21.100 113.500 24.800 ;
        RECT 113.900 24.200 114.200 24.800 ;
        RECT 115.000 24.400 115.400 25.200 ;
        RECT 113.800 23.800 114.200 24.200 ;
        RECT 115.800 21.100 116.200 25.800 ;
        RECT 117.400 25.500 120.200 25.600 ;
        RECT 117.400 25.400 120.300 25.500 ;
        RECT 117.400 25.300 122.300 25.400 ;
        RECT 117.400 21.100 117.800 25.300 ;
        RECT 119.900 25.100 122.300 25.300 ;
        RECT 119.000 24.500 121.700 24.800 ;
        RECT 119.000 24.400 119.400 24.500 ;
        RECT 121.300 24.400 121.700 24.500 ;
        RECT 122.000 24.500 122.300 25.100 ;
        RECT 123.000 25.200 123.300 25.800 ;
        RECT 124.500 25.700 124.900 25.800 ;
        RECT 126.200 25.700 126.600 27.400 ;
        RECT 127.400 27.200 127.800 27.400 ;
        RECT 129.400 27.200 129.700 27.900 ;
        RECT 127.000 26.900 127.800 27.200 ;
        RECT 128.500 27.100 129.800 27.200 ;
        RECT 130.200 27.100 130.600 27.200 ;
        RECT 127.000 26.800 127.400 26.900 ;
        RECT 128.500 26.800 130.600 27.100 ;
        RECT 127.800 25.800 128.200 26.600 ;
        RECT 124.500 25.400 126.600 25.700 ;
        RECT 123.000 24.900 124.200 25.200 ;
        RECT 122.700 24.500 123.100 24.600 ;
        RECT 122.000 24.200 123.100 24.500 ;
        RECT 123.900 24.400 124.200 24.900 ;
        RECT 123.900 24.000 124.600 24.400 ;
        RECT 120.700 23.700 121.100 23.800 ;
        RECT 122.100 23.700 122.500 23.800 ;
        RECT 119.000 23.100 119.400 23.500 ;
        RECT 120.700 23.400 122.500 23.700 ;
        RECT 121.800 23.100 122.100 23.400 ;
        RECT 123.800 23.100 124.200 23.500 ;
        RECT 119.000 22.800 120.000 23.100 ;
        RECT 119.600 21.100 120.000 22.800 ;
        RECT 121.800 21.100 122.200 23.100 ;
        RECT 123.900 21.100 124.500 23.100 ;
        RECT 126.200 21.100 126.600 25.400 ;
        RECT 128.500 25.100 128.800 26.800 ;
        RECT 131.000 26.100 131.400 27.900 ;
        RECT 131.800 26.800 132.200 27.600 ;
        RECT 132.600 27.500 133.000 29.900 ;
        RECT 134.800 29.200 135.200 29.900 ;
        RECT 134.200 28.900 135.200 29.200 ;
        RECT 137.000 28.900 137.400 29.900 ;
        RECT 139.100 29.200 139.700 29.900 ;
        RECT 139.000 28.900 139.700 29.200 ;
        RECT 134.200 28.500 134.600 28.900 ;
        RECT 137.000 28.600 137.300 28.900 ;
        RECT 135.000 28.200 135.400 28.600 ;
        RECT 135.900 28.300 137.300 28.600 ;
        RECT 139.000 28.500 139.400 28.900 ;
        RECT 135.900 28.200 136.300 28.300 ;
        RECT 133.000 27.100 133.800 27.200 ;
        RECT 135.100 27.100 135.400 28.200 ;
        RECT 139.900 27.700 140.300 27.800 ;
        RECT 141.400 27.700 141.800 29.900 ;
        RECT 142.200 27.900 142.600 29.900 ;
        RECT 143.000 28.000 143.400 29.900 ;
        RECT 144.600 28.000 145.000 29.900 ;
        RECT 143.000 27.900 145.000 28.000 ;
        RECT 145.400 28.500 145.800 29.500 ;
        RECT 147.500 29.200 147.900 29.500 ;
        RECT 147.000 28.800 147.900 29.200 ;
        RECT 139.900 27.400 141.800 27.700 ;
        RECT 137.900 27.100 138.300 27.200 ;
        RECT 133.000 26.800 138.500 27.100 ;
        RECT 134.500 26.700 134.900 26.800 ;
        RECT 129.400 25.800 131.400 26.100 ;
        RECT 133.700 26.200 134.100 26.300 ;
        RECT 135.000 26.200 135.400 26.300 ;
        RECT 133.700 25.900 136.200 26.200 ;
        RECT 135.800 25.800 136.200 25.900 ;
        RECT 129.400 25.200 129.700 25.800 ;
        RECT 129.400 25.100 129.800 25.200 ;
        RECT 128.300 24.800 128.800 25.100 ;
        RECT 129.100 24.800 129.800 25.100 ;
        RECT 128.300 21.100 128.700 24.800 ;
        RECT 129.100 24.200 129.400 24.800 ;
        RECT 130.200 24.400 130.600 25.200 ;
        RECT 129.000 23.800 129.400 24.200 ;
        RECT 131.000 21.100 131.400 25.800 ;
        RECT 132.600 25.500 135.400 25.600 ;
        RECT 132.600 25.400 135.500 25.500 ;
        RECT 132.600 25.300 137.500 25.400 ;
        RECT 132.600 21.100 133.000 25.300 ;
        RECT 135.100 25.100 137.500 25.300 ;
        RECT 134.200 24.500 136.900 24.800 ;
        RECT 134.200 24.400 134.600 24.500 ;
        RECT 136.500 24.400 136.900 24.500 ;
        RECT 137.200 24.500 137.500 25.100 ;
        RECT 138.200 25.200 138.500 26.800 ;
        RECT 139.000 26.400 139.400 26.500 ;
        RECT 139.000 26.100 140.900 26.400 ;
        RECT 140.500 26.000 140.900 26.100 ;
        RECT 139.700 25.700 140.100 25.800 ;
        RECT 141.400 25.700 141.800 27.400 ;
        RECT 142.300 27.200 142.600 27.900 ;
        RECT 143.100 27.700 144.900 27.900 ;
        RECT 145.400 27.400 145.700 28.500 ;
        RECT 147.500 28.000 147.900 28.800 ;
        RECT 151.800 28.500 152.200 29.500 ;
        RECT 153.900 29.200 154.300 29.500 ;
        RECT 153.400 28.800 154.300 29.200 ;
        RECT 147.500 27.700 148.300 28.000 ;
        RECT 147.900 27.500 148.300 27.700 ;
        RECT 144.200 27.200 144.600 27.400 ;
        RECT 142.200 26.800 143.500 27.200 ;
        RECT 144.200 26.900 145.000 27.200 ;
        RECT 145.400 27.100 147.500 27.400 ;
        RECT 144.600 26.800 145.000 26.900 ;
        RECT 147.000 26.900 147.500 27.100 ;
        RECT 148.000 27.200 148.300 27.500 ;
        RECT 151.800 27.400 152.100 28.500 ;
        RECT 153.900 28.000 154.300 28.800 ;
        RECT 153.900 27.700 154.700 28.000 ;
        RECT 154.300 27.500 154.700 27.700 ;
        RECT 139.700 25.400 141.800 25.700 ;
        RECT 138.200 24.900 139.400 25.200 ;
        RECT 137.900 24.500 138.300 24.600 ;
        RECT 137.200 24.200 138.300 24.500 ;
        RECT 139.100 24.400 139.400 24.900 ;
        RECT 139.100 24.000 139.800 24.400 ;
        RECT 135.900 23.700 136.300 23.800 ;
        RECT 137.300 23.700 137.700 23.800 ;
        RECT 134.200 23.100 134.600 23.500 ;
        RECT 135.900 23.400 137.700 23.700 ;
        RECT 137.000 23.100 137.300 23.400 ;
        RECT 139.000 23.100 139.400 23.500 ;
        RECT 134.200 22.800 135.200 23.100 ;
        RECT 134.800 21.100 135.200 22.800 ;
        RECT 137.000 21.100 137.400 23.100 ;
        RECT 139.100 21.100 139.700 23.100 ;
        RECT 141.400 21.100 141.800 25.400 ;
        RECT 142.200 25.100 142.600 25.200 ;
        RECT 143.200 25.100 143.500 26.800 ;
        RECT 143.800 25.800 144.200 26.600 ;
        RECT 145.400 25.800 145.800 26.600 ;
        RECT 146.200 25.800 146.600 26.600 ;
        RECT 147.000 26.500 147.700 26.900 ;
        RECT 148.000 26.800 149.000 27.200 ;
        RECT 151.800 27.100 153.900 27.400 ;
        RECT 153.400 26.900 153.900 27.100 ;
        RECT 154.400 27.200 154.700 27.500 ;
        RECT 156.600 27.600 157.000 29.900 ;
        RECT 158.200 28.200 158.600 29.900 ;
        RECT 161.100 28.200 161.500 29.900 ;
        RECT 158.200 27.900 158.700 28.200 ;
        RECT 156.600 27.300 157.900 27.600 ;
        RECT 147.000 25.500 147.300 26.500 ;
        RECT 145.400 25.200 147.300 25.500 ;
        RECT 142.200 24.800 142.900 25.100 ;
        RECT 143.200 24.800 143.700 25.100 ;
        RECT 142.600 24.200 142.900 24.800 ;
        RECT 142.600 23.800 143.000 24.200 ;
        RECT 143.300 21.100 143.700 24.800 ;
        RECT 145.400 23.500 145.700 25.200 ;
        RECT 148.000 24.900 148.300 26.800 ;
        RECT 148.600 25.400 149.000 26.200 ;
        RECT 151.800 25.800 152.200 26.600 ;
        RECT 152.600 25.800 153.000 26.600 ;
        RECT 153.400 26.500 154.100 26.900 ;
        RECT 154.400 26.800 155.400 27.200 ;
        RECT 153.400 25.500 153.700 26.500 ;
        RECT 147.500 24.600 148.300 24.900 ;
        RECT 151.800 25.200 153.700 25.500 ;
        RECT 145.400 21.500 145.800 23.500 ;
        RECT 147.500 21.100 147.900 24.600 ;
        RECT 151.800 23.500 152.100 25.200 ;
        RECT 154.400 24.900 154.700 26.800 ;
        RECT 156.700 26.200 157.100 26.600 ;
        RECT 155.000 25.400 155.400 26.200 ;
        RECT 155.800 26.100 156.200 26.200 ;
        RECT 156.600 26.100 157.100 26.200 ;
        RECT 155.800 25.800 157.100 26.100 ;
        RECT 157.600 26.500 157.900 27.300 ;
        RECT 158.400 27.200 158.700 27.900 ;
        RECT 160.600 27.900 161.500 28.200 ;
        RECT 162.200 27.900 162.600 29.900 ;
        RECT 163.000 28.000 163.400 29.900 ;
        RECT 164.600 28.000 165.000 29.900 ;
        RECT 163.000 27.900 165.000 28.000 ;
        RECT 158.200 26.800 158.700 27.200 ;
        RECT 159.800 27.100 160.200 27.600 ;
        RECT 157.600 26.100 158.100 26.500 ;
        RECT 157.600 25.100 157.900 26.100 ;
        RECT 158.400 25.100 158.700 26.800 ;
        RECT 159.000 26.800 160.200 27.100 ;
        RECT 159.000 26.200 159.300 26.800 ;
        RECT 159.000 25.800 159.400 26.200 ;
        RECT 160.600 26.100 161.000 27.900 ;
        RECT 162.300 27.200 162.600 27.900 ;
        RECT 163.100 27.700 164.900 27.900 ;
        RECT 165.400 27.600 165.800 29.900 ;
        RECT 167.000 28.200 167.400 29.900 ;
        RECT 167.000 27.900 167.500 28.200 ;
        RECT 168.600 27.900 169.000 29.900 ;
        RECT 169.400 28.000 169.800 29.900 ;
        RECT 171.000 28.000 171.400 29.900 ;
        RECT 169.400 27.900 171.400 28.000 ;
        RECT 164.200 27.200 164.600 27.400 ;
        RECT 165.400 27.300 166.700 27.600 ;
        RECT 162.200 26.800 163.500 27.200 ;
        RECT 164.200 26.900 165.000 27.200 ;
        RECT 164.600 26.800 165.000 26.900 ;
        RECT 160.600 25.800 162.500 26.100 ;
        RECT 153.900 24.600 154.700 24.900 ;
        RECT 156.600 24.800 157.900 25.100 ;
        RECT 151.800 21.500 152.200 23.500 ;
        RECT 153.900 21.100 154.300 24.600 ;
        RECT 156.600 21.100 157.000 24.800 ;
        RECT 158.200 24.600 158.700 25.100 ;
        RECT 158.200 21.100 158.600 24.600 ;
        RECT 160.600 21.100 161.000 25.800 ;
        RECT 162.200 25.200 162.500 25.800 ;
        RECT 161.400 24.400 161.800 25.200 ;
        RECT 162.200 25.100 162.600 25.200 ;
        RECT 163.200 25.100 163.500 26.800 ;
        RECT 163.800 25.800 164.200 26.600 ;
        RECT 166.400 26.500 166.700 27.300 ;
        RECT 167.200 27.200 167.500 27.900 ;
        RECT 168.700 27.200 169.000 27.900 ;
        RECT 169.500 27.700 171.300 27.900 ;
        RECT 171.800 27.700 172.200 29.900 ;
        RECT 173.900 29.200 174.500 29.900 ;
        RECT 173.900 28.900 174.600 29.200 ;
        RECT 176.200 28.900 176.600 29.900 ;
        RECT 178.400 29.200 178.800 29.900 ;
        RECT 178.400 28.900 179.400 29.200 ;
        RECT 174.200 28.500 174.600 28.900 ;
        RECT 176.300 28.600 176.600 28.900 ;
        RECT 176.300 28.300 177.700 28.600 ;
        RECT 177.300 28.200 177.700 28.300 ;
        RECT 178.200 28.200 178.600 28.600 ;
        RECT 179.000 28.500 179.400 28.900 ;
        RECT 173.300 27.700 173.700 27.800 ;
        RECT 171.800 27.400 173.700 27.700 ;
        RECT 170.600 27.200 171.000 27.400 ;
        RECT 167.000 26.800 167.500 27.200 ;
        RECT 168.600 26.800 169.900 27.200 ;
        RECT 170.600 26.900 171.400 27.200 ;
        RECT 171.000 26.800 171.400 26.900 ;
        RECT 166.400 26.100 166.900 26.500 ;
        RECT 166.400 25.100 166.700 26.100 ;
        RECT 167.200 25.100 167.500 26.800 ;
        RECT 167.800 26.100 168.200 26.200 ;
        RECT 167.800 25.800 168.900 26.100 ;
        RECT 162.200 24.800 162.900 25.100 ;
        RECT 163.200 24.800 163.700 25.100 ;
        RECT 162.600 24.200 162.900 24.800 ;
        RECT 162.600 23.800 163.000 24.200 ;
        RECT 163.300 21.100 163.700 24.800 ;
        RECT 165.400 24.800 166.700 25.100 ;
        RECT 165.400 21.100 165.800 24.800 ;
        RECT 167.000 24.600 167.500 25.100 ;
        RECT 168.600 25.200 168.900 25.800 ;
        RECT 168.600 25.100 169.000 25.200 ;
        RECT 169.600 25.100 169.900 26.800 ;
        RECT 170.200 25.800 170.600 26.600 ;
        RECT 171.800 25.700 172.200 27.400 ;
        RECT 175.300 27.100 175.700 27.200 ;
        RECT 176.600 27.100 177.000 27.200 ;
        RECT 178.200 27.100 178.500 28.200 ;
        RECT 180.600 27.500 181.000 29.900 ;
        RECT 182.700 28.200 183.100 29.900 ;
        RECT 182.200 27.900 183.100 28.200 ;
        RECT 183.800 27.900 184.200 29.900 ;
        RECT 184.600 28.000 185.000 29.900 ;
        RECT 186.200 28.000 186.600 29.900 ;
        RECT 184.600 27.900 186.600 28.000 ;
        RECT 179.800 27.100 180.600 27.200 ;
        RECT 175.100 26.800 180.600 27.100 ;
        RECT 181.400 26.800 181.800 27.600 ;
        RECT 174.200 26.400 174.600 26.500 ;
        RECT 172.700 26.100 174.600 26.400 ;
        RECT 172.700 26.000 173.100 26.100 ;
        RECT 173.500 25.700 173.900 25.800 ;
        RECT 171.800 25.400 173.900 25.700 ;
        RECT 168.600 24.800 169.300 25.100 ;
        RECT 169.600 24.800 170.100 25.100 ;
        RECT 167.000 21.100 167.400 24.600 ;
        RECT 169.000 24.200 169.300 24.800 ;
        RECT 169.000 23.800 169.400 24.200 ;
        RECT 169.700 21.100 170.100 24.800 ;
        RECT 171.800 21.100 172.200 25.400 ;
        RECT 175.100 25.200 175.400 26.800 ;
        RECT 178.700 26.700 179.100 26.800 ;
        RECT 179.500 26.200 179.900 26.300 ;
        RECT 177.400 25.900 179.900 26.200 ;
        RECT 182.200 26.100 182.600 27.900 ;
        RECT 183.900 27.200 184.200 27.900 ;
        RECT 184.700 27.700 186.500 27.900 ;
        RECT 187.000 27.700 187.400 29.900 ;
        RECT 189.100 29.200 189.700 29.900 ;
        RECT 189.100 28.900 189.800 29.200 ;
        RECT 191.400 28.900 191.800 29.900 ;
        RECT 193.600 29.200 194.000 29.900 ;
        RECT 193.600 28.900 194.600 29.200 ;
        RECT 189.400 28.500 189.800 28.900 ;
        RECT 191.500 28.600 191.800 28.900 ;
        RECT 191.500 28.300 192.900 28.600 ;
        RECT 192.500 28.200 192.900 28.300 ;
        RECT 193.400 28.200 193.800 28.600 ;
        RECT 194.200 28.500 194.600 28.900 ;
        RECT 188.500 27.700 188.900 27.800 ;
        RECT 187.000 27.400 188.900 27.700 ;
        RECT 185.800 27.200 186.200 27.400 ;
        RECT 183.800 26.800 185.100 27.200 ;
        RECT 185.800 26.900 186.600 27.200 ;
        RECT 186.200 26.800 186.600 26.900 ;
        RECT 177.400 25.800 177.800 25.900 ;
        RECT 182.200 25.800 184.100 26.100 ;
        RECT 178.200 25.500 181.000 25.600 ;
        RECT 178.100 25.400 181.000 25.500 ;
        RECT 174.200 24.900 175.400 25.200 ;
        RECT 176.100 25.300 181.000 25.400 ;
        RECT 176.100 25.100 178.500 25.300 ;
        RECT 174.200 24.400 174.500 24.900 ;
        RECT 173.800 24.000 174.500 24.400 ;
        RECT 175.300 24.500 175.700 24.600 ;
        RECT 176.100 24.500 176.400 25.100 ;
        RECT 175.300 24.200 176.400 24.500 ;
        RECT 176.700 24.500 179.400 24.800 ;
        RECT 176.700 24.400 177.100 24.500 ;
        RECT 179.000 24.400 179.400 24.500 ;
        RECT 175.900 23.700 176.300 23.800 ;
        RECT 177.300 23.700 177.700 23.800 ;
        RECT 174.200 23.100 174.600 23.500 ;
        RECT 175.900 23.400 177.700 23.700 ;
        RECT 176.300 23.100 176.600 23.400 ;
        RECT 179.000 23.100 179.400 23.500 ;
        RECT 173.900 21.100 174.500 23.100 ;
        RECT 176.200 21.100 176.600 23.100 ;
        RECT 178.400 22.800 179.400 23.100 ;
        RECT 178.400 21.100 178.800 22.800 ;
        RECT 180.600 21.100 181.000 25.300 ;
        RECT 182.200 21.100 182.600 25.800 ;
        RECT 183.800 25.200 184.100 25.800 ;
        RECT 184.800 25.200 185.100 26.800 ;
        RECT 185.400 25.800 185.800 26.600 ;
        RECT 187.000 25.700 187.400 27.400 ;
        RECT 190.500 27.100 190.900 27.200 ;
        RECT 193.400 27.100 193.700 28.200 ;
        RECT 195.800 27.500 196.200 29.900 ;
        RECT 196.600 28.500 197.000 29.500 ;
        RECT 198.700 29.200 199.100 29.500 ;
        RECT 198.200 28.800 199.100 29.200 ;
        RECT 196.600 27.400 196.900 28.500 ;
        RECT 198.700 28.000 199.100 28.800 ;
        RECT 198.700 27.700 199.500 28.000 ;
        RECT 199.100 27.500 199.500 27.700 ;
        RECT 195.000 27.100 195.800 27.200 ;
        RECT 196.600 27.100 198.700 27.400 ;
        RECT 190.300 26.800 195.800 27.100 ;
        RECT 198.200 26.900 198.700 27.100 ;
        RECT 199.200 27.200 199.500 27.500 ;
        RECT 203.000 27.600 203.400 29.900 ;
        RECT 204.600 28.200 205.000 29.900 ;
        RECT 207.500 28.200 207.900 29.900 ;
        RECT 204.600 27.900 205.100 28.200 ;
        RECT 203.000 27.300 204.300 27.600 ;
        RECT 189.400 26.400 189.800 26.500 ;
        RECT 187.900 26.100 189.800 26.400 ;
        RECT 190.300 26.200 190.600 26.800 ;
        RECT 193.900 26.700 194.300 26.800 ;
        RECT 194.700 26.200 195.100 26.300 ;
        RECT 187.900 26.000 188.300 26.100 ;
        RECT 190.200 25.800 190.600 26.200 ;
        RECT 192.600 25.900 195.100 26.200 ;
        RECT 192.600 25.800 193.000 25.900 ;
        RECT 196.600 25.800 197.000 26.600 ;
        RECT 197.400 25.800 197.800 26.600 ;
        RECT 198.200 26.500 198.900 26.900 ;
        RECT 199.200 26.800 200.200 27.200 ;
        RECT 188.700 25.700 189.100 25.800 ;
        RECT 187.000 25.400 189.100 25.700 ;
        RECT 183.000 24.400 183.400 25.200 ;
        RECT 183.800 25.100 184.200 25.200 ;
        RECT 183.800 24.800 184.500 25.100 ;
        RECT 184.800 24.800 185.800 25.200 ;
        RECT 184.200 24.200 184.500 24.800 ;
        RECT 184.200 23.800 184.600 24.200 ;
        RECT 184.900 21.100 185.300 24.800 ;
        RECT 187.000 21.100 187.400 25.400 ;
        RECT 190.300 25.200 190.600 25.800 ;
        RECT 193.400 25.500 196.200 25.600 ;
        RECT 198.200 25.500 198.500 26.500 ;
        RECT 193.300 25.400 196.200 25.500 ;
        RECT 189.400 24.900 190.600 25.200 ;
        RECT 191.300 25.300 196.200 25.400 ;
        RECT 191.300 25.100 193.700 25.300 ;
        RECT 189.400 24.400 189.700 24.900 ;
        RECT 189.000 24.000 189.700 24.400 ;
        RECT 190.500 24.500 190.900 24.600 ;
        RECT 191.300 24.500 191.600 25.100 ;
        RECT 190.500 24.200 191.600 24.500 ;
        RECT 191.900 24.500 194.600 24.800 ;
        RECT 191.900 24.400 192.300 24.500 ;
        RECT 194.200 24.400 194.600 24.500 ;
        RECT 191.100 23.700 191.500 23.800 ;
        RECT 192.500 23.700 192.900 23.800 ;
        RECT 189.400 23.100 189.800 23.500 ;
        RECT 191.100 23.400 192.900 23.700 ;
        RECT 191.500 23.100 191.800 23.400 ;
        RECT 194.200 23.100 194.600 23.500 ;
        RECT 189.100 21.100 189.700 23.100 ;
        RECT 191.400 21.100 191.800 23.100 ;
        RECT 193.600 22.800 194.600 23.100 ;
        RECT 193.600 21.100 194.000 22.800 ;
        RECT 195.800 21.100 196.200 25.300 ;
        RECT 196.600 25.200 198.500 25.500 ;
        RECT 196.600 23.500 196.900 25.200 ;
        RECT 199.200 24.900 199.500 26.800 ;
        RECT 204.000 26.500 204.300 27.300 ;
        RECT 204.800 27.200 205.100 27.900 ;
        RECT 207.000 27.900 207.900 28.200 ;
        RECT 208.600 27.900 209.000 29.900 ;
        RECT 209.400 28.000 209.800 29.900 ;
        RECT 211.000 28.000 211.400 29.900 ;
        RECT 209.400 27.900 211.400 28.000 ;
        RECT 211.800 28.000 212.200 29.900 ;
        RECT 213.400 28.000 213.800 29.900 ;
        RECT 211.800 27.900 213.800 28.000 ;
        RECT 214.200 27.900 214.600 29.900 ;
        RECT 215.800 28.200 216.200 29.900 ;
        RECT 215.700 27.900 216.200 28.200 ;
        RECT 204.600 26.800 205.100 27.200 ;
        RECT 205.400 27.100 205.800 27.200 ;
        RECT 206.200 27.100 206.600 27.600 ;
        RECT 205.400 26.800 206.600 27.100 ;
        RECT 199.800 25.400 200.200 26.200 ;
        RECT 204.000 26.100 204.500 26.500 ;
        RECT 204.000 25.100 204.300 26.100 ;
        RECT 204.800 25.100 205.100 26.800 ;
        RECT 198.700 24.600 199.500 24.900 ;
        RECT 203.000 24.800 204.300 25.100 ;
        RECT 196.600 21.500 197.000 23.500 ;
        RECT 198.700 21.100 199.100 24.600 ;
        RECT 203.000 21.100 203.400 24.800 ;
        RECT 204.600 24.600 205.100 25.100 ;
        RECT 207.000 26.100 207.400 27.900 ;
        RECT 208.700 27.200 209.000 27.900 ;
        RECT 209.500 27.700 211.300 27.900 ;
        RECT 211.900 27.700 213.700 27.900 ;
        RECT 210.600 27.200 211.000 27.400 ;
        RECT 212.200 27.200 212.600 27.400 ;
        RECT 214.200 27.200 214.500 27.900 ;
        RECT 215.700 27.200 216.000 27.900 ;
        RECT 217.400 27.600 217.800 29.900 ;
        RECT 216.500 27.300 217.800 27.600 ;
        RECT 218.200 27.700 218.600 29.900 ;
        RECT 220.300 29.200 220.900 29.900 ;
        RECT 220.300 28.900 221.000 29.200 ;
        RECT 222.600 28.900 223.000 29.900 ;
        RECT 224.800 29.200 225.200 29.900 ;
        RECT 224.800 28.900 225.800 29.200 ;
        RECT 220.600 28.500 221.000 28.900 ;
        RECT 222.700 28.600 223.000 28.900 ;
        RECT 222.700 28.300 224.100 28.600 ;
        RECT 223.700 28.200 224.100 28.300 ;
        RECT 224.600 28.200 225.000 28.600 ;
        RECT 225.400 28.500 225.800 28.900 ;
        RECT 219.700 27.700 220.100 27.800 ;
        RECT 218.200 27.400 220.100 27.700 ;
        RECT 208.600 26.800 209.900 27.200 ;
        RECT 210.600 27.100 211.400 27.200 ;
        RECT 211.800 27.100 212.600 27.200 ;
        RECT 210.600 26.900 212.600 27.100 ;
        RECT 211.000 26.800 212.200 26.900 ;
        RECT 213.300 26.800 214.600 27.200 ;
        RECT 215.000 27.100 215.400 27.200 ;
        RECT 215.700 27.100 216.200 27.200 ;
        RECT 215.000 26.800 216.200 27.100 ;
        RECT 207.000 25.800 208.900 26.100 ;
        RECT 204.600 21.100 205.000 24.600 ;
        RECT 207.000 21.100 207.400 25.800 ;
        RECT 208.600 25.200 208.900 25.800 ;
        RECT 207.800 24.400 208.200 25.200 ;
        RECT 208.600 25.100 209.000 25.200 ;
        RECT 209.600 25.100 209.900 26.800 ;
        RECT 210.200 25.800 210.600 26.600 ;
        RECT 212.600 25.800 213.000 26.600 ;
        RECT 213.300 26.100 213.600 26.800 ;
        RECT 215.000 26.100 215.400 26.200 ;
        RECT 213.300 25.800 215.400 26.100 ;
        RECT 213.300 25.100 213.600 25.800 ;
        RECT 214.200 25.100 214.600 25.200 ;
        RECT 208.600 24.800 209.300 25.100 ;
        RECT 209.600 24.800 210.100 25.100 ;
        RECT 209.000 24.200 209.300 24.800 ;
        RECT 209.000 23.800 209.400 24.200 ;
        RECT 209.700 21.100 210.100 24.800 ;
        RECT 213.100 24.800 213.600 25.100 ;
        RECT 213.900 24.800 214.600 25.100 ;
        RECT 215.700 25.100 216.000 26.800 ;
        RECT 216.500 26.500 216.800 27.300 ;
        RECT 216.300 26.100 216.800 26.500 ;
        RECT 216.500 25.100 216.800 26.100 ;
        RECT 217.300 26.200 217.700 26.600 ;
        RECT 217.300 25.800 217.800 26.200 ;
        RECT 218.200 25.700 218.600 27.400 ;
        RECT 221.700 27.100 222.100 27.200 ;
        RECT 224.600 27.100 224.900 28.200 ;
        RECT 227.000 27.500 227.400 29.900 ;
        RECT 229.100 29.200 229.500 29.900 ;
        RECT 228.600 28.800 229.500 29.200 ;
        RECT 229.100 28.200 229.500 28.800 ;
        RECT 228.600 27.900 229.500 28.200 ;
        RECT 226.200 27.100 227.000 27.200 ;
        RECT 221.500 26.800 227.000 27.100 ;
        RECT 227.800 26.800 228.200 27.600 ;
        RECT 220.600 26.400 221.000 26.500 ;
        RECT 219.100 26.100 221.000 26.400 ;
        RECT 221.500 26.100 221.800 26.800 ;
        RECT 225.100 26.700 225.500 26.800 ;
        RECT 225.900 26.200 226.300 26.300 ;
        RECT 222.200 26.100 222.600 26.200 ;
        RECT 219.100 26.000 219.500 26.100 ;
        RECT 221.400 25.800 222.600 26.100 ;
        RECT 223.800 25.900 226.300 26.200 ;
        RECT 223.800 25.800 224.200 25.900 ;
        RECT 219.900 25.700 220.300 25.800 ;
        RECT 218.200 25.400 220.300 25.700 ;
        RECT 213.100 21.100 213.500 24.800 ;
        RECT 213.900 24.200 214.200 24.800 ;
        RECT 215.700 24.600 216.200 25.100 ;
        RECT 216.500 24.800 217.800 25.100 ;
        RECT 213.800 23.800 214.200 24.200 ;
        RECT 215.800 21.100 216.200 24.600 ;
        RECT 217.400 21.100 217.800 24.800 ;
        RECT 218.200 21.100 218.600 25.400 ;
        RECT 221.500 25.200 221.800 25.800 ;
        RECT 224.600 25.500 227.400 25.600 ;
        RECT 224.500 25.400 227.400 25.500 ;
        RECT 220.600 24.900 221.800 25.200 ;
        RECT 222.500 25.300 227.400 25.400 ;
        RECT 222.500 25.100 224.900 25.300 ;
        RECT 220.600 24.400 220.900 24.900 ;
        RECT 220.200 24.000 220.900 24.400 ;
        RECT 221.700 24.500 222.100 24.600 ;
        RECT 222.500 24.500 222.800 25.100 ;
        RECT 221.700 24.200 222.800 24.500 ;
        RECT 223.100 24.500 225.800 24.800 ;
        RECT 223.100 24.400 223.500 24.500 ;
        RECT 225.400 24.400 225.800 24.500 ;
        RECT 222.300 23.700 222.700 23.800 ;
        RECT 223.700 23.700 224.100 23.800 ;
        RECT 220.600 23.100 221.000 23.500 ;
        RECT 222.300 23.400 224.100 23.700 ;
        RECT 222.700 23.100 223.000 23.400 ;
        RECT 225.400 23.100 225.800 23.500 ;
        RECT 220.300 21.100 220.900 23.100 ;
        RECT 222.600 21.100 223.000 23.100 ;
        RECT 224.800 22.800 225.800 23.100 ;
        RECT 224.800 21.100 225.200 22.800 ;
        RECT 227.000 21.100 227.400 25.300 ;
        RECT 228.600 21.100 229.000 27.900 ;
        RECT 230.200 27.700 230.600 29.900 ;
        RECT 232.300 29.200 232.900 29.900 ;
        RECT 232.300 28.900 233.000 29.200 ;
        RECT 234.600 28.900 235.000 29.900 ;
        RECT 236.800 29.200 237.200 29.900 ;
        RECT 236.800 28.900 237.800 29.200 ;
        RECT 232.600 28.500 233.000 28.900 ;
        RECT 234.700 28.600 235.000 28.900 ;
        RECT 234.700 28.300 236.100 28.600 ;
        RECT 235.700 28.200 236.100 28.300 ;
        RECT 236.600 28.200 237.000 28.600 ;
        RECT 237.400 28.500 237.800 28.900 ;
        RECT 231.700 27.700 232.100 27.800 ;
        RECT 230.200 27.400 232.100 27.700 ;
        RECT 230.200 25.700 230.600 27.400 ;
        RECT 236.600 27.200 236.900 28.200 ;
        RECT 239.000 27.500 239.400 29.900 ;
        RECT 239.800 27.700 240.200 29.900 ;
        RECT 241.900 29.200 242.500 29.900 ;
        RECT 241.900 28.900 242.600 29.200 ;
        RECT 244.200 28.900 244.600 29.900 ;
        RECT 246.400 29.200 246.800 29.900 ;
        RECT 246.400 28.900 247.400 29.200 ;
        RECT 242.200 28.500 242.600 28.900 ;
        RECT 244.300 28.600 244.600 28.900 ;
        RECT 244.300 28.300 245.700 28.600 ;
        RECT 245.300 28.200 245.700 28.300 ;
        RECT 246.200 27.800 246.600 28.600 ;
        RECT 247.000 28.500 247.400 28.900 ;
        RECT 241.300 27.700 241.700 27.800 ;
        RECT 239.800 27.400 241.700 27.700 ;
        RECT 233.700 27.100 234.100 27.200 ;
        RECT 236.600 27.100 237.000 27.200 ;
        RECT 238.200 27.100 239.000 27.200 ;
        RECT 233.500 26.800 239.000 27.100 ;
        RECT 232.600 26.400 233.000 26.500 ;
        RECT 231.100 26.100 233.000 26.400 ;
        RECT 231.100 26.000 231.500 26.100 ;
        RECT 231.900 25.700 232.300 25.800 ;
        RECT 230.200 25.400 232.300 25.700 ;
        RECT 229.400 24.400 229.800 25.200 ;
        RECT 230.200 21.100 230.600 25.400 ;
        RECT 233.500 25.200 233.800 26.800 ;
        RECT 237.100 26.700 237.500 26.800 ;
        RECT 237.900 26.200 238.300 26.300 ;
        RECT 235.800 25.900 238.300 26.200 ;
        RECT 235.800 25.800 236.200 25.900 ;
        RECT 239.800 25.700 240.200 27.400 ;
        RECT 243.300 27.100 243.700 27.200 ;
        RECT 246.200 27.100 246.500 27.800 ;
        RECT 248.600 27.500 249.000 29.900 ;
        RECT 249.400 28.000 249.800 29.900 ;
        RECT 251.000 28.000 251.400 29.900 ;
        RECT 249.400 27.900 251.400 28.000 ;
        RECT 251.800 27.900 252.200 29.900 ;
        RECT 249.500 27.700 251.300 27.900 ;
        RECT 249.800 27.200 250.200 27.400 ;
        RECT 251.800 27.200 252.100 27.900 ;
        RECT 247.800 27.100 248.600 27.200 ;
        RECT 243.100 26.800 248.600 27.100 ;
        RECT 249.400 26.900 250.200 27.200 ;
        RECT 249.400 26.800 249.800 26.900 ;
        RECT 250.900 26.800 252.200 27.200 ;
        RECT 242.200 26.400 242.600 26.500 ;
        RECT 240.700 26.100 242.600 26.400 ;
        RECT 243.100 26.100 243.400 26.800 ;
        RECT 246.700 26.700 247.100 26.800 ;
        RECT 247.500 26.200 247.900 26.300 ;
        RECT 243.800 26.100 244.200 26.200 ;
        RECT 240.700 26.000 241.100 26.100 ;
        RECT 243.000 25.800 244.200 26.100 ;
        RECT 245.400 25.900 247.900 26.200 ;
        RECT 245.400 25.800 245.800 25.900 ;
        RECT 250.200 25.800 250.600 26.600 ;
        RECT 241.500 25.700 241.900 25.800 ;
        RECT 236.600 25.500 239.400 25.600 ;
        RECT 236.500 25.400 239.400 25.500 ;
        RECT 232.600 24.900 233.800 25.200 ;
        RECT 234.500 25.300 239.400 25.400 ;
        RECT 234.500 25.100 236.900 25.300 ;
        RECT 232.600 24.400 232.900 24.900 ;
        RECT 232.200 24.000 232.900 24.400 ;
        RECT 233.700 24.500 234.100 24.600 ;
        RECT 234.500 24.500 234.800 25.100 ;
        RECT 233.700 24.200 234.800 24.500 ;
        RECT 235.100 24.500 237.800 24.800 ;
        RECT 235.100 24.400 235.500 24.500 ;
        RECT 237.400 24.400 237.800 24.500 ;
        RECT 234.300 23.700 234.700 23.800 ;
        RECT 235.700 23.700 236.100 23.800 ;
        RECT 232.600 23.100 233.000 23.500 ;
        RECT 234.300 23.400 236.100 23.700 ;
        RECT 234.700 23.100 235.000 23.400 ;
        RECT 237.400 23.100 237.800 23.500 ;
        RECT 232.300 21.100 232.900 23.100 ;
        RECT 234.600 21.100 235.000 23.100 ;
        RECT 236.800 22.800 237.800 23.100 ;
        RECT 236.800 21.100 237.200 22.800 ;
        RECT 239.000 21.100 239.400 25.300 ;
        RECT 239.800 25.400 241.900 25.700 ;
        RECT 239.800 21.100 240.200 25.400 ;
        RECT 243.100 25.200 243.400 25.800 ;
        RECT 246.200 25.500 249.000 25.600 ;
        RECT 246.100 25.400 249.000 25.500 ;
        RECT 242.200 24.900 243.400 25.200 ;
        RECT 244.100 25.300 249.000 25.400 ;
        RECT 244.100 25.100 246.500 25.300 ;
        RECT 242.200 24.400 242.500 24.900 ;
        RECT 241.800 24.000 242.500 24.400 ;
        RECT 243.300 24.500 243.700 24.600 ;
        RECT 244.100 24.500 244.400 25.100 ;
        RECT 243.300 24.200 244.400 24.500 ;
        RECT 244.700 24.500 247.400 24.800 ;
        RECT 244.700 24.400 245.100 24.500 ;
        RECT 247.000 24.400 247.400 24.500 ;
        RECT 243.900 23.700 244.300 23.800 ;
        RECT 245.300 23.700 245.700 23.800 ;
        RECT 242.200 23.100 242.600 23.500 ;
        RECT 243.900 23.400 245.700 23.700 ;
        RECT 244.300 23.100 244.600 23.400 ;
        RECT 247.000 23.100 247.400 23.500 ;
        RECT 241.900 21.100 242.500 23.100 ;
        RECT 244.200 21.100 244.600 23.100 ;
        RECT 246.400 22.800 247.400 23.100 ;
        RECT 246.400 21.100 246.800 22.800 ;
        RECT 248.600 21.100 249.000 25.300 ;
        RECT 250.900 25.100 251.200 26.800 ;
        RECT 251.800 25.100 252.200 25.200 ;
        RECT 250.700 24.800 251.200 25.100 ;
        RECT 251.500 24.800 252.200 25.100 ;
        RECT 250.700 21.100 251.100 24.800 ;
        RECT 251.500 24.200 251.800 24.800 ;
        RECT 251.400 23.800 251.800 24.200 ;
        RECT 0.600 15.600 1.000 19.900 ;
        RECT 2.700 17.900 3.300 19.900 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.200 18.200 7.600 19.900 ;
        RECT 7.200 17.900 8.200 18.200 ;
        RECT 3.000 17.500 3.400 17.900 ;
        RECT 5.100 17.600 5.400 17.900 ;
        RECT 4.700 17.300 6.500 17.600 ;
        RECT 7.800 17.500 8.200 17.900 ;
        RECT 4.700 17.200 5.100 17.300 ;
        RECT 6.100 17.200 6.500 17.300 ;
        RECT 2.600 16.600 3.300 17.000 ;
        RECT 3.000 16.100 3.300 16.600 ;
        RECT 4.100 16.500 5.200 16.800 ;
        RECT 4.100 16.400 4.500 16.500 ;
        RECT 3.000 15.800 4.200 16.100 ;
        RECT 0.600 15.300 2.700 15.600 ;
        RECT 0.600 13.600 1.000 15.300 ;
        RECT 2.300 15.200 2.700 15.300 ;
        RECT 1.500 14.900 1.900 15.000 ;
        RECT 1.500 14.600 3.400 14.900 ;
        RECT 3.000 14.500 3.400 14.600 ;
        RECT 3.900 14.200 4.200 15.800 ;
        RECT 4.900 15.900 5.200 16.500 ;
        RECT 5.500 16.500 5.900 16.600 ;
        RECT 7.800 16.500 8.200 16.600 ;
        RECT 5.500 16.200 8.200 16.500 ;
        RECT 4.900 15.700 7.300 15.900 ;
        RECT 9.400 15.700 9.800 19.900 ;
        RECT 4.900 15.600 9.800 15.700 ;
        RECT 6.900 15.500 9.800 15.600 ;
        RECT 7.000 15.400 9.800 15.500 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 11.000 15.100 11.400 19.900 ;
        RECT 13.000 16.800 13.400 17.200 ;
        RECT 11.800 15.800 12.200 16.600 ;
        RECT 13.000 16.200 13.300 16.800 ;
        RECT 13.700 16.200 14.100 19.900 ;
        RECT 12.600 15.900 13.300 16.200 ;
        RECT 13.600 15.900 14.100 16.200 ;
        RECT 12.600 15.800 13.000 15.900 ;
        RECT 12.600 15.100 12.900 15.800 ;
        RECT 6.200 14.800 8.700 15.100 ;
        RECT 7.000 14.700 7.400 14.800 ;
        RECT 8.300 14.700 8.700 14.800 ;
        RECT 11.000 14.800 12.900 15.100 ;
        RECT 7.500 14.200 7.900 14.300 ;
        RECT 3.900 13.900 9.400 14.200 ;
        RECT 4.100 13.800 4.500 13.900 ;
        RECT 0.600 13.300 2.500 13.600 ;
        RECT 0.600 11.100 1.000 13.300 ;
        RECT 2.100 13.200 2.500 13.300 ;
        RECT 7.000 13.200 7.300 13.900 ;
        RECT 8.600 13.800 9.400 13.900 ;
        RECT 6.100 12.700 6.500 12.800 ;
        RECT 3.000 12.100 3.400 12.500 ;
        RECT 5.100 12.400 6.500 12.700 ;
        RECT 7.000 12.400 7.400 13.200 ;
        RECT 5.100 12.100 5.400 12.400 ;
        RECT 7.800 12.100 8.200 12.500 ;
        RECT 2.700 11.800 3.400 12.100 ;
        RECT 2.700 11.100 3.300 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.200 11.800 8.200 12.100 ;
        RECT 7.200 11.100 7.600 11.800 ;
        RECT 9.400 11.100 9.800 13.500 ;
        RECT 10.200 13.400 10.600 14.200 ;
        RECT 11.000 13.100 11.400 14.800 ;
        RECT 13.600 14.200 13.900 15.900 ;
        RECT 15.800 15.800 16.200 16.600 ;
        RECT 14.200 14.400 14.600 15.200 ;
        RECT 12.600 13.800 13.900 14.200 ;
        RECT 15.000 14.100 15.400 14.200 ;
        RECT 14.600 13.800 15.400 14.100 ;
        RECT 12.700 13.100 13.000 13.800 ;
        RECT 14.600 13.600 15.000 13.800 ;
        RECT 13.500 13.100 15.300 13.300 ;
        RECT 16.600 13.100 17.000 19.900 ;
        RECT 18.200 16.200 18.600 19.900 ;
        RECT 19.800 16.200 20.200 19.900 ;
        RECT 18.200 15.900 20.200 16.200 ;
        RECT 20.600 15.900 21.000 19.900 ;
        RECT 21.700 16.300 22.100 19.900 ;
        RECT 21.700 15.900 22.600 16.300 ;
        RECT 18.600 15.200 19.000 15.400 ;
        RECT 20.600 15.200 20.900 15.900 ;
        RECT 17.400 15.100 17.800 15.200 ;
        RECT 18.200 15.100 19.000 15.200 ;
        RECT 17.400 14.900 19.000 15.100 ;
        RECT 19.800 14.900 21.000 15.200 ;
        RECT 17.400 14.800 18.600 14.900 ;
        RECT 17.400 13.400 17.800 14.200 ;
        RECT 19.000 13.800 19.400 14.600 ;
        RECT 11.000 12.800 11.900 13.100 ;
        RECT 11.500 11.100 11.900 12.800 ;
        RECT 12.600 11.100 13.000 13.100 ;
        RECT 13.400 13.000 15.400 13.100 ;
        RECT 13.400 11.100 13.800 13.000 ;
        RECT 15.000 11.100 15.400 13.000 ;
        RECT 16.100 12.800 17.000 13.100 ;
        RECT 19.800 13.100 20.100 14.900 ;
        RECT 20.600 14.800 21.000 14.900 ;
        RECT 21.400 14.800 21.800 15.600 ;
        RECT 20.600 14.200 20.900 14.800 ;
        RECT 22.200 14.200 22.500 15.900 ;
        RECT 23.800 15.700 24.200 19.900 ;
        RECT 26.000 18.200 26.400 19.900 ;
        RECT 25.400 17.900 26.400 18.200 ;
        RECT 28.200 17.900 28.600 19.900 ;
        RECT 30.300 17.900 30.900 19.900 ;
        RECT 25.400 17.500 25.800 17.900 ;
        RECT 28.200 17.600 28.500 17.900 ;
        RECT 27.100 17.300 28.900 17.600 ;
        RECT 30.200 17.500 30.600 17.900 ;
        RECT 27.100 17.200 27.500 17.300 ;
        RECT 28.500 17.200 28.900 17.300 ;
        RECT 25.400 16.500 25.800 16.600 ;
        RECT 27.700 16.500 28.100 16.600 ;
        RECT 25.400 16.200 28.100 16.500 ;
        RECT 28.400 16.500 29.500 16.800 ;
        RECT 28.400 15.900 28.700 16.500 ;
        RECT 29.100 16.400 29.500 16.500 ;
        RECT 30.300 16.600 31.000 17.000 ;
        RECT 30.300 16.100 30.600 16.600 ;
        RECT 26.300 15.700 28.700 15.900 ;
        RECT 23.800 15.600 28.700 15.700 ;
        RECT 29.400 15.800 30.600 16.100 ;
        RECT 23.800 15.500 26.700 15.600 ;
        RECT 23.800 15.400 26.600 15.500 ;
        RECT 27.000 15.100 27.400 15.200 ;
        RECT 24.900 14.800 27.400 15.100 ;
        RECT 24.900 14.700 25.300 14.800 ;
        RECT 26.200 14.700 26.600 14.800 ;
        RECT 25.700 14.200 26.100 14.300 ;
        RECT 29.400 14.200 29.700 15.800 ;
        RECT 32.600 15.600 33.000 19.900 ;
        RECT 30.900 15.300 33.000 15.600 ;
        RECT 30.900 15.200 31.300 15.300 ;
        RECT 31.700 14.900 32.100 15.000 ;
        RECT 30.200 14.600 32.100 14.900 ;
        RECT 30.200 14.500 30.600 14.600 ;
        RECT 20.600 13.800 21.000 14.200 ;
        RECT 22.200 13.800 22.600 14.200 ;
        RECT 24.200 13.900 29.700 14.200 ;
        RECT 24.200 13.800 25.000 13.900 ;
        RECT 20.600 13.100 21.000 13.200 ;
        RECT 22.200 13.100 22.500 13.800 ;
        RECT 16.100 12.200 16.500 12.800 ;
        RECT 16.100 11.800 17.000 12.200 ;
        RECT 16.100 11.100 16.500 11.800 ;
        RECT 19.800 11.100 20.200 13.100 ;
        RECT 20.600 12.800 22.500 13.100 ;
        RECT 20.500 12.400 20.900 12.800 ;
        RECT 22.200 12.100 22.500 12.800 ;
        RECT 23.000 12.400 23.400 13.200 ;
        RECT 22.200 11.100 22.600 12.100 ;
        RECT 23.800 11.100 24.200 13.500 ;
        RECT 26.300 12.800 26.600 13.900 ;
        RECT 29.100 13.800 29.500 13.900 ;
        RECT 32.600 13.600 33.000 15.300 ;
        RECT 34.200 15.600 34.600 19.900 ;
        RECT 35.800 15.600 36.200 19.900 ;
        RECT 37.400 15.600 37.800 19.900 ;
        RECT 39.000 15.600 39.400 19.900 ;
        RECT 41.400 15.600 41.800 19.900 ;
        RECT 43.000 15.600 43.400 19.900 ;
        RECT 46.500 19.200 46.900 19.900 ;
        RECT 46.500 18.800 47.400 19.200 ;
        RECT 46.500 16.400 46.900 18.800 ;
        RECT 48.600 17.500 49.000 19.500 ;
        RECT 46.100 16.100 46.900 16.400 ;
        RECT 34.200 15.200 35.100 15.600 ;
        RECT 35.800 15.200 36.900 15.600 ;
        RECT 37.400 15.200 38.500 15.600 ;
        RECT 39.000 15.200 40.200 15.600 ;
        RECT 34.700 14.500 35.100 15.200 ;
        RECT 36.500 14.500 36.900 15.200 ;
        RECT 38.100 14.500 38.500 15.200 ;
        RECT 33.400 14.100 34.300 14.500 ;
        RECT 34.700 14.100 36.000 14.500 ;
        RECT 36.500 14.100 37.700 14.500 ;
        RECT 38.100 14.100 39.400 14.500 ;
        RECT 33.400 13.800 33.800 14.100 ;
        RECT 34.700 13.800 35.100 14.100 ;
        RECT 36.500 13.800 36.900 14.100 ;
        RECT 38.100 13.800 38.500 14.100 ;
        RECT 39.800 13.800 40.200 15.200 ;
        RECT 31.100 13.300 33.000 13.600 ;
        RECT 31.100 13.200 31.500 13.300 ;
        RECT 25.400 12.100 25.800 12.500 ;
        RECT 26.200 12.400 26.600 12.800 ;
        RECT 27.100 12.700 27.500 12.800 ;
        RECT 27.100 12.400 28.500 12.700 ;
        RECT 28.200 12.100 28.500 12.400 ;
        RECT 30.200 12.100 30.600 12.500 ;
        RECT 25.400 11.800 26.400 12.100 ;
        RECT 26.000 11.100 26.400 11.800 ;
        RECT 28.200 11.100 28.600 12.100 ;
        RECT 30.200 11.800 30.900 12.100 ;
        RECT 30.300 11.100 30.900 11.800 ;
        RECT 32.600 11.100 33.000 13.300 ;
        RECT 34.200 13.400 35.100 13.800 ;
        RECT 35.800 13.400 36.900 13.800 ;
        RECT 37.400 13.400 38.500 13.800 ;
        RECT 39.000 13.400 40.200 13.800 ;
        RECT 41.400 15.200 43.400 15.600 ;
        RECT 41.400 13.800 41.800 15.200 ;
        RECT 44.600 15.100 45.000 15.200 ;
        RECT 45.400 15.100 45.800 15.600 ;
        RECT 44.600 14.800 45.800 15.100 ;
        RECT 46.100 14.200 46.400 16.100 ;
        RECT 48.700 15.800 49.000 17.500 ;
        RECT 51.000 16.200 51.400 19.900 ;
        RECT 51.000 15.900 52.100 16.200 ;
        RECT 47.100 15.500 49.000 15.800 ;
        RECT 51.800 15.600 52.100 15.900 ;
        RECT 54.200 15.600 54.600 19.900 ;
        RECT 55.800 15.600 56.200 19.900 ;
        RECT 57.400 15.600 57.800 19.900 ;
        RECT 59.000 15.600 59.400 19.900 ;
        RECT 47.100 14.500 47.400 15.500 ;
        RECT 51.800 15.200 52.400 15.600 ;
        RECT 54.200 15.200 55.100 15.600 ;
        RECT 55.800 15.200 56.900 15.600 ;
        RECT 57.400 15.200 58.500 15.600 ;
        RECT 59.000 15.200 60.200 15.600 ;
        RECT 45.400 13.800 46.400 14.200 ;
        RECT 46.700 14.100 47.400 14.500 ;
        RECT 47.800 14.400 48.200 15.200 ;
        RECT 48.600 14.400 49.000 15.200 ;
        RECT 51.000 14.400 51.400 15.200 ;
        RECT 41.400 13.400 43.400 13.800 ;
        RECT 34.200 11.100 34.600 13.400 ;
        RECT 35.800 11.100 36.200 13.400 ;
        RECT 37.400 11.100 37.800 13.400 ;
        RECT 39.000 11.100 39.400 13.400 ;
        RECT 41.400 11.100 41.800 13.400 ;
        RECT 43.000 11.100 43.400 13.400 ;
        RECT 46.100 13.500 46.400 13.800 ;
        RECT 46.900 13.900 47.400 14.100 ;
        RECT 46.900 13.600 49.000 13.900 ;
        RECT 51.800 13.700 52.100 15.200 ;
        RECT 54.700 14.500 55.100 15.200 ;
        RECT 56.500 14.500 56.900 15.200 ;
        RECT 58.100 14.500 58.500 15.200 ;
        RECT 53.400 14.100 54.300 14.500 ;
        RECT 54.700 14.100 56.000 14.500 ;
        RECT 56.500 14.100 57.700 14.500 ;
        RECT 58.100 14.100 59.400 14.500 ;
        RECT 53.400 13.800 53.800 14.100 ;
        RECT 54.700 13.800 55.100 14.100 ;
        RECT 56.500 13.800 56.900 14.100 ;
        RECT 58.100 13.800 58.500 14.100 ;
        RECT 59.800 13.800 60.200 15.200 ;
        RECT 61.400 15.100 61.800 19.900 ;
        RECT 63.400 16.800 63.800 17.200 ;
        RECT 62.200 15.800 62.600 16.600 ;
        RECT 63.400 16.200 63.700 16.800 ;
        RECT 64.100 16.200 64.500 19.900 ;
        RECT 68.100 19.200 68.500 19.900 ;
        RECT 67.800 18.800 68.500 19.200 ;
        RECT 68.100 16.400 68.500 18.800 ;
        RECT 70.200 17.500 70.600 19.500 ;
        RECT 63.000 15.900 63.700 16.200 ;
        RECT 64.000 15.900 64.500 16.200 ;
        RECT 67.700 16.100 68.500 16.400 ;
        RECT 63.000 15.800 63.400 15.900 ;
        RECT 63.000 15.100 63.300 15.800 ;
        RECT 61.400 14.800 63.300 15.100 ;
        RECT 46.100 13.300 46.500 13.500 ;
        RECT 46.100 13.000 46.900 13.300 ;
        RECT 46.500 11.500 46.900 13.000 ;
        RECT 48.700 12.500 49.000 13.600 ;
        RECT 48.600 11.500 49.000 12.500 ;
        RECT 51.000 13.400 52.100 13.700 ;
        RECT 54.200 13.400 55.100 13.800 ;
        RECT 55.800 13.400 56.900 13.800 ;
        RECT 57.400 13.400 58.500 13.800 ;
        RECT 59.000 13.400 60.200 13.800 ;
        RECT 60.600 13.400 61.000 14.200 ;
        RECT 51.000 11.100 51.400 13.400 ;
        RECT 54.200 11.100 54.600 13.400 ;
        RECT 55.800 11.100 56.200 13.400 ;
        RECT 57.400 11.100 57.800 13.400 ;
        RECT 59.000 11.100 59.400 13.400 ;
        RECT 61.400 13.100 61.800 14.800 ;
        RECT 64.000 14.200 64.300 15.900 ;
        RECT 64.600 14.400 65.000 15.200 ;
        RECT 65.400 15.100 65.800 15.200 ;
        RECT 67.000 15.100 67.400 15.600 ;
        RECT 65.400 14.800 67.400 15.100 ;
        RECT 67.700 14.200 68.000 16.100 ;
        RECT 70.300 15.800 70.600 17.500 ;
        RECT 68.700 15.500 70.600 15.800 ;
        RECT 71.000 15.700 71.400 19.900 ;
        RECT 73.200 18.200 73.600 19.900 ;
        RECT 72.600 17.900 73.600 18.200 ;
        RECT 75.400 17.900 75.800 19.900 ;
        RECT 77.500 17.900 78.100 19.900 ;
        RECT 72.600 17.500 73.000 17.900 ;
        RECT 75.400 17.600 75.700 17.900 ;
        RECT 74.300 17.300 76.100 17.600 ;
        RECT 77.400 17.500 77.800 17.900 ;
        RECT 74.300 17.200 74.700 17.300 ;
        RECT 75.700 17.200 76.100 17.300 ;
        RECT 77.900 17.000 78.600 17.200 ;
        RECT 77.500 16.800 78.600 17.000 ;
        RECT 79.800 17.100 80.200 19.900 ;
        RECT 80.600 17.100 81.000 17.200 ;
        RECT 79.800 16.800 81.000 17.100 ;
        RECT 72.600 16.500 73.000 16.600 ;
        RECT 74.900 16.500 75.300 16.600 ;
        RECT 72.600 16.200 75.300 16.500 ;
        RECT 75.600 16.500 76.700 16.800 ;
        RECT 75.600 15.900 75.900 16.500 ;
        RECT 76.300 16.400 76.700 16.500 ;
        RECT 77.500 16.600 78.200 16.800 ;
        RECT 77.500 16.100 77.800 16.600 ;
        RECT 73.500 15.700 75.900 15.900 ;
        RECT 71.000 15.600 75.900 15.700 ;
        RECT 76.600 15.800 77.800 16.100 ;
        RECT 71.000 15.500 73.900 15.600 ;
        RECT 68.700 14.500 69.000 15.500 ;
        RECT 71.000 15.400 73.800 15.500 ;
        RECT 63.000 13.800 64.300 14.200 ;
        RECT 65.400 14.100 65.800 14.200 ;
        RECT 65.000 13.800 65.800 14.100 ;
        RECT 67.000 13.800 68.000 14.200 ;
        RECT 68.300 14.100 69.000 14.500 ;
        RECT 69.400 14.400 69.800 15.200 ;
        RECT 70.200 14.400 70.600 15.200 ;
        RECT 74.200 15.100 74.600 15.200 ;
        RECT 72.100 14.800 74.600 15.100 ;
        RECT 72.100 14.700 72.500 14.800 ;
        RECT 72.900 14.200 73.300 14.300 ;
        RECT 76.600 14.200 76.900 15.800 ;
        RECT 79.800 15.600 80.200 16.800 ;
        RECT 78.100 15.300 80.200 15.600 ;
        RECT 78.100 15.200 78.500 15.300 ;
        RECT 78.900 14.900 79.300 15.000 ;
        RECT 77.400 14.600 79.300 14.900 ;
        RECT 77.400 14.500 77.800 14.600 ;
        RECT 63.100 13.100 63.400 13.800 ;
        RECT 65.000 13.600 65.400 13.800 ;
        RECT 67.700 13.500 68.000 13.800 ;
        RECT 68.500 13.900 69.000 14.100 ;
        RECT 71.400 13.900 76.900 14.200 ;
        RECT 68.500 13.600 70.600 13.900 ;
        RECT 71.400 13.800 72.200 13.900 ;
        RECT 67.700 13.300 68.100 13.500 ;
        RECT 63.900 13.100 65.700 13.300 ;
        RECT 61.400 12.800 62.300 13.100 ;
        RECT 61.900 11.100 62.300 12.800 ;
        RECT 63.000 11.100 63.400 13.100 ;
        RECT 63.800 13.000 65.800 13.100 ;
        RECT 67.700 13.000 68.500 13.300 ;
        RECT 63.800 11.100 64.200 13.000 ;
        RECT 65.400 11.100 65.800 13.000 ;
        RECT 68.100 11.500 68.500 13.000 ;
        RECT 70.300 12.500 70.600 13.600 ;
        RECT 70.200 11.500 70.600 12.500 ;
        RECT 71.000 11.100 71.400 13.500 ;
        RECT 73.500 12.800 73.800 13.900 ;
        RECT 76.300 13.800 76.700 13.900 ;
        RECT 79.800 13.600 80.200 15.300 ;
        RECT 81.400 15.100 81.800 19.900 ;
        RECT 83.400 16.800 83.800 17.200 ;
        RECT 82.200 15.800 82.600 16.600 ;
        RECT 83.400 16.200 83.700 16.800 ;
        RECT 84.100 16.200 84.500 19.900 ;
        RECT 83.000 15.900 83.700 16.200 ;
        RECT 84.000 15.900 84.500 16.200 ;
        RECT 83.000 15.800 83.400 15.900 ;
        RECT 83.000 15.100 83.300 15.800 ;
        RECT 81.400 14.800 83.300 15.100 ;
        RECT 78.300 13.300 80.200 13.600 ;
        RECT 80.600 13.400 81.000 14.200 ;
        RECT 78.300 13.200 78.700 13.300 ;
        RECT 72.600 12.100 73.000 12.500 ;
        RECT 73.400 12.400 73.800 12.800 ;
        RECT 74.300 12.700 74.700 12.800 ;
        RECT 74.300 12.400 75.700 12.700 ;
        RECT 75.400 12.100 75.700 12.400 ;
        RECT 77.400 12.100 77.800 12.500 ;
        RECT 72.600 11.800 73.600 12.100 ;
        RECT 73.200 11.100 73.600 11.800 ;
        RECT 75.400 11.100 75.800 12.100 ;
        RECT 77.400 11.800 78.100 12.100 ;
        RECT 77.500 11.100 78.100 11.800 ;
        RECT 79.800 11.100 80.200 13.300 ;
        RECT 81.400 13.100 81.800 14.800 ;
        RECT 84.000 14.200 84.300 15.900 ;
        RECT 87.000 15.600 87.400 19.900 ;
        RECT 88.600 15.600 89.000 19.900 ;
        RECT 87.000 15.200 89.000 15.600 ;
        RECT 91.000 15.600 91.400 19.900 ;
        RECT 92.600 15.600 93.000 19.900 ;
        RECT 94.200 15.600 94.600 19.900 ;
        RECT 95.800 15.600 96.200 19.900 ;
        RECT 100.900 16.400 101.300 19.900 ;
        RECT 103.000 17.500 103.400 19.500 ;
        RECT 100.500 16.100 101.300 16.400 ;
        RECT 91.000 15.200 91.900 15.600 ;
        RECT 92.600 15.200 93.700 15.600 ;
        RECT 94.200 15.200 95.300 15.600 ;
        RECT 95.800 15.200 97.000 15.600 ;
        RECT 84.600 14.400 85.000 15.200 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 83.000 14.100 84.300 14.200 ;
        RECT 85.400 14.100 85.800 14.200 ;
        RECT 86.200 14.100 86.600 14.200 ;
        RECT 82.200 13.800 84.300 14.100 ;
        RECT 85.000 13.800 86.600 14.100 ;
        RECT 87.000 13.800 87.400 15.200 ;
        RECT 91.500 14.500 91.900 15.200 ;
        RECT 93.300 14.500 93.700 15.200 ;
        RECT 94.900 14.500 95.300 15.200 ;
        RECT 91.500 14.100 92.800 14.500 ;
        RECT 93.300 14.100 94.500 14.500 ;
        RECT 94.900 14.100 96.200 14.500 ;
        RECT 91.500 13.800 91.900 14.100 ;
        RECT 93.300 13.800 93.700 14.100 ;
        RECT 94.900 13.800 95.300 14.100 ;
        RECT 96.600 13.800 97.000 15.200 ;
        RECT 99.800 14.800 100.200 15.600 ;
        RECT 100.500 14.200 100.800 16.100 ;
        RECT 103.100 15.800 103.400 17.500 ;
        RECT 105.700 16.400 106.100 19.900 ;
        RECT 107.800 17.500 108.200 19.500 ;
        RECT 101.500 15.500 103.400 15.800 ;
        RECT 105.300 16.100 106.100 16.400 ;
        RECT 101.500 14.500 101.800 15.500 ;
        RECT 99.800 13.800 100.800 14.200 ;
        RECT 101.100 14.100 101.800 14.500 ;
        RECT 102.200 14.400 102.600 15.200 ;
        RECT 103.000 14.400 103.400 15.200 ;
        RECT 103.800 15.100 104.200 15.200 ;
        RECT 104.600 15.100 105.000 15.600 ;
        RECT 103.800 14.800 105.000 15.100 ;
        RECT 105.300 14.200 105.600 16.100 ;
        RECT 107.900 15.800 108.200 17.500 ;
        RECT 106.300 15.500 108.200 15.800 ;
        RECT 106.300 14.500 106.600 15.500 ;
        RECT 83.100 13.100 83.400 13.800 ;
        RECT 85.000 13.600 85.400 13.800 ;
        RECT 87.000 13.400 89.000 13.800 ;
        RECT 83.900 13.100 85.700 13.300 ;
        RECT 81.400 12.800 82.300 13.100 ;
        RECT 81.900 11.100 82.300 12.800 ;
        RECT 83.000 11.100 83.400 13.100 ;
        RECT 83.800 13.000 85.800 13.100 ;
        RECT 83.800 11.100 84.200 13.000 ;
        RECT 85.400 11.100 85.800 13.000 ;
        RECT 87.000 11.100 87.400 13.400 ;
        RECT 88.600 11.100 89.000 13.400 ;
        RECT 91.000 13.400 91.900 13.800 ;
        RECT 92.600 13.400 93.700 13.800 ;
        RECT 94.200 13.400 95.300 13.800 ;
        RECT 95.800 13.400 97.000 13.800 ;
        RECT 100.500 13.500 100.800 13.800 ;
        RECT 101.300 13.900 101.800 14.100 ;
        RECT 101.300 13.600 103.400 13.900 ;
        RECT 104.600 13.800 105.600 14.200 ;
        RECT 105.900 14.100 106.600 14.500 ;
        RECT 107.000 14.400 107.400 15.200 ;
        RECT 107.800 14.400 108.200 15.200 ;
        RECT 109.400 15.100 109.800 19.900 ;
        RECT 111.400 16.800 111.800 17.200 ;
        RECT 110.200 15.800 110.600 16.600 ;
        RECT 111.400 16.200 111.700 16.800 ;
        RECT 112.100 16.200 112.500 19.900 ;
        RECT 111.000 15.900 111.700 16.200 ;
        RECT 112.000 15.900 112.500 16.200 ;
        RECT 111.000 15.800 111.400 15.900 ;
        RECT 111.000 15.100 111.300 15.800 ;
        RECT 112.000 15.200 112.300 15.900 ;
        RECT 114.200 15.600 114.600 19.900 ;
        RECT 116.300 17.900 116.900 19.900 ;
        RECT 118.600 17.900 119.000 19.900 ;
        RECT 120.800 18.200 121.200 19.900 ;
        RECT 120.800 17.900 121.800 18.200 ;
        RECT 116.600 17.500 117.000 17.900 ;
        RECT 118.700 17.600 119.000 17.900 ;
        RECT 118.300 17.300 120.100 17.600 ;
        RECT 121.400 17.500 121.800 17.900 ;
        RECT 118.300 17.200 118.700 17.300 ;
        RECT 119.700 17.200 120.100 17.300 ;
        RECT 115.800 17.000 116.500 17.200 ;
        RECT 115.800 16.800 116.900 17.000 ;
        RECT 116.200 16.600 116.900 16.800 ;
        RECT 116.600 16.100 116.900 16.600 ;
        RECT 117.700 16.500 118.800 16.800 ;
        RECT 117.700 16.400 118.100 16.500 ;
        RECT 116.600 15.800 117.800 16.100 ;
        RECT 114.200 15.300 116.300 15.600 ;
        RECT 109.400 14.800 111.300 15.100 ;
        RECT 111.800 14.800 112.300 15.200 ;
        RECT 91.000 11.100 91.400 13.400 ;
        RECT 92.600 11.100 93.000 13.400 ;
        RECT 94.200 11.100 94.600 13.400 ;
        RECT 95.800 11.100 96.200 13.400 ;
        RECT 100.500 13.300 100.900 13.500 ;
        RECT 100.500 13.200 101.300 13.300 ;
        RECT 100.500 13.000 101.800 13.200 ;
        RECT 100.900 12.800 101.800 13.000 ;
        RECT 100.900 11.500 101.300 12.800 ;
        RECT 103.100 12.500 103.400 13.600 ;
        RECT 105.300 13.500 105.600 13.800 ;
        RECT 106.100 13.900 106.600 14.100 ;
        RECT 106.100 13.600 108.200 13.900 ;
        RECT 105.300 13.300 105.700 13.500 ;
        RECT 105.300 13.000 106.100 13.300 ;
        RECT 103.000 11.500 103.400 12.500 ;
        RECT 105.700 11.500 106.100 13.000 ;
        RECT 107.900 12.500 108.200 13.600 ;
        RECT 108.600 13.400 109.000 14.200 ;
        RECT 109.400 13.100 109.800 14.800 ;
        RECT 112.000 14.200 112.300 14.800 ;
        RECT 112.600 14.400 113.000 15.200 ;
        RECT 111.000 13.800 112.300 14.200 ;
        RECT 113.400 14.100 113.800 14.200 ;
        RECT 113.000 13.800 113.800 14.100 ;
        RECT 111.100 13.100 111.400 13.800 ;
        RECT 113.000 13.600 113.400 13.800 ;
        RECT 114.200 13.600 114.600 15.300 ;
        RECT 115.900 15.200 116.300 15.300 ;
        RECT 115.100 14.900 115.500 15.000 ;
        RECT 115.100 14.600 117.000 14.900 ;
        RECT 116.600 14.500 117.000 14.600 ;
        RECT 117.500 14.200 117.800 15.800 ;
        RECT 118.500 15.900 118.800 16.500 ;
        RECT 119.100 16.500 119.500 16.600 ;
        RECT 121.400 16.500 121.800 16.600 ;
        RECT 119.100 16.200 121.800 16.500 ;
        RECT 118.500 15.700 120.900 15.900 ;
        RECT 123.000 15.700 123.400 19.900 ;
        RECT 118.500 15.600 123.400 15.700 ;
        RECT 120.500 15.500 123.400 15.600 ;
        RECT 123.800 17.500 124.200 19.500 ;
        RECT 125.900 19.200 126.300 19.900 ;
        RECT 125.900 18.800 126.600 19.200 ;
        RECT 123.800 15.800 124.100 17.500 ;
        RECT 125.900 16.400 126.300 18.800 ;
        RECT 125.900 16.100 126.700 16.400 ;
        RECT 123.800 15.500 125.700 15.800 ;
        RECT 120.600 15.400 123.400 15.500 ;
        RECT 119.800 15.100 120.200 15.200 ;
        RECT 119.800 14.800 122.300 15.100 ;
        RECT 121.900 14.700 122.300 14.800 ;
        RECT 123.800 14.400 124.200 15.200 ;
        RECT 124.600 14.400 125.000 15.200 ;
        RECT 125.400 14.500 125.700 15.500 ;
        RECT 121.100 14.200 121.500 14.300 ;
        RECT 117.500 13.900 123.000 14.200 ;
        RECT 125.400 14.100 126.100 14.500 ;
        RECT 126.400 14.200 126.700 16.100 ;
        RECT 128.600 15.600 129.000 19.900 ;
        RECT 130.700 17.900 131.300 19.900 ;
        RECT 133.000 17.900 133.400 19.900 ;
        RECT 135.200 18.200 135.600 19.900 ;
        RECT 135.200 17.900 136.200 18.200 ;
        RECT 131.000 17.500 131.400 17.900 ;
        RECT 133.100 17.600 133.400 17.900 ;
        RECT 132.700 17.300 134.500 17.600 ;
        RECT 135.800 17.500 136.200 17.900 ;
        RECT 132.700 17.200 133.100 17.300 ;
        RECT 134.100 17.200 134.500 17.300 ;
        RECT 130.600 16.600 131.300 17.000 ;
        RECT 131.000 16.100 131.300 16.600 ;
        RECT 132.100 16.500 133.200 16.800 ;
        RECT 132.100 16.400 132.500 16.500 ;
        RECT 131.000 15.800 132.200 16.100 ;
        RECT 127.000 15.100 127.400 15.600 ;
        RECT 128.600 15.300 130.700 15.600 ;
        RECT 127.800 15.100 128.200 15.200 ;
        RECT 127.000 14.800 128.200 15.100 ;
        RECT 125.400 13.900 125.900 14.100 ;
        RECT 117.700 13.800 118.100 13.900 ;
        RECT 114.200 13.300 116.100 13.600 ;
        RECT 111.900 13.100 113.700 13.300 ;
        RECT 109.400 12.800 110.300 13.100 ;
        RECT 107.800 11.500 108.200 12.500 ;
        RECT 109.900 11.100 110.300 12.800 ;
        RECT 111.000 11.100 111.400 13.100 ;
        RECT 111.800 13.000 113.800 13.100 ;
        RECT 111.800 11.100 112.200 13.000 ;
        RECT 113.400 11.100 113.800 13.000 ;
        RECT 114.200 11.100 114.600 13.300 ;
        RECT 115.700 13.200 116.100 13.300 ;
        RECT 120.600 12.800 120.900 13.900 ;
        RECT 122.200 13.800 123.000 13.900 ;
        RECT 123.800 13.600 125.900 13.900 ;
        RECT 126.400 13.800 127.400 14.200 ;
        RECT 119.700 12.700 120.100 12.800 ;
        RECT 116.600 12.100 117.000 12.500 ;
        RECT 118.700 12.400 120.100 12.700 ;
        RECT 120.600 12.400 121.000 12.800 ;
        RECT 118.700 12.100 119.000 12.400 ;
        RECT 121.400 12.100 121.800 12.500 ;
        RECT 116.300 11.800 117.000 12.100 ;
        RECT 116.300 11.100 116.900 11.800 ;
        RECT 118.600 11.100 119.000 12.100 ;
        RECT 120.800 11.800 121.800 12.100 ;
        RECT 120.800 11.100 121.200 11.800 ;
        RECT 123.000 11.100 123.400 13.500 ;
        RECT 123.800 12.500 124.100 13.600 ;
        RECT 126.400 13.500 126.700 13.800 ;
        RECT 126.300 13.300 126.700 13.500 ;
        RECT 125.900 13.000 126.700 13.300 ;
        RECT 128.600 13.600 129.000 15.300 ;
        RECT 130.300 15.200 130.700 15.300 ;
        RECT 129.500 14.900 129.900 15.000 ;
        RECT 129.500 14.600 131.400 14.900 ;
        RECT 131.000 14.500 131.400 14.600 ;
        RECT 131.900 14.200 132.200 15.800 ;
        RECT 132.900 15.900 133.200 16.500 ;
        RECT 133.500 16.500 133.900 16.600 ;
        RECT 135.800 16.500 136.200 16.600 ;
        RECT 133.500 16.200 136.200 16.500 ;
        RECT 132.900 15.700 135.300 15.900 ;
        RECT 137.400 15.700 137.800 19.900 ;
        RECT 132.900 15.600 137.800 15.700 ;
        RECT 134.900 15.500 137.800 15.600 ;
        RECT 135.000 15.400 137.800 15.500 ;
        RECT 134.200 15.100 134.600 15.200 ;
        RECT 139.000 15.100 139.400 19.900 ;
        RECT 141.000 16.800 141.400 17.200 ;
        RECT 139.800 15.800 140.200 16.600 ;
        RECT 141.000 16.200 141.300 16.800 ;
        RECT 141.700 16.200 142.100 19.900 ;
        RECT 140.600 15.900 141.300 16.200 ;
        RECT 141.600 15.900 142.100 16.200 ;
        RECT 140.600 15.800 141.000 15.900 ;
        RECT 140.600 15.100 140.900 15.800 ;
        RECT 134.200 14.800 136.700 15.100 ;
        RECT 136.300 14.700 136.700 14.800 ;
        RECT 139.000 14.800 140.900 15.100 ;
        RECT 135.500 14.200 135.900 14.300 ;
        RECT 131.900 13.900 137.400 14.200 ;
        RECT 132.100 13.800 133.000 13.900 ;
        RECT 128.600 13.300 130.500 13.600 ;
        RECT 123.800 11.500 124.200 12.500 ;
        RECT 125.900 11.500 126.300 13.000 ;
        RECT 128.600 11.100 129.000 13.300 ;
        RECT 130.100 13.200 130.500 13.300 ;
        RECT 135.000 12.800 135.300 13.900 ;
        RECT 136.600 13.800 137.400 13.900 ;
        RECT 134.100 12.700 134.500 12.800 ;
        RECT 131.000 12.100 131.400 12.500 ;
        RECT 133.100 12.400 134.500 12.700 ;
        RECT 135.000 12.400 135.400 12.800 ;
        RECT 133.100 12.100 133.400 12.400 ;
        RECT 135.800 12.100 136.200 12.500 ;
        RECT 130.700 11.800 131.400 12.100 ;
        RECT 130.700 11.100 131.300 11.800 ;
        RECT 133.000 11.100 133.400 12.100 ;
        RECT 135.200 11.800 136.200 12.100 ;
        RECT 135.200 11.100 135.600 11.800 ;
        RECT 137.400 11.100 137.800 13.500 ;
        RECT 138.200 13.400 138.600 14.200 ;
        RECT 139.000 13.100 139.400 14.800 ;
        RECT 141.600 14.200 141.900 15.900 ;
        RECT 143.800 15.800 144.200 16.600 ;
        RECT 142.200 14.400 142.600 15.200 ;
        RECT 139.800 14.100 140.200 14.200 ;
        RECT 140.600 14.100 141.900 14.200 ;
        RECT 143.000 14.100 143.400 14.200 ;
        RECT 139.800 13.800 141.900 14.100 ;
        RECT 142.600 13.800 143.400 14.100 ;
        RECT 140.700 13.100 141.000 13.800 ;
        RECT 142.600 13.600 143.000 13.800 ;
        RECT 141.500 13.100 143.300 13.300 ;
        RECT 144.600 13.100 145.000 19.900 ;
        RECT 146.200 15.800 146.600 16.600 ;
        RECT 145.400 13.400 145.800 14.200 ;
        RECT 147.000 13.100 147.400 19.900 ;
        RECT 152.100 16.400 152.500 19.900 ;
        RECT 154.200 17.500 154.600 19.500 ;
        RECT 151.700 16.100 152.500 16.400 ;
        RECT 151.000 14.800 151.400 15.600 ;
        RECT 151.700 14.200 152.000 16.100 ;
        RECT 154.300 15.800 154.600 17.500 ;
        RECT 152.700 15.500 154.600 15.800 ;
        RECT 152.700 14.500 153.000 15.500 ;
        RECT 147.800 13.400 148.200 14.200 ;
        RECT 149.400 14.100 149.800 14.200 ;
        RECT 151.000 14.100 152.000 14.200 ;
        RECT 152.300 14.100 153.000 14.500 ;
        RECT 153.400 14.400 153.800 15.200 ;
        RECT 154.200 14.400 154.600 15.200 ;
        RECT 155.800 15.100 156.200 19.900 ;
        RECT 158.500 18.200 158.900 19.900 ;
        RECT 158.500 17.800 159.400 18.200 ;
        RECT 157.800 16.800 158.200 17.200 ;
        RECT 156.600 15.800 157.000 16.600 ;
        RECT 157.800 16.200 158.100 16.800 ;
        RECT 158.500 16.200 158.900 17.800 ;
        RECT 157.400 15.900 158.100 16.200 ;
        RECT 158.400 15.900 158.900 16.200 ;
        RECT 157.400 15.800 157.800 15.900 ;
        RECT 157.400 15.100 157.700 15.800 ;
        RECT 155.800 14.800 157.700 15.100 ;
        RECT 149.400 13.800 152.000 14.100 ;
        RECT 151.700 13.500 152.000 13.800 ;
        RECT 152.500 13.900 153.000 14.100 ;
        RECT 152.500 13.600 154.600 13.900 ;
        RECT 139.000 12.800 139.900 13.100 ;
        RECT 139.500 11.100 139.900 12.800 ;
        RECT 140.600 11.100 141.000 13.100 ;
        RECT 141.400 13.000 143.400 13.100 ;
        RECT 141.400 11.100 141.800 13.000 ;
        RECT 143.000 11.100 143.400 13.000 ;
        RECT 144.100 12.800 145.000 13.100 ;
        RECT 146.500 12.800 147.400 13.100 ;
        RECT 151.700 13.300 152.100 13.500 ;
        RECT 151.700 13.000 152.500 13.300 ;
        RECT 144.100 12.200 144.500 12.800 ;
        RECT 146.500 12.200 146.900 12.800 ;
        RECT 143.800 11.800 144.500 12.200 ;
        RECT 146.200 11.800 146.900 12.200 ;
        RECT 144.100 11.100 144.500 11.800 ;
        RECT 146.500 11.100 146.900 11.800 ;
        RECT 152.100 11.500 152.500 13.000 ;
        RECT 154.300 12.500 154.600 13.600 ;
        RECT 155.000 13.400 155.400 14.200 ;
        RECT 155.800 13.100 156.200 14.800 ;
        RECT 158.400 14.200 158.700 15.900 ;
        RECT 160.600 15.700 161.000 19.900 ;
        RECT 162.800 18.200 163.200 19.900 ;
        RECT 162.200 17.900 163.200 18.200 ;
        RECT 165.000 17.900 165.400 19.900 ;
        RECT 167.100 17.900 167.700 19.900 ;
        RECT 162.200 17.500 162.600 17.900 ;
        RECT 165.000 17.600 165.300 17.900 ;
        RECT 163.900 17.300 165.700 17.600 ;
        RECT 167.000 17.500 167.400 17.900 ;
        RECT 163.900 17.200 164.300 17.300 ;
        RECT 165.300 17.200 165.700 17.300 ;
        RECT 162.200 16.500 162.600 16.600 ;
        RECT 164.500 16.500 164.900 16.600 ;
        RECT 162.200 16.200 164.900 16.500 ;
        RECT 165.200 16.500 166.300 16.800 ;
        RECT 165.200 15.900 165.500 16.500 ;
        RECT 165.900 16.400 166.300 16.500 ;
        RECT 167.100 16.600 167.800 17.000 ;
        RECT 167.100 16.100 167.400 16.600 ;
        RECT 163.100 15.700 165.500 15.900 ;
        RECT 160.600 15.600 165.500 15.700 ;
        RECT 166.200 15.800 167.400 16.100 ;
        RECT 160.600 15.500 163.500 15.600 ;
        RECT 160.600 15.400 163.400 15.500 ;
        RECT 159.000 14.400 159.400 15.200 ;
        RECT 163.800 15.100 164.200 15.200 ;
        RECT 161.700 14.800 164.200 15.100 ;
        RECT 161.700 14.700 162.100 14.800 ;
        RECT 163.000 14.700 163.400 14.800 ;
        RECT 162.500 14.200 162.900 14.300 ;
        RECT 166.200 14.200 166.500 15.800 ;
        RECT 169.400 15.600 169.800 19.900 ;
        RECT 170.200 15.800 170.600 16.600 ;
        RECT 171.000 16.100 171.400 19.900 ;
        RECT 173.000 16.800 173.400 17.200 ;
        RECT 173.000 16.200 173.300 16.800 ;
        RECT 173.700 16.200 174.100 19.900 ;
        RECT 172.600 16.100 173.300 16.200 ;
        RECT 171.000 15.900 173.300 16.100 ;
        RECT 173.600 15.900 174.100 16.200 ;
        RECT 171.000 15.800 173.000 15.900 ;
        RECT 167.700 15.300 169.800 15.600 ;
        RECT 167.700 15.200 168.100 15.300 ;
        RECT 168.500 14.900 168.900 15.000 ;
        RECT 167.000 14.600 168.900 14.900 ;
        RECT 167.000 14.500 167.400 14.600 ;
        RECT 157.400 13.800 158.700 14.200 ;
        RECT 159.800 14.100 160.200 14.200 ;
        RECT 159.400 13.800 160.200 14.100 ;
        RECT 161.000 13.900 166.500 14.200 ;
        RECT 161.000 13.800 161.800 13.900 ;
        RECT 157.500 13.100 157.800 13.800 ;
        RECT 159.400 13.600 159.800 13.800 ;
        RECT 158.300 13.100 160.100 13.300 ;
        RECT 155.800 12.800 156.700 13.100 ;
        RECT 154.200 11.500 154.600 12.500 ;
        RECT 156.300 11.100 156.700 12.800 ;
        RECT 157.400 11.100 157.800 13.100 ;
        RECT 158.200 13.000 160.200 13.100 ;
        RECT 158.200 11.100 158.600 13.000 ;
        RECT 159.800 11.100 160.200 13.000 ;
        RECT 160.600 11.100 161.000 13.500 ;
        RECT 163.100 12.800 163.400 13.900 ;
        RECT 165.900 13.800 166.300 13.900 ;
        RECT 169.400 13.600 169.800 15.300 ;
        RECT 167.900 13.300 169.800 13.600 ;
        RECT 167.900 13.200 168.300 13.300 ;
        RECT 162.200 12.100 162.600 12.500 ;
        RECT 163.000 12.400 163.400 12.800 ;
        RECT 163.900 12.700 164.300 12.800 ;
        RECT 163.900 12.400 165.300 12.700 ;
        RECT 165.000 12.100 165.300 12.400 ;
        RECT 167.000 12.100 167.400 12.500 ;
        RECT 162.200 11.800 163.200 12.100 ;
        RECT 162.800 11.100 163.200 11.800 ;
        RECT 165.000 11.100 165.400 12.100 ;
        RECT 167.000 11.800 167.700 12.100 ;
        RECT 167.100 11.100 167.700 11.800 ;
        RECT 169.400 11.100 169.800 13.300 ;
        RECT 171.000 13.100 171.400 15.800 ;
        RECT 173.600 15.200 173.900 15.900 ;
        RECT 175.800 15.600 176.200 19.900 ;
        RECT 177.900 17.900 178.500 19.900 ;
        RECT 180.200 17.900 180.600 19.900 ;
        RECT 182.400 18.200 182.800 19.900 ;
        RECT 182.400 17.900 183.400 18.200 ;
        RECT 178.200 17.500 178.600 17.900 ;
        RECT 180.300 17.600 180.600 17.900 ;
        RECT 179.900 17.300 181.700 17.600 ;
        RECT 183.000 17.500 183.400 17.900 ;
        RECT 179.900 17.200 180.300 17.300 ;
        RECT 181.300 17.200 181.700 17.300 ;
        RECT 177.800 16.600 178.500 17.000 ;
        RECT 178.200 16.100 178.500 16.600 ;
        RECT 179.300 16.500 180.400 16.800 ;
        RECT 179.300 16.400 179.700 16.500 ;
        RECT 178.200 15.800 179.400 16.100 ;
        RECT 175.800 15.300 177.900 15.600 ;
        RECT 173.400 14.800 173.900 15.200 ;
        RECT 173.600 14.200 173.900 14.800 ;
        RECT 174.200 14.400 174.600 15.200 ;
        RECT 171.800 13.400 172.200 14.200 ;
        RECT 172.600 13.800 173.900 14.200 ;
        RECT 175.000 14.100 175.400 14.200 ;
        RECT 174.600 13.800 175.400 14.100 ;
        RECT 172.700 13.100 173.000 13.800 ;
        RECT 174.600 13.600 175.000 13.800 ;
        RECT 175.800 13.600 176.200 15.300 ;
        RECT 177.500 15.200 177.900 15.300 ;
        RECT 176.700 14.900 177.100 15.000 ;
        RECT 176.700 14.600 178.600 14.900 ;
        RECT 178.200 14.500 178.600 14.600 ;
        RECT 179.100 14.200 179.400 15.800 ;
        RECT 180.100 15.900 180.400 16.500 ;
        RECT 180.700 16.500 181.100 16.600 ;
        RECT 183.000 16.500 183.400 16.600 ;
        RECT 180.700 16.200 183.400 16.500 ;
        RECT 180.100 15.700 182.500 15.900 ;
        RECT 184.600 15.700 185.000 19.900 ;
        RECT 186.700 16.200 187.100 19.900 ;
        RECT 187.400 16.800 187.800 17.200 ;
        RECT 187.500 16.200 187.800 16.800 ;
        RECT 186.700 15.900 187.200 16.200 ;
        RECT 187.500 15.900 188.200 16.200 ;
        RECT 180.100 15.600 185.000 15.700 ;
        RECT 182.100 15.500 185.000 15.600 ;
        RECT 182.200 15.400 185.000 15.500 ;
        RECT 180.600 15.100 181.000 15.200 ;
        RECT 181.400 15.100 181.800 15.200 ;
        RECT 180.600 14.800 183.900 15.100 ;
        RECT 183.500 14.700 183.900 14.800 ;
        RECT 186.200 14.400 186.600 15.200 ;
        RECT 182.700 14.200 183.100 14.300 ;
        RECT 186.900 14.200 187.200 15.900 ;
        RECT 187.800 15.800 188.200 15.900 ;
        RECT 188.600 15.800 189.000 16.600 ;
        RECT 187.800 15.100 188.100 15.800 ;
        RECT 189.400 15.100 189.800 19.900 ;
        RECT 191.000 15.700 191.400 19.900 ;
        RECT 193.200 18.200 193.600 19.900 ;
        RECT 192.600 17.900 193.600 18.200 ;
        RECT 195.400 17.900 195.800 19.900 ;
        RECT 197.500 17.900 198.100 19.900 ;
        RECT 192.600 17.500 193.000 17.900 ;
        RECT 195.400 17.600 195.700 17.900 ;
        RECT 194.300 17.300 196.100 17.600 ;
        RECT 197.400 17.500 197.800 17.900 ;
        RECT 194.300 17.200 194.700 17.300 ;
        RECT 195.700 17.200 196.100 17.300 ;
        RECT 192.600 16.500 193.000 16.600 ;
        RECT 194.900 16.500 195.300 16.600 ;
        RECT 192.600 16.200 195.300 16.500 ;
        RECT 195.600 16.500 196.700 16.800 ;
        RECT 195.600 15.900 195.900 16.500 ;
        RECT 196.300 16.400 196.700 16.500 ;
        RECT 197.500 16.600 198.200 17.000 ;
        RECT 197.500 16.100 197.800 16.600 ;
        RECT 193.500 15.700 195.900 15.900 ;
        RECT 191.000 15.600 195.900 15.700 ;
        RECT 196.600 15.800 197.800 16.100 ;
        RECT 191.000 15.500 193.900 15.600 ;
        RECT 191.000 15.400 193.800 15.500 ;
        RECT 194.200 15.100 194.600 15.200 ;
        RECT 187.800 14.800 189.800 15.100 ;
        RECT 179.100 13.900 184.600 14.200 ;
        RECT 179.300 13.800 179.700 13.900 ;
        RECT 175.800 13.300 177.700 13.600 ;
        RECT 173.500 13.100 175.300 13.300 ;
        RECT 170.500 12.800 171.400 13.100 ;
        RECT 170.500 11.100 170.900 12.800 ;
        RECT 172.600 11.100 173.000 13.100 ;
        RECT 173.400 13.000 175.400 13.100 ;
        RECT 173.400 11.100 173.800 13.000 ;
        RECT 175.000 11.100 175.400 13.000 ;
        RECT 175.800 11.100 176.200 13.300 ;
        RECT 177.300 13.200 177.700 13.300 ;
        RECT 182.200 12.800 182.500 13.900 ;
        RECT 183.800 13.800 184.600 13.900 ;
        RECT 185.400 14.100 185.800 14.200 ;
        RECT 185.400 13.800 186.200 14.100 ;
        RECT 186.900 13.800 188.200 14.200 ;
        RECT 185.800 13.600 186.200 13.800 ;
        RECT 181.300 12.700 181.700 12.800 ;
        RECT 178.200 12.100 178.600 12.500 ;
        RECT 180.300 12.400 181.700 12.700 ;
        RECT 182.200 12.400 182.600 12.800 ;
        RECT 180.300 12.100 180.600 12.400 ;
        RECT 183.000 12.100 183.400 12.500 ;
        RECT 177.900 11.800 178.600 12.100 ;
        RECT 177.900 11.100 178.500 11.800 ;
        RECT 180.200 11.100 180.600 12.100 ;
        RECT 182.400 11.800 183.400 12.100 ;
        RECT 182.400 11.100 182.800 11.800 ;
        RECT 184.600 11.100 185.000 13.500 ;
        RECT 185.500 13.100 187.300 13.300 ;
        RECT 187.800 13.200 188.100 13.800 ;
        RECT 185.400 13.000 187.400 13.100 ;
        RECT 185.400 11.100 185.800 13.000 ;
        RECT 187.000 11.100 187.400 13.000 ;
        RECT 187.800 11.100 188.200 13.200 ;
        RECT 189.400 13.100 189.800 14.800 ;
        RECT 192.100 14.800 194.600 15.100 ;
        RECT 192.100 14.700 192.500 14.800 ;
        RECT 192.900 14.200 193.300 14.300 ;
        RECT 196.600 14.200 196.900 15.800 ;
        RECT 199.800 15.600 200.200 19.900 ;
        RECT 204.100 16.400 204.500 19.900 ;
        RECT 206.200 17.500 206.600 19.500 ;
        RECT 203.700 16.100 204.500 16.400 ;
        RECT 198.100 15.300 200.200 15.600 ;
        RECT 198.100 15.200 198.500 15.300 ;
        RECT 199.800 15.100 200.200 15.300 ;
        RECT 203.000 15.100 203.400 15.600 ;
        RECT 198.900 14.900 199.300 15.000 ;
        RECT 197.400 14.600 199.300 14.900 ;
        RECT 199.800 14.800 203.400 15.100 ;
        RECT 197.400 14.500 197.800 14.600 ;
        RECT 190.200 13.400 190.600 14.200 ;
        RECT 191.400 13.900 196.900 14.200 ;
        RECT 191.400 13.800 192.200 13.900 ;
        RECT 188.900 12.800 189.800 13.100 ;
        RECT 188.900 11.100 189.300 12.800 ;
        RECT 191.000 11.100 191.400 13.500 ;
        RECT 193.500 12.800 193.800 13.900 ;
        RECT 196.300 13.800 196.700 13.900 ;
        RECT 199.800 13.600 200.200 14.800 ;
        RECT 203.700 14.200 204.000 16.100 ;
        RECT 206.300 15.800 206.600 17.500 ;
        RECT 207.800 16.400 208.200 19.900 ;
        RECT 204.700 15.500 206.600 15.800 ;
        RECT 207.700 15.900 208.200 16.400 ;
        RECT 209.400 16.200 209.800 19.900 ;
        RECT 208.500 15.900 209.800 16.200 ;
        RECT 210.200 17.500 210.600 19.500 ;
        RECT 212.300 19.200 212.700 19.900 ;
        RECT 211.800 18.800 212.700 19.200 ;
        RECT 204.700 14.500 205.000 15.500 ;
        RECT 201.400 14.100 201.800 14.200 ;
        RECT 203.000 14.100 204.000 14.200 ;
        RECT 204.300 14.100 205.000 14.500 ;
        RECT 205.400 14.400 205.800 15.200 ;
        RECT 206.200 14.400 206.600 15.200 ;
        RECT 207.700 14.200 208.000 15.900 ;
        RECT 208.500 14.900 208.800 15.900 ;
        RECT 210.200 15.800 210.500 17.500 ;
        RECT 212.300 16.400 212.700 18.800 ;
        RECT 212.300 16.100 213.100 16.400 ;
        RECT 210.200 15.500 212.100 15.800 ;
        RECT 208.300 14.500 208.800 14.900 ;
        RECT 201.400 13.800 204.000 14.100 ;
        RECT 198.300 13.300 200.200 13.600 ;
        RECT 198.300 13.200 198.700 13.300 ;
        RECT 192.600 12.100 193.000 12.500 ;
        RECT 193.400 12.400 193.800 12.800 ;
        RECT 194.300 12.700 194.700 12.800 ;
        RECT 194.300 12.400 195.700 12.700 ;
        RECT 195.400 12.100 195.700 12.400 ;
        RECT 197.400 12.100 197.800 12.500 ;
        RECT 192.600 11.800 193.600 12.100 ;
        RECT 193.200 11.100 193.600 11.800 ;
        RECT 195.400 11.100 195.800 12.100 ;
        RECT 197.400 11.800 198.100 12.100 ;
        RECT 197.500 11.100 198.100 11.800 ;
        RECT 199.800 11.100 200.200 13.300 ;
        RECT 203.700 13.500 204.000 13.800 ;
        RECT 204.500 13.900 205.000 14.100 ;
        RECT 207.000 14.100 207.400 14.200 ;
        RECT 207.700 14.100 208.200 14.200 ;
        RECT 204.500 13.600 206.600 13.900 ;
        RECT 207.000 13.800 208.200 14.100 ;
        RECT 203.700 13.300 204.100 13.500 ;
        RECT 203.700 13.000 204.500 13.300 ;
        RECT 204.100 11.500 204.500 13.000 ;
        RECT 206.300 12.500 206.600 13.600 ;
        RECT 207.700 13.100 208.000 13.800 ;
        RECT 208.500 13.700 208.800 14.500 ;
        RECT 209.300 14.800 209.800 15.200 ;
        RECT 209.300 14.400 209.700 14.800 ;
        RECT 210.200 14.400 210.600 15.200 ;
        RECT 211.000 14.400 211.400 15.200 ;
        RECT 211.800 14.500 212.100 15.500 ;
        RECT 211.800 14.100 212.500 14.500 ;
        RECT 212.800 14.200 213.100 16.100 ;
        RECT 216.300 16.200 216.700 19.900 ;
        RECT 217.000 16.800 217.400 17.200 ;
        RECT 217.100 16.200 217.400 16.800 ;
        RECT 216.300 15.900 216.800 16.200 ;
        RECT 217.100 15.900 217.800 16.200 ;
        RECT 213.400 14.800 213.800 15.600 ;
        RECT 215.800 14.400 216.200 15.200 ;
        RECT 216.500 14.200 216.800 15.900 ;
        RECT 217.400 15.800 217.800 15.900 ;
        RECT 218.200 15.800 218.600 16.600 ;
        RECT 217.400 15.100 217.700 15.800 ;
        RECT 219.000 15.100 219.400 19.900 ;
        RECT 221.900 16.200 222.300 19.900 ;
        RECT 222.600 16.800 223.000 17.200 ;
        RECT 222.700 16.200 223.000 16.800 ;
        RECT 221.900 15.900 222.400 16.200 ;
        RECT 222.700 15.900 223.400 16.200 ;
        RECT 217.400 14.800 219.400 15.100 ;
        RECT 211.800 13.900 212.300 14.100 ;
        RECT 208.500 13.400 209.800 13.700 ;
        RECT 207.700 12.800 208.200 13.100 ;
        RECT 206.200 11.500 206.600 12.500 ;
        RECT 207.800 11.100 208.200 12.800 ;
        RECT 209.400 11.100 209.800 13.400 ;
        RECT 210.200 13.600 212.300 13.900 ;
        RECT 212.800 13.800 213.800 14.200 ;
        RECT 215.000 14.100 215.400 14.200 ;
        RECT 215.000 13.800 215.800 14.100 ;
        RECT 216.500 13.800 217.800 14.200 ;
        RECT 210.200 12.500 210.500 13.600 ;
        RECT 212.800 13.500 213.100 13.800 ;
        RECT 215.400 13.600 215.800 13.800 ;
        RECT 212.700 13.300 213.100 13.500 ;
        RECT 212.300 13.000 213.100 13.300 ;
        RECT 215.100 13.100 216.900 13.300 ;
        RECT 217.400 13.100 217.700 13.800 ;
        RECT 219.000 13.100 219.400 14.800 ;
        RECT 221.400 14.400 221.800 15.200 ;
        RECT 222.100 14.200 222.400 15.900 ;
        RECT 223.000 15.800 223.400 15.900 ;
        RECT 223.800 15.800 224.200 16.600 ;
        RECT 223.000 15.100 223.300 15.800 ;
        RECT 224.600 15.100 225.000 19.900 ;
        RECT 225.400 17.100 225.800 17.200 ;
        RECT 226.200 17.100 226.600 19.900 ;
        RECT 228.300 17.900 228.900 19.900 ;
        RECT 230.600 17.900 231.000 19.900 ;
        RECT 232.800 18.200 233.200 19.900 ;
        RECT 232.800 17.900 233.800 18.200 ;
        RECT 228.600 17.500 229.000 17.900 ;
        RECT 230.700 17.600 231.000 17.900 ;
        RECT 230.300 17.300 232.100 17.600 ;
        RECT 233.400 17.500 233.800 17.900 ;
        RECT 230.300 17.200 230.700 17.300 ;
        RECT 231.700 17.200 232.100 17.300 ;
        RECT 225.400 16.800 226.600 17.100 ;
        RECT 223.000 14.800 225.000 15.100 ;
        RECT 219.800 13.400 220.200 14.200 ;
        RECT 220.600 14.100 221.000 14.200 ;
        RECT 222.100 14.100 223.400 14.200 ;
        RECT 223.800 14.100 224.200 14.200 ;
        RECT 220.600 13.800 221.400 14.100 ;
        RECT 222.100 13.800 224.200 14.100 ;
        RECT 221.000 13.600 221.400 13.800 ;
        RECT 220.700 13.100 222.500 13.300 ;
        RECT 223.000 13.100 223.300 13.800 ;
        RECT 224.600 13.100 225.000 14.800 ;
        RECT 226.200 15.600 226.600 16.800 ;
        RECT 228.200 16.600 228.900 17.000 ;
        RECT 228.600 16.100 228.900 16.600 ;
        RECT 229.700 16.500 230.800 16.800 ;
        RECT 229.700 16.400 230.100 16.500 ;
        RECT 228.600 15.800 229.800 16.100 ;
        RECT 226.200 15.300 228.300 15.600 ;
        RECT 225.400 13.400 225.800 14.200 ;
        RECT 226.200 13.600 226.600 15.300 ;
        RECT 227.900 15.200 228.300 15.300 ;
        RECT 227.100 14.900 227.500 15.000 ;
        RECT 227.100 14.600 229.000 14.900 ;
        RECT 228.600 14.500 229.000 14.600 ;
        RECT 229.500 14.200 229.800 15.800 ;
        RECT 230.500 15.900 230.800 16.500 ;
        RECT 231.100 16.500 231.500 16.600 ;
        RECT 233.400 16.500 233.800 16.600 ;
        RECT 231.100 16.200 233.800 16.500 ;
        RECT 230.500 15.700 232.900 15.900 ;
        RECT 235.000 15.700 235.400 19.900 ;
        RECT 230.500 15.600 235.400 15.700 ;
        RECT 236.600 15.600 237.000 19.900 ;
        RECT 238.200 15.600 238.600 19.900 ;
        RECT 239.800 15.600 240.200 19.900 ;
        RECT 241.400 15.600 241.800 19.900 ;
        RECT 243.800 15.600 244.200 19.900 ;
        RECT 245.400 15.600 245.800 19.900 ;
        RECT 247.000 15.600 247.400 19.900 ;
        RECT 248.600 15.600 249.000 19.900 ;
        RECT 250.200 15.800 250.600 16.600 ;
        RECT 232.500 15.500 235.400 15.600 ;
        RECT 232.600 15.400 235.400 15.500 ;
        RECT 235.800 15.200 237.000 15.600 ;
        RECT 237.500 15.200 238.600 15.600 ;
        RECT 239.100 15.200 240.200 15.600 ;
        RECT 240.900 15.200 241.800 15.600 ;
        RECT 243.000 15.200 244.200 15.600 ;
        RECT 244.700 15.200 245.800 15.600 ;
        RECT 246.300 15.200 247.400 15.600 ;
        RECT 248.100 15.200 249.000 15.600 ;
        RECT 231.800 15.100 232.200 15.200 ;
        RECT 231.800 14.800 234.300 15.100 ;
        RECT 233.900 14.700 234.300 14.800 ;
        RECT 233.100 14.200 233.500 14.300 ;
        RECT 229.500 13.900 235.000 14.200 ;
        RECT 229.700 13.800 230.100 13.900 ;
        RECT 215.000 13.000 217.000 13.100 ;
        RECT 210.200 11.500 210.600 12.500 ;
        RECT 212.300 11.500 212.700 13.000 ;
        RECT 215.000 11.100 215.400 13.000 ;
        RECT 216.600 11.100 217.000 13.000 ;
        RECT 217.400 11.100 217.800 13.100 ;
        RECT 218.500 12.800 219.400 13.100 ;
        RECT 220.600 13.000 222.600 13.100 ;
        RECT 218.500 11.100 218.900 12.800 ;
        RECT 220.600 11.100 221.000 13.000 ;
        RECT 222.200 11.100 222.600 13.000 ;
        RECT 223.000 11.100 223.400 13.100 ;
        RECT 224.100 12.800 225.000 13.100 ;
        RECT 226.200 13.300 228.100 13.600 ;
        RECT 224.100 11.100 224.500 12.800 ;
        RECT 226.200 11.100 226.600 13.300 ;
        RECT 227.700 13.200 228.100 13.300 ;
        RECT 232.600 12.800 232.900 13.900 ;
        RECT 234.200 13.800 235.000 13.900 ;
        RECT 235.800 13.800 236.200 15.200 ;
        RECT 237.500 14.500 237.900 15.200 ;
        RECT 239.100 14.500 239.500 15.200 ;
        RECT 240.900 14.500 241.300 15.200 ;
        RECT 236.600 14.100 237.900 14.500 ;
        RECT 238.300 14.100 239.500 14.500 ;
        RECT 240.000 14.100 241.300 14.500 ;
        RECT 241.700 14.100 242.600 14.500 ;
        RECT 237.500 13.800 237.900 14.100 ;
        RECT 239.100 13.800 239.500 14.100 ;
        RECT 240.900 13.800 241.300 14.100 ;
        RECT 242.200 13.800 242.600 14.100 ;
        RECT 243.000 13.800 243.400 15.200 ;
        RECT 244.700 14.500 245.100 15.200 ;
        RECT 246.300 14.500 246.700 15.200 ;
        RECT 248.100 14.500 248.500 15.200 ;
        RECT 243.800 14.100 245.100 14.500 ;
        RECT 245.500 14.100 246.700 14.500 ;
        RECT 247.200 14.100 248.500 14.500 ;
        RECT 244.700 13.800 245.100 14.100 ;
        RECT 246.300 13.800 246.700 14.100 ;
        RECT 248.100 13.800 248.500 14.100 ;
        RECT 231.700 12.700 232.100 12.800 ;
        RECT 228.600 12.100 229.000 12.500 ;
        RECT 230.700 12.400 232.100 12.700 ;
        RECT 232.600 12.400 233.000 12.800 ;
        RECT 230.700 12.100 231.000 12.400 ;
        RECT 233.400 12.100 233.800 12.500 ;
        RECT 228.300 11.800 229.000 12.100 ;
        RECT 228.300 11.100 228.900 11.800 ;
        RECT 230.600 11.100 231.000 12.100 ;
        RECT 232.800 11.800 233.800 12.100 ;
        RECT 232.800 11.100 233.200 11.800 ;
        RECT 235.000 11.100 235.400 13.500 ;
        RECT 235.800 13.400 237.000 13.800 ;
        RECT 237.500 13.400 238.600 13.800 ;
        RECT 239.100 13.400 240.200 13.800 ;
        RECT 240.900 13.400 241.800 13.800 ;
        RECT 243.000 13.400 244.200 13.800 ;
        RECT 244.700 13.400 245.800 13.800 ;
        RECT 246.300 13.400 247.400 13.800 ;
        RECT 248.100 13.400 249.000 13.800 ;
        RECT 236.600 11.100 237.000 13.400 ;
        RECT 238.200 11.100 238.600 13.400 ;
        RECT 239.800 11.100 240.200 13.400 ;
        RECT 241.400 11.100 241.800 13.400 ;
        RECT 243.800 11.100 244.200 13.400 ;
        RECT 245.400 11.100 245.800 13.400 ;
        RECT 247.000 11.100 247.400 13.400 ;
        RECT 248.600 11.100 249.000 13.400 ;
        RECT 251.000 13.100 251.400 19.900 ;
        RECT 251.800 13.400 252.200 14.200 ;
        RECT 250.500 12.800 251.400 13.100 ;
        RECT 250.500 11.100 250.900 12.800 ;
        RECT 1.400 7.600 1.800 9.900 ;
        RECT 3.000 7.600 3.400 9.900 ;
        RECT 4.600 7.600 5.000 9.900 ;
        RECT 6.200 7.600 6.600 9.900 ;
        RECT 8.600 7.600 9.000 9.900 ;
        RECT 10.200 7.600 10.600 9.900 ;
        RECT 11.800 7.600 12.200 9.900 ;
        RECT 13.400 7.600 13.800 9.900 ;
        RECT 15.000 8.000 15.400 9.900 ;
        RECT 16.600 8.000 17.000 9.900 ;
        RECT 15.000 7.900 17.000 8.000 ;
        RECT 17.400 7.900 17.800 9.900 ;
        RECT 15.100 7.700 16.900 7.900 ;
        RECT 1.400 7.200 2.300 7.600 ;
        RECT 3.000 7.200 4.100 7.600 ;
        RECT 4.600 7.200 5.700 7.600 ;
        RECT 6.200 7.200 7.400 7.600 ;
        RECT 8.600 7.200 9.500 7.600 ;
        RECT 10.200 7.200 11.300 7.600 ;
        RECT 11.800 7.200 12.900 7.600 ;
        RECT 13.400 7.200 14.600 7.600 ;
        RECT 15.400 7.200 15.800 7.400 ;
        RECT 17.400 7.200 17.700 7.900 ;
        RECT 18.200 7.500 18.600 9.900 ;
        RECT 20.400 9.200 20.800 9.900 ;
        RECT 19.800 8.900 20.800 9.200 ;
        RECT 22.600 8.900 23.000 9.900 ;
        RECT 24.700 9.200 25.300 9.900 ;
        RECT 24.600 8.900 25.300 9.200 ;
        RECT 19.800 8.500 20.200 8.900 ;
        RECT 22.600 8.600 22.900 8.900 ;
        RECT 20.600 8.200 21.000 8.600 ;
        RECT 21.500 8.300 22.900 8.600 ;
        RECT 24.600 8.500 25.000 8.900 ;
        RECT 21.500 8.200 21.900 8.300 ;
        RECT 1.900 6.900 2.300 7.200 ;
        RECT 3.700 6.900 4.100 7.200 ;
        RECT 5.300 6.900 5.700 7.200 ;
        RECT 1.900 6.500 3.200 6.900 ;
        RECT 3.700 6.500 4.900 6.900 ;
        RECT 5.300 6.500 6.600 6.900 ;
        RECT 1.900 5.800 2.300 6.500 ;
        RECT 3.700 5.800 4.100 6.500 ;
        RECT 5.300 5.800 5.700 6.500 ;
        RECT 7.000 5.800 7.400 7.200 ;
        RECT 7.800 6.900 8.200 7.200 ;
        RECT 9.100 6.900 9.500 7.200 ;
        RECT 10.900 6.900 11.300 7.200 ;
        RECT 12.500 6.900 12.900 7.200 ;
        RECT 7.800 6.500 8.700 6.900 ;
        RECT 9.100 6.500 10.400 6.900 ;
        RECT 10.900 6.500 12.100 6.900 ;
        RECT 12.500 6.500 13.800 6.900 ;
        RECT 9.100 5.800 9.500 6.500 ;
        RECT 10.900 5.800 11.300 6.500 ;
        RECT 12.500 5.800 12.900 6.500 ;
        RECT 14.200 6.100 14.600 7.200 ;
        RECT 15.000 6.900 15.800 7.200 ;
        RECT 15.000 6.800 15.400 6.900 ;
        RECT 16.500 6.800 17.800 7.200 ;
        RECT 18.600 7.100 19.400 7.200 ;
        RECT 20.700 7.100 21.000 8.200 ;
        RECT 25.500 7.700 25.900 7.800 ;
        RECT 27.000 7.700 27.400 9.900 ;
        RECT 25.500 7.400 27.400 7.700 ;
        RECT 23.500 7.100 23.900 7.200 ;
        RECT 18.600 6.800 24.100 7.100 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 14.200 5.800 15.400 6.100 ;
        RECT 15.800 5.800 16.200 6.600 ;
        RECT 16.500 6.200 16.800 6.800 ;
        RECT 20.100 6.700 20.500 6.800 ;
        RECT 19.300 6.200 19.700 6.300 ;
        RECT 20.600 6.200 21.000 6.300 ;
        RECT 16.500 5.800 17.000 6.200 ;
        RECT 19.300 5.900 21.800 6.200 ;
        RECT 21.400 5.800 21.800 5.900 ;
        RECT 1.400 5.400 2.300 5.800 ;
        RECT 3.000 5.400 4.100 5.800 ;
        RECT 4.600 5.400 5.700 5.800 ;
        RECT 6.200 5.400 7.400 5.800 ;
        RECT 8.600 5.400 9.500 5.800 ;
        RECT 10.200 5.400 11.300 5.800 ;
        RECT 11.800 5.400 12.900 5.800 ;
        RECT 13.400 5.400 14.600 5.800 ;
        RECT 1.400 1.100 1.800 5.400 ;
        RECT 3.000 1.100 3.400 5.400 ;
        RECT 4.600 1.100 5.000 5.400 ;
        RECT 6.200 1.100 6.600 5.400 ;
        RECT 8.600 1.100 9.000 5.400 ;
        RECT 10.200 1.100 10.600 5.400 ;
        RECT 11.800 1.100 12.200 5.400 ;
        RECT 13.400 1.100 13.800 5.400 ;
        RECT 16.500 5.100 16.800 5.800 ;
        RECT 18.200 5.500 21.000 5.600 ;
        RECT 18.200 5.400 21.100 5.500 ;
        RECT 18.200 5.300 23.100 5.400 ;
        RECT 17.400 5.100 17.800 5.200 ;
        RECT 16.300 4.800 16.800 5.100 ;
        RECT 17.100 4.800 17.800 5.100 ;
        RECT 16.300 1.100 16.700 4.800 ;
        RECT 17.100 4.200 17.400 4.800 ;
        RECT 17.000 3.800 17.400 4.200 ;
        RECT 18.200 1.100 18.600 5.300 ;
        RECT 20.700 5.100 23.100 5.300 ;
        RECT 19.800 4.500 22.500 4.800 ;
        RECT 19.800 4.400 20.200 4.500 ;
        RECT 22.100 4.400 22.500 4.500 ;
        RECT 22.800 4.500 23.100 5.100 ;
        RECT 23.800 5.200 24.100 6.800 ;
        RECT 24.600 6.400 25.000 6.500 ;
        RECT 24.600 6.100 26.500 6.400 ;
        RECT 26.100 6.000 26.500 6.100 ;
        RECT 25.300 5.700 25.700 5.800 ;
        RECT 27.000 5.700 27.400 7.400 ;
        RECT 28.600 8.900 29.000 9.900 ;
        RECT 28.600 7.200 28.900 8.900 ;
        RECT 29.400 7.800 29.800 8.600 ;
        RECT 30.300 8.200 30.700 8.600 ;
        RECT 30.200 7.800 30.600 8.200 ;
        RECT 31.000 7.900 31.400 9.900 ;
        RECT 28.600 7.100 29.000 7.200 ;
        RECT 30.200 7.100 30.500 7.800 ;
        RECT 28.600 6.800 30.500 7.100 ;
        RECT 25.300 5.400 27.400 5.700 ;
        RECT 27.800 5.400 28.200 6.200 ;
        RECT 23.800 4.900 25.000 5.200 ;
        RECT 23.500 4.500 23.900 4.600 ;
        RECT 22.800 4.200 23.900 4.500 ;
        RECT 24.700 4.400 25.000 4.900 ;
        RECT 24.700 4.000 25.400 4.400 ;
        RECT 21.500 3.700 21.900 3.800 ;
        RECT 22.900 3.700 23.300 3.800 ;
        RECT 19.800 3.100 20.200 3.500 ;
        RECT 21.500 3.400 23.300 3.700 ;
        RECT 22.600 3.100 22.900 3.400 ;
        RECT 24.600 3.100 25.000 3.500 ;
        RECT 19.800 2.800 20.800 3.100 ;
        RECT 20.400 1.100 20.800 2.800 ;
        RECT 22.600 1.100 23.000 3.100 ;
        RECT 24.700 1.100 25.300 3.100 ;
        RECT 27.000 1.100 27.400 5.400 ;
        RECT 28.600 5.100 28.900 6.800 ;
        RECT 31.100 6.200 31.400 7.900 ;
        RECT 33.400 7.500 33.800 9.900 ;
        RECT 35.600 9.200 36.000 9.900 ;
        RECT 35.000 8.900 36.000 9.200 ;
        RECT 37.800 8.900 38.200 9.900 ;
        RECT 39.900 9.200 40.500 9.900 ;
        RECT 39.800 8.900 40.500 9.200 ;
        RECT 35.000 8.500 35.400 8.900 ;
        RECT 37.800 8.600 38.100 8.900 ;
        RECT 35.800 8.200 36.200 8.600 ;
        RECT 36.700 8.300 38.100 8.600 ;
        RECT 39.800 8.500 40.200 8.900 ;
        RECT 36.700 8.200 37.100 8.300 ;
        RECT 31.800 6.400 32.200 7.200 ;
        RECT 33.800 7.100 34.600 7.200 ;
        RECT 35.900 7.100 36.200 8.200 ;
        RECT 40.700 7.700 41.100 7.800 ;
        RECT 42.200 7.700 42.600 9.900 ;
        RECT 43.000 8.000 43.400 9.900 ;
        RECT 44.600 8.000 45.000 9.900 ;
        RECT 43.000 7.900 45.000 8.000 ;
        RECT 45.400 7.900 45.800 9.900 ;
        RECT 46.500 8.200 46.900 9.900 ;
        RECT 49.400 9.100 49.800 9.200 ;
        RECT 50.200 9.100 50.600 9.900 ;
        RECT 49.400 8.800 50.600 9.100 ;
        RECT 52.300 9.200 52.900 9.900 ;
        RECT 52.300 8.900 53.000 9.200 ;
        RECT 54.600 8.900 55.000 9.900 ;
        RECT 56.800 9.200 57.200 9.900 ;
        RECT 56.800 8.900 57.800 9.200 ;
        RECT 46.500 7.900 47.400 8.200 ;
        RECT 43.100 7.700 44.900 7.900 ;
        RECT 40.700 7.400 42.600 7.700 ;
        RECT 38.700 7.100 39.100 7.200 ;
        RECT 33.800 6.800 39.300 7.100 ;
        RECT 35.300 6.700 35.700 6.800 ;
        RECT 34.500 6.200 34.900 6.300 ;
        RECT 35.800 6.200 36.200 6.300 ;
        RECT 30.200 6.100 30.600 6.200 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 32.600 6.100 33.000 6.200 ;
        RECT 30.200 5.800 31.400 6.100 ;
        RECT 32.200 5.800 33.000 6.100 ;
        RECT 34.500 5.900 37.000 6.200 ;
        RECT 36.600 5.800 37.000 5.900 ;
        RECT 30.300 5.100 30.600 5.800 ;
        RECT 32.200 5.600 32.600 5.800 ;
        RECT 33.400 5.500 36.200 5.600 ;
        RECT 33.400 5.400 36.300 5.500 ;
        RECT 33.400 5.300 38.300 5.400 ;
        RECT 28.100 4.700 29.000 5.100 ;
        RECT 28.100 1.100 28.500 4.700 ;
        RECT 30.200 1.100 30.600 5.100 ;
        RECT 31.000 4.800 33.000 5.100 ;
        RECT 31.000 1.100 31.400 4.800 ;
        RECT 32.600 1.100 33.000 4.800 ;
        RECT 33.400 1.100 33.800 5.300 ;
        RECT 35.900 5.100 38.300 5.300 ;
        RECT 35.000 4.500 37.700 4.800 ;
        RECT 35.000 4.400 35.400 4.500 ;
        RECT 37.300 4.400 37.700 4.500 ;
        RECT 38.000 4.500 38.300 5.100 ;
        RECT 39.000 5.200 39.300 6.800 ;
        RECT 39.800 6.400 40.200 6.500 ;
        RECT 39.800 6.100 41.700 6.400 ;
        RECT 41.300 6.000 41.700 6.100 ;
        RECT 40.500 5.700 40.900 5.800 ;
        RECT 42.200 5.700 42.600 7.400 ;
        RECT 43.400 7.200 43.800 7.400 ;
        RECT 45.400 7.200 45.700 7.900 ;
        RECT 43.000 6.900 43.800 7.200 ;
        RECT 44.500 7.100 45.800 7.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 43.000 6.800 43.400 6.900 ;
        RECT 44.500 6.800 46.600 7.100 ;
        RECT 43.800 5.800 44.200 6.600 ;
        RECT 40.500 5.400 42.600 5.700 ;
        RECT 39.000 4.900 40.200 5.200 ;
        RECT 38.700 4.500 39.100 4.600 ;
        RECT 38.000 4.200 39.100 4.500 ;
        RECT 39.900 4.400 40.200 4.900 ;
        RECT 39.900 4.000 40.600 4.400 ;
        RECT 36.700 3.700 37.100 3.800 ;
        RECT 38.100 3.700 38.500 3.800 ;
        RECT 35.000 3.100 35.400 3.500 ;
        RECT 36.700 3.400 38.500 3.700 ;
        RECT 37.800 3.100 38.100 3.400 ;
        RECT 39.800 3.100 40.200 3.500 ;
        RECT 35.000 2.800 36.000 3.100 ;
        RECT 35.600 1.100 36.000 2.800 ;
        RECT 37.800 1.100 38.200 3.100 ;
        RECT 39.900 1.100 40.500 3.100 ;
        RECT 42.200 1.100 42.600 5.400 ;
        RECT 44.500 5.100 44.800 6.800 ;
        RECT 47.000 6.100 47.400 7.900 ;
        RECT 50.200 7.700 50.600 8.800 ;
        RECT 52.600 8.500 53.000 8.900 ;
        RECT 54.700 8.600 55.000 8.900 ;
        RECT 54.700 8.300 56.100 8.600 ;
        RECT 55.700 8.200 56.100 8.300 ;
        RECT 56.600 8.200 57.000 8.600 ;
        RECT 57.400 8.500 57.800 8.900 ;
        RECT 51.700 7.700 52.100 7.800 ;
        RECT 47.800 7.100 48.200 7.600 ;
        RECT 50.200 7.400 52.100 7.700 ;
        RECT 49.400 7.100 49.800 7.200 ;
        RECT 47.800 6.800 49.800 7.100 ;
        RECT 45.400 5.800 47.400 6.100 ;
        RECT 45.400 5.200 45.700 5.800 ;
        RECT 45.400 5.100 45.800 5.200 ;
        RECT 44.300 4.800 44.800 5.100 ;
        RECT 45.100 4.800 45.800 5.100 ;
        RECT 44.300 1.100 44.700 4.800 ;
        RECT 45.100 4.200 45.400 4.800 ;
        RECT 46.200 4.400 46.600 5.200 ;
        RECT 45.000 3.800 45.400 4.200 ;
        RECT 47.000 1.100 47.400 5.800 ;
        RECT 50.200 5.700 50.600 7.400 ;
        RECT 53.400 7.100 54.100 7.200 ;
        RECT 56.600 7.100 56.900 8.200 ;
        RECT 59.000 7.500 59.400 9.900 ;
        RECT 59.800 7.700 60.200 9.900 ;
        RECT 61.900 9.200 62.500 9.900 ;
        RECT 61.900 8.900 62.600 9.200 ;
        RECT 64.200 8.900 64.600 9.900 ;
        RECT 66.400 9.200 66.800 9.900 ;
        RECT 66.400 8.900 67.400 9.200 ;
        RECT 62.200 8.500 62.600 8.900 ;
        RECT 64.300 8.600 64.600 8.900 ;
        RECT 64.300 8.300 65.700 8.600 ;
        RECT 65.300 8.200 65.700 8.300 ;
        RECT 66.200 7.800 66.600 8.600 ;
        RECT 67.000 8.500 67.400 8.900 ;
        RECT 61.300 7.700 61.700 7.800 ;
        RECT 59.800 7.400 61.700 7.700 ;
        RECT 58.200 7.100 59.000 7.200 ;
        RECT 53.400 6.800 59.000 7.100 ;
        RECT 52.600 6.400 53.000 6.500 ;
        RECT 51.100 6.100 53.000 6.400 ;
        RECT 51.100 6.000 51.500 6.100 ;
        RECT 51.900 5.700 52.300 5.800 ;
        RECT 50.200 5.400 52.300 5.700 ;
        RECT 50.200 1.100 50.600 5.400 ;
        RECT 53.500 5.200 53.800 6.800 ;
        RECT 57.100 6.700 57.500 6.800 ;
        RECT 57.900 6.200 58.300 6.300 ;
        RECT 55.800 5.900 58.300 6.200 ;
        RECT 55.800 5.800 56.200 5.900 ;
        RECT 59.800 5.700 60.200 7.400 ;
        RECT 63.300 7.100 63.700 7.200 ;
        RECT 66.200 7.100 66.500 7.800 ;
        RECT 68.600 7.500 69.000 9.900 ;
        RECT 69.400 7.600 69.800 9.900 ;
        RECT 71.000 8.200 71.400 9.900 ;
        RECT 71.000 7.900 71.500 8.200 ;
        RECT 69.400 7.300 70.700 7.600 ;
        RECT 67.800 7.100 68.600 7.200 ;
        RECT 63.100 6.800 68.600 7.100 ;
        RECT 62.200 6.400 62.600 6.500 ;
        RECT 60.700 6.100 62.600 6.400 ;
        RECT 60.700 6.000 61.100 6.100 ;
        RECT 61.500 5.700 61.900 5.800 ;
        RECT 56.600 5.500 59.400 5.600 ;
        RECT 56.500 5.400 59.400 5.500 ;
        RECT 52.600 4.900 53.800 5.200 ;
        RECT 54.500 5.300 59.400 5.400 ;
        RECT 54.500 5.100 56.900 5.300 ;
        RECT 52.600 4.400 52.900 4.900 ;
        RECT 52.200 4.000 52.900 4.400 ;
        RECT 53.700 4.500 54.100 4.600 ;
        RECT 54.500 4.500 54.800 5.100 ;
        RECT 53.700 4.200 54.800 4.500 ;
        RECT 55.100 4.500 57.800 4.800 ;
        RECT 55.100 4.400 55.500 4.500 ;
        RECT 57.400 4.400 57.800 4.500 ;
        RECT 54.300 3.700 54.700 3.800 ;
        RECT 55.700 3.700 56.100 3.800 ;
        RECT 52.600 3.100 53.000 3.500 ;
        RECT 54.300 3.400 56.100 3.700 ;
        RECT 54.700 3.100 55.000 3.400 ;
        RECT 57.400 3.100 57.800 3.500 ;
        RECT 52.300 1.100 52.900 3.100 ;
        RECT 54.600 1.100 55.000 3.100 ;
        RECT 56.800 2.800 57.800 3.100 ;
        RECT 56.800 1.100 57.200 2.800 ;
        RECT 59.000 1.100 59.400 5.300 ;
        RECT 59.800 5.400 61.900 5.700 ;
        RECT 59.800 1.100 60.200 5.400 ;
        RECT 63.100 5.200 63.400 6.800 ;
        RECT 66.700 6.700 67.100 6.800 ;
        RECT 67.500 6.200 67.900 6.300 ;
        RECT 69.500 6.200 69.900 6.600 ;
        RECT 63.800 6.100 64.200 6.200 ;
        RECT 65.400 6.100 67.900 6.200 ;
        RECT 63.800 5.900 67.900 6.100 ;
        RECT 63.800 5.800 65.800 5.900 ;
        RECT 69.400 5.800 69.900 6.200 ;
        RECT 70.400 6.500 70.700 7.300 ;
        RECT 71.200 7.200 71.500 7.900 ;
        RECT 72.600 7.500 73.000 9.900 ;
        RECT 74.800 9.200 75.200 9.900 ;
        RECT 74.200 8.900 75.200 9.200 ;
        RECT 77.000 8.900 77.400 9.900 ;
        RECT 79.100 9.200 79.700 9.900 ;
        RECT 79.000 8.900 79.700 9.200 ;
        RECT 74.200 8.500 74.600 8.900 ;
        RECT 77.000 8.600 77.300 8.900 ;
        RECT 75.000 8.200 75.400 8.600 ;
        RECT 75.900 8.300 77.300 8.600 ;
        RECT 79.000 8.500 79.400 8.900 ;
        RECT 75.900 8.200 76.300 8.300 ;
        RECT 71.000 6.800 71.500 7.200 ;
        RECT 73.000 7.100 73.800 7.200 ;
        RECT 75.100 7.100 75.400 8.200 ;
        RECT 78.200 8.100 78.600 8.200 ;
        RECT 78.200 7.800 80.200 8.100 ;
        RECT 79.800 7.700 80.300 7.800 ;
        RECT 81.400 7.700 81.800 9.900 ;
        RECT 83.500 8.200 83.900 9.900 ;
        RECT 79.800 7.400 81.800 7.700 ;
        RECT 83.000 7.900 83.900 8.200 ;
        RECT 84.600 7.900 85.000 9.900 ;
        RECT 85.400 8.000 85.800 9.900 ;
        RECT 87.000 8.000 87.400 9.900 ;
        RECT 85.400 7.900 87.400 8.000 ;
        RECT 77.900 7.100 78.300 7.200 ;
        RECT 81.400 7.100 81.800 7.400 ;
        RECT 82.200 7.100 82.600 7.600 ;
        RECT 73.000 6.800 78.500 7.100 ;
        RECT 70.400 6.100 70.900 6.500 ;
        RECT 66.200 5.500 69.000 5.600 ;
        RECT 66.100 5.400 69.000 5.500 ;
        RECT 62.200 4.900 63.400 5.200 ;
        RECT 64.100 5.300 69.000 5.400 ;
        RECT 64.100 5.100 66.500 5.300 ;
        RECT 62.200 4.400 62.500 4.900 ;
        RECT 61.800 4.000 62.500 4.400 ;
        RECT 63.300 4.500 63.700 4.600 ;
        RECT 64.100 4.500 64.400 5.100 ;
        RECT 63.300 4.200 64.400 4.500 ;
        RECT 64.700 4.500 67.400 4.800 ;
        RECT 64.700 4.400 65.100 4.500 ;
        RECT 67.000 4.400 67.400 4.500 ;
        RECT 63.900 3.700 64.300 3.800 ;
        RECT 65.300 3.700 65.700 3.800 ;
        RECT 62.200 3.100 62.600 3.500 ;
        RECT 63.900 3.400 65.700 3.700 ;
        RECT 64.300 3.100 64.600 3.400 ;
        RECT 67.000 3.100 67.400 3.500 ;
        RECT 61.900 1.100 62.500 3.100 ;
        RECT 64.200 1.100 64.600 3.100 ;
        RECT 66.400 2.800 67.400 3.100 ;
        RECT 66.400 1.100 66.800 2.800 ;
        RECT 68.600 1.100 69.000 5.300 ;
        RECT 70.400 5.100 70.700 6.100 ;
        RECT 71.200 5.100 71.500 6.800 ;
        RECT 74.500 6.700 74.900 6.800 ;
        RECT 73.700 6.200 74.100 6.300 ;
        RECT 73.700 5.900 76.200 6.200 ;
        RECT 75.800 5.800 76.200 5.900 ;
        RECT 69.400 4.800 70.700 5.100 ;
        RECT 69.400 1.100 69.800 4.800 ;
        RECT 71.000 4.600 71.500 5.100 ;
        RECT 72.600 5.500 75.400 5.600 ;
        RECT 72.600 5.400 75.500 5.500 ;
        RECT 72.600 5.300 77.500 5.400 ;
        RECT 71.000 1.100 71.400 4.600 ;
        RECT 72.600 1.100 73.000 5.300 ;
        RECT 75.100 5.100 77.500 5.300 ;
        RECT 74.200 4.500 76.900 4.800 ;
        RECT 74.200 4.400 74.600 4.500 ;
        RECT 76.500 4.400 76.900 4.500 ;
        RECT 77.200 4.500 77.500 5.100 ;
        RECT 78.200 5.200 78.500 6.800 ;
        RECT 81.400 6.800 82.600 7.100 ;
        RECT 79.000 6.400 79.400 6.500 ;
        RECT 79.000 6.100 80.900 6.400 ;
        RECT 80.500 6.000 80.900 6.100 ;
        RECT 79.700 5.700 80.100 5.800 ;
        RECT 81.400 5.700 81.800 6.800 ;
        RECT 79.700 5.400 81.800 5.700 ;
        RECT 78.200 4.900 79.400 5.200 ;
        RECT 77.900 4.500 78.300 4.600 ;
        RECT 77.200 4.200 78.300 4.500 ;
        RECT 79.100 4.400 79.400 4.900 ;
        RECT 79.100 4.000 79.800 4.400 ;
        RECT 75.900 3.700 76.300 3.800 ;
        RECT 77.300 3.700 77.700 3.800 ;
        RECT 74.200 3.100 74.600 3.500 ;
        RECT 75.900 3.400 77.700 3.700 ;
        RECT 77.000 3.100 77.300 3.400 ;
        RECT 79.000 3.100 79.400 3.500 ;
        RECT 74.200 2.800 75.200 3.100 ;
        RECT 74.800 1.100 75.200 2.800 ;
        RECT 77.000 1.100 77.400 3.100 ;
        RECT 79.100 1.100 79.700 3.100 ;
        RECT 81.400 1.100 81.800 5.400 ;
        RECT 83.000 6.100 83.400 7.900 ;
        RECT 84.700 7.200 85.000 7.900 ;
        RECT 85.500 7.700 87.300 7.900 ;
        RECT 87.800 7.600 88.200 9.900 ;
        RECT 89.400 8.200 89.800 9.900 ;
        RECT 89.400 7.900 89.900 8.200 ;
        RECT 86.600 7.200 87.000 7.400 ;
        RECT 87.800 7.300 89.100 7.600 ;
        RECT 83.800 7.100 84.200 7.200 ;
        RECT 84.600 7.100 85.900 7.200 ;
        RECT 83.800 6.800 85.900 7.100 ;
        RECT 86.600 6.900 87.400 7.200 ;
        RECT 87.000 6.800 87.400 6.900 ;
        RECT 83.000 5.800 84.900 6.100 ;
        RECT 83.000 1.100 83.400 5.800 ;
        RECT 84.600 5.200 84.900 5.800 ;
        RECT 83.800 4.400 84.200 5.200 ;
        RECT 84.600 5.100 85.000 5.200 ;
        RECT 85.600 5.100 85.900 6.800 ;
        RECT 86.200 5.800 86.600 6.600 ;
        RECT 87.900 6.200 88.300 6.600 ;
        RECT 87.800 5.800 88.300 6.200 ;
        RECT 88.800 6.500 89.100 7.300 ;
        RECT 89.600 7.200 89.900 7.900 ;
        RECT 89.400 6.800 89.900 7.200 ;
        RECT 88.800 6.100 89.300 6.500 ;
        RECT 88.800 5.100 89.100 6.100 ;
        RECT 89.600 5.100 89.900 6.800 ;
        RECT 84.600 4.800 85.300 5.100 ;
        RECT 85.600 4.800 86.100 5.100 ;
        RECT 85.000 4.200 85.300 4.800 ;
        RECT 85.000 3.800 85.400 4.200 ;
        RECT 85.700 1.100 86.100 4.800 ;
        RECT 87.800 4.800 89.100 5.100 ;
        RECT 87.800 1.100 88.200 4.800 ;
        RECT 89.400 4.600 89.900 5.100 ;
        RECT 91.000 7.700 91.400 9.900 ;
        RECT 93.100 9.200 93.700 9.900 ;
        RECT 93.100 8.900 93.800 9.200 ;
        RECT 95.400 8.900 95.800 9.900 ;
        RECT 97.600 9.200 98.000 9.900 ;
        RECT 97.600 8.900 98.600 9.200 ;
        RECT 93.400 8.500 93.800 8.900 ;
        RECT 95.500 8.600 95.800 8.900 ;
        RECT 95.500 8.300 96.900 8.600 ;
        RECT 96.500 8.200 96.900 8.300 ;
        RECT 97.400 8.200 97.800 8.600 ;
        RECT 98.200 8.500 98.600 8.900 ;
        RECT 92.500 7.700 92.900 7.800 ;
        RECT 91.000 7.400 92.900 7.700 ;
        RECT 91.000 5.700 91.400 7.400 ;
        RECT 94.500 7.100 94.900 7.200 ;
        RECT 95.800 7.100 96.200 7.200 ;
        RECT 97.400 7.100 97.700 8.200 ;
        RECT 99.800 7.500 100.200 9.900 ;
        RECT 103.500 8.200 103.900 9.900 ;
        RECT 103.000 7.900 103.900 8.200 ;
        RECT 104.600 7.900 105.000 9.900 ;
        RECT 105.400 8.000 105.800 9.900 ;
        RECT 107.000 8.000 107.400 9.900 ;
        RECT 105.400 7.900 107.400 8.000 ;
        RECT 99.000 7.100 99.800 7.200 ;
        RECT 94.300 6.800 99.800 7.100 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 102.200 7.100 102.600 7.600 ;
        RECT 100.600 6.800 102.600 7.100 ;
        RECT 93.400 6.400 93.800 6.500 ;
        RECT 91.900 6.100 93.800 6.400 ;
        RECT 91.900 6.000 92.300 6.100 ;
        RECT 92.700 5.700 93.100 5.800 ;
        RECT 91.000 5.400 93.100 5.700 ;
        RECT 89.400 1.100 89.800 4.600 ;
        RECT 91.000 1.100 91.400 5.400 ;
        RECT 94.300 5.200 94.600 6.800 ;
        RECT 97.900 6.700 98.300 6.800 ;
        RECT 97.400 6.200 97.800 6.300 ;
        RECT 98.700 6.200 99.100 6.300 ;
        RECT 96.600 5.900 99.100 6.200 ;
        RECT 103.000 6.100 103.400 7.900 ;
        RECT 104.700 7.200 105.000 7.900 ;
        RECT 105.500 7.700 107.300 7.900 ;
        RECT 108.600 7.600 109.000 9.900 ;
        RECT 110.200 7.600 110.600 9.900 ;
        RECT 111.800 7.600 112.200 9.900 ;
        RECT 113.400 7.600 113.800 9.900 ;
        RECT 106.600 7.200 107.000 7.400 ;
        RECT 108.600 7.200 109.500 7.600 ;
        RECT 110.200 7.200 111.300 7.600 ;
        RECT 111.800 7.200 112.900 7.600 ;
        RECT 113.400 7.200 114.600 7.600 ;
        RECT 115.000 7.500 115.400 9.900 ;
        RECT 117.200 9.200 117.600 9.900 ;
        RECT 116.600 8.900 117.600 9.200 ;
        RECT 119.400 8.900 119.800 9.900 ;
        RECT 121.500 9.200 122.100 9.900 ;
        RECT 121.400 8.900 122.100 9.200 ;
        RECT 116.600 8.500 117.000 8.900 ;
        RECT 119.400 8.600 119.700 8.900 ;
        RECT 117.400 8.200 117.800 8.600 ;
        RECT 118.300 8.300 119.700 8.600 ;
        RECT 121.400 8.500 121.800 8.900 ;
        RECT 118.300 8.200 118.700 8.300 ;
        RECT 103.800 7.100 104.200 7.200 ;
        RECT 104.600 7.100 105.900 7.200 ;
        RECT 103.800 6.800 105.900 7.100 ;
        RECT 106.600 6.900 107.400 7.200 ;
        RECT 107.000 6.800 107.400 6.900 ;
        RECT 107.800 6.900 108.200 7.200 ;
        RECT 109.100 6.900 109.500 7.200 ;
        RECT 110.900 6.900 111.300 7.200 ;
        RECT 112.500 6.900 112.900 7.200 ;
        RECT 96.600 5.800 97.000 5.900 ;
        RECT 103.000 5.800 104.900 6.100 ;
        RECT 97.400 5.500 100.200 5.600 ;
        RECT 97.300 5.400 100.200 5.500 ;
        RECT 93.400 4.900 94.600 5.200 ;
        RECT 95.300 5.300 100.200 5.400 ;
        RECT 95.300 5.100 97.700 5.300 ;
        RECT 93.400 4.400 93.700 4.900 ;
        RECT 93.000 4.000 93.700 4.400 ;
        RECT 94.500 4.500 94.900 4.600 ;
        RECT 95.300 4.500 95.600 5.100 ;
        RECT 94.500 4.200 95.600 4.500 ;
        RECT 95.900 4.500 98.600 4.800 ;
        RECT 95.900 4.400 96.300 4.500 ;
        RECT 98.200 4.400 98.600 4.500 ;
        RECT 95.100 3.700 95.500 3.800 ;
        RECT 96.500 3.700 96.900 3.800 ;
        RECT 93.400 3.100 93.800 3.500 ;
        RECT 95.100 3.400 96.900 3.700 ;
        RECT 95.500 3.100 95.800 3.400 ;
        RECT 98.200 3.100 98.600 3.500 ;
        RECT 93.100 1.100 93.700 3.100 ;
        RECT 95.400 1.100 95.800 3.100 ;
        RECT 97.600 2.800 98.600 3.100 ;
        RECT 97.600 1.100 98.000 2.800 ;
        RECT 99.800 1.100 100.200 5.300 ;
        RECT 103.000 1.100 103.400 5.800 ;
        RECT 104.600 5.200 104.900 5.800 ;
        RECT 103.800 4.400 104.200 5.200 ;
        RECT 104.600 5.100 105.000 5.200 ;
        RECT 105.600 5.100 105.900 6.800 ;
        RECT 106.200 5.800 106.600 6.600 ;
        RECT 107.800 6.500 108.700 6.900 ;
        RECT 109.100 6.500 110.400 6.900 ;
        RECT 110.900 6.500 112.100 6.900 ;
        RECT 112.500 6.500 113.800 6.900 ;
        RECT 109.100 5.800 109.500 6.500 ;
        RECT 110.900 5.800 111.300 6.500 ;
        RECT 112.500 5.800 112.900 6.500 ;
        RECT 114.200 5.800 114.600 7.200 ;
        RECT 115.400 7.100 116.200 7.200 ;
        RECT 117.500 7.100 117.800 8.200 ;
        RECT 120.600 8.100 121.000 8.200 ;
        RECT 120.600 7.800 122.600 8.100 ;
        RECT 122.200 7.700 122.700 7.800 ;
        RECT 123.800 7.700 124.200 9.900 ;
        RECT 125.900 8.200 126.300 9.900 ;
        RECT 122.200 7.400 124.200 7.700 ;
        RECT 125.400 7.900 126.300 8.200 ;
        RECT 127.000 7.900 127.400 9.900 ;
        RECT 127.800 8.000 128.200 9.900 ;
        RECT 129.400 8.000 129.800 9.900 ;
        RECT 127.800 7.900 129.800 8.000 ;
        RECT 119.800 7.100 120.700 7.200 ;
        RECT 123.800 7.100 124.200 7.400 ;
        RECT 124.600 7.100 125.000 7.600 ;
        RECT 115.400 6.800 120.900 7.100 ;
        RECT 116.900 6.700 117.300 6.800 ;
        RECT 116.100 6.200 116.500 6.300 ;
        RECT 116.100 5.900 118.600 6.200 ;
        RECT 118.200 5.800 118.600 5.900 ;
        RECT 108.600 5.400 109.500 5.800 ;
        RECT 110.200 5.400 111.300 5.800 ;
        RECT 111.800 5.400 112.900 5.800 ;
        RECT 113.400 5.400 114.600 5.800 ;
        RECT 115.000 5.500 117.800 5.600 ;
        RECT 115.000 5.400 117.900 5.500 ;
        RECT 104.600 4.800 105.300 5.100 ;
        RECT 105.600 4.800 106.100 5.100 ;
        RECT 105.000 4.200 105.300 4.800 ;
        RECT 105.000 3.800 105.400 4.200 ;
        RECT 105.700 1.100 106.100 4.800 ;
        RECT 108.600 1.100 109.000 5.400 ;
        RECT 110.200 1.100 110.600 5.400 ;
        RECT 111.800 1.100 112.200 5.400 ;
        RECT 113.400 1.100 113.800 5.400 ;
        RECT 115.000 5.300 119.900 5.400 ;
        RECT 115.000 1.100 115.400 5.300 ;
        RECT 117.500 5.100 119.900 5.300 ;
        RECT 116.600 4.500 119.300 4.800 ;
        RECT 116.600 4.400 117.000 4.500 ;
        RECT 118.900 4.400 119.300 4.500 ;
        RECT 119.600 4.500 119.900 5.100 ;
        RECT 120.600 5.200 120.900 6.800 ;
        RECT 123.800 6.800 125.000 7.100 ;
        RECT 121.400 6.400 121.800 6.500 ;
        RECT 121.400 6.100 123.300 6.400 ;
        RECT 122.900 6.000 123.300 6.100 ;
        RECT 122.100 5.700 122.500 5.800 ;
        RECT 123.800 5.700 124.200 6.800 ;
        RECT 122.100 5.400 124.200 5.700 ;
        RECT 120.600 4.900 121.800 5.200 ;
        RECT 120.300 4.500 120.700 4.600 ;
        RECT 119.600 4.200 120.700 4.500 ;
        RECT 121.500 4.400 121.800 4.900 ;
        RECT 121.500 4.000 122.200 4.400 ;
        RECT 118.300 3.700 118.700 3.800 ;
        RECT 119.700 3.700 120.100 3.800 ;
        RECT 116.600 3.100 117.000 3.500 ;
        RECT 118.300 3.400 120.100 3.700 ;
        RECT 119.400 3.100 119.700 3.400 ;
        RECT 121.400 3.100 121.800 3.500 ;
        RECT 116.600 2.800 117.600 3.100 ;
        RECT 117.200 1.100 117.600 2.800 ;
        RECT 119.400 1.100 119.800 3.100 ;
        RECT 121.500 1.100 122.100 3.100 ;
        RECT 123.800 1.100 124.200 5.400 ;
        RECT 125.400 6.100 125.800 7.900 ;
        RECT 127.100 7.200 127.400 7.900 ;
        RECT 127.900 7.700 129.700 7.900 ;
        RECT 130.200 7.500 130.600 9.900 ;
        RECT 132.400 9.200 132.800 9.900 ;
        RECT 131.800 8.900 132.800 9.200 ;
        RECT 134.600 8.900 135.000 9.900 ;
        RECT 136.700 9.200 137.300 9.900 ;
        RECT 136.600 8.900 137.300 9.200 ;
        RECT 131.800 8.500 132.200 8.900 ;
        RECT 134.600 8.600 134.900 8.900 ;
        RECT 132.600 7.800 133.000 8.600 ;
        RECT 133.500 8.300 134.900 8.600 ;
        RECT 136.600 8.500 137.000 8.900 ;
        RECT 133.500 8.200 133.900 8.300 ;
        RECT 129.000 7.200 129.400 7.400 ;
        RECT 126.200 7.100 126.600 7.200 ;
        RECT 127.000 7.100 128.300 7.200 ;
        RECT 126.200 6.800 128.300 7.100 ;
        RECT 129.000 6.900 129.800 7.200 ;
        RECT 129.400 6.800 129.800 6.900 ;
        RECT 130.600 7.100 131.400 7.200 ;
        RECT 132.700 7.100 133.000 7.800 ;
        RECT 137.500 7.700 137.900 7.800 ;
        RECT 139.000 7.700 139.400 9.900 ;
        RECT 139.800 7.900 140.200 9.900 ;
        RECT 140.600 8.000 141.000 9.900 ;
        RECT 142.200 8.000 142.600 9.900 ;
        RECT 140.600 7.900 142.600 8.000 ;
        RECT 143.000 8.000 143.400 9.900 ;
        RECT 144.600 8.000 145.000 9.900 ;
        RECT 143.000 7.900 145.000 8.000 ;
        RECT 145.400 7.900 145.800 9.900 ;
        RECT 137.500 7.400 139.400 7.700 ;
        RECT 135.500 7.100 135.900 7.200 ;
        RECT 130.600 6.800 136.100 7.100 ;
        RECT 125.400 5.800 127.300 6.100 ;
        RECT 125.400 1.100 125.800 5.800 ;
        RECT 127.000 5.200 127.300 5.800 ;
        RECT 126.200 4.400 126.600 5.200 ;
        RECT 127.000 5.100 127.400 5.200 ;
        RECT 128.000 5.100 128.300 6.800 ;
        RECT 132.100 6.700 132.500 6.800 ;
        RECT 128.600 5.800 129.000 6.600 ;
        RECT 131.300 6.200 131.700 6.300 ;
        RECT 131.300 5.900 133.800 6.200 ;
        RECT 133.400 5.800 133.800 5.900 ;
        RECT 130.200 5.500 133.000 5.600 ;
        RECT 130.200 5.400 133.100 5.500 ;
        RECT 130.200 5.300 135.100 5.400 ;
        RECT 127.000 4.800 127.700 5.100 ;
        RECT 128.000 4.800 128.500 5.100 ;
        RECT 127.400 4.200 127.700 4.800 ;
        RECT 127.400 3.800 127.800 4.200 ;
        RECT 128.100 1.100 128.500 4.800 ;
        RECT 130.200 1.100 130.600 5.300 ;
        RECT 132.700 5.100 135.100 5.300 ;
        RECT 131.800 4.500 134.500 4.800 ;
        RECT 131.800 4.400 132.200 4.500 ;
        RECT 134.100 4.400 134.500 4.500 ;
        RECT 134.800 4.500 135.100 5.100 ;
        RECT 135.800 5.200 136.100 6.800 ;
        RECT 136.600 6.400 137.000 6.500 ;
        RECT 136.600 6.100 138.500 6.400 ;
        RECT 138.100 6.000 138.500 6.100 ;
        RECT 137.300 5.700 137.700 5.800 ;
        RECT 139.000 5.700 139.400 7.400 ;
        RECT 139.900 7.200 140.200 7.900 ;
        RECT 140.700 7.700 142.500 7.900 ;
        RECT 143.100 7.700 144.900 7.900 ;
        RECT 141.800 7.200 142.200 7.400 ;
        RECT 143.400 7.200 143.800 7.400 ;
        RECT 145.400 7.200 145.700 7.900 ;
        RECT 147.800 7.700 148.200 9.900 ;
        RECT 149.900 9.200 150.500 9.900 ;
        RECT 149.900 8.900 150.600 9.200 ;
        RECT 152.200 8.900 152.600 9.900 ;
        RECT 154.400 9.200 154.800 9.900 ;
        RECT 154.400 8.900 155.400 9.200 ;
        RECT 150.200 8.500 150.600 8.900 ;
        RECT 152.300 8.600 152.600 8.900 ;
        RECT 152.300 8.300 153.700 8.600 ;
        RECT 153.300 8.200 153.700 8.300 ;
        RECT 154.200 8.200 154.600 8.600 ;
        RECT 155.000 8.500 155.400 8.900 ;
        RECT 149.300 7.700 149.700 7.800 ;
        RECT 147.800 7.400 149.700 7.700 ;
        RECT 139.800 6.800 141.100 7.200 ;
        RECT 141.800 7.100 142.600 7.200 ;
        RECT 143.000 7.100 143.800 7.200 ;
        RECT 141.800 6.900 143.800 7.100 ;
        RECT 142.200 6.800 143.400 6.900 ;
        RECT 144.500 6.800 145.800 7.200 ;
        RECT 147.000 6.800 147.400 7.200 ;
        RECT 137.300 5.400 139.400 5.700 ;
        RECT 135.800 4.900 137.000 5.200 ;
        RECT 135.500 4.500 135.900 4.600 ;
        RECT 134.800 4.200 135.900 4.500 ;
        RECT 136.700 4.400 137.000 4.900 ;
        RECT 136.700 4.000 137.400 4.400 ;
        RECT 133.500 3.700 133.900 3.800 ;
        RECT 134.900 3.700 135.300 3.800 ;
        RECT 131.800 3.100 132.200 3.500 ;
        RECT 133.500 3.400 135.300 3.700 ;
        RECT 134.600 3.100 134.900 3.400 ;
        RECT 136.600 3.100 137.000 3.500 ;
        RECT 131.800 2.800 132.800 3.100 ;
        RECT 132.400 1.100 132.800 2.800 ;
        RECT 134.600 1.100 135.000 3.100 ;
        RECT 136.700 1.100 137.300 3.100 ;
        RECT 139.000 1.100 139.400 5.400 ;
        RECT 139.800 5.100 140.200 5.200 ;
        RECT 140.800 5.100 141.100 6.800 ;
        RECT 141.400 5.800 141.800 6.600 ;
        RECT 143.800 5.800 144.200 6.600 ;
        RECT 144.500 6.100 144.800 6.800 ;
        RECT 147.000 6.100 147.300 6.800 ;
        RECT 144.500 5.800 147.300 6.100 ;
        RECT 144.500 5.100 144.800 5.800 ;
        RECT 147.800 5.700 148.200 7.400 ;
        RECT 151.300 7.100 151.700 7.200 ;
        RECT 154.200 7.100 154.500 8.200 ;
        RECT 156.600 7.500 157.000 9.900 ;
        RECT 158.200 7.600 158.600 9.900 ;
        RECT 159.800 7.600 160.200 9.900 ;
        RECT 161.400 7.600 161.800 9.900 ;
        RECT 163.000 7.600 163.400 9.900 ;
        RECT 164.600 8.000 165.000 9.900 ;
        RECT 166.200 8.000 166.600 9.900 ;
        RECT 164.600 7.900 166.600 8.000 ;
        RECT 167.000 7.900 167.400 9.900 ;
        RECT 169.100 8.200 169.500 9.900 ;
        RECT 168.600 7.900 169.500 8.200 ;
        RECT 164.700 7.700 166.500 7.900 ;
        RECT 157.400 7.200 158.600 7.600 ;
        RECT 159.100 7.200 160.200 7.600 ;
        RECT 160.700 7.200 161.800 7.600 ;
        RECT 162.500 7.200 163.400 7.600 ;
        RECT 165.000 7.200 165.400 7.400 ;
        RECT 167.000 7.200 167.300 7.900 ;
        RECT 155.800 7.100 156.600 7.200 ;
        RECT 151.100 6.800 156.600 7.100 ;
        RECT 150.200 6.400 150.600 6.500 ;
        RECT 148.700 6.100 150.600 6.400 ;
        RECT 148.700 6.000 149.100 6.100 ;
        RECT 149.500 5.700 149.900 5.800 ;
        RECT 147.800 5.400 149.900 5.700 ;
        RECT 145.400 5.100 145.800 5.200 ;
        RECT 146.200 5.100 146.600 5.200 ;
        RECT 139.800 4.800 140.500 5.100 ;
        RECT 140.800 4.800 141.300 5.100 ;
        RECT 140.200 4.200 140.500 4.800 ;
        RECT 140.200 3.800 140.600 4.200 ;
        RECT 140.900 1.100 141.300 4.800 ;
        RECT 144.300 4.800 144.800 5.100 ;
        RECT 145.100 4.800 146.600 5.100 ;
        RECT 144.300 1.100 144.700 4.800 ;
        RECT 145.100 4.200 145.400 4.800 ;
        RECT 145.000 3.800 145.400 4.200 ;
        RECT 147.800 1.100 148.200 5.400 ;
        RECT 151.100 5.200 151.400 6.800 ;
        RECT 154.700 6.700 155.100 6.800 ;
        RECT 155.500 6.200 155.900 6.300 ;
        RECT 153.400 5.900 155.900 6.200 ;
        RECT 153.400 5.800 153.800 5.900 ;
        RECT 157.400 5.800 157.800 7.200 ;
        RECT 159.100 6.900 159.500 7.200 ;
        RECT 160.700 6.900 161.100 7.200 ;
        RECT 162.500 6.900 162.900 7.200 ;
        RECT 163.800 6.900 164.200 7.200 ;
        RECT 158.200 6.500 159.500 6.900 ;
        RECT 159.900 6.500 161.100 6.900 ;
        RECT 161.600 6.500 162.900 6.900 ;
        RECT 163.300 6.500 164.200 6.900 ;
        RECT 164.600 6.900 165.400 7.200 ;
        RECT 164.600 6.800 165.000 6.900 ;
        RECT 166.100 6.800 167.400 7.200 ;
        RECT 167.800 6.800 168.200 7.600 ;
        RECT 159.100 5.800 159.500 6.500 ;
        RECT 160.700 5.800 161.100 6.500 ;
        RECT 162.500 5.800 162.900 6.500 ;
        RECT 165.400 5.800 165.800 6.600 ;
        RECT 154.200 5.500 157.000 5.600 ;
        RECT 154.100 5.400 157.000 5.500 ;
        RECT 157.400 5.400 158.600 5.800 ;
        RECT 159.100 5.400 160.200 5.800 ;
        RECT 160.700 5.400 161.800 5.800 ;
        RECT 162.500 5.400 163.400 5.800 ;
        RECT 150.200 4.900 151.400 5.200 ;
        RECT 152.100 5.300 157.000 5.400 ;
        RECT 152.100 5.100 154.500 5.300 ;
        RECT 150.200 4.400 150.500 4.900 ;
        RECT 149.800 4.000 150.500 4.400 ;
        RECT 151.300 4.500 151.700 4.600 ;
        RECT 152.100 4.500 152.400 5.100 ;
        RECT 151.300 4.200 152.400 4.500 ;
        RECT 152.700 4.500 155.400 4.800 ;
        RECT 152.700 4.400 153.100 4.500 ;
        RECT 155.000 4.400 155.400 4.500 ;
        RECT 151.900 3.700 152.300 3.800 ;
        RECT 153.300 3.700 153.700 3.800 ;
        RECT 150.200 3.100 150.600 3.500 ;
        RECT 151.900 3.400 153.700 3.700 ;
        RECT 152.300 3.100 152.600 3.400 ;
        RECT 155.000 3.100 155.400 3.500 ;
        RECT 149.900 1.100 150.500 3.100 ;
        RECT 152.200 1.100 152.600 3.100 ;
        RECT 154.400 2.800 155.400 3.100 ;
        RECT 154.400 1.100 154.800 2.800 ;
        RECT 156.600 1.100 157.000 5.300 ;
        RECT 158.200 1.100 158.600 5.400 ;
        RECT 159.800 1.100 160.200 5.400 ;
        RECT 161.400 1.100 161.800 5.400 ;
        RECT 163.000 1.100 163.400 5.400 ;
        RECT 166.100 5.100 166.400 6.800 ;
        RECT 167.000 6.200 167.300 6.800 ;
        RECT 167.000 5.800 167.400 6.200 ;
        RECT 167.000 5.100 167.400 5.200 ;
        RECT 168.600 5.100 169.000 7.900 ;
        RECT 170.200 7.700 170.600 9.900 ;
        RECT 172.300 9.200 172.900 9.900 ;
        RECT 172.300 8.900 173.000 9.200 ;
        RECT 174.600 8.900 175.000 9.900 ;
        RECT 176.800 9.200 177.200 9.900 ;
        RECT 176.800 8.900 177.800 9.200 ;
        RECT 172.600 8.500 173.000 8.900 ;
        RECT 174.700 8.600 175.000 8.900 ;
        RECT 174.700 8.300 176.100 8.600 ;
        RECT 175.700 8.200 176.100 8.300 ;
        RECT 176.600 7.800 177.000 8.600 ;
        RECT 177.400 8.500 177.800 8.900 ;
        RECT 171.700 7.700 172.100 7.800 ;
        RECT 170.200 7.400 172.100 7.700 ;
        RECT 170.200 5.700 170.600 7.400 ;
        RECT 173.700 7.100 174.100 7.200 ;
        RECT 176.600 7.100 176.900 7.800 ;
        RECT 179.000 7.500 179.400 9.900 ;
        RECT 180.100 8.200 180.500 9.900 ;
        RECT 180.100 7.900 181.000 8.200 ;
        RECT 182.200 7.900 182.600 9.900 ;
        RECT 183.000 8.000 183.400 9.900 ;
        RECT 184.600 8.000 185.000 9.900 ;
        RECT 183.000 7.900 185.000 8.000 ;
        RECT 178.200 7.100 179.000 7.200 ;
        RECT 173.500 6.800 179.000 7.100 ;
        RECT 172.600 6.400 173.000 6.500 ;
        RECT 171.100 6.100 173.000 6.400 ;
        RECT 171.100 6.000 171.500 6.100 ;
        RECT 171.900 5.700 172.300 5.800 ;
        RECT 170.200 5.400 172.300 5.700 ;
        RECT 165.900 4.800 166.400 5.100 ;
        RECT 166.700 4.800 169.000 5.100 ;
        RECT 165.900 1.100 166.300 4.800 ;
        RECT 166.700 4.200 167.000 4.800 ;
        RECT 166.600 3.800 167.000 4.200 ;
        RECT 168.600 1.100 169.000 4.800 ;
        RECT 169.400 4.400 169.800 5.200 ;
        RECT 170.200 1.100 170.600 5.400 ;
        RECT 173.500 5.200 173.800 6.800 ;
        RECT 177.100 6.700 177.500 6.800 ;
        RECT 177.900 6.200 178.300 6.300 ;
        RECT 175.800 5.900 178.300 6.200 ;
        RECT 175.800 5.800 176.200 5.900 ;
        RECT 176.600 5.500 179.400 5.600 ;
        RECT 176.500 5.400 179.400 5.500 ;
        RECT 172.600 4.900 173.800 5.200 ;
        RECT 174.500 5.300 179.400 5.400 ;
        RECT 174.500 5.100 176.900 5.300 ;
        RECT 172.600 4.400 172.900 4.900 ;
        RECT 172.200 4.000 172.900 4.400 ;
        RECT 173.700 4.500 174.100 4.600 ;
        RECT 174.500 4.500 174.800 5.100 ;
        RECT 173.700 4.200 174.800 4.500 ;
        RECT 175.100 4.500 177.800 4.800 ;
        RECT 175.100 4.400 175.500 4.500 ;
        RECT 177.400 4.400 177.800 4.500 ;
        RECT 174.300 3.700 174.700 3.800 ;
        RECT 175.700 3.700 176.100 3.800 ;
        RECT 172.600 3.100 173.000 3.500 ;
        RECT 174.300 3.400 176.100 3.700 ;
        RECT 174.700 3.100 175.000 3.400 ;
        RECT 177.400 3.100 177.800 3.500 ;
        RECT 172.300 1.100 172.900 3.100 ;
        RECT 174.600 1.100 175.000 3.100 ;
        RECT 176.800 2.800 177.800 3.100 ;
        RECT 176.800 1.100 177.200 2.800 ;
        RECT 179.000 1.100 179.400 5.300 ;
        RECT 179.800 4.400 180.200 5.200 ;
        RECT 180.600 5.100 181.000 7.900 ;
        RECT 181.400 6.800 181.800 7.600 ;
        RECT 182.300 7.200 182.600 7.900 ;
        RECT 183.100 7.700 184.900 7.900 ;
        RECT 185.400 7.500 185.800 9.900 ;
        RECT 187.600 9.200 188.000 9.900 ;
        RECT 187.000 8.900 188.000 9.200 ;
        RECT 189.800 8.900 190.200 9.900 ;
        RECT 191.900 9.200 192.500 9.900 ;
        RECT 191.800 8.900 192.500 9.200 ;
        RECT 187.000 8.500 187.400 8.900 ;
        RECT 189.800 8.600 190.100 8.900 ;
        RECT 187.800 8.200 188.200 8.600 ;
        RECT 188.700 8.300 190.100 8.600 ;
        RECT 191.800 8.500 192.200 8.900 ;
        RECT 188.700 8.200 189.100 8.300 ;
        RECT 184.200 7.200 184.600 7.400 ;
        RECT 182.200 6.800 183.500 7.200 ;
        RECT 184.200 6.900 185.000 7.200 ;
        RECT 184.600 6.800 185.000 6.900 ;
        RECT 185.800 7.100 186.600 7.200 ;
        RECT 187.900 7.100 188.200 8.200 ;
        RECT 192.700 7.700 193.100 7.800 ;
        RECT 194.200 7.700 194.600 9.900 ;
        RECT 195.000 8.000 195.400 9.900 ;
        RECT 196.600 8.000 197.000 9.900 ;
        RECT 195.000 7.900 197.000 8.000 ;
        RECT 197.400 7.900 197.800 9.900 ;
        RECT 198.500 8.200 198.900 9.900 ;
        RECT 198.500 7.900 199.400 8.200 ;
        RECT 195.100 7.700 196.900 7.900 ;
        RECT 192.700 7.400 194.600 7.700 ;
        RECT 189.400 7.100 189.800 7.200 ;
        RECT 190.700 7.100 191.100 7.200 ;
        RECT 185.800 6.800 191.300 7.100 ;
        RECT 183.200 5.200 183.500 6.800 ;
        RECT 187.300 6.700 187.700 6.800 ;
        RECT 183.800 5.800 184.200 6.600 ;
        RECT 186.500 6.200 186.900 6.300 ;
        RECT 187.800 6.200 188.200 6.300 ;
        RECT 186.500 5.900 189.000 6.200 ;
        RECT 188.600 5.800 189.000 5.900 ;
        RECT 185.400 5.500 188.200 5.600 ;
        RECT 185.400 5.400 188.300 5.500 ;
        RECT 185.400 5.300 190.300 5.400 ;
        RECT 182.200 5.100 182.600 5.200 ;
        RECT 180.600 4.800 182.900 5.100 ;
        RECT 183.200 4.800 184.200 5.200 ;
        RECT 180.600 1.100 181.000 4.800 ;
        RECT 182.600 4.200 182.900 4.800 ;
        RECT 182.600 3.800 183.000 4.200 ;
        RECT 183.300 1.100 183.700 4.800 ;
        RECT 185.400 1.100 185.800 5.300 ;
        RECT 187.900 5.100 190.300 5.300 ;
        RECT 187.000 4.500 189.700 4.800 ;
        RECT 187.000 4.400 187.400 4.500 ;
        RECT 189.300 4.400 189.700 4.500 ;
        RECT 190.000 4.500 190.300 5.100 ;
        RECT 191.000 5.200 191.300 6.800 ;
        RECT 191.800 6.400 192.200 6.500 ;
        RECT 191.800 6.100 193.700 6.400 ;
        RECT 193.300 6.000 193.700 6.100 ;
        RECT 192.500 5.700 192.900 5.800 ;
        RECT 194.200 5.700 194.600 7.400 ;
        RECT 195.400 7.200 195.800 7.400 ;
        RECT 197.400 7.200 197.700 7.900 ;
        RECT 195.000 6.900 195.800 7.200 ;
        RECT 196.500 7.100 197.800 7.200 ;
        RECT 198.200 7.100 198.600 7.200 ;
        RECT 195.000 6.800 195.400 6.900 ;
        RECT 196.500 6.800 198.600 7.100 ;
        RECT 195.800 5.800 196.200 6.600 ;
        RECT 192.500 5.400 194.600 5.700 ;
        RECT 191.000 4.900 192.200 5.200 ;
        RECT 190.700 4.500 191.100 4.600 ;
        RECT 190.000 4.200 191.100 4.500 ;
        RECT 191.900 4.400 192.200 4.900 ;
        RECT 191.900 4.000 192.600 4.400 ;
        RECT 188.700 3.700 189.100 3.800 ;
        RECT 190.100 3.700 190.500 3.800 ;
        RECT 187.000 3.100 187.400 3.500 ;
        RECT 188.700 3.400 190.500 3.700 ;
        RECT 189.800 3.100 190.100 3.400 ;
        RECT 191.800 3.100 192.200 3.500 ;
        RECT 187.000 2.800 188.000 3.100 ;
        RECT 187.600 1.100 188.000 2.800 ;
        RECT 189.800 1.100 190.200 3.100 ;
        RECT 191.900 1.100 192.500 3.100 ;
        RECT 194.200 1.100 194.600 5.400 ;
        RECT 196.500 5.100 196.800 6.800 ;
        RECT 199.000 6.100 199.400 7.900 ;
        RECT 199.800 7.100 200.200 7.600 ;
        RECT 202.200 7.500 202.600 9.900 ;
        RECT 204.400 9.200 204.800 9.900 ;
        RECT 203.800 8.900 204.800 9.200 ;
        RECT 206.600 8.900 207.000 9.900 ;
        RECT 208.700 9.200 209.300 9.900 ;
        RECT 208.600 8.900 209.300 9.200 ;
        RECT 203.800 8.500 204.200 8.900 ;
        RECT 206.600 8.600 206.900 8.900 ;
        RECT 204.600 8.200 205.000 8.600 ;
        RECT 205.500 8.300 206.900 8.600 ;
        RECT 208.600 8.500 209.000 8.900 ;
        RECT 205.500 8.200 205.900 8.300 ;
        RECT 200.600 7.100 201.000 7.200 ;
        RECT 199.800 6.800 201.000 7.100 ;
        RECT 202.600 7.100 203.400 7.200 ;
        RECT 204.700 7.100 205.000 8.200 ;
        RECT 209.500 7.700 209.900 7.800 ;
        RECT 211.000 7.700 211.400 9.900 ;
        RECT 209.500 7.400 211.400 7.700 ;
        RECT 211.800 7.500 212.200 9.900 ;
        RECT 214.000 9.200 214.400 9.900 ;
        RECT 213.400 8.900 214.400 9.200 ;
        RECT 216.200 8.900 216.600 9.900 ;
        RECT 218.300 9.200 218.900 9.900 ;
        RECT 218.200 8.900 218.900 9.200 ;
        RECT 213.400 8.500 213.800 8.900 ;
        RECT 216.200 8.600 216.500 8.900 ;
        RECT 214.200 8.200 214.600 8.600 ;
        RECT 215.100 8.300 216.500 8.600 ;
        RECT 218.200 8.500 218.600 8.900 ;
        RECT 215.100 8.200 215.500 8.300 ;
        RECT 206.200 7.100 206.600 7.200 ;
        RECT 207.500 7.100 207.900 7.200 ;
        RECT 202.600 6.800 208.100 7.100 ;
        RECT 204.100 6.700 204.500 6.800 ;
        RECT 197.400 5.800 199.400 6.100 ;
        RECT 203.300 6.200 203.700 6.300 ;
        RECT 204.600 6.200 205.000 6.300 ;
        RECT 203.300 5.900 205.800 6.200 ;
        RECT 205.400 5.800 205.800 5.900 ;
        RECT 197.400 5.200 197.700 5.800 ;
        RECT 197.400 5.100 197.800 5.200 ;
        RECT 196.300 4.800 196.800 5.100 ;
        RECT 197.100 4.800 197.800 5.100 ;
        RECT 196.300 1.100 196.700 4.800 ;
        RECT 197.100 4.200 197.400 4.800 ;
        RECT 198.200 4.400 198.600 5.200 ;
        RECT 197.000 3.800 197.400 4.200 ;
        RECT 199.000 1.100 199.400 5.800 ;
        RECT 202.200 5.500 205.000 5.600 ;
        RECT 202.200 5.400 205.100 5.500 ;
        RECT 202.200 5.300 207.100 5.400 ;
        RECT 202.200 1.100 202.600 5.300 ;
        RECT 204.700 5.100 207.100 5.300 ;
        RECT 203.800 4.500 206.500 4.800 ;
        RECT 203.800 4.400 204.200 4.500 ;
        RECT 206.100 4.400 206.500 4.500 ;
        RECT 206.800 4.500 207.100 5.100 ;
        RECT 207.800 5.200 208.100 6.800 ;
        RECT 208.600 6.400 209.000 6.500 ;
        RECT 208.600 6.100 210.500 6.400 ;
        RECT 210.100 6.000 210.500 6.100 ;
        RECT 209.300 5.700 209.700 5.800 ;
        RECT 211.000 5.700 211.400 7.400 ;
        RECT 212.200 7.100 213.000 7.200 ;
        RECT 214.300 7.100 214.600 8.200 ;
        RECT 219.100 7.700 219.500 7.800 ;
        RECT 220.600 7.700 221.000 9.900 ;
        RECT 221.400 8.000 221.800 9.900 ;
        RECT 223.000 8.000 223.400 9.900 ;
        RECT 221.400 7.900 223.400 8.000 ;
        RECT 223.800 7.900 224.200 9.900 ;
        RECT 224.900 8.200 225.300 9.900 ;
        RECT 224.900 7.900 225.800 8.200 ;
        RECT 221.500 7.700 223.300 7.900 ;
        RECT 219.100 7.400 221.000 7.700 ;
        RECT 215.800 7.100 216.200 7.200 ;
        RECT 217.100 7.100 217.500 7.200 ;
        RECT 212.200 6.800 217.700 7.100 ;
        RECT 213.700 6.700 214.100 6.800 ;
        RECT 212.900 6.200 213.300 6.300 ;
        RECT 212.900 6.100 215.400 6.200 ;
        RECT 216.600 6.100 217.000 6.200 ;
        RECT 212.900 5.900 217.000 6.100 ;
        RECT 215.000 5.800 217.000 5.900 ;
        RECT 209.300 5.400 211.400 5.700 ;
        RECT 207.800 4.900 209.000 5.200 ;
        RECT 207.500 4.500 207.900 4.600 ;
        RECT 206.800 4.200 207.900 4.500 ;
        RECT 208.700 4.400 209.000 4.900 ;
        RECT 208.700 4.000 209.400 4.400 ;
        RECT 205.500 3.700 205.900 3.800 ;
        RECT 206.900 3.700 207.300 3.800 ;
        RECT 203.800 3.100 204.200 3.500 ;
        RECT 205.500 3.400 207.300 3.700 ;
        RECT 206.600 3.100 206.900 3.400 ;
        RECT 208.600 3.100 209.000 3.500 ;
        RECT 203.800 2.800 204.800 3.100 ;
        RECT 204.400 1.100 204.800 2.800 ;
        RECT 206.600 1.100 207.000 3.100 ;
        RECT 208.700 1.100 209.300 3.100 ;
        RECT 211.000 1.100 211.400 5.400 ;
        RECT 211.800 5.500 214.600 5.600 ;
        RECT 211.800 5.400 214.700 5.500 ;
        RECT 211.800 5.300 216.700 5.400 ;
        RECT 211.800 1.100 212.200 5.300 ;
        RECT 214.300 5.100 216.700 5.300 ;
        RECT 213.400 4.500 216.100 4.800 ;
        RECT 213.400 4.400 213.800 4.500 ;
        RECT 215.700 4.400 216.100 4.500 ;
        RECT 216.400 4.500 216.700 5.100 ;
        RECT 217.400 5.200 217.700 6.800 ;
        RECT 218.200 6.400 218.600 6.500 ;
        RECT 218.200 6.100 220.100 6.400 ;
        RECT 219.700 6.000 220.100 6.100 ;
        RECT 218.900 5.700 219.300 5.800 ;
        RECT 220.600 5.700 221.000 7.400 ;
        RECT 221.800 7.200 222.200 7.400 ;
        RECT 223.800 7.200 224.100 7.900 ;
        RECT 221.400 6.900 222.200 7.200 ;
        RECT 222.900 7.100 224.200 7.200 ;
        RECT 224.600 7.100 225.000 7.200 ;
        RECT 221.400 6.800 221.800 6.900 ;
        RECT 222.900 6.800 225.000 7.100 ;
        RECT 222.200 5.800 222.600 6.600 ;
        RECT 218.900 5.400 221.000 5.700 ;
        RECT 217.400 4.900 218.600 5.200 ;
        RECT 217.100 4.500 217.500 4.600 ;
        RECT 216.400 4.200 217.500 4.500 ;
        RECT 218.300 4.400 218.600 4.900 ;
        RECT 218.300 4.000 219.000 4.400 ;
        RECT 215.100 3.700 215.500 3.800 ;
        RECT 216.500 3.700 216.900 3.800 ;
        RECT 213.400 3.100 213.800 3.500 ;
        RECT 215.100 3.400 216.900 3.700 ;
        RECT 216.200 3.100 216.500 3.400 ;
        RECT 218.200 3.100 218.600 3.500 ;
        RECT 213.400 2.800 214.400 3.100 ;
        RECT 214.000 1.100 214.400 2.800 ;
        RECT 216.200 1.100 216.600 3.100 ;
        RECT 218.300 1.100 218.900 3.100 ;
        RECT 220.600 1.100 221.000 5.400 ;
        RECT 222.900 5.100 223.200 6.800 ;
        RECT 225.400 6.100 225.800 7.900 ;
        RECT 227.000 7.700 227.400 9.900 ;
        RECT 229.100 9.200 229.700 9.900 ;
        RECT 229.100 8.900 229.800 9.200 ;
        RECT 231.400 8.900 231.800 9.900 ;
        RECT 233.600 9.200 234.000 9.900 ;
        RECT 233.600 8.900 234.600 9.200 ;
        RECT 229.400 8.500 229.800 8.900 ;
        RECT 231.500 8.600 231.800 8.900 ;
        RECT 231.500 8.300 232.900 8.600 ;
        RECT 232.500 8.200 232.900 8.300 ;
        RECT 233.400 8.200 233.800 8.600 ;
        RECT 234.200 8.500 234.600 8.900 ;
        RECT 228.500 7.700 228.900 7.800 ;
        RECT 226.200 7.100 226.600 7.600 ;
        RECT 227.000 7.400 228.900 7.700 ;
        RECT 227.000 7.100 227.400 7.400 ;
        RECT 230.500 7.100 230.900 7.200 ;
        RECT 233.400 7.100 233.700 8.200 ;
        RECT 235.800 7.500 236.200 9.900 ;
        RECT 237.400 7.600 237.800 9.900 ;
        RECT 239.000 7.600 239.400 9.900 ;
        RECT 240.600 7.600 241.000 9.900 ;
        RECT 242.200 7.600 242.600 9.900 ;
        RECT 244.600 7.600 245.000 9.900 ;
        RECT 246.200 7.600 246.600 9.900 ;
        RECT 237.400 7.200 238.300 7.600 ;
        RECT 239.000 7.200 240.100 7.600 ;
        RECT 240.600 7.200 241.700 7.600 ;
        RECT 242.200 7.200 243.400 7.600 ;
        RECT 235.000 7.100 235.800 7.200 ;
        RECT 226.200 6.800 227.400 7.100 ;
        RECT 223.800 5.800 225.800 6.100 ;
        RECT 223.800 5.200 224.100 5.800 ;
        RECT 223.800 5.100 224.200 5.200 ;
        RECT 222.700 4.800 223.200 5.100 ;
        RECT 223.500 4.800 224.200 5.100 ;
        RECT 222.700 1.100 223.100 4.800 ;
        RECT 223.500 4.200 223.800 4.800 ;
        RECT 224.600 4.400 225.000 5.200 ;
        RECT 223.400 3.800 223.800 4.200 ;
        RECT 225.400 1.100 225.800 5.800 ;
        RECT 227.000 5.700 227.400 6.800 ;
        RECT 230.300 6.800 235.800 7.100 ;
        RECT 237.900 6.900 238.300 7.200 ;
        RECT 239.700 6.900 240.100 7.200 ;
        RECT 241.300 6.900 241.700 7.200 ;
        RECT 229.400 6.400 229.800 6.500 ;
        RECT 227.900 6.100 229.800 6.400 ;
        RECT 227.900 6.000 228.300 6.100 ;
        RECT 228.700 5.700 229.100 5.800 ;
        RECT 227.000 5.400 229.100 5.700 ;
        RECT 227.000 1.100 227.400 5.400 ;
        RECT 230.300 5.200 230.600 6.800 ;
        RECT 233.900 6.700 234.300 6.800 ;
        RECT 237.900 6.500 239.200 6.900 ;
        RECT 239.700 6.500 240.900 6.900 ;
        RECT 241.300 6.500 242.600 6.900 ;
        RECT 234.700 6.200 235.100 6.300 ;
        RECT 232.600 5.900 235.100 6.200 ;
        RECT 232.600 5.800 233.000 5.900 ;
        RECT 237.900 5.800 238.300 6.500 ;
        RECT 239.700 5.800 240.100 6.500 ;
        RECT 241.300 5.800 241.700 6.500 ;
        RECT 243.000 5.800 243.400 7.200 ;
        RECT 233.400 5.500 236.200 5.600 ;
        RECT 233.300 5.400 236.200 5.500 ;
        RECT 229.400 4.900 230.600 5.200 ;
        RECT 231.300 5.300 236.200 5.400 ;
        RECT 231.300 5.100 233.700 5.300 ;
        RECT 229.400 4.400 229.700 4.900 ;
        RECT 229.000 4.000 229.700 4.400 ;
        RECT 230.500 4.500 230.900 4.600 ;
        RECT 231.300 4.500 231.600 5.100 ;
        RECT 230.500 4.200 231.600 4.500 ;
        RECT 231.900 4.500 234.600 4.800 ;
        RECT 231.900 4.400 232.300 4.500 ;
        RECT 234.200 4.400 234.600 4.500 ;
        RECT 231.100 3.700 231.500 3.800 ;
        RECT 232.500 3.700 232.900 3.800 ;
        RECT 229.400 3.100 229.800 3.500 ;
        RECT 231.100 3.400 232.900 3.700 ;
        RECT 231.500 3.100 231.800 3.400 ;
        RECT 234.200 3.100 234.600 3.500 ;
        RECT 229.100 1.100 229.700 3.100 ;
        RECT 231.400 1.100 231.800 3.100 ;
        RECT 233.600 2.800 234.600 3.100 ;
        RECT 233.600 1.100 234.000 2.800 ;
        RECT 235.800 1.100 236.200 5.300 ;
        RECT 237.400 5.400 238.300 5.800 ;
        RECT 239.000 5.400 240.100 5.800 ;
        RECT 240.600 5.400 241.700 5.800 ;
        RECT 242.200 5.400 243.400 5.800 ;
        RECT 244.600 7.200 246.600 7.600 ;
        RECT 248.600 7.600 249.000 9.900 ;
        RECT 250.200 7.600 250.600 9.900 ;
        RECT 248.600 7.200 250.600 7.600 ;
        RECT 244.600 5.800 245.000 7.200 ;
        RECT 248.600 5.800 249.000 7.200 ;
        RECT 244.600 5.400 246.600 5.800 ;
        RECT 237.400 1.100 237.800 5.400 ;
        RECT 239.000 1.100 239.400 5.400 ;
        RECT 240.600 1.100 241.000 5.400 ;
        RECT 242.200 1.100 242.600 5.400 ;
        RECT 244.600 1.100 245.000 5.400 ;
        RECT 246.200 1.100 246.600 5.400 ;
        RECT 248.600 5.400 250.600 5.800 ;
        RECT 248.600 1.100 249.000 5.400 ;
        RECT 250.200 1.100 250.600 5.400 ;
      LAYER via1 ;
        RECT 0.600 232.800 1.000 233.200 ;
        RECT 7.000 234.800 7.400 235.200 ;
        RECT 9.400 233.800 9.800 234.200 ;
        RECT 11.000 233.800 11.400 234.200 ;
        RECT 19.000 236.200 19.400 236.600 ;
        RECT 20.600 235.500 21.000 235.900 ;
        RECT 3.800 231.800 4.200 232.200 ;
        RECT 21.400 233.800 21.800 234.200 ;
        RECT 22.200 233.800 22.600 234.200 ;
        RECT 20.600 233.100 21.000 233.500 ;
        RECT 29.400 234.800 29.800 235.200 ;
        RECT 31.800 233.800 32.200 234.200 ;
        RECT 33.400 233.800 33.800 234.200 ;
        RECT 27.000 231.800 27.400 232.200 ;
        RECT 34.200 233.100 34.600 233.500 ;
        RECT 43.000 231.800 43.400 232.200 ;
        RECT 52.600 236.200 53.000 236.600 ;
        RECT 54.200 235.500 54.600 235.900 ;
        RECT 55.000 233.800 55.400 234.200 ;
        RECT 54.200 233.100 54.600 233.500 ;
        RECT 45.400 231.800 45.800 232.200 ;
        RECT 70.200 236.800 70.600 237.200 ;
        RECT 59.000 234.800 59.400 235.200 ;
        RECT 63.800 234.800 64.200 235.200 ;
        RECT 59.800 233.800 60.200 234.200 ;
        RECT 60.600 233.100 61.000 233.500 ;
        RECT 74.200 236.800 74.600 237.200 ;
        RECT 70.200 233.800 70.600 234.200 ;
        RECT 63.000 232.800 63.400 233.200 ;
        RECT 74.200 234.800 74.600 235.200 ;
        RECT 75.000 233.800 75.400 234.200 ;
        RECT 83.000 236.200 83.400 236.600 ;
        RECT 84.600 235.500 85.000 235.900 ;
        RECT 84.600 233.100 85.000 233.500 ;
        RECT 75.800 231.800 76.200 232.200 ;
        RECT 90.200 234.800 90.600 235.200 ;
        RECT 104.600 234.800 105.000 235.200 ;
        RECT 113.400 237.800 113.800 238.200 ;
        RECT 98.200 233.800 98.600 234.200 ;
        RECT 100.600 233.800 101.000 234.200 ;
        RECT 87.000 231.800 87.400 232.200 ;
        RECT 99.800 233.100 100.200 233.500 ;
        RECT 126.200 236.800 126.600 237.200 ;
        RECT 110.200 234.800 110.600 235.200 ;
        RECT 111.000 234.800 111.400 235.200 ;
        RECT 119.800 234.800 120.200 235.200 ;
        RECT 117.400 233.800 117.800 234.200 ;
        RECT 108.600 231.800 109.000 232.200 ;
        RECT 113.400 231.800 113.800 232.200 ;
        RECT 116.600 233.100 117.000 233.500 ;
        RECT 126.200 233.800 126.600 234.200 ;
        RECT 130.200 234.800 130.600 235.200 ;
        RECT 132.600 234.800 133.000 235.200 ;
        RECT 131.800 233.800 132.200 234.200 ;
        RECT 142.200 234.800 142.600 235.200 ;
        RECT 136.600 233.800 137.000 234.200 ;
        RECT 134.200 231.800 134.600 232.200 ;
        RECT 137.400 233.100 137.800 233.500 ;
        RECT 146.200 231.800 146.600 232.200 ;
        RECT 155.800 234.800 156.200 235.200 ;
        RECT 159.800 233.800 160.200 234.200 ;
        RECT 148.600 231.800 149.000 232.200 ;
        RECT 153.400 232.800 153.800 233.200 ;
        RECT 161.400 233.800 161.800 234.200 ;
        RECT 169.400 236.200 169.800 236.600 ;
        RECT 171.000 235.500 171.400 235.900 ;
        RECT 179.000 236.200 179.400 236.600 ;
        RECT 180.600 235.500 181.000 235.900 ;
        RECT 184.600 234.800 185.000 235.200 ;
        RECT 205.400 236.800 205.800 237.200 ;
        RECT 171.000 233.100 171.400 233.500 ;
        RECT 180.600 233.100 181.000 233.500 ;
        RECT 171.800 231.800 172.200 232.200 ;
        RECT 181.400 233.100 181.800 233.500 ;
        RECT 191.800 234.800 192.200 235.200 ;
        RECT 199.000 234.800 199.400 235.200 ;
        RECT 194.200 233.100 194.600 233.500 ;
        RECT 190.200 231.800 190.600 232.200 ;
        RECT 205.400 233.800 205.800 234.200 ;
        RECT 209.400 234.800 209.800 235.200 ;
        RECT 210.200 233.800 210.600 234.200 ;
        RECT 211.000 233.100 211.400 233.500 ;
        RECT 226.200 234.800 226.600 235.200 ;
        RECT 222.200 233.800 222.600 234.200 ;
        RECT 223.800 233.800 224.200 234.200 ;
        RECT 219.800 231.800 220.200 232.200 ;
        RECT 223.000 233.100 223.400 233.500 ;
        RECT 221.400 231.800 221.800 232.200 ;
        RECT 235.800 234.800 236.200 235.200 ;
        RECT 233.400 233.800 233.800 234.200 ;
        RECT 231.800 231.800 232.200 232.200 ;
        RECT 232.600 233.100 233.000 233.500 ;
        RECT 241.400 231.800 241.800 232.200 ;
        RECT 247.000 234.800 247.400 235.200 ;
        RECT 251.000 233.800 251.400 234.200 ;
        RECT 244.600 231.800 245.000 232.200 ;
        RECT 248.600 231.800 249.000 232.200 ;
        RECT 0.600 228.800 1.000 229.200 ;
        RECT 8.600 226.800 9.000 227.200 ;
        RECT 3.000 226.100 3.400 226.500 ;
        RECT 16.600 226.800 17.000 227.200 ;
        RECT 19.800 226.800 20.200 227.200 ;
        RECT 9.400 225.100 9.800 225.500 ;
        RECT 0.600 221.800 1.000 222.200 ;
        RECT 11.000 221.800 11.400 222.200 ;
        RECT 31.800 228.800 32.200 229.200 ;
        RECT 25.400 225.900 25.800 226.300 ;
        RECT 20.600 224.800 21.000 225.200 ;
        RECT 23.000 225.100 23.400 225.500 ;
        RECT 40.600 226.800 41.000 227.200 ;
        RECT 35.800 225.800 36.200 226.200 ;
        RECT 51.800 228.800 52.200 229.200 ;
        RECT 43.800 226.800 44.200 227.200 ;
        RECT 45.400 225.900 45.800 226.300 ;
        RECT 40.600 224.800 41.000 225.200 ;
        RECT 43.000 225.100 43.400 225.500 ;
        RECT 57.400 226.800 57.800 227.200 ;
        RECT 58.200 225.800 58.600 226.200 ;
        RECT 75.800 228.800 76.200 229.200 ;
        RECT 62.200 225.800 62.600 226.200 ;
        RECT 68.600 226.800 69.000 227.200 ;
        RECT 67.800 225.800 68.200 226.200 ;
        RECT 83.800 226.800 84.200 227.200 ;
        RECT 78.200 226.100 78.600 226.500 ;
        RECT 82.200 225.900 82.600 226.300 ;
        RECT 61.400 221.800 61.800 222.200 ;
        RECT 66.200 221.800 66.600 222.200 ;
        RECT 84.600 225.100 85.000 225.500 ;
        RECT 97.400 228.800 97.800 229.200 ;
        RECT 91.000 225.800 91.400 226.200 ;
        RECT 91.800 225.800 92.200 226.200 ;
        RECT 87.000 224.800 87.400 225.200 ;
        RECT 103.800 226.800 104.200 227.200 ;
        RECT 99.800 226.100 100.200 226.500 ;
        RECT 93.400 221.800 93.800 222.200 ;
        RECT 109.400 225.800 109.800 226.200 ;
        RECT 106.200 225.100 106.600 225.500 ;
        RECT 119.000 228.800 119.400 229.200 ;
        RECT 111.800 224.800 112.200 225.200 ;
        RECT 115.000 225.800 115.400 226.200 ;
        RECT 117.400 225.800 117.800 226.200 ;
        RECT 119.800 226.800 120.200 227.200 ;
        RECT 120.600 225.800 121.000 226.200 ;
        RECT 114.200 221.800 114.600 222.200 ;
        RECT 121.400 224.800 121.800 225.200 ;
        RECT 128.600 228.800 129.000 229.200 ;
        RECT 136.600 226.800 137.000 227.200 ;
        RECT 131.000 226.100 131.400 226.500 ;
        RECT 135.000 225.900 135.400 226.300 ;
        RECT 137.400 225.100 137.800 225.500 ;
        RECT 150.200 228.800 150.600 229.200 ;
        RECT 144.600 225.800 145.000 226.200 ;
        RECT 143.000 224.800 143.400 225.200 ;
        RECT 148.600 225.800 149.000 226.200 ;
        RECT 158.200 226.800 158.600 227.200 ;
        RECT 160.600 226.800 161.000 227.200 ;
        RECT 152.600 226.100 153.000 226.500 ;
        RECT 181.400 228.800 181.800 229.200 ;
        RECT 163.000 225.800 163.400 226.200 ;
        RECT 159.000 225.100 159.400 225.500 ;
        RECT 175.800 226.800 176.200 227.200 ;
        RECT 175.000 225.900 175.400 226.300 ;
        RECT 166.200 221.800 166.600 222.200 ;
        RECT 172.600 225.100 173.000 225.500 ;
        RECT 189.400 227.800 189.800 228.200 ;
        RECT 199.000 228.800 199.400 229.200 ;
        RECT 186.200 225.800 186.600 226.200 ;
        RECT 187.800 225.800 188.200 226.200 ;
        RECT 184.600 221.800 185.000 222.200 ;
        RECT 195.000 225.800 195.400 226.200 ;
        RECT 199.800 224.800 200.200 225.200 ;
        RECT 210.200 226.800 210.600 227.200 ;
        RECT 208.600 225.900 209.000 226.300 ;
        RECT 205.400 224.800 205.800 225.200 ;
        RECT 206.200 225.100 206.600 225.500 ;
        RECT 215.000 221.800 215.400 222.200 ;
        RECT 219.000 225.800 219.400 226.200 ;
        RECT 228.600 226.800 229.000 227.200 ;
        RECT 218.200 221.800 218.600 222.200 ;
        RECT 228.600 224.800 229.000 225.200 ;
        RECT 239.000 226.800 239.400 227.200 ;
        RECT 233.400 226.100 233.800 226.500 ;
        RECT 243.000 226.100 243.400 226.500 ;
        RECT 247.000 225.900 247.400 226.300 ;
        RECT 239.800 225.100 240.200 225.500 ;
        RECT 249.400 225.100 249.800 225.500 ;
        RECT 240.600 221.800 241.000 222.200 ;
        RECT 0.600 218.800 1.000 219.200 ;
        RECT 7.800 216.200 8.200 216.600 ;
        RECT 9.400 215.500 9.800 215.900 ;
        RECT 11.000 214.800 11.400 215.200 ;
        RECT 11.800 214.800 12.200 215.200 ;
        RECT 9.400 213.100 9.800 213.500 ;
        RECT 15.000 213.800 15.400 214.200 ;
        RECT 16.600 213.800 17.000 214.200 ;
        RECT 15.800 213.100 16.200 213.500 ;
        RECT 35.800 216.800 36.200 217.200 ;
        RECT 28.600 214.800 29.000 215.200 ;
        RECT 29.400 214.800 29.800 215.200 ;
        RECT 24.600 211.800 25.000 212.200 ;
        RECT 27.800 211.800 28.200 212.200 ;
        RECT 31.800 212.800 32.200 213.200 ;
        RECT 33.400 211.800 33.800 212.200 ;
        RECT 43.000 216.200 43.400 216.600 ;
        RECT 44.600 215.500 45.000 215.900 ;
        RECT 39.800 214.800 40.200 215.200 ;
        RECT 56.600 216.200 57.000 216.600 ;
        RECT 58.200 215.500 58.600 215.900 ;
        RECT 44.600 213.100 45.000 213.500 ;
        RECT 66.200 216.200 66.600 216.600 ;
        RECT 70.200 216.800 70.600 217.200 ;
        RECT 67.800 215.500 68.200 215.900 ;
        RECT 70.200 214.800 70.600 215.200 ;
        RECT 58.200 213.100 58.600 213.500 ;
        RECT 49.400 211.800 49.800 212.200 ;
        RECT 67.800 213.100 68.200 213.500 ;
        RECT 71.000 213.800 71.400 214.200 ;
        RECT 59.000 211.800 59.400 212.200 ;
        RECT 73.400 211.800 73.800 212.200 ;
        RECT 80.600 214.800 81.000 215.200 ;
        RECT 84.600 214.800 85.000 215.200 ;
        RECT 81.400 213.100 81.800 213.500 ;
        RECT 91.800 214.800 92.200 215.200 ;
        RECT 94.200 213.800 94.600 214.200 ;
        RECT 107.000 218.800 107.400 219.200 ;
        RECT 99.800 214.800 100.200 215.200 ;
        RECT 101.400 214.800 101.800 215.200 ;
        RECT 104.600 214.800 105.000 215.200 ;
        RECT 90.200 211.800 90.600 212.200 ;
        RECT 105.400 213.800 105.800 214.200 ;
        RECT 108.600 216.800 109.000 217.200 ;
        RECT 115.800 216.200 116.200 216.600 ;
        RECT 117.400 215.500 117.800 215.900 ;
        RECT 103.000 211.800 103.400 212.200 ;
        RECT 117.400 213.100 117.800 213.500 ;
        RECT 120.600 218.800 121.000 219.200 ;
        RECT 127.800 216.200 128.200 216.600 ;
        RECT 129.400 215.500 129.800 215.900 ;
        RECT 124.600 214.800 125.000 215.200 ;
        RECT 131.000 214.800 131.400 215.200 ;
        RECT 119.800 211.800 120.200 212.200 ;
        RECT 133.400 213.800 133.800 214.200 ;
        RECT 129.400 213.100 129.800 213.500 ;
        RECT 135.000 213.800 135.400 214.200 ;
        RECT 136.600 213.800 137.000 214.200 ;
        RECT 135.800 213.100 136.200 213.500 ;
        RECT 144.600 211.800 145.000 212.200 ;
        RECT 152.600 216.200 153.000 216.600 ;
        RECT 154.200 215.500 154.600 215.900 ;
        RECT 157.400 214.800 157.800 215.200 ;
        RECT 154.200 213.100 154.600 213.500 ;
        RECT 163.000 214.800 163.400 215.200 ;
        RECT 161.400 213.800 161.800 214.200 ;
        RECT 165.400 213.800 165.800 214.200 ;
        RECT 178.200 218.800 178.600 219.200 ;
        RECT 167.000 213.800 167.400 214.200 ;
        RECT 168.600 213.800 169.000 214.200 ;
        RECT 145.400 211.800 145.800 212.200 ;
        RECT 159.000 211.800 159.400 212.200 ;
        RECT 167.800 213.100 168.200 213.500 ;
        RECT 179.800 214.800 180.200 215.200 ;
        RECT 176.600 211.800 177.000 212.200 ;
        RECT 183.000 218.800 183.400 219.200 ;
        RECT 190.200 216.200 190.600 216.600 ;
        RECT 191.800 215.500 192.200 215.900 ;
        RECT 198.200 217.800 198.600 218.200 ;
        RECT 182.200 211.800 182.600 212.200 ;
        RECT 191.800 213.100 192.200 213.500 ;
        RECT 205.400 214.800 205.800 215.200 ;
        RECT 215.800 218.800 216.200 219.200 ;
        RECT 221.400 215.800 221.800 216.200 ;
        RECT 207.800 213.800 208.200 214.200 ;
        RECT 209.400 213.800 209.800 214.200 ;
        RECT 221.400 214.800 221.800 215.200 ;
        RECT 219.000 213.800 219.400 214.200 ;
        RECT 222.200 213.800 222.600 214.200 ;
        RECT 223.800 213.800 224.200 214.200 ;
        RECT 223.000 213.100 223.400 213.500 ;
        RECT 234.200 214.800 234.600 215.200 ;
        RECT 239.800 218.800 240.200 219.200 ;
        RECT 233.400 213.800 233.800 214.200 ;
        RECT 235.000 213.800 235.400 214.200 ;
        RECT 235.800 213.800 236.200 214.200 ;
        RECT 239.800 214.800 240.200 215.200 ;
        RECT 240.600 213.800 241.000 214.200 ;
        RECT 248.600 216.200 249.000 216.600 ;
        RECT 250.200 215.500 250.600 215.900 ;
        RECT 231.800 211.800 232.200 212.200 ;
        RECT 250.200 213.100 250.600 213.500 ;
        RECT 241.400 211.800 241.800 212.200 ;
        RECT 0.600 208.800 1.000 209.200 ;
        RECT 18.200 208.800 18.600 209.200 ;
        RECT 8.600 206.800 9.000 207.200 ;
        RECT 3.000 206.100 3.400 206.500 ;
        RECT 7.000 205.900 7.400 206.300 ;
        RECT 11.800 205.800 12.200 206.200 ;
        RECT 9.400 205.100 9.800 205.500 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 19.000 204.800 19.400 205.200 ;
        RECT 28.600 206.100 29.000 206.500 ;
        RECT 32.600 205.900 33.000 206.300 ;
        RECT 56.600 208.800 57.000 209.200 ;
        RECT 43.800 206.800 44.200 207.200 ;
        RECT 40.600 205.800 41.000 206.200 ;
        RECT 23.800 201.800 24.200 202.200 ;
        RECT 35.000 205.100 35.400 205.500 ;
        RECT 37.400 204.800 37.800 205.200 ;
        RECT 41.400 205.100 41.800 205.500 ;
        RECT 55.800 206.800 56.200 207.200 ;
        RECT 64.600 208.800 65.000 209.200 ;
        RECT 65.400 208.800 65.800 209.200 ;
        RECT 50.200 201.800 50.600 202.200 ;
        RECT 60.600 201.800 61.000 202.200 ;
        RECT 88.600 208.800 89.000 209.200 ;
        RECT 67.800 206.100 68.200 206.500 ;
        RECT 71.800 205.900 72.200 206.300 ;
        RECT 64.600 204.800 65.000 205.200 ;
        RECT 74.200 205.100 74.600 205.500 ;
        RECT 76.600 205.800 77.000 206.200 ;
        RECT 83.000 206.800 83.400 207.200 ;
        RECT 82.200 205.900 82.600 206.300 ;
        RECT 79.000 204.800 79.400 205.200 ;
        RECT 79.800 205.100 80.200 205.500 ;
        RECT 78.200 201.800 78.600 202.200 ;
        RECT 102.200 208.800 102.600 209.200 ;
        RECT 103.000 208.800 103.400 209.200 ;
        RECT 94.200 205.800 94.600 206.200 ;
        RECT 95.000 205.800 95.400 206.200 ;
        RECT 91.800 201.800 92.200 202.200 ;
        RECT 111.000 206.800 111.400 207.200 ;
        RECT 119.000 208.800 119.400 209.200 ;
        RECT 122.200 208.800 122.600 209.200 ;
        RECT 105.400 206.100 105.800 206.500 ;
        RECT 102.200 204.800 102.600 205.200 ;
        RECT 111.800 205.100 112.200 205.500 ;
        RECT 115.800 205.800 116.200 206.200 ;
        RECT 121.400 206.800 121.800 207.200 ;
        RECT 128.600 208.800 129.000 209.200 ;
        RECT 115.000 201.800 115.400 202.200 ;
        RECT 127.000 205.800 127.400 206.200 ;
        RECT 141.400 208.800 141.800 209.200 ;
        RECT 136.600 206.800 137.000 207.200 ;
        RECT 131.000 206.100 131.400 206.500 ;
        RECT 126.200 201.800 126.600 202.200 ;
        RECT 135.000 205.900 135.400 206.300 ;
        RECT 137.400 205.100 137.800 205.500 ;
        RECT 139.800 205.800 140.200 206.200 ;
        RECT 147.000 208.800 147.400 209.200 ;
        RECT 142.200 206.800 142.600 207.200 ;
        RECT 143.000 205.800 143.400 206.200 ;
        RECT 143.800 205.800 144.200 206.200 ;
        RECT 159.800 208.800 160.200 209.200 ;
        RECT 147.800 206.800 148.200 207.200 ;
        RECT 148.600 205.800 149.000 206.200 ;
        RECT 151.000 205.100 151.400 205.500 ;
        RECT 168.600 206.800 169.000 207.200 ;
        RECT 163.800 205.800 164.200 206.200 ;
        RECT 179.800 208.800 180.200 209.200 ;
        RECT 171.800 206.800 172.200 207.200 ;
        RECT 181.400 208.800 181.800 209.200 ;
        RECT 173.400 205.900 173.800 206.300 ;
        RECT 168.600 204.800 169.000 205.200 ;
        RECT 163.000 201.800 163.400 202.200 ;
        RECT 171.000 205.100 171.400 205.500 ;
        RECT 183.800 206.800 184.200 207.200 ;
        RECT 183.000 205.800 183.400 206.200 ;
        RECT 184.600 205.800 185.000 206.200 ;
        RECT 193.400 205.800 193.800 206.200 ;
        RECT 186.200 201.800 186.600 202.200 ;
        RECT 197.400 206.800 197.800 207.200 ;
        RECT 199.000 206.800 199.400 207.200 ;
        RECT 196.600 205.800 197.000 206.200 ;
        RECT 209.400 206.800 209.800 207.200 ;
        RECT 211.800 206.800 212.200 207.200 ;
        RECT 213.400 206.800 213.800 207.200 ;
        RECT 206.200 206.100 206.600 206.500 ;
        RECT 201.400 204.800 201.800 205.200 ;
        RECT 219.800 206.800 220.200 207.200 ;
        RECT 231.800 208.800 232.200 209.200 ;
        RECT 232.600 208.800 233.000 209.200 ;
        RECT 221.400 205.800 221.800 206.200 ;
        RECT 212.600 205.100 213.000 205.500 ;
        RECT 228.600 205.800 229.000 206.200 ;
        RECT 235.000 206.100 235.400 206.500 ;
        RECT 231.800 204.800 232.200 205.200 ;
        RECT 241.400 205.100 241.800 205.500 ;
        RECT 248.600 208.800 249.000 209.200 ;
        RECT 246.200 207.800 246.600 208.200 ;
        RECT 243.800 204.800 244.200 205.200 ;
        RECT 247.800 206.800 248.200 207.200 ;
        RECT 243.000 201.800 243.400 202.200 ;
        RECT 7.800 196.200 8.200 196.600 ;
        RECT 9.400 195.500 9.800 195.900 ;
        RECT 9.400 193.100 9.800 193.500 ;
        RECT 0.600 191.800 1.000 192.200 ;
        RECT 10.200 193.100 10.600 193.500 ;
        RECT 31.000 195.800 31.400 196.200 ;
        RECT 39.800 196.800 40.200 197.200 ;
        RECT 41.400 196.800 41.800 197.200 ;
        RECT 27.000 193.800 27.400 194.200 ;
        RECT 19.000 191.800 19.400 192.200 ;
        RECT 20.600 191.800 21.000 192.200 ;
        RECT 31.000 194.800 31.400 195.200 ;
        RECT 31.800 193.800 32.200 194.200 ;
        RECT 33.400 193.800 33.800 194.200 ;
        RECT 32.600 193.100 33.000 193.500 ;
        RECT 44.600 194.800 45.000 195.200 ;
        RECT 45.400 194.800 45.800 195.200 ;
        RECT 46.200 194.800 46.600 195.200 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 52.600 194.800 53.000 195.200 ;
        RECT 43.000 191.800 43.400 192.200 ;
        RECT 51.000 193.800 51.400 194.200 ;
        RECT 60.600 194.800 61.000 195.200 ;
        RECT 63.000 194.800 63.400 195.200 ;
        RECT 61.400 193.800 61.800 194.200 ;
        RECT 79.800 198.800 80.200 199.200 ;
        RECT 71.800 193.800 72.200 194.200 ;
        RECT 54.200 191.800 54.600 192.200 ;
        RECT 74.200 194.800 74.600 195.200 ;
        RECT 79.800 194.800 80.200 195.200 ;
        RECT 72.600 192.800 73.000 193.200 ;
        RECT 80.600 193.800 81.000 194.200 ;
        RECT 88.600 196.200 89.000 196.600 ;
        RECT 90.200 195.500 90.600 195.900 ;
        RECT 94.200 194.800 94.600 195.200 ;
        RECT 95.000 194.800 95.400 195.200 ;
        RECT 96.600 194.800 97.000 195.200 ;
        RECT 99.000 195.800 99.400 196.200 ;
        RECT 99.800 194.800 100.200 195.200 ;
        RECT 103.000 198.800 103.400 199.200 ;
        RECT 90.200 193.100 90.600 193.500 ;
        RECT 81.400 191.800 81.800 192.200 ;
        RECT 110.200 196.200 110.600 196.600 ;
        RECT 111.800 195.500 112.200 195.900 ;
        RECT 115.800 194.800 116.200 195.200 ;
        RECT 116.600 194.800 117.000 195.200 ;
        RECT 111.800 193.100 112.200 193.500 ;
        RECT 115.000 192.800 115.400 193.200 ;
        RECT 124.600 196.200 125.000 196.600 ;
        RECT 126.200 195.500 126.600 195.900 ;
        RECT 127.000 193.800 127.400 194.200 ;
        RECT 130.200 194.800 130.600 195.200 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 135.000 194.800 135.400 195.200 ;
        RECT 135.800 194.800 136.200 195.200 ;
        RECT 126.200 193.100 126.600 193.500 ;
        RECT 117.400 191.800 117.800 192.200 ;
        RECT 129.400 191.800 129.800 192.200 ;
        RECT 143.800 194.800 144.200 195.200 ;
        RECT 144.600 194.800 145.000 195.200 ;
        RECT 146.200 194.800 146.600 195.200 ;
        RECT 148.600 193.800 149.000 194.200 ;
        RECT 139.000 191.800 139.400 192.200 ;
        RECT 150.200 193.100 150.600 193.500 ;
        RECT 155.800 193.800 156.200 194.200 ;
        RECT 159.000 191.800 159.400 192.200 ;
        RECT 159.800 196.800 160.200 197.200 ;
        RECT 167.000 196.200 167.400 196.600 ;
        RECT 168.600 195.500 169.000 195.900 ;
        RECT 175.800 198.800 176.200 199.200 ;
        RECT 173.400 197.800 173.800 198.200 ;
        RECT 169.400 193.800 169.800 194.200 ;
        RECT 168.600 193.100 169.000 193.500 ;
        RECT 183.800 198.800 184.200 199.200 ;
        RECT 173.400 194.800 173.800 195.200 ;
        RECT 174.200 193.800 174.600 194.200 ;
        RECT 191.800 194.800 192.200 195.200 ;
        RECT 184.600 193.800 185.000 194.200 ;
        RECT 187.000 193.800 187.400 194.200 ;
        RECT 192.600 194.800 193.000 195.200 ;
        RECT 199.800 194.800 200.200 195.200 ;
        RECT 200.600 194.800 201.000 195.200 ;
        RECT 210.200 196.200 210.600 196.600 ;
        RECT 211.800 195.500 212.200 195.900 ;
        RECT 213.400 194.800 213.800 195.200 ;
        RECT 216.600 194.800 217.000 195.200 ;
        RECT 211.800 193.100 212.200 193.500 ;
        RECT 219.000 193.800 219.400 194.200 ;
        RECT 220.600 193.800 221.000 194.200 ;
        RECT 228.600 196.200 229.000 196.600 ;
        RECT 230.200 195.500 230.600 195.900 ;
        RECT 231.800 194.800 232.200 195.200 ;
        RECT 203.000 191.800 203.400 192.200 ;
        RECT 233.400 193.800 233.800 194.200 ;
        RECT 230.200 193.100 230.600 193.500 ;
        RECT 241.400 196.200 241.800 196.600 ;
        RECT 243.000 195.500 243.400 195.900 ;
        RECT 248.600 198.800 249.000 199.200 ;
        RECT 245.400 194.800 245.800 195.200 ;
        RECT 240.600 192.800 241.000 193.200 ;
        RECT 234.200 191.800 234.600 192.200 ;
        RECT 243.000 193.100 243.400 193.500 ;
        RECT 246.200 193.800 246.600 194.200 ;
        RECT 243.800 191.800 244.200 192.200 ;
        RECT 8.600 188.800 9.000 189.200 ;
        RECT 3.800 186.800 4.200 187.200 ;
        RECT 6.200 186.800 6.600 187.200 ;
        RECT 2.200 184.800 2.600 185.200 ;
        RECT 11.800 186.800 12.200 187.200 ;
        RECT 9.400 184.800 9.800 185.200 ;
        RECT 23.000 186.800 23.400 187.200 ;
        RECT 34.200 187.800 34.600 188.200 ;
        RECT 24.600 185.800 25.000 186.200 ;
        RECT 13.400 184.800 13.800 185.200 ;
        RECT 17.400 181.800 17.800 182.200 ;
        RECT 29.400 185.800 29.800 186.200 ;
        RECT 39.800 186.800 40.200 187.200 ;
        RECT 47.800 188.800 48.200 189.200 ;
        RECT 44.600 186.800 45.000 187.200 ;
        RECT 42.200 185.800 42.600 186.200 ;
        RECT 43.800 185.800 44.200 186.200 ;
        RECT 45.400 185.800 45.800 186.200 ;
        RECT 50.200 186.100 50.600 186.500 ;
        RECT 84.600 188.800 85.000 189.200 ;
        RECT 56.600 185.100 57.000 185.500 ;
        RECT 60.600 185.800 61.000 186.200 ;
        RECT 63.000 185.800 63.400 186.200 ;
        RECT 63.800 185.800 64.200 186.200 ;
        RECT 74.200 186.800 74.600 187.200 ;
        RECT 93.400 188.800 93.800 189.200 ;
        RECT 79.000 186.800 79.400 187.200 ;
        RECT 71.000 185.800 71.400 186.200 ;
        RECT 71.800 185.800 72.200 186.200 ;
        RECT 75.000 185.800 75.400 186.200 ;
        RECT 79.800 185.800 80.200 186.200 ;
        RECT 75.800 185.100 76.200 185.500 ;
        RECT 87.000 184.800 87.400 185.200 ;
        RECT 92.600 184.800 93.000 185.200 ;
        RECT 103.800 186.800 104.200 187.200 ;
        RECT 101.400 185.800 101.800 186.200 ;
        RECT 103.000 185.100 103.400 185.500 ;
        RECT 114.200 184.800 114.600 185.200 ;
        RECT 118.200 185.800 118.600 186.200 ;
        RECT 120.600 185.800 121.000 186.200 ;
        RECT 127.000 186.800 127.400 187.200 ;
        RECT 133.400 188.800 133.800 189.200 ;
        RECT 144.600 188.800 145.000 189.200 ;
        RECT 152.600 188.800 153.000 189.200 ;
        RECT 123.800 186.100 124.200 186.500 ;
        RECT 120.600 184.800 121.000 185.200 ;
        RECT 130.200 185.100 130.600 185.500 ;
        RECT 140.600 186.800 141.000 187.200 ;
        RECT 121.400 181.800 121.800 182.200 ;
        RECT 133.400 184.800 133.800 185.200 ;
        RECT 135.000 181.800 135.400 182.200 ;
        RECT 143.000 185.800 143.400 186.200 ;
        RECT 145.400 186.800 145.800 187.200 ;
        RECT 146.200 185.800 146.600 186.200 ;
        RECT 147.000 184.800 147.400 185.200 ;
        RECT 151.800 186.800 152.200 187.200 ;
        RECT 154.200 185.800 154.600 186.200 ;
        RECT 158.200 184.800 158.600 185.200 ;
        RECT 156.600 181.800 157.000 182.200 ;
        RECT 166.200 188.800 166.600 189.200 ;
        RECT 165.400 186.800 165.800 187.200 ;
        RECT 161.400 184.800 161.800 185.200 ;
        RECT 171.800 186.800 172.200 187.200 ;
        RECT 190.200 188.800 190.600 189.200 ;
        RECT 174.200 186.800 174.600 187.200 ;
        RECT 168.600 186.100 169.000 186.500 ;
        RECT 165.400 184.800 165.800 185.200 ;
        RECT 183.800 186.800 184.200 187.200 ;
        RECT 175.000 185.100 175.400 185.500 ;
        RECT 179.000 185.800 179.400 186.200 ;
        RECT 186.200 186.800 186.600 187.200 ;
        RECT 188.600 186.800 189.000 187.200 ;
        RECT 183.800 184.800 184.200 185.200 ;
        RECT 186.200 185.800 186.600 186.200 ;
        RECT 189.400 185.800 189.800 186.200 ;
        RECT 200.600 188.800 201.000 189.200 ;
        RECT 198.200 186.800 198.600 187.200 ;
        RECT 192.600 186.100 193.000 186.500 ;
        RECT 199.000 185.100 199.400 185.500 ;
        RECT 199.800 184.800 200.200 185.200 ;
        RECT 203.000 186.800 203.400 187.200 ;
        RECT 215.000 188.800 215.400 189.200 ;
        RECT 211.800 186.800 212.200 187.200 ;
        RECT 206.200 186.100 206.600 186.500 ;
        RECT 212.600 185.100 213.000 185.500 ;
        RECT 215.000 184.800 215.400 185.200 ;
        RECT 220.600 185.800 221.000 186.200 ;
        RECT 221.400 185.800 221.800 186.200 ;
        RECT 228.600 186.800 229.000 187.200 ;
        RECT 233.400 185.900 233.800 186.300 ;
        RECT 228.600 184.800 229.000 185.200 ;
        RECT 231.000 185.100 231.400 185.500 ;
        RECT 240.600 186.800 241.000 187.200 ;
        RECT 239.800 182.800 240.200 183.200 ;
        RECT 250.200 185.800 250.600 186.200 ;
        RECT 248.600 181.800 249.000 182.200 ;
        RECT 0.600 177.800 1.000 178.200 ;
        RECT 7.800 176.200 8.200 176.600 ;
        RECT 9.400 175.500 9.800 175.900 ;
        RECT 9.400 173.100 9.800 173.500 ;
        RECT 12.600 173.800 13.000 174.200 ;
        RECT 15.000 173.800 15.400 174.200 ;
        RECT 15.800 173.800 16.200 174.200 ;
        RECT 19.000 174.800 19.400 175.200 ;
        RECT 32.600 176.800 33.000 177.200 ;
        RECT 21.400 173.800 21.800 174.200 ;
        RECT 23.000 173.800 23.400 174.200 ;
        RECT 24.600 173.800 25.000 174.200 ;
        RECT 17.400 171.800 17.800 172.200 ;
        RECT 23.800 173.100 24.200 173.500 ;
        RECT 40.600 176.200 41.000 176.600 ;
        RECT 42.200 175.500 42.600 175.900 ;
        RECT 53.400 178.800 53.800 179.200 ;
        RECT 44.600 174.800 45.000 175.200 ;
        RECT 47.800 174.800 48.200 175.200 ;
        RECT 48.600 174.800 49.000 175.200 ;
        RECT 42.200 173.100 42.600 173.500 ;
        RECT 45.400 173.800 45.800 174.200 ;
        RECT 51.800 174.800 52.200 175.200 ;
        RECT 52.600 173.800 53.000 174.200 ;
        RECT 33.400 171.800 33.800 172.200 ;
        RECT 64.600 177.800 65.000 178.200 ;
        RECT 63.000 175.800 63.400 176.200 ;
        RECT 54.200 173.800 54.600 174.200 ;
        RECT 59.000 173.800 59.400 174.200 ;
        RECT 63.000 174.800 63.400 175.200 ;
        RECT 63.800 173.800 64.200 174.200 ;
        RECT 71.800 176.200 72.200 176.600 ;
        RECT 73.400 175.500 73.800 175.900 ;
        RECT 77.400 174.800 77.800 175.200 ;
        RECT 78.200 174.800 78.600 175.200 ;
        RECT 79.800 173.800 80.200 174.200 ;
        RECT 71.000 172.800 71.400 173.200 ;
        RECT 73.400 173.100 73.800 173.500 ;
        RECT 79.000 173.100 79.400 173.500 ;
        RECT 91.800 174.800 92.200 175.200 ;
        RECT 92.600 174.800 93.000 175.200 ;
        RECT 96.600 174.800 97.000 175.200 ;
        RECT 97.400 174.800 97.800 175.200 ;
        RECT 104.600 176.800 105.000 177.200 ;
        RECT 87.800 171.800 88.200 172.200 ;
        RECT 103.000 174.800 103.400 175.200 ;
        RECT 103.800 174.800 104.200 175.200 ;
        RECT 111.800 176.200 112.200 176.600 ;
        RECT 113.400 175.500 113.800 175.900 ;
        RECT 120.600 178.800 121.000 179.200 ;
        RECT 108.600 173.800 109.000 174.200 ;
        RECT 114.200 173.800 114.600 174.200 ;
        RECT 113.400 173.100 113.800 173.500 ;
        RECT 118.200 174.800 118.600 175.200 ;
        RECT 119.000 173.800 119.400 174.200 ;
        RECT 121.400 173.800 121.800 174.200 ;
        RECT 125.400 174.800 125.800 175.200 ;
        RECT 128.600 174.800 129.000 175.200 ;
        RECT 129.400 174.800 129.800 175.200 ;
        RECT 123.000 171.800 123.400 172.200 ;
        RECT 127.800 172.800 128.200 173.200 ;
        RECT 141.400 178.800 141.800 179.200 ;
        RECT 137.400 174.800 137.800 175.200 ;
        RECT 138.200 174.800 138.600 175.200 ;
        RECT 142.200 174.800 142.600 175.200 ;
        RECT 143.000 174.800 143.400 175.200 ;
        RECT 131.800 171.800 132.200 172.200 ;
        RECT 147.000 174.800 147.400 175.200 ;
        RECT 147.800 174.800 148.200 175.200 ;
        RECT 155.800 176.800 156.200 177.200 ;
        RECT 154.200 175.800 154.600 176.200 ;
        RECT 148.600 173.800 149.000 174.200 ;
        RECT 154.200 174.800 154.600 175.200 ;
        RECT 155.000 173.800 155.400 174.200 ;
        RECT 163.000 176.200 163.400 176.600 ;
        RECT 164.600 175.500 165.000 175.900 ;
        RECT 168.600 174.800 169.000 175.200 ;
        RECT 169.400 174.800 169.800 175.200 ;
        RECT 174.200 176.800 174.600 177.200 ;
        RECT 175.800 176.800 176.200 177.200 ;
        RECT 164.600 173.100 165.000 173.500 ;
        RECT 170.200 173.800 170.600 174.200 ;
        RECT 174.200 174.800 174.600 175.200 ;
        RECT 175.000 173.800 175.400 174.200 ;
        RECT 183.000 176.200 183.400 176.600 ;
        RECT 184.600 175.500 185.000 175.900 ;
        RECT 192.600 174.800 193.000 175.200 ;
        RECT 184.600 173.100 185.000 173.500 ;
        RECT 188.600 173.100 189.000 173.500 ;
        RECT 187.000 171.800 187.400 172.200 ;
        RECT 198.200 174.800 198.600 175.200 ;
        RECT 199.000 174.800 199.400 175.200 ;
        RECT 209.400 174.800 209.800 175.200 ;
        RECT 197.400 171.800 197.800 172.200 ;
        RECT 210.200 174.800 210.600 175.200 ;
        RECT 219.000 176.200 219.400 176.600 ;
        RECT 220.600 175.500 221.000 175.900 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 225.400 174.800 225.800 175.200 ;
        RECT 226.200 174.800 226.600 175.200 ;
        RECT 227.000 174.800 227.400 175.200 ;
        RECT 230.200 174.800 230.600 175.200 ;
        RECT 218.200 172.800 218.600 173.200 ;
        RECT 211.800 171.800 212.200 172.200 ;
        RECT 220.600 173.100 221.000 173.500 ;
        RECT 234.200 174.800 234.600 175.200 ;
        RECT 235.000 174.800 235.400 175.200 ;
        RECT 235.800 173.800 236.200 174.200 ;
        RECT 245.400 176.200 245.800 176.600 ;
        RECT 247.000 175.500 247.400 175.900 ;
        RECT 242.200 174.800 242.600 175.200 ;
        RECT 248.600 174.800 249.000 175.200 ;
        RECT 247.000 173.100 247.400 173.500 ;
        RECT 238.200 171.800 238.600 172.200 ;
        RECT 16.600 168.800 17.000 169.200 ;
        RECT 11.800 166.800 12.200 167.200 ;
        RECT 1.400 161.800 1.800 162.200 ;
        RECT 7.800 165.100 8.200 165.500 ;
        RECT 29.400 168.800 29.800 169.200 ;
        RECT 25.400 165.800 25.800 166.200 ;
        RECT 20.600 165.100 21.000 165.500 ;
        RECT 19.000 163.800 19.400 164.200 ;
        RECT 16.600 161.800 17.000 162.200 ;
        RECT 42.200 168.800 42.600 169.200 ;
        RECT 31.800 164.800 32.200 165.200 ;
        RECT 38.200 163.800 38.600 164.200 ;
        RECT 45.400 167.800 45.800 168.200 ;
        RECT 51.000 168.800 51.400 169.200 ;
        RECT 43.800 165.800 44.200 166.200 ;
        RECT 42.200 164.800 42.600 165.200 ;
        RECT 62.200 168.800 62.600 169.200 ;
        RECT 51.800 166.800 52.200 167.200 ;
        RECT 52.600 165.800 53.000 166.200 ;
        RECT 53.400 165.100 53.800 165.500 ;
        RECT 87.800 168.800 88.200 169.200 ;
        RECT 66.200 164.800 66.600 165.200 ;
        RECT 72.600 165.800 73.000 166.200 ;
        RECT 81.400 166.800 81.800 167.200 ;
        RECT 83.800 166.800 84.200 167.200 ;
        RECT 86.200 166.800 86.600 167.200 ;
        RECT 81.400 164.800 81.800 165.200 ;
        RECT 83.800 165.800 84.200 166.200 ;
        RECT 87.000 165.800 87.400 166.200 ;
        RECT 113.400 168.800 113.800 169.200 ;
        RECT 95.800 166.800 96.200 167.200 ;
        RECT 90.200 166.100 90.600 166.500 ;
        RECT 84.600 162.800 85.000 163.200 ;
        RECT 94.200 165.900 94.600 166.300 ;
        RECT 122.200 168.800 122.600 169.200 ;
        RECT 108.600 166.800 109.000 167.200 ;
        RECT 96.600 165.100 97.000 165.500 ;
        RECT 99.000 164.800 99.400 165.200 ;
        RECT 104.600 165.100 105.000 165.500 ;
        RECT 115.800 165.800 116.200 166.200 ;
        RECT 131.000 168.800 131.400 169.200 ;
        RECT 132.600 168.800 133.000 169.200 ;
        RECT 111.800 163.800 112.200 164.200 ;
        RECT 117.400 164.800 117.800 165.200 ;
        RECT 126.200 164.800 126.600 165.200 ;
        RECT 128.600 164.800 129.000 165.200 ;
        RECT 130.200 164.800 130.600 165.200 ;
        RECT 137.400 166.800 137.800 167.200 ;
        RECT 144.600 166.800 145.000 167.200 ;
        RECT 135.000 166.100 135.400 166.500 ;
        RECT 141.400 165.100 141.800 165.500 ;
        RECT 147.800 166.100 148.200 166.500 ;
        RECT 144.600 164.800 145.000 165.200 ;
        RECT 154.200 165.100 154.600 165.500 ;
        RECT 145.400 161.800 145.800 162.200 ;
        RECT 163.800 166.800 164.200 167.200 ;
        RECT 167.800 166.800 168.200 167.200 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 161.400 165.800 161.800 166.200 ;
        RECT 164.600 165.800 165.000 166.200 ;
        RECT 181.400 168.800 181.800 169.200 ;
        RECT 183.000 168.800 183.400 169.200 ;
        RECT 175.000 166.800 175.400 167.200 ;
        RECT 162.200 163.800 162.600 164.200 ;
        RECT 168.600 164.800 169.000 165.200 ;
        RECT 174.200 165.800 174.600 166.200 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 180.600 164.800 181.000 165.200 ;
        RECT 195.000 168.800 195.400 169.200 ;
        RECT 200.600 168.800 201.000 169.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 185.400 166.100 185.800 166.500 ;
        RECT 191.800 165.100 192.200 165.500 ;
        RECT 211.000 168.800 211.400 169.200 ;
        RECT 195.800 164.800 196.200 165.200 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 211.000 164.800 211.400 165.200 ;
        RECT 213.400 164.800 213.800 165.200 ;
        RECT 234.200 168.800 234.600 169.200 ;
        RECT 225.400 166.800 225.800 167.200 ;
        RECT 219.800 166.100 220.200 166.500 ;
        RECT 233.400 166.800 233.800 167.200 ;
        RECT 226.200 165.100 226.600 165.500 ;
        RECT 217.400 163.800 217.800 164.200 ;
        RECT 227.800 161.800 228.200 162.200 ;
        RECT 242.200 166.800 242.600 167.200 ;
        RECT 236.600 166.100 237.000 166.500 ;
        RECT 240.600 165.900 241.000 166.300 ;
        RECT 243.000 165.100 243.400 165.500 ;
        RECT 246.200 165.800 246.600 166.200 ;
        RECT 244.600 161.800 245.000 162.200 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 4.600 154.800 5.000 155.200 ;
        RECT 1.400 153.800 1.800 154.200 ;
        RECT 0.600 153.100 1.000 153.500 ;
        RECT 10.200 153.800 10.600 154.200 ;
        RECT 14.200 154.800 14.600 155.200 ;
        RECT 15.000 153.800 15.400 154.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 19.800 154.800 20.200 155.200 ;
        RECT 21.400 154.800 21.800 155.200 ;
        RECT 18.200 151.800 18.600 152.200 ;
        RECT 23.000 152.800 23.400 153.200 ;
        RECT 26.200 156.800 26.600 157.200 ;
        RECT 25.400 153.800 25.800 154.200 ;
        RECT 33.400 156.200 33.800 156.600 ;
        RECT 36.600 158.800 37.000 159.200 ;
        RECT 39.000 158.800 39.400 159.200 ;
        RECT 35.000 155.500 35.400 155.900 ;
        RECT 35.000 153.100 35.400 153.500 ;
        RECT 44.600 158.800 45.000 159.200 ;
        RECT 51.800 158.800 52.200 159.200 ;
        RECT 53.400 156.800 53.800 157.200 ;
        RECT 45.400 154.800 45.800 155.200 ;
        RECT 46.200 154.800 46.600 155.200 ;
        RECT 36.600 151.800 37.000 152.200 ;
        RECT 39.000 151.800 39.400 152.200 ;
        RECT 40.600 151.800 41.000 152.200 ;
        RECT 51.000 153.800 51.400 154.200 ;
        RECT 48.600 152.800 49.000 153.200 ;
        RECT 60.600 156.200 61.000 156.600 ;
        RECT 62.200 155.500 62.600 155.900 ;
        RECT 74.200 158.800 74.600 159.200 ;
        RECT 81.400 156.800 81.800 157.200 ;
        RECT 55.000 153.800 55.400 154.200 ;
        RECT 63.000 153.800 63.400 154.200 ;
        RECT 62.200 153.100 62.600 153.500 ;
        RECT 67.000 154.800 67.400 155.200 ;
        RECT 67.800 153.800 68.200 154.200 ;
        RECT 76.600 154.800 77.000 155.200 ;
        RECT 78.200 154.800 78.600 155.200 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 88.600 156.200 89.000 156.600 ;
        RECT 112.600 158.800 113.000 159.200 ;
        RECT 90.200 155.500 90.600 155.900 ;
        RECT 91.000 154.800 91.400 155.200 ;
        RECT 90.200 153.100 90.600 153.500 ;
        RECT 95.000 151.800 95.400 152.200 ;
        RECT 99.800 152.800 100.200 153.200 ;
        RECT 102.200 151.800 102.600 152.200 ;
        RECT 105.400 152.800 105.800 153.200 ;
        RECT 107.800 151.800 108.200 152.200 ;
        RECT 111.000 152.800 111.400 153.200 ;
        RECT 123.800 156.800 124.200 157.200 ;
        RECT 117.400 154.800 117.800 155.200 ;
        RECT 115.000 153.800 115.400 154.200 ;
        RECT 114.200 153.100 114.600 153.500 ;
        RECT 123.800 153.800 124.200 154.200 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 129.400 154.800 129.800 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 128.600 153.800 129.000 154.200 ;
        RECT 143.000 156.800 143.400 157.200 ;
        RECT 144.600 158.800 145.000 159.200 ;
        RECT 138.200 154.800 138.600 155.200 ;
        RECT 134.200 153.100 134.600 153.500 ;
        RECT 145.400 153.800 145.800 154.200 ;
        RECT 146.200 153.800 146.600 154.200 ;
        RECT 152.600 158.800 153.000 159.200 ;
        RECT 153.400 154.800 153.800 155.200 ;
        RECT 154.200 154.800 154.600 155.200 ;
        RECT 155.800 154.800 156.200 155.200 ;
        RECT 158.200 153.800 158.600 154.200 ;
        RECT 147.800 151.800 148.200 152.200 ;
        RECT 159.800 153.800 160.200 154.200 ;
        RECT 167.800 156.200 168.200 156.600 ;
        RECT 169.400 155.500 169.800 155.900 ;
        RECT 170.200 153.800 170.600 154.200 ;
        RECT 169.400 153.100 169.800 153.500 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 183.000 156.800 183.400 157.200 ;
        RECT 175.000 153.800 175.400 154.200 ;
        RECT 178.200 154.800 178.600 155.200 ;
        RECT 179.000 154.800 179.400 155.200 ;
        RECT 177.400 153.800 177.800 154.200 ;
        RECT 182.200 154.800 182.600 155.200 ;
        RECT 171.800 151.800 172.200 152.200 ;
        RECT 190.200 156.200 190.600 156.600 ;
        RECT 191.800 155.500 192.200 155.900 ;
        RECT 192.600 153.800 193.000 154.200 ;
        RECT 191.800 153.100 192.200 153.500 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 199.000 154.800 199.400 155.200 ;
        RECT 201.400 155.800 201.800 156.200 ;
        RECT 202.200 154.800 202.600 155.200 ;
        RECT 198.200 153.800 198.600 154.200 ;
        RECT 205.400 156.800 205.800 157.200 ;
        RECT 204.600 153.800 205.000 154.200 ;
        RECT 212.600 156.200 213.000 156.600 ;
        RECT 214.200 155.500 214.600 155.900 ;
        RECT 215.000 158.800 215.400 159.200 ;
        RECT 222.200 156.200 222.600 156.600 ;
        RECT 223.800 155.500 224.200 155.900 ;
        RECT 214.200 153.100 214.600 153.500 ;
        RECT 232.600 154.800 233.000 155.200 ;
        RECT 223.800 153.100 224.200 153.500 ;
        RECT 235.000 153.800 235.400 154.200 ;
        RECT 236.600 153.800 237.000 154.200 ;
        RECT 244.600 156.200 245.000 156.600 ;
        RECT 246.200 155.500 246.600 155.900 ;
        RECT 230.200 151.800 230.600 152.200 ;
        RECT 246.200 153.100 246.600 153.500 ;
        RECT 247.000 152.800 247.400 153.200 ;
        RECT 251.800 155.800 252.200 156.200 ;
        RECT 247.800 151.800 248.200 152.200 ;
        RECT 1.400 146.800 1.800 147.200 ;
        RECT 0.600 145.100 1.000 145.500 ;
        RECT 16.600 146.800 17.000 147.200 ;
        RECT 10.200 143.800 10.600 144.200 ;
        RECT 11.800 144.800 12.200 145.200 ;
        RECT 19.800 145.800 20.200 146.200 ;
        RECT 15.800 145.100 16.200 145.500 ;
        RECT 27.000 145.800 27.400 146.200 ;
        RECT 24.600 141.800 25.000 142.200 ;
        RECT 28.600 144.800 29.000 145.200 ;
        RECT 37.400 145.800 37.800 146.200 ;
        RECT 39.800 145.800 40.200 146.200 ;
        RECT 45.400 146.800 45.800 147.200 ;
        RECT 41.400 141.800 41.800 142.200 ;
        RECT 47.000 145.800 47.400 146.200 ;
        RECT 47.800 144.800 48.200 145.200 ;
        RECT 56.600 145.800 57.000 146.200 ;
        RECT 79.800 148.800 80.200 149.200 ;
        RECT 68.600 146.800 69.000 147.200 ;
        RECT 51.800 141.800 52.200 142.200 ;
        RECT 53.400 141.800 53.800 142.200 ;
        RECT 63.000 141.800 63.400 142.200 ;
        RECT 64.600 145.100 65.000 145.500 ;
        RECT 75.800 146.800 76.200 147.200 ;
        RECT 75.000 145.800 75.400 146.200 ;
        RECT 73.400 141.800 73.800 142.200 ;
        RECT 77.400 144.800 77.800 145.200 ;
        RECT 107.000 148.800 107.400 149.200 ;
        RECT 86.200 146.800 86.600 147.200 ;
        RECT 89.400 146.800 89.800 147.200 ;
        RECT 82.200 146.100 82.600 146.500 ;
        RECT 99.000 146.800 99.400 147.200 ;
        RECT 116.600 148.800 117.000 149.200 ;
        RECT 100.600 145.900 101.000 146.300 ;
        RECT 88.600 145.100 89.000 145.500 ;
        RECT 98.200 145.100 98.600 145.500 ;
        RECT 108.600 146.800 109.000 147.200 ;
        RECT 110.200 145.900 110.600 146.300 ;
        RECT 107.800 145.100 108.200 145.500 ;
        RECT 131.000 148.800 131.400 149.200 ;
        RECT 123.000 146.800 123.400 147.200 ;
        RECT 121.400 145.800 121.800 146.200 ;
        RECT 124.600 145.900 125.000 146.300 ;
        RECT 122.200 145.100 122.600 145.500 ;
        RECT 136.600 148.800 137.000 149.200 ;
        RECT 132.600 145.800 133.000 146.200 ;
        RECT 153.400 148.800 153.800 149.200 ;
        RECT 139.000 146.100 139.400 146.500 ;
        RECT 143.000 145.900 143.400 146.300 ;
        RECT 145.400 145.100 145.800 145.500 ;
        RECT 159.800 146.800 160.200 147.200 ;
        RECT 151.000 144.800 151.400 145.200 ;
        RECT 171.000 148.800 171.400 149.200 ;
        RECT 163.000 146.800 163.400 147.200 ;
        RECT 175.000 148.800 175.400 149.200 ;
        RECT 164.600 145.900 165.000 146.300 ;
        RECT 159.800 144.800 160.200 145.200 ;
        RECT 162.200 145.100 162.600 145.500 ;
        RECT 179.000 146.800 179.400 147.200 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 177.400 146.100 177.800 146.500 ;
        RECT 199.800 146.800 200.200 147.200 ;
        RECT 183.800 145.100 184.200 145.500 ;
        RECT 185.400 141.800 185.800 142.200 ;
        RECT 195.000 145.800 195.400 146.200 ;
        RECT 208.600 148.800 209.000 149.200 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 199.800 144.800 200.200 145.200 ;
        RECT 207.000 145.800 207.400 146.200 ;
        RECT 228.600 148.800 229.000 149.200 ;
        RECT 216.600 146.800 217.000 147.200 ;
        RECT 211.000 146.100 211.400 146.500 ;
        RECT 219.000 145.800 219.400 146.200 ;
        RECT 217.400 145.100 217.800 145.500 ;
        RECT 227.800 145.800 228.200 146.200 ;
        RECT 250.200 148.800 250.600 149.200 ;
        RECT 240.600 146.800 241.000 147.200 ;
        RECT 243.800 146.800 244.200 147.200 ;
        RECT 231.000 146.100 231.400 146.500 ;
        RECT 224.600 144.800 225.000 145.200 ;
        RECT 227.000 144.800 227.400 145.200 ;
        RECT 237.400 145.100 237.800 145.500 ;
        RECT 240.600 144.800 241.000 145.200 ;
        RECT 241.400 145.100 241.800 145.500 ;
        RECT 3.000 138.800 3.400 139.200 ;
        RECT 7.800 134.800 8.200 135.200 ;
        RECT 5.400 133.800 5.800 134.200 ;
        RECT 4.600 133.100 5.000 133.500 ;
        RECT 15.000 134.800 15.400 135.200 ;
        RECT 15.800 134.800 16.200 135.200 ;
        RECT 19.000 133.800 19.400 134.200 ;
        RECT 24.600 136.800 25.000 137.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 21.400 133.800 21.800 134.200 ;
        RECT 13.400 131.800 13.800 132.200 ;
        RECT 35.800 138.800 36.200 139.200 ;
        RECT 39.800 138.800 40.200 139.200 ;
        RECT 29.400 133.800 29.800 134.200 ;
        RECT 44.600 138.800 45.000 139.200 ;
        RECT 40.600 134.800 41.000 135.200 ;
        RECT 41.400 134.800 41.800 135.200 ;
        RECT 47.800 134.800 48.200 135.200 ;
        RECT 48.600 134.800 49.000 135.200 ;
        RECT 51.800 133.800 52.200 134.200 ;
        RECT 59.800 136.200 60.200 136.600 ;
        RECT 61.400 135.500 61.800 135.900 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 61.400 133.100 61.800 133.500 ;
        RECT 69.400 134.800 69.800 135.200 ;
        RECT 52.600 131.800 53.000 132.200 ;
        RECT 64.600 132.800 65.000 133.200 ;
        RECT 75.000 134.800 75.400 135.200 ;
        RECT 75.800 134.800 76.200 135.200 ;
        RECT 83.800 138.800 84.200 139.200 ;
        RECT 83.800 134.800 84.200 135.200 ;
        RECT 86.200 134.800 86.600 135.200 ;
        RECT 84.600 133.800 85.000 134.200 ;
        RECT 88.600 133.800 89.000 134.200 ;
        RECT 111.800 136.800 112.200 137.200 ;
        RECT 90.200 133.800 90.600 134.200 ;
        RECT 91.000 133.100 91.400 133.500 ;
        RECT 105.400 134.800 105.800 135.200 ;
        RECT 99.800 131.800 100.200 132.200 ;
        RECT 102.200 133.100 102.600 133.500 ;
        RECT 111.800 133.800 112.200 134.200 ;
        RECT 115.800 134.800 116.200 135.200 ;
        RECT 116.600 133.800 117.000 134.200 ;
        RECT 120.600 134.800 121.000 135.200 ;
        RECT 121.400 134.800 121.800 135.200 ;
        RECT 122.200 133.800 122.600 134.200 ;
        RECT 126.200 134.800 126.600 135.200 ;
        RECT 127.000 133.800 127.400 134.200 ;
        RECT 135.000 136.200 135.400 136.600 ;
        RECT 136.600 135.500 137.000 135.900 ;
        RECT 147.000 136.800 147.400 137.200 ;
        RECT 142.200 134.800 142.600 135.200 ;
        RECT 124.600 131.800 125.000 132.200 ;
        RECT 138.200 133.800 138.600 134.200 ;
        RECT 134.200 132.800 134.600 133.200 ;
        RECT 127.800 131.800 128.200 132.200 ;
        RECT 136.600 133.100 137.000 133.500 ;
        RECT 137.400 133.100 137.800 133.500 ;
        RECT 147.000 133.800 147.400 134.200 ;
        RECT 164.600 136.800 165.000 137.200 ;
        RECT 154.200 134.800 154.600 135.200 ;
        RECT 155.000 134.800 155.400 135.200 ;
        RECT 159.000 134.800 159.400 135.200 ;
        RECT 156.600 133.800 157.000 134.200 ;
        RECT 153.400 131.800 153.800 132.200 ;
        RECT 155.800 133.100 156.200 133.500 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 174.200 134.800 174.600 135.200 ;
        RECT 175.800 134.800 176.200 135.200 ;
        RECT 176.600 134.800 177.000 135.200 ;
        RECT 175.000 133.800 175.400 134.200 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 193.400 134.800 193.800 135.200 ;
        RECT 194.200 134.800 194.600 135.200 ;
        RECT 195.800 134.800 196.200 135.200 ;
        RECT 198.200 133.800 198.600 134.200 ;
        RECT 201.400 133.800 201.800 134.200 ;
        RECT 209.400 136.200 209.800 136.600 ;
        RECT 211.000 135.500 211.400 135.900 ;
        RECT 217.400 136.800 217.800 137.200 ;
        RECT 211.800 133.800 212.200 134.200 ;
        RECT 211.000 133.100 211.400 133.500 ;
        RECT 215.800 134.800 216.200 135.200 ;
        RECT 216.600 133.800 217.000 134.200 ;
        RECT 224.600 136.200 225.000 136.600 ;
        RECT 226.200 135.500 226.600 135.900 ;
        RECT 234.200 136.200 234.600 136.600 ;
        RECT 235.800 135.500 236.200 135.900 ;
        RECT 240.600 138.800 241.000 139.200 ;
        RECT 243.800 138.800 244.200 139.200 ;
        RECT 238.200 134.800 238.600 135.200 ;
        RECT 226.200 133.100 226.600 133.500 ;
        RECT 235.800 133.100 236.200 133.500 ;
        RECT 242.200 134.800 242.600 135.200 ;
        RECT 227.000 131.800 227.400 132.200 ;
        RECT 243.800 131.800 244.200 132.200 ;
        RECT 9.400 128.800 9.800 129.200 ;
        RECT 1.400 126.800 1.800 127.200 ;
        RECT 27.800 128.800 28.200 129.200 ;
        RECT 5.400 125.800 5.800 126.200 ;
        RECT 0.600 125.100 1.000 125.500 ;
        RECT 10.200 124.800 10.600 125.200 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 21.400 126.800 21.800 127.200 ;
        RECT 18.200 124.800 18.600 125.200 ;
        RECT 19.000 125.100 19.400 125.500 ;
        RECT 30.200 125.800 30.600 126.200 ;
        RECT 37.400 126.800 37.800 127.200 ;
        RECT 36.600 125.800 37.000 126.200 ;
        RECT 43.000 126.800 43.400 127.200 ;
        RECT 42.200 125.800 42.600 126.200 ;
        RECT 43.000 125.800 43.400 126.200 ;
        RECT 47.000 126.800 47.400 127.200 ;
        RECT 46.200 125.800 46.600 126.200 ;
        RECT 49.400 125.800 49.800 126.200 ;
        RECT 62.200 128.800 62.600 129.200 ;
        RECT 58.200 126.800 58.600 127.200 ;
        RECT 52.600 126.100 53.000 126.500 ;
        RECT 59.000 125.100 59.400 125.500 ;
        RECT 61.400 124.800 61.800 125.200 ;
        RECT 74.200 128.800 74.600 129.200 ;
        RECT 78.200 127.800 78.600 128.200 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 68.600 126.800 69.000 127.200 ;
        RECT 76.600 125.800 77.000 126.200 ;
        RECT 81.400 126.800 81.800 127.200 ;
        RECT 83.800 125.800 84.200 126.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 83.000 124.800 83.400 125.200 ;
        RECT 84.600 124.800 85.000 125.200 ;
        RECT 88.600 128.800 89.000 129.200 ;
        RECT 100.600 126.800 101.000 127.200 ;
        RECT 88.600 121.800 89.000 122.200 ;
        RECT 103.800 126.800 104.200 127.200 ;
        RECT 98.200 125.800 98.600 126.200 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 118.200 126.800 118.600 127.200 ;
        RECT 129.400 128.800 129.800 129.200 ;
        RECT 118.200 124.800 118.600 125.200 ;
        RECT 120.600 125.100 121.000 125.500 ;
        RECT 134.200 126.800 134.600 127.200 ;
        RECT 150.200 128.800 150.600 129.200 ;
        RECT 138.200 126.800 138.600 127.200 ;
        RECT 132.600 126.100 133.000 126.500 ;
        RECT 136.600 125.900 137.000 126.300 ;
        RECT 145.400 126.800 145.800 127.200 ;
        RECT 147.000 126.800 147.400 127.200 ;
        RECT 139.000 125.100 139.400 125.500 ;
        RECT 130.200 121.800 130.600 122.200 ;
        RECT 141.400 124.800 141.800 125.200 ;
        RECT 154.200 126.800 154.600 127.200 ;
        RECT 158.200 126.800 158.600 127.200 ;
        RECT 152.600 126.100 153.000 126.500 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 156.600 125.900 157.000 126.300 ;
        RECT 159.000 125.100 159.400 125.500 ;
        RECT 161.400 124.800 161.800 125.200 ;
        RECT 172.600 126.800 173.000 127.200 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 184.600 128.800 185.000 129.200 ;
        RECT 178.200 125.900 178.600 126.300 ;
        RECT 173.400 124.800 173.800 125.200 ;
        RECT 175.800 125.100 176.200 125.500 ;
        RECT 192.600 126.800 193.000 127.200 ;
        RECT 200.600 128.800 201.000 129.200 ;
        RECT 188.600 125.800 189.000 126.200 ;
        RECT 190.200 125.800 190.600 126.200 ;
        RECT 195.000 125.800 195.400 126.200 ;
        RECT 208.600 126.800 209.000 127.200 ;
        RECT 203.000 126.100 203.400 126.500 ;
        RECT 207.000 125.900 207.400 126.300 ;
        RECT 209.400 125.100 209.800 125.500 ;
        RECT 211.800 124.800 212.200 125.200 ;
        RECT 219.000 125.800 219.400 126.200 ;
        RECT 220.600 124.800 221.000 125.200 ;
        RECT 241.400 128.800 241.800 129.200 ;
        RECT 234.200 126.800 234.600 127.200 ;
        RECT 228.600 126.100 229.000 126.500 ;
        RECT 224.600 124.800 225.000 125.200 ;
        RECT 235.000 125.100 235.400 125.500 ;
        RECT 226.200 123.800 226.600 124.200 ;
        RECT 239.000 126.800 239.400 127.200 ;
        RECT 237.400 124.800 237.800 125.200 ;
        RECT 245.400 126.800 245.800 127.200 ;
        RECT 249.400 126.800 249.800 127.200 ;
        RECT 243.800 126.100 244.200 126.500 ;
        RECT 250.200 125.100 250.600 125.500 ;
        RECT 241.400 121.800 241.800 122.200 ;
        RECT 1.400 118.800 1.800 119.200 ;
        RECT 22.200 116.800 22.600 117.200 ;
        RECT 7.800 113.800 8.200 114.200 ;
        RECT 1.400 111.800 1.800 112.200 ;
        RECT 12.600 114.800 13.000 115.200 ;
        RECT 25.400 118.800 25.800 119.200 ;
        RECT 12.600 113.800 13.000 114.200 ;
        RECT 13.400 113.100 13.800 113.500 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 23.800 114.800 24.200 115.200 ;
        RECT 27.800 113.800 28.200 114.200 ;
        RECT 37.400 114.800 37.800 115.200 ;
        RECT 47.800 116.800 48.200 117.200 ;
        RECT 34.200 113.800 34.600 114.200 ;
        RECT 33.400 113.100 33.800 113.500 ;
        RECT 32.600 111.800 33.000 112.200 ;
        RECT 39.000 113.800 39.400 114.200 ;
        RECT 44.600 114.800 45.000 115.200 ;
        RECT 46.200 113.800 46.600 114.200 ;
        RECT 55.000 116.200 55.400 116.600 ;
        RECT 56.600 115.500 57.000 115.900 ;
        RECT 58.200 114.800 58.600 115.200 ;
        RECT 64.600 115.800 65.000 116.200 ;
        RECT 42.200 111.800 42.600 112.200 ;
        RECT 56.600 113.100 57.000 113.500 ;
        RECT 70.200 118.800 70.600 119.200 ;
        RECT 66.200 114.800 66.600 115.200 ;
        RECT 67.000 114.800 67.400 115.200 ;
        RECT 67.800 114.800 68.200 115.200 ;
        RECT 68.600 114.800 69.000 115.200 ;
        RECT 72.600 113.800 73.000 114.200 ;
        RECT 77.400 118.800 77.800 119.200 ;
        RECT 78.200 114.800 78.600 115.200 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 94.200 116.800 94.600 117.200 ;
        RECT 74.200 111.800 74.600 112.200 ;
        RECT 88.600 114.800 89.000 115.200 ;
        RECT 84.600 113.800 85.000 114.200 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 85.400 113.100 85.800 113.500 ;
        RECT 95.000 113.800 95.400 114.200 ;
        RECT 87.800 112.800 88.200 113.200 ;
        RECT 97.400 115.800 97.800 116.200 ;
        RECT 103.000 114.800 103.400 115.200 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 110.200 118.800 110.600 119.200 ;
        RECT 104.600 113.800 105.000 114.200 ;
        RECT 108.600 114.800 109.000 115.200 ;
        RECT 109.400 113.800 109.800 114.200 ;
        RECT 117.400 116.200 117.800 116.600 ;
        RECT 119.000 115.500 119.400 115.900 ;
        RECT 96.600 111.800 97.000 112.200 ;
        RECT 127.000 116.200 127.400 116.600 ;
        RECT 128.600 115.500 129.000 115.900 ;
        RECT 135.000 118.800 135.400 119.200 ;
        RECT 119.000 113.100 119.400 113.500 ;
        RECT 129.400 113.800 129.800 114.200 ;
        RECT 136.600 114.800 137.000 115.200 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 128.600 113.100 129.000 113.500 ;
        RECT 119.800 111.800 120.200 112.200 ;
        RECT 140.600 113.800 141.000 114.200 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 147.000 113.800 147.400 114.200 ;
        RECT 155.800 116.200 156.200 116.600 ;
        RECT 157.400 115.500 157.800 115.900 ;
        RECT 159.800 114.800 160.200 115.200 ;
        RECT 164.600 114.800 165.000 115.200 ;
        RECT 143.800 111.800 144.200 112.200 ;
        RECT 157.400 113.100 157.800 113.500 ;
        RECT 160.600 113.800 161.000 114.200 ;
        RECT 162.200 113.800 162.600 114.200 ;
        RECT 161.400 113.100 161.800 113.500 ;
        RECT 148.600 111.800 149.000 112.200 ;
        RECT 158.200 111.800 158.600 112.200 ;
        RECT 171.800 114.800 172.200 115.200 ;
        RECT 176.600 114.800 177.000 115.200 ;
        RECT 177.400 114.800 177.800 115.200 ;
        RECT 175.800 113.800 176.200 114.200 ;
        RECT 181.400 114.800 181.800 115.200 ;
        RECT 182.200 113.800 182.600 114.200 ;
        RECT 170.200 111.800 170.600 112.200 ;
        RECT 183.800 114.800 184.200 115.200 ;
        RECT 184.600 113.800 185.000 114.200 ;
        RECT 191.000 114.800 191.400 115.200 ;
        RECT 193.400 114.800 193.800 115.200 ;
        RECT 188.600 113.800 189.000 114.200 ;
        RECT 191.800 113.800 192.200 114.200 ;
        RECT 195.000 113.800 195.400 114.200 ;
        RECT 207.000 116.200 207.400 116.600 ;
        RECT 208.600 115.500 209.000 115.900 ;
        RECT 212.600 114.800 213.000 115.200 ;
        RECT 210.200 113.800 210.600 114.200 ;
        RECT 186.200 111.800 186.600 112.200 ;
        RECT 189.400 111.800 189.800 112.200 ;
        RECT 208.600 113.100 209.000 113.500 ;
        RECT 199.800 111.800 200.200 112.200 ;
        RECT 209.400 113.100 209.800 113.500 ;
        RECT 215.000 113.800 215.400 114.200 ;
        RECT 219.800 114.800 220.200 115.200 ;
        RECT 224.600 114.800 225.000 115.200 ;
        RECT 225.400 114.800 225.800 115.200 ;
        RECT 226.200 114.800 226.600 115.200 ;
        RECT 230.200 114.800 230.600 115.200 ;
        RECT 231.000 114.800 231.400 115.200 ;
        RECT 218.200 111.800 218.600 112.200 ;
        RECT 239.000 117.800 239.400 118.200 ;
        RECT 238.200 113.800 238.600 114.200 ;
        RECT 249.400 117.800 249.800 118.200 ;
        RECT 241.400 113.800 241.800 114.200 ;
        RECT 240.600 113.100 241.000 113.500 ;
        RECT 236.600 111.800 237.000 112.200 ;
        RECT 1.400 106.800 1.800 107.200 ;
        RECT 11.000 108.800 11.400 109.200 ;
        RECT 13.400 108.800 13.800 109.200 ;
        RECT 3.000 105.900 3.400 106.300 ;
        RECT 0.600 105.100 1.000 105.500 ;
        RECT 10.200 106.800 10.600 107.200 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 18.200 106.800 18.600 107.200 ;
        RECT 28.600 108.800 29.000 109.200 ;
        RECT 15.800 106.100 16.200 106.500 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 11.000 101.800 11.400 102.200 ;
        RECT 19.800 105.900 20.200 106.300 ;
        RECT 22.200 105.100 22.600 105.500 ;
        RECT 13.400 101.800 13.800 102.200 ;
        RECT 24.600 104.800 25.000 105.200 ;
        RECT 34.200 106.800 34.600 107.200 ;
        RECT 39.000 108.800 39.400 109.200 ;
        RECT 31.000 106.100 31.400 106.500 ;
        RECT 37.400 105.100 37.800 105.500 ;
        RECT 45.400 104.800 45.800 105.200 ;
        RECT 47.800 106.800 48.200 107.200 ;
        RECT 59.000 106.800 59.400 107.200 ;
        RECT 75.000 108.800 75.400 109.200 ;
        RECT 56.600 106.100 57.000 106.500 ;
        RECT 60.600 105.900 61.000 106.300 ;
        RECT 63.000 105.100 63.400 105.500 ;
        RECT 63.800 104.800 64.200 105.200 ;
        RECT 69.400 106.800 69.800 107.200 ;
        RECT 72.600 106.800 73.000 107.200 ;
        RECT 93.400 108.800 93.800 109.200 ;
        RECT 107.800 108.800 108.200 109.200 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 77.400 106.100 77.800 106.500 ;
        RECT 87.000 105.900 87.400 106.300 ;
        RECT 83.800 105.100 84.200 105.500 ;
        RECT 84.600 105.100 85.000 105.500 ;
        RECT 96.600 104.800 97.000 105.200 ;
        RECT 97.400 104.800 97.800 105.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 98.200 101.800 98.600 102.200 ;
        RECT 103.800 106.800 104.200 107.200 ;
        RECT 103.800 104.800 104.200 105.200 ;
        RECT 119.000 108.800 119.400 109.200 ;
        RECT 125.400 108.800 125.800 109.200 ;
        RECT 109.400 101.800 109.800 102.200 ;
        RECT 112.600 104.800 113.000 105.200 ;
        RECT 123.000 104.800 123.400 105.200 ;
        RECT 121.400 101.800 121.800 102.200 ;
        RECT 124.600 104.800 125.000 105.200 ;
        RECT 130.200 104.800 130.600 105.200 ;
        RECT 131.000 104.800 131.400 105.200 ;
        RECT 129.400 101.800 129.800 102.200 ;
        RECT 135.800 108.800 136.200 109.200 ;
        RECT 133.400 106.800 133.800 107.200 ;
        RECT 138.200 106.100 138.600 106.500 ;
        RECT 135.000 104.800 135.400 105.200 ;
        RECT 131.800 101.800 132.200 102.200 ;
        RECT 142.200 105.900 142.600 106.300 ;
        RECT 144.600 105.100 145.000 105.500 ;
        RECT 155.800 104.800 156.200 105.200 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 159.800 105.800 160.200 106.200 ;
        RECT 161.400 105.800 161.800 106.200 ;
        RECT 164.600 105.800 165.000 106.200 ;
        RECT 171.000 106.800 171.400 107.200 ;
        RECT 162.200 103.800 162.600 104.200 ;
        RECT 165.400 104.800 165.800 105.200 ;
        RECT 172.600 106.800 173.000 107.200 ;
        RECT 170.200 104.800 170.600 105.200 ;
        RECT 171.000 102.800 171.400 103.200 ;
        RECT 182.200 106.800 182.600 107.200 ;
        RECT 189.400 108.800 189.800 109.200 ;
        RECT 179.000 106.100 179.400 106.500 ;
        RECT 185.400 105.100 185.800 105.500 ;
        RECT 197.400 106.800 197.800 107.200 ;
        RECT 191.800 106.100 192.200 106.500 ;
        RECT 187.800 101.800 188.200 102.200 ;
        RECT 201.400 106.800 201.800 107.200 ;
        RECT 199.000 105.800 199.400 106.200 ;
        RECT 198.200 105.100 198.600 105.500 ;
        RECT 203.000 105.800 203.400 106.200 ;
        RECT 205.400 105.800 205.800 106.200 ;
        RECT 211.800 106.800 212.200 107.200 ;
        RECT 215.000 105.900 215.400 106.300 ;
        RECT 211.800 104.800 212.200 105.200 ;
        RECT 212.600 105.100 213.000 105.500 ;
        RECT 219.800 103.800 220.200 104.200 ;
        RECT 222.200 104.800 222.600 105.200 ;
        RECT 221.400 101.800 221.800 102.200 ;
        RECT 237.400 108.800 237.800 109.200 ;
        RECT 241.400 108.800 241.800 109.200 ;
        RECT 227.800 105.800 228.200 106.200 ;
        RECT 231.800 106.800 232.200 107.200 ;
        RECT 250.200 108.800 250.600 109.200 ;
        RECT 227.000 104.800 227.400 105.200 ;
        RECT 240.600 104.800 241.000 105.200 ;
        RECT 2.200 98.800 2.600 99.200 ;
        RECT 12.600 96.800 13.000 97.200 ;
        RECT 2.200 94.800 2.600 95.200 ;
        RECT 7.000 94.800 7.400 95.200 ;
        RECT 3.000 93.800 3.400 94.200 ;
        RECT 3.800 93.100 4.200 93.500 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 17.400 94.800 17.800 95.200 ;
        RECT 6.200 92.800 6.600 93.200 ;
        RECT 15.800 92.800 16.200 93.200 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 23.000 93.800 23.400 94.200 ;
        RECT 23.800 93.800 24.200 94.200 ;
        RECT 27.800 94.800 28.200 95.200 ;
        RECT 30.200 94.800 30.600 95.200 ;
        RECT 47.800 98.800 48.200 99.200 ;
        RECT 29.400 93.800 29.800 94.200 ;
        RECT 31.800 93.800 32.200 94.200 ;
        RECT 32.600 93.100 33.000 93.500 ;
        RECT 26.200 91.800 26.600 92.200 ;
        RECT 35.000 92.800 35.400 93.200 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 46.200 94.800 46.600 95.200 ;
        RECT 43.000 93.800 43.400 94.200 ;
        RECT 44.600 93.800 45.000 94.200 ;
        RECT 60.600 96.800 61.000 97.200 ;
        RECT 51.000 94.800 51.400 95.200 ;
        RECT 55.000 94.800 55.400 95.200 ;
        RECT 52.600 93.800 53.000 94.200 ;
        RECT 41.400 91.800 41.800 92.200 ;
        RECT 51.800 93.100 52.200 93.500 ;
        RECT 61.400 94.800 61.800 95.200 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 83.800 98.800 84.200 99.200 ;
        RECT 70.200 94.800 70.600 95.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 93.400 98.800 93.800 99.200 ;
        RECT 71.000 93.800 71.400 94.200 ;
        RECT 75.800 93.800 76.200 94.200 ;
        RECT 75.000 93.100 75.400 93.500 ;
        RECT 63.800 91.800 64.200 92.200 ;
        RECT 89.400 94.800 89.800 95.200 ;
        RECT 95.000 98.800 95.400 99.200 ;
        RECT 84.600 93.100 85.000 93.500 ;
        RECT 102.200 95.800 102.600 96.200 ;
        RECT 112.600 96.800 113.000 97.200 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 99.800 93.800 100.200 94.200 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 103.800 93.100 104.200 93.500 ;
        RECT 116.600 98.800 117.000 99.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 95.000 91.800 95.400 92.200 ;
        RECT 106.200 92.800 106.600 93.200 ;
        RECT 134.200 98.800 134.600 99.200 ;
        RECT 121.400 94.800 121.800 95.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 124.600 94.000 125.000 94.400 ;
        RECT 133.400 93.800 133.800 94.200 ;
        RECT 120.600 91.800 121.000 92.200 ;
        RECT 136.600 98.800 137.000 99.200 ;
        RECT 139.800 98.800 140.200 99.200 ;
        RECT 147.000 98.800 147.400 99.200 ;
        RECT 131.800 91.800 132.200 92.200 ;
        RECT 136.600 91.800 137.000 92.200 ;
        RECT 139.800 92.800 140.200 93.200 ;
        RECT 143.000 91.800 143.400 92.200 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 167.800 96.200 168.200 96.600 ;
        RECT 169.400 95.500 169.800 95.900 ;
        RECT 179.000 98.800 179.400 99.200 ;
        RECT 173.400 94.800 173.800 95.200 ;
        RECT 169.400 93.100 169.800 93.500 ;
        RECT 159.000 91.800 159.400 92.200 ;
        RECT 170.200 93.100 170.600 93.500 ;
        RECT 187.000 96.200 187.400 96.600 ;
        RECT 188.600 95.500 189.000 95.900 ;
        RECT 189.400 93.800 189.800 94.200 ;
        RECT 188.600 93.100 189.000 93.500 ;
        RECT 179.800 91.800 180.200 92.200 ;
        RECT 193.400 94.800 193.800 95.200 ;
        RECT 194.200 93.800 194.600 94.200 ;
        RECT 202.200 96.200 202.600 96.600 ;
        RECT 203.800 95.500 204.200 95.900 ;
        RECT 215.000 98.800 215.400 99.200 ;
        RECT 207.800 94.800 208.200 95.200 ;
        RECT 209.400 94.800 209.800 95.200 ;
        RECT 210.200 94.800 210.600 95.200 ;
        RECT 203.800 93.100 204.200 93.500 ;
        RECT 208.600 93.800 209.000 94.200 ;
        RECT 195.000 91.800 195.400 92.200 ;
        RECT 215.800 93.800 216.200 94.200 ;
        RECT 223.800 96.200 224.200 96.600 ;
        RECT 225.400 95.500 225.800 95.900 ;
        RECT 228.600 94.800 229.000 95.200 ;
        RECT 230.200 94.800 230.600 95.200 ;
        RECT 229.400 93.800 229.800 94.200 ;
        RECT 225.400 93.100 225.800 93.500 ;
        RECT 231.800 93.800 232.200 94.200 ;
        RECT 234.200 93.800 234.600 94.200 ;
        RECT 235.800 93.800 236.200 94.200 ;
        RECT 216.600 91.800 217.000 92.200 ;
        RECT 235.000 93.100 235.400 93.500 ;
        RECT 247.000 94.800 247.400 95.200 ;
        RECT 247.800 94.800 248.200 95.200 ;
        RECT 246.200 93.800 246.600 94.200 ;
        RECT 251.000 94.800 251.400 95.200 ;
        RECT 243.800 91.800 244.200 92.200 ;
        RECT 6.200 88.800 6.600 89.200 ;
        RECT 7.800 84.800 8.200 85.200 ;
        RECT 11.000 86.800 11.400 87.200 ;
        RECT 14.200 85.800 14.600 86.200 ;
        RECT 10.200 85.100 10.600 85.500 ;
        RECT 19.000 83.800 19.400 84.200 ;
        RECT 19.800 88.800 20.200 89.200 ;
        RECT 22.200 86.100 22.600 86.500 ;
        RECT 26.200 85.900 26.600 86.300 ;
        RECT 30.200 85.800 30.600 86.200 ;
        RECT 28.600 85.100 29.000 85.500 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 31.800 81.800 32.200 82.200 ;
        RECT 45.400 88.800 45.800 89.200 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 53.400 86.800 53.800 87.200 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 47.800 86.100 48.200 86.500 ;
        RECT 43.800 84.800 44.200 85.200 ;
        RECT 54.200 85.100 54.600 85.500 ;
        RECT 60.600 86.800 61.000 87.200 ;
        RECT 65.400 88.800 65.800 89.200 ;
        RECT 58.200 84.800 58.600 85.200 ;
        RECT 61.400 85.800 61.800 86.200 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 73.400 86.800 73.800 87.200 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 67.800 86.100 68.200 86.500 ;
        RECT 63.000 81.800 63.400 82.200 ;
        RECT 81.400 86.800 81.800 87.200 ;
        RECT 74.200 85.100 74.600 85.500 ;
        RECT 82.200 84.800 82.600 85.200 ;
        RECT 84.600 86.800 85.000 87.200 ;
        RECT 84.600 84.800 85.000 85.200 ;
        RECT 83.000 81.800 83.400 82.200 ;
        RECT 95.800 88.800 96.200 89.200 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 87.000 84.800 87.400 85.200 ;
        RECT 91.800 85.800 92.200 86.200 ;
        RECT 91.800 84.800 92.200 85.200 ;
        RECT 102.200 88.800 102.600 89.200 ;
        RECT 104.600 88.800 105.000 89.200 ;
        RECT 94.200 86.800 94.600 87.200 ;
        RECT 92.600 81.800 93.000 82.200 ;
        RECT 95.800 84.800 96.200 85.200 ;
        RECT 96.600 84.800 97.000 85.200 ;
        RECT 100.600 86.800 101.000 87.200 ;
        RECT 97.400 81.800 97.800 82.200 ;
        RECT 102.200 84.800 102.600 85.200 ;
        RECT 101.400 81.800 101.800 82.200 ;
        RECT 114.200 88.800 114.600 89.200 ;
        RECT 110.200 85.800 110.600 86.200 ;
        RECT 104.600 84.800 105.000 85.200 ;
        RECT 105.400 85.100 105.800 85.500 ;
        RECT 103.800 81.800 104.200 82.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 131.000 88.800 131.400 89.200 ;
        RECT 118.200 84.800 118.600 85.200 ;
        RECT 124.600 85.800 125.000 86.200 ;
        RECT 127.000 85.800 127.400 86.200 ;
        RECT 128.600 84.800 129.000 85.200 ;
        RECT 140.600 88.800 141.000 89.200 ;
        RECT 133.400 86.100 133.800 86.500 ;
        RECT 159.000 88.800 159.400 89.200 ;
        RECT 148.600 86.800 149.000 87.200 ;
        RECT 143.000 86.100 143.400 86.500 ;
        RECT 139.800 85.100 140.200 85.500 ;
        RECT 147.000 85.900 147.400 86.300 ;
        RECT 149.400 85.100 149.800 85.500 ;
        RECT 153.400 84.800 153.800 85.200 ;
        RECT 158.200 86.800 158.600 87.200 ;
        RECT 171.000 88.800 171.400 89.200 ;
        RECT 167.000 85.800 167.400 86.200 ;
        RECT 169.400 86.800 169.800 87.200 ;
        RECT 170.200 85.800 170.600 86.200 ;
        RECT 175.800 86.800 176.200 87.200 ;
        RECT 173.400 86.100 173.800 86.500 ;
        RECT 163.000 81.800 163.400 82.200 ;
        RECT 204.600 88.800 205.000 89.200 ;
        RECT 179.800 85.100 180.200 85.500 ;
        RECT 182.200 85.800 182.600 86.200 ;
        RECT 188.600 85.800 189.000 86.200 ;
        RECT 187.800 81.800 188.200 82.200 ;
        RECT 192.600 81.800 193.000 82.200 ;
        RECT 196.600 84.800 197.000 85.200 ;
        RECT 203.000 85.800 203.400 86.200 ;
        RECT 220.600 88.800 221.000 89.200 ;
        RECT 212.600 86.800 213.000 87.200 ;
        RECT 207.000 86.100 207.400 86.500 ;
        RECT 199.000 84.800 199.400 85.200 ;
        RECT 201.400 84.800 201.800 85.200 ;
        RECT 215.000 85.800 215.400 86.200 ;
        RECT 213.400 85.100 213.800 85.500 ;
        RECT 240.600 88.800 241.000 89.200 ;
        RECT 226.200 86.800 226.600 87.200 ;
        RECT 220.600 84.800 221.000 85.200 ;
        RECT 232.600 86.800 233.000 87.200 ;
        RECT 245.400 88.800 245.800 89.200 ;
        RECT 223.800 81.800 224.200 82.200 ;
        RECT 234.200 85.900 234.600 86.300 ;
        RECT 227.800 84.800 228.200 85.200 ;
        RECT 230.200 84.800 230.600 85.200 ;
        RECT 231.800 85.100 232.200 85.500 ;
        RECT 243.800 85.800 244.200 86.200 ;
        RECT 251.000 86.800 251.400 87.200 ;
        RECT 243.800 84.800 244.200 85.200 ;
        RECT 0.600 73.100 1.000 73.500 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 19.800 74.800 20.200 75.200 ;
        RECT 14.200 71.800 14.600 72.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 23.000 73.800 23.400 74.200 ;
        RECT 30.200 74.800 30.600 75.200 ;
        RECT 43.800 76.800 44.200 77.200 ;
        RECT 32.600 73.800 33.000 74.200 ;
        RECT 25.400 71.800 25.800 72.200 ;
        RECT 28.600 72.800 29.000 73.200 ;
        RECT 34.200 73.800 34.600 74.200 ;
        RECT 35.800 73.800 36.200 74.200 ;
        RECT 35.000 73.100 35.400 73.500 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 45.400 74.800 45.800 75.200 ;
        RECT 56.600 76.800 57.000 77.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 47.800 73.800 48.200 74.200 ;
        RECT 63.800 76.200 64.200 76.600 ;
        RECT 65.400 75.500 65.800 75.900 ;
        RECT 71.000 78.800 71.400 79.200 ;
        RECT 65.400 73.100 65.800 73.500 ;
        RECT 68.600 74.800 69.000 75.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 67.000 71.800 67.400 72.200 ;
        RECT 81.400 74.800 81.800 75.200 ;
        RECT 77.400 73.800 77.800 74.200 ;
        RECT 78.200 73.100 78.600 73.500 ;
        RECT 91.800 73.800 92.200 74.200 ;
        RECT 95.000 78.800 95.400 79.200 ;
        RECT 95.800 73.800 96.200 74.200 ;
        RECT 96.600 73.800 97.000 74.200 ;
        RECT 87.000 71.800 87.400 72.200 ;
        RECT 89.400 71.800 89.800 72.200 ;
        RECT 102.200 74.800 102.600 75.200 ;
        RECT 103.000 73.800 103.400 74.200 ;
        RECT 107.800 78.800 108.200 79.200 ;
        RECT 107.000 73.800 107.400 74.200 ;
        RECT 100.600 71.800 101.000 72.200 ;
        RECT 117.400 74.800 117.800 75.200 ;
        RECT 118.200 74.800 118.600 75.200 ;
        RECT 123.000 74.800 123.400 75.200 ;
        RECT 106.200 71.800 106.600 72.200 ;
        RECT 108.600 71.800 109.000 72.200 ;
        RECT 111.800 72.800 112.200 73.200 ;
        RECT 113.400 72.800 113.800 73.200 ;
        RECT 119.000 73.800 119.400 74.200 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 127.800 74.800 128.200 75.200 ;
        RECT 132.600 74.800 133.000 75.200 ;
        RECT 123.000 72.800 123.400 73.200 ;
        RECT 133.400 74.800 133.800 75.200 ;
        RECT 139.800 78.800 140.200 79.200 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 141.400 78.800 141.800 79.200 ;
        RECT 140.600 73.800 141.000 74.200 ;
        RECT 147.800 76.800 148.200 77.200 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 155.000 76.200 155.400 76.600 ;
        RECT 156.600 75.500 157.000 75.900 ;
        RECT 157.400 76.800 157.800 77.200 ;
        RECT 151.800 74.800 152.200 75.200 ;
        RECT 163.800 78.800 164.200 79.200 ;
        RECT 157.400 73.800 157.800 74.200 ;
        RECT 156.600 73.100 157.000 73.500 ;
        RECT 167.800 74.800 168.200 75.200 ;
        RECT 171.000 73.800 171.400 74.200 ;
        RECT 172.600 73.800 173.000 74.200 ;
        RECT 171.800 73.100 172.200 73.500 ;
        RECT 183.000 74.800 183.400 75.200 ;
        RECT 184.600 74.800 185.000 75.200 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 183.800 73.800 184.200 74.200 ;
        RECT 188.600 74.800 189.000 75.200 ;
        RECT 189.400 74.800 189.800 75.200 ;
        RECT 190.200 74.800 190.600 75.200 ;
        RECT 187.800 73.800 188.200 74.200 ;
        RECT 180.600 71.800 181.000 72.200 ;
        RECT 181.400 72.800 181.800 73.200 ;
        RECT 200.600 78.800 201.000 79.200 ;
        RECT 199.000 73.800 199.400 74.200 ;
        RECT 199.800 73.800 200.200 74.200 ;
        RECT 207.800 74.800 208.200 75.200 ;
        RECT 208.600 74.800 209.000 75.200 ;
        RECT 211.800 74.800 212.200 75.200 ;
        RECT 212.600 73.800 213.000 74.200 ;
        RECT 215.000 73.800 215.400 74.200 ;
        RECT 225.400 76.800 225.800 77.200 ;
        RECT 219.800 73.800 220.200 74.200 ;
        RECT 223.800 74.800 224.200 75.200 ;
        RECT 224.600 74.800 225.000 75.200 ;
        RECT 232.600 76.200 233.000 76.600 ;
        RECT 234.200 75.500 234.600 75.900 ;
        RECT 231.800 72.800 232.200 73.200 ;
        RECT 234.200 73.100 234.600 73.500 ;
        RECT 242.200 72.800 242.600 73.200 ;
        RECT 251.800 74.800 252.200 75.200 ;
        RECT 250.200 73.800 250.600 74.200 ;
        RECT 240.600 71.800 241.000 72.200 ;
        RECT 245.400 71.800 245.800 72.200 ;
        RECT 247.800 71.800 248.200 72.200 ;
        RECT 3.000 68.800 3.400 69.200 ;
        RECT 19.800 68.800 20.200 69.200 ;
        RECT 2.200 64.800 2.600 65.200 ;
        RECT 11.800 66.800 12.200 67.200 ;
        RECT 15.000 66.800 15.400 67.200 ;
        RECT 7.800 65.800 8.200 66.200 ;
        RECT 11.000 65.100 11.400 65.500 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 25.400 65.800 25.800 66.200 ;
        RECT 20.600 65.100 21.000 65.500 ;
        RECT 33.400 66.800 33.800 67.200 ;
        RECT 29.400 63.800 29.800 64.200 ;
        RECT 34.200 65.800 34.600 66.200 ;
        RECT 39.800 66.800 40.200 67.200 ;
        RECT 38.200 65.800 38.600 66.200 ;
        RECT 40.600 65.800 41.000 66.200 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 45.400 65.800 45.800 66.200 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 55.800 66.800 56.200 67.200 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 51.800 63.800 52.200 64.200 ;
        RECT 57.400 63.800 57.800 64.200 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 67.000 66.800 67.400 67.200 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 78.200 67.800 78.600 68.200 ;
        RECT 96.600 68.800 97.000 69.200 ;
        RECT 63.800 64.800 64.200 65.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 71.800 65.800 72.200 66.200 ;
        RECT 76.600 66.800 77.000 67.200 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 85.400 66.800 85.800 67.200 ;
        RECT 89.400 66.800 89.800 67.200 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 87.800 61.800 88.200 62.200 ;
        RECT 104.600 66.800 105.000 67.200 ;
        RECT 99.000 66.100 99.400 66.500 ;
        RECT 94.200 64.800 94.600 65.200 ;
        RECT 109.400 68.800 109.800 69.200 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 105.400 65.100 105.800 65.500 ;
        RECT 96.600 61.800 97.000 62.200 ;
        RECT 109.400 64.800 109.800 65.200 ;
        RECT 119.000 68.800 119.400 69.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 111.800 64.800 112.200 65.200 ;
        RECT 112.600 64.800 113.000 65.200 ;
        RECT 115.000 65.800 115.400 66.200 ;
        RECT 118.200 65.800 118.600 66.200 ;
        RECT 121.400 66.100 121.800 66.500 ;
        RECT 125.400 65.900 125.800 66.300 ;
        RECT 127.800 65.100 128.200 65.500 ;
        RECT 130.200 64.800 130.600 65.200 ;
        RECT 135.000 66.800 135.400 67.200 ;
        RECT 159.800 68.800 160.200 69.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 142.200 65.900 142.600 66.300 ;
        RECT 139.800 65.100 140.200 65.500 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 155.800 65.800 156.200 66.200 ;
        RECT 148.600 61.800 149.000 62.200 ;
        RECT 151.000 65.100 151.400 65.500 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 162.200 64.800 162.600 65.200 ;
        RECT 183.800 68.800 184.200 69.200 ;
        RECT 168.600 66.800 169.000 67.200 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 179.000 65.800 179.400 66.200 ;
        RECT 175.000 65.100 175.400 65.500 ;
        RECT 184.600 64.800 185.000 65.200 ;
        RECT 189.400 67.800 189.800 68.200 ;
        RECT 193.400 68.800 193.800 69.200 ;
        RECT 187.800 65.800 188.200 66.200 ;
        RECT 194.200 66.800 194.600 67.200 ;
        RECT 191.800 65.800 192.200 66.200 ;
        RECT 195.000 65.800 195.400 66.200 ;
        RECT 211.000 68.800 211.400 69.200 ;
        RECT 215.800 68.800 216.200 69.200 ;
        RECT 204.600 66.800 205.000 67.200 ;
        RECT 205.400 65.800 205.800 66.200 ;
        RECT 209.400 65.800 209.800 66.200 ;
        RECT 232.600 68.800 233.000 69.200 ;
        RECT 223.800 66.800 224.200 67.200 ;
        RECT 218.200 66.100 218.600 66.500 ;
        RECT 215.000 64.800 215.400 65.200 ;
        RECT 226.200 65.800 226.600 66.200 ;
        RECT 224.600 65.100 225.000 65.500 ;
        RECT 251.000 68.800 251.400 69.200 ;
        RECT 240.600 66.800 241.000 67.200 ;
        RECT 235.000 66.100 235.400 66.500 ;
        RECT 231.800 64.800 232.200 65.200 ;
        RECT 231.000 61.800 231.400 62.200 ;
        RECT 239.000 65.900 239.400 66.300 ;
        RECT 241.400 65.100 241.800 65.500 ;
        RECT 242.200 65.100 242.600 65.500 ;
        RECT 15.000 57.800 15.400 58.200 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 4.600 54.800 5.000 55.200 ;
        RECT 25.400 56.800 25.800 57.200 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 7.000 53.800 7.400 54.200 ;
        RECT 6.200 53.100 6.600 53.500 ;
        RECT 19.000 54.800 19.400 55.200 ;
        RECT 16.600 53.800 17.000 54.200 ;
        RECT 15.800 53.100 16.200 53.500 ;
        RECT 25.400 53.800 25.800 54.200 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 30.200 53.800 30.600 54.200 ;
        RECT 38.200 56.200 38.600 56.600 ;
        RECT 43.000 58.800 43.400 59.200 ;
        RECT 39.800 55.500 40.200 55.900 ;
        RECT 54.200 58.800 54.600 59.200 ;
        RECT 43.800 54.800 44.200 55.200 ;
        RECT 44.600 54.800 45.000 55.200 ;
        RECT 45.400 54.800 45.800 55.200 ;
        RECT 46.200 54.800 46.600 55.200 ;
        RECT 51.800 54.800 52.200 55.200 ;
        RECT 52.600 54.800 53.000 55.200 ;
        RECT 39.800 53.100 40.200 53.500 ;
        RECT 31.000 51.800 31.400 52.200 ;
        RECT 59.800 52.800 60.200 53.200 ;
        RECT 63.800 54.800 64.200 55.200 ;
        RECT 77.400 56.800 77.800 57.200 ;
        RECT 66.200 53.800 66.600 54.200 ;
        RECT 67.800 53.800 68.200 54.200 ;
        RECT 69.400 53.800 69.800 54.200 ;
        RECT 58.200 51.800 58.600 52.200 ;
        RECT 60.600 51.800 61.000 52.200 ;
        RECT 68.600 53.100 69.000 53.500 ;
        RECT 79.800 54.800 80.200 55.200 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 87.800 54.800 88.200 55.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 99.000 56.800 99.400 57.200 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 93.400 54.800 93.800 55.200 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 106.200 56.200 106.600 56.600 ;
        RECT 107.800 55.500 108.200 55.900 ;
        RECT 115.800 58.800 116.200 59.200 ;
        RECT 108.600 53.800 109.000 54.200 ;
        RECT 107.800 53.100 108.200 53.500 ;
        RECT 112.600 54.800 113.000 55.200 ;
        RECT 113.400 53.800 113.800 54.200 ;
        RECT 114.200 52.800 114.600 53.200 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 123.000 58.800 123.400 59.200 ;
        RECT 120.600 54.800 121.000 55.200 ;
        RECT 121.400 54.800 121.800 55.200 ;
        RECT 139.800 58.800 140.200 59.200 ;
        RECT 119.800 52.800 120.200 53.200 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 127.000 53.800 127.400 54.200 ;
        RECT 130.200 53.800 130.600 54.200 ;
        RECT 131.000 53.100 131.400 53.500 ;
        RECT 133.400 52.800 133.800 53.200 ;
        RECT 149.400 54.800 149.800 55.200 ;
        RECT 150.200 54.800 150.600 55.200 ;
        RECT 153.400 54.800 153.800 55.200 ;
        RECT 155.000 53.800 155.400 54.200 ;
        RECT 142.200 51.800 142.600 52.200 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 157.400 53.800 157.800 54.200 ;
        RECT 159.000 53.800 159.400 54.200 ;
        RECT 158.200 53.100 158.600 53.500 ;
        RECT 167.000 51.800 167.400 52.200 ;
        RECT 175.000 56.200 175.400 56.600 ;
        RECT 176.600 55.500 177.000 55.900 ;
        RECT 182.200 54.800 182.600 55.200 ;
        RECT 195.000 58.800 195.400 59.200 ;
        RECT 176.600 53.100 177.000 53.500 ;
        RECT 167.800 51.800 168.200 52.200 ;
        RECT 177.400 53.100 177.800 53.500 ;
        RECT 206.200 58.800 206.600 59.200 ;
        RECT 195.800 54.800 196.200 55.200 ;
        RECT 196.600 54.800 197.000 55.200 ;
        RECT 186.200 51.800 186.600 52.200 ;
        RECT 191.800 52.800 192.200 53.200 ;
        RECT 197.400 52.800 197.800 53.200 ;
        RECT 203.000 54.800 203.400 55.200 ;
        RECT 214.200 54.800 214.600 55.200 ;
        RECT 200.600 51.800 201.000 52.200 ;
        RECT 222.200 56.200 222.600 56.600 ;
        RECT 227.800 58.800 228.200 59.200 ;
        RECT 223.800 55.500 224.200 55.900 ;
        RECT 223.800 53.100 224.200 53.500 ;
        RECT 215.000 51.800 215.400 52.200 ;
        RECT 235.000 56.200 235.400 56.600 ;
        RECT 236.600 55.500 237.000 55.900 ;
        RECT 240.600 58.800 241.000 59.200 ;
        RECT 239.000 54.800 239.400 55.200 ;
        RECT 236.600 53.100 237.000 53.500 ;
        RECT 239.800 53.800 240.200 54.200 ;
        RECT 247.800 56.200 248.200 56.600 ;
        RECT 249.400 55.500 249.800 55.900 ;
        RECT 249.400 53.100 249.800 53.500 ;
        RECT 3.800 48.800 4.200 49.200 ;
        RECT 24.600 48.800 25.000 49.200 ;
        RECT 9.400 46.800 9.800 47.200 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 27.800 48.800 28.200 49.200 ;
        RECT 3.800 41.800 4.200 42.200 ;
        RECT 18.200 45.900 18.600 46.300 ;
        RECT 11.800 44.800 12.200 45.200 ;
        RECT 14.200 44.800 14.600 45.200 ;
        RECT 15.800 45.100 16.200 45.500 ;
        RECT 32.600 48.800 33.000 49.200 ;
        RECT 31.800 44.800 32.200 45.200 ;
        RECT 46.200 48.800 46.600 49.200 ;
        RECT 51.000 48.800 51.400 49.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 38.200 46.100 38.600 46.500 ;
        RECT 42.200 45.900 42.600 46.300 ;
        RECT 44.600 45.100 45.000 45.500 ;
        RECT 35.800 43.800 36.200 44.200 ;
        RECT 70.200 48.800 70.600 49.200 ;
        RECT 59.800 46.800 60.200 47.200 ;
        RECT 62.200 46.800 62.600 47.200 ;
        RECT 54.200 46.100 54.600 46.500 ;
        RECT 58.200 45.900 58.600 46.300 ;
        RECT 60.600 45.100 61.000 45.500 ;
        RECT 61.400 45.100 61.800 45.500 ;
        RECT 72.600 46.800 73.000 47.200 ;
        RECT 85.400 48.800 85.800 49.200 ;
        RECT 77.400 46.800 77.800 47.200 ;
        RECT 91.800 48.800 92.200 49.200 ;
        RECT 74.200 44.800 74.600 45.200 ;
        RECT 76.600 45.100 77.000 45.500 ;
        RECT 87.800 44.800 88.200 45.200 ;
        RECT 109.400 48.800 109.800 49.200 ;
        RECT 99.800 46.800 100.200 47.200 ;
        RECT 94.200 46.100 94.600 46.500 ;
        RECT 98.200 45.900 98.600 46.300 ;
        RECT 112.600 47.800 113.000 48.200 ;
        RECT 100.600 45.100 101.000 45.500 ;
        RECT 104.600 44.800 105.000 45.200 ;
        RECT 111.000 45.800 111.400 46.200 ;
        RECT 118.200 46.800 118.600 47.200 ;
        RECT 122.200 46.800 122.600 47.200 ;
        RECT 122.200 44.800 122.600 45.200 ;
        RECT 135.800 48.800 136.200 49.200 ;
        RECT 132.600 46.800 133.000 47.200 ;
        RECT 127.000 46.100 127.400 46.500 ;
        RECT 133.400 45.100 133.800 45.500 ;
        RECT 138.200 47.800 138.600 48.200 ;
        RECT 149.400 48.800 149.800 49.200 ;
        RECT 142.200 45.900 142.600 46.300 ;
        RECT 139.800 45.100 140.200 45.500 ;
        RECT 158.200 48.800 158.600 49.200 ;
        RECT 162.200 48.800 162.600 49.200 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 157.400 44.800 157.800 45.200 ;
        RECT 168.600 48.800 169.000 49.200 ;
        RECT 175.800 48.800 176.200 49.200 ;
        RECT 165.400 41.800 165.800 42.200 ;
        RECT 172.600 41.800 173.000 42.200 ;
        RECT 190.200 48.800 190.600 49.200 ;
        RECT 192.600 48.800 193.000 49.200 ;
        RECT 180.600 46.800 181.000 47.200 ;
        RECT 178.200 41.800 178.600 42.200 ;
        RECT 186.200 41.800 186.600 42.200 ;
        RECT 191.000 45.800 191.400 46.200 ;
        RECT 203.000 46.800 203.400 47.200 ;
        RECT 208.600 48.800 209.000 49.200 ;
        RECT 195.000 46.100 195.400 46.500 ;
        RECT 199.000 45.900 199.400 46.300 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 201.400 45.100 201.800 45.500 ;
        RECT 211.000 46.100 211.400 46.500 ;
        RECT 215.000 45.900 215.400 46.300 ;
        RECT 217.400 45.100 217.800 45.500 ;
        RECT 219.800 44.800 220.200 45.200 ;
        RECT 225.400 45.800 225.800 46.200 ;
        RECT 239.000 46.800 239.400 47.200 ;
        RECT 250.200 48.800 250.600 49.200 ;
        RECT 242.200 46.800 242.600 47.200 ;
        RECT 243.800 45.900 244.200 46.300 ;
        RECT 239.000 44.800 239.400 45.200 ;
        RECT 241.400 45.100 241.800 45.500 ;
        RECT 12.600 38.800 13.000 39.200 ;
        RECT 0.600 33.100 1.000 33.500 ;
        RECT 13.400 34.800 13.800 35.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 15.800 34.800 16.200 35.200 ;
        RECT 29.400 36.800 29.800 37.200 ;
        RECT 18.200 33.800 18.600 34.200 ;
        RECT 32.600 38.800 33.000 39.200 ;
        RECT 37.400 38.800 37.800 39.200 ;
        RECT 19.800 33.800 20.200 34.200 ;
        RECT 21.400 33.800 21.800 34.200 ;
        RECT 20.600 33.100 21.000 33.500 ;
        RECT 30.200 34.800 30.600 35.200 ;
        RECT 31.000 34.800 31.400 35.200 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 39.000 34.800 39.400 35.200 ;
        RECT 46.200 38.800 46.600 39.200 ;
        RECT 39.800 33.800 40.200 34.200 ;
        RECT 43.800 34.800 44.200 35.200 ;
        RECT 47.800 34.800 48.200 35.200 ;
        RECT 58.200 38.800 58.600 39.200 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 42.200 31.800 42.600 32.200 ;
        RECT 55.000 34.800 55.400 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 56.600 34.800 57.000 35.200 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 63.800 34.800 64.200 35.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 71.000 38.800 71.400 39.200 ;
        RECT 82.200 36.800 82.600 37.200 ;
        RECT 52.600 32.800 53.000 33.200 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 72.600 34.800 73.000 35.200 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 73.400 33.100 73.800 33.500 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 93.400 38.800 93.800 39.200 ;
        RECT 94.200 34.800 94.600 35.200 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 84.600 31.800 85.000 32.200 ;
        RECT 88.600 32.800 89.000 33.200 ;
        RECT 98.200 34.800 98.600 35.200 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 104.600 34.800 105.000 35.200 ;
        RECT 106.200 34.800 106.600 35.200 ;
        RECT 118.200 36.800 118.600 37.200 ;
        RECT 119.800 36.800 120.200 37.200 ;
        RECT 96.600 32.800 97.000 33.200 ;
        RECT 107.800 33.800 108.200 34.200 ;
        RECT 110.200 33.800 110.600 34.200 ;
        RECT 111.000 33.100 111.400 33.500 ;
        RECT 120.600 34.800 121.000 35.200 ;
        RECT 121.400 34.800 121.800 35.200 ;
        RECT 130.200 36.800 130.600 37.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 129.400 34.800 129.800 35.200 ;
        RECT 137.400 36.200 137.800 36.600 ;
        RECT 139.000 35.500 139.400 35.900 ;
        RECT 139.800 33.800 140.200 34.200 ;
        RECT 136.600 32.800 137.000 33.200 ;
        RECT 139.000 33.100 139.400 33.500 ;
        RECT 143.000 38.800 143.400 39.200 ;
        RECT 147.800 34.800 148.200 35.200 ;
        RECT 148.600 34.800 149.000 35.200 ;
        RECT 158.200 36.200 158.600 36.600 ;
        RECT 161.400 38.800 161.800 39.200 ;
        RECT 159.800 35.500 160.200 35.900 ;
        RECT 157.400 32.800 157.800 33.200 ;
        RECT 151.000 31.800 151.400 32.200 ;
        RECT 159.800 33.100 160.200 33.500 ;
        RECT 167.000 33.800 167.400 34.200 ;
        RECT 161.400 31.800 161.800 32.200 ;
        RECT 169.400 34.800 169.800 35.200 ;
        RECT 170.200 34.800 170.600 35.200 ;
        RECT 179.800 38.800 180.200 39.200 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 177.400 34.800 177.800 35.200 ;
        RECT 178.200 34.800 178.600 35.200 ;
        RECT 187.800 36.800 188.200 37.200 ;
        RECT 186.200 35.800 186.600 36.200 ;
        RECT 167.800 31.800 168.200 32.200 ;
        RECT 182.200 33.800 182.600 34.200 ;
        RECT 175.800 31.800 176.200 32.200 ;
        RECT 186.200 34.800 186.600 35.200 ;
        RECT 187.000 33.800 187.400 34.200 ;
        RECT 195.000 36.200 195.400 36.600 ;
        RECT 196.600 35.500 197.000 35.900 ;
        RECT 191.800 34.800 192.200 35.200 ;
        RECT 197.400 34.800 197.800 35.200 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 196.600 33.100 197.000 33.500 ;
        RECT 211.000 36.200 211.400 36.600 ;
        RECT 212.600 35.500 213.000 35.900 ;
        RECT 212.600 33.100 213.000 33.500 ;
        RECT 215.800 34.800 216.200 35.200 ;
        RECT 216.600 34.800 217.000 35.200 ;
        RECT 215.000 33.800 215.400 34.200 ;
        RECT 219.800 34.800 220.200 35.200 ;
        RECT 221.400 34.800 221.800 35.200 ;
        RECT 219.000 33.800 219.400 34.200 ;
        RECT 226.200 33.800 226.600 34.200 ;
        RECT 229.400 34.800 229.800 35.200 ;
        RECT 230.200 34.800 230.600 35.200 ;
        RECT 214.200 31.800 214.600 32.200 ;
        RECT 223.000 31.800 223.400 32.200 ;
        RECT 231.000 32.800 231.400 33.200 ;
        RECT 237.400 34.800 237.800 35.200 ;
        RECT 251.000 36.800 251.400 37.200 ;
        RECT 239.800 33.800 240.200 34.200 ;
        RECT 241.400 33.800 241.800 34.200 ;
        RECT 243.000 33.800 243.400 34.200 ;
        RECT 234.200 31.800 234.600 32.200 ;
        RECT 242.200 33.100 242.600 33.500 ;
        RECT 3.000 28.800 3.400 29.200 ;
        RECT 20.600 28.800 21.000 29.200 ;
        RECT 2.200 24.800 2.600 25.200 ;
        RECT 30.200 28.800 30.600 29.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 14.200 25.900 14.600 26.300 ;
        RECT 7.800 24.800 8.200 25.200 ;
        RECT 10.200 24.800 10.600 25.200 ;
        RECT 11.800 25.100 12.200 25.500 ;
        RECT 21.400 25.100 21.800 25.500 ;
        RECT 31.000 28.800 31.400 29.200 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 33.400 26.100 33.800 26.500 ;
        RECT 37.400 25.900 37.800 26.300 ;
        RECT 54.200 28.800 54.600 29.200 ;
        RECT 48.600 26.800 49.000 27.200 ;
        RECT 43.000 26.100 43.400 26.500 ;
        RECT 39.800 25.100 40.200 25.500 ;
        RECT 47.000 25.900 47.400 26.300 ;
        RECT 58.200 26.800 58.600 27.200 ;
        RECT 49.400 25.100 49.800 25.500 ;
        RECT 40.600 22.800 41.000 23.200 ;
        RECT 55.000 25.800 55.400 26.200 ;
        RECT 71.000 28.800 71.400 29.200 ;
        RECT 66.200 26.800 66.600 27.200 ;
        RECT 59.800 24.800 60.200 25.200 ;
        RECT 62.200 25.100 62.600 25.500 ;
        RECT 85.400 28.800 85.800 29.200 ;
        RECT 72.600 25.800 73.000 26.200 ;
        RECT 78.200 24.800 78.600 25.200 ;
        RECT 83.800 25.800 84.200 26.200 ;
        RECT 96.600 28.800 97.000 29.200 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 87.800 26.100 88.200 26.500 ;
        RECT 84.600 24.800 85.000 25.200 ;
        RECT 99.000 26.100 99.400 26.500 ;
        RECT 103.000 25.900 103.400 26.300 ;
        RECT 94.200 25.100 94.600 25.500 ;
        RECT 105.400 25.100 105.800 25.500 ;
        RECT 107.800 24.800 108.200 25.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 119.800 25.900 120.200 26.300 ;
        RECT 115.000 24.800 115.400 25.200 ;
        RECT 117.400 25.100 117.800 25.500 ;
        RECT 130.200 26.800 130.600 27.200 ;
        RECT 141.400 28.800 141.800 29.200 ;
        RECT 133.400 26.800 133.800 27.200 ;
        RECT 142.200 28.800 142.600 29.200 ;
        RECT 135.000 25.900 135.400 26.300 ;
        RECT 126.200 23.800 126.600 24.200 ;
        RECT 130.200 24.800 130.600 25.200 ;
        RECT 132.600 25.100 133.000 25.500 ;
        RECT 158.200 28.800 158.600 29.200 ;
        RECT 148.600 25.800 149.000 26.200 ;
        RECT 155.000 25.800 155.400 26.200 ;
        RECT 162.200 28.800 162.600 29.200 ;
        RECT 167.000 28.800 167.400 29.200 ;
        RECT 171.800 28.800 172.200 29.200 ;
        RECT 158.200 21.800 158.600 22.200 ;
        RECT 161.400 24.800 161.800 25.200 ;
        RECT 169.400 26.800 169.800 27.200 ;
        RECT 176.600 26.800 177.000 27.200 ;
        RECT 187.000 28.800 187.400 29.200 ;
        RECT 174.200 26.100 174.600 26.500 ;
        RECT 180.600 25.100 181.000 25.500 ;
        RECT 195.000 26.800 195.400 27.200 ;
        RECT 204.600 28.800 205.000 29.200 ;
        RECT 189.400 26.100 189.800 26.500 ;
        RECT 183.000 24.800 183.400 25.200 ;
        RECT 185.400 24.800 185.800 25.200 ;
        RECT 195.800 25.100 196.200 25.500 ;
        RECT 208.600 28.800 209.000 29.200 ;
        RECT 199.800 25.800 200.200 26.200 ;
        RECT 211.800 26.800 212.200 27.200 ;
        RECT 218.200 28.800 218.600 29.200 ;
        RECT 204.600 21.800 205.000 22.200 ;
        RECT 207.800 24.800 208.200 25.200 ;
        RECT 215.000 25.800 215.400 26.200 ;
        RECT 214.200 24.800 214.600 25.200 ;
        RECT 217.400 25.800 217.800 26.200 ;
        RECT 230.200 28.800 230.600 29.200 ;
        RECT 220.600 26.100 221.000 26.500 ;
        RECT 222.200 25.800 222.600 26.200 ;
        RECT 227.000 25.100 227.400 25.500 ;
        RECT 239.800 28.800 240.200 29.200 ;
        RECT 251.800 28.800 252.200 29.200 ;
        RECT 236.600 26.800 237.000 27.200 ;
        RECT 232.600 26.100 233.000 26.500 ;
        RECT 229.400 24.800 229.800 25.200 ;
        RECT 242.200 26.100 242.600 26.500 ;
        RECT 243.800 25.800 244.200 26.200 ;
        RECT 239.000 25.100 239.400 25.500 ;
        RECT 248.600 25.100 249.000 25.500 ;
        RECT 251.800 24.800 252.200 25.200 ;
        RECT 0.600 16.800 1.000 17.200 ;
        RECT 7.800 16.200 8.200 16.600 ;
        RECT 9.400 15.500 9.800 15.900 ;
        RECT 10.200 13.800 10.600 14.200 ;
        RECT 7.000 12.800 7.400 13.200 ;
        RECT 9.400 13.100 9.800 13.500 ;
        RECT 14.200 14.800 14.600 15.200 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 17.400 13.800 17.800 14.200 ;
        RECT 24.600 13.800 25.000 14.200 ;
        RECT 16.600 11.800 17.000 12.200 ;
        RECT 23.000 12.800 23.400 13.200 ;
        RECT 23.800 13.100 24.200 13.500 ;
        RECT 39.000 18.800 39.400 19.200 ;
        RECT 43.000 18.800 43.400 19.200 ;
        RECT 47.000 18.800 47.400 19.200 ;
        RECT 32.600 11.800 33.000 12.200 ;
        RECT 47.800 14.800 48.200 15.200 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 51.000 14.800 51.400 15.200 ;
        RECT 43.000 11.800 43.400 12.200 ;
        RECT 60.600 13.800 61.000 14.200 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 78.200 16.800 78.600 17.200 ;
        RECT 80.600 16.800 81.000 17.200 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 65.400 13.800 65.800 14.200 ;
        RECT 69.400 14.800 69.800 15.200 ;
        RECT 70.200 14.800 70.600 15.200 ;
        RECT 74.200 14.800 74.600 15.200 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 71.000 13.100 71.400 13.500 ;
        RECT 80.600 13.800 81.000 14.200 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 95.800 18.800 96.200 19.200 ;
        RECT 84.600 14.800 85.000 15.200 ;
        RECT 86.200 13.800 86.600 14.200 ;
        RECT 102.200 14.800 102.600 15.200 ;
        RECT 103.000 14.800 103.400 15.200 ;
        RECT 107.000 14.800 107.400 15.200 ;
        RECT 107.800 14.800 108.200 15.200 ;
        RECT 114.200 16.800 114.600 17.200 ;
        RECT 95.800 11.800 96.200 12.200 ;
        RECT 101.400 12.800 101.800 13.200 ;
        RECT 108.600 13.800 109.000 14.200 ;
        RECT 112.600 14.800 113.000 15.200 ;
        RECT 113.400 13.800 113.800 14.200 ;
        RECT 121.400 16.200 121.800 16.600 ;
        RECT 123.000 15.500 123.400 15.900 ;
        RECT 126.200 18.800 126.600 19.200 ;
        RECT 128.600 16.800 129.000 17.200 ;
        RECT 123.800 14.800 124.200 15.200 ;
        RECT 124.600 14.800 125.000 15.200 ;
        RECT 127.800 14.800 128.200 15.200 ;
        RECT 123.000 13.100 123.400 13.500 ;
        RECT 135.800 16.200 136.200 16.600 ;
        RECT 137.400 15.500 137.800 15.900 ;
        RECT 132.600 13.800 133.000 14.200 ;
        RECT 138.200 13.800 138.600 14.200 ;
        RECT 137.400 13.100 137.800 13.500 ;
        RECT 142.200 14.800 142.600 15.200 ;
        RECT 143.000 13.800 143.400 14.200 ;
        RECT 145.400 13.800 145.800 14.200 ;
        RECT 147.800 13.800 148.200 14.200 ;
        RECT 153.400 14.800 153.800 15.200 ;
        RECT 154.200 14.800 154.600 15.200 ;
        RECT 159.000 17.800 159.400 18.200 ;
        RECT 169.400 16.800 169.800 17.200 ;
        RECT 155.000 13.800 155.400 14.200 ;
        RECT 159.000 14.800 159.400 15.200 ;
        RECT 175.800 18.800 176.200 19.200 ;
        RECT 159.800 13.800 160.200 14.200 ;
        RECT 161.400 13.800 161.800 14.200 ;
        RECT 160.600 13.100 161.000 13.500 ;
        RECT 174.200 14.800 174.600 15.200 ;
        RECT 171.800 13.800 172.200 14.200 ;
        RECT 175.000 13.800 175.400 14.200 ;
        RECT 183.000 16.200 183.400 16.600 ;
        RECT 184.600 15.500 185.000 15.900 ;
        RECT 186.200 14.800 186.600 15.200 ;
        RECT 199.800 16.800 200.200 17.200 ;
        RECT 184.600 13.100 185.000 13.500 ;
        RECT 187.800 12.800 188.200 13.200 ;
        RECT 194.200 14.800 194.600 15.200 ;
        RECT 190.200 13.800 190.600 14.200 ;
        RECT 191.800 13.800 192.200 14.200 ;
        RECT 191.000 13.100 191.400 13.500 ;
        RECT 205.400 14.800 205.800 15.200 ;
        RECT 206.200 14.800 206.600 15.200 ;
        RECT 209.400 14.800 209.800 15.200 ;
        RECT 210.200 14.800 210.600 15.200 ;
        RECT 211.000 14.800 211.400 15.200 ;
        RECT 215.800 14.800 216.200 15.200 ;
        RECT 216.600 13.800 217.000 14.200 ;
        RECT 221.400 14.800 221.800 15.200 ;
        RECT 219.800 13.800 220.200 14.200 ;
        RECT 223.800 13.800 224.200 14.200 ;
        RECT 225.400 13.800 225.800 14.200 ;
        RECT 233.400 16.200 233.800 16.600 ;
        RECT 235.000 15.500 235.400 15.900 ;
        RECT 236.600 18.800 237.000 19.200 ;
        RECT 243.800 18.800 244.200 19.200 ;
        RECT 251.000 18.800 251.400 19.200 ;
        RECT 235.000 13.100 235.400 13.500 ;
        RECT 251.800 13.800 252.200 14.200 ;
        RECT 27.000 8.800 27.400 9.200 ;
        RECT 7.000 6.800 7.400 7.200 ;
        RECT 7.800 6.800 8.200 7.200 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 15.000 5.800 15.400 6.200 ;
        RECT 16.600 5.800 17.000 6.200 ;
        RECT 20.600 5.900 21.000 6.300 ;
        RECT 17.400 4.800 17.800 5.200 ;
        RECT 18.200 5.100 18.600 5.500 ;
        RECT 27.800 5.800 28.200 6.200 ;
        RECT 42.200 8.800 42.600 9.200 ;
        RECT 31.800 6.800 32.200 7.200 ;
        RECT 34.200 6.800 34.600 7.200 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 32.600 5.800 33.000 6.200 ;
        RECT 35.800 5.900 36.200 6.300 ;
        RECT 33.400 5.100 33.800 5.500 ;
        RECT 46.200 6.800 46.600 7.200 ;
        RECT 49.400 6.800 49.800 7.200 ;
        RECT 46.200 4.800 46.600 5.200 ;
        RECT 59.800 8.800 60.200 9.200 ;
        RECT 58.200 6.800 58.600 7.200 ;
        RECT 52.600 6.100 53.000 6.500 ;
        RECT 71.000 8.800 71.400 9.200 ;
        RECT 67.800 6.800 68.200 7.200 ;
        RECT 62.200 6.100 62.600 6.500 ;
        RECT 59.000 5.100 59.400 5.500 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 68.600 5.100 69.000 5.500 ;
        RECT 72.600 5.100 73.000 5.500 ;
        RECT 89.400 8.800 89.800 9.200 ;
        RECT 91.000 8.800 91.400 9.200 ;
        RECT 83.800 4.800 84.200 5.200 ;
        RECT 95.800 6.800 96.200 7.200 ;
        RECT 93.400 6.100 93.800 6.500 ;
        RECT 97.400 5.900 97.800 6.300 ;
        RECT 107.800 6.800 108.200 7.200 ;
        RECT 99.800 5.100 100.200 5.500 ;
        RECT 103.800 4.800 104.200 5.200 ;
        RECT 114.200 6.800 114.600 7.200 ;
        RECT 115.800 6.800 116.200 7.200 ;
        RECT 119.800 6.800 120.200 7.200 ;
        RECT 115.000 5.100 115.400 5.500 ;
        RECT 139.000 8.800 139.400 9.200 ;
        RECT 147.800 8.800 148.200 9.200 ;
        RECT 126.200 4.800 126.600 5.200 ;
        RECT 130.200 5.100 130.600 5.500 ;
        RECT 143.000 6.800 143.400 7.200 ;
        RECT 170.200 8.800 170.600 9.200 ;
        RECT 155.800 6.800 156.200 7.200 ;
        RECT 157.400 6.800 157.800 7.200 ;
        RECT 150.200 6.100 150.600 6.500 ;
        RECT 146.200 4.800 146.600 5.200 ;
        RECT 163.800 6.800 164.200 7.200 ;
        RECT 156.600 5.100 157.000 5.500 ;
        RECT 194.200 8.800 194.600 9.200 ;
        RECT 178.200 6.800 178.600 7.200 ;
        RECT 172.600 6.100 173.000 6.500 ;
        RECT 169.400 4.800 169.800 5.200 ;
        RECT 179.000 5.100 179.400 5.500 ;
        RECT 179.800 4.800 180.200 5.200 ;
        RECT 189.400 6.800 189.800 7.200 ;
        RECT 187.800 5.900 188.200 6.300 ;
        RECT 183.800 4.800 184.200 5.200 ;
        RECT 185.400 5.100 185.800 5.500 ;
        RECT 198.200 6.800 198.600 7.200 ;
        RECT 211.000 8.800 211.400 9.200 ;
        RECT 200.600 6.800 201.000 7.200 ;
        RECT 220.600 8.800 221.000 9.200 ;
        RECT 206.200 6.800 206.600 7.200 ;
        RECT 204.600 5.900 205.000 6.300 ;
        RECT 198.200 4.800 198.600 5.200 ;
        RECT 202.200 5.100 202.600 5.500 ;
        RECT 227.000 8.800 227.400 9.200 ;
        RECT 215.800 6.800 216.200 7.200 ;
        RECT 216.600 5.800 217.000 6.200 ;
        RECT 211.800 5.100 212.200 5.500 ;
        RECT 224.600 6.800 225.000 7.200 ;
        RECT 244.600 8.800 245.000 9.200 ;
        RECT 224.600 4.800 225.000 5.200 ;
        RECT 235.000 6.800 235.400 7.200 ;
        RECT 229.400 6.100 229.800 6.500 ;
        RECT 243.000 6.800 243.400 7.200 ;
        RECT 235.800 5.100 236.200 5.500 ;
        RECT 248.600 8.800 249.000 9.200 ;
      LAYER metal2 ;
        RECT 11.000 236.800 11.400 237.200 ;
        RECT 7.000 235.800 7.400 236.200 ;
        RECT 8.600 236.100 9.000 236.200 ;
        RECT 9.400 236.100 9.800 236.200 ;
        RECT 8.600 235.800 9.800 236.100 ;
        RECT 7.000 235.200 7.300 235.800 ;
        RECT 2.200 234.800 2.600 235.200 ;
        RECT 7.000 234.800 7.400 235.200 ;
        RECT 9.400 234.800 9.800 235.200 ;
        RECT 2.200 234.200 2.500 234.800 ;
        RECT 2.200 233.800 2.600 234.200 ;
        RECT 4.600 234.100 5.000 234.200 ;
        RECT 5.400 234.100 5.800 234.200 ;
        RECT 4.600 233.800 5.800 234.100 ;
        RECT 6.200 233.800 6.600 234.200 ;
        RECT 6.200 233.200 6.500 233.800 ;
        RECT 0.600 232.800 1.000 233.200 ;
        RECT 6.200 232.800 6.600 233.200 ;
        RECT 0.600 229.200 0.900 232.800 ;
        RECT 3.800 232.100 4.200 232.200 ;
        RECT 3.800 231.800 4.900 232.100 ;
        RECT 0.600 228.800 1.000 229.200 ;
        RECT 3.000 223.100 3.400 228.900 ;
        RECT 4.600 226.200 4.900 231.800 ;
        RECT 4.600 225.800 5.000 226.200 ;
        RECT 0.600 222.100 1.000 222.200 ;
        RECT 1.400 222.100 1.800 222.200 ;
        RECT 0.600 221.800 1.800 222.100 ;
        RECT 7.000 221.200 7.300 234.800 ;
        RECT 9.400 234.200 9.700 234.800 ;
        RECT 11.000 234.200 11.300 236.800 ;
        RECT 9.400 233.800 9.800 234.200 ;
        RECT 11.000 233.800 11.400 234.200 ;
        RECT 7.800 223.100 8.200 228.900 ;
        RECT 8.600 226.800 9.000 227.200 ;
        RECT 8.600 224.200 8.900 226.800 ;
        RECT 9.400 225.100 9.800 227.900 ;
        RECT 11.000 227.200 11.300 233.800 ;
        RECT 14.200 232.100 14.600 237.900 ;
        RECT 16.600 235.100 17.000 235.200 ;
        RECT 17.400 235.100 17.800 235.200 ;
        RECT 16.600 234.800 17.800 235.100 ;
        RECT 17.400 232.800 17.800 233.200 ;
        RECT 17.400 227.200 17.700 232.800 ;
        RECT 19.000 232.100 19.400 237.900 ;
        RECT 20.600 233.100 21.000 235.900 ;
        RECT 29.400 235.800 29.800 236.200 ;
        RECT 31.000 236.100 31.400 236.200 ;
        RECT 31.800 236.100 32.200 236.200 ;
        RECT 31.000 235.800 32.200 236.100 ;
        RECT 29.400 235.200 29.700 235.800 ;
        RECT 28.600 235.100 29.000 235.200 ;
        RECT 29.400 235.100 29.800 235.200 ;
        RECT 28.600 234.800 29.800 235.100 ;
        RECT 31.800 234.800 32.200 235.200 ;
        RECT 31.800 234.200 32.100 234.800 ;
        RECT 21.400 233.800 21.800 234.200 ;
        RECT 22.200 233.800 22.600 234.200 ;
        RECT 27.800 234.100 28.200 234.200 ;
        RECT 28.600 234.100 29.000 234.200 ;
        RECT 27.800 233.800 29.000 234.100 ;
        RECT 31.800 233.800 32.200 234.200 ;
        RECT 33.400 233.800 33.800 234.200 ;
        RECT 11.000 226.800 11.400 227.200 ;
        RECT 16.600 226.800 17.000 227.200 ;
        RECT 17.400 226.800 17.800 227.200 ;
        RECT 19.800 226.800 20.200 227.200 ;
        RECT 16.600 224.200 16.900 226.800 ;
        RECT 18.200 226.100 18.600 226.200 ;
        RECT 19.000 226.100 19.400 226.200 ;
        RECT 18.200 225.800 19.400 226.100 ;
        RECT 19.800 225.200 20.100 226.800 ;
        RECT 20.600 225.800 21.000 226.200 ;
        RECT 20.600 225.200 20.900 225.800 ;
        RECT 19.800 224.800 20.200 225.200 ;
        RECT 20.600 224.800 21.000 225.200 ;
        RECT 8.600 223.800 9.000 224.200 ;
        RECT 16.600 223.800 17.000 224.200 ;
        RECT 13.400 222.800 13.800 223.200 ;
        RECT 11.000 221.800 11.400 222.200 ;
        RECT 7.000 220.800 7.400 221.200 ;
        RECT 0.600 219.100 1.000 219.200 ;
        RECT 1.400 219.100 1.800 219.200 ;
        RECT 0.600 218.800 1.800 219.100 ;
        RECT 3.000 212.100 3.400 217.900 ;
        RECT 7.000 215.800 7.400 216.200 ;
        RECT 7.000 215.100 7.300 215.800 ;
        RECT 7.000 214.700 7.400 215.100 ;
        RECT 7.800 212.100 8.200 217.900 ;
        RECT 11.000 217.200 11.300 221.800 ;
        RECT 8.600 216.800 9.000 217.200 ;
        RECT 11.000 216.800 11.400 217.200 ;
        RECT 8.600 214.200 8.900 216.800 ;
        RECT 13.400 216.200 13.700 222.800 ;
        RECT 19.000 220.800 19.400 221.200 ;
        RECT 15.000 218.800 15.400 219.200 ;
        RECT 14.200 216.800 14.600 217.200 ;
        RECT 8.600 213.800 9.000 214.200 ;
        RECT 9.400 213.100 9.800 215.900 ;
        RECT 11.800 215.800 12.200 216.200 ;
        RECT 13.400 215.800 13.800 216.200 ;
        RECT 11.800 215.200 12.100 215.800 ;
        RECT 13.400 215.200 13.700 215.800 ;
        RECT 10.200 215.100 10.600 215.200 ;
        RECT 11.000 215.100 11.400 215.200 ;
        RECT 10.200 214.800 11.400 215.100 ;
        RECT 11.800 214.800 12.200 215.200 ;
        RECT 13.400 214.800 13.800 215.200 ;
        RECT 10.200 213.800 10.600 214.200 ;
        RECT 10.200 211.200 10.500 213.800 ;
        RECT 10.200 210.800 10.600 211.200 ;
        RECT 0.600 209.100 1.000 209.200 ;
        RECT 1.400 209.100 1.800 209.200 ;
        RECT 0.600 208.800 1.800 209.100 ;
        RECT 3.000 203.100 3.400 208.900 ;
        RECT 6.200 206.100 6.600 206.200 ;
        RECT 7.000 206.100 7.400 206.300 ;
        RECT 6.200 205.900 7.400 206.100 ;
        RECT 6.200 205.800 7.300 205.900 ;
        RECT 7.800 203.100 8.200 208.900 ;
        RECT 8.600 207.800 9.000 208.200 ;
        RECT 8.600 207.200 8.900 207.800 ;
        RECT 8.600 206.800 9.000 207.200 ;
        RECT 9.400 205.100 9.800 207.900 ;
        RECT 10.200 207.200 10.500 210.800 ;
        RECT 10.200 206.800 10.600 207.200 ;
        RECT 0.600 191.800 1.000 192.200 ;
        RECT 3.000 192.100 3.400 197.900 ;
        RECT 6.200 196.800 6.600 197.200 ;
        RECT 4.600 194.800 5.000 195.200 ;
        RECT 0.600 187.200 0.900 191.800 ;
        RECT 0.600 187.100 1.000 187.200 ;
        RECT 1.400 187.100 1.800 187.200 ;
        RECT 0.600 186.800 1.800 187.100 ;
        RECT 3.800 187.100 4.200 187.200 ;
        RECT 4.600 187.100 4.900 194.800 ;
        RECT 3.800 186.800 4.900 187.100 ;
        RECT 6.200 187.200 6.500 196.800 ;
        RECT 7.800 192.100 8.200 197.900 ;
        RECT 10.200 197.200 10.500 206.800 ;
        RECT 11.000 205.800 11.400 206.200 ;
        RECT 11.800 206.100 12.200 206.200 ;
        RECT 12.600 206.100 13.000 206.200 ;
        RECT 11.800 205.800 13.000 206.100 ;
        RECT 11.000 205.200 11.300 205.800 ;
        RECT 11.000 204.800 11.400 205.200 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 13.400 204.200 13.700 204.800 ;
        RECT 13.400 203.800 13.800 204.200 ;
        RECT 10.200 196.800 10.600 197.200 ;
        RECT 8.600 194.800 9.000 195.200 ;
        RECT 8.600 189.200 8.900 194.800 ;
        RECT 9.400 193.100 9.800 195.900 ;
        RECT 10.200 193.100 10.600 195.900 ;
        RECT 11.800 192.100 12.200 197.900 ;
        RECT 12.600 194.700 13.000 195.100 ;
        RECT 12.600 194.200 12.900 194.700 ;
        RECT 14.200 194.200 14.500 216.800 ;
        RECT 15.000 214.200 15.300 218.800 ;
        RECT 16.600 216.800 17.000 217.200 ;
        RECT 15.000 213.800 15.400 214.200 ;
        RECT 15.800 213.100 16.200 215.900 ;
        RECT 16.600 214.200 16.900 216.800 ;
        RECT 16.600 213.800 17.000 214.200 ;
        RECT 17.400 212.100 17.800 217.900 ;
        RECT 18.200 214.700 18.600 215.100 ;
        RECT 15.800 210.800 16.200 211.200 ;
        RECT 15.000 207.800 15.400 208.200 ;
        RECT 15.000 207.200 15.300 207.800 ;
        RECT 15.800 207.200 16.100 210.800 ;
        RECT 18.200 209.200 18.500 214.700 ;
        RECT 18.200 208.800 18.600 209.200 ;
        RECT 15.000 206.800 15.400 207.200 ;
        RECT 15.800 206.800 16.200 207.200 ;
        RECT 19.000 206.200 19.300 220.800 ;
        RECT 20.600 215.200 20.900 224.800 ;
        RECT 20.600 214.800 21.000 215.200 ;
        RECT 21.400 213.200 21.700 233.800 ;
        RECT 22.200 233.200 22.500 233.800 ;
        RECT 28.600 233.200 28.900 233.800 ;
        RECT 22.200 232.800 22.600 233.200 ;
        RECT 28.600 232.800 29.000 233.200 ;
        RECT 33.400 232.200 33.700 233.800 ;
        RECT 34.200 233.100 34.600 235.900 ;
        RECT 27.000 231.800 27.400 232.200 ;
        RECT 33.400 231.800 33.800 232.200 ;
        RECT 35.800 232.100 36.200 237.900 ;
        RECT 36.600 235.800 37.000 236.200 ;
        RECT 36.600 235.100 36.900 235.800 ;
        RECT 36.600 234.700 37.000 235.100 ;
        RECT 37.400 233.800 37.800 234.200 ;
        RECT 36.600 232.800 37.000 233.200 ;
        RECT 22.200 228.800 22.600 229.200 ;
        RECT 22.200 227.200 22.500 228.800 ;
        RECT 22.200 226.800 22.600 227.200 ;
        RECT 23.000 225.100 23.400 227.900 ;
        RECT 24.600 223.100 25.000 228.900 ;
        RECT 25.400 225.900 25.800 226.300 ;
        RECT 25.400 225.200 25.700 225.900 ;
        RECT 25.400 224.800 25.800 225.200 ;
        RECT 25.400 221.800 25.800 222.200 ;
        RECT 21.400 212.800 21.800 213.200 ;
        RECT 20.600 211.800 21.000 212.200 ;
        RECT 22.200 212.100 22.600 217.900 ;
        RECT 25.400 215.200 25.700 221.800 ;
        RECT 25.400 214.800 25.800 215.200 ;
        RECT 23.800 212.100 24.200 212.200 ;
        RECT 24.600 212.100 25.000 212.200 ;
        RECT 23.800 211.800 25.000 212.100 ;
        RECT 20.600 207.200 20.900 211.800 ;
        RECT 24.600 210.200 24.900 211.800 ;
        RECT 24.600 209.800 25.000 210.200 ;
        RECT 20.600 206.800 21.000 207.200 ;
        RECT 22.200 206.800 22.600 207.200 ;
        RECT 22.200 206.200 22.500 206.800 ;
        RECT 16.600 206.100 17.000 206.200 ;
        RECT 17.400 206.100 17.800 206.200 ;
        RECT 16.600 205.800 17.800 206.100 ;
        RECT 19.000 205.800 19.400 206.200 ;
        RECT 21.400 205.800 21.800 206.200 ;
        RECT 22.200 205.800 22.600 206.200 ;
        RECT 19.000 205.200 19.300 205.800 ;
        RECT 19.000 204.800 19.400 205.200 ;
        RECT 19.000 199.200 19.300 204.800 ;
        RECT 19.000 198.800 19.400 199.200 ;
        RECT 12.600 193.800 13.000 194.200 ;
        RECT 14.200 193.800 14.600 194.200 ;
        RECT 16.600 192.100 17.000 197.900 ;
        RECT 21.400 192.200 21.700 205.800 ;
        RECT 23.800 201.800 24.200 202.200 ;
        RECT 19.000 191.800 19.400 192.200 ;
        RECT 20.600 191.800 21.000 192.200 ;
        RECT 21.400 191.800 21.800 192.200 ;
        RECT 8.600 188.800 9.000 189.200 ;
        RECT 6.200 186.800 6.600 187.200 ;
        RECT 11.000 186.800 11.400 187.200 ;
        RECT 11.800 186.800 12.200 187.200 ;
        RECT 11.000 186.200 11.300 186.800 ;
        RECT 11.800 186.200 12.100 186.800 ;
        RECT 19.000 186.200 19.300 191.800 ;
        RECT 20.600 187.200 20.900 191.800 ;
        RECT 20.600 186.800 21.000 187.200 ;
        RECT 22.200 187.100 22.600 187.200 ;
        RECT 23.000 187.100 23.400 187.200 ;
        RECT 22.200 186.800 23.400 187.100 ;
        RECT 4.600 185.800 5.000 186.200 ;
        RECT 7.000 186.100 7.400 186.200 ;
        RECT 7.800 186.100 8.200 186.200 ;
        RECT 7.000 185.800 8.200 186.100 ;
        RECT 9.400 185.800 9.800 186.200 ;
        RECT 11.000 185.800 11.400 186.200 ;
        RECT 11.800 185.800 12.200 186.200 ;
        RECT 14.200 186.100 14.600 186.200 ;
        RECT 15.000 186.100 15.400 186.200 ;
        RECT 14.200 185.800 15.400 186.100 ;
        RECT 15.800 185.800 16.200 186.200 ;
        RECT 19.000 185.800 19.400 186.200 ;
        RECT 4.600 185.200 4.900 185.800 ;
        RECT 9.400 185.200 9.700 185.800 ;
        RECT 2.200 185.100 2.600 185.200 ;
        RECT 3.000 185.100 3.400 185.200 ;
        RECT 2.200 184.800 3.400 185.100 ;
        RECT 4.600 184.800 5.000 185.200 ;
        RECT 9.400 184.800 9.800 185.200 ;
        RECT 13.400 184.800 13.800 185.200 ;
        RECT 0.600 178.100 1.000 178.200 ;
        RECT 1.400 178.100 1.800 178.200 ;
        RECT 0.600 177.800 1.800 178.100 ;
        RECT 3.000 172.100 3.400 177.900 ;
        RECT 4.600 165.200 4.900 184.800 ;
        RECT 9.400 180.200 9.700 184.800 ;
        RECT 13.400 184.200 13.700 184.800 ;
        RECT 15.800 184.200 16.100 185.800 ;
        RECT 13.400 183.800 13.800 184.200 ;
        RECT 15.800 183.800 16.200 184.200 ;
        RECT 17.400 181.800 17.800 182.200 ;
        RECT 9.400 179.800 9.800 180.200 ;
        RECT 7.000 175.800 7.400 176.200 ;
        RECT 7.000 175.100 7.300 175.800 ;
        RECT 7.000 174.700 7.400 175.100 ;
        RECT 7.800 172.100 8.200 177.900 ;
        RECT 15.000 177.800 15.400 178.200 ;
        RECT 8.600 176.800 9.000 177.200 ;
        RECT 8.600 174.200 8.900 176.800 ;
        RECT 8.600 173.800 9.000 174.200 ;
        RECT 9.400 173.100 9.800 175.900 ;
        RECT 10.200 175.800 10.600 176.200 ;
        RECT 13.400 176.100 13.800 176.200 ;
        RECT 14.200 176.100 14.600 176.200 ;
        RECT 13.400 175.800 14.600 176.100 ;
        RECT 10.200 174.200 10.500 175.800 ;
        RECT 11.000 175.100 11.400 175.200 ;
        RECT 11.800 175.100 12.200 175.200 ;
        RECT 11.000 174.800 12.200 175.100 ;
        RECT 15.000 174.200 15.300 177.800 ;
        RECT 17.400 177.200 17.700 181.800 ;
        RECT 17.400 176.800 17.800 177.200 ;
        RECT 17.400 176.100 17.800 176.200 ;
        RECT 18.200 176.100 18.600 176.200 ;
        RECT 17.400 175.800 18.600 176.100 ;
        RECT 18.200 175.100 18.600 175.200 ;
        RECT 19.000 175.100 19.400 175.200 ;
        RECT 18.200 174.800 19.400 175.100 ;
        RECT 10.200 173.800 10.600 174.200 ;
        RECT 12.600 173.800 13.000 174.200 ;
        RECT 13.400 174.100 13.800 174.200 ;
        RECT 14.200 174.100 14.600 174.200 ;
        RECT 13.400 173.800 14.600 174.100 ;
        RECT 15.000 173.800 15.400 174.200 ;
        RECT 15.800 173.800 16.200 174.200 ;
        RECT 18.200 173.800 18.600 174.200 ;
        RECT 12.600 173.200 12.900 173.800 ;
        RECT 12.600 172.800 13.000 173.200 ;
        RECT 4.600 164.800 5.000 165.200 ;
        RECT 7.800 165.100 8.200 167.900 ;
        RECT 9.400 163.100 9.800 168.900 ;
        RECT 11.800 168.800 12.200 169.200 ;
        RECT 15.800 169.100 16.100 173.800 ;
        RECT 18.200 173.200 18.500 173.800 ;
        RECT 18.200 172.800 18.600 173.200 ;
        RECT 17.400 171.800 17.800 172.200 ;
        RECT 16.600 169.100 17.000 169.200 ;
        RECT 11.800 167.200 12.100 168.800 ;
        RECT 11.800 166.800 12.200 167.200 ;
        RECT 11.000 166.100 11.400 166.200 ;
        RECT 11.800 166.100 12.200 166.200 ;
        RECT 11.000 165.800 12.200 166.100 ;
        RECT 14.200 163.100 14.600 168.900 ;
        RECT 15.800 168.800 17.000 169.100 ;
        RECT 15.000 166.800 15.400 167.200 ;
        RECT 1.400 161.800 1.800 162.200 ;
        RECT 0.600 153.100 1.000 155.900 ;
        RECT 1.400 154.200 1.700 161.800 ;
        RECT 1.400 153.800 1.800 154.200 ;
        RECT 0.600 145.100 1.000 147.900 ;
        RECT 1.400 147.200 1.700 153.800 ;
        RECT 2.200 152.100 2.600 157.900 ;
        RECT 4.600 155.100 5.000 155.200 ;
        RECT 5.400 155.100 5.800 155.200 ;
        RECT 4.600 154.800 5.800 155.100 ;
        RECT 7.000 152.100 7.400 157.900 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 10.200 154.200 10.500 156.800 ;
        RECT 11.000 156.100 11.400 156.200 ;
        RECT 11.800 156.100 12.200 156.200 ;
        RECT 11.000 155.800 12.200 156.100 ;
        RECT 14.200 155.800 14.600 156.200 ;
        RECT 14.200 155.200 14.500 155.800 ;
        RECT 12.600 155.100 13.000 155.200 ;
        RECT 13.400 155.100 13.800 155.200 ;
        RECT 12.600 154.800 13.800 155.100 ;
        RECT 14.200 154.800 14.600 155.200 ;
        RECT 15.000 154.200 15.300 166.800 ;
        RECT 17.400 165.200 17.700 171.800 ;
        RECT 20.600 169.200 20.900 186.800 ;
        RECT 23.800 186.200 24.100 201.800 ;
        RECT 27.000 199.200 27.300 231.800 ;
        RECT 31.000 229.100 31.400 229.200 ;
        RECT 31.800 229.100 32.200 229.200 ;
        RECT 28.600 225.800 29.000 226.200 ;
        RECT 28.600 224.200 28.900 225.800 ;
        RECT 28.600 223.800 29.000 224.200 ;
        RECT 29.400 223.100 29.800 228.900 ;
        RECT 31.000 228.800 32.200 229.100 ;
        RECT 33.400 228.800 33.800 229.200 ;
        RECT 33.400 226.200 33.700 228.800 ;
        RECT 36.600 227.200 36.900 232.800 ;
        RECT 35.800 226.800 36.200 227.200 ;
        RECT 36.600 226.800 37.000 227.200 ;
        RECT 35.800 226.200 36.100 226.800 ;
        RECT 32.600 225.800 33.000 226.200 ;
        RECT 33.400 225.800 33.800 226.200 ;
        RECT 35.000 225.800 35.400 226.200 ;
        RECT 35.800 225.800 36.200 226.200 ;
        RECT 32.600 222.200 32.900 225.800 ;
        RECT 35.000 225.200 35.300 225.800 ;
        RECT 35.000 224.800 35.400 225.200 ;
        RECT 37.400 224.200 37.700 233.800 ;
        RECT 40.600 232.100 41.000 237.900 ;
        RECT 45.400 233.800 45.800 234.200 ;
        RECT 45.400 232.200 45.700 233.800 ;
        RECT 42.200 232.100 42.600 232.200 ;
        RECT 43.000 232.100 43.400 232.200 ;
        RECT 42.200 231.800 43.400 232.100 ;
        RECT 45.400 231.800 45.800 232.200 ;
        RECT 47.800 232.100 48.200 237.900 ;
        RECT 51.000 235.100 51.400 235.200 ;
        RECT 51.000 234.800 52.200 235.100 ;
        RECT 51.800 234.700 52.200 234.800 ;
        RECT 52.600 232.100 53.000 237.900 ;
        RECT 55.000 237.100 55.400 237.200 ;
        RECT 55.800 237.100 56.200 237.200 ;
        RECT 55.000 236.800 56.200 237.100 ;
        RECT 57.400 236.800 57.800 237.200 ;
        RECT 57.400 236.200 57.700 236.800 ;
        RECT 55.800 236.100 56.200 236.200 ;
        RECT 56.600 236.100 57.000 236.200 ;
        RECT 53.400 233.800 53.800 234.200 ;
        RECT 53.400 233.200 53.700 233.800 ;
        RECT 53.400 232.800 53.800 233.200 ;
        RECT 54.200 233.100 54.600 235.900 ;
        RECT 55.800 235.800 57.000 236.100 ;
        RECT 57.400 235.800 57.800 236.200 ;
        RECT 59.000 235.800 59.400 236.200 ;
        RECT 59.000 235.200 59.300 235.800 ;
        RECT 55.800 235.100 56.200 235.200 ;
        RECT 56.600 235.100 57.000 235.200 ;
        RECT 55.800 234.800 57.000 235.100 ;
        RECT 59.000 234.800 59.400 235.200 ;
        RECT 59.800 234.800 60.200 235.200 ;
        RECT 59.800 234.200 60.100 234.800 ;
        RECT 55.000 234.100 55.400 234.200 ;
        RECT 55.800 234.100 56.200 234.200 ;
        RECT 55.000 233.800 56.200 234.100 ;
        RECT 58.200 233.800 58.600 234.200 ;
        RECT 59.800 233.800 60.200 234.200 ;
        RECT 42.200 228.800 42.600 229.200 ;
        RECT 51.000 229.100 51.400 229.200 ;
        RECT 51.800 229.100 52.200 229.200 ;
        RECT 42.200 227.200 42.500 228.800 ;
        RECT 40.600 226.800 41.000 227.200 ;
        RECT 42.200 226.800 42.600 227.200 ;
        RECT 40.600 226.200 40.900 226.800 ;
        RECT 38.200 225.800 38.600 226.200 ;
        RECT 40.600 225.800 41.000 226.200 ;
        RECT 38.200 225.200 38.500 225.800 ;
        RECT 38.200 224.800 38.600 225.200 ;
        RECT 40.600 225.100 41.000 225.200 ;
        RECT 41.400 225.100 41.800 225.200 ;
        RECT 43.000 225.100 43.400 227.900 ;
        RECT 43.800 226.800 44.200 227.200 ;
        RECT 40.600 224.800 41.800 225.100 ;
        RECT 37.400 223.800 37.800 224.200 ;
        RECT 32.600 221.800 33.000 222.200 ;
        RECT 37.400 217.200 37.700 223.800 ;
        RECT 35.000 216.800 35.400 217.200 ;
        RECT 35.800 216.800 36.200 217.200 ;
        RECT 37.400 216.800 37.800 217.200 ;
        RECT 28.600 215.800 29.000 216.200 ;
        RECT 31.800 215.800 32.200 216.200 ;
        RECT 28.600 215.200 28.900 215.800 ;
        RECT 28.600 214.800 29.000 215.200 ;
        RECT 29.400 214.800 29.800 215.200 ;
        RECT 30.200 214.800 30.600 215.200 ;
        RECT 27.800 211.800 28.200 212.200 ;
        RECT 27.800 209.200 28.100 211.800 ;
        RECT 27.800 208.800 28.200 209.200 ;
        RECT 27.800 207.800 28.200 208.200 ;
        RECT 27.800 207.200 28.100 207.800 ;
        RECT 27.800 206.800 28.200 207.200 ;
        RECT 27.800 205.800 28.200 206.200 ;
        RECT 27.000 198.800 27.400 199.200 ;
        RECT 27.000 196.800 27.400 197.200 ;
        RECT 27.000 194.200 27.300 196.800 ;
        RECT 27.000 193.800 27.400 194.200 ;
        RECT 27.800 186.200 28.100 205.800 ;
        RECT 28.600 203.100 29.000 208.900 ;
        RECT 29.400 207.200 29.700 214.800 ;
        RECT 30.200 214.200 30.500 214.800 ;
        RECT 30.200 213.800 30.600 214.200 ;
        RECT 31.800 213.200 32.100 215.800 ;
        RECT 35.000 215.200 35.300 216.800 ;
        RECT 35.800 216.200 36.100 216.800 ;
        RECT 35.800 215.800 36.200 216.200 ;
        RECT 35.000 214.800 35.400 215.200 ;
        RECT 34.200 213.800 34.600 214.200 ;
        RECT 31.800 212.800 32.200 213.200 ;
        RECT 32.600 212.100 33.000 212.200 ;
        RECT 33.400 212.100 33.800 212.200 ;
        RECT 32.600 211.800 33.800 212.100 ;
        RECT 29.400 206.800 29.800 207.200 ;
        RECT 29.400 205.800 29.800 206.200 ;
        RECT 32.600 205.900 33.000 206.300 ;
        RECT 28.600 195.800 29.000 196.200 ;
        RECT 28.600 195.200 28.900 195.800 ;
        RECT 28.600 194.800 29.000 195.200 ;
        RECT 29.400 187.200 29.700 205.800 ;
        RECT 32.600 205.200 32.900 205.900 ;
        RECT 32.600 204.800 33.000 205.200 ;
        RECT 33.400 203.100 33.800 208.900 ;
        RECT 34.200 202.200 34.500 213.800 ;
        RECT 38.200 212.100 38.600 217.900 ;
        RECT 39.800 214.800 40.200 215.200 ;
        RECT 41.400 214.800 41.800 215.200 ;
        RECT 35.000 205.100 35.400 207.900 ;
        RECT 35.800 207.800 36.200 208.200 ;
        RECT 35.800 207.200 36.100 207.800 ;
        RECT 35.800 206.800 36.200 207.200 ;
        RECT 37.400 205.800 37.800 206.200 ;
        RECT 39.000 205.800 39.400 206.200 ;
        RECT 37.400 205.200 37.700 205.800 ;
        RECT 39.000 205.200 39.300 205.800 ;
        RECT 37.400 204.800 37.800 205.200 ;
        RECT 39.000 204.800 39.400 205.200 ;
        RECT 34.200 201.800 34.600 202.200 ;
        RECT 31.000 196.100 31.400 196.200 ;
        RECT 31.800 196.100 32.200 196.200 ;
        RECT 31.000 195.800 32.200 196.100 ;
        RECT 31.000 194.800 31.400 195.200 ;
        RECT 29.400 186.800 29.800 187.200 ;
        RECT 23.800 185.800 24.200 186.200 ;
        RECT 24.600 185.800 25.000 186.200 ;
        RECT 27.000 185.800 27.400 186.200 ;
        RECT 27.800 185.800 28.200 186.200 ;
        RECT 29.400 185.800 29.800 186.200 ;
        RECT 24.600 178.200 24.900 185.800 ;
        RECT 25.400 181.800 25.800 182.200 ;
        RECT 25.400 179.200 25.700 181.800 ;
        RECT 25.400 178.800 25.800 179.200 ;
        RECT 24.600 177.800 25.000 178.200 ;
        RECT 24.600 176.800 25.000 177.200 ;
        RECT 21.400 175.800 21.800 176.200 ;
        RECT 23.000 175.800 23.400 176.200 ;
        RECT 21.400 175.200 21.700 175.800 ;
        RECT 21.400 174.800 21.800 175.200 ;
        RECT 23.000 174.200 23.300 175.800 ;
        RECT 21.400 174.100 21.800 174.200 ;
        RECT 22.200 174.100 22.600 174.200 ;
        RECT 21.400 173.800 22.600 174.100 ;
        RECT 23.000 173.800 23.400 174.200 ;
        RECT 23.800 173.100 24.200 175.900 ;
        RECT 24.600 174.200 24.900 176.800 ;
        RECT 24.600 173.800 25.000 174.200 ;
        RECT 23.800 170.800 24.200 171.200 ;
        RECT 20.600 168.800 21.000 169.200 ;
        RECT 19.000 167.100 19.400 167.200 ;
        RECT 19.800 167.100 20.200 167.200 ;
        RECT 19.000 166.800 20.200 167.100 ;
        RECT 19.000 166.100 19.400 166.200 ;
        RECT 19.800 166.100 20.200 166.200 ;
        RECT 19.000 165.800 20.200 166.100 ;
        RECT 17.400 164.800 17.800 165.200 ;
        RECT 20.600 165.100 21.000 167.900 ;
        RECT 19.000 163.800 19.400 164.200 ;
        RECT 19.000 163.200 19.300 163.800 ;
        RECT 19.000 162.800 19.400 163.200 ;
        RECT 22.200 163.100 22.600 168.900 ;
        RECT 23.000 168.800 23.400 169.200 ;
        RECT 23.000 168.200 23.300 168.800 ;
        RECT 23.000 167.800 23.400 168.200 ;
        RECT 16.600 161.800 17.000 162.200 ;
        RECT 16.600 155.200 16.900 161.800 ;
        RECT 23.800 156.200 24.100 170.800 ;
        RECT 24.600 168.200 24.900 173.800 ;
        RECT 25.400 172.100 25.800 177.900 ;
        RECT 27.000 176.200 27.300 185.800 ;
        RECT 27.000 175.800 27.400 176.200 ;
        RECT 26.200 174.700 26.600 175.100 ;
        RECT 26.200 174.200 26.500 174.700 ;
        RECT 26.200 173.800 26.600 174.200 ;
        RECT 24.600 167.800 25.000 168.200 ;
        RECT 25.400 166.800 25.800 167.200 ;
        RECT 25.400 166.200 25.700 166.800 ;
        RECT 25.400 165.800 25.800 166.200 ;
        RECT 27.000 163.100 27.400 168.900 ;
        RECT 27.800 159.200 28.100 185.800 ;
        RECT 29.400 185.200 29.700 185.800 ;
        RECT 29.400 184.800 29.800 185.200 ;
        RECT 30.200 181.800 30.600 182.200 ;
        RECT 30.200 179.200 30.500 181.800 ;
        RECT 30.200 178.800 30.600 179.200 ;
        RECT 28.600 175.100 29.000 175.200 ;
        RECT 29.400 175.100 29.800 175.200 ;
        RECT 28.600 174.800 29.800 175.100 ;
        RECT 30.200 172.100 30.600 177.900 ;
        RECT 31.000 177.200 31.300 194.800 ;
        RECT 31.800 193.800 32.200 194.200 ;
        RECT 31.800 193.200 32.100 193.800 ;
        RECT 31.800 192.800 32.200 193.200 ;
        RECT 32.600 193.100 33.000 195.900 ;
        RECT 33.400 193.800 33.800 194.200 ;
        RECT 33.400 187.200 33.700 193.800 ;
        RECT 34.200 192.100 34.600 197.900 ;
        RECT 35.000 195.800 35.400 196.200 ;
        RECT 35.000 195.100 35.300 195.800 ;
        RECT 35.000 194.700 35.400 195.100 ;
        RECT 34.200 188.800 34.600 189.200 ;
        RECT 34.200 188.200 34.500 188.800 ;
        RECT 34.200 187.800 34.600 188.200 ;
        RECT 33.400 186.800 33.800 187.200 ;
        RECT 31.800 185.800 32.200 186.200 ;
        RECT 32.600 186.100 33.000 186.200 ;
        RECT 33.400 186.100 33.800 186.200 ;
        RECT 32.600 185.800 33.800 186.100 ;
        RECT 31.800 185.200 32.100 185.800 ;
        RECT 31.800 184.800 32.200 185.200 ;
        RECT 31.000 176.800 31.400 177.200 ;
        RECT 32.600 176.800 33.000 177.200 ;
        RECT 32.600 176.200 32.900 176.800 ;
        RECT 32.600 175.800 33.000 176.200 ;
        RECT 35.000 172.800 35.400 173.200 ;
        RECT 33.400 171.800 33.800 172.200 ;
        RECT 29.400 168.800 29.800 169.200 ;
        RECT 29.400 168.100 29.700 168.800 ;
        RECT 30.200 168.100 30.600 168.200 ;
        RECT 29.400 167.800 30.600 168.100 ;
        RECT 30.200 167.200 30.500 167.800 ;
        RECT 33.400 167.200 33.700 171.800 ;
        RECT 35.000 169.200 35.300 172.800 ;
        RECT 35.800 172.100 36.200 177.900 ;
        RECT 36.600 174.800 37.000 175.200 ;
        RECT 36.600 174.200 36.900 174.800 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 37.400 171.200 37.700 204.800 ;
        RECT 39.000 192.100 39.400 197.900 ;
        RECT 39.800 197.200 40.100 214.800 ;
        RECT 40.600 213.800 41.000 214.200 ;
        RECT 40.600 211.200 40.900 213.800 ;
        RECT 41.400 212.200 41.700 214.800 ;
        RECT 41.400 211.800 41.800 212.200 ;
        RECT 43.000 212.100 43.400 217.900 ;
        RECT 43.800 216.200 44.100 226.800 ;
        RECT 44.600 223.100 45.000 228.900 ;
        RECT 45.400 225.900 45.800 226.300 ;
        RECT 45.400 225.200 45.700 225.900 ;
        RECT 45.400 224.800 45.800 225.200 ;
        RECT 49.400 223.100 49.800 228.900 ;
        RECT 51.000 228.800 52.200 229.100 ;
        RECT 55.000 228.800 55.400 229.200 ;
        RECT 55.000 226.200 55.300 228.800 ;
        RECT 56.600 227.100 57.000 227.200 ;
        RECT 57.400 227.100 57.800 227.200 ;
        RECT 56.600 226.800 57.800 227.100 ;
        RECT 58.200 226.200 58.500 233.800 ;
        RECT 60.600 233.100 61.000 235.900 ;
        RECT 62.200 232.100 62.600 237.900 ;
        RECT 63.800 236.800 64.200 237.200 ;
        RECT 63.800 235.200 64.100 236.800 ;
        RECT 63.800 234.800 64.200 235.200 ;
        RECT 63.000 232.800 63.400 233.200 ;
        RECT 62.200 226.800 62.600 227.200 ;
        RECT 62.200 226.200 62.500 226.800 ;
        RECT 63.000 226.200 63.300 232.800 ;
        RECT 64.600 231.800 65.000 232.200 ;
        RECT 67.000 232.100 67.400 237.900 ;
        RECT 74.200 237.800 74.600 238.200 ;
        RECT 74.200 237.200 74.500 237.800 ;
        RECT 70.200 236.800 70.600 237.200 ;
        RECT 74.200 236.800 74.600 237.200 ;
        RECT 70.200 234.200 70.500 236.800 ;
        RECT 71.800 235.800 72.200 236.200 ;
        RECT 71.800 235.200 72.100 235.800 ;
        RECT 71.800 234.800 72.200 235.200 ;
        RECT 74.200 235.100 74.600 235.200 ;
        RECT 75.000 235.100 75.400 235.200 ;
        RECT 74.200 234.800 75.400 235.100 ;
        RECT 70.200 233.800 70.600 234.200 ;
        RECT 75.000 234.100 75.400 234.200 ;
        RECT 75.800 234.100 76.200 234.200 ;
        RECT 75.000 233.800 76.200 234.100 ;
        RECT 76.600 233.800 77.000 234.200 ;
        RECT 70.200 232.200 70.500 233.800 ;
        RECT 70.200 231.800 70.600 232.200 ;
        RECT 75.800 231.800 76.200 232.200 ;
        RECT 64.600 226.200 64.900 231.800 ;
        RECT 75.800 231.200 76.100 231.800 ;
        RECT 75.800 230.800 76.200 231.200 ;
        RECT 75.800 228.800 76.200 229.200 ;
        RECT 75.800 228.200 76.100 228.800 ;
        RECT 67.800 227.800 68.200 228.200 ;
        RECT 75.800 227.800 76.200 228.200 ;
        RECT 67.800 226.200 68.100 227.800 ;
        RECT 68.600 226.800 69.000 227.200 ;
        RECT 54.200 225.800 54.600 226.200 ;
        RECT 55.000 225.800 55.400 226.200 ;
        RECT 58.200 225.800 58.600 226.200 ;
        RECT 59.000 225.800 59.400 226.200 ;
        RECT 59.800 225.800 60.200 226.200 ;
        RECT 62.200 225.800 62.600 226.200 ;
        RECT 63.000 225.800 63.400 226.200 ;
        RECT 63.800 225.800 64.200 226.200 ;
        RECT 64.600 225.800 65.000 226.200 ;
        RECT 67.800 225.800 68.200 226.200 ;
        RECT 43.800 215.800 44.200 216.200 ;
        RECT 43.800 214.200 44.100 215.800 ;
        RECT 43.800 213.800 44.200 214.200 ;
        RECT 43.800 212.800 44.200 213.200 ;
        RECT 44.600 213.100 45.000 215.900 ;
        RECT 40.600 210.800 41.000 211.200 ;
        RECT 40.600 207.200 40.900 210.800 ;
        RECT 40.600 206.800 41.000 207.200 ;
        RECT 40.600 205.800 41.000 206.200 ;
        RECT 40.600 205.200 40.900 205.800 ;
        RECT 40.600 204.800 41.000 205.200 ;
        RECT 41.400 205.100 41.800 207.900 ;
        RECT 43.000 203.100 43.400 208.900 ;
        RECT 43.800 207.200 44.100 212.800 ;
        RECT 49.400 211.800 49.800 212.200 ;
        RECT 51.800 212.100 52.200 217.900 ;
        RECT 52.600 214.800 53.000 215.200 ;
        RECT 52.600 213.200 52.900 214.800 ;
        RECT 52.600 212.800 53.000 213.200 ;
        RECT 43.800 206.800 44.200 207.200 ;
        RECT 39.800 196.800 40.200 197.200 ;
        RECT 40.600 197.100 41.000 197.200 ;
        RECT 41.400 197.100 41.800 197.200 ;
        RECT 40.600 196.800 41.800 197.100 ;
        RECT 43.000 193.800 43.400 194.200 ;
        RECT 43.000 192.200 43.300 193.800 ;
        RECT 43.000 191.800 43.400 192.200 ;
        RECT 40.600 188.800 41.000 189.200 ;
        RECT 40.600 188.200 40.900 188.800 ;
        RECT 40.600 187.800 41.000 188.200 ;
        RECT 39.000 187.100 39.400 187.200 ;
        RECT 39.800 187.100 40.200 187.200 ;
        RECT 39.000 186.800 40.200 187.100 ;
        RECT 43.000 186.200 43.300 191.800 ;
        RECT 43.800 188.200 44.100 206.800 ;
        RECT 44.600 205.800 45.000 206.200 ;
        RECT 44.600 205.200 44.900 205.800 ;
        RECT 44.600 204.800 45.000 205.200 ;
        RECT 47.800 203.100 48.200 208.900 ;
        RECT 49.400 206.200 49.700 211.800 ;
        RECT 54.200 211.200 54.500 225.800 ;
        RECT 59.000 224.200 59.300 225.800 ;
        RECT 59.800 225.200 60.100 225.800 ;
        RECT 59.800 224.800 60.200 225.200 ;
        RECT 59.000 223.800 59.400 224.200 ;
        RECT 63.800 222.200 64.100 225.800 ;
        RECT 61.400 221.800 61.800 222.200 ;
        RECT 63.800 221.800 64.200 222.200 ;
        RECT 66.200 221.800 66.600 222.200 ;
        RECT 61.400 220.200 61.700 221.800 ;
        RECT 66.200 220.200 66.500 221.800 ;
        RECT 68.600 221.200 68.900 226.800 ;
        RECT 74.200 226.100 74.600 226.200 ;
        RECT 75.000 226.100 75.400 226.200 ;
        RECT 74.200 225.800 75.400 226.100 ;
        RECT 67.000 220.800 67.400 221.200 ;
        RECT 68.600 220.800 69.000 221.200 ;
        RECT 61.400 219.800 61.800 220.200 ;
        RECT 63.800 219.800 64.200 220.200 ;
        RECT 66.200 219.800 66.600 220.200 ;
        RECT 55.800 214.700 56.200 215.100 ;
        RECT 54.200 210.800 54.600 211.200 ;
        RECT 55.800 211.100 56.100 214.700 ;
        RECT 56.600 212.100 57.000 217.900 ;
        RECT 58.200 213.100 58.600 215.900 ;
        RECT 59.000 211.800 59.400 212.200 ;
        RECT 61.400 212.100 61.800 217.900 ;
        RECT 62.200 215.800 62.600 216.200 ;
        RECT 62.200 215.200 62.500 215.800 ;
        RECT 62.200 214.800 62.600 215.200 ;
        RECT 55.800 210.800 56.900 211.100 ;
        RECT 56.600 209.200 56.900 210.800 ;
        RECT 58.200 209.800 58.600 210.200 ;
        RECT 54.200 208.800 54.600 209.200 ;
        RECT 56.600 208.800 57.000 209.200 ;
        RECT 57.400 208.800 57.800 209.200 ;
        RECT 49.400 205.800 49.800 206.200 ;
        RECT 51.000 205.800 51.400 206.200 ;
        RECT 51.000 205.200 51.300 205.800 ;
        RECT 51.000 204.800 51.400 205.200 ;
        RECT 50.200 201.800 50.600 202.200 ;
        RECT 44.600 198.800 45.000 199.200 ;
        RECT 44.600 195.200 44.900 198.800 ;
        RECT 50.200 198.200 50.500 201.800 ;
        RECT 50.200 197.800 50.600 198.200 ;
        RECT 46.200 196.800 46.600 197.200 ;
        RECT 46.200 195.200 46.500 196.800 ;
        RECT 51.000 195.800 51.400 196.200 ;
        RECT 52.600 195.800 53.000 196.200 ;
        RECT 44.600 194.800 45.000 195.200 ;
        RECT 45.400 194.800 45.800 195.200 ;
        RECT 46.200 194.800 46.600 195.200 ;
        RECT 48.600 194.800 49.000 195.200 ;
        RECT 45.400 194.200 45.700 194.800 ;
        RECT 45.400 193.800 45.800 194.200 ;
        RECT 48.600 189.200 48.900 194.800 ;
        RECT 51.000 194.200 51.300 195.800 ;
        RECT 52.600 195.200 52.900 195.800 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 52.600 194.800 53.000 195.200 ;
        RECT 54.200 195.100 54.500 208.800 ;
        RECT 57.400 208.200 57.700 208.800 ;
        RECT 57.400 207.800 57.800 208.200 ;
        RECT 55.800 206.800 56.200 207.200 ;
        RECT 55.800 204.200 56.100 206.800 ;
        RECT 58.200 206.200 58.500 209.800 ;
        RECT 59.000 206.200 59.300 211.800 ;
        RECT 62.200 206.800 62.600 207.200 ;
        RECT 63.000 206.800 63.400 207.200 ;
        RECT 62.200 206.200 62.500 206.800 ;
        RECT 63.000 206.200 63.300 206.800 ;
        RECT 58.200 205.800 58.600 206.200 ;
        RECT 59.000 205.800 59.400 206.200 ;
        RECT 60.600 206.100 61.000 206.200 ;
        RECT 61.400 206.100 61.800 206.200 ;
        RECT 60.600 205.800 61.800 206.100 ;
        RECT 62.200 205.800 62.600 206.200 ;
        RECT 63.000 205.800 63.400 206.200 ;
        RECT 59.000 204.800 59.400 205.200 ;
        RECT 55.800 203.800 56.200 204.200 ;
        RECT 55.800 197.800 56.200 198.200 ;
        RECT 55.000 195.100 55.400 195.200 ;
        RECT 54.200 194.800 55.400 195.100 ;
        RECT 51.800 194.200 52.100 194.800 ;
        RECT 55.800 194.200 56.100 197.800 ;
        RECT 58.200 195.800 58.600 196.200 ;
        RECT 58.200 195.200 58.500 195.800 ;
        RECT 58.200 194.800 58.600 195.200 ;
        RECT 59.000 194.200 59.300 204.800 ;
        RECT 63.000 203.800 63.400 204.200 ;
        RECT 60.600 201.800 61.000 202.200 ;
        RECT 60.600 201.200 60.900 201.800 ;
        RECT 60.600 200.800 61.000 201.200 ;
        RECT 63.000 199.200 63.300 203.800 ;
        RECT 63.000 198.800 63.400 199.200 ;
        RECT 60.600 194.800 61.000 195.200 ;
        RECT 62.200 195.100 62.600 195.200 ;
        RECT 63.000 195.100 63.400 195.200 ;
        RECT 62.200 194.800 63.400 195.100 ;
        RECT 63.800 195.100 64.100 219.800 ;
        RECT 65.400 216.800 65.800 217.200 ;
        RECT 64.600 215.800 65.000 216.200 ;
        RECT 64.600 209.200 64.900 215.800 ;
        RECT 65.400 215.100 65.700 216.800 ;
        RECT 65.400 214.700 65.800 215.100 ;
        RECT 66.200 212.100 66.600 217.900 ;
        RECT 67.000 214.200 67.300 220.800 ;
        RECT 70.200 217.800 70.600 218.200 ;
        RECT 70.200 217.200 70.500 217.800 ;
        RECT 70.200 216.800 70.600 217.200 ;
        RECT 68.600 216.100 69.000 216.200 ;
        RECT 69.400 216.100 69.800 216.200 ;
        RECT 67.000 213.800 67.400 214.200 ;
        RECT 66.200 210.800 66.600 211.200 ;
        RECT 64.600 208.800 65.000 209.200 ;
        RECT 65.400 208.800 65.800 209.200 ;
        RECT 65.400 208.200 65.700 208.800 ;
        RECT 65.400 207.800 65.800 208.200 ;
        RECT 64.600 204.800 65.000 205.200 ;
        RECT 64.600 202.200 64.900 204.800 ;
        RECT 64.600 201.800 65.000 202.200 ;
        RECT 64.600 196.100 65.000 196.200 ;
        RECT 65.400 196.100 65.800 196.200 ;
        RECT 64.600 195.800 65.800 196.100 ;
        RECT 64.600 195.100 65.000 195.200 ;
        RECT 63.800 194.800 65.000 195.100 ;
        RECT 60.600 194.200 60.900 194.800 ;
        RECT 51.000 193.800 51.400 194.200 ;
        RECT 51.800 193.800 52.200 194.200 ;
        RECT 55.800 193.800 56.200 194.200 ;
        RECT 59.000 193.800 59.400 194.200 ;
        RECT 60.600 193.800 61.000 194.200 ;
        RECT 61.400 193.800 61.800 194.200 ;
        RECT 62.200 193.800 62.600 194.200 ;
        RECT 64.600 194.100 65.000 194.200 ;
        RECT 65.400 194.100 65.800 194.200 ;
        RECT 64.600 193.800 65.800 194.100 ;
        RECT 54.200 191.800 54.600 192.200 ;
        RECT 54.200 189.200 54.500 191.800 ;
        RECT 47.000 189.100 47.400 189.200 ;
        RECT 47.800 189.100 48.200 189.200 ;
        RECT 47.000 188.800 48.200 189.100 ;
        RECT 48.600 188.800 49.000 189.200 ;
        RECT 43.800 187.800 44.200 188.200 ;
        RECT 44.600 186.800 45.000 187.200 ;
        RECT 45.400 186.800 45.800 187.200 ;
        RECT 42.200 185.800 42.600 186.200 ;
        RECT 43.000 185.800 43.400 186.200 ;
        RECT 43.800 185.800 44.200 186.200 ;
        RECT 42.200 182.200 42.500 185.800 ;
        RECT 43.800 185.200 44.100 185.800 ;
        RECT 43.800 184.800 44.200 185.200 ;
        RECT 44.600 182.200 44.900 186.800 ;
        RECT 45.400 186.200 45.700 186.800 ;
        RECT 45.400 185.800 45.800 186.200 ;
        RECT 42.200 181.800 42.600 182.200 ;
        RECT 44.600 181.800 45.000 182.200 ;
        RECT 44.600 179.800 45.000 180.200 ;
        RECT 39.800 175.800 40.200 176.200 ;
        RECT 39.800 175.100 40.100 175.800 ;
        RECT 39.800 174.700 40.200 175.100 ;
        RECT 40.600 172.100 41.000 177.900 ;
        RECT 41.400 173.800 41.800 174.200 ;
        RECT 37.400 170.800 37.800 171.200 ;
        RECT 35.000 168.800 35.400 169.200 ;
        RECT 35.000 167.200 35.300 168.800 ;
        RECT 41.400 168.200 41.700 173.800 ;
        RECT 42.200 173.100 42.600 175.900 ;
        RECT 43.000 175.800 43.400 176.200 ;
        RECT 43.000 172.100 43.300 175.800 ;
        RECT 44.600 175.200 44.900 179.800 ;
        RECT 43.800 174.800 44.200 175.200 ;
        RECT 44.600 174.800 45.000 175.200 ;
        RECT 43.800 174.200 44.100 174.800 ;
        RECT 43.800 173.800 44.200 174.200 ;
        RECT 42.200 171.800 43.300 172.100 ;
        RECT 42.200 169.200 42.500 171.800 ;
        RECT 42.200 168.800 42.600 169.200 ;
        RECT 35.800 167.800 36.200 168.200 ;
        RECT 41.400 167.800 41.800 168.200 ;
        RECT 30.200 166.800 30.600 167.200 ;
        RECT 31.800 167.100 32.200 167.200 ;
        RECT 32.600 167.100 33.000 167.200 ;
        RECT 31.800 166.800 33.000 167.100 ;
        RECT 33.400 166.800 33.800 167.200 ;
        RECT 35.000 166.800 35.400 167.200 ;
        RECT 35.800 166.200 36.100 167.800 ;
        RECT 39.000 166.800 39.400 167.200 ;
        RECT 40.600 166.800 41.000 167.200 ;
        RECT 39.000 166.200 39.300 166.800 ;
        RECT 40.600 166.200 40.900 166.800 ;
        RECT 34.200 165.800 34.600 166.200 ;
        RECT 35.800 165.800 36.200 166.200 ;
        RECT 39.000 165.800 39.400 166.200 ;
        RECT 39.800 165.800 40.200 166.200 ;
        RECT 40.600 165.800 41.000 166.200 ;
        RECT 43.800 165.800 44.200 166.200 ;
        RECT 34.200 165.200 34.500 165.800 ;
        RECT 31.800 164.800 32.200 165.200 ;
        RECT 34.200 164.800 34.600 165.200 ;
        RECT 27.800 158.800 28.200 159.200 ;
        RECT 26.200 156.800 26.600 157.200 ;
        RECT 19.800 155.800 20.200 156.200 ;
        RECT 23.800 155.800 24.200 156.200 ;
        RECT 19.800 155.200 20.100 155.800 ;
        RECT 23.800 155.200 24.100 155.800 ;
        RECT 15.800 154.800 16.200 155.200 ;
        RECT 16.600 154.800 17.000 155.200 ;
        RECT 18.200 155.100 18.600 155.200 ;
        RECT 19.000 155.100 19.400 155.200 ;
        RECT 18.200 154.800 19.400 155.100 ;
        RECT 19.800 154.800 20.200 155.200 ;
        RECT 20.600 154.800 21.000 155.200 ;
        RECT 21.400 155.100 21.800 155.200 ;
        RECT 22.200 155.100 22.600 155.200 ;
        RECT 21.400 154.800 22.600 155.100 ;
        RECT 23.800 154.800 24.200 155.200 ;
        RECT 15.800 154.200 16.100 154.800 ;
        RECT 20.600 154.200 20.900 154.800 ;
        RECT 10.200 154.100 10.600 154.200 ;
        RECT 11.000 154.100 11.400 154.200 ;
        RECT 10.200 153.800 11.400 154.100 ;
        RECT 15.000 153.800 15.400 154.200 ;
        RECT 15.800 153.800 16.200 154.200 ;
        RECT 20.600 153.800 21.000 154.200 ;
        RECT 1.400 146.800 1.800 147.200 ;
        RECT 2.200 143.100 2.600 148.900 ;
        RECT 3.800 146.800 4.200 147.200 ;
        RECT 3.800 146.200 4.100 146.800 ;
        RECT 3.800 145.800 4.200 146.200 ;
        RECT 5.400 145.800 5.800 146.200 ;
        RECT 5.400 144.200 5.700 145.800 ;
        RECT 5.400 143.800 5.800 144.200 ;
        RECT 3.000 139.100 3.400 139.200 ;
        RECT 3.800 139.100 4.200 139.200 ;
        RECT 3.000 138.800 4.200 139.100 ;
        RECT 4.600 133.100 5.000 135.900 ;
        RECT 5.400 134.200 5.700 143.800 ;
        RECT 7.000 143.100 7.400 148.900 ;
        RECT 15.000 147.200 15.300 153.800 ;
        RECT 22.200 153.100 22.600 153.200 ;
        RECT 23.000 153.100 23.400 153.200 ;
        RECT 22.200 152.800 23.400 153.100 ;
        RECT 17.400 152.100 17.800 152.200 ;
        RECT 18.200 152.100 18.600 152.200 ;
        RECT 17.400 151.800 18.600 152.100 ;
        RECT 10.200 146.800 10.600 147.200 ;
        RECT 11.800 147.100 12.200 147.200 ;
        RECT 12.600 147.100 13.000 147.200 ;
        RECT 11.800 146.800 13.000 147.100 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 15.000 147.100 15.400 147.200 ;
        RECT 14.200 146.800 15.400 147.100 ;
        RECT 10.200 144.200 10.500 146.800 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 15.000 146.100 15.400 146.200 ;
        RECT 14.200 145.800 15.400 146.100 ;
        RECT 11.800 145.200 12.100 145.800 ;
        RECT 11.800 144.800 12.200 145.200 ;
        RECT 15.800 145.100 16.200 147.900 ;
        RECT 16.600 146.800 17.000 147.200 ;
        RECT 16.600 144.200 16.900 146.800 ;
        RECT 10.200 143.800 10.600 144.200 ;
        RECT 16.600 143.800 17.000 144.200 ;
        RECT 10.200 140.200 10.500 143.800 ;
        RECT 17.400 143.100 17.800 148.900 ;
        RECT 19.800 146.100 20.200 146.200 ;
        RECT 20.600 146.100 21.000 146.200 ;
        RECT 19.800 145.800 21.000 146.100 ;
        RECT 21.400 142.800 21.800 143.200 ;
        RECT 22.200 143.100 22.600 148.900 ;
        RECT 10.200 139.800 10.600 140.200 ;
        RECT 5.400 133.800 5.800 134.200 ;
        RECT 6.200 132.100 6.600 137.900 ;
        RECT 7.800 135.100 8.200 135.200 ;
        RECT 8.600 135.100 9.000 135.200 ;
        RECT 7.800 134.800 9.000 135.100 ;
        RECT 11.000 132.100 11.400 137.900 ;
        RECT 15.000 137.800 15.400 138.200 ;
        RECT 17.400 137.800 17.800 138.200 ;
        RECT 15.000 135.200 15.300 137.800 ;
        RECT 17.400 136.200 17.700 137.800 ;
        RECT 17.400 135.800 17.800 136.200 ;
        RECT 19.800 135.800 20.200 136.200 ;
        RECT 19.800 135.200 20.100 135.800 ;
        RECT 21.400 135.200 21.700 142.800 ;
        RECT 23.000 139.800 23.400 140.200 ;
        RECT 23.000 135.200 23.300 139.800 ;
        RECT 15.000 134.800 15.400 135.200 ;
        RECT 15.800 135.100 16.200 135.200 ;
        RECT 16.600 135.100 17.000 135.200 ;
        RECT 15.800 134.800 17.000 135.100 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 21.400 134.800 21.800 135.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 14.200 134.100 14.600 134.200 ;
        RECT 15.000 134.100 15.400 134.200 ;
        RECT 14.200 133.800 15.400 134.100 ;
        RECT 15.800 133.800 16.200 134.200 ;
        RECT 19.000 133.800 19.400 134.200 ;
        RECT 21.400 133.800 21.800 134.200 ;
        RECT 13.400 132.800 13.800 133.200 ;
        RECT 13.400 132.200 13.700 132.800 ;
        RECT 13.400 131.800 13.800 132.200 ;
        RECT 14.200 131.800 14.600 132.200 ;
        RECT 0.600 125.100 1.000 127.900 ;
        RECT 1.400 126.800 1.800 127.200 ;
        RECT 1.400 119.200 1.700 126.800 ;
        RECT 2.200 123.100 2.600 128.900 ;
        RECT 5.400 126.800 5.800 127.200 ;
        RECT 5.400 126.200 5.700 126.800 ;
        RECT 5.400 125.800 5.800 126.200 ;
        RECT 7.000 123.100 7.400 128.900 ;
        RECT 9.400 128.800 9.800 129.200 ;
        RECT 9.400 128.200 9.700 128.800 ;
        RECT 9.400 127.800 9.800 128.200 ;
        RECT 11.800 127.800 12.200 128.200 ;
        RECT 11.800 127.200 12.100 127.800 ;
        RECT 11.800 126.800 12.200 127.200 ;
        RECT 12.600 126.800 13.000 127.200 ;
        RECT 12.600 126.200 12.900 126.800 ;
        RECT 14.200 126.200 14.500 131.800 ;
        RECT 15.800 127.200 16.100 133.800 ;
        RECT 19.000 133.200 19.300 133.800 ;
        RECT 21.400 133.200 21.700 133.800 ;
        RECT 19.000 132.800 19.400 133.200 ;
        RECT 21.400 132.800 21.800 133.200 ;
        RECT 19.000 129.200 19.300 132.800 ;
        RECT 19.800 131.800 20.200 132.200 ;
        RECT 19.000 128.800 19.400 129.200 ;
        RECT 15.000 126.800 15.400 127.200 ;
        RECT 15.800 126.800 16.200 127.200 ;
        RECT 17.400 127.100 17.800 127.200 ;
        RECT 18.200 127.100 18.600 127.200 ;
        RECT 17.400 126.800 18.600 127.100 ;
        RECT 12.600 125.800 13.000 126.200 ;
        RECT 14.200 125.800 14.600 126.200 ;
        RECT 14.200 125.200 14.500 125.800 ;
        RECT 10.200 125.100 10.600 125.200 ;
        RECT 11.000 125.100 11.400 125.200 ;
        RECT 10.200 124.800 11.400 125.100 ;
        RECT 14.200 124.800 14.600 125.200 ;
        RECT 10.200 123.800 10.600 124.200 ;
        RECT 15.000 124.100 15.300 126.800 ;
        RECT 16.600 126.100 17.000 126.200 ;
        RECT 17.400 126.100 17.800 126.200 ;
        RECT 16.600 125.800 17.800 126.100 ;
        RECT 18.200 125.800 18.600 126.200 ;
        RECT 18.200 125.200 18.500 125.800 ;
        RECT 18.200 124.800 18.600 125.200 ;
        RECT 19.000 125.100 19.400 127.900 ;
        RECT 19.800 125.200 20.100 131.800 ;
        RECT 19.800 124.800 20.200 125.200 ;
        RECT 14.200 123.800 15.300 124.100 ;
        RECT 1.400 118.800 1.800 119.200 ;
        RECT 9.400 116.800 9.800 117.200 ;
        RECT 9.400 116.200 9.700 116.800 ;
        RECT 7.800 115.800 8.200 116.200 ;
        RECT 9.400 115.800 9.800 116.200 ;
        RECT 7.800 114.200 8.100 115.800 ;
        RECT 7.000 113.800 7.400 114.200 ;
        RECT 7.800 113.800 8.200 114.200 ;
        RECT 7.000 113.200 7.300 113.800 ;
        RECT 7.000 112.800 7.400 113.200 ;
        RECT 1.400 111.800 1.800 112.200 ;
        RECT 1.400 109.200 1.700 111.800 ;
        RECT 1.400 108.800 1.800 109.200 ;
        RECT 0.600 105.100 1.000 107.900 ;
        RECT 1.400 107.200 1.700 108.800 ;
        RECT 1.400 106.800 1.800 107.200 ;
        RECT 2.200 103.100 2.600 108.900 ;
        RECT 3.000 105.900 3.400 106.300 ;
        RECT 3.000 102.100 3.300 105.900 ;
        RECT 7.000 103.100 7.400 108.900 ;
        RECT 10.200 107.200 10.500 123.800 ;
        RECT 12.600 121.800 13.000 122.200 ;
        RECT 12.600 117.200 12.900 121.800 ;
        RECT 12.600 116.800 13.000 117.200 ;
        RECT 12.600 115.200 12.900 116.800 ;
        RECT 11.000 115.100 11.400 115.200 ;
        RECT 11.800 115.100 12.200 115.200 ;
        RECT 11.000 114.800 12.200 115.100 ;
        RECT 12.600 114.800 13.000 115.200 ;
        RECT 11.000 113.800 11.400 114.200 ;
        RECT 11.800 114.100 12.200 114.200 ;
        RECT 12.600 114.100 13.000 114.200 ;
        RECT 11.800 113.800 13.000 114.100 ;
        RECT 11.000 109.200 11.300 113.800 ;
        RECT 13.400 113.100 13.800 115.900 ;
        RECT 14.200 114.200 14.500 123.800 ;
        RECT 20.600 123.100 21.000 128.900 ;
        RECT 23.800 127.200 24.100 154.800 ;
        RECT 26.200 154.200 26.500 156.800 ;
        RECT 25.400 154.100 25.800 154.200 ;
        RECT 26.200 154.100 26.600 154.200 ;
        RECT 25.400 153.800 26.600 154.100 ;
        RECT 28.600 152.100 29.000 157.900 ;
        RECT 30.200 154.800 30.600 155.200 ;
        RECT 30.200 153.200 30.500 154.800 ;
        RECT 30.200 152.800 30.600 153.200 ;
        RECT 25.400 146.800 25.800 147.200 ;
        RECT 30.200 146.800 30.600 147.200 ;
        RECT 25.400 143.100 25.700 146.800 ;
        RECT 26.200 145.800 26.600 146.200 ;
        RECT 27.000 146.100 27.400 146.200 ;
        RECT 27.800 146.100 28.200 146.200 ;
        RECT 27.000 145.800 28.200 146.100 ;
        RECT 26.200 144.200 26.500 145.800 ;
        RECT 28.600 144.800 29.000 145.200 ;
        RECT 28.600 144.200 28.900 144.800 ;
        RECT 26.200 143.800 26.600 144.200 ;
        RECT 28.600 143.800 29.000 144.200 ;
        RECT 25.400 142.800 26.500 143.100 ;
        RECT 24.600 142.100 25.000 142.200 ;
        RECT 25.400 142.100 25.800 142.200 ;
        RECT 24.600 141.800 25.800 142.100 ;
        RECT 24.600 136.800 25.000 137.200 ;
        RECT 24.600 136.200 24.900 136.800 ;
        RECT 24.600 135.800 25.000 136.200 ;
        RECT 25.400 134.800 25.800 135.200 ;
        RECT 25.400 133.200 25.700 134.800 ;
        RECT 26.200 134.200 26.500 142.800 ;
        RECT 30.200 142.200 30.500 146.800 ;
        RECT 30.200 141.800 30.600 142.200 ;
        RECT 27.000 138.800 27.400 139.200 ;
        RECT 27.000 136.200 27.300 138.800 ;
        RECT 27.000 135.800 27.400 136.200 ;
        RECT 27.000 135.200 27.300 135.800 ;
        RECT 27.000 134.800 27.400 135.200 ;
        RECT 26.200 133.800 26.600 134.200 ;
        RECT 28.600 134.100 29.000 134.200 ;
        RECT 29.400 134.100 29.800 134.200 ;
        RECT 28.600 133.800 29.800 134.100 ;
        RECT 25.400 132.800 25.800 133.200 ;
        RECT 27.800 132.800 28.200 133.200 ;
        RECT 27.800 129.200 28.100 132.800 ;
        RECT 31.800 132.200 32.100 164.800 ;
        RECT 37.400 164.100 37.800 164.200 ;
        RECT 38.200 164.100 38.600 164.200 ;
        RECT 37.400 163.800 38.600 164.100 ;
        RECT 36.600 162.800 37.000 163.200 ;
        RECT 36.600 159.200 36.900 162.800 ;
        RECT 39.000 161.800 39.400 162.200 ;
        RECT 39.000 159.200 39.300 161.800 ;
        RECT 39.800 161.200 40.100 165.800 ;
        RECT 42.200 165.100 42.600 165.200 ;
        RECT 43.000 165.100 43.400 165.200 ;
        RECT 42.200 164.800 43.400 165.100 ;
        RECT 43.800 164.200 44.100 165.800 ;
        RECT 44.600 165.200 44.900 174.800 ;
        RECT 45.400 174.200 45.700 185.800 ;
        RECT 50.200 183.100 50.600 188.900 ;
        RECT 54.200 188.800 54.600 189.200 ;
        RECT 51.000 187.800 51.400 188.200 ;
        RECT 51.000 186.200 51.300 187.800 ;
        RECT 51.000 185.800 51.400 186.200 ;
        RECT 53.400 185.800 53.800 186.200 ;
        RECT 53.400 185.200 53.700 185.800 ;
        RECT 53.400 184.800 53.800 185.200 ;
        RECT 53.400 183.800 53.800 184.200 ;
        RECT 53.400 179.200 53.700 183.800 ;
        RECT 55.000 183.100 55.400 188.900 ;
        RECT 55.800 188.200 56.100 193.800 ;
        RECT 61.400 193.200 61.700 193.800 ;
        RECT 61.400 192.800 61.800 193.200 ;
        RECT 55.800 187.800 56.200 188.200 ;
        RECT 56.600 185.100 57.000 187.900 ;
        RECT 60.600 186.800 61.000 187.200 ;
        RECT 60.600 186.200 60.900 186.800 ;
        RECT 57.400 185.800 57.800 186.200 ;
        RECT 58.200 185.800 58.600 186.200 ;
        RECT 60.600 185.800 61.000 186.200 ;
        RECT 57.400 185.200 57.700 185.800 ;
        RECT 57.400 184.800 57.800 185.200 ;
        RECT 57.400 182.800 57.800 183.200 ;
        RECT 51.800 178.800 52.200 179.200 ;
        RECT 53.400 178.800 53.800 179.200 ;
        RECT 48.600 177.800 49.000 178.200 ;
        RECT 48.600 175.200 48.900 177.800 ;
        RECT 51.000 175.800 51.400 176.200 ;
        RECT 47.000 175.100 47.400 175.200 ;
        RECT 47.800 175.100 48.200 175.200 ;
        RECT 47.000 174.800 48.200 175.100 ;
        RECT 48.600 174.800 49.000 175.200 ;
        RECT 45.400 173.800 45.800 174.200 ;
        RECT 45.400 169.200 45.700 173.800 ;
        RECT 51.000 169.200 51.300 175.800 ;
        RECT 51.800 175.200 52.100 178.800 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 52.600 176.200 52.900 176.800 ;
        RECT 52.600 175.800 53.000 176.200 ;
        RECT 51.800 174.800 52.200 175.200 ;
        RECT 52.600 174.800 53.000 175.200 ;
        RECT 54.200 175.100 54.600 175.200 ;
        RECT 55.000 175.100 55.400 175.200 ;
        RECT 54.200 174.800 55.400 175.100 ;
        RECT 52.600 174.200 52.900 174.800 ;
        RECT 57.400 174.200 57.700 182.800 ;
        RECT 58.200 178.100 58.500 185.800 ;
        RECT 62.200 184.200 62.500 193.800 ;
        RECT 63.000 187.800 63.400 188.200 ;
        RECT 65.400 187.800 65.800 188.200 ;
        RECT 63.000 186.200 63.300 187.800 ;
        RECT 65.400 186.200 65.700 187.800 ;
        RECT 66.200 186.200 66.500 210.800 ;
        RECT 67.000 206.200 67.300 213.800 ;
        RECT 67.800 213.100 68.200 215.900 ;
        RECT 68.600 215.800 69.800 216.100 ;
        RECT 76.600 215.200 76.900 233.800 ;
        RECT 78.200 232.100 78.600 237.900 ;
        RECT 82.200 234.700 82.600 235.100 ;
        RECT 80.600 230.800 81.000 231.200 ;
        RECT 78.200 223.100 78.600 228.900 ;
        RECT 79.000 226.800 79.400 227.200 ;
        RECT 79.000 226.200 79.300 226.800 ;
        RECT 79.000 225.800 79.400 226.200 ;
        RECT 80.600 215.200 80.900 230.800 ;
        RECT 82.200 230.200 82.500 234.700 ;
        RECT 83.000 232.100 83.400 237.900 ;
        RECT 85.400 237.800 85.800 238.200 ;
        RECT 112.600 238.100 113.000 238.200 ;
        RECT 113.400 238.100 113.800 238.200 ;
        RECT 83.800 233.800 84.200 234.200 ;
        RECT 83.800 233.200 84.100 233.800 ;
        RECT 83.800 232.800 84.200 233.200 ;
        RECT 84.600 233.100 85.000 235.900 ;
        RECT 85.400 235.200 85.700 237.800 ;
        RECT 85.400 234.800 85.800 235.200 ;
        RECT 90.200 234.800 90.600 235.200 ;
        RECT 85.400 231.200 85.700 234.800 ;
        RECT 87.000 231.800 87.400 232.200 ;
        RECT 85.400 230.800 85.800 231.200 ;
        RECT 82.200 229.800 82.600 230.200 ;
        RECT 87.000 229.200 87.300 231.800 ;
        RECT 81.400 226.100 81.800 226.200 ;
        RECT 82.200 226.100 82.600 226.300 ;
        RECT 81.400 225.900 82.600 226.100 ;
        RECT 81.400 225.800 82.500 225.900 ;
        RECT 83.000 223.100 83.400 228.900 ;
        RECT 87.000 228.800 87.400 229.200 ;
        RECT 90.200 228.200 90.500 234.800 ;
        RECT 91.000 233.800 91.400 234.200 ;
        RECT 97.400 234.100 97.800 234.200 ;
        RECT 98.200 234.100 98.600 234.200 ;
        RECT 97.400 233.800 98.600 234.100 ;
        RECT 83.800 226.800 84.200 227.200 ;
        RECT 70.200 214.800 70.600 215.200 ;
        RECT 71.800 215.100 72.200 215.200 ;
        RECT 72.600 215.100 73.000 215.200 ;
        RECT 71.800 214.800 73.000 215.100 ;
        RECT 75.000 214.800 75.400 215.200 ;
        RECT 76.600 214.800 77.000 215.200 ;
        RECT 80.600 214.800 81.000 215.200 ;
        RECT 67.000 205.800 67.400 206.200 ;
        RECT 67.000 204.800 67.400 205.200 ;
        RECT 67.000 187.200 67.300 204.800 ;
        RECT 67.800 203.100 68.200 208.900 ;
        RECT 68.600 206.100 69.000 206.200 ;
        RECT 69.400 206.100 69.800 206.200 ;
        RECT 68.600 205.800 69.800 206.100 ;
        RECT 70.200 202.200 70.500 214.800 ;
        RECT 71.000 214.100 71.400 214.200 ;
        RECT 71.800 214.100 72.200 214.200 ;
        RECT 71.000 213.800 72.200 214.100 ;
        RECT 72.600 213.800 73.000 214.200 ;
        RECT 72.600 211.200 72.900 213.800 ;
        RECT 75.000 213.200 75.300 214.800 ;
        RECT 76.600 214.200 76.900 214.800 ;
        RECT 76.600 213.800 77.000 214.200 ;
        RECT 77.400 214.100 77.800 214.200 ;
        RECT 78.200 214.100 78.600 214.200 ;
        RECT 77.400 213.800 78.600 214.100 ;
        RECT 74.200 212.800 74.600 213.200 ;
        RECT 75.000 212.800 75.400 213.200 ;
        RECT 81.400 213.100 81.800 215.900 ;
        RECT 74.200 212.200 74.500 212.800 ;
        RECT 73.400 211.800 73.800 212.200 ;
        RECT 74.200 211.800 74.600 212.200 ;
        RECT 75.800 211.800 76.200 212.200 ;
        RECT 83.000 212.100 83.400 217.900 ;
        RECT 83.800 214.200 84.100 226.800 ;
        RECT 84.600 225.100 85.000 227.900 ;
        RECT 85.400 227.800 85.800 228.200 ;
        RECT 90.200 227.800 90.600 228.200 ;
        RECT 85.400 227.200 85.700 227.800 ;
        RECT 91.000 227.200 91.300 233.800 ;
        RECT 99.800 233.100 100.200 235.900 ;
        RECT 100.600 233.800 101.000 234.200 ;
        RECT 100.600 233.200 100.900 233.800 ;
        RECT 100.600 232.800 101.000 233.200 ;
        RECT 91.800 231.800 92.200 232.200 ;
        RECT 101.400 232.100 101.800 237.900 ;
        RECT 104.600 236.800 105.000 237.200 ;
        RECT 104.600 235.200 104.900 236.800 ;
        RECT 104.600 234.800 105.000 235.200 ;
        RECT 106.200 232.100 106.600 237.900 ;
        RECT 112.600 237.800 113.800 238.100 ;
        RECT 111.000 236.800 111.400 237.200 ;
        RECT 110.200 235.800 110.600 236.200 ;
        RECT 110.200 235.200 110.500 235.800 ;
        RECT 111.000 235.200 111.300 236.800 ;
        RECT 111.800 236.100 112.200 236.200 ;
        RECT 112.600 236.100 113.000 236.200 ;
        RECT 111.800 235.800 113.000 236.100 ;
        RECT 110.200 234.800 110.600 235.200 ;
        RECT 111.000 234.800 111.400 235.200 ;
        RECT 110.200 234.200 110.500 234.800 ;
        RECT 109.400 233.800 109.800 234.200 ;
        RECT 110.200 233.800 110.600 234.200 ;
        RECT 108.600 231.800 109.000 232.200 ;
        RECT 85.400 226.800 85.800 227.200 ;
        RECT 90.200 226.800 90.600 227.200 ;
        RECT 91.000 226.800 91.400 227.200 ;
        RECT 86.200 226.100 86.600 226.200 ;
        RECT 87.000 226.100 87.400 226.200 ;
        RECT 86.200 225.800 87.400 226.100 ;
        RECT 87.800 225.800 88.200 226.200 ;
        RECT 87.800 225.200 88.100 225.800 ;
        RECT 85.400 225.100 85.800 225.200 ;
        RECT 86.200 225.100 86.600 225.200 ;
        RECT 85.400 224.800 86.600 225.100 ;
        RECT 87.000 224.800 87.400 225.200 ;
        RECT 87.800 224.800 88.200 225.200 ;
        RECT 87.000 223.200 87.300 224.800 ;
        RECT 87.000 222.800 87.400 223.200 ;
        RECT 87.000 220.200 87.300 222.800 ;
        RECT 89.400 221.800 89.800 222.200 ;
        RECT 87.000 219.800 87.400 220.200 ;
        RECT 84.600 215.800 85.000 216.200 ;
        RECT 84.600 215.200 84.900 215.800 ;
        RECT 84.600 214.800 85.000 215.200 ;
        RECT 83.800 213.800 84.200 214.200 ;
        RECT 87.800 212.100 88.200 217.900 ;
        RECT 72.600 210.800 73.000 211.200 ;
        RECT 71.800 205.900 72.200 206.300 ;
        RECT 71.800 205.200 72.100 205.900 ;
        RECT 71.800 204.800 72.200 205.200 ;
        RECT 72.600 203.100 73.000 208.900 ;
        RECT 73.400 206.200 73.700 211.800 ;
        RECT 75.800 209.200 76.100 211.800 ;
        RECT 76.600 210.800 77.000 211.200 ;
        RECT 79.000 210.800 79.400 211.200 ;
        RECT 75.800 208.800 76.200 209.200 ;
        RECT 73.400 205.800 73.800 206.200 ;
        RECT 74.200 205.100 74.600 207.900 ;
        RECT 75.000 207.800 75.400 208.200 ;
        RECT 75.000 207.200 75.300 207.800 ;
        RECT 75.000 206.800 75.400 207.200 ;
        RECT 76.600 206.200 76.900 210.800 ;
        RECT 77.400 207.800 77.800 208.200 ;
        RECT 77.400 207.200 77.700 207.800 ;
        RECT 77.400 206.800 77.800 207.200 ;
        RECT 76.600 205.800 77.000 206.200 ;
        RECT 70.200 201.800 70.600 202.200 ;
        RECT 76.600 200.200 76.900 205.800 ;
        RECT 79.000 205.200 79.300 210.800 ;
        RECT 79.000 204.800 79.400 205.200 ;
        RECT 79.800 205.100 80.200 207.900 ;
        RECT 78.200 201.800 78.600 202.200 ;
        RECT 76.600 199.800 77.000 200.200 ;
        RECT 74.200 198.800 74.600 199.200 ;
        RECT 67.800 196.800 68.200 197.200 ;
        RECT 67.800 196.200 68.100 196.800 ;
        RECT 67.800 195.800 68.200 196.200 ;
        RECT 68.600 196.100 69.000 196.200 ;
        RECT 69.400 196.100 69.800 196.200 ;
        RECT 68.600 195.800 69.800 196.100 ;
        RECT 71.000 195.800 71.400 196.200 ;
        RECT 68.600 194.800 69.000 195.200 ;
        RECT 69.400 195.100 69.800 195.200 ;
        RECT 70.200 195.100 70.600 195.200 ;
        RECT 69.400 194.800 70.600 195.100 ;
        RECT 68.600 194.200 68.900 194.800 ;
        RECT 67.800 193.800 68.200 194.200 ;
        RECT 68.600 193.800 69.000 194.200 ;
        RECT 67.800 192.200 68.100 193.800 ;
        RECT 67.800 191.800 68.200 192.200 ;
        RECT 67.000 186.800 67.400 187.200 ;
        RECT 67.800 186.800 68.200 187.200 ;
        RECT 67.800 186.200 68.100 186.800 ;
        RECT 71.000 186.200 71.300 195.800 ;
        RECT 74.200 195.200 74.500 198.800 ;
        RECT 78.200 196.200 78.500 201.800 ;
        RECT 78.200 195.800 78.600 196.200 ;
        RECT 74.200 194.800 74.600 195.200 ;
        RECT 77.400 194.800 77.800 195.200 ;
        RECT 79.000 195.100 79.300 204.800 ;
        RECT 79.800 203.800 80.200 204.200 ;
        RECT 79.800 199.200 80.100 203.800 ;
        RECT 81.400 203.100 81.800 208.900 ;
        RECT 83.000 206.800 83.400 207.200 ;
        RECT 82.200 205.900 82.600 206.300 ;
        RECT 82.200 204.200 82.500 205.900 ;
        RECT 82.200 203.800 82.600 204.200 ;
        RECT 79.800 198.800 80.200 199.200 ;
        RECT 83.000 197.200 83.300 206.800 ;
        RECT 86.200 203.100 86.600 208.900 ;
        RECT 88.600 208.800 89.000 209.200 ;
        RECT 88.600 208.200 88.900 208.800 ;
        RECT 88.600 207.800 89.000 208.200 ;
        RECT 89.400 206.200 89.700 221.800 ;
        RECT 90.200 215.200 90.500 226.800 ;
        RECT 91.800 226.200 92.100 231.800 ;
        RECT 108.600 231.200 108.900 231.800 ;
        RECT 108.600 230.800 109.000 231.200 ;
        RECT 109.400 229.200 109.700 233.800 ;
        RECT 116.600 233.100 117.000 235.900 ;
        RECT 117.400 233.800 117.800 234.200 ;
        RECT 117.400 233.200 117.700 233.800 ;
        RECT 117.400 232.800 117.800 233.200 ;
        RECT 113.400 231.800 113.800 232.200 ;
        RECT 118.200 232.100 118.600 237.900 ;
        RECT 121.400 235.800 121.800 236.200 ;
        RECT 119.800 234.800 120.200 235.200 ;
        RECT 119.800 234.200 120.100 234.800 ;
        RECT 119.800 233.800 120.200 234.200 ;
        RECT 119.000 231.800 119.400 232.200 ;
        RECT 97.400 228.800 97.800 229.200 ;
        RECT 97.400 228.200 97.700 228.800 ;
        RECT 94.200 227.800 94.600 228.200 ;
        RECT 97.400 227.800 97.800 228.200 ;
        RECT 94.200 226.200 94.500 227.800 ;
        RECT 91.000 225.800 91.400 226.200 ;
        RECT 91.800 225.800 92.200 226.200 ;
        RECT 94.200 225.800 94.600 226.200 ;
        RECT 95.000 226.100 95.400 226.200 ;
        RECT 95.800 226.100 96.200 226.200 ;
        RECT 95.000 225.800 96.200 226.100 ;
        RECT 91.000 220.200 91.300 225.800 ;
        RECT 99.800 223.100 100.200 228.900 ;
        RECT 100.600 227.800 101.000 228.200 ;
        RECT 100.600 227.200 100.900 227.800 ;
        RECT 100.600 226.800 101.000 227.200 ;
        RECT 103.000 226.800 103.400 227.200 ;
        RECT 103.800 226.800 104.200 227.200 ;
        RECT 103.000 226.200 103.300 226.800 ;
        RECT 101.400 225.800 101.800 226.200 ;
        RECT 103.000 225.800 103.400 226.200 ;
        RECT 93.400 221.800 93.800 222.200 ;
        RECT 91.000 219.800 91.400 220.200 ;
        RECT 91.800 216.800 92.200 217.200 ;
        RECT 91.800 216.200 92.100 216.800 ;
        RECT 91.800 215.800 92.200 216.200 ;
        RECT 90.200 214.800 90.600 215.200 ;
        RECT 91.000 214.800 91.400 215.200 ;
        RECT 91.800 215.100 92.200 215.200 ;
        RECT 92.600 215.100 93.000 215.200 ;
        RECT 91.800 214.800 93.000 215.100 ;
        RECT 91.000 214.200 91.300 214.800 ;
        RECT 91.000 213.800 91.400 214.200 ;
        RECT 90.200 212.100 90.600 212.200 ;
        RECT 91.000 212.100 91.400 212.200 ;
        RECT 90.200 211.800 91.400 212.100 ;
        RECT 90.200 207.800 90.600 208.200 ;
        RECT 90.200 206.200 90.500 207.800 ;
        RECT 89.400 205.800 89.800 206.200 ;
        RECT 90.200 205.800 90.600 206.200 ;
        RECT 89.400 204.200 89.700 205.800 ;
        RECT 89.400 203.800 89.800 204.200 ;
        RECT 91.800 201.800 92.200 202.200 ;
        RECT 83.000 196.800 83.400 197.200 ;
        RECT 79.800 195.100 80.200 195.200 ;
        RECT 80.600 195.100 81.000 195.200 ;
        RECT 79.000 194.800 81.000 195.100 ;
        RECT 77.400 194.200 77.700 194.800 ;
        RECT 71.800 193.800 72.200 194.200 ;
        RECT 72.600 193.800 73.000 194.200 ;
        RECT 77.400 193.800 77.800 194.200 ;
        RECT 79.800 194.100 80.200 194.200 ;
        RECT 80.600 194.100 81.000 194.200 ;
        RECT 79.800 193.800 81.000 194.100 ;
        RECT 71.800 192.100 72.100 193.800 ;
        RECT 72.600 193.200 72.900 193.800 ;
        RECT 72.600 192.800 73.000 193.200 ;
        RECT 71.800 191.800 72.900 192.100 ;
        RECT 72.600 189.200 72.900 191.800 ;
        RECT 80.600 190.200 80.900 193.800 ;
        RECT 81.400 191.800 81.800 192.200 ;
        RECT 83.800 192.100 84.200 197.900 ;
        RECT 87.800 194.700 88.200 195.100 ;
        RECT 80.600 189.800 81.000 190.200 ;
        RECT 71.800 188.800 72.200 189.200 ;
        RECT 72.600 188.800 73.000 189.200 ;
        RECT 71.800 187.200 72.100 188.800 ;
        RECT 71.800 186.800 72.200 187.200 ;
        RECT 73.400 187.100 73.800 187.200 ;
        RECT 74.200 187.100 74.600 187.200 ;
        RECT 73.400 186.800 74.600 187.100 ;
        RECT 63.000 185.800 63.400 186.200 ;
        RECT 63.800 185.800 64.200 186.200 ;
        RECT 65.400 185.800 65.800 186.200 ;
        RECT 66.200 185.800 66.600 186.200 ;
        RECT 67.000 185.800 67.400 186.200 ;
        RECT 67.800 185.800 68.200 186.200 ;
        RECT 71.000 185.800 71.400 186.200 ;
        RECT 71.800 185.800 72.200 186.200 ;
        RECT 75.000 185.800 75.400 186.200 ;
        RECT 63.800 185.200 64.100 185.800 ;
        RECT 63.800 184.800 64.200 185.200 ;
        RECT 66.200 184.200 66.500 185.800 ;
        RECT 67.000 185.200 67.300 185.800 ;
        RECT 71.800 185.200 72.100 185.800 ;
        RECT 67.000 184.800 67.400 185.200 ;
        RECT 71.800 184.800 72.200 185.200 ;
        RECT 62.200 183.800 62.600 184.200 ;
        RECT 66.200 183.800 66.600 184.200 ;
        RECT 68.600 183.100 69.000 183.200 ;
        RECT 69.400 183.100 69.800 183.200 ;
        RECT 68.600 182.800 69.800 183.100 ;
        RECT 59.000 181.800 59.400 182.200 ;
        RECT 59.000 179.200 59.300 181.800 ;
        RECT 59.000 178.800 59.400 179.200 ;
        RECT 59.000 178.100 59.400 178.200 ;
        RECT 58.200 177.800 59.400 178.100 ;
        RECT 63.800 178.100 64.200 178.200 ;
        RECT 64.600 178.100 65.000 178.200 ;
        RECT 63.800 177.800 65.000 178.100 ;
        RECT 58.200 174.800 58.600 175.200 ;
        RECT 52.600 173.800 53.000 174.200 ;
        RECT 54.200 173.800 54.600 174.200 ;
        RECT 55.000 173.800 55.400 174.200 ;
        RECT 56.600 173.800 57.000 174.200 ;
        RECT 57.400 173.800 57.800 174.200 ;
        RECT 54.200 173.200 54.500 173.800 ;
        RECT 54.200 172.800 54.600 173.200 ;
        RECT 55.000 172.100 55.300 173.800 ;
        RECT 56.600 173.200 56.900 173.800 ;
        RECT 56.600 172.800 57.000 173.200 ;
        RECT 54.200 171.800 55.300 172.100 ;
        RECT 52.600 169.800 53.000 170.200 ;
        RECT 45.400 168.800 45.800 169.200 ;
        RECT 51.000 168.800 51.400 169.200 ;
        RECT 45.400 167.800 45.800 168.200 ;
        RECT 45.400 167.200 45.700 167.800 ;
        RECT 45.400 166.800 45.800 167.200 ;
        RECT 49.400 167.100 49.800 167.200 ;
        RECT 50.200 167.100 50.600 167.200 ;
        RECT 49.400 166.800 50.600 167.100 ;
        RECT 51.800 166.800 52.200 167.200 ;
        RECT 46.200 165.800 46.600 166.200 ;
        RECT 47.000 165.800 47.400 166.200 ;
        RECT 47.800 165.800 48.200 166.200 ;
        RECT 44.600 164.800 45.000 165.200 ;
        RECT 46.200 164.200 46.500 165.800 ;
        RECT 47.000 165.200 47.300 165.800 ;
        RECT 47.000 164.800 47.400 165.200 ;
        RECT 43.800 163.800 44.200 164.200 ;
        RECT 44.600 163.800 45.000 164.200 ;
        RECT 46.200 163.800 46.600 164.200 ;
        RECT 39.800 160.800 40.200 161.200 ;
        RECT 44.600 159.200 44.900 163.800 ;
        RECT 47.800 162.200 48.100 165.800 ;
        RECT 51.000 163.800 51.400 164.200 ;
        RECT 47.800 161.800 48.200 162.200 ;
        RECT 36.600 158.800 37.000 159.200 ;
        RECT 39.000 158.800 39.400 159.200 ;
        RECT 44.600 158.800 45.000 159.200 ;
        RECT 33.400 152.100 33.800 157.900 ;
        RECT 45.400 156.800 45.800 157.200 ;
        RECT 34.200 153.800 34.600 154.200 ;
        RECT 34.200 153.200 34.500 153.800 ;
        RECT 34.200 152.800 34.600 153.200 ;
        RECT 35.000 153.100 35.400 155.900 ;
        RECT 45.400 155.200 45.700 156.800 ;
        RECT 35.800 154.800 36.200 155.200 ;
        RECT 36.600 155.100 37.000 155.200 ;
        RECT 37.400 155.100 37.800 155.200 ;
        RECT 36.600 154.800 37.800 155.100 ;
        RECT 42.200 154.800 42.600 155.200 ;
        RECT 45.400 154.800 45.800 155.200 ;
        RECT 46.200 154.800 46.600 155.200 ;
        RECT 47.000 155.100 47.400 155.200 ;
        RECT 47.800 155.100 48.200 155.200 ;
        RECT 47.000 154.800 48.200 155.100 ;
        RECT 48.600 155.100 49.000 155.200 ;
        RECT 49.400 155.100 49.800 155.200 ;
        RECT 48.600 154.800 49.800 155.100 ;
        RECT 32.600 149.100 33.000 149.200 ;
        RECT 33.400 149.100 33.800 149.200 ;
        RECT 32.600 148.800 33.800 149.100 ;
        RECT 34.200 147.200 34.500 152.800 ;
        RECT 35.000 150.800 35.400 151.200 ;
        RECT 35.000 149.200 35.300 150.800 ;
        RECT 35.800 149.200 36.100 154.800 ;
        RECT 42.200 154.200 42.500 154.800 ;
        RECT 46.200 154.200 46.500 154.800 ;
        RECT 42.200 153.800 42.600 154.200 ;
        RECT 46.200 153.800 46.600 154.200 ;
        RECT 36.600 151.800 37.000 152.200 ;
        RECT 39.000 151.800 39.400 152.200 ;
        RECT 40.600 151.800 41.000 152.200 ;
        RECT 42.200 151.800 42.600 152.200 ;
        RECT 35.000 148.800 35.400 149.200 ;
        RECT 35.800 148.800 36.200 149.200 ;
        RECT 34.200 146.800 34.600 147.200 ;
        RECT 35.800 146.800 36.200 147.200 ;
        RECT 32.600 145.800 33.000 146.200 ;
        RECT 34.200 145.800 34.600 146.200 ;
        RECT 32.600 145.200 32.900 145.800 ;
        RECT 34.200 145.200 34.500 145.800 ;
        RECT 32.600 144.800 33.000 145.200 ;
        RECT 34.200 144.800 34.600 145.200 ;
        RECT 35.800 139.200 36.100 146.800 ;
        RECT 36.600 141.200 36.900 151.800 ;
        RECT 37.400 146.800 37.800 147.200 ;
        RECT 37.400 146.200 37.700 146.800 ;
        RECT 37.400 145.800 37.800 146.200 ;
        RECT 37.400 141.800 37.800 142.200 ;
        RECT 36.600 140.800 37.000 141.200 ;
        RECT 35.800 138.800 36.200 139.200 ;
        RECT 37.400 135.200 37.700 141.800 ;
        RECT 37.400 134.800 37.800 135.200 ;
        RECT 39.000 132.200 39.300 151.800 ;
        RECT 40.600 148.200 40.900 151.800 ;
        RECT 40.600 147.800 41.000 148.200 ;
        RECT 42.200 146.200 42.500 151.800 ;
        RECT 47.000 151.200 47.300 154.800 ;
        RECT 51.000 154.200 51.300 163.800 ;
        RECT 51.800 163.200 52.100 166.800 ;
        RECT 52.600 166.200 52.900 169.800 ;
        RECT 52.600 165.800 53.000 166.200 ;
        RECT 53.400 165.100 53.800 167.900 ;
        RECT 51.800 162.800 52.200 163.200 ;
        RECT 54.200 162.200 54.500 171.800 ;
        RECT 55.000 163.100 55.400 168.900 ;
        RECT 55.800 168.800 56.200 169.200 ;
        RECT 55.800 168.200 56.100 168.800 ;
        RECT 55.800 167.800 56.200 168.200 ;
        RECT 56.600 165.800 57.000 166.200 ;
        RECT 56.600 165.200 56.900 165.800 ;
        RECT 56.600 164.800 57.000 165.200 ;
        RECT 58.200 164.200 58.500 174.800 ;
        RECT 59.000 174.200 59.300 177.800 ;
        RECT 63.000 176.800 63.400 177.200 ;
        RECT 63.000 176.200 63.300 176.800 ;
        RECT 60.600 175.800 61.000 176.200 ;
        RECT 63.000 175.800 63.400 176.200 ;
        RECT 59.000 173.800 59.400 174.200 ;
        RECT 60.600 172.200 60.900 175.800 ;
        RECT 63.000 174.800 63.400 175.200 ;
        RECT 63.800 174.800 64.200 175.200 ;
        RECT 63.000 172.200 63.300 174.800 ;
        RECT 63.800 174.200 64.100 174.800 ;
        RECT 63.800 173.800 64.200 174.200 ;
        RECT 60.600 171.800 61.000 172.200 ;
        RECT 63.000 171.800 63.400 172.200 ;
        RECT 62.200 169.100 62.600 169.200 ;
        RECT 63.000 169.100 63.400 169.200 ;
        RECT 58.200 163.800 58.600 164.200 ;
        RECT 59.800 163.100 60.200 168.900 ;
        RECT 62.200 168.800 63.400 169.100 ;
        RECT 63.800 168.200 64.100 173.800 ;
        RECT 67.000 172.100 67.400 177.900 ;
        RECT 70.200 175.800 70.600 176.200 ;
        RECT 70.200 175.200 70.500 175.800 ;
        RECT 70.200 174.800 70.600 175.200 ;
        RECT 71.000 172.800 71.400 173.200 ;
        RECT 68.600 171.800 69.000 172.200 ;
        RECT 67.800 168.800 68.200 169.200 ;
        RECT 63.800 167.800 64.200 168.200 ;
        RECT 63.000 167.100 63.400 167.200 ;
        RECT 63.800 167.100 64.100 167.800 ;
        RECT 63.000 166.800 64.100 167.100 ;
        RECT 67.800 167.200 68.100 168.800 ;
        RECT 67.800 166.800 68.200 167.200 ;
        RECT 68.600 166.200 68.900 171.800 ;
        RECT 70.200 169.800 70.600 170.200 ;
        RECT 70.200 169.200 70.500 169.800 ;
        RECT 70.200 168.800 70.600 169.200 ;
        RECT 71.000 166.200 71.300 172.800 ;
        RECT 71.800 172.100 72.200 177.900 ;
        RECT 72.600 175.800 73.000 176.200 ;
        RECT 72.600 166.200 72.900 175.800 ;
        RECT 73.400 173.100 73.800 175.900 ;
        RECT 74.200 174.800 74.600 175.200 ;
        RECT 73.400 168.800 73.800 169.200 ;
        RECT 73.400 166.200 73.700 168.800 ;
        RECT 74.200 167.200 74.500 174.800 ;
        RECT 75.000 174.200 75.300 185.800 ;
        RECT 75.800 185.100 76.200 187.900 ;
        RECT 77.400 183.100 77.800 188.900 ;
        RECT 81.400 188.200 81.700 191.800 ;
        RECT 87.800 189.200 88.100 194.700 ;
        RECT 88.600 192.100 89.000 197.900 ;
        RECT 89.400 193.800 89.800 194.200 ;
        RECT 89.400 193.200 89.700 193.800 ;
        RECT 89.400 192.800 89.800 193.200 ;
        RECT 90.200 193.100 90.600 195.900 ;
        RECT 91.800 195.200 92.100 201.800 ;
        RECT 91.800 194.800 92.200 195.200 ;
        RECT 93.400 195.100 93.700 221.800 ;
        RECT 96.600 218.800 97.000 219.200 ;
        RECT 95.800 215.800 96.200 216.200 ;
        RECT 95.800 215.200 96.100 215.800 ;
        RECT 96.600 215.200 96.900 218.800 ;
        RECT 99.800 217.800 100.200 218.200 ;
        RECT 99.800 215.200 100.100 217.800 ;
        RECT 101.400 215.200 101.700 225.800 ;
        RECT 103.800 221.200 104.100 226.800 ;
        RECT 104.600 223.100 105.000 228.900 ;
        RECT 109.400 228.800 109.800 229.200 ;
        RECT 105.400 226.800 105.800 227.200 ;
        RECT 103.800 220.800 104.200 221.200 ;
        RECT 102.200 215.800 102.600 216.200 ;
        RECT 95.800 214.800 96.200 215.200 ;
        RECT 96.600 214.800 97.000 215.200 ;
        RECT 99.800 214.800 100.200 215.200 ;
        RECT 101.400 214.800 101.800 215.200 ;
        RECT 94.200 213.800 94.600 214.200 ;
        RECT 94.200 212.200 94.500 213.800 ;
        RECT 94.200 211.800 94.600 212.200 ;
        RECT 98.200 212.100 98.600 212.200 ;
        RECT 99.000 212.100 99.400 212.200 ;
        RECT 98.200 211.800 99.400 212.100 ;
        RECT 94.200 206.200 94.500 211.800 ;
        RECT 97.400 207.800 97.800 208.200 ;
        RECT 100.600 207.800 101.000 208.200 ;
        RECT 97.400 206.200 97.700 207.800 ;
        RECT 100.600 207.200 100.900 207.800 ;
        RECT 100.600 206.800 101.000 207.200 ;
        RECT 101.400 206.200 101.700 214.800 ;
        RECT 102.200 209.200 102.500 215.800 ;
        RECT 105.400 215.200 105.700 226.800 ;
        RECT 106.200 225.100 106.600 227.900 ;
        RECT 110.200 227.800 110.600 228.200 ;
        RECT 110.200 227.200 110.500 227.800 ;
        RECT 107.000 227.100 107.400 227.200 ;
        RECT 107.800 227.100 108.200 227.200 ;
        RECT 107.000 226.800 108.200 227.100 ;
        RECT 110.200 226.800 110.600 227.200 ;
        RECT 107.800 225.800 108.200 226.200 ;
        RECT 108.600 226.100 109.000 226.200 ;
        RECT 109.400 226.100 109.800 226.200 ;
        RECT 108.600 225.800 109.800 226.100 ;
        RECT 107.800 225.200 108.100 225.800 ;
        RECT 107.800 224.800 108.200 225.200 ;
        RECT 111.000 225.100 111.400 225.200 ;
        RECT 111.800 225.100 112.200 225.200 ;
        RECT 111.000 224.800 112.200 225.100 ;
        RECT 112.600 224.800 113.000 225.200 ;
        RECT 112.600 224.200 112.900 224.800 ;
        RECT 107.000 223.800 107.400 224.200 ;
        RECT 112.600 223.800 113.000 224.200 ;
        RECT 107.000 219.200 107.300 223.800 ;
        RECT 107.000 218.800 107.400 219.200 ;
        RECT 106.200 217.800 106.600 218.200 ;
        RECT 106.200 215.200 106.500 217.800 ;
        RECT 108.600 216.800 109.000 217.200 ;
        RECT 107.800 215.800 108.200 216.200 ;
        RECT 104.600 214.800 105.000 215.200 ;
        RECT 105.400 214.800 105.800 215.200 ;
        RECT 106.200 214.800 106.600 215.200 ;
        RECT 103.000 211.800 103.400 212.200 ;
        RECT 103.000 210.200 103.300 211.800 ;
        RECT 103.000 209.800 103.400 210.200 ;
        RECT 102.200 208.800 102.600 209.200 ;
        RECT 103.000 208.800 103.400 209.200 ;
        RECT 103.000 208.200 103.300 208.800 ;
        RECT 103.000 207.800 103.400 208.200 ;
        RECT 104.600 206.200 104.900 214.800 ;
        RECT 105.400 214.200 105.700 214.800 ;
        RECT 106.200 214.200 106.500 214.800 ;
        RECT 105.400 213.800 105.800 214.200 ;
        RECT 106.200 213.800 106.600 214.200 ;
        RECT 107.800 213.200 108.100 215.800 ;
        RECT 108.600 214.200 108.900 216.800 ;
        RECT 108.600 213.800 109.000 214.200 ;
        RECT 107.800 212.800 108.200 213.200 ;
        RECT 111.000 212.100 111.400 217.900 ;
        RECT 111.800 213.800 112.200 214.200 ;
        RECT 107.800 209.800 108.200 210.200 ;
        RECT 94.200 205.800 94.600 206.200 ;
        RECT 95.000 205.800 95.400 206.200 ;
        RECT 97.400 205.800 97.800 206.200 ;
        RECT 98.200 205.800 98.600 206.200 ;
        RECT 101.400 205.800 101.800 206.200 ;
        RECT 102.200 205.800 102.600 206.200 ;
        RECT 104.600 205.800 105.000 206.200 ;
        RECT 95.000 203.200 95.300 205.800 ;
        RECT 98.200 205.200 98.500 205.800 ;
        RECT 102.200 205.200 102.500 205.800 ;
        RECT 98.200 204.800 98.600 205.200 ;
        RECT 102.200 204.800 102.600 205.200 ;
        RECT 95.000 202.800 95.400 203.200 ;
        RECT 95.800 201.800 96.200 202.200 ;
        RECT 95.800 196.200 96.100 201.800 ;
        RECT 95.800 195.800 96.200 196.200 ;
        RECT 96.600 195.800 97.000 196.200 ;
        RECT 99.000 195.800 99.400 196.200 ;
        RECT 100.600 196.100 101.000 196.200 ;
        RECT 101.400 196.100 101.800 196.200 ;
        RECT 100.600 195.800 101.800 196.100 ;
        RECT 96.600 195.200 96.900 195.800 ;
        RECT 94.200 195.100 94.600 195.200 ;
        RECT 93.400 194.800 94.600 195.100 ;
        RECT 95.000 195.100 95.400 195.200 ;
        RECT 95.800 195.100 96.200 195.200 ;
        RECT 95.000 194.800 96.200 195.100 ;
        RECT 96.600 194.800 97.000 195.200 ;
        RECT 95.800 193.800 96.200 194.200 ;
        RECT 92.600 192.100 93.000 192.200 ;
        RECT 93.400 192.100 93.800 192.200 ;
        RECT 92.600 191.800 93.800 192.100 ;
        RECT 95.800 190.200 96.100 193.800 ;
        RECT 96.600 193.200 96.900 194.800 ;
        RECT 99.000 194.200 99.300 195.800 ;
        RECT 99.800 195.100 100.200 195.200 ;
        RECT 100.600 195.100 101.000 195.200 ;
        RECT 99.800 194.800 101.000 195.100 ;
        RECT 99.000 193.800 99.400 194.200 ;
        RECT 96.600 192.800 97.000 193.200 ;
        RECT 90.200 189.800 90.600 190.200 ;
        RECT 95.800 189.800 96.200 190.200 ;
        RECT 81.400 187.800 81.800 188.200 ;
        RECT 79.000 186.800 79.400 187.200 ;
        RECT 79.000 185.100 79.300 186.800 ;
        RECT 79.800 186.100 80.200 186.200 ;
        RECT 80.600 186.100 81.000 186.200 ;
        RECT 79.800 185.800 81.000 186.100 ;
        RECT 79.000 184.800 80.100 185.100 ;
        RECT 79.800 183.200 80.100 184.800 ;
        RECT 79.800 182.800 80.200 183.200 ;
        RECT 82.200 183.100 82.600 188.900 ;
        RECT 84.600 188.800 85.000 189.200 ;
        RECT 87.800 188.800 88.200 189.200 ;
        RECT 84.600 187.200 84.900 188.800 ;
        RECT 90.200 187.200 90.500 189.800 ;
        RECT 92.600 189.100 93.000 189.200 ;
        RECT 93.400 189.100 93.800 189.200 ;
        RECT 92.600 188.800 93.800 189.100 ;
        RECT 95.800 188.200 96.100 189.800 ;
        RECT 91.000 187.800 91.400 188.200 ;
        RECT 95.800 187.800 96.200 188.200 ;
        RECT 91.000 187.200 91.300 187.800 ;
        RECT 95.800 187.200 96.100 187.800 ;
        RECT 84.600 186.800 85.000 187.200 ;
        RECT 85.400 187.100 85.800 187.200 ;
        RECT 86.200 187.100 86.600 187.200 ;
        RECT 85.400 186.800 86.600 187.100 ;
        RECT 87.800 186.800 88.200 187.200 ;
        RECT 90.200 186.800 90.600 187.200 ;
        RECT 91.000 186.800 91.400 187.200 ;
        RECT 95.800 186.800 96.200 187.200 ;
        RECT 96.600 186.800 97.000 187.200 ;
        RECT 99.800 186.800 100.200 187.200 ;
        RECT 87.800 186.200 88.100 186.800 ;
        RECT 96.600 186.200 96.900 186.800 ;
        RECT 99.800 186.200 100.100 186.800 ;
        RECT 87.800 185.800 88.200 186.200 ;
        RECT 89.400 185.800 89.800 186.200 ;
        RECT 95.000 185.800 95.400 186.200 ;
        RECT 96.600 185.800 97.000 186.200 ;
        RECT 99.800 185.800 100.200 186.200 ;
        RECT 101.400 185.800 101.800 186.200 ;
        RECT 89.400 185.200 89.700 185.800 ;
        RECT 87.000 185.100 87.400 185.200 ;
        RECT 87.800 185.100 88.200 185.200 ;
        RECT 87.000 184.800 88.200 185.100 ;
        RECT 89.400 184.800 89.800 185.200 ;
        RECT 92.600 184.800 93.000 185.200 ;
        RECT 77.400 174.800 77.800 175.200 ;
        RECT 78.200 174.800 78.600 175.200 ;
        RECT 75.000 173.800 75.400 174.200 ;
        RECT 77.400 173.200 77.700 174.800 ;
        RECT 78.200 174.200 78.500 174.800 ;
        RECT 78.200 173.800 78.600 174.200 ;
        RECT 77.400 172.800 77.800 173.200 ;
        RECT 79.000 173.100 79.400 175.900 ;
        RECT 79.800 174.200 80.100 182.800 ;
        RECT 79.800 173.800 80.200 174.200 ;
        RECT 75.800 167.800 76.200 168.200 ;
        RECT 78.200 167.800 78.600 168.200 ;
        RECT 74.200 166.800 74.600 167.200 ;
        RECT 63.800 166.100 64.200 166.200 ;
        RECT 64.600 166.100 65.000 166.200 ;
        RECT 63.800 165.800 65.000 166.100 ;
        RECT 66.200 165.800 66.600 166.200 ;
        RECT 68.600 165.800 69.000 166.200 ;
        RECT 69.400 166.100 69.800 166.200 ;
        RECT 70.200 166.100 70.600 166.200 ;
        RECT 69.400 165.800 70.600 166.100 ;
        RECT 71.000 165.800 71.400 166.200 ;
        RECT 72.600 165.800 73.000 166.200 ;
        RECT 73.400 165.800 73.800 166.200 ;
        RECT 74.200 165.800 74.600 166.200 ;
        RECT 66.200 165.200 66.500 165.800 ;
        RECT 63.800 164.800 64.200 165.200 ;
        RECT 66.200 164.800 66.600 165.200 ;
        RECT 63.800 164.200 64.100 164.800 ;
        RECT 63.800 163.800 64.200 164.200 ;
        RECT 51.800 161.800 52.200 162.200 ;
        RECT 54.200 161.800 54.600 162.200 ;
        RECT 51.800 159.200 52.100 161.800 ;
        RECT 66.200 161.200 66.500 164.800 ;
        RECT 66.200 160.800 66.600 161.200 ;
        RECT 51.800 158.800 52.200 159.200 ;
        RECT 68.600 158.200 68.900 165.800 ;
        RECT 71.800 159.800 72.200 160.200 ;
        RECT 52.600 157.100 53.000 157.200 ;
        RECT 53.400 157.100 53.800 157.200 ;
        RECT 52.600 156.800 53.800 157.100 ;
        RECT 51.000 153.800 51.400 154.200 ;
        RECT 54.200 154.100 54.600 154.200 ;
        RECT 55.000 154.100 55.400 154.200 ;
        RECT 54.200 153.800 55.400 154.100 ;
        RECT 48.600 152.800 49.000 153.200 ;
        RECT 47.000 150.800 47.400 151.200 ;
        RECT 48.600 148.200 48.900 152.800 ;
        RECT 48.600 147.800 49.000 148.200 ;
        RECT 44.600 147.100 45.000 147.200 ;
        RECT 45.400 147.100 45.800 147.200 ;
        RECT 44.600 146.800 45.800 147.100 ;
        RECT 39.800 145.800 40.200 146.200 ;
        RECT 42.200 145.800 42.600 146.200 ;
        RECT 43.000 146.100 43.400 146.200 ;
        RECT 43.800 146.100 44.200 146.200 ;
        RECT 43.000 145.800 44.200 146.100 ;
        RECT 47.000 146.100 47.400 146.200 ;
        RECT 47.800 146.100 48.200 146.200 ;
        RECT 47.000 145.800 48.200 146.100 ;
        RECT 39.800 139.200 40.100 145.800 ;
        RECT 47.000 145.100 47.400 145.200 ;
        RECT 47.800 145.100 48.200 145.200 ;
        RECT 47.000 144.800 48.200 145.100 ;
        RECT 41.400 141.800 41.800 142.200 ;
        RECT 39.800 138.800 40.200 139.200 ;
        RECT 41.400 136.100 41.700 141.800 ;
        RECT 51.000 141.200 51.300 153.800 ;
        RECT 55.800 152.100 56.200 157.900 ;
        RECT 59.800 156.800 60.200 157.200 ;
        RECT 56.600 154.800 57.000 155.200 ;
        RECT 59.800 155.100 60.100 156.800 ;
        RECT 56.600 153.200 56.900 154.800 ;
        RECT 59.800 154.700 60.200 155.100 ;
        RECT 56.600 152.800 57.000 153.200 ;
        RECT 60.600 152.100 61.000 157.900 ;
        RECT 68.600 157.800 69.000 158.200 ;
        RECT 66.200 156.800 66.600 157.200 ;
        RECT 64.600 156.100 65.000 156.200 ;
        RECT 65.400 156.100 65.800 156.200 ;
        RECT 62.200 153.100 62.600 155.900 ;
        RECT 64.600 155.800 65.800 156.100 ;
        RECT 66.200 155.200 66.500 156.800 ;
        RECT 67.000 155.800 67.400 156.200 ;
        RECT 67.800 155.800 68.200 156.200 ;
        RECT 67.000 155.200 67.300 155.800 ;
        RECT 63.000 154.800 63.400 155.200 ;
        RECT 66.200 154.800 66.600 155.200 ;
        RECT 67.000 154.800 67.400 155.200 ;
        RECT 63.000 154.200 63.300 154.800 ;
        RECT 63.000 153.800 63.400 154.200 ;
        RECT 55.800 150.800 56.200 151.200 ;
        RECT 55.800 149.200 56.100 150.800 ;
        RECT 67.000 149.200 67.300 154.800 ;
        RECT 67.800 154.200 68.100 155.800 ;
        RECT 67.800 153.800 68.200 154.200 ;
        RECT 68.600 153.800 69.000 154.200 ;
        RECT 68.600 153.200 68.900 153.800 ;
        RECT 68.600 152.800 69.000 153.200 ;
        RECT 55.800 148.800 56.200 149.200 ;
        RECT 54.200 147.800 54.600 148.200 ;
        RECT 56.600 147.800 57.000 148.200 ;
        RECT 58.200 147.800 58.600 148.200 ;
        RECT 54.200 147.200 54.500 147.800 ;
        RECT 56.600 147.200 56.900 147.800 ;
        RECT 58.200 147.200 58.500 147.800 ;
        RECT 51.800 146.800 52.200 147.200 ;
        RECT 54.200 146.800 54.600 147.200 ;
        RECT 56.600 146.800 57.000 147.200 ;
        RECT 58.200 146.800 58.600 147.200 ;
        RECT 51.800 146.200 52.100 146.800 ;
        RECT 56.600 146.200 56.900 146.800 ;
        RECT 51.800 145.800 52.200 146.200 ;
        RECT 56.600 145.800 57.000 146.200 ;
        RECT 64.600 145.100 65.000 147.900 ;
        RECT 66.200 143.100 66.600 148.900 ;
        RECT 67.000 148.800 67.400 149.200 ;
        RECT 68.600 147.200 68.900 152.800 ;
        RECT 68.600 146.800 69.000 147.200 ;
        RECT 69.400 146.800 69.800 147.200 ;
        RECT 67.800 145.800 68.200 146.200 ;
        RECT 67.800 145.200 68.100 145.800 ;
        RECT 67.800 144.800 68.200 145.200 ;
        RECT 51.800 141.800 52.200 142.200 ;
        RECT 53.400 141.800 53.800 142.200 ;
        RECT 63.000 141.800 63.400 142.200 ;
        RECT 43.000 140.800 43.400 141.200 ;
        RECT 51.000 140.800 51.400 141.200 ;
        RECT 41.400 135.800 42.500 136.100 ;
        RECT 42.200 135.200 42.500 135.800 ;
        RECT 43.000 135.200 43.300 140.800 ;
        RECT 51.800 140.200 52.100 141.800 ;
        RECT 51.800 139.800 52.200 140.200 ;
        RECT 44.600 139.100 45.000 139.200 ;
        RECT 45.400 139.100 45.800 139.200 ;
        RECT 44.600 138.800 45.800 139.100 ;
        RECT 48.600 136.800 49.000 137.200 ;
        RECT 48.600 135.200 48.900 136.800 ;
        RECT 40.600 134.800 41.000 135.200 ;
        RECT 41.400 134.800 41.800 135.200 ;
        RECT 42.200 134.800 42.600 135.200 ;
        RECT 43.000 134.800 43.400 135.200 ;
        RECT 45.400 134.800 45.800 135.200 ;
        RECT 47.000 135.100 47.400 135.200 ;
        RECT 47.800 135.100 48.200 135.200 ;
        RECT 47.000 134.800 48.200 135.100 ;
        RECT 48.600 134.800 49.000 135.200 ;
        RECT 51.000 134.800 51.400 135.200 ;
        RECT 51.800 134.800 52.200 135.200 ;
        RECT 40.600 134.200 40.900 134.800 ;
        RECT 40.600 133.800 41.000 134.200 ;
        RECT 31.800 131.800 32.200 132.200 ;
        RECT 39.000 131.800 39.400 132.200 ;
        RECT 37.400 130.800 37.800 131.200 ;
        RECT 32.600 129.800 33.000 130.200 ;
        RECT 21.400 126.800 21.800 127.200 ;
        RECT 22.200 126.800 22.600 127.200 ;
        RECT 23.800 126.800 24.200 127.200 ;
        RECT 21.400 119.200 21.700 126.800 ;
        RECT 22.200 126.200 22.500 126.800 ;
        RECT 22.200 125.800 22.600 126.200 ;
        RECT 25.400 123.100 25.800 128.900 ;
        RECT 27.800 128.800 28.200 129.200 ;
        RECT 28.600 127.800 29.000 128.200 ;
        RECT 28.600 126.200 28.900 127.800 ;
        RECT 29.400 126.800 29.800 127.200 ;
        RECT 28.600 125.800 29.000 126.200 ;
        RECT 25.400 120.800 25.800 121.200 ;
        RECT 25.400 119.200 25.700 120.800 ;
        RECT 18.200 118.800 18.600 119.200 ;
        RECT 21.400 118.800 21.800 119.200 ;
        RECT 25.400 118.800 25.800 119.200 ;
        RECT 14.200 113.800 14.600 114.200 ;
        RECT 15.000 112.100 15.400 117.900 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 15.800 114.800 17.000 115.100 ;
        RECT 15.800 114.700 16.200 114.800 ;
        RECT 17.400 113.800 17.800 114.200 ;
        RECT 17.400 113.200 17.700 113.800 ;
        RECT 17.400 112.800 17.800 113.200 ;
        RECT 18.200 109.200 18.500 118.800 ;
        RECT 19.800 112.100 20.200 117.900 ;
        RECT 21.400 116.800 21.800 117.200 ;
        RECT 22.200 117.100 22.600 117.200 ;
        RECT 23.000 117.100 23.400 117.200 ;
        RECT 22.200 116.800 23.400 117.100 ;
        RECT 23.800 116.800 24.200 117.200 ;
        RECT 11.000 108.800 11.400 109.200 ;
        RECT 13.400 108.800 13.800 109.200 ;
        RECT 13.400 107.200 13.700 108.800 ;
        RECT 10.200 106.800 10.600 107.200 ;
        RECT 12.600 106.800 13.000 107.200 ;
        RECT 13.400 106.800 13.800 107.200 ;
        RECT 12.600 106.200 12.900 106.800 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 15.800 103.100 16.200 108.900 ;
        RECT 18.200 108.800 18.600 109.200 ;
        RECT 18.200 107.200 18.500 108.800 ;
        RECT 18.200 106.800 18.600 107.200 ;
        RECT 19.000 106.200 19.400 106.300 ;
        RECT 19.800 106.200 20.200 106.300 ;
        RECT 19.000 105.900 20.200 106.200 ;
        RECT 20.600 103.100 21.000 108.900 ;
        RECT 2.200 101.800 3.300 102.100 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 11.000 101.800 11.400 102.200 ;
        RECT 13.400 101.800 13.800 102.200 ;
        RECT 2.200 99.200 2.500 101.800 ;
        RECT 2.200 98.800 2.600 99.200 ;
        RECT 2.200 97.800 2.600 98.200 ;
        RECT 0.600 95.800 1.000 96.200 ;
        RECT 0.600 93.200 0.900 95.800 ;
        RECT 2.200 95.200 2.500 97.800 ;
        RECT 2.200 94.800 2.600 95.200 ;
        RECT 3.000 94.800 3.400 95.200 ;
        RECT 0.600 92.800 1.000 93.200 ;
        RECT 2.200 85.200 2.500 94.800 ;
        RECT 3.000 94.200 3.300 94.800 ;
        RECT 3.000 93.800 3.400 94.200 ;
        RECT 3.800 93.100 4.200 95.900 ;
        RECT 5.400 92.100 5.800 97.900 ;
        RECT 7.000 95.100 7.400 95.200 ;
        RECT 7.800 95.100 8.200 95.200 ;
        RECT 7.000 94.800 8.200 95.100 ;
        RECT 6.200 92.800 6.600 93.200 ;
        RECT 7.800 92.800 8.200 93.200 ;
        RECT 6.200 89.200 6.500 92.800 ;
        RECT 7.800 89.200 8.100 92.800 ;
        RECT 6.200 88.800 6.600 89.200 ;
        RECT 7.800 88.800 8.200 89.200 ;
        RECT 6.200 88.200 6.500 88.800 ;
        RECT 6.200 87.800 6.600 88.200 ;
        RECT 9.400 87.200 9.700 101.800 ;
        RECT 10.200 92.100 10.600 97.900 ;
        RECT 11.000 94.200 11.300 101.800 ;
        RECT 12.600 96.800 13.000 97.200 ;
        RECT 12.600 94.200 12.900 96.800 ;
        RECT 13.400 95.200 13.700 101.800 ;
        RECT 19.800 96.100 20.200 96.200 ;
        RECT 20.600 96.100 21.000 96.200 ;
        RECT 19.800 95.800 21.000 96.100 ;
        RECT 13.400 94.800 13.800 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 17.400 94.800 17.800 95.200 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 19.800 94.800 20.200 95.200 ;
        RECT 16.600 94.200 16.900 94.800 ;
        RECT 11.000 93.800 11.400 94.200 ;
        RECT 12.600 93.800 13.000 94.200 ;
        RECT 16.600 93.800 17.000 94.200 ;
        RECT 15.000 93.100 15.400 93.200 ;
        RECT 15.800 93.100 16.200 93.200 ;
        RECT 15.000 92.800 16.200 93.100 ;
        RECT 9.400 86.800 9.800 87.200 ;
        RECT 2.200 84.800 2.600 85.200 ;
        RECT 7.800 85.100 8.200 85.200 ;
        RECT 8.600 85.100 9.000 85.200 ;
        RECT 10.200 85.100 10.600 87.900 ;
        RECT 11.000 87.800 11.400 88.200 ;
        RECT 11.000 87.200 11.300 87.800 ;
        RECT 11.000 86.800 11.400 87.200 ;
        RECT 7.800 84.800 9.000 85.100 ;
        RECT 11.800 83.100 12.200 88.900 ;
        RECT 14.200 85.800 14.600 86.200 ;
        RECT 15.000 85.800 15.400 86.200 ;
        RECT 0.600 73.100 1.000 75.900 ;
        RECT 2.200 72.100 2.600 77.900 ;
        RECT 3.000 74.700 3.400 75.100 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 3.000 69.200 3.300 74.700 ;
        RECT 5.400 73.800 5.800 74.200 ;
        RECT 3.000 68.800 3.400 69.200 ;
        RECT 4.600 68.100 5.000 68.200 ;
        RECT 5.400 68.100 5.700 73.800 ;
        RECT 4.600 67.800 5.700 68.100 ;
        RECT 6.200 68.100 6.500 74.800 ;
        RECT 7.000 72.100 7.400 77.900 ;
        RECT 14.200 77.200 14.500 85.800 ;
        RECT 14.200 76.800 14.600 77.200 ;
        RECT 11.800 75.800 12.200 76.200 ;
        RECT 11.800 75.200 12.100 75.800 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 12.600 74.800 13.000 75.200 ;
        RECT 13.400 74.800 13.800 75.200 ;
        RECT 12.600 74.200 12.900 74.800 ;
        RECT 13.400 74.200 13.700 74.800 ;
        RECT 12.600 73.800 13.000 74.200 ;
        RECT 13.400 73.800 13.800 74.200 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 14.200 71.800 14.600 72.200 ;
        RECT 6.200 67.800 7.300 68.100 ;
        RECT 5.400 67.200 5.700 67.800 ;
        RECT 0.600 67.100 1.000 67.200 ;
        RECT 1.400 67.100 1.800 67.200 ;
        RECT 0.600 66.800 1.800 67.100 ;
        RECT 5.400 66.800 5.800 67.200 ;
        RECT 6.200 66.800 6.600 67.200 ;
        RECT 6.200 66.200 6.500 66.800 ;
        RECT 2.200 65.800 2.600 66.200 ;
        RECT 4.600 66.100 5.000 66.200 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 4.600 65.800 5.800 66.100 ;
        RECT 6.200 65.800 6.600 66.200 ;
        RECT 2.200 65.200 2.500 65.800 ;
        RECT 2.200 64.800 2.600 65.200 ;
        RECT 0.600 57.800 1.000 58.200 ;
        RECT 0.600 54.200 0.900 57.800 ;
        RECT 2.200 56.800 2.600 57.200 ;
        RECT 2.200 56.200 2.500 56.800 ;
        RECT 2.200 55.800 2.600 56.200 ;
        RECT 4.600 55.800 5.000 56.200 ;
        RECT 4.600 55.200 4.900 55.800 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 4.600 54.800 5.000 55.200 ;
        RECT 3.800 54.200 4.100 54.800 ;
        RECT 0.600 53.800 1.000 54.200 ;
        RECT 3.800 53.800 4.200 54.200 ;
        RECT 4.600 54.100 5.000 54.200 ;
        RECT 5.400 54.100 5.800 54.200 ;
        RECT 4.600 53.800 5.800 54.100 ;
        RECT 3.800 52.800 4.200 53.200 ;
        RECT 6.200 53.100 6.600 55.900 ;
        RECT 7.000 54.200 7.300 67.800 ;
        RECT 9.400 67.200 9.700 71.800 ;
        RECT 10.200 68.800 10.600 69.200 ;
        RECT 9.400 66.800 9.800 67.200 ;
        RECT 10.200 66.200 10.500 68.800 ;
        RECT 7.800 65.800 8.200 66.200 ;
        RECT 9.400 65.800 9.800 66.200 ;
        RECT 10.200 65.800 10.600 66.200 ;
        RECT 7.800 65.200 8.100 65.800 ;
        RECT 7.800 64.800 8.200 65.200 ;
        RECT 9.400 58.200 9.700 65.800 ;
        RECT 11.000 65.100 11.400 67.900 ;
        RECT 11.800 66.800 12.200 67.200 ;
        RECT 7.000 53.800 7.400 54.200 ;
        RECT 7.000 53.200 7.300 53.800 ;
        RECT 7.000 52.800 7.400 53.200 ;
        RECT 3.800 49.200 4.100 52.800 ;
        RECT 7.800 52.100 8.200 57.900 ;
        RECT 9.400 57.800 9.800 58.200 ;
        RECT 8.600 55.800 9.000 56.200 ;
        RECT 8.600 55.100 8.900 55.800 ;
        RECT 8.600 54.700 9.000 55.100 ;
        RECT 11.800 50.200 12.100 66.800 ;
        RECT 12.600 63.100 13.000 68.900 ;
        RECT 14.200 66.200 14.500 71.800 ;
        RECT 15.000 67.200 15.300 85.800 ;
        RECT 16.600 83.100 17.000 88.900 ;
        RECT 17.400 83.200 17.700 94.800 ;
        RECT 18.200 94.200 18.500 94.800 ;
        RECT 19.800 94.200 20.100 94.800 ;
        RECT 18.200 93.800 18.600 94.200 ;
        RECT 19.800 93.800 20.200 94.200 ;
        RECT 19.800 89.100 20.200 89.200 ;
        RECT 20.600 89.100 21.000 89.200 ;
        RECT 19.800 88.800 21.000 89.100 ;
        RECT 19.000 84.100 19.400 84.200 ;
        RECT 19.800 84.100 20.200 84.200 ;
        RECT 19.000 83.800 20.200 84.100 ;
        RECT 17.400 82.800 17.800 83.200 ;
        RECT 19.800 76.800 20.200 77.200 ;
        RECT 19.000 75.800 19.400 76.200 ;
        RECT 19.000 75.200 19.300 75.800 ;
        RECT 19.800 75.200 20.100 76.800 ;
        RECT 21.400 76.200 21.700 116.800 ;
        RECT 22.200 116.200 22.500 116.800 ;
        RECT 22.200 115.800 22.600 116.200 ;
        RECT 23.800 115.200 24.100 116.800 ;
        RECT 29.400 116.200 29.700 126.800 ;
        RECT 32.600 126.200 32.900 129.800 ;
        RECT 37.400 127.200 37.700 130.800 ;
        RECT 39.000 128.800 39.400 129.200 ;
        RECT 37.400 126.800 37.800 127.200 ;
        RECT 39.000 126.200 39.300 128.800 ;
        RECT 30.200 125.800 30.600 126.200 ;
        RECT 31.800 125.800 32.200 126.200 ;
        RECT 32.600 125.800 33.000 126.200 ;
        RECT 33.400 125.800 33.800 126.200 ;
        RECT 34.200 125.800 34.600 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 36.600 126.100 37.000 126.200 ;
        RECT 35.800 125.800 37.000 126.100 ;
        RECT 38.200 125.800 38.600 126.200 ;
        RECT 39.000 125.800 39.400 126.200 ;
        RECT 30.200 125.200 30.500 125.800 ;
        RECT 30.200 124.800 30.600 125.200 ;
        RECT 31.800 124.200 32.100 125.800 ;
        RECT 33.400 125.200 33.700 125.800 ;
        RECT 33.400 124.800 33.800 125.200 ;
        RECT 31.800 123.800 32.200 124.200 ;
        RECT 34.200 121.200 34.500 125.800 ;
        RECT 38.200 125.200 38.500 125.800 ;
        RECT 38.200 124.800 38.600 125.200 ;
        RECT 34.200 120.800 34.600 121.200 ;
        RECT 27.800 116.100 28.200 116.200 ;
        RECT 28.600 116.100 29.000 116.200 ;
        RECT 27.800 115.800 29.000 116.100 ;
        RECT 29.400 115.800 29.800 116.200 ;
        RECT 31.800 116.100 32.200 116.200 ;
        RECT 32.600 116.100 33.000 116.200 ;
        RECT 31.800 115.800 33.000 116.100 ;
        RECT 29.400 115.200 29.700 115.800 ;
        RECT 23.000 114.800 23.400 115.200 ;
        RECT 23.800 114.800 24.200 115.200 ;
        RECT 29.400 114.800 29.800 115.200 ;
        RECT 30.200 114.800 30.600 115.200 ;
        RECT 23.000 109.200 23.300 114.800 ;
        RECT 27.800 113.800 28.200 114.200 ;
        RECT 23.000 108.800 23.400 109.200 ;
        RECT 27.800 109.100 28.100 113.800 ;
        RECT 28.600 109.100 29.000 109.200 ;
        RECT 27.800 108.800 29.000 109.100 ;
        RECT 22.200 105.100 22.600 107.900 ;
        RECT 23.000 106.800 23.400 107.200 ;
        RECT 24.600 106.800 25.000 107.200 ;
        RECT 27.000 107.100 27.400 107.200 ;
        RECT 27.800 107.100 28.200 107.200 ;
        RECT 27.000 106.800 28.200 107.100 ;
        RECT 23.000 106.200 23.300 106.800 ;
        RECT 24.600 106.200 24.900 106.800 ;
        RECT 23.000 105.800 23.400 106.200 ;
        RECT 24.600 105.800 25.000 106.200 ;
        RECT 27.000 105.800 27.400 106.200 ;
        RECT 24.600 104.800 25.000 105.200 ;
        RECT 24.600 104.200 24.900 104.800 ;
        RECT 27.000 104.200 27.300 105.800 ;
        RECT 24.600 103.800 25.000 104.200 ;
        RECT 27.000 103.800 27.400 104.200 ;
        RECT 22.200 102.800 22.600 103.200 ;
        RECT 22.200 96.200 22.500 102.800 ;
        RECT 27.800 97.200 28.100 106.800 ;
        RECT 23.000 96.800 23.400 97.200 ;
        RECT 27.800 96.800 28.200 97.200 ;
        RECT 22.200 95.800 22.600 96.200 ;
        RECT 22.200 95.200 22.500 95.800 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 23.000 94.200 23.300 96.800 ;
        RECT 29.400 96.200 29.700 114.800 ;
        RECT 30.200 114.200 30.500 114.800 ;
        RECT 30.200 113.800 30.600 114.200 ;
        RECT 30.200 107.200 30.500 113.800 ;
        RECT 33.400 113.100 33.800 115.900 ;
        RECT 34.200 113.800 34.600 114.200 ;
        RECT 34.200 113.200 34.500 113.800 ;
        RECT 34.200 112.800 34.600 113.200 ;
        RECT 32.600 111.800 33.000 112.200 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 31.000 103.100 31.400 108.900 ;
        RECT 32.600 106.200 32.900 111.800 ;
        RECT 34.200 107.200 34.500 112.800 ;
        RECT 35.000 112.100 35.400 117.900 ;
        RECT 37.400 115.100 37.800 115.200 ;
        RECT 38.200 115.100 38.600 115.200 ;
        RECT 37.400 114.800 38.600 115.100 ;
        RECT 39.000 113.800 39.400 114.200 ;
        RECT 39.000 109.200 39.300 113.800 ;
        RECT 39.800 112.100 40.200 117.900 ;
        RECT 34.200 106.800 34.600 107.200 ;
        RECT 32.600 105.800 33.000 106.200 ;
        RECT 35.800 103.100 36.200 108.900 ;
        RECT 36.600 108.800 37.000 109.200 ;
        RECT 39.000 108.800 39.400 109.200 ;
        RECT 30.200 96.800 30.600 97.200 ;
        RECT 25.400 96.100 25.800 96.200 ;
        RECT 26.200 96.100 26.600 96.200 ;
        RECT 25.400 95.800 26.600 96.100 ;
        RECT 27.800 95.800 28.200 96.200 ;
        RECT 29.400 95.800 29.800 96.200 ;
        RECT 27.800 95.200 28.100 95.800 ;
        RECT 30.200 95.200 30.500 96.800 ;
        RECT 31.800 95.800 32.200 96.200 ;
        RECT 31.800 95.200 32.100 95.800 ;
        RECT 27.800 94.800 28.200 95.200 ;
        RECT 30.200 94.800 30.600 95.200 ;
        RECT 31.800 94.800 32.200 95.200 ;
        RECT 23.000 93.800 23.400 94.200 ;
        RECT 23.800 94.100 24.200 94.200 ;
        RECT 24.600 94.100 25.000 94.200 ;
        RECT 23.800 93.800 25.000 94.100 ;
        RECT 23.800 89.200 24.100 93.800 ;
        RECT 26.200 91.800 26.600 92.200 ;
        RECT 22.200 83.100 22.600 88.900 ;
        RECT 23.800 88.800 24.200 89.200 ;
        RECT 23.000 87.800 23.400 88.200 ;
        RECT 23.000 86.200 23.300 87.800 ;
        RECT 26.200 86.300 26.500 91.800 ;
        RECT 23.000 85.800 23.400 86.200 ;
        RECT 26.200 85.900 26.600 86.300 ;
        RECT 26.200 85.800 26.500 85.900 ;
        RECT 23.000 83.800 23.400 84.200 ;
        RECT 21.400 75.800 21.800 76.200 ;
        RECT 21.400 75.200 21.700 75.800 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 15.800 74.800 17.000 75.100 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 19.800 74.800 20.200 75.200 ;
        RECT 21.400 74.800 21.800 75.200 ;
        RECT 23.000 74.200 23.300 83.800 ;
        RECT 27.000 83.100 27.400 88.900 ;
        RECT 27.800 82.200 28.100 94.800 ;
        RECT 29.400 93.800 29.800 94.200 ;
        RECT 30.200 93.800 30.600 94.200 ;
        RECT 31.000 94.100 31.400 94.200 ;
        RECT 31.800 94.100 32.200 94.200 ;
        RECT 31.000 93.800 32.200 94.100 ;
        RECT 28.600 85.100 29.000 87.900 ;
        RECT 29.400 87.200 29.700 93.800 ;
        RECT 29.400 86.800 29.800 87.200 ;
        RECT 30.200 86.200 30.500 93.800 ;
        RECT 32.600 93.100 33.000 95.900 ;
        RECT 33.400 95.800 33.800 96.200 ;
        RECT 33.400 91.100 33.700 95.800 ;
        RECT 34.200 92.100 34.600 97.900 ;
        RECT 35.000 94.700 35.400 95.100 ;
        RECT 35.000 94.200 35.300 94.700 ;
        RECT 35.000 93.800 35.400 94.200 ;
        RECT 35.000 92.800 35.400 93.200 ;
        RECT 33.400 90.800 34.500 91.100 ;
        RECT 34.200 89.200 34.500 90.800 ;
        RECT 34.200 88.800 34.600 89.200 ;
        RECT 35.000 88.200 35.300 92.800 ;
        RECT 35.000 87.800 35.400 88.200 ;
        RECT 30.200 85.800 30.600 86.200 ;
        RECT 32.600 85.800 33.000 86.200 ;
        RECT 33.400 85.800 33.800 86.200 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 32.600 84.200 32.900 85.800 ;
        RECT 33.400 85.200 33.700 85.800 ;
        RECT 34.200 85.200 34.500 85.800 ;
        RECT 33.400 84.800 33.800 85.200 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 32.600 83.800 33.000 84.200 ;
        RECT 27.800 81.800 28.200 82.200 ;
        RECT 31.800 81.800 32.200 82.200 ;
        RECT 30.200 75.800 30.600 76.200 ;
        RECT 30.200 75.200 30.500 75.800 ;
        RECT 23.800 75.100 24.200 75.200 ;
        RECT 24.600 75.100 25.000 75.200 ;
        RECT 23.800 74.800 25.000 75.100 ;
        RECT 27.000 74.800 27.400 75.200 ;
        RECT 29.400 74.800 29.800 75.200 ;
        RECT 30.200 74.800 30.600 75.200 ;
        RECT 23.800 74.200 24.100 74.800 ;
        RECT 27.000 74.200 27.300 74.800 ;
        RECT 29.400 74.200 29.700 74.800 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 18.200 73.800 19.400 74.100 ;
        RECT 23.000 73.800 23.400 74.200 ;
        RECT 23.800 73.800 24.200 74.200 ;
        RECT 24.600 74.100 25.000 74.200 ;
        RECT 25.400 74.100 25.800 74.200 ;
        RECT 24.600 73.800 25.800 74.100 ;
        RECT 27.000 73.800 27.400 74.200 ;
        RECT 29.400 73.800 29.800 74.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 28.600 72.800 29.000 73.200 ;
        RECT 17.400 70.200 17.700 72.800 ;
        RECT 25.400 71.800 25.800 72.200 ;
        RECT 17.400 69.800 17.800 70.200 ;
        RECT 19.800 69.800 20.200 70.200 ;
        RECT 19.800 69.200 20.100 69.800 ;
        RECT 15.000 66.800 15.400 67.200 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 17.400 63.100 17.800 68.900 ;
        RECT 19.800 68.800 20.200 69.200 ;
        RECT 20.600 65.100 21.000 67.900 ;
        RECT 21.400 67.800 21.800 68.200 ;
        RECT 21.400 67.200 21.700 67.800 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 22.200 63.100 22.600 68.900 ;
        RECT 25.400 66.200 25.700 71.800 ;
        RECT 25.400 65.800 25.800 66.200 ;
        RECT 26.200 65.800 26.600 66.200 ;
        RECT 14.200 58.100 14.600 58.200 ;
        RECT 15.000 58.100 15.400 58.200 ;
        RECT 12.600 52.100 13.000 57.900 ;
        RECT 14.200 57.800 15.400 58.100 ;
        RECT 15.800 53.100 16.200 55.900 ;
        RECT 16.600 53.800 17.000 54.200 ;
        RECT 9.400 49.800 9.800 50.200 ;
        RECT 11.800 49.800 12.200 50.200 ;
        RECT 3.800 48.800 4.200 49.200 ;
        RECT 9.400 47.200 9.700 49.800 ;
        RECT 10.200 48.800 10.600 49.200 ;
        RECT 10.200 47.200 10.500 48.800 ;
        RECT 15.000 47.800 15.400 48.200 ;
        RECT 15.000 47.200 15.300 47.800 ;
        RECT 9.400 46.800 9.800 47.200 ;
        RECT 10.200 46.800 10.600 47.200 ;
        RECT 15.000 46.800 15.400 47.200 ;
        RECT 2.200 45.800 2.600 46.200 ;
        RECT 11.800 45.800 12.200 46.200 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 15.000 46.100 15.400 46.200 ;
        RECT 14.200 45.800 15.400 46.100 ;
        RECT 2.200 44.200 2.500 45.800 ;
        RECT 11.800 45.200 12.100 45.800 ;
        RECT 11.800 44.800 12.200 45.200 ;
        RECT 14.200 45.100 14.600 45.200 ;
        RECT 15.000 45.100 15.400 45.200 ;
        RECT 15.800 45.100 16.200 47.900 ;
        RECT 16.600 47.200 16.900 53.800 ;
        RECT 17.400 52.100 17.800 57.900 ;
        RECT 19.000 54.800 19.400 55.200 ;
        RECT 19.000 54.200 19.300 54.800 ;
        RECT 19.000 53.800 19.400 54.200 ;
        RECT 22.200 52.100 22.600 57.900 ;
        RECT 25.400 56.800 25.800 57.200 ;
        RECT 25.400 55.200 25.700 56.800 ;
        RECT 25.400 54.800 25.800 55.200 ;
        RECT 25.400 54.200 25.700 54.800 ;
        RECT 25.400 53.800 25.800 54.200 ;
        RECT 23.800 49.100 24.200 49.200 ;
        RECT 24.600 49.100 25.000 49.200 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 14.200 44.800 15.400 45.100 ;
        RECT 2.200 43.800 2.600 44.200 ;
        RECT 12.600 42.800 13.000 43.200 ;
        RECT 3.800 41.800 4.200 42.200 ;
        RECT 0.600 33.100 1.000 35.900 ;
        RECT 2.200 32.100 2.600 37.900 ;
        RECT 3.000 34.700 3.400 35.100 ;
        RECT 2.200 29.800 2.600 30.200 ;
        RECT 0.600 27.100 1.000 27.200 ;
        RECT 1.400 27.100 1.800 27.200 ;
        RECT 0.600 26.800 1.800 27.100 ;
        RECT 2.200 25.200 2.500 29.800 ;
        RECT 3.000 29.200 3.300 34.700 ;
        RECT 3.800 34.200 4.100 41.800 ;
        RECT 12.600 39.200 12.900 42.800 ;
        RECT 12.600 38.800 13.000 39.200 ;
        RECT 15.800 38.800 16.200 39.200 ;
        RECT 5.400 36.800 5.800 37.200 ;
        RECT 3.800 33.800 4.200 34.200 ;
        RECT 3.800 33.200 4.100 33.800 ;
        RECT 3.800 32.800 4.200 33.200 ;
        RECT 4.600 29.800 5.000 30.200 ;
        RECT 3.000 28.800 3.400 29.200 ;
        RECT 4.600 26.200 4.900 29.800 ;
        RECT 5.400 27.200 5.700 36.800 ;
        RECT 7.000 32.100 7.400 37.900 ;
        RECT 15.000 36.800 15.400 37.200 ;
        RECT 10.200 35.800 10.600 36.200 ;
        RECT 7.800 32.800 8.200 33.200 ;
        RECT 6.200 28.800 6.600 29.200 ;
        RECT 6.200 27.200 6.500 28.800 ;
        RECT 7.800 27.200 8.100 32.800 ;
        RECT 5.400 26.800 5.800 27.200 ;
        RECT 6.200 26.800 6.600 27.200 ;
        RECT 7.800 26.800 8.200 27.200 ;
        RECT 10.200 26.200 10.500 35.800 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 13.400 35.100 13.800 35.200 ;
        RECT 12.600 34.800 13.800 35.100 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 14.200 34.200 14.500 34.800 ;
        RECT 15.000 34.200 15.300 36.800 ;
        RECT 15.800 35.200 16.100 38.800 ;
        RECT 15.800 34.800 16.200 35.200 ;
        RECT 14.200 33.800 14.600 34.200 ;
        RECT 15.000 33.800 15.400 34.200 ;
        RECT 11.000 27.800 11.400 28.200 ;
        RECT 11.000 27.200 11.300 27.800 ;
        RECT 11.000 26.800 11.400 27.200 ;
        RECT 4.600 25.800 5.000 26.200 ;
        RECT 7.800 25.800 8.200 26.200 ;
        RECT 10.200 25.800 10.600 26.200 ;
        RECT 7.800 25.200 8.100 25.800 ;
        RECT 2.200 24.800 2.600 25.200 ;
        RECT 7.800 24.800 8.200 25.200 ;
        RECT 10.200 25.100 10.600 25.200 ;
        RECT 11.000 25.100 11.400 25.200 ;
        RECT 11.800 25.100 12.200 27.900 ;
        RECT 10.200 24.800 11.400 25.100 ;
        RECT 13.400 23.100 13.800 28.900 ;
        RECT 14.200 25.900 14.600 26.300 ;
        RECT 14.200 25.200 14.500 25.900 ;
        RECT 14.200 24.800 14.600 25.200 ;
        RECT 0.600 16.800 1.000 17.200 ;
        RECT 0.600 15.200 0.900 16.800 ;
        RECT 0.600 14.800 1.000 15.200 ;
        RECT 3.000 12.100 3.400 17.900 ;
        RECT 7.000 15.800 7.400 16.200 ;
        RECT 7.000 15.100 7.300 15.800 ;
        RECT 7.000 14.700 7.400 15.100 ;
        RECT 7.000 12.800 7.400 13.200 ;
        RECT 7.000 7.200 7.300 12.800 ;
        RECT 7.800 12.100 8.200 17.900 ;
        RECT 15.000 16.200 15.300 33.800 ;
        RECT 16.600 27.200 16.900 46.800 ;
        RECT 17.400 43.100 17.800 48.900 ;
        RECT 18.200 45.900 18.600 46.300 ;
        RECT 18.200 45.200 18.500 45.900 ;
        RECT 18.200 44.800 18.600 45.200 ;
        RECT 22.200 43.100 22.600 48.900 ;
        RECT 23.800 48.800 25.000 49.100 ;
        RECT 25.400 45.800 25.800 46.200 ;
        RECT 18.200 38.800 18.600 39.200 ;
        RECT 18.200 36.200 18.500 38.800 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 19.800 34.800 20.200 35.200 ;
        RECT 19.800 34.200 20.100 34.800 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 18.200 34.100 18.600 34.200 ;
        RECT 17.400 33.800 18.600 34.100 ;
        RECT 19.800 33.800 20.200 34.200 ;
        RECT 20.600 33.100 21.000 35.900 ;
        RECT 21.400 33.800 21.800 34.200 ;
        RECT 21.400 33.200 21.700 33.800 ;
        RECT 21.400 32.800 21.800 33.200 ;
        RECT 22.200 32.100 22.600 37.900 ;
        RECT 25.400 35.200 25.700 45.800 ;
        RECT 23.000 34.700 23.400 35.100 ;
        RECT 25.400 34.800 25.800 35.200 ;
        RECT 23.000 34.200 23.300 34.700 ;
        RECT 23.000 33.800 23.400 34.200 ;
        RECT 24.600 32.800 25.000 33.200 ;
        RECT 20.600 30.800 21.000 31.200 ;
        RECT 20.600 29.200 20.900 30.800 ;
        RECT 19.800 29.100 20.200 29.200 ;
        RECT 20.600 29.100 21.000 29.200 ;
        RECT 16.600 26.800 17.000 27.200 ;
        RECT 17.400 25.800 17.800 26.200 ;
        RECT 17.400 22.200 17.700 25.800 ;
        RECT 18.200 23.100 18.600 28.900 ;
        RECT 19.800 28.800 21.000 29.100 ;
        RECT 21.400 25.100 21.800 27.900 ;
        RECT 23.000 23.100 23.400 28.900 ;
        RECT 24.600 26.200 24.900 32.800 ;
        RECT 26.200 26.200 26.500 65.800 ;
        RECT 27.000 63.100 27.400 68.900 ;
        RECT 28.600 64.100 28.900 72.800 ;
        RECT 29.400 69.200 29.700 73.800 ;
        RECT 29.400 68.800 29.800 69.200 ;
        RECT 31.800 68.200 32.100 81.800 ;
        RECT 34.200 76.800 34.600 77.200 ;
        RECT 35.000 77.100 35.300 87.800 ;
        RECT 35.800 86.800 36.200 87.200 ;
        RECT 35.800 86.200 36.100 86.800 ;
        RECT 36.600 86.200 36.900 108.800 ;
        RECT 37.400 105.100 37.800 107.900 ;
        RECT 41.400 102.200 41.700 134.800 ;
        RECT 43.000 134.200 43.300 134.800 ;
        RECT 43.000 133.800 43.400 134.200 ;
        RECT 44.600 133.800 45.000 134.200 ;
        RECT 43.000 132.800 43.400 133.200 ;
        RECT 43.000 127.200 43.300 132.800 ;
        RECT 44.600 131.200 44.900 133.800 ;
        RECT 45.400 132.200 45.700 134.800 ;
        RECT 51.000 133.200 51.300 134.800 ;
        RECT 51.800 134.200 52.100 134.800 ;
        RECT 51.800 133.800 52.200 134.200 ;
        RECT 52.600 133.800 53.000 134.200 ;
        RECT 51.000 132.800 51.400 133.200 ;
        RECT 52.600 132.200 52.900 133.800 ;
        RECT 45.400 131.800 45.800 132.200 ;
        RECT 52.600 131.800 53.000 132.200 ;
        RECT 52.600 131.200 52.900 131.800 ;
        RECT 44.600 130.800 45.000 131.200 ;
        RECT 52.600 130.800 53.000 131.200 ;
        RECT 53.400 130.200 53.700 141.800 ;
        RECT 63.000 138.200 63.300 141.800 ;
        RECT 66.200 140.800 66.600 141.200 ;
        RECT 54.200 132.800 54.600 133.200 ;
        RECT 53.400 129.800 53.800 130.200 ;
        RECT 43.800 128.800 44.200 129.200 ;
        RECT 45.400 128.800 45.800 129.200 ;
        RECT 48.600 128.800 49.000 129.200 ;
        RECT 43.800 128.200 44.100 128.800 ;
        RECT 45.400 128.200 45.700 128.800 ;
        RECT 43.800 127.800 44.200 128.200 ;
        RECT 44.600 127.800 45.000 128.200 ;
        RECT 45.400 127.800 45.800 128.200 ;
        RECT 42.200 126.800 42.600 127.200 ;
        RECT 43.000 126.800 43.400 127.200 ;
        RECT 42.200 126.200 42.500 126.800 ;
        RECT 44.600 126.200 44.900 127.800 ;
        RECT 47.000 126.800 47.400 127.200 ;
        RECT 42.200 125.800 42.600 126.200 ;
        RECT 43.000 125.800 43.400 126.200 ;
        RECT 44.600 125.800 45.000 126.200 ;
        RECT 46.200 125.800 46.600 126.200 ;
        RECT 43.000 124.200 43.300 125.800 ;
        RECT 46.200 125.200 46.500 125.800 ;
        RECT 46.200 124.800 46.600 125.200 ;
        RECT 47.000 124.200 47.300 126.800 ;
        RECT 48.600 126.200 48.900 128.800 ;
        RECT 49.400 126.800 49.800 127.200 ;
        RECT 49.400 126.200 49.700 126.800 ;
        RECT 48.600 125.800 49.000 126.200 ;
        RECT 49.400 125.800 49.800 126.200 ;
        RECT 43.000 123.800 43.400 124.200 ;
        RECT 47.000 123.800 47.400 124.200 ;
        RECT 49.400 123.200 49.700 125.800 ;
        RECT 46.200 122.800 46.600 123.200 ;
        RECT 49.400 122.800 49.800 123.200 ;
        RECT 52.600 123.100 53.000 128.900 ;
        RECT 43.000 116.100 43.400 116.200 ;
        RECT 43.800 116.100 44.200 116.200 ;
        RECT 43.000 115.800 44.200 116.100 ;
        RECT 45.400 115.800 45.800 116.200 ;
        RECT 43.000 115.100 43.400 115.200 ;
        RECT 43.800 115.100 44.200 115.200 ;
        RECT 43.000 114.800 44.200 115.100 ;
        RECT 44.600 114.800 45.000 115.200 ;
        RECT 44.600 113.200 44.900 114.800 ;
        RECT 44.600 112.800 45.000 113.200 ;
        RECT 42.200 111.800 42.600 112.200 ;
        RECT 42.200 107.200 42.500 111.800 ;
        RECT 45.400 109.200 45.700 115.800 ;
        RECT 46.200 114.200 46.500 122.800 ;
        RECT 47.800 117.100 48.200 117.200 ;
        RECT 48.600 117.100 49.000 117.200 ;
        RECT 47.800 116.800 49.000 117.100 ;
        RECT 46.200 113.800 46.600 114.200 ;
        RECT 46.200 112.800 46.600 113.200 ;
        RECT 45.400 108.800 45.800 109.200 ;
        RECT 42.200 106.800 42.600 107.200 ;
        RECT 43.800 105.800 44.200 106.200 ;
        RECT 41.400 101.800 41.800 102.200 ;
        RECT 38.200 93.800 38.600 94.200 ;
        RECT 38.200 93.200 38.500 93.800 ;
        RECT 38.200 92.800 38.600 93.200 ;
        RECT 38.200 91.800 38.600 92.200 ;
        RECT 39.000 92.100 39.400 97.900 ;
        RECT 42.200 95.800 42.600 96.200 ;
        RECT 40.600 92.100 41.000 92.200 ;
        RECT 41.400 92.100 41.800 92.200 ;
        RECT 40.600 91.800 41.800 92.100 ;
        RECT 38.200 86.200 38.500 91.800 ;
        RECT 42.200 89.200 42.500 95.800 ;
        RECT 43.800 95.200 44.100 105.800 ;
        RECT 45.400 105.100 45.800 105.200 ;
        RECT 46.200 105.100 46.500 112.800 ;
        RECT 50.200 112.100 50.600 117.900 ;
        RECT 53.400 115.800 53.800 116.200 ;
        RECT 53.400 115.200 53.700 115.800 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 54.200 114.200 54.500 132.800 ;
        RECT 55.000 132.100 55.400 137.900 ;
        RECT 58.200 134.800 58.600 135.200 ;
        RECT 58.200 129.200 58.500 134.800 ;
        RECT 59.800 132.100 60.200 137.900 ;
        RECT 63.000 137.800 63.400 138.200 ;
        RECT 64.600 136.800 65.000 137.200 ;
        RECT 60.600 133.800 61.000 134.200 ;
        RECT 60.600 133.200 60.900 133.800 ;
        RECT 60.600 132.800 61.000 133.200 ;
        RECT 61.400 133.100 61.800 135.900 ;
        RECT 62.200 135.100 62.600 135.200 ;
        RECT 63.000 135.100 63.400 135.200 ;
        RECT 62.200 134.800 63.400 135.100 ;
        RECT 64.600 134.200 64.900 136.800 ;
        RECT 66.200 135.200 66.500 140.800 ;
        RECT 67.800 138.800 68.200 139.200 ;
        RECT 67.800 136.200 68.100 138.800 ;
        RECT 67.800 135.800 68.200 136.200 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 63.000 134.100 63.400 134.200 ;
        RECT 63.800 134.100 64.200 134.200 ;
        RECT 63.000 133.800 64.200 134.100 ;
        RECT 64.600 133.800 65.000 134.200 ;
        RECT 65.400 133.800 65.800 134.200 ;
        RECT 64.600 133.100 65.000 133.200 ;
        RECT 65.400 133.100 65.700 133.800 ;
        RECT 64.600 132.800 65.700 133.100 ;
        RECT 59.800 130.800 60.200 131.200 ;
        RECT 55.800 125.800 56.200 126.200 ;
        RECT 55.800 125.200 56.100 125.800 ;
        RECT 55.800 124.800 56.200 125.200 ;
        RECT 57.400 123.100 57.800 128.900 ;
        RECT 58.200 128.800 58.600 129.200 ;
        RECT 58.200 126.800 58.600 127.200 ;
        RECT 58.200 126.200 58.500 126.800 ;
        RECT 58.200 125.800 58.600 126.200 ;
        RECT 59.000 125.100 59.400 127.900 ;
        RECT 59.800 127.200 60.100 130.800 ;
        RECT 62.200 128.800 62.600 129.200 ;
        RECT 62.200 128.200 62.500 128.800 ;
        RECT 62.200 127.800 62.600 128.200 ;
        RECT 59.800 126.800 60.200 127.200 ;
        RECT 64.600 127.100 65.000 127.200 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 64.600 126.800 65.800 127.100 ;
        RECT 63.800 125.800 64.200 126.200 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 63.800 125.200 64.100 125.800 ;
        RECT 65.400 125.200 65.700 125.800 ;
        RECT 61.400 125.100 61.800 125.200 ;
        RECT 62.200 125.100 62.600 125.200 ;
        RECT 61.400 124.800 62.600 125.100 ;
        RECT 63.800 124.800 64.200 125.200 ;
        RECT 65.400 124.800 65.800 125.200 ;
        RECT 63.800 120.200 64.100 124.800 ;
        RECT 66.200 120.200 66.500 134.800 ;
        RECT 68.600 127.200 68.900 146.800 ;
        RECT 69.400 139.200 69.700 146.800 ;
        RECT 71.000 143.100 71.400 148.900 ;
        RECT 69.400 138.800 69.800 139.200 ;
        RECT 70.200 136.800 70.600 137.200 ;
        RECT 69.400 134.800 69.800 135.200 ;
        RECT 69.400 128.200 69.700 134.800 ;
        RECT 69.400 127.800 69.800 128.200 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 67.800 127.100 68.200 127.200 ;
        RECT 67.000 126.800 68.200 127.100 ;
        RECT 68.600 126.800 69.000 127.200 ;
        RECT 69.400 126.800 69.800 127.200 ;
        RECT 68.600 126.200 68.900 126.800 ;
        RECT 68.600 125.800 69.000 126.200 ;
        RECT 63.800 119.800 64.200 120.200 ;
        RECT 66.200 119.800 66.600 120.200 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 49.400 110.800 49.800 111.200 ;
        RECT 47.800 107.100 48.200 107.200 ;
        RECT 48.600 107.100 49.000 107.200 ;
        RECT 47.800 106.800 49.000 107.100 ;
        RECT 49.400 106.200 49.700 110.800 ;
        RECT 54.200 109.200 54.500 113.800 ;
        RECT 55.000 112.100 55.400 117.900 ;
        RECT 62.200 116.800 62.600 117.200 ;
        RECT 64.600 116.800 65.000 117.200 ;
        RECT 58.200 116.100 58.600 116.200 ;
        RECT 59.000 116.100 59.400 116.200 ;
        RECT 56.600 113.100 57.000 115.900 ;
        RECT 58.200 115.800 59.400 116.100 ;
        RECT 60.600 115.800 61.000 116.200 ;
        RECT 60.600 115.200 60.900 115.800 ;
        RECT 57.400 114.800 57.800 115.200 ;
        RECT 58.200 115.100 58.600 115.200 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 58.200 114.800 59.400 115.100 ;
        RECT 60.600 114.800 61.000 115.200 ;
        RECT 57.400 114.200 57.700 114.800 ;
        RECT 57.400 113.800 57.800 114.200 ;
        RECT 60.600 109.200 60.900 114.800 ;
        RECT 62.200 114.200 62.500 116.800 ;
        RECT 64.600 116.200 64.900 116.800 ;
        RECT 64.600 115.800 65.000 116.200 ;
        RECT 68.600 115.800 69.000 116.200 ;
        RECT 68.600 115.200 68.900 115.800 ;
        RECT 66.200 114.800 66.600 115.200 ;
        RECT 67.000 114.800 67.400 115.200 ;
        RECT 67.800 114.800 68.200 115.200 ;
        RECT 68.600 114.800 69.000 115.200 ;
        RECT 62.200 113.800 62.600 114.200 ;
        RECT 66.200 112.200 66.500 114.800 ;
        RECT 66.200 111.800 66.600 112.200 ;
        RECT 67.000 111.200 67.300 114.800 ;
        RECT 67.800 114.200 68.100 114.800 ;
        RECT 67.800 113.800 68.200 114.200 ;
        RECT 67.000 110.800 67.400 111.200 ;
        RECT 54.200 108.800 54.600 109.200 ;
        RECT 50.200 106.800 50.600 107.200 ;
        RECT 55.000 107.100 55.400 107.200 ;
        RECT 55.800 107.100 56.200 107.200 ;
        RECT 55.000 106.800 56.200 107.100 ;
        RECT 50.200 106.200 50.500 106.800 ;
        RECT 49.400 105.800 49.800 106.200 ;
        RECT 50.200 105.800 50.600 106.200 ;
        RECT 45.400 104.800 46.500 105.100 ;
        RECT 45.400 97.200 45.700 104.800 ;
        RECT 55.800 103.800 56.200 104.200 ;
        RECT 51.000 101.800 51.400 102.200 ;
        RECT 47.000 99.100 47.400 99.200 ;
        RECT 47.800 99.100 48.200 99.200 ;
        RECT 47.000 98.800 48.200 99.100 ;
        RECT 45.400 96.800 45.800 97.200 ;
        RECT 51.000 95.200 51.300 101.800 ;
        RECT 43.800 94.800 44.200 95.200 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 46.200 94.800 46.600 95.200 ;
        RECT 51.000 94.800 51.400 95.200 ;
        RECT 43.000 93.800 43.400 94.200 ;
        RECT 43.000 92.200 43.300 93.800 ;
        RECT 43.000 91.800 43.400 92.200 ;
        RECT 41.400 88.800 41.800 89.200 ;
        RECT 42.200 88.800 42.600 89.200 ;
        RECT 41.400 87.200 41.700 88.800 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 41.400 86.800 41.800 87.200 ;
        RECT 40.600 86.200 40.900 86.800 ;
        RECT 35.800 85.800 36.200 86.200 ;
        RECT 36.600 85.800 37.000 86.200 ;
        RECT 37.400 86.100 37.800 86.200 ;
        RECT 38.200 86.100 38.600 86.200 ;
        RECT 37.400 85.800 38.600 86.100 ;
        RECT 40.600 85.800 41.000 86.200 ;
        RECT 36.600 79.200 36.900 85.800 ;
        RECT 43.800 85.200 44.100 94.800 ;
        RECT 44.600 93.800 45.000 94.200 ;
        RECT 44.600 87.200 44.900 93.800 ;
        RECT 45.400 91.200 45.700 94.800 ;
        RECT 46.200 93.200 46.500 94.800 ;
        RECT 46.200 92.800 46.600 93.200 ;
        RECT 51.800 93.100 52.200 95.900 ;
        RECT 52.600 94.800 53.000 95.200 ;
        RECT 52.600 94.200 52.900 94.800 ;
        RECT 52.600 93.800 53.000 94.200 ;
        RECT 49.400 91.800 49.800 92.200 ;
        RECT 53.400 92.100 53.800 97.900 ;
        RECT 55.000 96.800 55.400 97.200 ;
        RECT 55.000 95.200 55.300 96.800 ;
        RECT 55.000 94.800 55.400 95.200 ;
        RECT 45.400 90.800 45.800 91.200 ;
        RECT 45.400 88.800 45.800 89.200 ;
        RECT 45.400 88.200 45.700 88.800 ;
        RECT 45.400 87.800 45.800 88.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 43.800 84.800 44.200 85.200 ;
        RECT 44.600 83.800 45.000 84.200 ;
        RECT 36.600 78.800 37.000 79.200 ;
        RECT 35.000 76.800 36.100 77.100 ;
        RECT 32.600 76.100 33.000 76.200 ;
        RECT 33.400 76.100 33.800 76.200 ;
        RECT 32.600 75.800 33.800 76.100 ;
        RECT 32.600 74.800 33.000 75.200 ;
        RECT 32.600 74.200 32.900 74.800 ;
        RECT 34.200 74.200 34.500 76.800 ;
        RECT 32.600 73.800 33.000 74.200 ;
        RECT 34.200 73.800 34.600 74.200 ;
        RECT 35.000 73.100 35.400 75.900 ;
        RECT 35.800 74.200 36.100 76.800 ;
        RECT 35.800 73.800 36.200 74.200 ;
        RECT 36.600 72.100 37.000 77.900 ;
        RECT 37.400 74.700 37.800 75.100 ;
        RECT 37.400 74.200 37.700 74.700 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 41.400 72.100 41.800 77.900 ;
        RECT 43.000 77.100 43.400 77.200 ;
        RECT 43.800 77.100 44.200 77.200 ;
        RECT 43.000 76.800 44.200 77.100 ;
        RECT 44.600 75.200 44.900 83.800 ;
        RECT 47.800 83.100 48.200 88.900 ;
        RECT 49.400 86.200 49.700 91.800 ;
        RECT 49.400 85.800 49.800 86.200 ;
        RECT 52.600 83.100 53.000 88.900 ;
        RECT 55.800 88.200 56.100 103.800 ;
        RECT 56.600 103.100 57.000 108.900 ;
        RECT 59.000 108.800 59.400 109.200 ;
        RECT 60.600 108.800 61.000 109.200 ;
        RECT 59.000 107.200 59.300 108.800 ;
        RECT 59.000 106.800 59.400 107.200 ;
        RECT 60.600 105.900 61.000 106.300 ;
        RECT 60.600 105.200 60.900 105.900 ;
        RECT 60.600 104.800 61.000 105.200 ;
        RECT 61.400 103.100 61.800 108.900 ;
        RECT 63.000 105.100 63.400 107.900 ;
        RECT 69.400 107.200 69.700 126.800 ;
        RECT 70.200 119.200 70.500 136.800 ;
        RECT 71.000 136.100 71.400 136.200 ;
        RECT 71.800 136.100 72.100 159.800 ;
        RECT 74.200 159.200 74.500 165.800 ;
        RECT 74.200 158.800 74.600 159.200 ;
        RECT 75.800 156.200 76.100 167.800 ;
        RECT 78.200 167.200 78.500 167.800 ;
        RECT 78.200 166.800 78.600 167.200 ;
        RECT 79.800 166.200 80.100 173.800 ;
        RECT 80.600 172.100 81.000 177.900 ;
        RECT 81.400 174.700 81.800 175.100 ;
        RECT 81.400 167.200 81.700 174.700 ;
        RECT 83.800 171.800 84.200 172.200 ;
        RECT 85.400 172.100 85.800 177.900 ;
        RECT 88.600 173.800 89.000 174.200 ;
        RECT 88.600 173.200 88.900 173.800 ;
        RECT 88.600 172.800 89.000 173.200 ;
        RECT 87.000 172.100 87.400 172.200 ;
        RECT 87.800 172.100 88.200 172.200 ;
        RECT 87.000 171.800 88.200 172.100 ;
        RECT 83.800 167.200 84.100 171.800 ;
        RECT 84.600 170.800 85.000 171.200 ;
        RECT 84.600 167.200 84.900 170.800 ;
        RECT 87.000 169.800 87.400 170.200 ;
        RECT 81.400 166.800 81.800 167.200 ;
        RECT 83.800 166.800 84.200 167.200 ;
        RECT 84.600 166.800 85.000 167.200 ;
        RECT 85.400 167.100 85.800 167.200 ;
        RECT 86.200 167.100 86.600 167.200 ;
        RECT 85.400 166.800 86.600 167.100 ;
        RECT 87.000 166.200 87.300 169.800 ;
        RECT 87.800 168.800 88.200 169.200 ;
        RECT 87.800 168.200 88.100 168.800 ;
        RECT 87.800 167.800 88.200 168.200 ;
        RECT 76.600 165.800 77.000 166.200 ;
        RECT 77.400 165.800 77.800 166.200 ;
        RECT 79.000 165.800 79.400 166.200 ;
        RECT 79.800 165.800 80.200 166.200 ;
        RECT 83.800 165.800 84.200 166.200 ;
        RECT 87.000 165.800 87.400 166.200 ;
        RECT 76.600 159.200 76.900 165.800 ;
        RECT 76.600 158.800 77.000 159.200 ;
        RECT 75.800 155.800 76.200 156.200 ;
        RECT 75.800 154.200 76.100 155.800 ;
        RECT 77.400 155.200 77.700 165.800 ;
        RECT 79.000 165.200 79.300 165.800 ;
        RECT 83.800 165.200 84.100 165.800 ;
        RECT 79.000 164.800 79.400 165.200 ;
        RECT 81.400 164.800 81.800 165.200 ;
        RECT 83.800 164.800 84.200 165.200 ;
        RECT 79.000 158.800 79.400 159.200 ;
        RECT 78.200 155.800 78.600 156.200 ;
        RECT 78.200 155.200 78.500 155.800 ;
        RECT 79.000 155.200 79.300 158.800 ;
        RECT 81.400 158.200 81.700 164.800 ;
        RECT 89.400 164.200 89.700 184.800 ;
        RECT 92.600 182.200 92.900 184.800 ;
        RECT 95.000 182.200 95.300 185.800 ;
        RECT 92.600 181.800 93.000 182.200 ;
        RECT 95.000 181.800 95.400 182.200 ;
        RECT 98.200 181.800 98.600 182.200 ;
        RECT 91.800 177.800 92.200 178.200 ;
        RECT 91.800 175.200 92.100 177.800 ;
        RECT 98.200 176.200 98.500 181.800 ;
        RECT 101.400 176.200 101.700 185.800 ;
        RECT 98.200 175.800 98.600 176.200 ;
        RECT 101.400 175.800 101.800 176.200 ;
        RECT 91.800 174.800 92.200 175.200 ;
        RECT 92.600 174.800 93.000 175.200 ;
        RECT 94.200 174.800 94.600 175.200 ;
        RECT 95.800 175.100 96.200 175.200 ;
        RECT 96.600 175.100 97.000 175.200 ;
        RECT 95.800 174.800 97.000 175.100 ;
        RECT 97.400 174.800 97.800 175.200 ;
        RECT 100.600 174.800 101.000 175.200 ;
        RECT 84.600 163.800 85.000 164.200 ;
        RECT 89.400 163.800 89.800 164.200 ;
        RECT 84.600 163.200 84.900 163.800 ;
        RECT 84.600 162.800 85.000 163.200 ;
        RECT 90.200 163.100 90.600 168.900 ;
        RECT 92.600 167.200 92.900 174.800 ;
        RECT 94.200 173.200 94.500 174.800 ;
        RECT 97.400 174.200 97.700 174.800 ;
        RECT 97.400 173.800 97.800 174.200 ;
        RECT 98.200 173.800 98.600 174.200 ;
        RECT 94.200 172.800 94.600 173.200 ;
        RECT 97.400 172.200 97.700 173.800 ;
        RECT 98.200 173.200 98.500 173.800 ;
        RECT 98.200 172.800 98.600 173.200 ;
        RECT 95.000 171.800 95.400 172.200 ;
        RECT 97.400 171.800 97.800 172.200 ;
        RECT 95.000 170.200 95.300 171.800 ;
        RECT 95.000 169.800 95.400 170.200 ;
        RECT 92.600 166.800 93.000 167.200 ;
        RECT 93.400 166.100 93.800 166.200 ;
        RECT 94.200 166.100 94.600 166.300 ;
        RECT 93.400 165.900 94.600 166.100 ;
        RECT 93.400 165.800 94.500 165.900 ;
        RECT 95.000 163.100 95.400 168.900 ;
        RECT 95.800 168.800 96.200 169.200 ;
        RECT 95.800 167.200 96.100 168.800 ;
        RECT 100.600 168.200 100.900 174.800 ;
        RECT 102.200 170.200 102.500 204.800 ;
        RECT 104.600 204.200 104.900 205.800 ;
        RECT 104.600 203.800 105.000 204.200 ;
        RECT 103.000 202.800 103.400 203.200 ;
        RECT 105.400 203.100 105.800 208.900 ;
        RECT 107.800 206.200 108.100 209.800 ;
        RECT 111.800 209.100 112.100 213.800 ;
        RECT 113.400 211.200 113.700 231.800 ;
        RECT 119.000 229.200 119.300 231.800 ;
        RECT 121.400 229.200 121.700 235.800 ;
        RECT 123.000 232.100 123.400 237.900 ;
        RECT 126.200 236.800 126.600 237.200 ;
        RECT 126.200 234.200 126.500 236.800 ;
        RECT 127.800 236.100 128.200 236.200 ;
        RECT 128.600 236.100 129.000 236.200 ;
        RECT 127.800 235.800 129.000 236.100 ;
        RECT 130.200 235.800 130.600 236.200 ;
        RECT 132.600 235.800 133.000 236.200 ;
        RECT 134.200 236.100 134.600 236.200 ;
        RECT 135.000 236.100 135.400 236.200 ;
        RECT 134.200 235.800 135.400 236.100 ;
        RECT 127.800 235.200 128.100 235.800 ;
        RECT 130.200 235.200 130.500 235.800 ;
        RECT 132.600 235.200 132.900 235.800 ;
        RECT 127.800 234.800 128.200 235.200 ;
        RECT 130.200 234.800 130.600 235.200 ;
        RECT 132.600 234.800 133.000 235.200 ;
        RECT 126.200 233.800 126.600 234.200 ;
        RECT 127.800 234.100 128.200 234.200 ;
        RECT 128.600 234.100 129.000 234.200 ;
        RECT 127.800 233.800 129.000 234.100 ;
        RECT 124.600 232.800 125.000 233.200 ;
        RECT 123.000 230.800 123.400 231.200 ;
        RECT 115.000 228.800 115.400 229.200 ;
        RECT 119.000 228.800 119.400 229.200 ;
        RECT 120.600 228.800 121.000 229.200 ;
        RECT 121.400 228.800 121.800 229.200 ;
        RECT 115.000 227.200 115.300 228.800 ;
        RECT 115.800 227.800 116.200 228.200 ;
        RECT 115.000 226.800 115.400 227.200 ;
        RECT 115.000 225.800 115.400 226.200 ;
        RECT 114.200 221.800 114.600 222.200 ;
        RECT 114.200 215.200 114.500 221.800 ;
        RECT 114.200 214.800 114.600 215.200 ;
        RECT 115.000 213.200 115.300 225.800 ;
        RECT 115.800 222.200 116.100 227.800 ;
        RECT 119.800 226.800 120.200 227.200 ;
        RECT 119.800 226.200 120.100 226.800 ;
        RECT 120.600 226.200 120.900 228.800 ;
        RECT 123.000 227.200 123.300 230.800 ;
        RECT 123.000 226.800 123.400 227.200 ;
        RECT 123.800 226.800 124.200 227.200 ;
        RECT 117.400 226.100 117.800 226.200 ;
        RECT 118.200 226.100 118.600 226.200 ;
        RECT 117.400 225.800 118.600 226.100 ;
        RECT 119.800 225.800 120.200 226.200 ;
        RECT 120.600 225.800 121.000 226.200 ;
        RECT 121.400 224.800 121.800 225.200 ;
        RECT 116.600 223.800 117.000 224.200 ;
        RECT 115.800 221.800 116.200 222.200 ;
        RECT 116.600 221.200 116.900 223.800 ;
        RECT 120.600 222.800 121.000 223.200 ;
        RECT 116.600 220.800 117.000 221.200 ;
        RECT 115.000 212.800 115.400 213.200 ;
        RECT 115.800 212.100 116.200 217.900 ;
        RECT 116.600 214.200 116.900 220.800 ;
        RECT 120.600 219.200 120.900 222.800 ;
        RECT 121.400 222.200 121.700 224.800 ;
        RECT 121.400 221.800 121.800 222.200 ;
        RECT 120.600 218.800 121.000 219.200 ;
        RECT 116.600 213.800 117.000 214.200 ;
        RECT 117.400 213.100 117.800 215.900 ;
        RECT 122.200 214.800 122.600 215.200 ;
        RECT 119.000 213.800 119.400 214.200 ;
        RECT 113.400 210.800 113.800 211.200 ;
        RECT 117.400 210.800 117.800 211.200 ;
        RECT 107.800 205.800 108.200 206.200 ;
        RECT 110.200 203.100 110.600 208.900 ;
        RECT 111.000 208.800 112.100 209.100 ;
        RECT 111.000 207.200 111.300 208.800 ;
        RECT 111.000 206.800 111.400 207.200 ;
        RECT 103.000 199.200 103.300 202.800 ;
        RECT 103.000 198.800 103.400 199.200 ;
        RECT 105.400 192.100 105.800 197.900 ;
        RECT 107.800 195.100 108.200 195.200 ;
        RECT 108.600 195.100 109.000 195.200 ;
        RECT 107.800 194.800 109.000 195.100 ;
        RECT 106.200 193.800 106.600 194.200 ;
        RECT 106.200 193.200 106.500 193.800 ;
        RECT 106.200 192.800 106.600 193.200 ;
        RECT 110.200 192.100 110.600 197.900 ;
        RECT 111.000 195.200 111.300 206.800 ;
        RECT 111.800 205.100 112.200 207.900 ;
        RECT 115.800 207.800 116.200 208.200 ;
        RECT 115.800 206.200 116.100 207.800 ;
        RECT 117.400 206.200 117.700 210.800 ;
        RECT 119.000 209.200 119.300 213.800 ;
        RECT 119.800 211.800 120.200 212.200 ;
        RECT 119.000 208.800 119.400 209.200 ;
        RECT 119.800 206.200 120.100 211.800 ;
        RECT 122.200 209.200 122.500 214.800 ;
        RECT 123.000 212.100 123.400 217.900 ;
        RECT 122.200 208.800 122.600 209.200 ;
        RECT 123.000 208.800 123.400 209.200 ;
        RECT 123.000 208.200 123.300 208.800 ;
        RECT 123.800 208.200 124.100 226.800 ;
        RECT 124.600 218.200 124.900 232.800 ;
        RECT 126.200 231.200 126.500 233.800 ;
        RECT 130.200 232.200 130.500 234.800 ;
        RECT 131.800 233.800 132.200 234.200 ;
        RECT 130.200 231.800 130.600 232.200 ;
        RECT 126.200 230.800 126.600 231.200 ;
        RECT 131.800 229.200 132.100 233.800 ;
        RECT 128.600 228.800 129.000 229.200 ;
        RECT 128.600 228.200 128.900 228.800 ;
        RECT 127.000 227.800 127.400 228.200 ;
        RECT 128.600 227.800 129.000 228.200 ;
        RECT 127.000 226.200 127.300 227.800 ;
        RECT 127.000 225.800 127.400 226.200 ;
        RECT 127.800 225.800 128.200 226.200 ;
        RECT 127.800 223.200 128.100 225.800 ;
        RECT 127.800 222.800 128.200 223.200 ;
        RECT 131.000 223.100 131.400 228.900 ;
        RECT 131.800 228.800 132.200 229.200 ;
        RECT 132.600 225.200 132.900 234.800 ;
        RECT 136.600 233.800 137.000 234.200 ;
        RECT 134.200 231.800 134.600 232.200 ;
        RECT 134.200 230.200 134.500 231.800 ;
        RECT 136.600 230.200 136.900 233.800 ;
        RECT 137.400 233.100 137.800 235.900 ;
        RECT 139.000 232.100 139.400 237.900 ;
        RECT 142.200 234.800 142.600 235.200 ;
        RECT 140.600 233.800 141.000 234.200 ;
        RECT 134.200 229.800 134.600 230.200 ;
        RECT 136.600 229.800 137.000 230.200 ;
        RECT 135.000 225.900 135.400 226.300 ;
        RECT 135.000 225.200 135.300 225.900 ;
        RECT 132.600 224.800 133.000 225.200 ;
        RECT 135.000 224.800 135.400 225.200 ;
        RECT 135.800 223.100 136.200 228.900 ;
        RECT 138.200 228.800 138.600 229.200 ;
        RECT 136.600 226.800 137.000 227.200 ;
        RECT 136.600 224.200 136.900 226.800 ;
        RECT 137.400 225.100 137.800 227.900 ;
        RECT 138.200 227.200 138.500 228.800 ;
        RECT 138.200 226.800 138.600 227.200 ;
        RECT 138.200 226.100 138.600 226.200 ;
        RECT 139.000 226.100 139.400 226.200 ;
        RECT 138.200 225.800 139.400 226.100 ;
        RECT 140.600 225.200 140.900 233.800 ;
        RECT 142.200 228.200 142.500 234.800 ;
        RECT 143.800 232.100 144.200 237.900 ;
        RECT 161.400 236.800 161.800 237.200 ;
        RECT 159.800 235.800 160.200 236.200 ;
        RECT 159.800 235.200 160.100 235.800 ;
        RECT 147.000 234.800 147.400 235.200 ;
        RECT 147.800 234.800 148.200 235.200 ;
        RECT 151.000 235.100 151.400 235.200 ;
        RECT 151.800 235.100 152.200 235.200 ;
        RECT 151.000 234.800 152.200 235.100 ;
        RECT 155.800 234.800 156.200 235.200 ;
        RECT 156.600 235.100 157.000 235.200 ;
        RECT 157.400 235.100 157.800 235.200 ;
        RECT 156.600 234.800 157.800 235.100 ;
        RECT 159.800 234.800 160.200 235.200 ;
        RECT 147.000 234.200 147.300 234.800 ;
        RECT 147.800 234.200 148.100 234.800 ;
        RECT 147.000 233.800 147.400 234.200 ;
        RECT 147.800 233.800 148.200 234.200 ;
        RECT 146.200 231.800 146.600 232.200 ;
        RECT 144.600 230.800 145.000 231.200 ;
        RECT 141.400 227.800 141.800 228.200 ;
        RECT 142.200 227.800 142.600 228.200 ;
        RECT 141.400 227.200 141.700 227.800 ;
        RECT 141.400 226.800 141.800 227.200 ;
        RECT 144.600 226.200 144.900 230.800 ;
        RECT 146.200 226.200 146.500 231.800 ;
        RECT 147.000 229.800 147.400 230.200 ;
        RECT 147.000 226.200 147.300 229.800 ;
        RECT 147.800 227.200 148.100 233.800 ;
        RECT 153.400 232.800 153.800 233.200 ;
        RECT 148.600 231.800 149.000 232.200 ;
        RECT 148.600 231.200 148.900 231.800 ;
        RECT 148.600 230.800 149.000 231.200 ;
        RECT 150.200 229.800 150.600 230.200 ;
        RECT 150.200 229.200 150.500 229.800 ;
        RECT 153.400 229.200 153.700 232.800 ;
        RECT 150.200 228.800 150.600 229.200 ;
        RECT 147.800 226.800 148.200 227.200 ;
        RECT 143.000 225.800 143.400 226.200 ;
        RECT 144.600 225.800 145.000 226.200 ;
        RECT 146.200 225.800 146.600 226.200 ;
        RECT 147.000 225.800 147.400 226.200 ;
        RECT 148.600 225.800 149.000 226.200 ;
        RECT 143.000 225.200 143.300 225.800 ;
        RECT 139.000 225.100 139.400 225.200 ;
        RECT 139.800 225.100 140.200 225.200 ;
        RECT 139.000 224.800 140.200 225.100 ;
        RECT 140.600 224.800 141.000 225.200 ;
        RECT 143.000 224.800 143.400 225.200 ;
        RECT 136.600 223.800 137.000 224.200 ;
        RECT 145.400 221.800 145.800 222.200 ;
        RECT 124.600 217.800 125.000 218.200 ;
        RECT 124.600 215.200 124.900 217.800 ;
        RECT 124.600 214.800 125.000 215.200 ;
        RECT 125.400 215.100 125.800 215.200 ;
        RECT 126.200 215.100 126.600 215.200 ;
        RECT 125.400 214.800 126.600 215.100 ;
        RECT 124.600 211.800 125.000 212.200 ;
        RECT 127.800 212.100 128.200 217.900 ;
        RECT 136.600 217.800 137.000 218.200 ;
        RECT 129.400 213.100 129.800 215.900 ;
        RECT 133.400 215.800 133.800 216.200 ;
        RECT 133.400 215.200 133.700 215.800 ;
        RECT 130.200 215.100 130.600 215.200 ;
        RECT 131.000 215.100 131.400 215.200 ;
        RECT 130.200 214.800 131.400 215.100 ;
        RECT 133.400 214.800 133.800 215.200 ;
        RECT 130.200 214.100 130.600 214.200 ;
        RECT 131.000 214.100 131.400 214.200 ;
        RECT 130.200 213.800 131.400 214.100 ;
        RECT 132.600 214.100 133.000 214.200 ;
        RECT 133.400 214.100 133.800 214.200 ;
        RECT 132.600 213.800 133.800 214.100 ;
        RECT 135.000 213.800 135.400 214.200 ;
        RECT 123.000 207.800 123.400 208.200 ;
        RECT 123.800 207.800 124.200 208.200 ;
        RECT 121.400 206.800 121.800 207.200 ;
        RECT 123.800 206.800 124.200 207.200 ;
        RECT 112.600 205.800 113.000 206.200 ;
        RECT 113.400 205.800 113.800 206.200 ;
        RECT 115.800 205.800 116.200 206.200 ;
        RECT 117.400 205.800 117.800 206.200 ;
        RECT 119.800 205.800 120.200 206.200 ;
        RECT 112.600 205.200 112.900 205.800 ;
        RECT 112.600 204.800 113.000 205.200 ;
        RECT 113.400 204.100 113.700 205.800 ;
        RECT 112.600 203.800 113.700 204.100 ;
        RECT 112.600 201.200 112.900 203.800 ;
        RECT 113.400 202.800 113.800 203.200 ;
        RECT 112.600 200.800 113.000 201.200 ;
        RECT 111.000 194.800 111.400 195.200 ;
        RECT 111.000 194.200 111.300 194.800 ;
        RECT 111.000 193.800 111.400 194.200 ;
        RECT 111.800 193.100 112.200 195.900 ;
        RECT 113.400 195.200 113.700 202.800 ;
        RECT 115.000 201.800 115.400 202.200 ;
        RECT 115.000 201.200 115.300 201.800 ;
        RECT 115.000 200.800 115.400 201.200 ;
        RECT 113.400 194.800 113.800 195.200 ;
        RECT 115.800 194.800 116.200 195.200 ;
        RECT 116.600 194.800 117.000 195.200 ;
        RECT 115.000 193.800 115.400 194.200 ;
        RECT 115.000 193.200 115.300 193.800 ;
        RECT 115.000 192.800 115.400 193.200 ;
        RECT 115.800 192.200 116.100 194.800 ;
        RECT 115.800 191.800 116.200 192.200 ;
        RECT 103.000 185.100 103.400 187.900 ;
        RECT 103.800 186.800 104.200 187.200 ;
        RECT 103.800 183.200 104.100 186.800 ;
        RECT 103.800 182.800 104.200 183.200 ;
        RECT 104.600 183.100 105.000 188.900 ;
        RECT 106.200 186.100 106.600 186.200 ;
        RECT 107.000 186.100 107.400 186.200 ;
        RECT 106.200 185.800 107.400 186.100 ;
        RECT 109.400 183.100 109.800 188.900 ;
        RECT 116.600 187.200 116.900 194.800 ;
        RECT 117.400 193.200 117.700 205.800 ;
        RECT 121.400 205.200 121.700 206.800 ;
        RECT 123.800 206.200 124.100 206.800 ;
        RECT 124.600 206.200 124.900 211.800 ;
        RECT 131.000 211.200 131.300 213.800 ;
        RECT 135.000 212.200 135.300 213.800 ;
        RECT 135.800 213.100 136.200 215.900 ;
        RECT 136.600 214.200 136.900 217.800 ;
        RECT 136.600 213.800 137.000 214.200 ;
        RECT 135.000 211.800 135.400 212.200 ;
        RECT 137.400 212.100 137.800 217.900 ;
        RECT 138.200 214.700 138.600 215.100 ;
        RECT 138.200 214.200 138.500 214.700 ;
        RECT 138.200 213.800 138.600 214.200 ;
        RECT 142.200 212.100 142.600 217.900 ;
        RECT 145.400 214.200 145.700 221.800 ;
        RECT 148.600 218.200 148.900 225.800 ;
        RECT 152.600 223.100 153.000 228.900 ;
        RECT 153.400 228.800 153.800 229.200 ;
        RECT 155.000 226.800 155.400 227.200 ;
        RECT 155.000 226.200 155.300 226.800 ;
        RECT 155.000 225.800 155.400 226.200 ;
        RECT 155.800 223.200 156.100 234.800 ;
        RECT 161.400 234.200 161.700 236.800 ;
        RECT 156.600 233.800 157.000 234.200 ;
        RECT 159.000 234.100 159.400 234.200 ;
        RECT 159.800 234.100 160.200 234.200 ;
        RECT 159.000 233.800 160.200 234.100 ;
        RECT 161.400 233.800 161.800 234.200 ;
        RECT 155.800 222.800 156.200 223.200 ;
        RECT 156.600 222.200 156.900 233.800 ;
        RECT 161.400 230.200 161.700 233.800 ;
        RECT 164.600 232.100 165.000 237.900 ;
        RECT 167.800 234.800 168.200 235.200 ;
        RECT 167.800 234.200 168.100 234.800 ;
        RECT 167.800 233.800 168.200 234.200 ;
        RECT 169.400 232.100 169.800 237.900 ;
        RECT 170.200 234.800 170.600 235.200 ;
        RECT 170.200 234.200 170.500 234.800 ;
        RECT 170.200 233.800 170.600 234.200 ;
        RECT 171.000 233.100 171.400 235.900 ;
        RECT 171.800 231.800 172.200 232.200 ;
        RECT 174.200 232.100 174.600 237.900 ;
        RECT 178.200 234.700 178.600 235.100 ;
        RECT 178.200 233.200 178.500 234.700 ;
        RECT 178.200 232.800 178.600 233.200 ;
        RECT 179.000 232.100 179.400 237.900 ;
        RECT 180.600 233.100 181.000 235.900 ;
        RECT 181.400 233.100 181.800 235.900 ;
        RECT 183.000 232.100 183.400 237.900 ;
        RECT 184.600 235.800 185.000 236.200 ;
        RECT 184.600 235.200 184.900 235.800 ;
        RECT 184.600 234.800 185.000 235.200 ;
        RECT 185.400 233.800 185.800 234.200 ;
        RECT 161.400 229.800 161.800 230.200 ;
        RECT 157.400 223.100 157.800 228.900 ;
        RECT 171.800 228.200 172.100 231.800 ;
        RECT 175.000 230.800 175.400 231.200 ;
        RECT 161.400 228.100 161.800 228.200 ;
        RECT 162.200 228.100 162.600 228.200 ;
        RECT 158.200 226.800 158.600 227.200 ;
        RECT 158.200 225.200 158.500 226.800 ;
        RECT 158.200 224.800 158.600 225.200 ;
        RECT 159.000 225.100 159.400 227.900 ;
        RECT 161.400 227.800 162.600 228.100 ;
        RECT 164.600 227.800 165.000 228.200 ;
        RECT 171.800 227.800 172.200 228.200 ;
        RECT 160.600 226.800 161.000 227.200 ;
        RECT 159.800 225.800 160.200 226.200 ;
        RECT 159.800 222.200 160.100 225.800 ;
        RECT 160.600 224.200 160.900 226.800 ;
        RECT 164.600 226.200 164.900 227.800 ;
        RECT 163.000 225.800 163.400 226.200 ;
        RECT 164.600 225.800 165.000 226.200 ;
        RECT 163.000 224.200 163.300 225.800 ;
        RECT 172.600 225.100 173.000 227.900 ;
        RECT 160.600 223.800 161.000 224.200 ;
        RECT 163.000 223.800 163.400 224.200 ;
        RECT 174.200 223.100 174.600 228.900 ;
        RECT 175.000 226.300 175.300 230.800 ;
        RECT 181.400 229.100 181.800 229.200 ;
        RECT 182.200 229.100 182.600 229.200 ;
        RECT 175.800 226.800 176.200 227.200 ;
        RECT 175.000 225.900 175.400 226.300 ;
        RECT 175.000 225.800 175.300 225.900 ;
        RECT 175.800 225.200 176.100 226.800 ;
        RECT 175.800 224.800 176.200 225.200 ;
        RECT 156.600 221.800 157.000 222.200 ;
        RECT 159.800 221.800 160.200 222.200 ;
        RECT 166.200 221.800 166.600 222.200 ;
        RECT 159.800 218.800 160.200 219.200 ;
        RECT 147.000 214.800 147.400 215.200 ;
        RECT 145.400 213.800 145.800 214.200 ;
        RECT 143.800 212.100 144.200 212.200 ;
        RECT 144.600 212.100 145.000 212.200 ;
        RECT 143.800 211.800 145.000 212.100 ;
        RECT 145.400 212.100 145.800 212.200 ;
        RECT 146.200 212.100 146.600 212.200 ;
        RECT 145.400 211.800 146.600 212.100 ;
        RECT 131.000 210.800 131.400 211.200 ;
        RECT 143.000 210.800 143.400 211.200 ;
        RECT 135.000 209.800 135.400 210.200 ;
        RECT 141.400 209.800 141.800 210.200 ;
        RECT 128.600 208.800 129.000 209.200 ;
        RECT 128.600 206.200 128.900 208.800 ;
        RECT 123.800 205.800 124.200 206.200 ;
        RECT 124.600 205.800 125.000 206.200 ;
        RECT 127.000 206.100 127.400 206.200 ;
        RECT 127.800 206.100 128.200 206.200 ;
        RECT 127.000 205.800 128.200 206.100 ;
        RECT 128.600 205.800 129.000 206.200 ;
        RECT 121.400 204.800 121.800 205.200 ;
        RECT 131.000 203.100 131.400 208.900 ;
        RECT 135.000 206.300 135.300 209.800 ;
        RECT 141.400 209.200 141.700 209.800 ;
        RECT 135.000 205.900 135.400 206.300 ;
        RECT 133.400 204.800 133.800 205.200 ;
        RECT 126.200 201.800 126.600 202.200 ;
        RECT 126.200 198.200 126.500 201.800 ;
        RECT 127.000 199.800 127.400 200.200 ;
        RECT 132.600 199.800 133.000 200.200 ;
        RECT 127.000 198.200 127.300 199.800 ;
        RECT 117.400 192.800 117.800 193.200 ;
        RECT 117.400 192.100 117.800 192.200 ;
        RECT 118.200 192.100 118.600 192.200 ;
        RECT 119.800 192.100 120.200 197.900 ;
        RECT 120.600 195.800 121.000 196.200 ;
        RECT 120.600 195.200 120.900 195.800 ;
        RECT 120.600 194.800 121.000 195.200 ;
        RECT 123.800 194.700 124.200 195.100 ;
        RECT 117.400 191.800 118.600 192.100 ;
        RECT 123.800 190.200 124.100 194.700 ;
        RECT 124.600 192.100 125.000 197.900 ;
        RECT 126.200 197.800 126.600 198.200 ;
        RECT 127.000 197.800 127.400 198.200 ;
        RECT 125.400 192.800 125.800 193.200 ;
        RECT 126.200 193.100 126.600 195.900 ;
        RECT 132.600 195.200 132.900 199.800 ;
        RECT 127.800 194.800 128.200 195.200 ;
        RECT 130.200 194.800 130.600 195.200 ;
        RECT 131.000 194.800 131.400 195.200 ;
        RECT 131.800 194.800 132.200 195.200 ;
        RECT 132.600 194.800 133.000 195.200 ;
        RECT 127.800 194.200 128.100 194.800 ;
        RECT 130.200 194.200 130.500 194.800 ;
        RECT 127.000 193.800 127.400 194.200 ;
        RECT 127.800 193.800 128.200 194.200 ;
        RECT 130.200 193.800 130.600 194.200 ;
        RECT 123.800 189.800 124.200 190.200 ;
        RECT 117.400 187.800 117.800 188.200 ;
        RECT 117.400 187.200 117.700 187.800 ;
        RECT 110.200 187.100 110.600 187.200 ;
        RECT 111.000 187.100 111.400 187.200 ;
        RECT 110.200 186.800 111.400 187.100 ;
        RECT 114.200 186.800 114.600 187.200 ;
        RECT 116.600 186.800 117.000 187.200 ;
        RECT 117.400 186.800 117.800 187.200 ;
        RECT 114.200 186.200 114.500 186.800 ;
        RECT 114.200 185.800 114.600 186.200 ;
        RECT 118.200 185.800 118.600 186.200 ;
        RECT 119.000 185.800 119.400 186.200 ;
        RECT 119.800 186.100 120.200 186.200 ;
        RECT 120.600 186.100 121.000 186.200 ;
        RECT 119.800 185.800 121.000 186.100 ;
        RECT 118.200 185.200 118.500 185.800 ;
        RECT 114.200 185.100 114.600 185.200 ;
        RECT 115.000 185.100 115.400 185.200 ;
        RECT 114.200 184.800 115.400 185.100 ;
        RECT 118.200 184.800 118.600 185.200 ;
        RECT 119.000 185.100 119.300 185.800 ;
        RECT 119.000 184.800 120.100 185.100 ;
        RECT 112.600 178.800 113.000 179.200 ;
        RECT 103.000 176.800 103.400 177.200 ;
        RECT 104.600 177.100 105.000 177.200 ;
        RECT 105.400 177.100 105.800 177.200 ;
        RECT 104.600 176.800 105.800 177.100 ;
        RECT 103.000 175.200 103.300 176.800 ;
        RECT 103.000 174.800 103.400 175.200 ;
        RECT 103.800 174.800 104.200 175.200 ;
        RECT 103.800 174.200 104.100 174.800 ;
        RECT 103.800 173.800 104.200 174.200 ;
        RECT 107.000 172.100 107.400 177.900 ;
        RECT 110.200 175.000 110.600 175.100 ;
        RECT 111.000 175.000 111.400 175.100 ;
        RECT 110.200 174.700 111.400 175.000 ;
        RECT 108.600 173.800 109.000 174.200 ;
        RECT 103.800 170.800 104.200 171.200 ;
        RECT 102.200 169.800 102.600 170.200 ;
        RECT 95.800 166.800 96.200 167.200 ;
        RECT 96.600 165.100 97.000 167.900 ;
        RECT 97.400 167.800 97.800 168.200 ;
        RECT 100.600 167.800 101.000 168.200 ;
        RECT 97.400 167.200 97.700 167.800 ;
        RECT 103.800 167.200 104.100 170.800 ;
        RECT 108.600 169.200 108.900 173.800 ;
        RECT 111.800 172.100 112.200 177.900 ;
        RECT 112.600 174.200 112.900 178.800 ;
        RECT 114.200 176.800 114.600 177.200 ;
        RECT 112.600 173.800 113.000 174.200 ;
        RECT 113.400 173.100 113.800 175.900 ;
        RECT 114.200 174.200 114.500 176.800 ;
        RECT 118.200 176.200 118.500 184.800 ;
        RECT 119.800 177.200 120.100 184.800 ;
        RECT 120.600 184.800 121.000 185.200 ;
        RECT 120.600 179.200 120.900 184.800 ;
        RECT 123.800 183.100 124.200 188.900 ;
        RECT 125.400 188.200 125.700 192.800 ;
        RECT 125.400 187.800 125.800 188.200 ;
        RECT 121.400 181.800 121.800 182.200 ;
        RECT 120.600 178.800 121.000 179.200 ;
        RECT 121.400 178.200 121.700 181.800 ;
        RECT 121.400 177.800 121.800 178.200 ;
        RECT 119.800 176.800 120.200 177.200 ;
        RECT 119.800 176.200 120.100 176.800 ;
        RECT 115.800 176.100 116.200 176.200 ;
        RECT 116.600 176.100 117.000 176.200 ;
        RECT 115.800 175.800 117.000 176.100 ;
        RECT 118.200 175.800 118.600 176.200 ;
        RECT 119.800 175.800 120.200 176.200 ;
        RECT 118.200 175.200 118.500 175.800 ;
        RECT 115.800 174.800 116.200 175.200 ;
        RECT 118.200 174.800 118.600 175.200 ;
        RECT 115.800 174.200 116.100 174.800 ;
        RECT 114.200 173.800 114.600 174.200 ;
        RECT 115.800 173.800 116.200 174.200 ;
        RECT 114.200 170.800 114.600 171.200 ;
        RECT 97.400 166.800 97.800 167.200 ;
        RECT 101.400 166.800 101.800 167.200 ;
        RECT 103.800 166.800 104.200 167.200 ;
        RECT 101.400 166.200 101.700 166.800 ;
        RECT 101.400 165.800 101.800 166.200 ;
        RECT 103.000 165.800 103.400 166.200 ;
        RECT 99.000 164.800 99.400 165.200 ;
        RECT 99.000 164.200 99.300 164.800 ;
        RECT 103.000 164.200 103.300 165.800 ;
        RECT 104.600 165.100 105.000 167.900 ;
        RECT 99.000 163.800 99.400 164.200 ;
        RECT 103.000 163.800 103.400 164.200 ;
        RECT 106.200 163.100 106.600 168.900 ;
        RECT 108.600 168.800 109.000 169.200 ;
        RECT 108.600 167.200 108.900 168.800 ;
        RECT 108.600 166.800 109.000 167.200 ;
        RECT 107.800 166.100 108.200 166.200 ;
        RECT 108.600 166.100 109.000 166.200 ;
        RECT 107.800 165.800 109.000 166.100 ;
        RECT 111.000 163.100 111.400 168.900 ;
        RECT 113.400 168.800 113.800 169.200 ;
        RECT 113.400 168.200 113.700 168.800 ;
        RECT 113.400 167.800 113.800 168.200 ;
        RECT 114.200 167.200 114.500 170.800 ;
        RECT 114.200 166.800 114.600 167.200 ;
        RECT 114.200 165.800 114.600 166.200 ;
        RECT 115.800 166.100 116.200 166.200 ;
        RECT 116.600 166.100 117.000 166.200 ;
        RECT 115.800 165.800 117.000 166.100 ;
        RECT 111.800 163.800 112.200 164.200 ;
        RECT 87.800 160.800 88.200 161.200 ;
        RECT 81.400 157.800 81.800 158.200 ;
        RECT 81.400 156.800 81.800 157.200 ;
        RECT 80.600 155.800 81.000 156.200 ;
        RECT 76.600 154.800 77.000 155.200 ;
        RECT 77.400 154.800 77.800 155.200 ;
        RECT 78.200 154.800 78.600 155.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 75.800 153.800 76.200 154.200 ;
        RECT 76.600 152.200 76.900 154.800 ;
        RECT 76.600 151.800 77.000 152.200 ;
        RECT 77.400 151.100 77.700 154.800 ;
        RECT 79.000 154.200 79.300 154.800 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 76.600 150.800 77.700 151.100 ;
        RECT 80.600 152.200 80.900 155.800 ;
        RECT 81.400 155.200 81.700 156.800 ;
        RECT 81.400 154.800 81.800 155.200 ;
        RECT 80.600 151.800 81.000 152.200 ;
        RECT 83.800 152.100 84.200 157.900 ;
        RECT 87.000 155.800 87.400 156.200 ;
        RECT 87.000 155.200 87.300 155.800 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 87.000 154.800 87.400 155.200 ;
        RECT 84.600 154.200 84.900 154.800 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 73.400 148.100 73.800 148.200 ;
        RECT 74.200 148.100 74.600 148.200 ;
        RECT 73.400 147.800 74.600 148.100 ;
        RECT 75.000 147.100 75.400 147.200 ;
        RECT 75.800 147.100 76.200 147.200 ;
        RECT 75.000 146.800 76.200 147.100 ;
        RECT 75.000 146.100 75.400 146.200 ;
        RECT 75.800 146.100 76.200 146.200 ;
        RECT 75.000 145.800 76.200 146.100 ;
        RECT 76.600 142.200 76.900 150.800 ;
        RECT 77.400 148.800 77.800 149.200 ;
        RECT 79.800 148.800 80.200 149.200 ;
        RECT 77.400 145.200 77.700 148.800 ;
        RECT 79.800 148.200 80.100 148.800 ;
        RECT 79.800 147.800 80.200 148.200 ;
        RECT 77.400 144.800 77.800 145.200 ;
        RECT 73.400 141.800 73.800 142.200 ;
        RECT 75.000 141.800 75.400 142.200 ;
        RECT 76.600 141.800 77.000 142.200 ;
        RECT 73.400 140.200 73.700 141.800 ;
        RECT 73.400 139.800 73.800 140.200 ;
        RECT 71.000 135.800 72.100 136.100 ;
        RECT 73.400 136.800 73.800 137.200 ;
        RECT 73.400 136.200 73.700 136.800 ;
        RECT 73.400 135.800 73.800 136.200 ;
        RECT 71.000 134.800 71.400 135.200 ;
        RECT 71.000 129.200 71.300 134.800 ;
        RECT 71.000 128.800 71.400 129.200 ;
        RECT 71.000 125.200 71.300 128.800 ;
        RECT 71.000 124.800 71.400 125.200 ;
        RECT 71.000 122.800 71.400 123.200 ;
        RECT 70.200 118.800 70.600 119.200 ;
        RECT 71.000 115.200 71.300 122.800 ;
        RECT 71.000 114.800 71.400 115.200 ;
        RECT 71.000 113.800 71.400 114.200 ;
        RECT 64.600 107.100 65.000 107.200 ;
        RECT 65.400 107.100 65.800 107.200 ;
        RECT 64.600 106.800 65.800 107.100 ;
        RECT 66.200 106.800 66.600 107.200 ;
        RECT 69.400 106.800 69.800 107.200 ;
        RECT 63.800 105.800 64.200 106.200 ;
        RECT 63.800 105.200 64.100 105.800 ;
        RECT 66.200 105.200 66.500 106.800 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 67.800 105.800 69.000 106.100 ;
        RECT 63.800 104.800 64.200 105.200 ;
        RECT 66.200 104.800 66.600 105.200 ;
        RECT 67.800 102.800 68.200 103.200 ;
        RECT 61.400 101.800 61.800 102.200 ;
        RECT 58.200 92.100 58.600 97.900 ;
        RECT 60.600 96.800 61.000 97.200 ;
        RECT 60.600 96.200 60.900 96.800 ;
        RECT 60.600 95.800 61.000 96.200 ;
        RECT 61.400 95.200 61.700 101.800 ;
        RECT 67.800 97.200 68.100 102.800 ;
        RECT 67.800 96.800 68.200 97.200 ;
        RECT 67.800 96.200 68.100 96.800 ;
        RECT 62.200 95.800 62.600 96.200 ;
        RECT 65.400 95.800 65.800 96.200 ;
        RECT 67.800 95.800 68.200 96.200 ;
        RECT 68.600 95.800 69.000 96.200 ;
        RECT 62.200 95.200 62.500 95.800 ;
        RECT 60.600 95.100 61.000 95.200 ;
        RECT 61.400 95.100 61.800 95.200 ;
        RECT 60.600 94.800 61.800 95.100 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 63.800 91.800 64.200 92.200 ;
        RECT 60.600 88.800 61.000 89.200 ;
        RECT 53.400 86.800 53.800 87.200 ;
        RECT 53.400 80.200 53.700 86.800 ;
        RECT 54.200 85.100 54.600 87.900 ;
        RECT 55.000 87.800 55.400 88.200 ;
        RECT 55.800 87.800 56.200 88.200 ;
        RECT 58.200 87.800 58.600 88.200 ;
        RECT 55.000 87.200 55.300 87.800 ;
        RECT 55.000 86.800 55.400 87.200 ;
        RECT 53.400 79.800 53.800 80.200 ;
        RECT 45.400 76.800 45.800 77.200 ;
        RECT 49.400 76.800 49.800 77.200 ;
        RECT 45.400 75.200 45.700 76.800 ;
        RECT 49.400 75.200 49.700 76.800 ;
        RECT 44.600 74.800 45.000 75.200 ;
        RECT 45.400 74.800 45.800 75.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 52.600 74.800 53.000 75.200 ;
        RECT 53.400 75.100 53.800 75.200 ;
        RECT 54.200 75.100 54.600 75.200 ;
        RECT 53.400 74.800 54.600 75.100 ;
        RECT 55.000 75.100 55.300 86.800 ;
        RECT 55.800 86.200 56.100 87.800 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 55.800 85.800 56.200 86.200 ;
        RECT 57.400 85.200 57.700 86.800 ;
        RECT 58.200 85.200 58.500 87.800 ;
        RECT 60.600 87.200 60.900 88.800 ;
        RECT 60.600 86.800 61.000 87.200 ;
        RECT 63.800 86.200 64.100 91.800 ;
        RECT 64.600 89.200 64.900 94.800 ;
        RECT 65.400 94.200 65.700 95.800 ;
        RECT 68.600 94.200 68.900 95.800 ;
        RECT 69.400 95.200 69.700 106.800 ;
        RECT 70.200 105.800 70.600 106.200 ;
        RECT 70.200 105.200 70.500 105.800 ;
        RECT 70.200 104.800 70.600 105.200 ;
        RECT 70.200 96.800 70.600 97.200 ;
        RECT 70.200 95.200 70.500 96.800 ;
        RECT 71.000 95.200 71.300 113.800 ;
        RECT 71.800 110.200 72.100 135.800 ;
        RECT 75.000 135.200 75.300 141.800 ;
        RECT 75.800 139.800 76.200 140.200 ;
        RECT 78.200 139.800 78.600 140.200 ;
        RECT 75.800 135.200 76.100 139.800 ;
        RECT 78.200 135.200 78.500 139.800 ;
        RECT 75.000 134.800 75.400 135.200 ;
        RECT 75.800 134.800 76.200 135.200 ;
        RECT 78.200 134.800 78.600 135.200 ;
        RECT 79.000 134.800 79.400 135.200 ;
        RECT 74.200 132.800 74.600 133.200 ;
        RECT 75.000 133.100 75.300 134.800 ;
        RECT 75.800 134.200 76.100 134.800 ;
        RECT 79.000 134.200 79.300 134.800 ;
        RECT 80.600 134.200 80.900 151.800 ;
        RECT 82.200 143.100 82.600 148.900 ;
        RECT 86.200 146.800 86.600 147.200 ;
        RECT 86.200 146.200 86.500 146.800 ;
        RECT 84.600 146.100 85.000 146.200 ;
        RECT 85.400 146.100 85.800 146.200 ;
        RECT 84.600 145.800 85.800 146.100 ;
        RECT 86.200 145.800 86.600 146.200 ;
        RECT 83.800 144.800 84.200 145.200 ;
        RECT 83.800 139.200 84.100 144.800 ;
        RECT 87.000 143.100 87.400 148.900 ;
        RECT 83.800 138.800 84.200 139.200 ;
        RECT 85.400 138.800 85.800 139.200 ;
        RECT 85.400 136.200 85.700 138.800 ;
        RECT 87.800 136.200 88.100 160.800 ;
        RECT 88.600 152.100 89.000 157.900 ;
        RECT 103.000 156.800 103.400 157.200 ;
        RECT 89.400 153.800 89.800 154.200 ;
        RECT 89.400 148.200 89.700 153.800 ;
        RECT 90.200 153.100 90.600 155.900 ;
        RECT 91.000 154.800 91.400 155.200 ;
        RECT 93.400 154.800 93.800 155.200 ;
        RECT 96.600 154.800 97.000 155.200 ;
        RECT 99.800 155.100 100.200 155.200 ;
        RECT 100.600 155.100 101.000 155.200 ;
        RECT 99.800 154.800 101.000 155.100 ;
        RECT 91.000 149.200 91.300 154.800 ;
        RECT 91.000 148.800 91.400 149.200 ;
        RECT 88.600 145.100 89.000 147.900 ;
        RECT 89.400 147.800 89.800 148.200 ;
        RECT 89.400 147.200 89.700 147.800 ;
        RECT 89.400 146.800 89.800 147.200 ;
        RECT 81.400 135.800 81.800 136.200 ;
        RECT 85.400 135.800 85.800 136.200 ;
        RECT 86.200 135.800 86.600 136.200 ;
        RECT 87.800 136.100 88.200 136.200 ;
        RECT 88.600 136.100 89.000 136.200 ;
        RECT 87.800 135.800 89.000 136.100 ;
        RECT 81.400 135.200 81.700 135.800 ;
        RECT 81.400 134.800 81.800 135.200 ;
        RECT 83.800 135.100 84.200 135.200 ;
        RECT 84.600 135.100 85.000 135.200 ;
        RECT 83.800 134.800 85.000 135.100 ;
        RECT 85.400 134.200 85.700 135.800 ;
        RECT 86.200 135.200 86.500 135.800 ;
        RECT 86.200 134.800 86.600 135.200 ;
        RECT 88.600 134.800 89.000 135.200 ;
        RECT 88.600 134.200 88.900 134.800 ;
        RECT 75.800 133.800 76.200 134.200 ;
        RECT 79.000 133.800 79.400 134.200 ;
        RECT 80.600 133.800 81.000 134.200 ;
        RECT 84.600 133.800 85.000 134.200 ;
        RECT 85.400 133.800 85.800 134.200 ;
        RECT 88.600 133.800 89.000 134.200 ;
        RECT 84.600 133.200 84.900 133.800 ;
        RECT 75.000 132.800 76.100 133.100 ;
        RECT 84.600 132.800 85.000 133.200 ;
        RECT 88.600 132.800 89.000 133.200 ;
        RECT 74.200 129.200 74.500 132.800 ;
        RECT 74.200 128.800 74.600 129.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 74.200 118.200 74.500 121.800 ;
        RECT 74.200 117.800 74.600 118.200 ;
        RECT 74.200 116.100 74.600 116.200 ;
        RECT 75.000 116.100 75.400 116.200 ;
        RECT 74.200 115.800 75.400 116.100 ;
        RECT 74.200 114.200 74.500 115.800 ;
        RECT 75.000 114.800 75.400 115.200 ;
        RECT 72.600 113.800 73.000 114.200 ;
        RECT 74.200 113.800 74.600 114.200 ;
        RECT 72.600 112.200 72.900 113.800 ;
        RECT 72.600 111.800 73.000 112.200 ;
        RECT 74.200 111.800 74.600 112.200 ;
        RECT 71.800 109.800 72.200 110.200 ;
        RECT 72.600 106.800 73.000 107.200 ;
        RECT 72.600 106.200 72.900 106.800 ;
        RECT 72.600 105.800 73.000 106.200 ;
        RECT 72.600 105.100 73.000 105.200 ;
        RECT 73.400 105.100 73.800 105.200 ;
        RECT 72.600 104.800 73.800 105.100 ;
        RECT 74.200 96.200 74.500 111.800 ;
        RECT 75.000 109.200 75.300 114.800 ;
        RECT 75.000 108.800 75.400 109.200 ;
        RECT 75.800 102.200 76.100 132.800 ;
        RECT 76.600 131.800 77.000 132.200 ;
        RECT 76.600 126.200 76.900 131.800 ;
        RECT 79.800 130.800 80.200 131.200 ;
        RECT 78.200 127.800 78.600 128.200 ;
        RECT 78.200 127.200 78.500 127.800 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 79.800 126.200 80.100 130.800 ;
        RECT 88.600 129.200 88.900 132.800 ;
        RECT 89.400 129.200 89.700 146.800 ;
        RECT 93.400 142.200 93.700 154.800 ;
        RECT 96.600 154.200 96.900 154.800 ;
        RECT 94.200 153.800 94.600 154.200 ;
        RECT 96.600 153.800 97.000 154.200 ;
        RECT 101.400 154.100 101.800 154.200 ;
        RECT 102.200 154.100 102.600 154.200 ;
        RECT 101.400 153.800 102.600 154.100 ;
        RECT 93.400 141.800 93.800 142.200 ;
        RECT 93.400 139.200 93.700 141.800 ;
        RECT 94.200 141.200 94.500 153.800 ;
        RECT 99.800 152.800 100.200 153.200 ;
        RECT 99.800 152.200 100.100 152.800 ;
        RECT 95.000 151.800 95.400 152.200 ;
        RECT 99.800 151.800 100.200 152.200 ;
        RECT 102.200 151.800 102.600 152.200 ;
        RECT 95.000 147.200 95.300 151.800 ;
        RECT 95.000 146.800 95.400 147.200 ;
        RECT 95.800 145.800 96.200 146.200 ;
        RECT 95.000 143.800 95.400 144.200 ;
        RECT 94.200 140.800 94.600 141.200 ;
        RECT 93.400 138.800 93.800 139.200 ;
        RECT 90.200 133.800 90.600 134.200 ;
        RECT 90.200 132.200 90.500 133.800 ;
        RECT 91.000 133.100 91.400 135.900 ;
        RECT 90.200 131.800 90.600 132.200 ;
        RECT 92.600 132.100 93.000 137.900 ;
        RECT 93.400 135.800 93.800 136.200 ;
        RECT 93.400 135.100 93.700 135.800 ;
        RECT 93.400 134.700 93.800 135.100 ;
        RECT 87.000 128.800 87.400 129.200 ;
        RECT 88.600 128.800 89.000 129.200 ;
        RECT 89.400 128.800 89.800 129.200 ;
        RECT 91.000 128.800 91.400 129.200 ;
        RECT 93.400 128.800 93.800 129.200 ;
        RECT 84.600 127.800 85.000 128.200 ;
        RECT 86.200 127.800 86.600 128.200 ;
        RECT 84.600 127.200 84.900 127.800 ;
        RECT 86.200 127.200 86.500 127.800 ;
        RECT 81.400 126.800 81.800 127.200 ;
        RECT 82.200 127.100 82.600 127.200 ;
        RECT 83.000 127.100 83.400 127.200 ;
        RECT 82.200 126.800 83.400 127.100 ;
        RECT 84.600 126.800 85.000 127.200 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 76.600 125.800 77.000 126.200 ;
        RECT 77.400 125.800 77.800 126.200 ;
        RECT 78.200 126.100 78.600 126.200 ;
        RECT 79.000 126.100 79.400 126.200 ;
        RECT 78.200 125.800 79.400 126.100 ;
        RECT 79.800 125.800 80.200 126.200 ;
        RECT 80.600 125.800 81.000 126.200 ;
        RECT 77.400 119.200 77.700 125.800 ;
        RECT 80.600 120.200 80.900 125.800 ;
        RECT 81.400 125.200 81.700 126.800 ;
        RECT 87.000 126.200 87.300 128.800 ;
        RECT 89.400 126.800 89.800 127.200 ;
        RECT 83.000 126.100 83.400 126.200 ;
        RECT 83.800 126.100 84.200 126.200 ;
        RECT 83.000 125.800 84.200 126.100 ;
        RECT 87.000 125.800 87.400 126.200 ;
        RECT 81.400 124.800 81.800 125.200 ;
        RECT 83.000 125.100 83.400 125.200 ;
        RECT 84.600 125.100 85.000 125.200 ;
        RECT 83.000 124.800 85.000 125.100 ;
        RECT 89.400 123.200 89.700 126.800 ;
        RECT 90.200 125.800 90.600 126.200 ;
        RECT 89.400 122.800 89.800 123.200 ;
        RECT 88.600 121.800 89.000 122.200 ;
        RECT 80.600 119.800 81.000 120.200 ;
        RECT 77.400 118.800 77.800 119.200 ;
        RECT 79.000 118.800 79.400 119.200 ;
        RECT 79.000 115.200 79.300 118.800 ;
        RECT 81.400 117.800 81.800 118.200 ;
        RECT 79.800 116.800 80.200 117.200 ;
        RECT 78.200 114.800 78.600 115.200 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 78.200 114.200 78.500 114.800 ;
        RECT 79.800 114.200 80.100 116.800 ;
        RECT 80.600 114.800 81.000 115.200 ;
        RECT 78.200 113.800 78.600 114.200 ;
        RECT 79.800 113.800 80.200 114.200 ;
        RECT 77.400 103.100 77.800 108.900 ;
        RECT 79.000 106.100 79.400 106.200 ;
        RECT 79.800 106.100 80.200 106.200 ;
        RECT 79.000 105.800 80.200 106.100 ;
        RECT 75.800 101.800 76.200 102.200 ;
        RECT 74.200 95.800 74.600 96.200 ;
        RECT 69.400 94.800 69.800 95.200 ;
        RECT 70.200 94.800 70.600 95.200 ;
        RECT 71.000 94.800 71.400 95.200 ;
        RECT 71.800 94.800 72.200 95.200 ;
        RECT 73.400 95.100 73.800 95.200 ;
        RECT 74.200 95.100 74.600 95.200 ;
        RECT 73.400 94.800 74.600 95.100 ;
        RECT 71.800 94.200 72.100 94.800 ;
        RECT 65.400 93.800 65.800 94.200 ;
        RECT 68.600 93.800 69.000 94.200 ;
        RECT 71.000 93.800 71.400 94.200 ;
        RECT 71.800 93.800 72.200 94.200 ;
        RECT 64.600 89.100 65.000 89.200 ;
        RECT 65.400 89.100 65.800 89.200 ;
        RECT 64.600 88.800 65.800 89.100 ;
        RECT 60.600 86.100 61.000 86.200 ;
        RECT 61.400 86.100 61.800 86.200 ;
        RECT 60.600 85.800 61.800 86.100 ;
        RECT 63.800 85.800 64.200 86.200 ;
        RECT 64.600 86.100 65.000 86.200 ;
        RECT 65.400 86.100 65.800 86.200 ;
        RECT 64.600 85.800 65.800 86.100 ;
        RECT 57.400 84.800 57.800 85.200 ;
        RECT 58.200 84.800 58.600 85.200 ;
        RECT 67.000 83.800 67.400 84.200 ;
        RECT 63.000 81.800 63.400 82.200 ;
        RECT 58.200 79.800 58.600 80.200 ;
        RECT 58.200 77.200 58.500 79.800 ;
        RECT 63.000 78.200 63.300 81.800 ;
        RECT 55.800 77.100 56.200 77.200 ;
        RECT 56.600 77.100 57.000 77.200 ;
        RECT 55.800 76.800 57.000 77.100 ;
        RECT 58.200 76.800 58.600 77.200 ;
        RECT 55.800 75.100 56.200 75.200 ;
        RECT 55.000 74.800 56.200 75.100 ;
        RECT 44.600 74.200 44.900 74.800 ;
        RECT 44.600 73.800 45.000 74.200 ;
        RECT 47.800 73.800 48.200 74.200 ;
        RECT 44.600 71.800 45.000 72.200 ;
        RECT 34.200 69.800 34.600 70.200 ;
        RECT 31.800 67.800 32.200 68.200 ;
        RECT 32.600 67.100 33.000 67.200 ;
        RECT 33.400 67.100 33.800 67.200 ;
        RECT 32.600 66.800 33.800 67.100 ;
        RECT 34.200 66.200 34.500 69.800 ;
        RECT 35.800 67.800 36.200 68.200 ;
        RECT 39.800 67.800 40.200 68.200 ;
        RECT 35.000 66.800 35.400 67.200 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 35.800 66.200 36.100 67.800 ;
        RECT 39.800 67.200 40.100 67.800 ;
        RECT 39.800 66.800 40.200 67.200 ;
        RECT 44.600 66.200 44.900 71.800 ;
        RECT 45.400 66.800 45.800 67.200 ;
        RECT 46.200 66.800 46.600 67.200 ;
        RECT 45.400 66.200 45.700 66.800 ;
        RECT 46.200 66.200 46.500 66.800 ;
        RECT 47.800 66.200 48.100 73.800 ;
        RECT 49.400 73.200 49.700 74.800 ;
        RECT 52.600 74.200 52.900 74.800 ;
        RECT 52.600 73.800 53.000 74.200 ;
        RECT 54.200 74.100 54.600 74.200 ;
        RECT 55.000 74.100 55.400 74.200 ;
        RECT 54.200 73.800 55.400 74.100 ;
        RECT 49.400 72.800 49.800 73.200 ;
        RECT 51.800 67.800 52.200 68.200 ;
        RECT 51.800 67.200 52.100 67.800 ;
        RECT 51.000 66.800 51.400 67.200 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 51.000 66.200 51.300 66.800 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 30.200 66.100 30.600 66.200 ;
        RECT 29.400 65.800 30.600 66.100 ;
        RECT 31.000 65.800 31.400 66.200 ;
        RECT 34.200 65.800 34.600 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 35.800 65.800 36.200 66.200 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 37.400 65.800 38.600 66.100 ;
        RECT 39.800 66.100 40.200 66.200 ;
        RECT 40.600 66.100 41.000 66.200 ;
        RECT 39.800 65.800 41.000 66.100 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 45.400 65.800 45.800 66.200 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 47.000 65.800 47.400 66.200 ;
        RECT 47.800 65.800 48.200 66.200 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 31.000 65.200 31.300 65.800 ;
        RECT 41.400 65.200 41.700 65.800 ;
        RECT 29.400 64.800 29.800 65.200 ;
        RECT 31.000 64.800 31.400 65.200 ;
        RECT 41.400 64.800 41.800 65.200 ;
        RECT 29.400 64.200 29.700 64.800 ;
        RECT 29.400 64.100 29.800 64.200 ;
        RECT 28.600 63.800 29.800 64.100 ;
        RECT 34.200 62.800 34.600 63.200 ;
        RECT 27.000 58.800 27.400 59.200 ;
        RECT 29.400 58.800 29.800 59.200 ;
        RECT 27.000 56.200 27.300 58.800 ;
        RECT 27.000 55.800 27.400 56.200 ;
        RECT 27.000 39.200 27.300 55.800 ;
        RECT 29.400 55.200 29.700 58.800 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 27.800 54.100 28.200 54.200 ;
        RECT 28.600 54.100 29.000 54.200 ;
        RECT 27.800 53.800 29.000 54.100 ;
        RECT 30.200 53.800 30.600 54.200 ;
        RECT 32.600 53.800 33.000 54.200 ;
        RECT 27.800 52.800 28.200 53.200 ;
        RECT 27.800 49.200 28.100 52.800 ;
        RECT 28.600 49.800 29.000 50.200 ;
        RECT 27.800 48.800 28.200 49.200 ;
        RECT 28.600 46.200 28.900 49.800 ;
        RECT 30.200 48.200 30.500 53.800 ;
        RECT 31.000 51.800 31.400 52.200 ;
        RECT 31.000 50.200 31.300 51.800 ;
        RECT 31.000 49.800 31.400 50.200 ;
        RECT 30.200 47.800 30.600 48.200 ;
        RECT 29.400 46.800 29.800 47.200 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 31.000 47.100 31.300 49.800 ;
        RECT 32.600 49.200 32.900 53.800 ;
        RECT 33.400 52.100 33.800 57.900 ;
        RECT 32.600 48.800 33.000 49.200 ;
        RECT 30.200 46.800 31.300 47.100 ;
        RECT 29.400 46.200 29.700 46.800 ;
        RECT 34.200 46.200 34.500 62.800 ;
        RECT 43.000 59.200 43.300 65.800 ;
        RECT 44.600 65.100 44.900 65.800 ;
        RECT 44.600 64.800 45.700 65.100 ;
        RECT 43.000 58.800 43.400 59.200 ;
        RECT 36.600 54.800 37.000 55.200 ;
        RECT 36.600 54.200 36.900 54.800 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 38.200 52.100 38.600 57.900 ;
        RECT 45.400 56.200 45.700 64.800 ;
        RECT 47.000 59.200 47.300 65.800 ;
        RECT 50.200 61.200 50.500 65.800 ;
        RECT 51.800 64.800 52.200 65.200 ;
        RECT 51.800 64.200 52.100 64.800 ;
        RECT 51.800 63.800 52.200 64.200 ;
        RECT 52.600 62.200 52.900 73.800 ;
        RECT 59.000 72.100 59.400 77.900 ;
        RECT 63.000 77.800 63.400 78.200 ;
        RECT 61.400 75.100 61.800 75.200 ;
        RECT 62.200 75.100 62.600 75.200 ;
        RECT 61.400 74.800 62.600 75.100 ;
        RECT 63.000 73.800 63.400 74.200 ;
        RECT 53.400 70.800 53.800 71.200 ;
        RECT 53.400 67.200 53.700 70.800 ;
        RECT 55.800 67.800 56.200 68.200 ;
        RECT 55.800 67.200 56.100 67.800 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 55.800 66.800 56.200 67.200 ;
        RECT 57.400 67.100 57.800 67.200 ;
        RECT 58.200 67.100 58.600 67.200 ;
        RECT 57.400 66.800 58.600 67.100 ;
        RECT 59.000 66.800 59.400 67.200 ;
        RECT 63.000 67.100 63.300 73.800 ;
        RECT 63.800 72.100 64.200 77.900 ;
        RECT 64.600 74.800 65.000 75.200 ;
        RECT 64.600 74.200 64.900 74.800 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 65.400 73.100 65.800 75.900 ;
        RECT 67.000 75.200 67.300 83.800 ;
        RECT 67.800 83.100 68.200 88.900 ;
        RECT 71.000 87.200 71.300 93.800 ;
        RECT 75.000 93.100 75.400 95.900 ;
        RECT 75.800 93.800 76.200 94.200 ;
        RECT 75.800 93.200 76.100 93.800 ;
        RECT 75.800 92.800 76.200 93.200 ;
        RECT 76.600 92.100 77.000 97.900 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 77.400 94.800 78.600 95.100 ;
        RECT 77.400 94.700 77.800 94.800 ;
        RECT 80.600 92.200 80.900 114.800 ;
        RECT 81.400 108.200 81.700 117.800 ;
        RECT 83.000 115.800 83.400 116.200 ;
        RECT 83.000 115.200 83.300 115.800 ;
        RECT 83.000 114.800 83.400 115.200 ;
        RECT 84.600 113.800 85.000 114.200 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 82.200 110.200 82.500 111.800 ;
        RECT 82.200 109.800 82.600 110.200 ;
        RECT 84.600 109.200 84.900 113.800 ;
        RECT 85.400 113.100 85.800 115.900 ;
        RECT 87.000 112.100 87.400 117.900 ;
        RECT 88.600 117.200 88.900 121.800 ;
        RECT 90.200 120.200 90.500 125.800 ;
        RECT 90.200 119.800 90.600 120.200 ;
        RECT 88.600 116.800 89.000 117.200 ;
        RECT 88.600 114.800 89.000 115.200 ;
        RECT 88.600 113.200 88.900 114.800 ;
        RECT 87.800 112.800 88.200 113.200 ;
        RECT 88.600 112.800 89.000 113.200 ;
        RECT 87.000 109.800 87.400 110.200 ;
        RECT 81.400 107.800 81.800 108.200 ;
        RECT 82.200 103.100 82.600 108.900 ;
        RECT 83.000 108.800 83.400 109.200 ;
        RECT 84.600 108.800 85.000 109.200 ;
        RECT 80.600 91.800 81.000 92.200 ;
        RECT 81.400 92.100 81.800 97.900 ;
        RECT 83.000 89.200 83.300 108.800 ;
        RECT 83.800 105.100 84.200 107.900 ;
        RECT 84.600 105.100 85.000 107.900 ;
        RECT 86.200 103.100 86.600 108.900 ;
        RECT 87.000 106.300 87.300 109.800 ;
        RECT 87.000 105.900 87.400 106.300 ;
        RECT 83.800 99.800 84.200 100.200 ;
        RECT 83.800 99.200 84.100 99.800 ;
        RECT 83.800 98.800 84.200 99.200 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 84.600 93.100 85.000 95.900 ;
        RECT 84.600 91.800 85.000 92.200 ;
        RECT 86.200 92.100 86.600 97.900 ;
        RECT 84.600 89.200 84.900 91.800 ;
        RECT 71.000 86.800 71.400 87.200 ;
        RECT 70.200 85.800 70.600 86.200 ;
        RECT 70.200 85.200 70.500 85.800 ;
        RECT 70.200 84.800 70.600 85.200 ;
        RECT 70.200 83.800 70.600 84.200 ;
        RECT 67.000 74.800 67.400 75.200 ;
        RECT 68.600 74.800 69.000 75.200 ;
        RECT 68.600 72.200 68.900 74.800 ;
        RECT 67.000 71.800 67.400 72.200 ;
        RECT 68.600 71.800 69.000 72.200 ;
        RECT 67.000 69.200 67.300 71.800 ;
        RECT 67.000 68.800 67.400 69.200 ;
        RECT 66.200 68.100 66.600 68.200 ;
        RECT 66.200 67.800 68.900 68.100 ;
        RECT 68.600 67.200 68.900 67.800 ;
        RECT 70.200 67.200 70.500 83.800 ;
        RECT 71.000 79.200 71.300 86.800 ;
        RECT 72.600 83.100 73.000 88.900 ;
        RECT 81.400 88.800 81.800 89.200 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 73.400 86.800 73.800 87.200 ;
        RECT 73.400 86.200 73.700 86.800 ;
        RECT 73.400 85.800 73.800 86.200 ;
        RECT 74.200 85.100 74.600 87.900 ;
        RECT 81.400 87.200 81.700 88.800 ;
        RECT 75.000 86.800 75.400 87.200 ;
        RECT 81.400 86.800 81.800 87.200 ;
        RECT 84.600 86.800 85.000 87.200 ;
        RECT 85.400 87.100 85.800 87.200 ;
        RECT 86.200 87.100 86.600 87.200 ;
        RECT 85.400 86.800 86.600 87.100 ;
        RECT 75.000 86.200 75.300 86.800 ;
        RECT 75.000 85.800 75.400 86.200 ;
        RECT 80.600 85.800 81.000 86.200 ;
        RECT 79.000 82.800 79.400 83.200 ;
        RECT 71.000 78.800 71.400 79.200 ;
        RECT 74.200 76.800 74.600 77.200 ;
        RECT 74.200 75.200 74.500 76.800 ;
        RECT 75.800 75.800 76.200 76.200 ;
        RECT 76.600 75.800 77.000 76.200 ;
        RECT 75.800 75.200 76.100 75.800 ;
        RECT 72.600 75.100 73.000 75.200 ;
        RECT 73.400 75.100 73.800 75.200 ;
        RECT 72.600 74.800 73.800 75.100 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 75.800 74.800 76.200 75.200 ;
        RECT 71.800 72.800 72.200 73.200 ;
        RECT 71.000 69.800 71.400 70.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 65.400 67.100 65.800 67.200 ;
        RECT 63.000 66.800 64.100 67.100 ;
        RECT 64.600 66.800 65.800 67.100 ;
        RECT 67.000 67.100 67.400 67.200 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 67.000 66.800 68.200 67.100 ;
        RECT 68.600 66.800 69.000 67.200 ;
        RECT 70.200 66.800 70.600 67.200 ;
        RECT 55.000 66.200 55.300 66.800 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 55.000 65.800 55.400 66.200 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 52.600 61.800 53.000 62.200 ;
        RECT 50.200 60.800 50.600 61.200 ;
        RECT 51.800 59.800 52.200 60.200 ;
        RECT 47.000 58.800 47.400 59.200 ;
        RECT 51.800 58.200 52.100 59.800 ;
        RECT 54.200 59.200 54.500 65.800 ;
        RECT 58.200 65.200 58.500 65.800 ;
        RECT 57.400 64.800 57.800 65.200 ;
        RECT 58.200 64.800 58.600 65.200 ;
        RECT 57.400 64.200 57.700 64.800 ;
        RECT 59.000 64.200 59.300 66.800 ;
        RECT 63.800 66.200 64.100 66.800 ;
        RECT 71.000 66.200 71.300 69.800 ;
        RECT 71.800 66.200 72.100 72.800 ;
        RECT 76.600 68.200 76.900 75.800 ;
        RECT 77.400 73.800 77.800 74.200 ;
        RECT 77.400 73.200 77.700 73.800 ;
        RECT 77.400 72.800 77.800 73.200 ;
        RECT 78.200 73.100 78.600 75.900 ;
        RECT 76.600 67.800 77.000 68.200 ;
        RECT 77.400 68.100 77.800 68.200 ;
        RECT 78.200 68.100 78.600 68.200 ;
        RECT 77.400 67.800 78.600 68.100 ;
        RECT 76.600 67.200 76.900 67.800 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 76.600 66.800 77.000 67.200 ;
        RECT 78.200 66.800 78.600 67.200 ;
        RECT 75.000 66.200 75.300 66.800 ;
        RECT 62.200 66.100 62.600 66.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 62.200 65.800 63.400 66.100 ;
        RECT 63.800 65.800 64.200 66.200 ;
        RECT 67.800 66.100 68.200 66.200 ;
        RECT 67.000 65.800 68.200 66.100 ;
        RECT 68.600 65.800 69.000 66.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 71.800 65.800 72.200 66.200 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 73.400 65.800 74.600 66.100 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 75.800 65.800 77.000 66.100 ;
        RECT 60.600 64.800 61.000 65.200 ;
        RECT 63.800 64.800 64.200 65.200 ;
        RECT 60.600 64.200 60.900 64.800 ;
        RECT 63.800 64.200 64.100 64.800 ;
        RECT 57.400 63.800 57.800 64.200 ;
        RECT 59.000 63.800 59.400 64.200 ;
        RECT 60.600 63.800 61.000 64.200 ;
        RECT 63.800 63.800 64.200 64.200 ;
        RECT 62.200 61.800 62.600 62.200 ;
        RECT 54.200 58.800 54.600 59.200 ;
        RECT 51.800 57.800 52.200 58.200 ;
        RECT 39.000 53.800 39.400 54.200 ;
        RECT 37.400 49.800 37.800 50.200 ;
        RECT 35.000 47.100 35.400 47.200 ;
        RECT 35.800 47.100 36.200 47.200 ;
        RECT 35.000 46.800 36.200 47.100 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 29.400 46.100 29.800 46.200 ;
        RECT 29.400 45.800 30.500 46.100 ;
        RECT 27.000 38.800 27.400 39.200 ;
        RECT 27.000 32.100 27.400 37.900 ;
        RECT 29.400 36.800 29.800 37.200 ;
        RECT 29.400 35.200 29.700 36.800 ;
        RECT 30.200 35.200 30.500 45.800 ;
        RECT 31.800 45.800 32.200 46.200 ;
        RECT 34.200 45.800 34.600 46.200 ;
        RECT 31.800 45.200 32.100 45.800 ;
        RECT 31.800 44.800 32.200 45.200 ;
        RECT 32.600 44.800 33.000 45.200 ;
        RECT 32.600 39.200 32.900 44.800 ;
        RECT 32.600 38.800 33.000 39.200 ;
        RECT 35.000 37.200 35.300 46.800 ;
        RECT 35.800 44.100 36.200 44.200 ;
        RECT 36.600 44.100 37.000 44.200 ;
        RECT 35.800 43.800 37.000 44.100 ;
        RECT 37.400 39.200 37.700 49.800 ;
        RECT 38.200 43.100 38.600 48.900 ;
        RECT 39.000 46.200 39.300 53.800 ;
        RECT 39.800 53.100 40.200 55.900 ;
        RECT 44.600 55.800 45.000 56.200 ;
        RECT 45.400 55.800 45.800 56.200 ;
        RECT 44.600 55.200 44.900 55.800 ;
        RECT 45.400 55.200 45.700 55.800 ;
        RECT 51.800 55.200 52.100 57.800 ;
        RECT 55.000 56.800 55.400 57.200 ;
        RECT 55.000 55.200 55.300 56.800 ;
        RECT 62.200 56.200 62.500 61.800 ;
        RECT 66.200 60.800 66.600 61.200 ;
        RECT 66.200 56.200 66.500 60.800 ;
        RECT 57.400 55.800 57.800 56.200 ;
        RECT 62.200 55.800 62.600 56.200 ;
        RECT 63.800 55.800 64.200 56.200 ;
        RECT 66.200 55.800 66.600 56.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 41.400 55.100 41.800 55.200 ;
        RECT 40.600 54.800 41.800 55.100 ;
        RECT 43.800 54.800 44.200 55.200 ;
        RECT 44.600 54.800 45.000 55.200 ;
        RECT 45.400 54.800 45.800 55.200 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 46.200 54.800 47.400 55.100 ;
        RECT 48.600 54.800 49.000 55.200 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 51.800 54.800 52.200 55.200 ;
        RECT 52.600 54.800 53.000 55.200 ;
        RECT 55.000 54.800 55.400 55.200 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 42.200 51.800 42.600 52.200 ;
        RECT 42.200 46.300 42.500 51.800 ;
        RECT 43.800 49.200 44.100 54.800 ;
        RECT 46.200 53.800 46.600 54.200 ;
        RECT 46.200 49.200 46.500 53.800 ;
        RECT 48.600 50.200 48.900 54.800 ;
        RECT 48.600 49.800 49.000 50.200 ;
        RECT 51.000 49.200 51.300 54.800 ;
        RECT 39.000 45.800 39.400 46.200 ;
        RECT 42.200 45.900 42.600 46.300 ;
        RECT 37.400 38.800 37.800 39.200 ;
        RECT 39.000 37.200 39.300 45.800 ;
        RECT 43.000 43.100 43.400 48.900 ;
        RECT 43.800 48.800 44.200 49.200 ;
        RECT 45.400 48.800 45.800 49.200 ;
        RECT 46.200 48.800 46.600 49.200 ;
        RECT 51.000 48.800 51.400 49.200 ;
        RECT 44.600 45.100 45.000 47.900 ;
        RECT 45.400 47.200 45.700 48.800 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 46.200 46.800 46.600 47.200 ;
        RECT 45.400 44.800 45.800 45.200 ;
        RECT 45.400 44.200 45.700 44.800 ;
        RECT 45.400 43.800 45.800 44.200 ;
        RECT 46.200 39.200 46.500 46.800 ;
        RECT 51.000 43.800 51.400 44.200 ;
        RECT 46.200 38.800 46.600 39.200 ;
        RECT 35.000 36.800 35.400 37.200 ;
        RECT 37.400 36.800 37.800 37.200 ;
        RECT 39.000 36.800 39.400 37.200 ;
        RECT 29.400 34.800 29.800 35.200 ;
        RECT 30.200 34.800 30.600 35.200 ;
        RECT 31.000 34.800 31.400 35.200 ;
        RECT 33.400 34.800 33.800 35.200 ;
        RECT 35.800 34.800 36.200 35.200 ;
        RECT 31.000 31.200 31.300 34.800 ;
        RECT 33.400 32.200 33.700 34.800 ;
        RECT 33.400 31.800 33.800 32.200 ;
        RECT 31.000 30.800 31.400 31.200 ;
        RECT 30.200 29.800 30.600 30.200 ;
        RECT 31.000 29.800 31.400 30.200 ;
        RECT 30.200 29.200 30.500 29.800 ;
        RECT 31.000 29.200 31.300 29.800 ;
        RECT 24.600 25.800 25.000 26.200 ;
        RECT 26.200 25.800 26.600 26.200 ;
        RECT 17.400 21.800 17.800 22.200 ;
        RECT 15.800 16.800 16.200 17.200 ;
        RECT 15.800 16.200 16.100 16.800 ;
        RECT 9.400 13.100 9.800 15.900 ;
        RECT 11.800 15.800 12.200 16.200 ;
        RECT 12.600 15.800 13.000 16.200 ;
        RECT 15.000 15.800 15.400 16.200 ;
        RECT 15.800 15.800 16.200 16.200 ;
        RECT 17.400 15.800 17.800 16.200 ;
        RECT 11.800 15.200 12.100 15.800 ;
        RECT 10.200 14.800 10.600 15.200 ;
        RECT 11.800 14.800 12.200 15.200 ;
        RECT 10.200 14.200 10.500 14.800 ;
        RECT 12.600 14.200 12.900 15.800 ;
        RECT 14.200 15.100 14.600 15.200 ;
        RECT 15.000 15.100 15.400 15.200 ;
        RECT 14.200 14.800 15.400 15.100 ;
        RECT 10.200 13.800 10.600 14.200 ;
        RECT 12.600 13.800 13.000 14.200 ;
        RECT 14.200 14.100 14.600 14.200 ;
        RECT 15.000 14.100 15.400 14.200 ;
        RECT 14.200 13.800 15.400 14.100 ;
        RECT 7.000 7.100 7.400 7.200 ;
        RECT 7.800 7.100 8.200 7.200 ;
        RECT 7.000 6.800 8.200 7.100 ;
        RECT 14.200 7.100 14.600 7.200 ;
        RECT 15.000 7.100 15.400 7.200 ;
        RECT 14.200 6.800 15.400 7.100 ;
        RECT 15.800 6.200 16.100 15.800 ;
        RECT 17.400 15.200 17.700 15.800 ;
        RECT 17.400 14.800 17.800 15.200 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 20.600 14.200 20.900 14.800 ;
        RECT 21.400 14.200 21.700 14.800 ;
        RECT 17.400 13.800 17.800 14.200 ;
        RECT 19.000 14.100 19.400 14.200 ;
        RECT 19.800 14.100 20.200 14.200 ;
        RECT 19.000 13.800 20.200 14.100 ;
        RECT 20.600 13.800 21.000 14.200 ;
        RECT 21.400 13.800 21.800 14.200 ;
        RECT 16.600 11.800 17.000 12.200 ;
        RECT 16.600 7.100 16.900 11.800 ;
        RECT 17.400 10.200 17.700 13.800 ;
        RECT 17.400 9.800 17.800 10.200 ;
        RECT 16.600 6.800 17.700 7.100 ;
        RECT 14.200 6.100 14.600 6.200 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 14.200 5.800 15.400 6.100 ;
        RECT 15.800 5.800 16.200 6.200 ;
        RECT 16.600 5.800 17.000 6.200 ;
        RECT 16.600 5.200 16.900 5.800 ;
        RECT 17.400 5.200 17.700 6.800 ;
        RECT 16.600 4.800 17.000 5.200 ;
        RECT 17.400 4.800 17.800 5.200 ;
        RECT 18.200 5.100 18.600 7.900 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 19.000 6.200 19.300 6.800 ;
        RECT 19.000 5.800 19.400 6.200 ;
        RECT 19.800 3.100 20.200 8.900 ;
        RECT 21.400 8.200 21.700 13.800 ;
        RECT 23.000 12.800 23.400 13.200 ;
        RECT 23.800 13.100 24.200 15.900 ;
        RECT 24.600 13.800 25.000 14.200 ;
        RECT 24.600 13.200 24.900 13.800 ;
        RECT 24.600 12.800 25.000 13.200 ;
        RECT 23.000 12.200 23.300 12.800 ;
        RECT 23.000 11.800 23.400 12.200 ;
        RECT 25.400 12.100 25.800 17.900 ;
        RECT 26.200 17.200 26.500 25.800 ;
        RECT 27.800 23.100 28.200 28.900 ;
        RECT 30.200 28.800 30.600 29.200 ;
        RECT 31.000 28.800 31.400 29.200 ;
        RECT 33.400 23.100 33.800 28.900 ;
        RECT 26.200 16.800 26.600 17.200 ;
        RECT 26.200 15.800 26.600 16.200 ;
        RECT 26.200 15.100 26.500 15.800 ;
        RECT 26.200 14.700 26.600 15.100 ;
        RECT 30.200 12.100 30.600 17.900 ;
        RECT 33.400 16.800 33.800 17.200 ;
        RECT 33.400 14.200 33.700 16.800 ;
        RECT 33.400 13.800 33.800 14.200 ;
        RECT 34.200 12.800 34.600 13.200 ;
        RECT 31.800 12.100 32.200 12.200 ;
        RECT 32.600 12.100 33.000 12.200 ;
        RECT 31.800 11.800 33.000 12.100 ;
        RECT 27.000 9.800 27.400 10.200 ;
        RECT 27.000 9.200 27.300 9.800 ;
        RECT 21.400 7.800 21.800 8.200 ;
        RECT 20.600 5.900 21.000 6.300 ;
        RECT 20.600 5.200 20.900 5.900 ;
        RECT 20.600 4.800 21.000 5.200 ;
        RECT 24.600 3.100 25.000 8.900 ;
        RECT 27.000 8.800 27.400 9.200 ;
        RECT 29.400 8.800 29.800 9.200 ;
        RECT 29.400 8.200 29.700 8.800 ;
        RECT 27.800 7.800 28.200 8.200 ;
        RECT 29.400 7.800 29.800 8.200 ;
        RECT 31.800 7.800 32.200 8.200 ;
        RECT 27.800 6.200 28.100 7.800 ;
        RECT 31.800 7.200 32.100 7.800 ;
        RECT 31.800 6.800 32.200 7.200 ;
        RECT 32.600 6.800 33.000 7.200 ;
        RECT 32.600 6.200 32.900 6.800 ;
        RECT 27.800 5.800 28.200 6.200 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 32.600 5.800 33.000 6.200 ;
        RECT 31.000 5.200 31.300 5.800 ;
        RECT 31.000 4.800 31.400 5.200 ;
        RECT 33.400 5.100 33.800 7.900 ;
        RECT 34.200 7.200 34.500 12.800 ;
        RECT 35.800 12.200 36.100 34.800 ;
        RECT 37.400 28.200 37.700 36.800 ;
        RECT 41.400 35.800 41.800 36.200 ;
        RECT 47.800 35.800 48.200 36.200 ;
        RECT 41.400 35.200 41.700 35.800 ;
        RECT 47.800 35.200 48.100 35.800 ;
        RECT 38.200 34.800 38.600 35.200 ;
        RECT 39.000 35.100 39.400 35.200 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 39.000 34.800 40.200 35.100 ;
        RECT 41.400 34.800 41.800 35.200 ;
        RECT 43.800 35.100 44.200 35.200 ;
        RECT 44.600 35.100 45.000 35.200 ;
        RECT 43.800 34.800 45.000 35.100 ;
        RECT 47.800 34.800 48.200 35.200 ;
        RECT 38.200 34.200 38.500 34.800 ;
        RECT 38.200 33.800 38.600 34.200 ;
        RECT 39.800 34.100 40.200 34.200 ;
        RECT 40.600 34.100 41.000 34.200 ;
        RECT 39.800 33.800 41.000 34.100 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 38.200 30.200 38.500 33.800 ;
        RECT 42.200 31.800 42.600 32.200 ;
        RECT 38.200 29.800 38.600 30.200 ;
        RECT 37.400 27.800 37.800 28.200 ;
        RECT 36.600 26.200 37.000 26.300 ;
        RECT 37.400 26.200 37.800 26.300 ;
        RECT 36.600 25.900 37.800 26.200 ;
        RECT 38.200 23.100 38.600 28.900 ;
        RECT 39.000 26.800 39.400 27.200 ;
        RECT 39.000 19.200 39.300 26.800 ;
        RECT 39.800 25.100 40.200 27.900 ;
        RECT 42.200 26.200 42.500 31.800 ;
        RECT 50.200 29.200 50.500 33.800 ;
        RECT 42.200 25.800 42.600 26.200 ;
        RECT 40.600 23.100 41.000 23.200 ;
        RECT 41.400 23.100 41.800 23.200 ;
        RECT 43.000 23.100 43.400 28.900 ;
        RECT 47.000 26.800 47.400 27.200 ;
        RECT 47.000 26.300 47.300 26.800 ;
        RECT 47.000 25.900 47.400 26.300 ;
        RECT 47.800 23.100 48.200 28.900 ;
        RECT 50.200 28.800 50.600 29.200 ;
        RECT 48.600 27.800 49.000 28.200 ;
        RECT 48.600 27.200 48.900 27.800 ;
        RECT 48.600 26.800 49.000 27.200 ;
        RECT 49.400 25.100 49.800 27.900 ;
        RECT 50.200 26.200 50.500 28.800 ;
        RECT 50.200 25.800 50.600 26.200 ;
        RECT 40.600 22.800 41.800 23.100 ;
        RECT 47.000 21.800 47.400 22.200 ;
        RECT 47.000 19.200 47.300 21.800 ;
        RECT 39.000 18.800 39.400 19.200 ;
        RECT 43.000 19.100 43.400 19.200 ;
        RECT 43.800 19.100 44.200 19.200 ;
        RECT 43.000 18.800 44.200 19.100 ;
        RECT 47.000 18.800 47.400 19.200 ;
        RECT 48.600 17.800 49.000 18.200 ;
        RECT 48.600 15.200 48.900 17.800 ;
        RECT 51.000 15.200 51.300 43.800 ;
        RECT 52.600 43.200 52.900 54.800 ;
        RECT 56.600 54.200 56.900 54.800 ;
        RECT 57.400 54.200 57.700 55.800 ;
        RECT 63.800 55.200 64.100 55.800 ;
        RECT 61.400 55.100 61.800 55.200 ;
        RECT 62.200 55.100 62.600 55.200 ;
        RECT 61.400 54.800 62.600 55.100 ;
        RECT 63.800 54.800 64.200 55.200 ;
        RECT 66.200 54.800 66.600 55.200 ;
        RECT 66.200 54.200 66.500 54.800 ;
        RECT 56.600 53.800 57.000 54.200 ;
        RECT 57.400 53.800 57.800 54.200 ;
        RECT 61.400 54.100 61.800 54.200 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 61.400 53.800 62.600 54.100 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 63.000 53.800 64.200 54.100 ;
        RECT 66.200 53.800 66.600 54.200 ;
        RECT 58.200 52.800 58.600 53.200 ;
        RECT 59.800 53.100 60.200 53.200 ;
        RECT 60.600 53.100 61.000 53.200 ;
        RECT 59.800 52.800 61.000 53.100 ;
        RECT 58.200 52.200 58.500 52.800 ;
        RECT 58.200 51.800 58.600 52.200 ;
        RECT 60.600 51.800 61.000 52.200 ;
        RECT 60.600 50.200 60.900 51.800 ;
        RECT 58.200 49.800 58.600 50.200 ;
        RECT 60.600 49.800 61.000 50.200 ;
        RECT 53.400 46.800 53.800 47.200 ;
        RECT 52.600 42.800 53.000 43.200 ;
        RECT 51.800 36.800 52.200 37.200 ;
        RECT 51.800 36.200 52.100 36.800 ;
        RECT 51.800 35.800 52.200 36.200 ;
        RECT 51.800 34.800 52.200 35.200 ;
        RECT 51.800 26.200 52.100 34.800 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 52.600 33.200 52.900 33.800 ;
        RECT 52.600 32.800 53.000 33.200 ;
        RECT 51.800 25.800 52.200 26.200 ;
        RECT 52.600 25.800 53.000 26.200 ;
        RECT 52.600 25.200 52.900 25.800 ;
        RECT 52.600 24.800 53.000 25.200 ;
        RECT 53.400 17.200 53.700 46.800 ;
        RECT 54.200 43.100 54.600 48.900 ;
        RECT 58.200 46.300 58.500 49.800 ;
        RECT 58.200 45.900 58.600 46.300 ;
        RECT 58.200 43.800 58.600 44.200 ;
        RECT 55.000 41.800 55.400 42.200 ;
        RECT 55.000 37.200 55.300 41.800 ;
        RECT 58.200 39.200 58.500 43.800 ;
        RECT 59.000 43.100 59.400 48.900 ;
        RECT 59.800 46.800 60.200 47.200 ;
        RECT 59.800 45.200 60.100 46.800 ;
        RECT 59.800 44.800 60.200 45.200 ;
        RECT 60.600 45.100 61.000 47.900 ;
        RECT 61.400 45.100 61.800 47.900 ;
        RECT 62.200 46.800 62.600 47.200 ;
        RECT 62.200 46.200 62.500 46.800 ;
        RECT 62.200 45.800 62.600 46.200 ;
        RECT 63.000 43.100 63.400 48.900 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 64.600 46.200 64.900 46.800 ;
        RECT 64.600 45.800 65.000 46.200 ;
        RECT 67.000 39.200 67.300 65.800 ;
        RECT 68.600 65.200 68.900 65.800 ;
        RECT 68.600 64.800 69.000 65.200 ;
        RECT 72.600 61.800 73.000 62.200 ;
        RECT 67.800 55.800 68.200 56.200 ;
        RECT 67.800 54.200 68.100 55.800 ;
        RECT 67.800 53.800 68.200 54.200 ;
        RECT 68.600 53.100 69.000 55.900 ;
        RECT 69.400 53.800 69.800 54.200 ;
        RECT 69.400 49.200 69.700 53.800 ;
        RECT 70.200 52.100 70.600 57.900 ;
        RECT 72.600 57.200 72.900 61.800 ;
        RECT 78.200 59.200 78.500 66.800 ;
        RECT 79.000 66.200 79.300 82.800 ;
        RECT 79.800 72.100 80.200 77.900 ;
        RECT 80.600 74.200 80.900 85.800 ;
        RECT 84.600 85.200 84.900 86.800 ;
        RECT 82.200 84.800 82.600 85.200 ;
        RECT 84.600 85.100 85.000 85.200 ;
        RECT 85.400 85.100 85.800 85.200 ;
        RECT 84.600 84.800 85.800 85.100 ;
        RECT 82.200 83.200 82.500 84.800 ;
        RECT 86.200 84.200 86.500 86.800 ;
        RECT 87.000 85.200 87.300 98.800 ;
        RECT 87.800 94.200 88.100 112.800 ;
        RECT 89.400 100.800 89.800 101.200 ;
        RECT 89.400 95.200 89.700 100.800 ;
        RECT 90.200 100.200 90.500 119.800 ;
        RECT 91.000 115.200 91.300 128.800 ;
        RECT 93.400 126.200 93.700 128.800 ;
        RECT 94.200 126.800 94.600 127.200 ;
        RECT 94.200 126.200 94.500 126.800 ;
        RECT 95.000 126.200 95.300 143.800 ;
        RECT 95.800 135.200 96.100 145.800 ;
        RECT 98.200 145.100 98.600 147.900 ;
        RECT 99.000 146.800 99.400 147.200 ;
        RECT 99.000 146.200 99.300 146.800 ;
        RECT 99.000 145.800 99.400 146.200 ;
        RECT 99.800 143.100 100.200 148.900 ;
        RECT 100.600 146.800 101.000 147.200 ;
        RECT 100.600 146.300 100.900 146.800 ;
        RECT 100.600 145.900 101.000 146.300 ;
        RECT 102.200 146.200 102.500 151.800 ;
        RECT 102.200 145.800 102.600 146.200 ;
        RECT 95.800 134.800 96.200 135.200 ;
        RECT 97.400 132.100 97.800 137.900 ;
        RECT 102.200 133.100 102.600 135.900 ;
        RECT 103.000 134.200 103.300 156.800 ;
        RECT 111.800 155.200 112.100 163.800 ;
        RECT 114.200 161.200 114.500 165.800 ;
        RECT 118.200 165.200 118.500 174.800 ;
        RECT 119.000 173.800 119.400 174.200 ;
        RECT 119.000 171.200 119.300 173.800 ;
        RECT 119.000 170.800 119.400 171.200 ;
        RECT 119.000 168.800 119.400 169.200 ;
        RECT 119.000 167.200 119.300 168.800 ;
        RECT 119.000 166.800 119.400 167.200 ;
        RECT 117.400 164.800 117.800 165.200 ;
        RECT 118.200 164.800 118.600 165.200 ;
        RECT 117.400 161.200 117.700 164.800 ;
        RECT 114.200 160.800 114.600 161.200 ;
        RECT 117.400 160.800 117.800 161.200 ;
        RECT 112.600 159.800 113.000 160.200 ;
        RECT 112.600 159.200 112.900 159.800 ;
        RECT 112.600 158.800 113.000 159.200 ;
        RECT 118.200 158.200 118.500 164.800 ;
        RECT 103.800 154.800 104.200 155.200 ;
        RECT 105.400 155.100 105.800 155.200 ;
        RECT 106.200 155.100 106.600 155.200 ;
        RECT 105.400 154.800 106.600 155.100 ;
        RECT 109.400 154.800 109.800 155.200 ;
        RECT 111.800 154.800 112.200 155.200 ;
        RECT 103.800 154.200 104.100 154.800 ;
        RECT 109.400 154.200 109.700 154.800 ;
        RECT 103.800 153.800 104.200 154.200 ;
        RECT 107.000 154.100 107.400 154.200 ;
        RECT 107.800 154.100 108.200 154.200 ;
        RECT 107.000 153.800 108.200 154.100 ;
        RECT 109.400 153.800 109.800 154.200 ;
        RECT 105.400 152.800 105.800 153.200 ;
        RECT 111.000 152.800 111.400 153.200 ;
        RECT 114.200 153.100 114.600 155.900 ;
        RECT 115.000 154.800 115.400 155.200 ;
        RECT 115.000 154.200 115.300 154.800 ;
        RECT 115.000 153.800 115.400 154.200 ;
        RECT 105.400 150.200 105.700 152.800 ;
        RECT 107.000 151.800 107.400 152.200 ;
        RECT 107.800 152.100 108.200 152.200 ;
        RECT 108.600 152.100 109.000 152.200 ;
        RECT 107.800 151.800 109.000 152.100 ;
        RECT 105.400 149.800 105.800 150.200 ;
        RECT 107.000 149.200 107.300 151.800 ;
        RECT 111.000 151.200 111.300 152.800 ;
        RECT 115.800 152.100 116.200 157.900 ;
        RECT 118.200 157.800 118.600 158.200 ;
        RECT 117.400 155.100 117.800 155.200 ;
        RECT 118.200 155.100 118.600 155.200 ;
        RECT 117.400 154.800 118.600 155.100 ;
        RECT 111.000 150.800 111.400 151.200 ;
        RECT 116.600 149.800 117.000 150.200 ;
        RECT 118.200 149.800 118.600 150.200 ;
        RECT 116.600 149.200 116.900 149.800 ;
        RECT 104.600 143.100 105.000 148.900 ;
        RECT 107.000 148.800 107.400 149.200 ;
        RECT 107.800 145.100 108.200 147.900 ;
        RECT 108.600 147.800 109.000 148.200 ;
        RECT 108.600 147.200 108.900 147.800 ;
        RECT 108.600 146.800 109.000 147.200 ;
        RECT 109.400 143.100 109.800 148.900 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 110.200 146.300 110.500 146.800 ;
        RECT 110.200 145.900 110.600 146.300 ;
        RECT 114.200 143.100 114.600 148.900 ;
        RECT 116.600 148.800 117.000 149.200 ;
        RECT 118.200 146.200 118.500 149.800 ;
        RECT 117.400 145.800 117.800 146.200 ;
        RECT 118.200 145.800 118.600 146.200 ;
        RECT 117.400 143.200 117.700 145.800 ;
        RECT 117.400 142.800 117.800 143.200 ;
        RECT 116.600 141.800 117.000 142.200 ;
        RECT 119.000 141.800 119.400 142.200 ;
        RECT 111.800 139.800 112.200 140.200 ;
        RECT 107.000 138.800 107.400 139.200 ;
        RECT 103.000 133.800 103.400 134.200 ;
        RECT 99.000 132.100 99.400 132.200 ;
        RECT 99.800 132.100 100.200 132.200 ;
        RECT 99.000 131.800 100.200 132.100 ;
        RECT 102.200 129.100 102.600 129.200 ;
        RECT 101.400 128.800 102.600 129.100 ;
        RECT 101.400 128.200 101.700 128.800 ;
        RECT 101.400 127.800 101.800 128.200 ;
        RECT 102.200 127.800 102.600 128.200 ;
        RECT 102.200 127.200 102.500 127.800 ;
        RECT 100.600 126.800 101.000 127.200 ;
        RECT 101.400 126.800 101.800 127.200 ;
        RECT 102.200 126.800 102.600 127.200 ;
        RECT 100.600 126.200 100.900 126.800 ;
        RECT 101.400 126.200 101.700 126.800 ;
        RECT 93.400 125.800 93.800 126.200 ;
        RECT 94.200 125.800 94.600 126.200 ;
        RECT 95.000 125.800 95.400 126.200 ;
        RECT 95.800 125.800 96.200 126.200 ;
        RECT 97.400 126.100 97.800 126.200 ;
        RECT 98.200 126.100 98.600 126.200 ;
        RECT 97.400 125.800 98.600 126.100 ;
        RECT 100.600 125.800 101.000 126.200 ;
        RECT 101.400 125.800 101.800 126.200 ;
        RECT 92.600 124.800 93.000 125.200 ;
        RECT 91.000 114.800 91.400 115.200 ;
        RECT 91.800 112.100 92.200 117.900 ;
        RECT 92.600 109.200 92.900 124.800 ;
        RECT 94.200 119.200 94.500 125.800 ;
        RECT 95.000 123.200 95.300 125.800 ;
        RECT 95.000 122.800 95.400 123.200 ;
        RECT 95.000 119.800 95.400 120.200 ;
        RECT 94.200 118.800 94.600 119.200 ;
        RECT 93.400 116.800 93.800 117.200 ;
        RECT 94.200 116.800 94.600 117.200 ;
        RECT 93.400 112.100 93.700 116.800 ;
        RECT 94.200 115.200 94.500 116.800 ;
        RECT 94.200 114.800 94.600 115.200 ;
        RECT 95.000 114.200 95.300 119.800 ;
        RECT 95.800 115.200 96.100 125.800 ;
        RECT 101.400 120.200 101.700 125.800 ;
        RECT 103.000 123.200 103.300 133.800 ;
        RECT 103.800 132.100 104.200 137.900 ;
        RECT 104.600 134.800 105.000 135.200 ;
        RECT 105.400 135.100 105.800 135.200 ;
        RECT 106.200 135.100 106.600 135.200 ;
        RECT 105.400 134.800 106.600 135.100 ;
        RECT 104.600 134.200 104.900 134.800 ;
        RECT 104.600 133.800 105.000 134.200 ;
        RECT 103.800 126.800 104.200 127.200 ;
        RECT 103.000 122.800 103.400 123.200 ;
        RECT 101.400 119.800 101.800 120.200 ;
        RECT 97.400 115.800 97.800 116.200 ;
        RECT 99.000 115.800 99.400 116.200 ;
        RECT 95.800 114.800 96.200 115.200 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 96.600 114.200 96.900 114.800 ;
        RECT 95.000 113.800 95.400 114.200 ;
        RECT 96.600 113.800 97.000 114.200 ;
        RECT 93.400 111.800 94.500 112.100 ;
        RECT 92.600 109.100 93.000 109.200 ;
        RECT 93.400 109.100 93.800 109.200 ;
        RECT 91.000 103.100 91.400 108.900 ;
        RECT 92.600 108.800 93.800 109.100 ;
        RECT 94.200 107.200 94.500 111.800 ;
        RECT 96.600 111.800 97.000 112.200 ;
        RECT 94.200 106.800 94.600 107.200 ;
        RECT 95.000 106.800 95.400 107.200 ;
        RECT 95.000 106.200 95.300 106.800 ;
        RECT 91.800 105.800 92.200 106.200 ;
        RECT 95.000 105.800 95.400 106.200 ;
        RECT 90.200 99.800 90.600 100.200 ;
        RECT 90.200 95.800 90.600 96.200 ;
        RECT 89.400 94.800 89.800 95.200 ;
        RECT 87.800 93.800 88.200 94.200 ;
        RECT 87.800 93.200 88.100 93.800 ;
        RECT 87.800 92.800 88.200 93.200 ;
        RECT 87.800 89.200 88.100 92.800 ;
        RECT 90.200 89.200 90.500 95.800 ;
        RECT 91.000 92.100 91.400 97.900 ;
        RECT 87.800 88.800 88.200 89.200 ;
        RECT 90.200 88.800 90.600 89.200 ;
        RECT 90.200 88.200 90.500 88.800 ;
        RECT 90.200 87.800 90.600 88.200 ;
        RECT 89.400 86.800 89.800 87.200 ;
        RECT 88.600 85.800 89.000 86.200 ;
        RECT 88.600 85.200 88.900 85.800 ;
        RECT 89.400 85.200 89.700 86.800 ;
        RECT 91.800 86.200 92.100 105.800 ;
        RECT 96.600 105.200 96.900 111.800 ;
        RECT 97.400 107.200 97.700 115.800 ;
        RECT 99.000 115.200 99.300 115.800 ;
        RECT 103.000 115.200 103.300 122.800 ;
        RECT 103.800 122.200 104.100 126.800 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 105.400 126.100 105.800 126.200 ;
        RECT 104.600 125.800 105.800 126.100 ;
        RECT 103.800 121.800 104.200 122.200 ;
        RECT 105.400 121.800 105.800 122.200 ;
        RECT 99.000 114.800 99.400 115.200 ;
        RECT 102.200 115.100 102.600 115.200 ;
        RECT 103.000 115.100 103.400 115.200 ;
        RECT 102.200 114.800 103.400 115.100 ;
        RECT 99.800 113.100 100.200 113.200 ;
        RECT 100.600 113.100 101.000 113.200 ;
        RECT 99.800 112.800 101.000 113.100 ;
        RECT 103.800 112.200 104.100 121.800 ;
        RECT 104.600 116.800 105.000 117.200 ;
        RECT 104.600 115.200 104.900 116.800 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 104.600 114.100 105.000 114.200 ;
        RECT 105.400 114.100 105.700 121.800 ;
        RECT 107.000 116.200 107.300 138.800 ;
        RECT 108.600 132.100 109.000 137.900 ;
        RECT 111.800 137.200 112.100 139.800 ;
        RECT 109.400 136.800 109.800 137.200 ;
        RECT 111.800 136.800 112.200 137.200 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 108.600 126.200 108.900 126.800 ;
        RECT 109.400 126.200 109.700 136.800 ;
        RECT 111.800 134.200 112.100 136.800 ;
        RECT 113.400 136.100 113.800 136.200 ;
        RECT 114.200 136.100 114.600 136.200 ;
        RECT 113.400 135.800 114.600 136.100 ;
        RECT 115.800 135.800 116.200 136.200 ;
        RECT 115.800 135.200 116.100 135.800 ;
        RECT 113.400 134.800 113.800 135.200 ;
        RECT 115.800 134.800 116.200 135.200 ;
        RECT 113.400 134.200 113.700 134.800 ;
        RECT 111.800 133.800 112.200 134.200 ;
        RECT 113.400 133.800 113.800 134.200 ;
        RECT 113.400 131.800 113.800 132.200 ;
        RECT 110.200 126.800 110.600 127.200 ;
        RECT 110.200 126.200 110.500 126.800 ;
        RECT 113.400 126.200 113.700 131.800 ;
        RECT 115.800 130.200 116.100 134.800 ;
        RECT 116.600 134.200 116.900 141.800 ;
        RECT 118.200 135.100 118.600 135.200 ;
        RECT 119.000 135.100 119.300 141.800 ;
        RECT 119.800 136.200 120.100 175.800 ;
        RECT 121.400 174.200 121.700 177.800 ;
        RECT 125.400 175.200 125.700 187.800 ;
        RECT 127.000 187.200 127.300 193.800 ;
        RECT 129.400 191.800 129.800 192.200 ;
        RECT 129.400 191.200 129.700 191.800 ;
        RECT 129.400 190.800 129.800 191.200 ;
        RECT 131.000 189.200 131.300 194.800 ;
        RECT 131.800 194.200 132.100 194.800 ;
        RECT 131.800 193.800 132.200 194.200 ;
        RECT 133.400 189.200 133.700 204.800 ;
        RECT 135.800 203.100 136.200 208.900 ;
        RECT 141.400 208.800 141.800 209.200 ;
        RECT 136.600 207.800 137.000 208.200 ;
        RECT 136.600 207.200 136.900 207.800 ;
        RECT 136.600 206.800 137.000 207.200 ;
        RECT 137.400 205.100 137.800 207.900 ;
        RECT 138.200 207.800 138.600 208.200 ;
        RECT 138.200 206.200 138.500 207.800 ;
        RECT 142.200 206.800 142.600 207.200 ;
        RECT 142.200 206.200 142.500 206.800 ;
        RECT 143.000 206.200 143.300 210.800 ;
        RECT 147.000 209.200 147.300 214.800 ;
        RECT 147.800 212.100 148.200 217.900 ;
        RECT 148.600 217.800 149.000 218.200 ;
        RECT 150.200 215.100 150.600 215.200 ;
        RECT 151.000 215.100 151.400 215.200 ;
        RECT 150.200 214.800 151.400 215.100 ;
        RECT 152.600 212.100 153.000 217.900 ;
        RECT 159.800 216.200 160.100 218.800 ;
        RECT 163.000 216.800 163.400 217.200 ;
        RECT 165.400 216.800 165.800 217.200 ;
        RECT 153.400 214.800 153.800 215.200 ;
        RECT 153.400 214.200 153.700 214.800 ;
        RECT 153.400 213.800 153.800 214.200 ;
        RECT 148.600 210.800 149.000 211.200 ;
        RECT 144.600 209.100 145.000 209.200 ;
        RECT 144.600 208.800 146.500 209.100 ;
        RECT 147.000 208.800 147.400 209.200 ;
        RECT 146.200 208.200 146.500 208.800 ;
        RECT 144.600 208.100 145.000 208.200 ;
        RECT 145.400 208.100 145.800 208.200 ;
        RECT 144.600 207.800 145.800 208.100 ;
        RECT 146.200 207.800 146.600 208.200 ;
        RECT 138.200 205.800 138.600 206.200 ;
        RECT 139.800 205.800 140.200 206.200 ;
        RECT 142.200 205.800 142.600 206.200 ;
        RECT 143.000 205.800 143.400 206.200 ;
        RECT 143.800 205.800 144.200 206.200 ;
        RECT 136.600 200.800 137.000 201.200 ;
        RECT 135.000 196.800 135.400 197.200 ;
        RECT 135.000 195.200 135.300 196.800 ;
        RECT 136.600 195.200 136.900 200.800 ;
        RECT 139.800 198.200 140.100 205.800 ;
        RECT 143.800 202.200 144.100 205.800 ;
        RECT 143.800 201.800 144.200 202.200 ;
        RECT 144.600 200.200 144.900 207.800 ;
        RECT 147.800 206.800 148.200 207.200 ;
        RECT 147.800 206.200 148.100 206.800 ;
        RECT 148.600 206.200 148.900 210.800 ;
        RECT 149.400 207.100 149.800 207.200 ;
        RECT 150.200 207.100 150.600 207.200 ;
        RECT 149.400 206.800 150.600 207.100 ;
        RECT 147.800 205.800 148.200 206.200 ;
        RECT 148.600 205.800 149.000 206.200 ;
        RECT 147.800 202.200 148.100 205.800 ;
        RECT 151.000 205.100 151.400 207.900 ;
        RECT 152.600 203.100 153.000 208.900 ;
        RECT 147.800 201.800 148.200 202.200 ;
        RECT 144.600 199.800 145.000 200.200 ;
        RECT 139.800 197.800 140.200 198.200 ;
        RECT 141.400 197.800 141.800 198.200 ;
        RECT 141.400 195.200 141.700 197.800 ;
        RECT 147.800 195.800 148.200 196.200 ;
        RECT 135.000 194.800 135.400 195.200 ;
        RECT 135.800 194.800 136.200 195.200 ;
        RECT 136.600 194.800 137.000 195.200 ;
        RECT 139.800 195.100 140.200 195.200 ;
        RECT 140.600 195.100 141.000 195.200 ;
        RECT 139.800 194.800 141.000 195.100 ;
        RECT 141.400 194.800 141.800 195.200 ;
        RECT 143.000 195.100 143.400 195.200 ;
        RECT 143.800 195.100 144.200 195.200 ;
        RECT 143.000 194.800 144.200 195.100 ;
        RECT 144.600 194.800 145.000 195.200 ;
        RECT 146.200 195.100 146.600 195.200 ;
        RECT 147.000 195.100 147.400 195.200 ;
        RECT 146.200 194.800 147.400 195.100 ;
        RECT 126.200 186.800 126.600 187.200 ;
        RECT 127.000 186.800 127.400 187.200 ;
        RECT 126.200 186.200 126.500 186.800 ;
        RECT 126.200 185.800 126.600 186.200 ;
        RECT 128.600 183.100 129.000 188.900 ;
        RECT 131.000 188.800 131.400 189.200 ;
        RECT 131.800 188.800 132.200 189.200 ;
        RECT 133.400 188.800 133.800 189.200 ;
        RECT 130.200 185.100 130.600 187.900 ;
        RECT 131.000 186.800 131.400 187.200 ;
        RECT 131.000 186.200 131.300 186.800 ;
        RECT 131.800 186.200 132.100 188.800 ;
        RECT 131.000 185.800 131.400 186.200 ;
        RECT 131.800 185.800 132.200 186.200 ;
        RECT 132.600 185.100 133.000 185.200 ;
        RECT 133.400 185.100 133.800 185.200 ;
        RECT 132.600 184.800 133.800 185.100 ;
        RECT 135.000 181.800 135.400 182.200 ;
        RECT 135.000 179.200 135.300 181.800 ;
        RECT 135.000 178.800 135.400 179.200 ;
        RECT 126.200 175.800 126.600 176.200 ;
        RECT 129.400 175.800 129.800 176.200 ;
        RECT 135.000 175.800 135.400 176.200 ;
        RECT 126.200 175.200 126.500 175.800 ;
        RECT 129.400 175.200 129.700 175.800 ;
        RECT 135.000 175.200 135.300 175.800 ;
        RECT 125.400 174.800 125.800 175.200 ;
        RECT 126.200 174.800 126.600 175.200 ;
        RECT 128.600 174.800 129.000 175.200 ;
        RECT 129.400 174.800 129.800 175.200 ;
        RECT 130.200 174.800 130.600 175.200 ;
        RECT 133.400 174.800 133.800 175.200 ;
        RECT 135.000 174.800 135.400 175.200 ;
        RECT 121.400 173.800 121.800 174.200 ;
        RECT 127.800 173.800 128.200 174.200 ;
        RECT 127.800 173.200 128.100 173.800 ;
        RECT 127.800 172.800 128.200 173.200 ;
        RECT 123.000 171.800 123.400 172.200 ;
        RECT 123.000 171.200 123.300 171.800 ;
        RECT 123.000 170.800 123.400 171.200 ;
        RECT 122.200 169.800 122.600 170.200 ;
        RECT 122.200 169.200 122.500 169.800 ;
        RECT 122.200 168.800 122.600 169.200 ;
        RECT 124.600 168.800 125.000 169.200 ;
        RECT 124.600 167.200 124.900 168.800 ;
        RECT 128.600 168.200 128.900 174.800 ;
        RECT 130.200 174.200 130.500 174.800 ;
        RECT 130.200 173.800 130.600 174.200 ;
        RECT 131.000 174.100 131.400 174.200 ;
        RECT 131.800 174.100 132.200 174.200 ;
        RECT 131.000 173.800 132.200 174.100 ;
        RECT 131.000 171.800 131.400 172.200 ;
        RECT 131.800 171.800 132.200 172.200 ;
        RECT 129.400 170.800 129.800 171.200 ;
        RECT 128.600 167.800 129.000 168.200 ;
        RECT 129.400 167.200 129.700 170.800 ;
        RECT 131.000 169.200 131.300 171.800 ;
        RECT 131.000 168.800 131.400 169.200 ;
        RECT 131.000 167.800 131.400 168.200 ;
        RECT 123.800 166.800 124.200 167.200 ;
        RECT 124.600 166.800 125.000 167.200 ;
        RECT 129.400 166.800 129.800 167.200 ;
        RECT 123.800 166.200 124.100 166.800 ;
        RECT 124.600 166.200 124.900 166.800 ;
        RECT 122.200 166.100 122.600 166.200 ;
        RECT 123.000 166.100 123.400 166.200 ;
        RECT 122.200 165.800 123.400 166.100 ;
        RECT 123.800 165.800 124.200 166.200 ;
        RECT 124.600 165.800 125.000 166.200 ;
        RECT 126.200 165.800 126.600 166.200 ;
        RECT 127.800 166.100 128.200 166.200 ;
        RECT 128.600 166.100 129.000 166.200 ;
        RECT 127.800 165.800 129.000 166.100 ;
        RECT 123.800 162.200 124.100 165.800 ;
        RECT 126.200 165.200 126.500 165.800 ;
        RECT 126.200 164.800 126.600 165.200 ;
        RECT 128.600 164.800 129.000 165.200 ;
        RECT 123.800 161.800 124.200 162.200 ;
        RECT 120.600 152.100 121.000 157.900 ;
        RECT 126.200 157.200 126.500 164.800 ;
        RECT 128.600 164.200 128.900 164.800 ;
        RECT 128.600 163.800 129.000 164.200 ;
        RECT 129.400 160.100 129.700 166.800 ;
        RECT 130.200 164.800 130.600 165.200 ;
        RECT 130.200 163.200 130.500 164.800 ;
        RECT 130.200 162.800 130.600 163.200 ;
        RECT 128.600 159.800 129.700 160.100 ;
        RECT 123.800 156.800 124.200 157.200 ;
        RECT 126.200 156.800 126.600 157.200 ;
        RECT 123.800 155.200 124.100 156.800 ;
        RECT 124.600 156.100 125.000 156.200 ;
        RECT 125.400 156.100 125.800 156.200 ;
        RECT 124.600 155.800 125.800 156.100 ;
        RECT 127.800 155.800 128.200 156.200 ;
        RECT 127.800 155.200 128.100 155.800 ;
        RECT 123.800 154.800 124.200 155.200 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 123.800 154.200 124.100 154.800 ;
        RECT 128.600 154.200 128.900 159.800 ;
        RECT 131.000 159.200 131.300 167.800 ;
        RECT 131.800 167.200 132.100 171.800 ;
        RECT 132.600 169.800 133.000 170.200 ;
        RECT 132.600 169.200 132.900 169.800 ;
        RECT 132.600 168.800 133.000 169.200 ;
        RECT 131.800 166.800 132.200 167.200 ;
        RECT 133.400 159.200 133.700 174.800 ;
        RECT 135.000 163.100 135.400 168.900 ;
        RECT 135.800 159.200 136.100 194.800 ;
        RECT 144.600 194.200 144.900 194.800 ;
        RECT 137.400 193.800 137.800 194.200 ;
        RECT 144.600 193.800 145.000 194.200 ;
        RECT 145.400 194.100 145.800 194.200 ;
        RECT 145.400 193.800 146.500 194.100 ;
        RECT 137.400 193.200 137.700 193.800 ;
        RECT 137.400 192.800 137.800 193.200 ;
        RECT 139.000 191.800 139.400 192.200 ;
        RECT 141.400 191.800 141.800 192.200 ;
        RECT 139.000 184.200 139.300 191.800 ;
        RECT 141.400 188.200 141.700 191.800 ;
        RECT 144.600 189.800 145.000 190.200 ;
        RECT 144.600 189.200 144.900 189.800 ;
        RECT 144.600 188.800 145.000 189.200 ;
        RECT 141.400 187.800 141.800 188.200 ;
        RECT 139.800 187.100 140.200 187.200 ;
        RECT 140.600 187.100 141.000 187.200 ;
        RECT 139.800 186.800 141.000 187.100 ;
        RECT 143.000 186.800 143.400 187.200 ;
        RECT 144.600 187.100 145.000 187.200 ;
        RECT 145.400 187.100 145.800 187.200 ;
        RECT 144.600 186.800 145.800 187.100 ;
        RECT 143.000 186.200 143.300 186.800 ;
        RECT 146.200 186.200 146.500 193.800 ;
        RECT 147.800 193.200 148.100 195.800 ;
        RECT 148.600 194.100 149.000 194.200 ;
        RECT 149.400 194.100 149.800 194.200 ;
        RECT 148.600 193.800 149.800 194.100 ;
        RECT 147.800 192.800 148.200 193.200 ;
        RECT 150.200 193.100 150.600 195.900 ;
        RECT 151.800 192.100 152.200 197.900 ;
        RECT 152.600 194.700 153.000 195.100 ;
        RECT 152.600 194.200 152.900 194.700 ;
        RECT 153.400 194.200 153.700 213.800 ;
        RECT 154.200 213.100 154.600 215.900 ;
        RECT 157.400 215.800 157.800 216.200 ;
        RECT 159.000 216.100 159.400 216.200 ;
        RECT 159.800 216.100 160.200 216.200 ;
        RECT 159.000 215.800 160.200 216.100 ;
        RECT 157.400 215.200 157.700 215.800 ;
        RECT 163.000 215.200 163.300 216.800 ;
        RECT 165.400 216.200 165.700 216.800 ;
        RECT 165.400 215.800 165.800 216.200 ;
        RECT 166.200 215.200 166.500 221.800 ;
        RECT 157.400 214.800 157.800 215.200 ;
        RECT 163.000 214.800 163.400 215.200 ;
        RECT 166.200 214.800 166.600 215.200 ;
        RECT 156.600 213.800 157.000 214.200 ;
        RECT 161.400 213.800 161.800 214.200 ;
        RECT 162.200 213.800 162.600 214.200 ;
        RECT 164.600 214.100 165.000 214.200 ;
        RECT 165.400 214.100 165.800 214.200 ;
        RECT 164.600 213.800 165.800 214.100 ;
        RECT 167.000 213.800 167.400 214.200 ;
        RECT 156.600 211.200 156.900 213.800 ;
        RECT 159.000 211.800 159.400 212.200 ;
        RECT 156.600 210.800 157.000 211.200 ;
        RECT 154.200 206.800 154.600 207.200 ;
        RECT 154.200 206.200 154.500 206.800 ;
        RECT 154.200 205.800 154.600 206.200 ;
        RECT 156.600 205.800 157.000 206.200 ;
        RECT 156.600 201.200 156.900 205.800 ;
        RECT 157.400 203.100 157.800 208.900 ;
        RECT 159.000 207.200 159.300 211.800 ;
        RECT 160.600 209.800 161.000 210.200 ;
        RECT 159.800 208.800 160.200 209.200 ;
        RECT 159.800 208.200 160.100 208.800 ;
        RECT 159.800 207.800 160.200 208.200 ;
        RECT 159.000 206.800 159.400 207.200 ;
        RECT 160.600 206.200 160.900 209.800 ;
        RECT 161.400 208.200 161.700 213.800 ;
        RECT 162.200 211.200 162.500 213.800 ;
        RECT 167.000 212.200 167.300 213.800 ;
        RECT 167.800 213.100 168.200 215.900 ;
        RECT 168.600 214.800 169.000 215.200 ;
        RECT 168.600 214.200 168.900 214.800 ;
        RECT 168.600 213.800 169.000 214.200 ;
        RECT 167.000 211.800 167.400 212.200 ;
        RECT 169.400 212.100 169.800 217.900 ;
        RECT 170.200 214.700 170.600 215.100 ;
        RECT 170.200 214.200 170.500 214.700 ;
        RECT 170.200 213.800 170.600 214.200 ;
        RECT 174.200 212.100 174.600 217.900 ;
        RECT 162.200 210.800 162.600 211.200 ;
        RECT 165.400 210.800 165.800 211.200 ;
        RECT 161.400 207.800 161.800 208.200 ;
        RECT 161.400 206.200 161.700 207.800 ;
        RECT 165.400 207.200 165.700 210.800 ;
        RECT 167.000 207.200 167.300 211.800 ;
        RECT 170.200 207.800 170.600 208.200 ;
        RECT 170.200 207.200 170.500 207.800 ;
        RECT 163.800 206.800 164.200 207.200 ;
        RECT 165.400 206.800 165.800 207.200 ;
        RECT 167.000 206.800 167.400 207.200 ;
        RECT 167.800 207.100 168.200 207.200 ;
        RECT 168.600 207.100 169.000 207.200 ;
        RECT 167.800 206.800 169.000 207.100 ;
        RECT 170.200 206.800 170.600 207.200 ;
        RECT 163.800 206.200 164.100 206.800 ;
        RECT 160.600 205.800 161.000 206.200 ;
        RECT 161.400 205.800 161.800 206.200 ;
        RECT 163.800 205.800 164.200 206.200 ;
        RECT 166.200 205.800 166.600 206.200 ;
        RECT 156.600 200.800 157.000 201.200 ;
        RECT 160.600 199.200 160.900 205.800 ;
        RECT 166.200 204.200 166.500 205.800 ;
        RECT 168.600 204.800 169.000 205.200 ;
        RECT 171.000 205.100 171.400 207.900 ;
        RECT 171.800 206.800 172.200 207.200 ;
        RECT 168.600 204.200 168.900 204.800 ;
        RECT 166.200 203.800 166.600 204.200 ;
        RECT 168.600 203.800 169.000 204.200 ;
        RECT 163.000 201.800 163.400 202.200 ;
        RECT 161.400 200.800 161.800 201.200 ;
        RECT 160.600 198.800 161.000 199.200 ;
        RECT 152.600 193.800 153.000 194.200 ;
        RECT 153.400 193.800 153.800 194.200 ;
        RECT 155.800 193.800 156.200 194.200 ;
        RECT 153.400 190.800 153.800 191.200 ;
        RECT 147.000 189.100 147.400 189.200 ;
        RECT 147.800 189.100 148.200 189.200 ;
        RECT 147.000 188.800 148.200 189.100 ;
        RECT 148.600 188.800 149.000 189.200 ;
        RECT 151.800 189.100 152.200 189.200 ;
        RECT 152.600 189.100 153.000 189.200 ;
        RECT 151.800 188.800 153.000 189.100 ;
        RECT 148.600 187.200 148.900 188.800 ;
        RECT 153.400 187.200 153.700 190.800 ;
        RECT 155.000 187.800 155.400 188.200 ;
        RECT 148.600 186.800 149.000 187.200 ;
        RECT 151.800 187.100 152.200 187.200 ;
        RECT 152.600 187.100 153.000 187.200 ;
        RECT 151.800 186.800 153.000 187.100 ;
        RECT 153.400 186.800 153.800 187.200 ;
        RECT 154.200 186.800 154.600 187.200 ;
        RECT 154.200 186.200 154.500 186.800 ;
        RECT 155.000 186.200 155.300 187.800 ;
        RECT 141.400 185.800 141.800 186.200 ;
        RECT 143.000 185.800 143.400 186.200 ;
        RECT 146.200 185.800 146.600 186.200 ;
        RECT 150.200 186.100 150.600 186.200 ;
        RECT 151.000 186.100 151.400 186.200 ;
        RECT 150.200 185.800 151.400 186.100 ;
        RECT 154.200 185.800 154.600 186.200 ;
        RECT 155.000 185.800 155.400 186.200 ;
        RECT 139.000 183.800 139.400 184.200 ;
        RECT 138.200 179.800 138.600 180.200 ;
        RECT 138.200 175.200 138.500 179.800 ;
        RECT 141.400 179.200 141.700 185.800 ;
        RECT 143.000 181.200 143.300 185.800 ;
        RECT 146.200 185.200 146.500 185.800 ;
        RECT 146.200 184.800 146.600 185.200 ;
        RECT 147.000 184.800 147.400 185.200 ;
        RECT 147.000 184.200 147.300 184.800 ;
        RECT 147.000 183.800 147.400 184.200 ;
        RECT 147.800 183.800 148.200 184.200 ;
        RECT 143.000 180.800 143.400 181.200 ;
        RECT 141.400 178.800 141.800 179.200 ;
        RECT 147.800 176.100 148.100 183.800 ;
        RECT 155.800 179.200 156.100 193.800 ;
        RECT 156.600 192.100 157.000 197.900 ;
        RECT 161.400 197.200 161.700 200.800 ;
        RECT 163.000 198.200 163.300 201.800 ;
        RECT 159.800 197.100 160.200 197.200 ;
        RECT 160.600 197.100 161.000 197.200 ;
        RECT 159.800 196.800 161.000 197.100 ;
        RECT 161.400 196.800 161.800 197.200 ;
        RECT 157.400 194.800 157.800 195.200 ;
        RECT 157.400 185.200 157.700 194.800 ;
        RECT 158.200 192.800 158.600 193.200 ;
        RECT 158.200 189.200 158.500 192.800 ;
        RECT 159.000 192.100 159.400 192.200 ;
        RECT 162.200 192.100 162.600 197.900 ;
        RECT 163.000 197.800 163.400 198.200 ;
        RECT 166.200 197.800 166.600 198.200 ;
        RECT 166.200 195.100 166.500 197.800 ;
        RECT 166.200 194.700 166.600 195.100 ;
        RECT 167.000 192.100 167.400 197.900 ;
        RECT 169.400 196.800 169.800 197.200 ;
        RECT 167.800 193.800 168.200 194.200 ;
        RECT 159.000 191.800 160.100 192.100 ;
        RECT 158.200 188.800 158.600 189.200 ;
        RECT 159.800 187.200 160.100 191.800 ;
        RECT 160.600 188.800 161.000 189.200 ;
        RECT 165.400 189.100 165.800 189.200 ;
        RECT 166.200 189.100 166.600 189.200 ;
        RECT 165.400 188.800 166.600 189.100 ;
        RECT 160.600 187.200 160.900 188.800 ;
        RECT 158.200 186.800 158.600 187.200 ;
        RECT 159.800 186.800 160.200 187.200 ;
        RECT 160.600 186.800 161.000 187.200 ;
        RECT 162.200 187.100 162.600 187.200 ;
        RECT 163.000 187.100 163.400 187.200 ;
        RECT 162.200 186.800 163.400 187.100 ;
        RECT 165.400 186.800 165.800 187.200 ;
        RECT 158.200 186.200 158.500 186.800 ;
        RECT 158.200 185.800 158.600 186.200 ;
        RECT 156.600 184.800 157.000 185.200 ;
        RECT 157.400 185.100 157.800 185.200 ;
        RECT 158.200 185.100 158.600 185.200 ;
        RECT 157.400 184.800 158.600 185.100 ;
        RECT 156.600 182.200 156.900 184.800 ;
        RECT 156.600 181.800 157.000 182.200 ;
        RECT 151.800 178.800 152.200 179.200 ;
        RECT 155.800 178.800 156.200 179.200 ;
        RECT 147.000 175.800 148.100 176.100 ;
        RECT 149.400 176.100 149.800 176.200 ;
        RECT 150.200 176.100 150.600 176.200 ;
        RECT 149.400 175.800 150.600 176.100 ;
        RECT 147.000 175.200 147.300 175.800 ;
        RECT 137.400 174.800 137.800 175.200 ;
        RECT 138.200 174.800 138.600 175.200 ;
        RECT 139.800 174.800 140.200 175.200 ;
        RECT 142.200 174.800 142.600 175.200 ;
        RECT 143.000 174.800 143.400 175.200 ;
        RECT 143.800 174.800 144.200 175.200 ;
        RECT 144.600 175.100 145.000 175.200 ;
        RECT 145.400 175.100 145.800 175.200 ;
        RECT 144.600 174.800 145.800 175.100 ;
        RECT 147.000 174.800 147.400 175.200 ;
        RECT 147.800 174.800 148.200 175.200 ;
        RECT 148.600 174.800 149.000 175.200 ;
        RECT 137.400 174.200 137.700 174.800 ;
        RECT 137.400 173.800 137.800 174.200 ;
        RECT 139.800 172.200 140.100 174.800 ;
        RECT 142.200 173.200 142.500 174.800 ;
        RECT 142.200 172.800 142.600 173.200 ;
        RECT 139.800 171.800 140.200 172.200 ;
        RECT 137.400 166.800 137.800 167.200 ;
        RECT 129.400 158.800 129.800 159.200 ;
        RECT 131.000 158.800 131.400 159.200 ;
        RECT 133.400 158.800 133.800 159.200 ;
        RECT 135.800 158.800 136.200 159.200 ;
        RECT 129.400 155.200 129.700 158.800 ;
        RECT 130.200 155.800 130.600 156.200 ;
        RECT 130.200 155.200 130.500 155.800 ;
        RECT 129.400 154.800 129.800 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 132.600 155.100 133.000 155.200 ;
        RECT 133.400 155.100 133.800 155.200 ;
        RECT 132.600 154.800 133.800 155.100 ;
        RECT 123.800 153.800 124.200 154.200 ;
        RECT 125.400 154.100 125.800 154.200 ;
        RECT 126.200 154.100 126.600 154.200 ;
        RECT 125.400 153.800 126.600 154.100 ;
        RECT 128.600 153.800 129.000 154.200 ;
        RECT 124.600 151.800 125.000 152.200 ;
        RECT 121.400 149.800 121.800 150.200 ;
        RECT 121.400 146.200 121.700 149.800 ;
        RECT 121.400 145.800 121.800 146.200 ;
        RECT 121.400 144.800 121.800 145.200 ;
        RECT 122.200 145.100 122.600 147.900 ;
        RECT 123.000 147.800 123.400 148.200 ;
        RECT 123.000 147.200 123.300 147.800 ;
        RECT 123.000 146.800 123.400 147.200 ;
        RECT 120.600 137.800 121.000 138.200 ;
        RECT 119.800 135.800 120.200 136.200 ;
        RECT 118.200 134.800 119.300 135.100 ;
        RECT 120.600 135.200 120.900 137.800 ;
        RECT 121.400 135.200 121.700 144.800 ;
        RECT 120.600 134.800 121.000 135.200 ;
        RECT 121.400 134.800 121.800 135.200 ;
        RECT 116.600 133.800 117.000 134.200 ;
        RECT 119.000 131.800 119.400 132.200 ;
        RECT 115.800 129.800 116.200 130.200 ;
        RECT 119.000 128.200 119.300 131.800 ;
        RECT 119.800 128.800 120.200 129.200 ;
        RECT 119.000 127.800 119.400 128.200 ;
        RECT 119.800 127.200 120.100 128.800 ;
        RECT 114.200 127.100 114.600 127.200 ;
        RECT 115.000 127.100 115.400 127.200 ;
        RECT 114.200 126.800 115.400 127.100 ;
        RECT 118.200 126.800 118.600 127.200 ;
        RECT 119.800 126.800 120.200 127.200 ;
        RECT 118.200 126.200 118.500 126.800 ;
        RECT 108.600 125.800 109.000 126.200 ;
        RECT 109.400 125.800 109.800 126.200 ;
        RECT 110.200 125.800 110.600 126.200 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 114.200 125.800 114.600 126.200 ;
        RECT 115.000 125.800 115.400 126.200 ;
        RECT 118.200 125.800 118.600 126.200 ;
        RECT 111.000 125.200 111.300 125.800 ;
        RECT 111.000 124.800 111.400 125.200 ;
        RECT 110.200 121.800 110.600 122.200 ;
        RECT 110.200 119.200 110.500 121.800 ;
        RECT 114.200 119.200 114.500 125.800 ;
        RECT 115.000 125.200 115.300 125.800 ;
        RECT 115.000 124.800 115.400 125.200 ;
        RECT 117.400 125.100 117.800 125.200 ;
        RECT 118.200 125.100 118.600 125.200 ;
        RECT 120.600 125.100 121.000 127.900 ;
        RECT 117.400 124.800 118.600 125.100 ;
        RECT 110.200 118.800 110.600 119.200 ;
        RECT 114.200 118.800 114.600 119.200 ;
        RECT 109.400 117.800 109.800 118.200 ;
        RECT 106.200 116.100 106.600 116.200 ;
        RECT 107.000 116.100 107.400 116.200 ;
        RECT 106.200 115.800 107.400 116.100 ;
        RECT 108.600 115.800 109.000 116.200 ;
        RECT 108.600 115.200 108.900 115.800 ;
        RECT 104.600 113.800 105.700 114.100 ;
        RECT 107.800 114.800 108.200 115.200 ;
        RECT 108.600 114.800 109.000 115.200 ;
        RECT 107.800 114.200 108.100 114.800 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 104.600 112.800 105.000 113.200 ;
        RECT 100.600 111.800 101.000 112.200 ;
        RECT 103.800 111.800 104.200 112.200 ;
        RECT 100.600 109.200 100.900 111.800 ;
        RECT 103.800 110.800 104.200 111.200 ;
        RECT 100.600 108.800 101.000 109.200 ;
        RECT 103.800 107.200 104.100 110.800 ;
        RECT 97.400 106.800 97.800 107.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 103.800 106.800 104.200 107.200 ;
        RECT 96.600 104.800 97.000 105.200 ;
        RECT 97.400 104.800 97.800 105.200 ;
        RECT 98.200 105.100 98.600 105.200 ;
        RECT 99.000 105.100 99.400 105.200 ;
        RECT 98.200 104.800 99.400 105.100 ;
        RECT 95.000 101.800 95.400 102.200 ;
        RECT 95.000 101.200 95.300 101.800 ;
        RECT 95.000 100.800 95.400 101.200 ;
        RECT 93.400 99.800 93.800 100.200 ;
        RECT 95.000 99.800 95.400 100.200 ;
        RECT 93.400 99.200 93.700 99.800 ;
        RECT 95.000 99.200 95.300 99.800 ;
        RECT 93.400 98.800 93.800 99.200 ;
        RECT 95.000 98.800 95.400 99.200 ;
        RECT 94.200 95.800 94.600 96.200 ;
        RECT 95.800 96.100 96.200 96.200 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 95.800 95.800 97.000 96.100 ;
        RECT 94.200 89.200 94.500 95.800 ;
        RECT 95.800 94.800 96.200 95.200 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 95.000 91.800 95.400 92.200 ;
        RECT 94.200 88.800 94.600 89.200 ;
        RECT 94.200 87.200 94.500 88.800 ;
        RECT 94.200 86.800 94.600 87.200 ;
        RECT 91.800 85.800 92.200 86.200 ;
        RECT 94.200 85.800 94.600 86.200 ;
        RECT 87.000 84.800 87.400 85.200 ;
        RECT 88.600 84.800 89.000 85.200 ;
        RECT 89.400 84.800 89.800 85.200 ;
        RECT 91.800 84.800 92.200 85.200 ;
        RECT 86.200 83.800 86.600 84.200 ;
        RECT 82.200 82.800 82.600 83.200 ;
        RECT 83.000 81.800 83.400 82.200 ;
        RECT 81.400 76.800 81.800 77.200 ;
        RECT 81.400 75.200 81.700 76.800 ;
        RECT 81.400 74.800 81.800 75.200 ;
        RECT 80.600 73.800 81.000 74.200 ;
        RECT 83.000 71.200 83.300 81.800 ;
        RECT 84.600 72.100 85.000 77.900 ;
        RECT 85.400 72.800 85.800 73.200 ;
        RECT 87.000 73.100 87.300 84.800 ;
        RECT 88.600 82.200 88.900 84.800 ;
        RECT 88.600 81.800 89.000 82.200 ;
        RECT 87.800 77.800 88.200 78.200 ;
        RECT 88.600 77.800 89.000 78.200 ;
        RECT 87.800 75.200 88.100 77.800 ;
        RECT 87.800 74.800 88.200 75.200 ;
        RECT 88.600 74.200 88.900 77.800 ;
        RECT 89.400 74.200 89.700 84.800 ;
        RECT 91.000 83.800 91.400 84.200 ;
        RECT 91.000 78.200 91.300 83.800 ;
        RECT 91.000 77.800 91.400 78.200 ;
        RECT 91.000 76.800 91.400 77.200 ;
        RECT 91.000 75.200 91.300 76.800 ;
        RECT 91.800 76.200 92.100 84.800 ;
        RECT 92.600 81.800 93.000 82.200 ;
        RECT 92.600 81.200 92.900 81.800 ;
        RECT 92.600 80.800 93.000 81.200 ;
        RECT 94.200 77.200 94.500 85.800 ;
        RECT 95.000 82.200 95.300 91.800 ;
        RECT 95.800 89.200 96.100 94.800 ;
        RECT 96.600 94.200 96.900 94.800 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 96.600 92.200 96.900 93.800 ;
        RECT 96.600 91.800 97.000 92.200 ;
        RECT 96.600 89.800 97.000 90.200 ;
        RECT 96.600 89.200 96.900 89.800 ;
        RECT 97.400 89.200 97.700 104.800 ;
        RECT 98.200 101.800 98.600 102.200 ;
        RECT 98.200 98.200 98.500 101.800 ;
        RECT 99.800 99.200 100.100 106.800 ;
        RECT 103.800 106.200 104.100 106.800 ;
        RECT 103.800 105.800 104.200 106.200 ;
        RECT 100.600 104.800 101.000 105.200 ;
        RECT 103.000 105.100 103.400 105.200 ;
        RECT 103.800 105.100 104.200 105.200 ;
        RECT 103.000 104.800 104.200 105.100 ;
        RECT 99.800 98.800 100.200 99.200 ;
        RECT 98.200 97.800 98.600 98.200 ;
        RECT 98.200 94.200 98.500 97.800 ;
        RECT 99.800 96.800 100.200 97.200 ;
        RECT 99.800 94.200 100.100 96.800 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 99.800 93.800 100.200 94.200 ;
        RECT 95.800 88.800 96.200 89.200 ;
        RECT 96.600 88.800 97.000 89.200 ;
        RECT 97.400 88.800 97.800 89.200 ;
        RECT 95.800 87.100 96.100 88.800 ;
        RECT 100.600 87.200 100.900 104.800 ;
        RECT 101.400 103.800 101.800 104.200 ;
        RECT 101.400 95.200 101.700 103.800 ;
        RECT 102.200 95.800 102.600 96.200 ;
        RECT 103.000 95.800 103.400 96.200 ;
        RECT 102.200 95.200 102.500 95.800 ;
        RECT 103.000 95.200 103.300 95.800 ;
        RECT 101.400 94.800 101.800 95.200 ;
        RECT 102.200 94.800 102.600 95.200 ;
        RECT 103.000 94.800 103.400 95.200 ;
        RECT 102.200 94.100 102.600 94.200 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 102.200 93.800 103.400 94.100 ;
        RECT 103.800 93.100 104.200 95.900 ;
        RECT 102.200 90.800 102.600 91.200 ;
        RECT 102.200 89.200 102.500 90.800 ;
        RECT 104.600 89.200 104.900 112.800 ;
        RECT 105.400 111.800 105.800 112.200 ;
        RECT 107.800 111.800 108.200 112.200 ;
        RECT 105.400 110.200 105.700 111.800 ;
        RECT 105.400 109.800 105.800 110.200 ;
        RECT 105.400 107.200 105.700 109.800 ;
        RECT 107.800 109.200 108.100 111.800 ;
        RECT 108.600 109.200 108.900 114.800 ;
        RECT 109.400 114.200 109.700 117.800 ;
        RECT 109.400 113.800 109.800 114.200 ;
        RECT 112.600 112.100 113.000 117.900 ;
        RECT 113.400 115.100 113.800 115.200 ;
        RECT 114.200 115.100 114.600 115.200 ;
        RECT 113.400 114.800 114.600 115.100 ;
        RECT 115.000 113.200 115.300 124.800 ;
        RECT 115.800 121.800 116.200 122.200 ;
        RECT 115.800 121.200 116.100 121.800 ;
        RECT 121.400 121.200 121.700 134.800 ;
        RECT 122.200 133.800 122.600 134.200 ;
        RECT 122.200 132.200 122.500 133.800 ;
        RECT 122.200 131.800 122.600 132.200 ;
        RECT 122.200 123.100 122.600 128.900 ;
        RECT 123.000 128.200 123.300 146.800 ;
        RECT 123.800 143.100 124.200 148.900 ;
        RECT 124.600 146.300 124.900 151.800 ;
        RECT 124.600 145.900 125.000 146.300 ;
        RECT 124.600 145.800 124.900 145.900 ;
        RECT 128.600 143.100 129.000 148.900 ;
        RECT 129.400 147.200 129.700 154.800 ;
        RECT 134.200 153.100 134.600 155.900 ;
        RECT 135.800 152.100 136.200 157.900 ;
        RECT 137.400 154.200 137.700 166.800 ;
        RECT 138.200 165.800 138.600 166.200 ;
        RECT 138.200 165.200 138.500 165.800 ;
        RECT 138.200 164.800 138.600 165.200 ;
        RECT 139.800 163.100 140.200 168.900 ;
        RECT 141.400 165.100 141.800 167.900 ;
        RECT 142.200 167.800 142.600 168.200 ;
        RECT 142.200 167.200 142.500 167.800 ;
        RECT 142.200 166.800 142.600 167.200 ;
        RECT 142.200 165.800 142.600 166.200 ;
        RECT 142.200 165.200 142.500 165.800 ;
        RECT 142.200 164.800 142.600 165.200 ;
        RECT 138.200 154.800 138.600 155.200 ;
        RECT 139.800 154.800 140.200 155.200 ;
        RECT 137.400 153.800 137.800 154.200 ;
        RECT 135.800 150.800 136.200 151.200 ;
        RECT 131.000 149.800 131.400 150.200 ;
        RECT 131.000 149.200 131.300 149.800 ;
        RECT 131.000 148.800 131.400 149.200 ;
        RECT 132.600 148.800 133.000 149.200 ;
        RECT 129.400 146.800 129.800 147.200 ;
        RECT 132.600 146.200 132.900 148.800 ;
        RECT 135.000 147.800 135.400 148.200 ;
        RECT 135.000 146.200 135.300 147.800 ;
        RECT 135.800 146.200 136.100 150.800 ;
        RECT 138.200 149.200 138.500 154.800 ;
        RECT 139.800 151.200 140.100 154.800 ;
        RECT 140.600 152.100 141.000 157.900 ;
        RECT 142.200 156.200 142.500 164.800 ;
        RECT 143.000 163.200 143.300 174.800 ;
        RECT 143.800 174.200 144.100 174.800 ;
        RECT 143.800 173.800 144.200 174.200 ;
        RECT 147.800 171.200 148.100 174.800 ;
        RECT 148.600 174.200 148.900 174.800 ;
        RECT 148.600 173.800 149.000 174.200 ;
        RECT 147.800 170.800 148.200 171.200 ;
        RECT 144.600 166.800 145.000 167.200 ;
        RECT 144.600 166.200 144.900 166.800 ;
        RECT 144.600 165.800 145.000 166.200 ;
        RECT 144.600 164.800 145.000 165.200 ;
        RECT 143.000 162.800 143.400 163.200 ;
        RECT 144.600 159.200 144.900 164.800 ;
        RECT 147.800 163.100 148.200 168.900 ;
        RECT 151.800 168.200 152.100 178.800 ;
        RECT 155.800 176.800 156.200 177.200 ;
        RECT 154.200 176.100 154.600 176.200 ;
        RECT 155.000 176.100 155.400 176.200 ;
        RECT 154.200 175.800 155.400 176.100 ;
        RECT 153.400 175.100 153.800 175.200 ;
        RECT 154.200 175.100 154.600 175.200 ;
        RECT 153.400 174.800 154.600 175.100 ;
        RECT 155.000 174.800 155.400 175.200 ;
        RECT 155.000 174.200 155.300 174.800 ;
        RECT 155.800 174.200 156.100 176.800 ;
        RECT 156.600 175.200 156.900 181.800 ;
        RECT 159.000 178.800 159.400 179.200 ;
        RECT 156.600 174.800 157.000 175.200 ;
        RECT 155.000 173.800 155.400 174.200 ;
        RECT 155.800 173.800 156.200 174.200 ;
        RECT 158.200 172.100 158.600 177.900 ;
        RECT 159.000 175.200 159.300 178.800 ;
        RECT 159.800 176.200 160.100 186.800 ;
        RECT 160.600 184.200 160.900 186.800 ;
        RECT 165.400 186.200 165.700 186.800 ;
        RECT 161.400 185.800 161.800 186.200 ;
        RECT 165.400 185.800 165.800 186.200 ;
        RECT 161.400 185.200 161.700 185.800 ;
        RECT 161.400 184.800 161.800 185.200 ;
        RECT 164.600 185.100 165.000 185.200 ;
        RECT 165.400 185.100 165.800 185.200 ;
        RECT 164.600 184.800 165.800 185.100 ;
        RECT 167.800 184.200 168.100 193.800 ;
        RECT 168.600 193.100 169.000 195.900 ;
        RECT 169.400 194.200 169.700 196.800 ;
        RECT 171.000 195.800 171.400 196.200 ;
        RECT 171.000 195.200 171.300 195.800 ;
        RECT 171.000 194.800 171.400 195.200 ;
        RECT 169.400 193.800 169.800 194.200 ;
        RECT 160.600 183.800 161.000 184.200 ;
        RECT 162.200 183.800 162.600 184.200 ;
        RECT 167.800 183.800 168.200 184.200 ;
        RECT 162.200 182.200 162.500 183.800 ;
        RECT 168.600 183.100 169.000 188.900 ;
        RECT 169.400 186.100 169.800 186.200 ;
        RECT 170.200 186.100 170.600 186.200 ;
        RECT 169.400 185.800 170.600 186.100 ;
        RECT 162.200 181.800 162.600 182.200 ;
        RECT 159.800 175.800 160.200 176.200 ;
        RECT 159.000 174.800 159.400 175.200 ;
        RECT 160.600 175.100 161.000 175.200 ;
        RECT 161.400 175.100 161.800 175.200 ;
        RECT 160.600 174.800 161.800 175.100 ;
        RECT 163.000 172.100 163.400 177.900 ;
        RECT 164.600 173.100 165.000 175.900 ;
        RECT 166.200 175.800 166.600 176.200 ;
        RECT 168.600 175.800 169.000 176.200 ;
        RECT 166.200 175.200 166.500 175.800 ;
        RECT 168.600 175.200 168.900 175.800 ;
        RECT 166.200 174.800 166.600 175.200 ;
        RECT 168.600 174.800 169.000 175.200 ;
        RECT 169.400 174.800 169.800 175.200 ;
        RECT 170.200 174.800 170.600 175.200 ;
        RECT 165.400 173.800 165.800 174.200 ;
        RECT 165.400 173.200 165.700 173.800 ;
        RECT 169.400 173.200 169.700 174.800 ;
        RECT 170.200 174.200 170.500 174.800 ;
        RECT 171.000 174.200 171.300 194.800 ;
        RECT 171.800 187.200 172.100 206.800 ;
        RECT 172.600 203.100 173.000 208.900 ;
        RECT 173.400 206.800 173.800 207.200 ;
        RECT 173.400 206.300 173.700 206.800 ;
        RECT 173.400 205.900 173.800 206.300 ;
        RECT 172.600 200.800 173.000 201.200 ;
        RECT 172.600 195.200 172.900 200.800 ;
        RECT 175.800 199.200 176.100 224.800 ;
        RECT 179.000 223.100 179.400 228.900 ;
        RECT 181.400 228.800 182.600 229.100 ;
        RECT 183.000 226.800 183.400 227.200 ;
        RECT 183.000 226.200 183.300 226.800 ;
        RECT 182.200 225.800 182.600 226.200 ;
        RECT 183.000 225.800 183.400 226.200 ;
        RECT 182.200 225.200 182.500 225.800 ;
        RECT 182.200 224.800 182.600 225.200 ;
        RECT 185.400 224.200 185.700 233.800 ;
        RECT 187.800 232.100 188.200 237.900 ;
        RECT 191.800 236.800 192.200 237.200 ;
        RECT 191.800 236.200 192.100 236.800 ;
        RECT 191.800 235.800 192.200 236.200 ;
        RECT 193.400 235.800 193.800 236.200 ;
        RECT 193.400 235.200 193.700 235.800 ;
        RECT 191.000 235.100 191.400 235.200 ;
        RECT 191.800 235.100 192.200 235.200 ;
        RECT 191.000 234.800 192.200 235.100 ;
        RECT 193.400 234.800 193.800 235.200 ;
        RECT 188.600 233.800 189.000 234.200 ;
        RECT 191.000 233.800 191.400 234.200 ;
        RECT 187.800 229.800 188.200 230.200 ;
        RECT 186.200 228.800 186.600 229.200 ;
        RECT 186.200 226.200 186.500 228.800 ;
        RECT 187.800 226.200 188.100 229.800 ;
        RECT 186.200 225.800 186.600 226.200 ;
        RECT 187.800 225.800 188.200 226.200 ;
        RECT 185.400 223.800 185.800 224.200 ;
        RECT 183.000 222.800 183.400 223.200 ;
        RECT 178.200 221.800 178.600 222.200 ;
        RECT 178.200 219.200 178.500 221.800 ;
        RECT 183.000 219.200 183.300 222.800 ;
        RECT 184.600 221.800 185.000 222.200 ;
        RECT 178.200 218.800 178.600 219.200 ;
        RECT 183.000 218.800 183.400 219.200 ;
        RECT 179.800 215.100 180.200 215.200 ;
        RECT 180.600 215.100 181.000 215.200 ;
        RECT 179.800 214.800 181.000 215.100 ;
        RECT 181.400 213.800 181.800 214.200 ;
        RECT 176.600 211.800 177.000 212.200 ;
        RECT 176.600 211.200 176.900 211.800 ;
        RECT 176.600 210.800 177.000 211.200 ;
        RECT 181.400 209.200 181.700 213.800 ;
        RECT 182.200 211.800 182.600 212.200 ;
        RECT 176.600 207.800 177.000 208.200 ;
        RECT 175.800 198.800 176.200 199.200 ;
        RECT 173.400 197.800 173.800 198.200 ;
        RECT 173.400 197.200 173.700 197.800 ;
        RECT 173.400 196.800 173.800 197.200 ;
        RECT 172.600 195.100 173.000 195.200 ;
        RECT 173.400 195.100 173.800 195.200 ;
        RECT 172.600 194.800 173.800 195.100 ;
        RECT 174.200 193.800 174.600 194.200 ;
        RECT 171.800 186.800 172.200 187.200 ;
        RECT 173.400 183.100 173.800 188.900 ;
        RECT 174.200 188.200 174.500 193.800 ;
        RECT 174.200 187.800 174.600 188.200 ;
        RECT 174.200 186.800 174.600 187.200 ;
        RECT 174.200 181.200 174.500 186.800 ;
        RECT 175.000 185.100 175.400 187.900 ;
        RECT 176.600 186.200 176.900 207.800 ;
        RECT 177.400 203.100 177.800 208.900 ;
        RECT 179.800 208.800 180.200 209.200 ;
        RECT 181.400 208.800 181.800 209.200 ;
        RECT 179.800 208.200 180.100 208.800 ;
        RECT 179.800 207.800 180.200 208.200 ;
        RECT 180.600 207.800 181.000 208.200 ;
        RECT 180.600 205.200 180.900 207.800 ;
        RECT 182.200 206.100 182.500 211.800 ;
        RECT 183.800 206.800 184.200 207.200 ;
        RECT 183.000 206.100 183.400 206.200 ;
        RECT 182.200 205.800 183.400 206.100 ;
        RECT 180.600 204.800 181.000 205.200 ;
        RECT 183.800 199.200 184.100 206.800 ;
        RECT 184.600 206.200 184.900 221.800 ;
        RECT 185.400 212.100 185.800 217.900 ;
        RECT 187.800 214.800 188.200 215.200 ;
        RECT 187.800 214.200 188.100 214.800 ;
        RECT 188.600 214.200 188.900 233.800 ;
        RECT 190.200 231.800 190.600 232.200 ;
        RECT 190.200 229.200 190.500 231.800 ;
        RECT 191.000 231.200 191.300 233.800 ;
        RECT 194.200 233.100 194.600 235.900 ;
        RECT 195.800 232.100 196.200 237.900 ;
        RECT 199.000 235.800 199.400 236.200 ;
        RECT 199.000 235.200 199.300 235.800 ;
        RECT 199.000 234.800 199.400 235.200 ;
        RECT 198.200 234.100 198.600 234.200 ;
        RECT 199.000 234.100 199.400 234.200 ;
        RECT 198.200 233.800 199.400 234.100 ;
        RECT 199.000 232.800 199.400 233.200 ;
        RECT 191.000 230.800 191.400 231.200 ;
        RECT 195.800 230.800 196.200 231.200 ;
        RECT 190.200 228.800 190.600 229.200 ;
        RECT 189.400 227.800 189.800 228.200 ;
        RECT 190.200 227.800 190.600 228.200 ;
        RECT 189.400 226.200 189.700 227.800 ;
        RECT 190.200 226.200 190.500 227.800 ;
        RECT 195.800 227.200 196.100 230.800 ;
        RECT 199.000 229.200 199.300 232.800 ;
        RECT 200.600 232.100 201.000 237.900 ;
        RECT 205.400 236.800 205.800 237.200 ;
        RECT 204.600 234.800 205.000 235.200 ;
        RECT 204.600 229.200 204.900 234.800 ;
        RECT 205.400 234.200 205.700 236.800 ;
        RECT 207.000 235.800 207.400 236.200 ;
        RECT 208.600 235.800 209.000 236.200 ;
        RECT 209.400 235.800 209.800 236.200 ;
        RECT 207.000 235.200 207.300 235.800 ;
        RECT 208.600 235.200 208.900 235.800 ;
        RECT 209.400 235.200 209.700 235.800 ;
        RECT 207.000 234.800 207.400 235.200 ;
        RECT 208.600 234.800 209.000 235.200 ;
        RECT 209.400 234.800 209.800 235.200 ;
        RECT 205.400 233.800 205.800 234.200 ;
        RECT 210.200 233.800 210.600 234.200 ;
        RECT 205.400 232.200 205.700 233.800 ;
        RECT 210.200 233.200 210.500 233.800 ;
        RECT 210.200 232.800 210.600 233.200 ;
        RECT 211.000 233.100 211.400 235.900 ;
        RECT 205.400 231.800 205.800 232.200 ;
        RECT 212.600 232.100 213.000 237.900 ;
        RECT 213.400 234.700 213.800 235.100 ;
        RECT 199.000 228.800 199.400 229.200 ;
        RECT 204.600 228.800 205.000 229.200 ;
        RECT 201.400 227.800 201.800 228.200 ;
        RECT 203.800 227.800 204.200 228.200 ;
        RECT 201.400 227.200 201.700 227.800 ;
        RECT 203.800 227.200 204.100 227.800 ;
        RECT 192.600 226.800 193.000 227.200 ;
        RECT 195.000 226.800 195.400 227.200 ;
        RECT 195.800 226.800 196.200 227.200 ;
        RECT 201.400 226.800 201.800 227.200 ;
        RECT 203.800 226.800 204.200 227.200 ;
        RECT 192.600 226.200 192.900 226.800 ;
        RECT 195.000 226.200 195.300 226.800 ;
        RECT 189.400 225.800 189.800 226.200 ;
        RECT 190.200 225.800 190.600 226.200 ;
        RECT 191.000 225.800 191.400 226.200 ;
        RECT 191.800 225.800 192.200 226.200 ;
        RECT 192.600 225.800 193.000 226.200 ;
        RECT 195.000 225.800 195.400 226.200 ;
        RECT 187.800 213.800 188.200 214.200 ;
        RECT 188.600 213.800 189.000 214.200 ;
        RECT 190.200 212.100 190.600 217.900 ;
        RECT 191.000 210.200 191.300 225.800 ;
        RECT 191.800 218.200 192.100 225.800 ;
        RECT 195.800 222.200 196.100 226.800 ;
        RECT 196.600 226.100 197.000 226.200 ;
        RECT 197.400 226.100 197.800 226.200 ;
        RECT 196.600 225.800 197.800 226.100 ;
        RECT 199.800 225.800 200.200 226.200 ;
        RECT 199.800 225.200 200.100 225.800 ;
        RECT 199.800 224.800 200.200 225.200 ;
        RECT 204.600 225.100 205.000 225.200 ;
        RECT 205.400 225.100 205.800 225.200 ;
        RECT 206.200 225.100 206.600 227.900 ;
        RECT 204.600 224.800 205.800 225.100 ;
        RECT 197.400 223.800 197.800 224.200 ;
        RECT 199.800 223.800 200.200 224.200 ;
        RECT 193.400 221.800 193.800 222.200 ;
        RECT 195.800 221.800 196.200 222.200 ;
        RECT 191.800 217.800 192.200 218.200 ;
        RECT 191.800 213.100 192.200 215.900 ;
        RECT 191.000 209.800 191.400 210.200 ;
        RECT 193.400 209.200 193.700 221.800 ;
        RECT 197.400 218.200 197.700 223.800 ;
        RECT 199.000 221.800 199.400 222.200 ;
        RECT 197.400 218.100 197.800 218.200 ;
        RECT 198.200 218.100 198.600 218.200 ;
        RECT 197.400 217.800 198.600 218.100 ;
        RECT 191.000 208.800 191.400 209.200 ;
        RECT 193.400 208.800 193.800 209.200 ;
        RECT 194.200 209.100 194.600 209.200 ;
        RECT 195.000 209.100 195.400 209.200 ;
        RECT 194.200 208.800 195.400 209.100 ;
        RECT 195.800 208.800 196.200 209.200 ;
        RECT 188.600 207.800 189.000 208.200 ;
        RECT 187.000 206.800 187.400 207.200 ;
        RECT 187.000 206.200 187.300 206.800 ;
        RECT 188.600 206.200 188.900 207.800 ;
        RECT 189.400 207.100 189.800 207.200 ;
        RECT 190.200 207.100 190.600 207.200 ;
        RECT 189.400 206.800 190.600 207.100 ;
        RECT 184.600 205.800 185.000 206.200 ;
        RECT 187.000 205.800 187.400 206.200 ;
        RECT 187.800 205.800 188.200 206.200 ;
        RECT 188.600 205.800 189.000 206.200 ;
        RECT 187.800 203.200 188.100 205.800 ;
        RECT 187.800 202.800 188.200 203.200 ;
        RECT 186.200 201.800 186.600 202.200 ;
        RECT 183.800 198.800 184.200 199.200 ;
        RECT 186.200 198.200 186.500 201.800 ;
        RECT 186.200 197.800 186.600 198.200 ;
        RECT 181.400 196.100 181.800 196.200 ;
        RECT 182.200 196.100 182.600 196.200 ;
        RECT 181.400 195.800 182.600 196.100 ;
        RECT 185.400 196.100 185.800 196.200 ;
        RECT 188.600 196.100 189.000 196.200 ;
        RECT 185.400 195.800 189.000 196.100 ;
        RECT 191.000 195.200 191.300 208.800 ;
        RECT 195.800 208.200 196.100 208.800 ;
        RECT 195.000 207.800 195.400 208.200 ;
        RECT 195.800 207.800 196.200 208.200 ;
        RECT 195.000 207.200 195.300 207.800 ;
        RECT 199.000 207.200 199.300 221.800 ;
        RECT 199.800 215.200 200.100 223.800 ;
        RECT 207.800 223.100 208.200 228.900 ;
        RECT 210.200 226.800 210.600 227.200 ;
        RECT 208.600 225.900 209.000 226.300 ;
        RECT 205.400 215.800 205.800 216.200 ;
        RECT 207.800 215.800 208.200 216.200 ;
        RECT 205.400 215.200 205.700 215.800 ;
        RECT 207.800 215.200 208.100 215.800 ;
        RECT 199.800 214.800 200.200 215.200 ;
        RECT 204.600 214.800 205.000 215.200 ;
        RECT 205.400 214.800 205.800 215.200 ;
        RECT 207.800 214.800 208.200 215.200 ;
        RECT 204.600 214.200 204.900 214.800 ;
        RECT 204.600 213.800 205.000 214.200 ;
        RECT 202.200 208.800 202.600 209.200 ;
        RECT 202.200 208.200 202.500 208.800 ;
        RECT 202.200 207.800 202.600 208.200 ;
        RECT 191.800 206.800 192.200 207.200 ;
        RECT 195.000 206.800 195.400 207.200 ;
        RECT 197.400 206.800 197.800 207.200 ;
        RECT 199.000 206.800 199.400 207.200 ;
        RECT 191.800 206.200 192.100 206.800 ;
        RECT 197.400 206.200 197.700 206.800 ;
        RECT 191.800 205.800 192.200 206.200 ;
        RECT 192.600 205.800 193.000 206.200 ;
        RECT 193.400 206.100 193.800 206.200 ;
        RECT 194.200 206.100 194.600 206.200 ;
        RECT 193.400 205.800 194.600 206.100 ;
        RECT 196.600 205.800 197.000 206.200 ;
        RECT 197.400 205.800 197.800 206.200 ;
        RECT 199.000 206.100 199.400 206.200 ;
        RECT 199.800 206.100 200.200 206.200 ;
        RECT 199.000 205.800 200.200 206.100 ;
        RECT 192.600 205.200 192.900 205.800 ;
        RECT 196.600 205.200 196.900 205.800 ;
        RECT 192.600 204.800 193.000 205.200 ;
        RECT 196.600 204.800 197.000 205.200 ;
        RECT 201.400 204.800 201.800 205.200 ;
        RECT 199.800 201.800 200.200 202.200 ;
        RECT 195.000 199.800 195.400 200.200 ;
        RECT 195.000 195.200 195.300 199.800 ;
        RECT 199.800 196.200 200.100 201.800 ;
        RECT 199.800 195.800 200.200 196.200 ;
        RECT 187.800 194.800 188.200 195.200 ;
        RECT 191.000 194.800 191.400 195.200 ;
        RECT 191.800 194.800 192.200 195.200 ;
        RECT 192.600 195.100 193.000 195.200 ;
        RECT 193.400 195.100 193.800 195.200 ;
        RECT 192.600 194.800 193.800 195.100 ;
        RECT 195.000 194.800 195.400 195.200 ;
        RECT 195.800 194.800 196.200 195.200 ;
        RECT 197.400 194.800 197.800 195.200 ;
        RECT 199.800 194.800 200.200 195.200 ;
        RECT 200.600 194.800 201.000 195.200 ;
        RECT 184.600 193.800 185.000 194.200 ;
        RECT 187.000 193.800 187.400 194.200 ;
        RECT 179.000 188.800 179.400 189.200 ;
        RECT 179.000 186.200 179.300 188.800 ;
        RECT 179.800 187.100 180.200 187.200 ;
        RECT 180.600 187.100 181.000 187.200 ;
        RECT 179.800 186.800 181.000 187.100 ;
        RECT 183.000 187.100 183.400 187.200 ;
        RECT 183.800 187.100 184.200 187.200 ;
        RECT 183.000 186.800 184.200 187.100 ;
        RECT 175.800 185.800 176.200 186.200 ;
        RECT 176.600 185.800 177.000 186.200 ;
        RECT 179.000 185.800 179.400 186.200 ;
        RECT 181.400 185.800 181.800 186.200 ;
        RECT 174.200 180.800 174.600 181.200 ;
        RECT 171.800 178.800 172.200 179.200 ;
        RECT 171.800 177.200 172.100 178.800 ;
        RECT 175.800 178.200 176.100 185.800 ;
        RECT 181.400 184.200 181.700 185.800 ;
        RECT 183.800 184.800 184.200 185.200 ;
        RECT 183.800 184.200 184.100 184.800 ;
        RECT 181.400 183.800 181.800 184.200 ;
        RECT 183.800 183.800 184.200 184.200 ;
        RECT 177.400 183.100 177.800 183.200 ;
        RECT 178.200 183.100 178.600 183.200 ;
        RECT 177.400 182.800 178.600 183.100 ;
        RECT 184.600 181.200 184.900 193.800 ;
        RECT 187.000 189.200 187.300 193.800 ;
        RECT 187.800 192.200 188.100 194.800 ;
        RECT 188.600 193.800 189.000 194.200 ;
        RECT 190.200 193.800 190.600 194.200 ;
        RECT 188.600 192.200 188.900 193.800 ;
        RECT 187.800 191.800 188.200 192.200 ;
        RECT 188.600 191.800 189.000 192.200 ;
        RECT 190.200 191.200 190.500 193.800 ;
        RECT 191.800 193.200 192.100 194.800 ;
        RECT 195.800 194.200 196.100 194.800 ;
        RECT 195.800 193.800 196.200 194.200 ;
        RECT 191.800 192.800 192.200 193.200 ;
        RECT 197.400 192.200 197.700 194.800 ;
        RECT 193.400 192.100 193.800 192.200 ;
        RECT 194.200 192.100 194.600 192.200 ;
        RECT 193.400 191.800 194.600 192.100 ;
        RECT 197.400 191.800 197.800 192.200 ;
        RECT 190.200 190.800 190.600 191.200 ;
        RECT 199.800 189.200 200.100 194.800 ;
        RECT 200.600 194.200 200.900 194.800 ;
        RECT 200.600 193.800 201.000 194.200 ;
        RECT 201.400 193.100 201.700 204.800 ;
        RECT 205.400 204.200 205.700 214.800 ;
        RECT 207.800 214.100 208.200 214.200 ;
        RECT 208.600 214.100 208.900 225.900 ;
        RECT 207.800 213.800 208.900 214.100 ;
        RECT 209.400 221.800 209.800 222.200 ;
        RECT 209.400 214.200 209.700 221.800 ;
        RECT 210.200 218.200 210.500 226.800 ;
        RECT 212.600 223.100 213.000 228.900 ;
        RECT 213.400 221.200 213.700 234.700 ;
        RECT 214.200 233.800 214.600 234.200 ;
        RECT 214.200 225.200 214.500 233.800 ;
        RECT 217.400 232.100 217.800 237.900 ;
        RECT 220.600 236.100 221.000 236.200 ;
        RECT 221.400 236.100 221.800 236.200 ;
        RECT 220.600 235.800 221.800 236.100 ;
        RECT 221.400 234.100 221.800 234.200 ;
        RECT 222.200 234.100 222.600 234.200 ;
        RECT 221.400 233.800 222.600 234.100 ;
        RECT 223.000 233.100 223.400 235.900 ;
        RECT 223.800 234.800 224.200 235.200 ;
        RECT 223.800 234.200 224.100 234.800 ;
        RECT 223.800 233.800 224.200 234.200 ;
        RECT 219.800 231.800 220.200 232.200 ;
        RECT 220.600 231.800 221.000 232.200 ;
        RECT 221.400 231.800 221.800 232.200 ;
        RECT 224.600 232.100 225.000 237.900 ;
        RECT 226.200 235.100 226.600 235.200 ;
        RECT 227.000 235.100 227.400 235.200 ;
        RECT 226.200 234.800 227.400 235.100 ;
        RECT 225.400 232.800 225.800 233.200 ;
        RECT 219.000 227.800 219.400 228.200 ;
        RECT 219.000 226.200 219.300 227.800 ;
        RECT 215.000 226.100 215.400 226.200 ;
        RECT 215.800 226.100 216.200 226.200 ;
        RECT 215.000 225.800 216.200 226.100 ;
        RECT 216.600 225.800 217.000 226.200 ;
        RECT 219.000 225.800 219.400 226.200 ;
        RECT 214.200 224.800 214.600 225.200 ;
        RECT 215.800 224.800 216.200 225.200 ;
        RECT 214.200 222.100 214.600 222.200 ;
        RECT 215.000 222.100 215.400 222.200 ;
        RECT 214.200 221.800 215.400 222.100 ;
        RECT 213.400 220.800 213.800 221.200 ;
        RECT 215.800 220.200 216.100 224.800 ;
        RECT 216.600 222.200 216.900 225.800 ;
        RECT 216.600 221.800 217.000 222.200 ;
        RECT 218.200 221.800 218.600 222.200 ;
        RECT 215.800 219.800 216.200 220.200 ;
        RECT 215.800 219.200 216.100 219.800 ;
        RECT 215.800 218.800 216.200 219.200 ;
        RECT 210.200 217.800 210.600 218.200 ;
        RECT 210.200 214.200 210.500 217.800 ;
        RECT 217.400 216.800 217.800 217.200 ;
        RECT 217.400 216.200 217.700 216.800 ;
        RECT 217.400 215.800 217.800 216.200 ;
        RECT 217.400 215.200 217.700 215.800 ;
        RECT 217.400 214.800 217.800 215.200 ;
        RECT 209.400 213.800 209.800 214.200 ;
        RECT 210.200 213.800 210.600 214.200 ;
        RECT 215.800 213.800 216.200 214.200 ;
        RECT 205.400 203.800 205.800 204.200 ;
        RECT 206.200 203.100 206.600 208.900 ;
        RECT 209.400 206.800 209.800 207.200 ;
        RECT 208.600 205.800 209.000 206.200 ;
        RECT 208.600 205.200 208.900 205.800 ;
        RECT 208.600 204.800 209.000 205.200 ;
        RECT 200.600 192.800 201.700 193.100 ;
        RECT 200.600 189.200 200.900 192.800 ;
        RECT 203.000 192.100 203.400 192.200 ;
        RECT 203.800 192.100 204.200 192.200 ;
        RECT 205.400 192.100 205.800 197.900 ;
        RECT 209.400 197.200 209.700 206.800 ;
        RECT 211.000 203.100 211.400 208.900 ;
        RECT 211.800 206.800 212.200 207.200 ;
        RECT 211.800 206.200 212.100 206.800 ;
        RECT 211.800 205.800 212.200 206.200 ;
        RECT 212.600 205.100 213.000 207.900 ;
        RECT 213.400 206.800 213.800 207.200 ;
        RECT 213.400 206.200 213.700 206.800 ;
        RECT 213.400 205.800 213.800 206.200 ;
        RECT 209.400 196.800 209.800 197.200 ;
        RECT 207.800 195.800 208.200 196.200 ;
        RECT 208.600 195.800 209.000 196.200 ;
        RECT 203.000 191.800 204.200 192.100 ;
        RECT 186.200 188.800 186.600 189.200 ;
        RECT 187.000 188.800 187.400 189.200 ;
        RECT 189.400 189.100 189.800 189.200 ;
        RECT 190.200 189.100 190.600 189.200 ;
        RECT 189.400 188.800 190.600 189.100 ;
        RECT 186.200 187.200 186.500 188.800 ;
        RECT 187.000 187.800 187.400 188.200 ;
        RECT 187.000 187.200 187.300 187.800 ;
        RECT 186.200 186.800 186.600 187.200 ;
        RECT 187.000 186.800 187.400 187.200 ;
        RECT 188.600 186.800 189.000 187.200 ;
        RECT 188.600 186.200 188.900 186.800 ;
        RECT 185.400 185.800 185.800 186.200 ;
        RECT 186.200 185.800 186.600 186.200 ;
        RECT 188.600 185.800 189.000 186.200 ;
        RECT 189.400 185.800 189.800 186.200 ;
        RECT 177.400 180.800 177.800 181.200 ;
        RECT 181.400 180.800 181.800 181.200 ;
        RECT 184.600 180.800 185.000 181.200 ;
        RECT 174.200 177.800 174.600 178.200 ;
        RECT 175.800 177.800 176.200 178.200 ;
        RECT 174.200 177.200 174.500 177.800 ;
        RECT 177.400 177.200 177.700 180.800 ;
        RECT 171.800 176.800 172.200 177.200 ;
        RECT 174.200 176.800 174.600 177.200 ;
        RECT 175.800 176.800 176.200 177.200 ;
        RECT 177.400 176.800 177.800 177.200 ;
        RECT 171.800 176.200 172.100 176.800 ;
        RECT 175.800 176.200 176.100 176.800 ;
        RECT 171.800 175.800 172.200 176.200 ;
        RECT 175.800 175.800 176.200 176.200 ;
        RECT 171.800 175.200 172.100 175.800 ;
        RECT 171.800 174.800 172.200 175.200 ;
        RECT 173.400 175.100 173.800 175.200 ;
        RECT 174.200 175.100 174.600 175.200 ;
        RECT 173.400 174.800 174.600 175.100 ;
        RECT 175.000 174.800 175.400 175.200 ;
        RECT 175.000 174.200 175.300 174.800 ;
        RECT 170.200 173.800 170.600 174.200 ;
        RECT 171.000 173.800 171.400 174.200 ;
        RECT 175.000 173.800 175.400 174.200 ;
        RECT 165.400 172.800 165.800 173.200 ;
        RECT 169.400 172.800 169.800 173.200 ;
        RECT 178.200 172.100 178.600 177.900 ;
        RECT 180.600 176.800 181.000 177.200 ;
        RECT 180.600 175.200 180.900 176.800 ;
        RECT 180.600 174.800 181.000 175.200 ;
        RECT 165.400 169.800 165.800 170.200 ;
        RECT 172.600 169.800 173.000 170.200 ;
        RECT 151.800 167.800 152.200 168.200 ;
        RECT 149.400 166.100 149.800 166.200 ;
        RECT 150.200 166.100 150.600 166.200 ;
        RECT 149.400 165.800 150.600 166.100 ;
        RECT 152.600 163.100 153.000 168.900 ;
        RECT 164.600 168.800 165.000 169.200 ;
        RECT 154.200 165.100 154.600 167.900 ;
        RECT 163.800 166.800 164.200 167.200 ;
        RECT 155.800 166.100 156.200 166.200 ;
        RECT 156.600 166.100 157.000 166.200 ;
        RECT 155.800 165.800 157.000 166.100 ;
        RECT 157.400 165.800 157.800 166.200 ;
        RECT 159.800 166.100 160.200 166.200 ;
        RECT 160.600 166.100 161.000 166.200 ;
        RECT 159.800 165.800 161.000 166.100 ;
        RECT 161.400 165.800 161.800 166.200 ;
        RECT 145.400 161.800 145.800 162.200 ;
        RECT 154.200 161.800 154.600 162.200 ;
        RECT 144.600 158.800 145.000 159.200 ;
        RECT 143.000 156.800 143.400 157.200 ;
        RECT 142.200 155.800 142.600 156.200 ;
        RECT 143.000 154.200 143.300 156.800 ;
        RECT 143.800 156.100 144.200 156.200 ;
        RECT 144.600 156.100 145.000 156.200 ;
        RECT 143.800 155.800 145.000 156.100 ;
        RECT 145.400 155.200 145.700 161.800 ;
        RECT 152.600 160.800 153.000 161.200 ;
        RECT 152.600 159.200 152.900 160.800 ;
        RECT 152.600 158.800 153.000 159.200 ;
        RECT 147.800 156.100 148.200 156.200 ;
        RECT 148.600 156.100 149.000 156.200 ;
        RECT 147.800 155.800 149.000 156.100 ;
        RECT 154.200 155.200 154.500 161.800 ;
        RECT 157.400 161.200 157.700 165.800 ;
        RECT 161.400 165.200 161.700 165.800 ;
        RECT 161.400 164.800 161.800 165.200 ;
        RECT 162.200 164.800 162.600 165.200 ;
        RECT 162.200 164.200 162.500 164.800 ;
        RECT 162.200 163.800 162.600 164.200 ;
        RECT 159.800 161.800 160.200 162.200 ;
        RECT 157.400 160.800 157.800 161.200 ;
        RECT 159.800 157.200 160.100 161.800 ;
        RECT 159.800 156.800 160.200 157.200 ;
        RECT 155.800 155.800 156.200 156.200 ;
        RECT 158.200 156.100 158.600 156.200 ;
        RECT 159.000 156.100 159.400 156.200 ;
        RECT 158.200 155.800 159.400 156.100 ;
        RECT 155.800 155.200 156.100 155.800 ;
        RECT 145.400 154.800 145.800 155.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 153.400 154.800 153.800 155.200 ;
        RECT 154.200 154.800 154.600 155.200 ;
        RECT 155.800 154.800 156.200 155.200 ;
        RECT 145.400 154.200 145.700 154.800 ;
        RECT 147.800 154.200 148.100 154.800 ;
        RECT 143.000 153.800 143.400 154.200 ;
        RECT 145.400 153.800 145.800 154.200 ;
        RECT 146.200 154.100 146.600 154.200 ;
        RECT 147.000 154.100 147.400 154.200 ;
        RECT 146.200 153.800 147.400 154.100 ;
        RECT 147.800 153.800 148.200 154.200 ;
        RECT 153.400 153.200 153.700 154.800 ;
        RECT 153.400 152.800 153.800 153.200 ;
        RECT 147.800 151.800 148.200 152.200 ;
        RECT 139.800 150.800 140.200 151.200 ;
        RECT 136.600 148.800 137.000 149.200 ;
        RECT 138.200 148.800 138.600 149.200 ;
        RECT 136.600 148.200 136.900 148.800 ;
        RECT 136.600 147.800 137.000 148.200 ;
        RECT 132.600 145.800 133.000 146.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 133.400 141.800 133.800 142.200 ;
        RECT 127.000 140.800 127.400 141.200 ;
        RECT 123.800 135.800 124.200 136.200 ;
        RECT 123.800 135.200 124.100 135.800 ;
        RECT 123.800 134.800 124.200 135.200 ;
        RECT 125.400 135.100 125.800 135.200 ;
        RECT 126.200 135.100 126.600 135.200 ;
        RECT 125.400 134.800 126.600 135.100 ;
        RECT 127.000 134.200 127.300 140.800 ;
        RECT 133.400 138.200 133.700 141.800 ;
        RECT 126.200 134.100 126.600 134.200 ;
        RECT 127.000 134.100 127.400 134.200 ;
        RECT 126.200 133.800 127.400 134.100 ;
        RECT 124.600 131.800 125.000 132.200 ;
        RECT 127.000 132.100 127.400 132.200 ;
        RECT 127.800 132.100 128.200 132.200 ;
        RECT 130.200 132.100 130.600 137.900 ;
        RECT 133.400 137.800 133.800 138.200 ;
        RECT 133.400 134.800 133.800 135.200 ;
        RECT 127.000 131.800 128.200 132.100 ;
        RECT 131.800 131.800 132.200 132.200 ;
        RECT 124.600 131.200 124.900 131.800 ;
        RECT 124.600 130.800 125.000 131.200 ;
        RECT 131.000 129.800 131.400 130.200 ;
        RECT 128.600 129.100 129.000 129.200 ;
        RECT 129.400 129.100 129.800 129.200 ;
        RECT 123.000 127.800 123.400 128.200 ;
        RECT 115.800 120.800 116.200 121.200 ;
        RECT 121.400 120.800 121.800 121.200 ;
        RECT 115.000 112.800 115.400 113.200 ;
        RECT 111.000 110.800 111.400 111.200 ;
        RECT 114.200 110.800 114.600 111.200 ;
        RECT 107.800 108.800 108.200 109.200 ;
        RECT 108.600 108.800 109.000 109.200 ;
        RECT 111.000 107.200 111.300 110.800 ;
        RECT 105.400 106.800 105.800 107.200 ;
        RECT 106.200 106.800 106.600 107.200 ;
        RECT 110.200 106.800 110.600 107.200 ;
        RECT 111.000 106.800 111.400 107.200 ;
        RECT 105.400 105.800 105.800 106.200 ;
        RECT 105.400 105.200 105.700 105.800 ;
        RECT 105.400 104.800 105.800 105.200 ;
        RECT 106.200 104.200 106.500 106.800 ;
        RECT 110.200 105.200 110.500 106.800 ;
        RECT 107.000 105.100 107.400 105.200 ;
        RECT 107.800 105.100 108.200 105.200 ;
        RECT 107.000 104.800 108.200 105.100 ;
        RECT 110.200 104.800 110.600 105.200 ;
        RECT 111.000 105.100 111.400 105.200 ;
        RECT 111.800 105.100 112.200 105.200 ;
        RECT 111.000 104.800 112.200 105.100 ;
        RECT 112.600 104.800 113.000 105.200 ;
        RECT 106.200 103.800 106.600 104.200 ;
        RECT 107.800 102.200 108.100 104.800 ;
        RECT 107.800 101.800 108.200 102.200 ;
        RECT 109.400 101.800 109.800 102.200 ;
        RECT 105.400 92.100 105.800 97.900 ;
        RECT 106.200 95.000 106.600 95.100 ;
        RECT 107.000 95.000 107.400 95.100 ;
        RECT 106.200 94.700 107.400 95.000 ;
        RECT 106.200 92.800 106.600 93.200 ;
        RECT 107.800 92.800 108.200 93.200 ;
        RECT 102.200 88.800 102.600 89.200 ;
        RECT 103.000 88.800 103.400 89.200 ;
        RECT 104.600 88.800 105.000 89.200 ;
        RECT 103.000 87.200 103.300 88.800 ;
        RECT 96.600 87.100 97.000 87.200 ;
        RECT 95.800 86.800 97.000 87.100 ;
        RECT 100.600 86.800 101.000 87.200 ;
        RECT 103.000 86.800 103.400 87.200 ;
        RECT 95.800 85.800 96.200 86.200 ;
        RECT 95.800 85.200 96.100 85.800 ;
        RECT 95.800 84.800 96.200 85.200 ;
        RECT 96.600 84.800 97.000 85.200 ;
        RECT 101.400 85.100 101.800 85.200 ;
        RECT 102.200 85.100 102.600 85.200 ;
        RECT 101.400 84.800 102.600 85.100 ;
        RECT 96.600 84.200 96.900 84.800 ;
        RECT 96.600 83.800 97.000 84.200 ;
        RECT 95.000 81.800 95.400 82.200 ;
        RECT 97.400 81.800 97.800 82.200 ;
        RECT 101.400 81.800 101.800 82.200 ;
        RECT 95.000 79.800 95.400 80.200 ;
        RECT 95.000 79.200 95.300 79.800 ;
        RECT 95.000 78.800 95.400 79.200 ;
        RECT 94.200 76.800 94.600 77.200 ;
        RECT 94.200 76.200 94.500 76.800 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 92.600 76.100 93.000 76.200 ;
        RECT 93.400 76.100 93.800 76.200 ;
        RECT 92.600 75.800 93.800 76.100 ;
        RECT 94.200 75.800 94.600 76.200 ;
        RECT 91.000 74.800 91.400 75.200 ;
        RECT 88.600 73.800 89.000 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 91.800 74.100 92.200 74.200 ;
        RECT 92.600 74.100 93.000 74.200 ;
        RECT 91.800 73.800 93.000 74.100 ;
        RECT 94.200 73.800 94.600 74.200 ;
        RECT 95.000 74.100 95.400 74.200 ;
        RECT 95.800 74.100 96.200 74.200 ;
        RECT 95.000 73.800 96.200 74.100 ;
        RECT 96.600 73.800 97.000 74.200 ;
        RECT 87.000 72.800 88.100 73.100 ;
        RECT 83.000 70.800 83.400 71.200 ;
        RECT 83.000 67.800 83.400 68.200 ;
        RECT 83.000 67.200 83.300 67.800 ;
        RECT 85.400 67.200 85.700 72.800 ;
        RECT 86.200 72.100 86.600 72.200 ;
        RECT 87.000 72.100 87.400 72.200 ;
        RECT 86.200 71.800 87.400 72.100 ;
        RECT 87.800 68.200 88.100 72.800 ;
        RECT 90.200 72.200 90.500 73.800 ;
        RECT 89.400 71.800 89.800 72.200 ;
        RECT 90.200 71.800 90.600 72.200 ;
        RECT 92.600 71.800 93.000 72.200 ;
        RECT 89.400 70.200 89.700 71.800 ;
        RECT 92.600 70.200 92.900 71.800 ;
        RECT 89.400 69.800 89.800 70.200 ;
        RECT 92.600 69.800 93.000 70.200 ;
        RECT 91.000 68.800 91.400 69.200 ;
        RECT 87.800 67.800 88.200 68.200 ;
        RECT 91.000 67.200 91.300 68.800 ;
        RECT 91.800 67.800 92.200 68.200 ;
        RECT 83.000 66.800 83.400 67.200 ;
        RECT 85.400 66.800 85.800 67.200 ;
        RECT 89.400 67.100 89.800 67.200 ;
        RECT 90.200 67.100 90.600 67.200 ;
        RECT 89.400 66.800 90.600 67.100 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 91.800 66.200 92.100 67.800 ;
        RECT 92.600 67.100 93.000 67.200 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 92.600 66.800 93.800 67.100 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 79.800 65.800 80.200 66.200 ;
        RECT 80.600 65.800 81.000 66.200 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 82.200 66.100 82.600 66.200 ;
        RECT 81.400 65.800 82.600 66.100 ;
        RECT 84.600 65.800 85.000 66.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 88.600 66.100 89.000 66.200 ;
        RECT 90.200 66.100 90.600 66.200 ;
        RECT 91.000 66.100 91.400 66.200 ;
        RECT 88.600 65.800 89.700 66.100 ;
        RECT 90.200 65.800 91.400 66.100 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 79.000 65.200 79.300 65.800 ;
        RECT 79.800 65.200 80.100 65.800 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 79.800 64.800 80.200 65.200 ;
        RECT 78.200 58.800 78.600 59.200 ;
        RECT 80.600 58.200 80.900 65.800 ;
        RECT 84.600 65.200 84.900 65.800 ;
        RECT 86.200 65.200 86.500 65.800 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 86.200 64.800 86.600 65.200 ;
        RECT 87.800 62.800 88.200 63.200 ;
        RECT 87.800 62.200 88.100 62.800 ;
        RECT 87.800 61.800 88.200 62.200 ;
        RECT 87.800 59.800 88.200 60.200 ;
        RECT 84.600 59.100 85.000 59.200 ;
        RECT 85.400 59.100 85.800 59.200 ;
        RECT 84.600 58.800 85.800 59.100 ;
        RECT 72.600 56.800 73.000 57.200 ;
        RECT 71.000 55.000 71.400 55.100 ;
        RECT 71.800 55.000 72.200 55.100 ;
        RECT 71.000 54.700 72.200 55.000 ;
        RECT 75.000 52.100 75.400 57.900 ;
        RECT 80.600 57.800 81.000 58.200 ;
        RECT 77.400 56.800 77.800 57.200 ;
        RECT 81.400 56.800 81.800 57.200 ;
        RECT 77.400 56.200 77.700 56.800 ;
        RECT 77.400 55.800 77.800 56.200 ;
        RECT 81.400 55.200 81.700 56.800 ;
        RECT 87.000 55.800 87.400 56.200 ;
        RECT 87.000 55.200 87.300 55.800 ;
        RECT 87.800 55.200 88.100 59.800 ;
        RECT 89.400 59.200 89.700 65.800 ;
        RECT 94.200 65.200 94.500 73.800 ;
        RECT 96.600 69.200 96.900 73.800 ;
        RECT 95.800 68.800 96.200 69.200 ;
        RECT 96.600 68.800 97.000 69.200 ;
        RECT 95.800 68.200 96.100 68.800 ;
        RECT 95.800 67.800 96.200 68.200 ;
        RECT 93.400 65.100 93.800 65.200 ;
        RECT 94.200 65.100 94.600 65.200 ;
        RECT 93.400 64.800 94.600 65.100 ;
        RECT 94.200 59.200 94.500 64.800 ;
        RECT 96.600 61.800 97.000 62.200 ;
        RECT 89.400 58.800 89.800 59.200 ;
        RECT 94.200 58.800 94.600 59.200 ;
        RECT 96.600 55.200 96.900 61.800 ;
        RECT 79.000 54.800 79.400 55.200 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 80.600 55.100 81.000 55.200 ;
        RECT 79.800 54.800 81.000 55.100 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 83.000 55.100 83.400 55.200 ;
        RECT 83.800 55.100 84.200 55.200 ;
        RECT 83.000 54.800 84.200 55.100 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 87.800 54.800 88.200 55.200 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 91.000 55.100 91.400 55.200 ;
        RECT 91.800 55.100 92.200 55.200 ;
        RECT 91.000 54.800 92.200 55.100 ;
        RECT 92.600 54.800 93.000 55.200 ;
        RECT 93.400 54.800 93.800 55.200 ;
        RECT 95.000 55.100 95.400 55.200 ;
        RECT 95.800 55.100 96.200 55.200 ;
        RECT 95.000 54.800 96.200 55.100 ;
        RECT 96.600 54.800 97.000 55.200 ;
        RECT 79.000 49.200 79.300 54.800 ;
        RECT 67.800 43.100 68.200 48.900 ;
        RECT 69.400 48.800 69.800 49.200 ;
        RECT 70.200 49.100 70.600 49.200 ;
        RECT 71.000 49.100 71.400 49.200 ;
        RECT 70.200 48.800 71.400 49.100 ;
        RECT 75.800 48.800 76.200 49.200 ;
        RECT 71.000 47.800 71.400 48.200 ;
        RECT 71.000 47.200 71.300 47.800 ;
        RECT 75.800 47.200 76.100 48.800 ;
        RECT 71.000 46.800 71.400 47.200 ;
        RECT 72.600 47.100 73.000 47.200 ;
        RECT 73.400 47.100 73.800 47.200 ;
        RECT 72.600 46.800 73.800 47.100 ;
        RECT 75.800 46.800 76.200 47.200 ;
        RECT 71.000 39.200 71.300 46.800 ;
        RECT 71.800 46.100 72.200 46.200 ;
        RECT 72.600 46.100 73.000 46.200 ;
        RECT 71.800 45.800 73.000 46.100 ;
        RECT 74.200 45.800 74.600 46.200 ;
        RECT 74.200 45.200 74.500 45.800 ;
        RECT 74.200 44.800 74.600 45.200 ;
        RECT 76.600 45.100 77.000 47.900 ;
        RECT 77.400 46.800 77.800 47.200 ;
        RECT 77.400 45.200 77.700 46.800 ;
        RECT 77.400 44.800 77.800 45.200 ;
        RECT 58.200 38.800 58.600 39.200 ;
        RECT 67.000 38.800 67.400 39.200 ;
        RECT 71.000 38.800 71.400 39.200 ;
        RECT 72.600 37.800 73.000 38.200 ;
        RECT 55.000 36.800 55.400 37.200 ;
        RECT 55.000 35.200 55.300 36.800 ;
        RECT 55.800 35.800 56.200 36.200 ;
        RECT 55.800 35.200 56.100 35.800 ;
        RECT 72.600 35.200 72.900 37.800 ;
        RECT 55.000 34.800 55.400 35.200 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 56.600 34.800 57.000 35.200 ;
        RECT 61.400 34.800 61.800 35.200 ;
        RECT 63.800 34.800 64.200 35.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 66.200 35.100 66.600 35.200 ;
        RECT 67.000 35.100 67.400 35.200 ;
        RECT 66.200 34.800 67.400 35.100 ;
        RECT 67.800 34.800 68.200 35.200 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 69.400 35.100 69.800 35.200 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 69.400 34.800 70.600 35.100 ;
        RECT 72.600 34.800 73.000 35.200 ;
        RECT 56.600 34.200 56.900 34.800 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 56.600 33.800 57.000 34.200 ;
        RECT 54.200 29.200 54.500 33.800 ;
        RECT 55.000 33.200 55.300 33.800 ;
        RECT 55.000 32.800 55.400 33.200 ;
        RECT 56.600 32.800 57.000 33.200 ;
        RECT 54.200 28.800 54.600 29.200 ;
        RECT 56.600 27.200 56.900 32.800 ;
        RECT 61.400 30.200 61.700 34.800 ;
        RECT 63.800 32.200 64.100 34.800 ;
        RECT 63.800 31.800 64.200 32.200 ;
        RECT 61.400 29.800 61.800 30.200 ;
        RECT 56.600 26.800 57.000 27.200 ;
        RECT 58.200 27.100 58.600 27.200 ;
        RECT 59.000 27.100 59.400 27.200 ;
        RECT 58.200 26.800 59.400 27.100 ;
        RECT 61.400 26.800 61.800 27.200 ;
        RECT 55.000 25.800 55.400 26.200 ;
        RECT 55.000 24.200 55.300 25.800 ;
        RECT 55.000 23.800 55.400 24.200 ;
        RECT 53.400 16.800 53.800 17.200 ;
        RECT 44.600 14.800 45.000 15.200 ;
        RECT 47.800 14.800 48.200 15.200 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 51.000 14.800 51.400 15.200 ;
        RECT 35.800 11.800 36.200 12.200 ;
        RECT 43.000 11.800 43.400 12.200 ;
        RECT 43.000 9.200 43.300 11.800 ;
        RECT 44.600 10.200 44.900 14.800 ;
        RECT 44.600 9.800 45.000 10.200 ;
        RECT 41.400 9.100 41.800 9.200 ;
        RECT 42.200 9.100 42.600 9.200 ;
        RECT 34.200 6.800 34.600 7.200 ;
        RECT 35.000 3.100 35.400 8.900 ;
        RECT 35.800 5.900 36.200 6.300 ;
        RECT 35.800 5.200 36.100 5.900 ;
        RECT 35.800 4.800 36.200 5.200 ;
        RECT 39.800 3.100 40.200 8.900 ;
        RECT 41.400 8.800 42.600 9.100 ;
        RECT 43.000 8.800 43.400 9.200 ;
        RECT 47.800 7.200 48.100 14.800 ;
        RECT 53.400 14.200 53.700 16.800 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 49.400 7.200 49.700 8.800 ;
        RECT 43.000 7.100 43.400 7.200 ;
        RECT 43.800 7.100 44.200 7.200 ;
        RECT 43.000 6.800 44.200 7.100 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 45.400 6.800 46.600 7.100 ;
        RECT 47.800 6.800 48.200 7.200 ;
        RECT 49.400 6.800 49.800 7.200 ;
        RECT 43.000 6.100 43.400 6.200 ;
        RECT 43.800 6.100 44.200 6.200 ;
        RECT 43.000 5.800 44.200 6.100 ;
        RECT 46.200 5.800 46.600 6.200 ;
        RECT 46.200 5.200 46.500 5.800 ;
        RECT 46.200 4.800 46.600 5.200 ;
        RECT 52.600 3.100 53.000 8.900 ;
        RECT 53.400 7.200 53.700 13.800 ;
        RECT 56.600 12.200 56.900 26.800 ;
        RECT 57.400 26.100 57.800 26.200 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 57.400 25.800 58.600 26.100 ;
        RECT 59.800 25.100 60.200 25.200 ;
        RECT 60.600 25.100 61.000 25.200 ;
        RECT 59.800 24.800 61.000 25.100 ;
        RECT 60.600 23.800 61.000 24.200 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 59.800 14.200 60.100 14.800 ;
        RECT 60.600 14.200 60.900 23.800 ;
        RECT 61.400 23.200 61.700 26.800 ;
        RECT 62.200 25.100 62.600 27.900 ;
        RECT 61.400 22.800 61.800 23.200 ;
        RECT 63.800 23.100 64.200 28.900 ;
        RECT 64.600 23.200 64.900 34.800 ;
        RECT 66.200 27.800 66.600 28.200 ;
        RECT 66.200 27.200 66.500 27.800 ;
        RECT 65.400 26.800 65.800 27.200 ;
        RECT 66.200 26.800 66.600 27.200 ;
        RECT 65.400 26.200 65.700 26.800 ;
        RECT 65.400 25.800 65.800 26.200 ;
        RECT 64.600 22.800 65.000 23.200 ;
        RECT 61.400 15.200 61.700 22.800 ;
        RECT 64.600 18.200 64.900 22.800 ;
        RECT 64.600 17.800 65.000 18.200 ;
        RECT 62.200 16.800 62.600 17.200 ;
        RECT 64.600 16.800 65.000 17.200 ;
        RECT 62.200 16.200 62.500 16.800 ;
        RECT 62.200 15.800 62.600 16.200 ;
        RECT 64.600 15.200 64.900 16.800 ;
        RECT 65.400 15.800 65.800 16.200 ;
        RECT 65.400 15.200 65.700 15.800 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 64.600 14.800 65.000 15.200 ;
        RECT 65.400 14.800 65.800 15.200 ;
        RECT 59.800 13.800 60.200 14.200 ;
        RECT 60.600 13.800 61.000 14.200 ;
        RECT 63.800 13.800 64.200 14.200 ;
        RECT 65.400 13.800 65.800 14.200 ;
        RECT 56.600 11.800 57.000 12.200 ;
        RECT 59.800 9.100 60.200 9.200 ;
        RECT 60.600 9.100 60.900 13.800 ;
        RECT 53.400 6.800 53.800 7.200 ;
        RECT 55.800 6.800 56.200 7.200 ;
        RECT 55.800 6.200 56.100 6.800 ;
        RECT 55.800 5.800 56.200 6.200 ;
        RECT 57.400 3.100 57.800 8.900 ;
        RECT 59.800 8.800 60.900 9.100 ;
        RECT 58.200 7.800 58.600 8.200 ;
        RECT 58.200 7.200 58.500 7.800 ;
        RECT 58.200 6.800 58.600 7.200 ;
        RECT 59.000 5.100 59.400 7.900 ;
        RECT 62.200 3.100 62.600 8.900 ;
        RECT 63.800 6.200 64.100 13.800 ;
        RECT 65.400 12.200 65.700 13.800 ;
        RECT 65.400 11.800 65.800 12.200 ;
        RECT 66.200 8.200 66.500 26.800 ;
        RECT 67.800 19.200 68.100 34.800 ;
        RECT 68.600 31.200 68.900 34.800 ;
        RECT 73.400 33.100 73.800 35.900 ;
        RECT 75.000 32.100 75.400 37.900 ;
        RECT 76.600 34.800 77.000 35.200 ;
        RECT 76.600 34.200 76.900 34.800 ;
        RECT 77.400 34.200 77.700 44.800 ;
        RECT 78.200 43.100 78.600 48.900 ;
        RECT 79.000 48.800 79.400 49.200 ;
        RECT 79.800 46.800 80.200 47.200 ;
        RECT 79.800 46.200 80.100 46.800 ;
        RECT 79.800 45.800 80.200 46.200 ;
        RECT 82.200 44.200 82.500 54.800 ;
        RECT 86.200 54.200 86.500 54.800 ;
        RECT 86.200 53.800 86.600 54.200 ;
        RECT 85.400 52.800 85.800 53.200 ;
        RECT 85.400 49.200 85.700 52.800 ;
        RECT 82.200 43.800 82.600 44.200 ;
        RECT 83.000 43.100 83.400 48.900 ;
        RECT 85.400 48.800 85.800 49.200 ;
        RECT 84.600 44.800 85.000 45.200 ;
        RECT 76.600 33.800 77.000 34.200 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 68.600 30.800 69.000 31.200 ;
        RECT 73.400 30.800 73.800 31.200 ;
        RECT 73.400 29.200 73.700 30.800 ;
        RECT 68.600 23.100 69.000 28.900 ;
        RECT 71.000 28.800 71.400 29.200 ;
        RECT 73.400 28.800 73.800 29.200 ;
        RECT 71.000 26.200 71.300 28.800 ;
        RECT 75.800 27.800 76.200 28.200 ;
        RECT 75.800 26.200 76.100 27.800 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 76.600 26.200 76.900 26.800 ;
        RECT 71.000 25.800 71.400 26.200 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 73.400 26.100 73.800 26.200 ;
        RECT 72.600 25.800 73.800 26.100 ;
        RECT 75.000 25.800 75.400 26.200 ;
        RECT 75.800 25.800 76.200 26.200 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 70.200 20.800 70.600 21.200 ;
        RECT 67.800 18.800 68.200 19.200 ;
        RECT 70.200 15.200 70.500 20.800 ;
        RECT 69.400 14.800 69.800 15.200 ;
        RECT 70.200 14.800 70.600 15.200 ;
        RECT 69.400 13.200 69.700 14.800 ;
        RECT 69.400 12.800 69.800 13.200 ;
        RECT 71.000 13.100 71.400 15.900 ;
        RECT 71.800 14.800 72.200 15.200 ;
        RECT 71.800 14.200 72.100 14.800 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 71.000 11.800 71.400 12.200 ;
        RECT 72.600 12.100 73.000 17.900 ;
        RECT 74.200 14.800 74.600 15.200 ;
        RECT 74.200 14.200 74.500 14.800 ;
        RECT 74.200 13.800 74.600 14.200 ;
        RECT 75.000 12.200 75.300 25.800 ;
        RECT 77.400 24.100 77.700 33.800 ;
        RECT 79.800 32.100 80.200 37.900 ;
        RECT 82.200 36.800 82.600 37.200 ;
        RECT 82.200 35.200 82.500 36.800 ;
        RECT 84.600 36.200 84.900 44.800 ;
        RECT 86.200 40.800 86.600 41.200 ;
        RECT 85.400 36.800 85.800 37.200 ;
        RECT 84.600 35.800 85.000 36.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 83.000 34.100 83.400 34.200 ;
        RECT 83.000 33.800 84.100 34.100 ;
        RECT 83.000 32.800 83.400 33.200 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 78.200 27.100 78.600 27.200 ;
        RECT 79.000 27.100 79.400 27.200 ;
        RECT 78.200 26.800 79.400 27.100 ;
        RECT 80.600 26.800 81.000 27.200 ;
        RECT 81.400 26.800 81.800 27.200 ;
        RECT 80.600 26.200 80.900 26.800 ;
        RECT 78.200 25.800 78.600 26.200 ;
        RECT 80.600 25.800 81.000 26.200 ;
        RECT 78.200 25.200 78.500 25.800 ;
        RECT 78.200 24.800 78.600 25.200 ;
        RECT 77.400 23.800 78.500 24.100 ;
        RECT 75.000 11.800 75.400 12.200 ;
        RECT 77.400 12.100 77.800 17.900 ;
        RECT 78.200 17.200 78.500 23.800 ;
        RECT 78.200 16.800 78.600 17.200 ;
        RECT 80.600 16.800 81.000 17.200 ;
        RECT 80.600 16.200 80.900 16.800 ;
        RECT 80.600 15.800 81.000 16.200 ;
        RECT 80.600 14.200 80.900 15.800 ;
        RECT 80.600 13.800 81.000 14.200 ;
        RECT 78.200 12.800 78.600 13.200 ;
        RECT 71.000 9.200 71.300 11.800 ;
        RECT 66.200 7.800 66.600 8.200 ;
        RECT 63.800 5.800 64.200 6.200 ;
        RECT 67.000 3.100 67.400 8.900 ;
        RECT 69.400 8.800 69.800 9.200 ;
        RECT 71.000 8.800 71.400 9.200 ;
        RECT 67.800 6.800 68.200 7.200 ;
        RECT 67.800 6.200 68.100 6.800 ;
        RECT 67.800 5.800 68.200 6.200 ;
        RECT 68.600 5.100 69.000 7.900 ;
        RECT 69.400 6.200 69.700 8.800 ;
        RECT 69.400 5.800 69.800 6.200 ;
        RECT 72.600 5.100 73.000 7.900 ;
        RECT 73.400 7.800 73.800 8.200 ;
        RECT 73.400 7.200 73.700 7.800 ;
        RECT 73.400 6.800 73.800 7.200 ;
        RECT 74.200 3.100 74.600 8.900 ;
        RECT 78.200 8.200 78.500 12.800 ;
        RECT 81.400 9.200 81.700 26.800 ;
        RECT 82.200 16.200 82.500 28.800 ;
        RECT 83.000 26.200 83.300 32.800 ;
        RECT 83.800 29.200 84.100 33.800 ;
        RECT 84.600 33.200 84.900 35.800 ;
        RECT 85.400 35.200 85.700 36.800 ;
        RECT 85.400 34.800 85.800 35.200 ;
        RECT 84.600 32.800 85.000 33.200 ;
        RECT 84.600 31.800 85.000 32.200 ;
        RECT 83.800 28.800 84.200 29.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 83.800 26.200 84.100 26.800 ;
        RECT 83.000 25.800 83.400 26.200 ;
        RECT 83.800 25.800 84.200 26.200 ;
        RECT 84.600 25.200 84.900 31.800 ;
        RECT 85.400 31.100 85.700 34.800 ;
        RECT 86.200 34.200 86.500 40.800 ;
        RECT 87.000 36.200 87.300 54.800 ;
        RECT 88.600 54.200 88.900 54.800 ;
        RECT 92.600 54.200 92.900 54.800 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 92.600 53.800 93.000 54.200 ;
        RECT 92.600 51.200 92.900 53.800 ;
        RECT 93.400 53.200 93.700 54.800 ;
        RECT 93.400 52.800 93.800 53.200 ;
        RECT 92.600 50.800 93.000 51.200 ;
        RECT 91.800 49.100 92.200 49.200 ;
        RECT 92.600 49.100 93.000 49.200 ;
        RECT 91.800 48.800 93.000 49.100 ;
        RECT 87.800 47.100 88.200 47.200 ;
        RECT 88.600 47.100 89.000 47.200 ;
        RECT 87.800 46.800 89.000 47.100 ;
        RECT 91.000 47.100 91.400 47.200 ;
        RECT 91.000 46.800 92.100 47.100 ;
        RECT 87.800 45.800 88.200 46.200 ;
        RECT 90.200 46.100 90.600 46.200 ;
        RECT 91.000 46.100 91.400 46.200 ;
        RECT 90.200 45.800 91.400 46.100 ;
        RECT 87.800 45.200 88.100 45.800 ;
        RECT 87.800 44.800 88.200 45.200 ;
        RECT 90.200 40.800 90.600 41.200 ;
        RECT 87.000 35.800 87.400 36.200 ;
        RECT 90.200 35.200 90.500 40.800 ;
        RECT 91.800 37.200 92.100 46.800 ;
        RECT 91.800 36.800 92.200 37.200 ;
        RECT 92.600 35.200 92.900 48.800 ;
        RECT 93.400 44.800 93.800 45.200 ;
        RECT 93.400 39.200 93.700 44.800 ;
        RECT 94.200 43.100 94.600 48.900 ;
        RECT 95.000 42.800 95.400 43.200 ;
        RECT 93.400 38.800 93.800 39.200 ;
        RECT 95.000 35.200 95.300 42.800 ;
        RECT 97.400 42.200 97.700 81.800 ;
        RECT 98.200 77.800 98.600 78.200 ;
        RECT 98.200 76.200 98.500 77.800 ;
        RECT 98.200 75.800 98.600 76.200 ;
        RECT 98.200 75.200 98.500 75.800 ;
        RECT 98.200 74.800 98.600 75.200 ;
        RECT 100.600 71.800 101.000 72.200 ;
        RECT 99.000 63.100 99.400 68.900 ;
        RECT 100.600 66.200 100.900 71.800 ;
        RECT 100.600 65.800 101.000 66.200 ;
        RECT 101.400 64.200 101.700 81.800 ;
        RECT 102.200 79.200 102.500 84.800 ;
        RECT 102.200 78.800 102.600 79.200 ;
        RECT 102.200 77.800 102.600 78.200 ;
        RECT 102.200 75.200 102.500 77.800 ;
        RECT 103.000 76.200 103.300 86.800 ;
        RECT 104.600 84.800 105.000 85.200 ;
        RECT 105.400 85.100 105.800 87.900 ;
        RECT 104.600 84.200 104.900 84.800 ;
        RECT 104.600 83.800 105.000 84.200 ;
        RECT 103.800 81.800 104.200 82.200 ;
        RECT 103.800 77.200 104.100 81.800 ;
        RECT 103.800 76.800 104.200 77.200 ;
        RECT 103.000 75.800 103.400 76.200 ;
        RECT 104.600 75.800 105.000 76.200 ;
        RECT 104.600 75.200 104.900 75.800 ;
        RECT 102.200 74.800 102.600 75.200 ;
        RECT 103.800 75.100 104.200 75.200 ;
        RECT 103.000 74.800 104.200 75.100 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 103.000 74.200 103.300 74.800 ;
        RECT 106.200 74.200 106.500 92.800 ;
        RECT 107.000 83.100 107.400 88.900 ;
        RECT 107.800 88.200 108.100 92.800 ;
        RECT 107.800 87.800 108.200 88.200 ;
        RECT 107.800 84.800 108.200 85.200 ;
        RECT 107.800 79.200 108.100 84.800 ;
        RECT 107.800 78.800 108.200 79.200 ;
        RECT 109.400 76.200 109.700 101.800 ;
        RECT 111.000 100.200 111.300 104.800 ;
        RECT 112.600 102.200 112.900 104.800 ;
        RECT 112.600 101.800 113.000 102.200 ;
        RECT 114.200 101.200 114.500 110.800 ;
        RECT 115.000 109.200 115.300 112.800 ;
        RECT 115.000 108.800 115.400 109.200 ;
        RECT 115.000 101.800 115.400 102.200 ;
        RECT 114.200 100.800 114.600 101.200 ;
        RECT 111.000 99.800 111.400 100.200 ;
        RECT 113.400 98.800 113.800 99.200 ;
        RECT 110.200 92.100 110.600 97.900 ;
        RECT 111.800 97.100 112.200 97.200 ;
        RECT 112.600 97.100 113.000 97.200 ;
        RECT 111.800 96.800 113.000 97.100 ;
        RECT 113.400 94.200 113.700 98.800 ;
        RECT 115.000 96.200 115.300 101.800 ;
        RECT 115.000 95.800 115.400 96.200 ;
        RECT 115.000 94.200 115.300 95.800 ;
        RECT 115.800 95.200 116.100 120.800 ;
        RECT 117.400 112.100 117.800 117.900 ;
        RECT 118.200 114.800 118.600 115.200 ;
        RECT 118.200 114.200 118.500 114.800 ;
        RECT 118.200 113.800 118.600 114.200 ;
        RECT 119.000 113.100 119.400 115.900 ;
        RECT 120.600 112.800 121.000 113.200 ;
        RECT 119.800 111.800 120.200 112.200 ;
        RECT 119.800 111.200 120.100 111.800 ;
        RECT 119.800 110.800 120.200 111.200 ;
        RECT 119.000 109.800 119.400 110.200 ;
        RECT 119.000 109.200 119.300 109.800 ;
        RECT 119.000 108.800 119.400 109.200 ;
        RECT 116.600 99.800 117.000 100.200 ;
        RECT 116.600 99.200 116.900 99.800 ;
        RECT 116.600 98.800 117.000 99.200 ;
        RECT 119.000 96.800 119.400 97.200 ;
        RECT 117.400 95.800 117.800 96.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 112.600 93.800 113.000 94.200 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 115.000 93.800 115.400 94.200 ;
        RECT 110.200 85.800 110.600 86.200 ;
        RECT 110.200 85.200 110.500 85.800 ;
        RECT 110.200 84.800 110.600 85.200 ;
        RECT 111.800 83.100 112.200 88.900 ;
        RECT 110.200 76.800 110.600 77.200 ;
        RECT 108.600 75.800 109.000 76.200 ;
        RECT 109.400 75.800 109.800 76.200 ;
        RECT 108.600 74.200 108.900 75.800 ;
        RECT 109.400 74.800 109.800 75.200 ;
        RECT 103.000 73.800 103.400 74.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 104.600 73.800 105.000 74.200 ;
        RECT 106.200 73.800 106.600 74.200 ;
        RECT 107.000 74.100 107.400 74.200 ;
        RECT 107.800 74.100 108.200 74.200 ;
        RECT 107.000 73.800 108.200 74.100 ;
        RECT 108.600 73.800 109.000 74.200 ;
        RECT 102.200 71.800 102.600 72.200 ;
        RECT 101.400 63.800 101.800 64.200 ;
        RECT 99.000 57.100 99.400 57.200 ;
        RECT 99.800 57.100 100.200 57.200 ;
        RECT 99.000 56.800 100.200 57.100 ;
        RECT 101.400 52.100 101.800 57.900 ;
        RECT 98.200 46.800 98.600 47.200 ;
        RECT 98.200 46.300 98.500 46.800 ;
        RECT 98.200 45.900 98.600 46.300 ;
        RECT 99.000 43.100 99.400 48.900 ;
        RECT 101.400 48.800 101.800 49.200 ;
        RECT 99.800 47.800 100.200 48.200 ;
        RECT 99.800 47.200 100.100 47.800 ;
        RECT 99.800 46.800 100.200 47.200 ;
        RECT 100.600 45.100 101.000 47.900 ;
        RECT 101.400 47.200 101.700 48.800 ;
        RECT 101.400 46.800 101.800 47.200 ;
        RECT 97.400 41.800 97.800 42.200 ;
        RECT 96.600 36.800 97.000 37.200 ;
        RECT 88.600 34.800 89.000 35.200 ;
        RECT 90.200 34.800 90.600 35.200 ;
        RECT 91.800 34.800 92.200 35.200 ;
        RECT 92.600 34.800 93.000 35.200 ;
        RECT 93.400 35.100 93.800 35.200 ;
        RECT 94.200 35.100 94.600 35.200 ;
        RECT 93.400 34.800 94.600 35.100 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 87.000 33.800 87.400 34.200 ;
        RECT 87.000 33.200 87.300 33.800 ;
        RECT 88.600 33.200 88.900 34.800 ;
        RECT 91.800 33.200 92.100 34.800 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 88.600 33.100 89.000 33.200 ;
        RECT 89.400 33.100 89.800 33.200 ;
        RECT 88.600 32.800 89.800 33.100 ;
        RECT 91.800 32.800 92.200 33.200 ;
        RECT 85.400 30.800 86.500 31.100 ;
        RECT 85.400 29.800 85.800 30.200 ;
        RECT 85.400 29.200 85.700 29.800 ;
        RECT 85.400 28.800 85.800 29.200 ;
        RECT 84.600 24.800 85.000 25.200 ;
        RECT 82.200 15.800 82.600 16.200 ;
        RECT 82.200 15.200 82.500 15.800 ;
        RECT 82.200 14.800 82.600 15.200 ;
        RECT 83.800 15.100 84.200 15.200 ;
        RECT 84.600 15.100 85.000 15.200 ;
        RECT 83.800 14.800 85.000 15.100 ;
        RECT 86.200 14.200 86.500 30.800 ;
        RECT 87.800 23.100 88.200 28.900 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 90.200 26.100 90.600 26.200 ;
        RECT 89.400 25.800 90.600 26.100 ;
        RECT 92.600 23.100 93.000 28.900 ;
        RECT 94.200 25.100 94.600 27.900 ;
        RECT 95.000 21.200 95.300 34.800 ;
        RECT 96.600 34.200 96.900 36.800 ;
        RECT 97.400 35.200 97.700 41.800 ;
        RECT 102.200 39.200 102.500 71.800 ;
        RECT 103.000 53.200 103.300 73.800 ;
        RECT 103.800 73.200 104.100 73.800 ;
        RECT 103.800 72.800 104.200 73.200 ;
        RECT 103.800 63.100 104.200 68.900 ;
        RECT 104.600 68.200 104.900 73.800 ;
        RECT 106.200 71.800 106.600 72.200 ;
        RECT 108.600 71.800 109.000 72.200 ;
        RECT 106.200 70.200 106.500 71.800 ;
        RECT 106.200 69.800 106.600 70.200 ;
        RECT 104.600 67.800 105.000 68.200 ;
        RECT 106.200 68.100 106.600 68.200 ;
        RECT 107.000 68.100 107.400 68.200 ;
        RECT 104.600 67.200 104.900 67.800 ;
        RECT 104.600 66.800 105.000 67.200 ;
        RECT 105.400 65.100 105.800 67.900 ;
        RECT 106.200 67.800 107.400 68.100 ;
        RECT 107.800 66.800 108.200 67.200 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 107.000 65.200 107.300 65.800 ;
        RECT 107.800 65.200 108.100 66.800 ;
        RECT 107.000 64.800 107.400 65.200 ;
        RECT 107.800 64.800 108.200 65.200 ;
        RECT 108.600 58.200 108.900 71.800 ;
        RECT 109.400 69.200 109.700 74.800 ;
        RECT 109.400 68.800 109.800 69.200 ;
        RECT 109.400 66.800 109.800 67.200 ;
        RECT 109.400 66.200 109.700 66.800 ;
        RECT 109.400 65.800 109.800 66.200 ;
        RECT 109.400 65.200 109.700 65.800 ;
        RECT 109.400 64.800 109.800 65.200 ;
        RECT 105.400 55.800 105.800 56.200 ;
        RECT 105.400 55.100 105.700 55.800 ;
        RECT 105.400 54.700 105.800 55.100 ;
        RECT 103.000 52.800 103.400 53.200 ;
        RECT 106.200 52.100 106.600 57.900 ;
        RECT 108.600 57.800 109.000 58.200 ;
        RECT 110.200 57.200 110.500 76.800 ;
        RECT 112.600 76.200 112.900 93.800 ;
        RECT 113.400 80.200 113.700 93.800 ;
        RECT 114.200 88.800 114.600 89.200 ;
        RECT 114.200 87.200 114.500 88.800 ;
        RECT 115.000 87.800 115.400 88.200 ;
        RECT 115.000 87.200 115.300 87.800 ;
        RECT 114.200 86.800 114.600 87.200 ;
        RECT 115.000 86.800 115.400 87.200 ;
        RECT 115.800 86.200 116.100 94.800 ;
        RECT 117.400 93.200 117.700 95.800 ;
        RECT 119.000 95.200 119.300 96.800 ;
        RECT 119.800 95.200 120.100 110.800 ;
        RECT 120.600 107.200 120.900 112.800 ;
        RECT 122.200 112.100 122.600 117.900 ;
        RECT 123.000 115.200 123.300 127.800 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 123.800 126.200 124.100 126.800 ;
        RECT 123.800 125.800 124.200 126.200 ;
        RECT 127.000 123.100 127.400 128.900 ;
        RECT 128.600 128.800 129.800 129.100 ;
        RECT 130.200 121.800 130.600 122.200 ;
        RECT 123.000 114.800 123.400 115.200 ;
        RECT 125.400 114.800 125.800 115.200 ;
        RECT 123.000 113.800 123.400 114.200 ;
        RECT 122.200 110.800 122.600 111.200 ;
        RECT 122.200 107.200 122.500 110.800 ;
        RECT 123.000 110.200 123.300 113.800 ;
        RECT 123.000 109.800 123.400 110.200 ;
        RECT 125.400 109.200 125.700 114.800 ;
        RECT 127.000 112.100 127.400 117.900 ;
        RECT 130.200 116.200 130.500 121.800 ;
        RECT 128.600 113.100 129.000 115.900 ;
        RECT 130.200 115.800 130.600 116.200 ;
        RECT 129.400 113.800 129.800 114.200 ;
        RECT 129.400 112.200 129.700 113.800 ;
        RECT 129.400 111.800 129.800 112.200 ;
        RECT 128.600 109.800 129.000 110.200 ;
        RECT 125.400 108.800 125.800 109.200 ;
        RECT 128.600 107.200 128.900 109.800 ;
        RECT 131.000 109.200 131.300 129.800 ;
        RECT 131.000 108.800 131.400 109.200 ;
        RECT 120.600 106.800 121.000 107.200 ;
        RECT 122.200 106.800 122.600 107.200 ;
        RECT 127.800 106.800 128.200 107.200 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 127.000 105.800 127.400 106.200 ;
        RECT 127.000 105.200 127.300 105.800 ;
        RECT 123.000 104.800 123.400 105.200 ;
        RECT 123.800 105.100 124.200 105.200 ;
        RECT 124.600 105.100 125.000 105.200 ;
        RECT 123.800 104.800 125.000 105.100 ;
        RECT 127.000 104.800 127.400 105.200 ;
        RECT 121.400 101.800 121.800 102.200 ;
        RECT 122.200 101.800 122.600 102.200 ;
        RECT 121.400 99.200 121.700 101.800 ;
        RECT 121.400 98.800 121.800 99.200 ;
        RECT 122.200 95.200 122.500 101.800 ;
        RECT 119.000 94.800 119.400 95.200 ;
        RECT 119.800 94.800 120.200 95.200 ;
        RECT 120.600 95.100 121.000 95.200 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 120.600 94.800 121.800 95.100 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 117.400 92.800 117.800 93.200 ;
        RECT 116.600 91.800 117.000 92.200 ;
        RECT 116.600 89.200 116.900 91.800 ;
        RECT 117.400 90.200 117.700 92.800 ;
        RECT 122.200 92.200 122.500 94.800 ;
        RECT 123.000 94.100 123.300 104.800 ;
        RECT 127.000 98.200 127.300 104.800 ;
        RECT 127.000 97.800 127.400 98.200 ;
        RECT 127.800 97.100 128.100 106.800 ;
        RECT 131.800 105.200 132.100 131.800 ;
        RECT 133.400 131.200 133.700 134.800 ;
        RECT 134.200 132.800 134.600 133.200 ;
        RECT 133.400 130.800 133.800 131.200 ;
        RECT 132.600 123.100 133.000 128.900 ;
        RECT 134.200 127.200 134.500 132.800 ;
        RECT 135.000 132.100 135.400 137.900 ;
        RECT 135.800 136.200 136.100 145.800 ;
        RECT 139.000 143.100 139.400 148.900 ;
        RECT 143.000 146.800 143.400 147.200 ;
        RECT 143.000 146.300 143.300 146.800 ;
        RECT 139.800 145.800 140.200 146.200 ;
        RECT 143.000 145.900 143.400 146.300 ;
        RECT 135.800 135.800 136.200 136.200 ;
        RECT 136.600 133.100 137.000 135.900 ;
        RECT 137.400 133.100 137.800 135.900 ;
        RECT 138.200 133.800 138.600 134.200 ;
        RECT 138.200 131.200 138.500 133.800 ;
        RECT 139.000 132.100 139.400 137.900 ;
        RECT 135.000 130.800 135.400 131.200 ;
        RECT 138.200 130.800 138.600 131.200 ;
        RECT 134.200 126.800 134.600 127.200 ;
        RECT 135.000 119.200 135.300 130.800 ;
        RECT 139.800 129.200 140.100 145.800 ;
        RECT 143.800 143.100 144.200 148.900 ;
        RECT 145.400 145.100 145.800 147.900 ;
        RECT 146.200 146.800 146.600 147.200 ;
        RECT 143.000 141.800 143.400 142.200 ;
        RECT 142.200 134.800 142.600 135.200 ;
        RECT 136.600 126.800 137.000 127.200 ;
        RECT 136.600 126.300 136.900 126.800 ;
        RECT 136.600 125.900 137.000 126.300 ;
        RECT 136.600 125.800 136.900 125.900 ;
        RECT 137.400 123.100 137.800 128.900 ;
        RECT 138.200 128.800 138.600 129.200 ;
        RECT 139.800 128.800 140.200 129.200 ;
        RECT 138.200 127.200 138.500 128.800 ;
        RECT 142.200 128.200 142.500 134.800 ;
        RECT 138.200 126.800 138.600 127.200 ;
        RECT 139.000 125.100 139.400 127.900 ;
        RECT 142.200 127.800 142.600 128.200 ;
        RECT 139.800 126.800 140.200 127.200 ;
        RECT 141.400 127.100 141.800 127.200 ;
        RECT 142.200 127.100 142.600 127.200 ;
        RECT 141.400 126.800 142.600 127.100 ;
        RECT 139.000 120.800 139.400 121.200 ;
        RECT 135.000 118.800 135.400 119.200 ;
        RECT 137.400 115.800 137.800 116.200 ;
        RECT 137.400 115.200 137.700 115.800 ;
        RECT 136.600 114.800 137.000 115.200 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 136.600 114.200 136.900 114.800 ;
        RECT 136.600 113.800 137.000 114.200 ;
        RECT 134.200 112.800 134.600 113.200 ;
        RECT 133.400 109.800 133.800 110.200 ;
        RECT 133.400 107.200 133.700 109.800 ;
        RECT 134.200 109.200 134.500 112.800 ;
        RECT 135.800 110.800 136.200 111.200 ;
        RECT 135.000 109.800 135.400 110.200 ;
        RECT 134.200 108.800 134.600 109.200 ;
        RECT 133.400 106.800 133.800 107.200 ;
        RECT 134.200 106.800 134.600 107.200 ;
        RECT 130.200 104.800 130.600 105.200 ;
        RECT 131.000 105.100 131.400 105.200 ;
        RECT 131.800 105.100 132.200 105.200 ;
        RECT 131.000 104.800 132.200 105.100 ;
        RECT 127.000 96.800 128.100 97.100 ;
        RECT 129.400 102.800 129.800 103.200 ;
        RECT 129.400 102.200 129.700 102.800 ;
        RECT 129.400 101.800 129.800 102.200 ;
        RECT 123.800 94.300 124.200 94.400 ;
        RECT 124.600 94.300 125.000 94.400 ;
        RECT 123.800 94.100 125.000 94.300 ;
        RECT 123.000 94.000 125.000 94.100 ;
        RECT 123.000 93.800 124.100 94.000 ;
        RECT 120.600 91.800 121.000 92.200 ;
        RECT 122.200 91.800 122.600 92.200 ;
        RECT 123.000 91.800 123.400 92.200 ;
        RECT 120.600 90.200 120.900 91.800 ;
        RECT 117.400 89.800 117.800 90.200 ;
        RECT 120.600 89.800 121.000 90.200 ;
        RECT 123.000 89.200 123.300 91.800 ;
        RECT 116.600 88.800 117.000 89.200 ;
        RECT 123.000 88.800 123.400 89.200 ;
        RECT 119.800 86.800 120.200 87.200 ;
        RECT 120.600 86.800 121.000 87.200 ;
        RECT 115.800 85.800 116.200 86.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 118.200 85.800 118.600 86.200 ;
        RECT 116.600 85.200 116.900 85.800 ;
        RECT 118.200 85.200 118.500 85.800 ;
        RECT 119.800 85.200 120.100 86.800 ;
        RECT 120.600 86.200 120.900 86.800 ;
        RECT 120.600 85.800 121.000 86.200 ;
        RECT 121.400 85.800 121.800 86.200 ;
        RECT 121.400 85.200 121.700 85.800 ;
        RECT 116.600 84.800 117.000 85.200 ;
        RECT 118.200 84.800 118.600 85.200 ;
        RECT 119.800 84.800 120.200 85.200 ;
        RECT 121.400 84.800 121.800 85.200 ;
        RECT 120.600 82.800 121.000 83.200 ;
        RECT 118.200 80.800 118.600 81.200 ;
        RECT 113.400 79.800 113.800 80.200 ;
        RECT 112.600 75.800 113.000 76.200 ;
        RECT 117.400 75.800 117.800 76.200 ;
        RECT 117.400 75.200 117.700 75.800 ;
        RECT 118.200 75.200 118.500 80.800 ;
        RECT 120.600 76.200 120.900 82.800 ;
        RECT 122.200 81.800 122.600 82.200 ;
        RECT 120.600 75.800 121.000 76.200 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 115.000 75.100 115.400 75.200 ;
        RECT 115.800 75.100 116.200 75.200 ;
        RECT 115.000 74.800 116.200 75.100 ;
        RECT 117.400 74.800 117.800 75.200 ;
        RECT 118.200 74.800 118.600 75.200 ;
        RECT 111.000 69.200 111.300 74.800 ;
        RECT 117.400 73.800 117.800 74.200 ;
        RECT 111.800 72.800 112.200 73.200 ;
        RECT 113.400 72.800 113.800 73.200 ;
        RECT 115.000 72.800 115.400 73.200 ;
        RECT 111.800 72.200 112.100 72.800 ;
        RECT 113.400 72.200 113.700 72.800 ;
        RECT 111.800 71.800 112.200 72.200 ;
        RECT 113.400 71.800 113.800 72.200 ;
        RECT 111.000 68.800 111.400 69.200 ;
        RECT 111.800 66.100 112.200 66.200 ;
        RECT 112.600 66.100 113.000 66.200 ;
        RECT 111.800 65.800 113.000 66.100 ;
        RECT 113.400 66.100 113.700 71.800 ;
        RECT 114.200 67.800 114.600 68.200 ;
        RECT 114.200 67.200 114.500 67.800 ;
        RECT 114.200 66.800 114.600 67.200 ;
        RECT 115.000 66.200 115.300 72.800 ;
        RECT 115.800 71.800 116.200 72.200 ;
        RECT 115.800 71.200 116.100 71.800 ;
        RECT 115.800 70.800 116.200 71.200 ;
        RECT 115.800 68.100 116.200 68.200 ;
        RECT 116.600 68.100 117.000 68.200 ;
        RECT 115.800 67.800 117.000 68.100 ;
        RECT 117.400 67.200 117.700 73.800 ;
        RECT 118.200 69.200 118.500 74.800 ;
        RECT 119.000 74.100 119.400 74.200 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 119.000 73.800 120.200 74.100 ;
        RECT 118.200 68.800 118.600 69.200 ;
        RECT 119.000 69.100 119.400 69.200 ;
        RECT 119.800 69.100 120.200 69.200 ;
        RECT 119.000 68.800 120.200 69.100 ;
        RECT 115.800 66.800 116.200 67.200 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 113.400 65.800 114.500 66.100 ;
        RECT 115.000 65.800 115.400 66.200 ;
        RECT 111.800 64.800 112.200 65.200 ;
        RECT 112.600 65.100 113.000 65.200 ;
        RECT 113.400 65.100 113.800 65.200 ;
        RECT 112.600 64.800 113.800 65.100 ;
        RECT 108.600 56.800 109.000 57.200 ;
        RECT 110.200 56.800 110.600 57.200 ;
        RECT 107.000 53.800 107.400 54.200 ;
        RECT 107.000 47.200 107.300 53.800 ;
        RECT 107.800 53.100 108.200 55.900 ;
        RECT 108.600 54.200 108.900 56.800 ;
        RECT 110.200 56.200 110.500 56.800 ;
        RECT 111.800 56.200 112.100 64.800 ;
        RECT 112.600 56.800 113.000 57.200 ;
        RECT 110.200 55.800 110.600 56.200 ;
        RECT 111.800 55.800 112.200 56.200 ;
        RECT 112.600 55.200 112.900 56.800 ;
        RECT 110.200 54.800 110.600 55.200 ;
        RECT 112.600 54.800 113.000 55.200 ;
        RECT 110.200 54.200 110.500 54.800 ;
        RECT 108.600 53.800 109.000 54.200 ;
        RECT 110.200 53.800 110.600 54.200 ;
        RECT 113.400 53.800 113.800 54.200 ;
        RECT 109.400 52.800 109.800 53.200 ;
        RECT 107.800 50.800 108.200 51.200 ;
        RECT 107.800 47.200 108.100 50.800 ;
        RECT 109.400 49.200 109.700 52.800 ;
        RECT 113.400 51.200 113.700 53.800 ;
        RECT 114.200 53.200 114.500 65.800 ;
        RECT 115.800 64.200 116.100 66.800 ;
        RECT 118.200 65.800 118.600 66.200 ;
        RECT 118.200 65.200 118.500 65.800 ;
        RECT 118.200 64.800 118.600 65.200 ;
        RECT 115.800 63.800 116.200 64.200 ;
        RECT 120.600 61.200 120.900 75.800 ;
        RECT 122.200 75.200 122.500 81.800 ;
        RECT 123.800 76.100 124.100 93.800 ;
        RECT 125.400 93.800 125.800 94.200 ;
        RECT 125.400 93.200 125.700 93.800 ;
        RECT 125.400 92.800 125.800 93.200 ;
        RECT 126.200 91.800 126.600 92.200 ;
        RECT 125.400 87.800 125.800 88.200 ;
        RECT 125.400 87.200 125.700 87.800 ;
        RECT 124.600 86.800 125.000 87.200 ;
        RECT 125.400 86.800 125.800 87.200 ;
        RECT 124.600 86.200 124.900 86.800 ;
        RECT 126.200 86.200 126.500 91.800 ;
        RECT 127.000 88.200 127.300 96.800 ;
        RECT 127.800 89.800 128.200 90.200 ;
        RECT 127.000 87.800 127.400 88.200 ;
        RECT 124.600 85.800 125.000 86.200 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 125.400 85.800 126.600 86.100 ;
        RECT 127.000 85.800 127.400 86.200 ;
        RECT 127.000 85.200 127.300 85.800 ;
        RECT 127.000 84.800 127.400 85.200 ;
        RECT 123.000 75.800 124.100 76.100 ;
        RECT 127.800 76.200 128.100 89.800 ;
        RECT 129.400 88.200 129.700 101.800 ;
        RECT 130.200 101.200 130.500 104.800 ;
        RECT 132.600 103.800 133.000 104.200 ;
        RECT 131.800 101.800 132.200 102.200 ;
        RECT 130.200 100.800 130.600 101.200 ;
        RECT 131.800 93.200 132.100 101.800 ;
        RECT 131.800 92.800 132.200 93.200 ;
        RECT 131.800 91.800 132.200 92.200 ;
        RECT 131.000 88.800 131.400 89.200 ;
        RECT 129.400 87.800 129.800 88.200 ;
        RECT 131.000 87.200 131.300 88.800 ;
        RECT 129.400 87.100 129.800 87.200 ;
        RECT 130.200 87.100 130.600 87.200 ;
        RECT 129.400 86.800 130.600 87.100 ;
        RECT 131.000 86.800 131.400 87.200 ;
        RECT 131.800 86.200 132.100 91.800 ;
        RECT 132.600 91.200 132.900 103.800 ;
        RECT 133.400 94.200 133.700 106.800 ;
        RECT 134.200 99.200 134.500 106.800 ;
        RECT 135.000 105.200 135.300 109.800 ;
        RECT 135.800 109.200 136.100 110.800 ;
        RECT 139.000 110.100 139.300 120.800 ;
        RECT 139.800 116.200 140.100 126.800 ;
        RECT 141.400 124.800 141.800 125.200 ;
        RECT 141.400 122.200 141.700 124.800 ;
        RECT 141.400 121.800 141.800 122.200 ;
        RECT 143.000 116.200 143.300 141.800 ;
        RECT 146.200 141.200 146.500 146.800 ;
        RECT 147.000 145.800 147.400 146.200 ;
        RECT 147.000 145.200 147.300 145.800 ;
        RECT 147.800 145.200 148.100 151.800 ;
        RECT 152.600 149.100 153.000 149.200 ;
        RECT 153.400 149.100 153.800 149.200 ;
        RECT 152.600 148.800 153.800 149.100 ;
        RECT 149.400 147.800 149.800 148.200 ;
        RECT 149.400 147.200 149.700 147.800 ;
        RECT 148.600 146.800 149.000 147.200 ;
        RECT 149.400 146.800 149.800 147.200 ;
        RECT 148.600 146.200 148.900 146.800 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 151.000 145.800 151.400 146.200 ;
        RECT 151.000 145.200 151.300 145.800 ;
        RECT 147.000 144.800 147.400 145.200 ;
        RECT 147.800 144.800 148.200 145.200 ;
        RECT 151.000 144.800 151.400 145.200 ;
        RECT 152.600 145.100 153.000 145.200 ;
        RECT 153.400 145.100 153.800 145.200 ;
        RECT 152.600 144.800 153.800 145.100 ;
        RECT 146.200 140.800 146.600 141.200 ;
        RECT 154.200 141.100 154.500 154.800 ;
        RECT 159.800 154.200 160.100 156.800 ;
        RECT 160.600 155.800 161.000 156.200 ;
        RECT 155.000 153.800 155.400 154.200 ;
        RECT 157.400 154.100 157.800 154.200 ;
        RECT 158.200 154.100 158.600 154.200 ;
        RECT 157.400 153.800 158.600 154.100 ;
        RECT 159.800 153.800 160.200 154.200 ;
        RECT 155.000 148.100 155.300 153.800 ;
        RECT 155.800 148.100 156.200 148.200 ;
        RECT 155.000 147.800 156.200 148.100 ;
        RECT 155.800 147.200 156.100 147.800 ;
        RECT 155.800 146.800 156.200 147.200 ;
        RECT 156.600 146.800 157.000 147.200 ;
        RECT 159.000 147.100 159.400 147.200 ;
        RECT 159.800 147.100 160.200 147.200 ;
        RECT 159.000 146.800 160.200 147.100 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 155.800 145.800 156.200 146.200 ;
        RECT 155.000 142.200 155.300 145.800 ;
        RECT 155.800 145.200 156.100 145.800 ;
        RECT 155.800 144.800 156.200 145.200 ;
        RECT 155.000 141.800 155.400 142.200 ;
        RECT 154.200 140.800 155.300 141.100 ;
        RECT 155.000 138.200 155.300 140.800 ;
        RECT 155.800 139.200 156.100 144.800 ;
        RECT 155.800 138.800 156.200 139.200 ;
        RECT 143.800 132.100 144.200 137.900 ;
        RECT 155.000 137.800 155.400 138.200 ;
        RECT 147.000 136.800 147.400 137.200 ;
        RECT 146.200 135.800 146.600 136.200 ;
        RECT 145.400 129.800 145.800 130.200 ;
        RECT 145.400 127.200 145.700 129.800 ;
        RECT 143.800 126.800 144.200 127.200 ;
        RECT 145.400 126.800 145.800 127.200 ;
        RECT 143.800 126.200 144.100 126.800 ;
        RECT 146.200 126.200 146.500 135.800 ;
        RECT 147.000 134.200 147.300 136.800 ;
        RECT 147.800 136.100 148.200 136.200 ;
        RECT 148.600 136.100 149.000 136.200 ;
        RECT 147.800 135.800 149.000 136.100 ;
        RECT 155.000 135.200 155.300 137.800 ;
        RECT 148.600 134.800 149.000 135.200 ;
        RECT 150.200 134.800 150.600 135.200 ;
        RECT 153.400 135.100 153.800 135.200 ;
        RECT 154.200 135.100 154.600 135.200 ;
        RECT 153.400 134.800 154.600 135.100 ;
        RECT 155.000 134.800 155.400 135.200 ;
        RECT 148.600 134.200 148.900 134.800 ;
        RECT 147.000 134.100 147.400 134.200 ;
        RECT 147.800 134.100 148.200 134.200 ;
        RECT 147.000 133.800 148.200 134.100 ;
        RECT 148.600 133.800 149.000 134.200 ;
        RECT 147.800 131.800 148.200 132.200 ;
        RECT 147.000 127.800 147.400 128.200 ;
        RECT 147.000 127.200 147.300 127.800 ;
        RECT 147.000 126.800 147.400 127.200 ;
        RECT 143.800 125.800 144.200 126.200 ;
        RECT 146.200 125.800 146.600 126.200 ;
        RECT 143.800 122.200 144.100 125.800 ;
        RECT 143.800 121.800 144.200 122.200 ;
        RECT 146.200 117.200 146.500 125.800 ;
        RECT 147.800 125.200 148.100 131.800 ;
        RECT 150.200 129.200 150.500 134.800 ;
        RECT 155.000 134.200 155.300 134.800 ;
        RECT 155.000 133.800 155.400 134.200 ;
        RECT 155.800 133.100 156.200 135.900 ;
        RECT 156.600 135.200 156.900 146.800 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 159.800 145.100 160.200 145.200 ;
        RECT 159.000 144.800 160.200 145.100 ;
        RECT 158.200 141.800 158.600 142.200 ;
        RECT 156.600 134.800 157.000 135.200 ;
        RECT 156.600 133.800 157.000 134.200 ;
        RECT 153.400 131.800 153.800 132.200 ;
        RECT 151.800 130.800 152.200 131.200 ;
        RECT 150.200 128.800 150.600 129.200 ;
        RECT 150.200 128.200 150.500 128.800 ;
        RECT 150.200 127.800 150.600 128.200 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 146.200 116.800 146.600 117.200 ;
        RECT 139.800 115.800 140.200 116.200 ;
        RECT 143.000 116.100 143.400 116.200 ;
        RECT 143.800 116.100 144.200 116.200 ;
        RECT 143.000 115.800 144.200 116.100 ;
        RECT 146.200 115.800 146.600 116.200 ;
        RECT 146.200 115.200 146.500 115.800 ;
        RECT 139.800 114.800 140.200 115.200 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 139.800 111.200 140.100 114.800 ;
        RECT 140.600 113.800 141.000 114.200 ;
        RECT 139.800 110.800 140.200 111.200 ;
        RECT 139.000 109.800 140.100 110.100 ;
        RECT 135.800 108.800 136.200 109.200 ;
        RECT 135.000 104.800 135.400 105.200 ;
        RECT 136.600 104.800 137.000 105.200 ;
        RECT 135.000 104.200 135.300 104.800 ;
        RECT 135.000 103.800 135.400 104.200 ;
        RECT 136.600 99.200 136.900 104.800 ;
        RECT 138.200 103.100 138.600 108.900 ;
        RECT 139.800 99.200 140.100 109.800 ;
        RECT 140.600 104.200 140.900 113.800 ;
        RECT 142.200 111.800 142.600 112.200 ;
        RECT 143.800 111.800 144.200 112.200 ;
        RECT 142.200 108.200 142.500 111.800 ;
        RECT 142.200 107.800 142.600 108.200 ;
        RECT 142.200 105.900 142.600 106.300 ;
        RECT 142.200 105.200 142.500 105.900 ;
        RECT 142.200 104.800 142.600 105.200 ;
        RECT 140.600 103.800 141.000 104.200 ;
        RECT 143.000 103.100 143.400 108.900 ;
        RECT 143.800 105.200 144.100 111.800 ;
        RECT 143.800 104.800 144.200 105.200 ;
        RECT 144.600 105.100 145.000 107.900 ;
        RECT 134.200 98.800 134.600 99.200 ;
        RECT 136.600 98.800 137.000 99.200 ;
        RECT 139.800 98.800 140.200 99.200 ;
        RECT 135.000 95.800 135.400 96.200 ;
        RECT 135.000 95.200 135.300 95.800 ;
        RECT 135.000 94.800 135.400 95.200 ;
        RECT 133.400 94.100 133.800 94.200 ;
        RECT 134.200 94.100 134.600 94.200 ;
        RECT 133.400 93.800 134.600 94.100 ;
        RECT 139.000 93.800 139.400 94.200 ;
        RECT 139.800 93.800 140.200 94.200 ;
        RECT 141.400 93.800 141.800 94.200 ;
        RECT 136.600 91.800 137.000 92.200 ;
        RECT 132.600 90.800 133.000 91.200 ;
        RECT 132.600 89.800 133.000 90.200 ;
        RECT 128.600 85.800 129.000 86.200 ;
        RECT 131.800 85.800 132.200 86.200 ;
        RECT 128.600 85.200 128.900 85.800 ;
        RECT 128.600 84.800 129.000 85.200 ;
        RECT 131.000 76.800 131.400 77.200 ;
        RECT 127.800 75.800 128.200 76.200 ;
        RECT 123.000 75.200 123.300 75.800 ;
        RECT 122.200 74.800 122.600 75.200 ;
        RECT 123.000 74.800 123.400 75.200 ;
        RECT 123.800 74.800 124.200 75.200 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 127.800 74.800 128.200 75.200 ;
        RECT 128.600 75.100 129.000 75.200 ;
        RECT 129.400 75.100 129.800 75.200 ;
        RECT 128.600 74.800 129.800 75.100 ;
        RECT 123.000 72.800 123.400 73.200 ;
        RECT 123.000 72.200 123.300 72.800 ;
        RECT 123.000 71.800 123.400 72.200 ;
        RECT 123.800 69.200 124.100 74.800 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 124.600 73.200 124.900 73.800 ;
        RECT 124.600 72.800 125.000 73.200 ;
        RECT 121.400 63.100 121.800 68.900 ;
        RECT 123.800 68.800 124.200 69.200 ;
        RECT 122.200 66.800 122.600 67.200 ;
        RECT 125.400 66.800 125.800 67.200 ;
        RECT 122.200 66.200 122.500 66.800 ;
        RECT 125.400 66.300 125.700 66.800 ;
        RECT 122.200 65.800 122.600 66.200 ;
        RECT 125.400 65.900 125.800 66.300 ;
        RECT 125.400 65.800 125.700 65.900 ;
        RECT 120.600 60.800 121.000 61.200 ;
        RECT 115.000 59.100 115.400 59.200 ;
        RECT 115.800 59.100 116.200 59.200 ;
        RECT 115.000 58.800 116.200 59.100 ;
        RECT 115.000 57.800 115.400 58.200 ;
        RECT 114.200 52.800 114.600 53.200 ;
        RECT 113.400 50.800 113.800 51.200 ;
        RECT 114.200 50.200 114.500 52.800 ;
        RECT 114.200 49.800 114.600 50.200 ;
        RECT 109.400 48.800 109.800 49.200 ;
        RECT 112.600 48.800 113.000 49.200 ;
        RECT 112.600 48.200 112.900 48.800 ;
        RECT 112.600 47.800 113.000 48.200 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 103.800 46.800 105.000 47.100 ;
        RECT 107.000 46.800 107.400 47.200 ;
        RECT 107.800 46.800 108.200 47.200 ;
        RECT 103.800 46.200 104.100 46.800 ;
        RECT 103.800 45.800 104.200 46.200 ;
        RECT 104.600 45.800 105.000 46.200 ;
        RECT 107.000 46.100 107.400 46.200 ;
        RECT 107.800 46.100 108.200 46.200 ;
        RECT 107.000 45.800 108.200 46.100 ;
        RECT 111.000 45.800 111.400 46.200 ;
        RECT 104.600 45.200 104.900 45.800 ;
        RECT 104.600 44.800 105.000 45.200 ;
        RECT 111.000 44.200 111.300 45.800 ;
        RECT 111.000 43.800 111.400 44.200 ;
        RECT 102.200 38.800 102.600 39.200 ;
        RECT 111.000 38.200 111.300 43.800 ;
        RECT 98.200 37.800 98.600 38.200 ;
        RECT 111.000 37.800 111.400 38.200 ;
        RECT 98.200 35.200 98.500 37.800 ;
        RECT 110.200 36.800 110.600 37.200 ;
        RECT 107.800 35.800 108.200 36.200 ;
        RECT 108.600 35.800 109.000 36.200 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 98.200 34.800 98.600 35.200 ;
        RECT 101.400 34.800 101.800 35.200 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 104.600 34.800 105.000 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 106.200 35.100 106.600 35.200 ;
        RECT 105.400 34.800 106.600 35.100 ;
        RECT 96.600 33.800 97.000 34.200 ;
        RECT 96.600 33.200 96.900 33.800 ;
        RECT 96.600 32.800 97.000 33.200 ;
        RECT 101.400 32.200 101.700 34.800 ;
        RECT 103.800 33.100 104.100 34.800 ;
        RECT 104.600 34.200 104.900 34.800 ;
        RECT 107.800 34.200 108.100 35.800 ;
        RECT 108.600 35.200 108.900 35.800 ;
        RECT 108.600 34.800 109.000 35.200 ;
        RECT 110.200 34.200 110.500 36.800 ;
        RECT 104.600 33.800 105.000 34.200 ;
        RECT 105.400 33.800 105.800 34.200 ;
        RECT 107.800 33.800 108.200 34.200 ;
        RECT 110.200 33.800 110.600 34.200 ;
        RECT 105.400 33.200 105.700 33.800 ;
        RECT 103.800 32.800 104.900 33.100 ;
        RECT 105.400 32.800 105.800 33.200 ;
        RECT 111.000 33.100 111.400 35.900 ;
        RECT 111.800 32.800 112.200 33.200 ;
        RECT 96.600 31.800 97.000 32.200 ;
        RECT 101.400 31.800 101.800 32.200 ;
        RECT 96.600 29.200 96.900 31.800 ;
        RECT 96.600 29.100 97.000 29.200 ;
        RECT 97.400 29.100 97.800 29.200 ;
        RECT 96.600 28.800 97.800 29.100 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 95.800 26.200 96.100 26.800 ;
        RECT 95.800 25.800 96.200 26.200 ;
        RECT 95.000 20.800 95.400 21.200 ;
        RECT 88.600 19.800 89.000 20.200 ;
        RECT 88.600 19.200 88.900 19.800 ;
        RECT 95.800 19.200 96.100 25.800 ;
        RECT 99.000 23.100 99.400 28.900 ;
        RECT 99.800 26.800 100.200 27.200 ;
        RECT 103.000 26.800 103.400 27.200 ;
        RECT 99.800 26.200 100.100 26.800 ;
        RECT 103.000 26.300 103.300 26.800 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 103.000 25.900 103.400 26.300 ;
        RECT 103.800 23.100 104.200 28.900 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 95.800 18.800 96.200 19.200 ;
        RECT 99.800 15.800 100.200 16.200 ;
        RECT 103.000 15.800 103.400 16.200 ;
        RECT 99.800 15.200 100.100 15.800 ;
        RECT 103.000 15.200 103.300 15.800 ;
        RECT 99.800 14.800 100.200 15.200 ;
        RECT 102.200 14.800 102.600 15.200 ;
        RECT 103.000 14.800 103.400 15.200 ;
        RECT 103.800 14.800 104.200 15.200 ;
        RECT 102.200 14.200 102.500 14.800 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 83.000 14.100 83.400 14.200 ;
        RECT 82.200 13.800 83.400 14.100 ;
        RECT 86.200 13.800 86.600 14.200 ;
        RECT 102.200 13.800 102.600 14.200 ;
        RECT 100.600 13.100 101.000 13.200 ;
        RECT 101.400 13.100 101.800 13.200 ;
        RECT 100.600 12.800 101.800 13.100 ;
        RECT 103.800 12.200 104.100 14.800 ;
        RECT 104.600 14.200 104.900 32.800 ;
        RECT 106.200 28.800 106.600 29.200 ;
        RECT 105.400 25.100 105.800 27.900 ;
        RECT 106.200 27.200 106.500 28.800 ;
        RECT 111.000 27.800 111.400 28.200 ;
        RECT 111.000 27.200 111.300 27.800 ;
        RECT 111.800 27.200 112.100 32.800 ;
        RECT 112.600 32.100 113.000 37.900 ;
        RECT 113.400 35.800 113.800 36.200 ;
        RECT 113.400 35.100 113.700 35.800 ;
        RECT 113.400 34.700 113.800 35.100 ;
        RECT 114.200 28.800 114.600 29.200 ;
        RECT 114.200 28.200 114.500 28.800 ;
        RECT 114.200 27.800 114.600 28.200 ;
        RECT 106.200 26.800 106.600 27.200 ;
        RECT 107.800 27.100 108.200 27.200 ;
        RECT 108.600 27.100 109.000 27.200 ;
        RECT 107.800 26.800 109.000 27.100 ;
        RECT 110.200 26.800 110.600 27.200 ;
        RECT 111.000 26.800 111.400 27.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 110.200 26.200 110.500 26.800 ;
        RECT 107.800 25.800 108.200 26.200 ;
        RECT 110.200 25.800 110.600 26.200 ;
        RECT 111.000 25.800 111.400 26.200 ;
        RECT 107.800 25.200 108.100 25.800 ;
        RECT 107.800 24.800 108.200 25.200 ;
        RECT 107.800 22.800 108.200 23.200 ;
        RECT 107.000 17.800 107.400 18.200 ;
        RECT 107.000 15.200 107.300 17.800 ;
        RECT 107.800 15.200 108.100 22.800 ;
        RECT 108.600 16.800 109.000 17.200 ;
        RECT 108.600 15.200 108.900 16.800 ;
        RECT 109.400 16.100 109.800 16.200 ;
        RECT 110.200 16.100 110.600 16.200 ;
        RECT 109.400 15.800 110.600 16.100 ;
        RECT 107.000 14.800 107.400 15.200 ;
        RECT 107.800 14.800 108.200 15.200 ;
        RECT 108.600 14.800 109.000 15.200 ;
        RECT 108.600 14.200 108.900 14.800 ;
        RECT 104.600 13.800 105.000 14.200 ;
        RECT 108.600 13.800 109.000 14.200 ;
        RECT 91.000 11.800 91.400 12.200 ;
        RECT 95.800 11.800 96.200 12.200 ;
        RECT 100.600 11.800 101.000 12.200 ;
        RECT 103.800 11.800 104.200 12.200 ;
        RECT 91.000 9.200 91.300 11.800 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 75.800 6.800 76.200 7.200 ;
        RECT 75.800 6.200 76.100 6.800 ;
        RECT 75.800 5.800 76.200 6.200 ;
        RECT 79.000 3.100 79.400 8.900 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 87.000 8.800 87.400 9.200 ;
        RECT 89.400 8.800 89.800 9.200 ;
        RECT 91.000 8.800 91.400 9.200 ;
        RECT 87.000 7.200 87.300 8.800 ;
        RECT 89.400 8.200 89.700 8.800 ;
        RECT 89.400 7.800 89.800 8.200 ;
        RECT 83.800 7.100 84.200 7.200 ;
        RECT 84.600 7.100 85.000 7.200 ;
        RECT 83.800 6.800 85.000 7.100 ;
        RECT 86.200 6.800 86.600 7.200 ;
        RECT 87.000 6.800 87.400 7.200 ;
        RECT 86.200 6.200 86.500 6.800 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 87.000 6.100 87.400 6.200 ;
        RECT 87.800 6.100 88.200 6.200 ;
        RECT 87.000 5.800 88.200 6.100 ;
        RECT 86.200 5.200 86.500 5.800 ;
        RECT 83.800 5.100 84.200 5.200 ;
        RECT 84.600 5.100 85.000 5.200 ;
        RECT 83.800 4.800 85.000 5.100 ;
        RECT 86.200 4.800 86.600 5.200 ;
        RECT 93.400 3.100 93.800 8.900 ;
        RECT 95.800 8.200 96.100 11.800 ;
        RECT 95.800 7.800 96.200 8.200 ;
        RECT 95.800 7.200 96.100 7.800 ;
        RECT 95.800 6.800 96.200 7.200 ;
        RECT 96.600 6.200 97.000 6.300 ;
        RECT 97.400 6.200 97.800 6.300 ;
        RECT 96.600 5.900 97.800 6.200 ;
        RECT 98.200 3.100 98.600 8.900 ;
        RECT 99.800 5.100 100.200 7.900 ;
        RECT 100.600 7.200 100.900 11.800 ;
        RECT 107.000 8.800 107.400 9.200 ;
        RECT 107.000 7.200 107.300 8.800 ;
        RECT 107.800 7.800 108.200 8.200 ;
        RECT 107.800 7.200 108.100 7.800 ;
        RECT 111.000 7.200 111.300 25.800 ;
        RECT 111.800 19.200 112.100 26.800 ;
        RECT 115.000 26.200 115.300 57.800 ;
        RECT 118.200 56.800 118.600 57.200 ;
        RECT 120.600 56.800 121.000 57.200 ;
        RECT 118.200 56.200 118.500 56.800 ;
        RECT 116.600 56.100 117.000 56.200 ;
        RECT 117.400 56.100 117.800 56.200 ;
        RECT 116.600 55.800 117.800 56.100 ;
        RECT 118.200 55.800 118.600 56.200 ;
        RECT 120.600 55.200 120.900 56.800 ;
        RECT 120.600 54.800 121.000 55.200 ;
        RECT 121.400 54.800 121.800 55.200 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 118.200 53.200 118.500 53.800 ;
        RECT 118.200 52.800 118.600 53.200 ;
        RECT 119.800 53.100 120.200 53.200 ;
        RECT 120.600 53.100 121.000 53.200 ;
        RECT 119.800 52.800 121.000 53.100 ;
        RECT 119.800 51.800 120.200 52.200 ;
        RECT 121.400 52.100 121.700 54.800 ;
        RECT 120.600 51.800 121.700 52.100 ;
        RECT 119.000 50.800 119.400 51.200 ;
        RECT 119.000 47.200 119.300 50.800 ;
        RECT 118.200 46.800 118.600 47.200 ;
        RECT 119.000 46.800 119.400 47.200 ;
        RECT 115.800 34.800 116.200 35.200 ;
        RECT 112.600 26.100 113.000 26.200 ;
        RECT 113.400 26.100 113.800 26.200 ;
        RECT 112.600 25.800 113.800 26.100 ;
        RECT 115.000 25.800 115.400 26.200 ;
        RECT 115.000 25.200 115.300 25.800 ;
        RECT 115.000 24.800 115.400 25.200 ;
        RECT 111.800 18.800 112.200 19.200 ;
        RECT 115.800 17.200 116.100 34.800 ;
        RECT 117.400 32.100 117.800 37.900 ;
        RECT 118.200 37.200 118.500 46.800 ;
        RECT 119.800 46.200 120.100 51.800 ;
        RECT 119.800 45.800 120.200 46.200 ;
        RECT 120.600 45.200 120.900 51.800 ;
        RECT 122.200 48.200 122.500 65.800 ;
        RECT 123.000 63.800 123.400 64.200 ;
        RECT 123.000 59.200 123.300 63.800 ;
        RECT 126.200 63.100 126.600 68.900 ;
        RECT 127.000 64.200 127.300 74.800 ;
        RECT 127.800 72.200 128.100 74.800 ;
        RECT 131.000 74.200 131.300 76.800 ;
        RECT 132.600 75.200 132.900 89.800 ;
        RECT 133.400 83.100 133.800 88.900 ;
        RECT 135.800 88.800 136.200 89.200 ;
        RECT 134.200 86.800 134.600 87.200 ;
        RECT 134.200 86.200 134.500 86.800 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 135.000 85.800 135.400 86.200 ;
        RECT 135.000 85.200 135.300 85.800 ;
        RECT 135.000 84.800 135.400 85.200 ;
        RECT 133.400 75.800 133.800 76.200 ;
        RECT 133.400 75.200 133.700 75.800 ;
        RECT 131.800 74.800 132.200 75.200 ;
        RECT 132.600 74.800 133.000 75.200 ;
        RECT 133.400 74.800 133.800 75.200 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 135.000 75.100 135.400 75.200 ;
        RECT 134.200 74.800 135.400 75.100 ;
        RECT 131.800 74.200 132.100 74.800 ;
        RECT 129.400 73.800 129.800 74.200 ;
        RECT 131.000 73.800 131.400 74.200 ;
        RECT 131.800 73.800 132.200 74.200 ;
        RECT 129.400 73.200 129.700 73.800 ;
        RECT 129.400 72.800 129.800 73.200 ;
        RECT 127.800 71.800 128.200 72.200 ;
        RECT 129.400 71.800 129.800 72.200 ;
        RECT 129.400 71.200 129.700 71.800 ;
        RECT 129.400 70.800 129.800 71.200 ;
        RECT 132.600 70.800 133.000 71.200 ;
        RECT 128.600 68.800 129.000 69.200 ;
        RECT 127.800 65.100 128.200 67.900 ;
        RECT 128.600 67.200 128.900 68.800 ;
        RECT 128.600 66.800 129.000 67.200 ;
        RECT 130.200 67.100 130.600 67.200 ;
        RECT 131.000 67.100 131.400 67.200 ;
        RECT 130.200 66.800 131.400 67.100 ;
        RECT 132.600 66.200 132.900 70.800 ;
        RECT 133.400 67.800 133.800 68.200 ;
        RECT 133.400 67.200 133.700 67.800 ;
        RECT 135.800 67.200 136.100 88.800 ;
        RECT 136.600 78.200 136.900 91.800 ;
        RECT 138.200 83.100 138.600 88.900 ;
        RECT 137.400 78.800 137.800 79.200 ;
        RECT 136.600 77.800 137.000 78.200 ;
        RECT 136.600 75.800 137.000 76.200 ;
        RECT 136.600 75.200 136.900 75.800 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 137.400 74.200 137.700 78.800 ;
        RECT 139.000 75.200 139.300 93.800 ;
        RECT 139.800 93.200 140.100 93.800 ;
        RECT 139.800 92.800 140.200 93.200 ;
        RECT 140.600 88.800 141.000 89.200 ;
        RECT 139.800 85.100 140.200 87.900 ;
        RECT 140.600 87.200 140.900 88.800 ;
        RECT 140.600 86.800 141.000 87.200 ;
        RECT 140.600 84.100 141.000 84.200 ;
        RECT 139.800 83.800 141.000 84.100 ;
        RECT 139.800 79.200 140.100 83.800 ;
        RECT 141.400 79.200 141.700 93.800 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 143.000 92.200 143.300 92.800 ;
        RECT 146.200 92.200 146.500 114.800 ;
        RECT 147.000 114.100 147.400 114.200 ;
        RECT 147.800 114.100 148.200 114.200 ;
        RECT 147.000 113.800 148.200 114.100 ;
        RECT 148.600 112.100 149.000 112.200 ;
        RECT 149.400 112.100 149.800 112.200 ;
        RECT 151.000 112.100 151.400 117.900 ;
        RECT 151.800 115.200 152.100 130.800 ;
        RECT 152.600 123.100 153.000 128.900 ;
        RECT 153.400 124.200 153.700 131.800 ;
        RECT 156.600 131.200 156.900 133.800 ;
        RECT 157.400 132.100 157.800 137.900 ;
        RECT 156.600 130.800 157.000 131.200 ;
        RECT 154.200 128.800 154.600 129.200 ;
        RECT 154.200 127.200 154.500 128.800 ;
        RECT 154.200 126.800 154.600 127.200 ;
        RECT 155.800 126.200 156.200 126.300 ;
        RECT 156.600 126.200 157.000 126.300 ;
        RECT 155.800 125.900 157.000 126.200 ;
        RECT 153.400 123.800 153.800 124.200 ;
        RECT 157.400 123.100 157.800 128.900 ;
        RECT 158.200 127.200 158.500 141.800 ;
        RECT 159.000 134.800 159.400 135.200 ;
        RECT 159.000 134.200 159.300 134.800 ;
        RECT 159.000 133.800 159.400 134.200 ;
        RECT 158.200 126.800 158.600 127.200 ;
        RECT 159.000 125.100 159.400 127.900 ;
        RECT 159.800 127.800 160.200 128.200 ;
        RECT 159.800 127.200 160.100 127.800 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 160.600 125.200 160.900 155.800 ;
        RECT 163.000 152.100 163.400 157.900 ;
        RECT 163.800 156.200 164.100 166.800 ;
        RECT 164.600 166.200 164.900 168.800 ;
        RECT 165.400 167.200 165.700 169.800 ;
        RECT 165.400 166.800 165.800 167.200 ;
        RECT 167.800 167.100 168.200 167.200 ;
        RECT 168.600 167.100 169.000 167.200 ;
        RECT 167.800 166.800 169.000 167.100 ;
        RECT 170.200 166.800 170.600 167.200 ;
        RECT 171.000 166.800 171.400 167.200 ;
        RECT 170.200 166.200 170.500 166.800 ;
        RECT 171.000 166.200 171.300 166.800 ;
        RECT 164.600 165.800 165.000 166.200 ;
        RECT 165.400 165.800 165.800 166.200 ;
        RECT 170.200 165.800 170.600 166.200 ;
        RECT 171.000 165.800 171.400 166.200 ;
        RECT 171.800 165.800 172.200 166.200 ;
        RECT 165.400 165.200 165.700 165.800 ;
        RECT 165.400 164.800 165.800 165.200 ;
        RECT 167.800 165.100 168.200 165.200 ;
        RECT 168.600 165.100 169.000 165.200 ;
        RECT 167.800 164.800 169.000 165.100 ;
        RECT 163.800 155.800 164.200 156.200 ;
        RECT 163.000 150.800 163.400 151.200 ;
        RECT 161.400 148.800 161.800 149.200 ;
        RECT 161.400 147.200 161.700 148.800 ;
        RECT 161.400 146.800 161.800 147.200 ;
        RECT 162.200 145.100 162.600 147.900 ;
        RECT 163.000 147.200 163.300 150.800 ;
        RECT 163.000 146.800 163.400 147.200 ;
        RECT 163.800 143.100 164.200 148.900 ;
        RECT 164.600 146.800 165.000 147.200 ;
        RECT 164.600 146.300 164.900 146.800 ;
        RECT 164.600 145.900 165.000 146.300 ;
        RECT 162.200 132.100 162.600 137.900 ;
        RECT 164.600 136.800 165.000 137.200 ;
        RECT 164.600 135.200 164.900 136.800 ;
        RECT 165.400 136.200 165.700 164.800 ;
        RECT 171.800 162.200 172.100 165.800 ;
        RECT 171.800 161.800 172.200 162.200 ;
        RECT 166.200 154.800 166.600 155.200 ;
        RECT 166.200 154.200 166.500 154.800 ;
        RECT 166.200 153.800 166.600 154.200 ;
        RECT 167.800 152.100 168.200 157.900 ;
        RECT 168.600 153.800 169.000 154.200 ;
        RECT 168.600 150.200 168.900 153.800 ;
        RECT 169.400 153.100 169.800 155.900 ;
        RECT 171.800 155.800 172.200 156.200 ;
        RECT 171.800 154.200 172.100 155.800 ;
        RECT 172.600 154.200 172.900 169.800 ;
        RECT 181.400 169.200 181.700 180.800 ;
        RECT 183.000 172.100 183.400 177.900 ;
        RECT 183.800 174.800 184.200 175.200 ;
        RECT 183.800 174.200 184.100 174.800 ;
        RECT 183.800 173.800 184.200 174.200 ;
        RECT 177.400 169.100 177.800 169.200 ;
        RECT 178.200 169.100 178.600 169.200 ;
        RECT 177.400 168.800 178.600 169.100 ;
        RECT 181.400 168.800 181.800 169.200 ;
        RECT 182.200 168.800 182.600 169.200 ;
        RECT 183.000 168.800 183.400 169.200 ;
        RECT 174.200 167.800 174.600 168.200 ;
        RECT 174.200 166.200 174.500 167.800 ;
        RECT 182.200 167.200 182.500 168.800 ;
        RECT 183.000 168.200 183.300 168.800 ;
        RECT 183.000 167.800 183.400 168.200 ;
        RECT 175.000 166.800 175.400 167.200 ;
        RECT 182.200 166.800 182.600 167.200 ;
        RECT 175.000 166.200 175.300 166.800 ;
        RECT 173.400 166.100 173.800 166.200 ;
        RECT 174.200 166.100 174.600 166.200 ;
        RECT 173.400 165.800 174.600 166.100 ;
        RECT 175.000 165.800 175.400 166.200 ;
        RECT 175.800 165.800 176.200 166.200 ;
        RECT 176.600 166.100 177.000 166.200 ;
        RECT 177.400 166.100 177.800 166.200 ;
        RECT 176.600 165.800 177.800 166.100 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 175.800 165.200 176.100 165.800 ;
        RECT 175.800 164.800 176.200 165.200 ;
        RECT 179.800 159.200 180.100 165.800 ;
        RECT 180.600 164.800 181.000 165.200 ;
        RECT 180.600 164.200 180.900 164.800 ;
        RECT 180.600 163.800 181.000 164.200 ;
        RECT 179.800 158.800 180.200 159.200 ;
        RECT 173.400 156.800 173.800 157.200 ;
        RECT 175.800 156.800 176.200 157.200 ;
        RECT 183.000 156.800 183.400 157.200 ;
        RECT 173.400 155.200 173.700 156.800 ;
        RECT 175.800 156.200 176.100 156.800 ;
        RECT 175.000 155.800 175.400 156.200 ;
        RECT 175.800 155.800 176.200 156.200 ;
        RECT 182.200 155.800 182.600 156.200 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 175.000 154.200 175.300 155.800 ;
        RECT 182.200 155.200 182.500 155.800 ;
        RECT 177.400 155.100 177.800 155.200 ;
        RECT 178.200 155.100 178.600 155.200 ;
        RECT 177.400 154.800 178.600 155.100 ;
        RECT 179.000 154.800 179.400 155.200 ;
        RECT 182.200 154.800 182.600 155.200 ;
        RECT 179.000 154.200 179.300 154.800 ;
        RECT 183.000 154.200 183.300 156.800 ;
        RECT 170.200 153.800 170.600 154.200 ;
        RECT 171.800 153.800 172.200 154.200 ;
        RECT 172.600 153.800 173.000 154.200 ;
        RECT 173.400 153.800 173.800 154.200 ;
        RECT 175.000 153.800 175.400 154.200 ;
        RECT 177.400 154.100 177.800 154.200 ;
        RECT 178.200 154.100 178.600 154.200 ;
        RECT 177.400 153.800 178.600 154.100 ;
        RECT 179.000 153.800 179.400 154.200 ;
        RECT 183.000 153.800 183.400 154.200 ;
        RECT 170.200 153.200 170.500 153.800 ;
        RECT 170.200 152.800 170.600 153.200 ;
        RECT 171.800 151.800 172.200 152.200 ;
        RECT 168.600 149.800 169.000 150.200 ;
        RECT 166.200 148.800 166.600 149.200 ;
        RECT 170.200 149.100 170.600 149.200 ;
        RECT 171.000 149.100 171.400 149.200 ;
        RECT 165.400 135.800 165.800 136.200 ;
        RECT 166.200 135.200 166.500 148.800 ;
        RECT 167.800 146.800 168.200 147.200 ;
        RECT 167.800 146.200 168.100 146.800 ;
        RECT 167.800 145.800 168.200 146.200 ;
        RECT 168.600 143.100 169.000 148.900 ;
        RECT 170.200 148.800 171.400 149.100 ;
        RECT 171.800 145.200 172.100 151.800 ;
        RECT 172.600 148.200 172.900 153.800 ;
        RECT 172.600 147.800 173.000 148.200 ;
        RECT 173.400 146.200 173.700 153.800 ;
        RECT 175.000 152.800 175.400 153.200 ;
        RECT 175.000 149.200 175.300 152.800 ;
        RECT 178.200 149.800 178.600 150.200 ;
        RECT 175.000 148.800 175.400 149.200 ;
        RECT 174.200 147.800 174.600 148.200 ;
        RECT 174.200 147.200 174.500 147.800 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 172.600 145.800 173.000 146.200 ;
        RECT 173.400 145.800 173.800 146.200 ;
        RECT 172.600 145.200 172.900 145.800 ;
        RECT 171.800 144.800 172.200 145.200 ;
        RECT 172.600 144.800 173.000 145.200 ;
        RECT 167.800 136.800 168.200 137.200 ;
        RECT 167.800 136.200 168.100 136.800 ;
        RECT 167.800 135.800 168.200 136.200 ;
        RECT 171.800 135.800 172.200 136.200 ;
        RECT 171.800 135.200 172.100 135.800 ;
        RECT 164.600 134.800 165.000 135.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 168.600 135.100 169.000 135.200 ;
        RECT 169.400 135.100 169.800 135.200 ;
        RECT 168.600 134.800 169.800 135.100 ;
        RECT 171.800 134.800 172.200 135.200 ;
        RECT 164.600 129.800 165.000 130.200 ;
        RECT 164.600 127.200 164.900 129.800 ;
        RECT 165.400 129.200 165.700 134.800 ;
        RECT 171.800 134.100 172.200 134.200 ;
        RECT 172.600 134.100 173.000 134.200 ;
        RECT 171.800 133.800 173.000 134.100 ;
        RECT 169.400 130.800 169.800 131.200 ;
        RECT 165.400 128.800 165.800 129.200 ;
        RECT 161.400 126.800 161.800 127.200 ;
        RECT 164.600 126.800 165.000 127.200 ;
        RECT 161.400 126.200 161.700 126.800 ;
        RECT 161.400 125.800 161.800 126.200 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 165.400 125.800 165.800 126.200 ;
        RECT 166.200 125.800 166.600 126.200 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 163.800 125.200 164.100 125.800 ;
        RECT 160.600 125.100 161.000 125.200 ;
        RECT 161.400 125.100 161.800 125.200 ;
        RECT 160.600 124.800 161.800 125.100 ;
        RECT 163.800 124.800 164.200 125.200 ;
        RECT 154.200 115.800 154.600 116.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 148.600 111.800 149.800 112.100 ;
        RECT 153.400 111.800 153.800 112.200 ;
        RECT 148.600 110.800 149.000 111.200 ;
        RECT 147.000 102.800 147.400 103.200 ;
        RECT 147.000 99.200 147.300 102.800 ;
        RECT 147.000 98.800 147.400 99.200 ;
        RECT 148.600 94.200 148.900 110.800 ;
        RECT 153.400 107.200 153.700 111.800 ;
        RECT 153.400 106.800 153.800 107.200 ;
        RECT 151.800 105.800 152.200 106.200 ;
        RECT 148.600 93.800 149.000 94.200 ;
        RECT 143.000 91.800 143.400 92.200 ;
        RECT 146.200 91.800 146.600 92.200 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 143.000 90.200 143.300 91.800 ;
        RECT 146.200 90.200 146.500 91.800 ;
        RECT 147.000 91.200 147.300 91.800 ;
        RECT 147.000 90.800 147.400 91.200 ;
        RECT 143.000 89.800 143.400 90.200 ;
        RECT 146.200 89.800 146.600 90.200 ;
        RECT 143.000 83.100 143.400 88.900 ;
        RECT 146.200 86.200 146.600 86.300 ;
        RECT 147.000 86.200 147.400 86.300 ;
        RECT 144.600 85.800 145.000 86.200 ;
        RECT 146.200 85.900 147.400 86.200 ;
        RECT 142.200 79.800 142.600 80.200 ;
        RECT 139.800 78.800 140.200 79.200 ;
        RECT 141.400 78.800 141.800 79.200 ;
        RECT 142.200 76.200 142.500 79.800 ;
        RECT 143.800 77.800 144.200 78.200 ;
        RECT 142.200 75.800 142.600 76.200 ;
        RECT 138.200 75.100 138.600 75.200 ;
        RECT 139.000 75.100 139.400 75.200 ;
        RECT 138.200 74.800 139.400 75.100 ;
        RECT 140.600 74.800 141.000 75.200 ;
        RECT 140.600 74.200 140.900 74.800 ;
        RECT 137.400 73.800 137.800 74.200 ;
        RECT 140.600 73.800 141.000 74.200 ;
        RECT 141.400 71.800 141.800 72.200 ;
        RECT 141.400 71.200 141.700 71.800 ;
        RECT 142.200 71.200 142.500 75.800 ;
        RECT 141.400 70.800 141.800 71.200 ;
        RECT 142.200 70.800 142.600 71.200 ;
        RECT 143.800 70.200 144.100 77.800 ;
        RECT 143.800 69.800 144.200 70.200 ;
        RECT 139.000 67.800 139.400 68.200 ;
        RECT 133.400 66.800 133.800 67.200 ;
        RECT 135.000 67.100 135.400 67.200 ;
        RECT 135.800 67.100 136.200 67.200 ;
        RECT 135.000 66.800 136.200 67.100 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 137.400 66.200 137.700 66.800 ;
        RECT 130.200 65.800 130.600 66.200 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 136.600 66.100 137.000 66.200 ;
        RECT 135.800 65.800 137.000 66.100 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 130.200 65.200 130.500 65.800 ;
        RECT 130.200 64.800 130.600 65.200 ;
        RECT 127.000 63.800 127.400 64.200 ;
        RECT 125.400 59.800 125.800 60.200 ;
        RECT 123.000 58.800 123.400 59.200 ;
        RECT 125.400 56.200 125.700 59.800 ;
        RECT 125.400 55.800 125.800 56.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 123.800 53.200 124.100 54.800 ;
        RECT 127.000 54.200 127.300 63.800 ;
        RECT 129.400 62.800 129.800 63.200 ;
        RECT 129.400 60.200 129.700 62.800 ;
        RECT 129.400 59.800 129.800 60.200 ;
        RECT 129.400 55.200 129.700 59.800 ;
        RECT 137.400 59.200 137.700 65.800 ;
        RECT 139.000 61.200 139.300 67.800 ;
        RECT 139.800 65.100 140.200 67.900 ;
        RECT 139.800 63.800 140.200 64.200 ;
        RECT 139.000 60.800 139.400 61.200 ;
        RECT 139.800 59.200 140.100 63.800 ;
        RECT 141.400 63.100 141.800 68.900 ;
        RECT 142.200 66.100 142.600 66.300 ;
        RECT 143.000 66.100 143.400 66.200 ;
        RECT 142.200 65.800 143.400 66.100 ;
        RECT 143.000 63.800 143.400 64.200 ;
        RECT 137.400 58.800 137.800 59.200 ;
        RECT 139.800 58.800 140.200 59.200 ;
        RECT 127.800 55.100 128.200 55.200 ;
        RECT 128.600 55.100 129.000 55.200 ;
        RECT 127.800 54.800 129.000 55.100 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 127.000 53.800 127.400 54.200 ;
        RECT 129.400 53.800 129.800 54.200 ;
        RECT 130.200 53.800 130.600 54.200 ;
        RECT 123.800 52.800 124.200 53.200 ;
        RECT 122.200 47.800 122.600 48.200 ;
        RECT 121.400 47.100 121.800 47.200 ;
        RECT 122.200 47.100 122.600 47.200 ;
        RECT 121.400 46.800 122.600 47.100 ;
        RECT 123.800 46.800 124.200 47.200 ;
        RECT 122.200 45.800 122.600 46.200 ;
        RECT 122.200 45.200 122.500 45.800 ;
        RECT 120.600 44.800 121.000 45.200 ;
        RECT 122.200 44.800 122.600 45.200 ;
        RECT 123.800 44.200 124.100 46.800 ;
        RECT 123.800 43.800 124.200 44.200 ;
        RECT 120.600 41.800 121.000 42.200 ;
        RECT 118.200 36.800 118.600 37.200 ;
        RECT 119.000 37.100 119.400 37.200 ;
        RECT 119.800 37.100 120.200 37.200 ;
        RECT 119.000 36.800 120.200 37.100 ;
        RECT 120.600 35.200 120.900 41.800 ;
        RECT 122.200 39.800 122.600 40.200 ;
        RECT 122.200 39.200 122.500 39.800 ;
        RECT 122.200 38.800 122.600 39.200 ;
        RECT 121.400 36.800 121.800 37.200 ;
        RECT 121.400 35.200 121.700 36.800 ;
        RECT 123.800 35.200 124.100 43.800 ;
        RECT 127.000 43.100 127.400 48.900 ;
        RECT 127.800 47.800 128.200 48.200 ;
        RECT 127.800 46.200 128.100 47.800 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 128.600 36.800 129.000 37.200 ;
        RECT 128.600 35.200 128.900 36.800 ;
        RECT 129.400 35.200 129.700 53.800 ;
        RECT 130.200 51.200 130.500 53.800 ;
        RECT 131.000 53.100 131.400 55.900 ;
        RECT 132.600 52.100 133.000 57.900 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 133.400 55.100 133.700 55.800 ;
        RECT 133.400 54.700 133.800 55.100 ;
        RECT 133.400 52.800 133.800 53.200 ;
        RECT 130.200 50.800 130.600 51.200 ;
        RECT 133.400 51.100 133.700 52.800 ;
        RECT 137.400 52.100 137.800 57.900 ;
        RECT 140.600 54.800 141.000 55.200 ;
        RECT 140.600 51.200 140.900 54.800 ;
        RECT 141.400 54.100 141.800 54.200 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 141.400 53.800 142.600 54.100 ;
        RECT 142.200 51.800 142.600 52.200 ;
        RECT 132.600 50.800 133.700 51.100 ;
        RECT 135.800 50.800 136.200 51.200 ;
        RECT 140.600 50.800 141.000 51.200 ;
        RECT 130.200 46.800 130.600 47.200 ;
        RECT 130.200 46.200 130.500 46.800 ;
        RECT 130.200 45.800 130.600 46.200 ;
        RECT 131.800 43.100 132.200 48.900 ;
        RECT 132.600 47.200 132.900 50.800 ;
        RECT 135.800 49.200 136.100 50.800 ;
        RECT 138.200 49.800 138.600 50.200 ;
        RECT 135.800 48.800 136.200 49.200 ;
        RECT 138.200 48.200 138.500 49.800 ;
        RECT 132.600 46.800 133.000 47.200 ;
        RECT 133.400 45.100 133.800 47.900 ;
        RECT 138.200 47.800 138.600 48.200 ;
        RECT 139.000 46.800 139.400 47.200 ;
        RECT 134.200 45.800 134.600 46.200 ;
        RECT 139.000 46.100 139.300 46.800 ;
        RECT 138.200 45.800 139.300 46.100 ;
        RECT 134.200 44.200 134.500 45.800 ;
        RECT 134.200 43.800 134.600 44.200 ;
        RECT 134.200 38.200 134.500 43.800 ;
        RECT 130.200 37.100 130.600 37.200 ;
        RECT 131.000 37.100 131.400 37.200 ;
        RECT 130.200 36.800 131.400 37.100 ;
        RECT 120.600 34.800 121.000 35.200 ;
        RECT 121.400 34.800 121.800 35.200 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 126.200 34.800 126.600 35.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 129.400 35.100 129.800 35.200 ;
        RECT 130.200 35.100 130.600 35.200 ;
        RECT 129.400 34.800 130.600 35.100 ;
        RECT 126.200 29.200 126.500 34.800 ;
        RECT 127.000 32.100 127.400 32.200 ;
        RECT 127.800 32.100 128.200 32.200 ;
        RECT 132.600 32.100 133.000 37.900 ;
        RECT 134.200 37.800 134.600 38.200 ;
        RECT 136.600 34.700 137.000 35.100 ;
        RECT 136.600 34.200 136.900 34.700 ;
        RECT 136.600 33.800 137.000 34.200 ;
        RECT 136.600 32.800 137.000 33.200 ;
        RECT 127.000 31.800 128.200 32.100 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 116.600 24.200 116.900 26.800 ;
        RECT 117.400 25.100 117.800 27.900 ;
        RECT 116.600 23.800 117.000 24.200 ;
        RECT 119.000 23.100 119.400 28.900 ;
        RECT 119.800 27.800 120.200 28.200 ;
        RECT 119.800 26.300 120.100 27.800 ;
        RECT 119.800 25.900 120.200 26.300 ;
        RECT 122.200 25.800 122.600 26.200 ;
        RECT 113.400 17.100 113.800 17.200 ;
        RECT 114.200 17.100 114.600 17.200 ;
        RECT 113.400 16.800 114.600 17.100 ;
        RECT 115.800 16.800 116.200 17.200 ;
        RECT 112.600 15.800 113.000 16.200 ;
        RECT 112.600 15.200 112.900 15.800 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 112.600 14.800 113.000 15.200 ;
        RECT 111.800 14.200 112.100 14.800 ;
        RECT 111.800 13.800 112.200 14.200 ;
        RECT 112.600 14.100 113.000 14.200 ;
        RECT 113.400 14.100 113.800 14.200 ;
        RECT 112.600 13.800 113.800 14.100 ;
        RECT 116.600 12.100 117.000 17.900 ;
        RECT 119.000 15.100 119.400 15.200 ;
        RECT 119.800 15.100 120.200 15.200 ;
        RECT 119.000 14.800 120.200 15.100 ;
        RECT 120.600 11.800 121.000 12.200 ;
        RECT 121.400 12.100 121.800 17.900 ;
        RECT 122.200 14.200 122.500 25.800 ;
        RECT 123.800 23.100 124.200 28.900 ;
        RECT 126.200 28.800 126.600 29.200 ;
        RECT 131.800 28.800 132.200 29.200 ;
        RECT 131.800 27.200 132.100 28.800 ;
        RECT 127.000 26.800 127.400 27.200 ;
        RECT 127.800 26.800 128.200 27.200 ;
        RECT 129.400 27.100 129.800 27.200 ;
        RECT 130.200 27.100 130.600 27.200 ;
        RECT 129.400 26.800 130.600 27.100 ;
        RECT 131.800 26.800 132.200 27.200 ;
        RECT 125.400 24.100 125.800 24.200 ;
        RECT 126.200 24.100 126.600 24.200 ;
        RECT 125.400 23.800 126.600 24.100 ;
        RECT 126.200 21.800 126.600 22.200 ;
        RECT 126.200 19.200 126.500 21.800 ;
        RECT 126.200 18.800 126.600 19.200 ;
        RECT 122.200 13.800 122.600 14.200 ;
        RECT 122.200 12.200 122.500 13.800 ;
        RECT 123.000 13.100 123.400 15.900 ;
        RECT 123.800 14.800 124.200 15.200 ;
        RECT 124.600 14.800 125.000 15.200 ;
        RECT 123.800 14.200 124.100 14.800 ;
        RECT 123.800 13.800 124.200 14.200 ;
        RECT 124.600 13.200 124.900 14.800 ;
        RECT 124.600 12.800 125.000 13.200 ;
        RECT 122.200 11.800 122.600 12.200 ;
        RECT 119.800 10.800 120.200 11.200 ;
        RECT 100.600 6.800 101.000 7.200 ;
        RECT 103.800 6.800 104.200 7.200 ;
        RECT 107.000 6.800 107.400 7.200 ;
        RECT 107.800 6.800 108.200 7.200 ;
        RECT 111.000 6.800 111.400 7.200 ;
        RECT 114.200 6.800 114.600 7.200 ;
        RECT 103.800 6.200 104.100 6.800 ;
        RECT 103.800 5.800 104.200 6.200 ;
        RECT 106.200 6.100 106.600 6.200 ;
        RECT 107.000 6.100 107.400 6.200 ;
        RECT 106.200 5.800 107.400 6.100 ;
        RECT 106.200 5.200 106.500 5.800 ;
        RECT 103.800 5.100 104.200 5.200 ;
        RECT 104.600 5.100 105.000 5.200 ;
        RECT 103.800 4.800 105.000 5.100 ;
        RECT 106.200 4.800 106.600 5.200 ;
        RECT 111.000 3.200 111.300 6.800 ;
        RECT 114.200 6.200 114.500 6.800 ;
        RECT 114.200 5.800 114.600 6.200 ;
        RECT 115.000 5.100 115.400 7.900 ;
        RECT 115.800 6.800 116.200 7.200 ;
        RECT 115.800 6.200 116.100 6.800 ;
        RECT 115.800 5.800 116.200 6.200 ;
        RECT 111.000 2.800 111.400 3.200 ;
        RECT 116.600 3.100 117.000 8.900 ;
        RECT 119.800 7.200 120.100 10.800 ;
        RECT 120.600 8.200 120.900 11.800 ;
        RECT 127.000 9.200 127.300 26.800 ;
        RECT 127.800 26.200 128.100 26.800 ;
        RECT 127.800 25.800 128.200 26.200 ;
        RECT 130.200 25.800 130.600 26.200 ;
        RECT 130.200 25.200 130.500 25.800 ;
        RECT 130.200 24.800 130.600 25.200 ;
        RECT 132.600 25.100 133.000 27.900 ;
        RECT 133.400 26.800 133.800 27.200 ;
        RECT 128.600 17.800 129.000 18.200 ;
        RECT 128.600 17.200 128.900 17.800 ;
        RECT 128.600 17.100 129.000 17.200 ;
        RECT 129.400 17.100 129.800 17.200 ;
        RECT 128.600 16.800 129.800 17.100 ;
        RECT 127.800 14.800 128.200 15.200 ;
        RECT 127.800 13.200 128.100 14.800 ;
        RECT 127.800 12.800 128.200 13.200 ;
        RECT 131.000 12.100 131.400 17.900 ;
        RECT 132.600 13.800 133.000 14.200 ;
        RECT 132.600 12.200 132.900 13.800 ;
        RECT 132.600 11.800 133.000 12.200 ;
        RECT 128.600 9.800 129.000 10.200 ;
        RECT 120.600 7.800 121.000 8.200 ;
        RECT 118.200 6.800 118.600 7.200 ;
        RECT 119.800 6.800 120.200 7.200 ;
        RECT 118.200 6.200 118.500 6.800 ;
        RECT 118.200 5.800 118.600 6.200 ;
        RECT 121.400 3.100 121.800 8.900 ;
        RECT 127.000 8.800 127.400 9.200 ;
        RECT 126.200 7.100 126.600 7.200 ;
        RECT 127.000 7.100 127.400 7.200 ;
        RECT 126.200 6.800 127.400 7.100 ;
        RECT 128.600 6.200 128.900 9.800 ;
        RECT 129.400 8.800 129.800 9.200 ;
        RECT 129.400 7.200 129.700 8.800 ;
        RECT 129.400 6.800 129.800 7.200 ;
        RECT 126.200 5.800 126.600 6.200 ;
        RECT 128.600 5.800 129.000 6.200 ;
        RECT 126.200 5.200 126.500 5.800 ;
        RECT 126.200 4.800 126.600 5.200 ;
        RECT 130.200 5.100 130.600 7.900 ;
        RECT 131.800 3.100 132.200 8.900 ;
        RECT 132.600 8.200 132.900 11.800 ;
        RECT 133.400 11.200 133.700 26.800 ;
        RECT 134.200 23.100 134.600 28.900 ;
        RECT 135.000 26.800 135.400 27.200 ;
        RECT 135.000 26.300 135.300 26.800 ;
        RECT 135.000 25.900 135.400 26.300 ;
        RECT 134.200 14.800 134.600 15.200 ;
        RECT 134.200 14.200 134.500 14.800 ;
        RECT 134.200 13.800 134.600 14.200 ;
        RECT 135.800 12.100 136.200 17.900 ;
        RECT 136.600 14.200 136.900 32.800 ;
        RECT 137.400 32.100 137.800 37.900 ;
        RECT 138.200 34.200 138.500 45.800 ;
        RECT 139.800 45.100 140.200 47.900 ;
        RECT 141.400 43.100 141.800 48.900 ;
        RECT 142.200 46.300 142.500 51.800 ;
        RECT 142.200 45.900 142.600 46.300 ;
        RECT 143.000 39.200 143.300 63.800 ;
        RECT 143.800 55.200 144.100 69.800 ;
        RECT 144.600 67.200 144.900 85.800 ;
        RECT 147.800 83.100 148.200 88.900 ;
        RECT 151.800 88.200 152.100 105.800 ;
        RECT 153.400 95.200 153.700 106.800 ;
        RECT 154.200 106.200 154.500 115.800 ;
        RECT 155.000 114.700 155.400 115.100 ;
        RECT 155.000 112.200 155.300 114.700 ;
        RECT 155.000 111.800 155.400 112.200 ;
        RECT 155.800 112.100 156.200 117.900 ;
        RECT 158.200 116.800 158.600 117.200 ;
        RECT 158.200 116.200 158.500 116.800 ;
        RECT 156.600 114.800 157.000 115.200 ;
        RECT 156.600 114.200 156.900 114.800 ;
        RECT 156.600 113.800 157.000 114.200 ;
        RECT 157.400 113.100 157.800 115.900 ;
        RECT 158.200 115.800 158.600 116.200 ;
        RECT 159.800 115.100 160.200 115.200 ;
        RECT 159.000 114.800 160.200 115.100 ;
        RECT 157.400 112.100 157.800 112.200 ;
        RECT 158.200 112.100 158.600 112.200 ;
        RECT 157.400 111.800 158.600 112.100 ;
        RECT 154.200 105.800 154.600 106.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 157.400 105.800 157.800 106.200 ;
        RECT 155.800 104.800 156.200 105.200 ;
        RECT 155.000 100.800 155.400 101.200 ;
        RECT 155.000 99.200 155.300 100.800 ;
        RECT 155.000 98.800 155.400 99.200 ;
        RECT 153.400 94.800 153.800 95.200 ;
        RECT 155.800 94.200 156.100 104.800 ;
        RECT 156.600 103.200 156.900 105.800 ;
        RECT 157.400 104.200 157.700 105.800 ;
        RECT 159.000 105.200 159.300 114.800 ;
        RECT 159.800 114.100 160.200 114.200 ;
        RECT 160.600 114.100 161.000 114.200 ;
        RECT 159.800 113.800 161.000 114.100 ;
        RECT 161.400 113.100 161.800 115.900 ;
        RECT 162.200 114.800 162.600 115.200 ;
        RECT 162.200 114.200 162.500 114.800 ;
        RECT 162.200 113.800 162.600 114.200 ;
        RECT 161.400 111.800 161.800 112.200 ;
        RECT 163.000 112.100 163.400 117.900 ;
        RECT 164.600 116.800 165.000 117.200 ;
        RECT 164.600 115.200 164.900 116.800 ;
        RECT 164.600 114.800 165.000 115.200 ;
        RECT 164.600 111.800 165.000 112.200 ;
        RECT 161.400 106.200 161.700 111.800 ;
        RECT 163.800 109.800 164.200 110.200 ;
        RECT 163.800 107.200 164.100 109.800 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 164.600 106.200 164.900 111.800 ;
        RECT 165.400 111.200 165.700 125.800 ;
        RECT 166.200 124.200 166.500 125.800 ;
        RECT 168.600 124.200 168.900 125.800 ;
        RECT 166.200 123.800 166.600 124.200 ;
        RECT 168.600 123.800 169.000 124.200 ;
        RECT 167.000 121.800 167.400 122.200 ;
        RECT 167.000 112.200 167.300 121.800 ;
        RECT 167.000 111.800 167.400 112.200 ;
        RECT 167.800 112.100 168.200 117.900 ;
        RECT 165.400 110.800 165.800 111.200 ;
        RECT 167.000 106.800 167.400 107.200 ;
        RECT 159.800 105.800 160.200 106.200 ;
        RECT 161.400 105.800 161.800 106.200 ;
        RECT 164.600 105.800 165.000 106.200 ;
        RECT 159.000 104.800 159.400 105.200 ;
        RECT 157.400 103.800 157.800 104.200 ;
        RECT 156.600 102.800 157.000 103.200 ;
        RECT 156.600 97.200 156.900 102.800 ;
        RECT 159.800 101.200 160.100 105.800 ;
        RECT 159.800 100.800 160.200 101.200 ;
        RECT 156.600 96.800 157.000 97.200 ;
        RECT 157.400 95.800 157.800 96.200 ;
        RECT 157.400 95.200 157.700 95.800 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 158.200 94.800 158.600 95.200 ;
        RECT 155.800 93.800 156.200 94.200 ;
        RECT 148.600 87.800 149.000 88.200 ;
        RECT 148.600 87.200 148.900 87.800 ;
        RECT 148.600 86.800 149.000 87.200 ;
        RECT 149.400 85.100 149.800 87.900 ;
        RECT 151.800 87.800 152.200 88.200 ;
        RECT 150.200 87.100 150.600 87.200 ;
        RECT 151.000 87.100 151.400 87.200 ;
        RECT 150.200 86.800 151.400 87.100 ;
        RECT 147.800 77.100 148.200 77.200 ;
        RECT 148.600 77.100 149.000 77.200 ;
        RECT 147.800 76.800 149.000 77.100 ;
        RECT 147.000 73.800 147.400 74.200 ;
        RECT 144.600 66.800 145.000 67.200 ;
        RECT 144.600 66.200 144.900 66.800 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 143.800 54.800 144.200 55.200 ;
        RECT 143.800 54.200 144.100 54.800 ;
        RECT 143.800 53.800 144.200 54.200 ;
        RECT 144.600 46.200 144.900 65.800 ;
        RECT 146.200 63.100 146.600 68.900 ;
        RECT 146.200 60.800 146.600 61.200 ;
        RECT 146.200 55.200 146.500 60.800 ;
        RECT 146.200 54.800 146.600 55.200 ;
        RECT 145.400 53.800 145.800 54.200 ;
        RECT 146.200 53.800 146.600 54.200 ;
        RECT 145.400 53.200 145.700 53.800 ;
        RECT 146.200 53.200 146.500 53.800 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 146.200 52.800 146.600 53.200 ;
        RECT 144.600 45.800 145.000 46.200 ;
        RECT 146.200 43.100 146.600 48.900 ;
        RECT 146.200 40.800 146.600 41.200 ;
        RECT 146.200 39.200 146.500 40.800 ;
        RECT 141.400 38.800 141.800 39.200 ;
        RECT 143.000 38.800 143.400 39.200 ;
        RECT 143.800 38.800 144.200 39.200 ;
        RECT 146.200 38.800 146.600 39.200 ;
        RECT 139.800 36.800 140.200 37.200 ;
        RECT 138.200 33.800 138.600 34.200 ;
        RECT 139.000 33.100 139.400 35.900 ;
        RECT 139.800 34.200 140.100 36.800 ;
        RECT 141.400 36.200 141.700 38.800 ;
        RECT 141.400 35.800 141.800 36.200 ;
        RECT 139.800 33.800 140.200 34.200 ;
        RECT 141.400 33.800 141.800 34.200 ;
        RECT 140.600 31.800 141.000 32.200 ;
        RECT 141.400 32.100 141.700 33.800 ;
        RECT 141.400 31.800 142.500 32.100 ;
        RECT 140.600 30.200 140.900 31.800 ;
        RECT 140.600 29.800 141.000 30.200 ;
        RECT 142.200 29.200 142.500 31.800 ;
        RECT 140.600 29.100 141.000 29.200 ;
        RECT 141.400 29.100 141.800 29.200 ;
        RECT 139.000 23.100 139.400 28.900 ;
        RECT 140.600 28.800 141.800 29.100 ;
        RECT 142.200 28.800 142.600 29.200 ;
        RECT 142.200 26.800 142.600 27.200 ;
        RECT 142.200 25.200 142.500 26.800 ;
        RECT 143.800 26.200 144.100 38.800 ;
        RECT 147.000 36.200 147.300 73.800 ;
        RECT 150.200 72.100 150.600 77.900 ;
        RECT 151.800 75.200 152.100 87.800 ;
        RECT 153.400 86.800 153.800 87.200 ;
        RECT 153.400 86.200 153.700 86.800 ;
        RECT 153.400 85.800 153.800 86.200 ;
        RECT 155.800 85.800 156.200 86.200 ;
        RECT 155.800 85.200 156.100 85.800 ;
        RECT 152.600 85.100 153.000 85.200 ;
        RECT 153.400 85.100 153.800 85.200 ;
        RECT 152.600 84.800 153.800 85.100 ;
        RECT 155.800 84.800 156.200 85.200 ;
        RECT 156.600 80.200 156.900 94.800 ;
        RECT 158.200 89.200 158.500 94.800 ;
        RECT 159.800 92.800 160.200 93.200 ;
        RECT 159.000 91.800 159.400 92.200 ;
        RECT 159.000 91.200 159.300 91.800 ;
        RECT 159.000 90.800 159.400 91.200 ;
        RECT 159.800 91.100 160.100 92.800 ;
        RECT 159.800 90.800 160.900 91.100 ;
        RECT 158.200 88.800 158.600 89.200 ;
        RECT 159.000 89.100 159.400 89.200 ;
        RECT 159.800 89.100 160.200 89.200 ;
        RECT 159.000 88.800 160.200 89.100 ;
        RECT 158.200 87.200 158.500 88.800 ;
        RECT 159.000 88.100 159.400 88.200 ;
        RECT 159.800 88.100 160.200 88.200 ;
        RECT 159.000 87.800 160.200 88.100 ;
        RECT 158.200 86.800 158.600 87.200 ;
        RECT 160.600 86.200 160.900 90.800 ;
        RECT 157.400 86.100 157.800 86.200 ;
        RECT 158.200 86.100 158.600 86.200 ;
        RECT 157.400 85.800 158.600 86.100 ;
        RECT 160.600 85.800 161.000 86.200 ;
        RECT 161.400 85.200 161.700 105.800 ;
        RECT 162.200 104.800 162.600 105.200 ;
        RECT 165.400 104.800 165.800 105.200 ;
        RECT 162.200 104.200 162.500 104.800 ;
        RECT 165.400 104.200 165.700 104.800 ;
        RECT 167.000 104.200 167.300 106.800 ;
        RECT 168.600 106.100 169.000 106.200 ;
        RECT 169.400 106.100 169.700 130.800 ;
        RECT 173.400 127.200 173.700 145.800 ;
        RECT 177.400 143.100 177.800 148.900 ;
        RECT 176.600 135.800 177.000 136.200 ;
        RECT 176.600 135.200 176.900 135.800 ;
        RECT 174.200 134.800 174.600 135.200 ;
        RECT 175.800 134.800 176.200 135.200 ;
        RECT 176.600 134.800 177.000 135.200 ;
        RECT 174.200 128.200 174.500 134.800 ;
        RECT 175.800 134.200 176.100 134.800 ;
        RECT 175.000 133.800 175.400 134.200 ;
        RECT 175.800 133.800 176.200 134.200 ;
        RECT 175.000 130.200 175.300 133.800 ;
        RECT 175.000 129.800 175.400 130.200 ;
        RECT 175.000 128.800 175.400 129.200 ;
        RECT 174.200 127.800 174.600 128.200 ;
        RECT 175.000 127.200 175.300 128.800 ;
        RECT 170.200 126.800 170.600 127.200 ;
        RECT 172.600 126.800 173.000 127.200 ;
        RECT 173.400 126.800 173.800 127.200 ;
        RECT 175.000 126.800 175.400 127.200 ;
        RECT 170.200 114.200 170.500 126.800 ;
        RECT 171.000 125.800 171.400 126.200 ;
        RECT 171.000 123.200 171.300 125.800 ;
        RECT 172.600 125.200 172.900 126.800 ;
        RECT 172.600 124.800 173.000 125.200 ;
        RECT 173.400 124.800 173.800 125.200 ;
        RECT 175.800 125.100 176.200 127.900 ;
        RECT 173.400 123.200 173.700 124.800 ;
        RECT 171.000 122.800 171.400 123.200 ;
        RECT 173.400 122.800 173.800 123.200 ;
        RECT 177.400 123.100 177.800 128.900 ;
        RECT 178.200 128.200 178.500 149.800 ;
        RECT 183.800 149.100 184.100 173.800 ;
        RECT 184.600 173.100 185.000 175.900 ;
        RECT 185.400 175.200 185.700 185.800 ;
        RECT 186.200 184.200 186.500 185.800 ;
        RECT 189.400 184.200 189.700 185.800 ;
        RECT 186.200 183.800 186.600 184.200 ;
        RECT 189.400 183.800 189.800 184.200 ;
        RECT 191.800 183.800 192.200 184.200 ;
        RECT 185.400 174.800 185.800 175.200 ;
        RECT 185.400 163.100 185.800 168.900 ;
        RECT 185.400 152.100 185.800 157.900 ;
        RECT 186.200 151.200 186.500 183.800 ;
        RECT 188.600 173.100 189.000 175.900 ;
        RECT 187.000 171.800 187.400 172.200 ;
        RECT 190.200 172.100 190.600 177.900 ;
        RECT 191.800 175.200 192.100 183.800 ;
        RECT 192.600 183.100 193.000 188.900 ;
        RECT 195.800 186.800 196.200 187.200 ;
        RECT 195.800 186.200 196.100 186.800 ;
        RECT 195.800 185.800 196.200 186.200 ;
        RECT 197.400 183.100 197.800 188.900 ;
        RECT 199.800 188.800 200.200 189.200 ;
        RECT 200.600 188.800 201.000 189.200 ;
        RECT 203.000 188.800 203.400 189.200 ;
        RECT 198.200 186.800 198.600 187.200 ;
        RECT 198.200 186.200 198.500 186.800 ;
        RECT 198.200 185.800 198.600 186.200 ;
        RECT 199.000 185.100 199.400 187.900 ;
        RECT 203.000 187.200 203.300 188.800 ;
        RECT 203.000 186.800 203.400 187.200 ;
        RECT 199.800 185.800 200.200 186.200 ;
        RECT 199.800 185.200 200.100 185.800 ;
        RECT 199.800 184.800 200.200 185.200 ;
        RECT 199.800 183.800 200.200 184.200 ;
        RECT 199.000 180.800 199.400 181.200 ;
        RECT 191.800 174.800 192.200 175.200 ;
        RECT 192.600 174.800 193.000 175.200 ;
        RECT 191.800 174.200 192.100 174.800 ;
        RECT 191.800 173.800 192.200 174.200 ;
        RECT 187.000 170.200 187.300 171.800 ;
        RECT 192.600 170.200 192.900 174.800 ;
        RECT 195.000 172.100 195.400 177.900 ;
        RECT 199.000 175.200 199.300 180.800 ;
        RECT 199.800 179.200 200.100 183.800 ;
        RECT 206.200 183.100 206.600 188.900 ;
        RECT 207.000 187.800 207.400 188.200 ;
        RECT 207.000 187.200 207.300 187.800 ;
        RECT 207.000 186.800 207.400 187.200 ;
        RECT 207.800 186.200 208.100 195.800 ;
        RECT 208.600 195.200 208.900 195.800 ;
        RECT 208.600 194.800 209.000 195.200 ;
        RECT 209.400 194.200 209.700 196.800 ;
        RECT 208.600 193.800 209.000 194.200 ;
        RECT 209.400 193.800 209.800 194.200 ;
        RECT 207.800 185.800 208.200 186.200 ;
        RECT 199.800 178.800 200.200 179.200 ;
        RECT 206.200 175.800 206.600 176.200 ;
        RECT 198.200 174.800 198.600 175.200 ;
        RECT 199.000 174.800 199.400 175.200 ;
        RECT 201.400 175.100 201.800 175.200 ;
        RECT 200.600 174.800 201.800 175.100 ;
        RECT 203.800 175.100 204.200 175.200 ;
        RECT 204.600 175.100 205.000 175.200 ;
        RECT 206.200 175.100 206.500 175.800 ;
        RECT 203.800 174.800 205.000 175.100 ;
        RECT 205.400 174.800 206.500 175.100 ;
        RECT 207.800 174.800 208.200 175.200 ;
        RECT 198.200 174.200 198.500 174.800 ;
        RECT 198.200 173.800 198.600 174.200 ;
        RECT 197.400 171.800 197.800 172.200 ;
        RECT 187.000 169.800 187.400 170.200 ;
        RECT 192.600 169.800 193.000 170.200 ;
        RECT 195.000 169.800 195.400 170.200 ;
        RECT 187.000 168.200 187.300 169.800 ;
        RECT 195.000 169.200 195.300 169.800 ;
        RECT 187.000 167.800 187.400 168.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 187.000 165.200 187.300 165.800 ;
        RECT 187.000 164.800 187.400 165.200 ;
        RECT 189.400 158.200 189.700 166.800 ;
        RECT 190.200 163.100 190.600 168.900 ;
        RECT 195.000 168.800 195.400 169.200 ;
        RECT 191.800 165.100 192.200 167.900 ;
        RECT 192.600 167.800 193.000 168.200 ;
        RECT 192.600 167.200 192.900 167.800 ;
        RECT 197.400 167.200 197.700 171.800 ;
        RECT 200.600 169.200 200.900 174.800 ;
        RECT 205.400 174.200 205.700 174.800 ;
        RECT 203.800 173.800 204.200 174.200 ;
        RECT 205.400 173.800 205.800 174.200 ;
        RECT 206.200 174.100 206.600 174.200 ;
        RECT 207.000 174.100 207.400 174.200 ;
        RECT 206.200 173.800 207.400 174.100 ;
        RECT 200.600 168.800 201.000 169.200 ;
        RECT 192.600 166.800 193.000 167.200 ;
        RECT 197.400 167.100 197.800 167.200 ;
        RECT 197.400 166.800 199.300 167.100 ;
        RECT 199.000 166.200 199.300 166.800 ;
        RECT 192.600 166.100 193.000 166.200 ;
        RECT 193.400 166.100 193.800 166.200 ;
        RECT 192.600 165.800 193.800 166.100 ;
        RECT 195.800 165.800 196.200 166.200 ;
        RECT 198.200 165.800 198.600 166.200 ;
        RECT 199.000 165.800 199.400 166.200 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 195.800 165.200 196.100 165.800 ;
        RECT 195.800 164.800 196.200 165.200 ;
        RECT 198.200 161.200 198.500 165.800 ;
        RECT 198.200 160.800 198.600 161.200 ;
        RECT 198.200 159.800 198.600 160.200 ;
        RECT 189.400 157.800 189.800 158.200 ;
        RECT 187.800 155.100 188.200 155.200 ;
        RECT 188.600 155.100 189.000 155.200 ;
        RECT 187.800 154.800 189.000 155.100 ;
        RECT 189.400 154.200 189.700 157.800 ;
        RECT 189.400 153.800 189.800 154.200 ;
        RECT 190.200 152.100 190.600 157.900 ;
        RECT 191.800 153.100 192.200 155.900 ;
        RECT 192.600 155.800 193.000 156.200 ;
        RECT 194.200 155.800 194.600 156.200 ;
        RECT 195.800 155.800 196.200 156.200 ;
        RECT 192.600 154.200 192.900 155.800 ;
        RECT 194.200 155.200 194.500 155.800 ;
        RECT 195.800 155.200 196.100 155.800 ;
        RECT 194.200 154.800 194.600 155.200 ;
        RECT 195.800 154.800 196.200 155.200 ;
        RECT 196.600 154.800 197.000 155.200 ;
        RECT 192.600 153.800 193.000 154.200 ;
        RECT 186.200 150.800 186.600 151.200 ;
        RECT 190.200 150.800 190.600 151.200 ;
        RECT 179.000 147.100 179.400 147.200 ;
        RECT 179.800 147.100 180.200 147.200 ;
        RECT 179.000 146.800 180.200 147.100 ;
        RECT 179.000 146.100 179.400 146.200 ;
        RECT 179.800 146.100 180.200 146.200 ;
        RECT 179.000 145.800 180.200 146.100 ;
        RECT 182.200 143.100 182.600 148.900 ;
        RECT 183.000 148.800 184.100 149.100 ;
        RECT 183.000 147.200 183.300 148.800 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 183.800 145.100 184.200 147.900 ;
        RECT 184.600 142.100 185.000 142.200 ;
        RECT 185.400 142.100 185.800 142.200 ;
        RECT 184.600 141.800 185.800 142.100 ;
        RECT 183.800 140.800 184.200 141.200 ;
        RECT 182.200 135.800 182.600 136.200 ;
        RECT 182.200 135.200 182.500 135.800 ;
        RECT 183.800 135.200 184.100 140.800 ;
        RECT 184.600 136.800 185.000 137.200 ;
        RECT 184.600 136.200 184.900 136.800 ;
        RECT 184.600 135.800 185.000 136.200 ;
        RECT 179.000 135.100 179.400 135.200 ;
        RECT 179.800 135.100 180.200 135.200 ;
        RECT 179.000 134.800 180.200 135.100 ;
        RECT 180.600 134.800 181.000 135.200 ;
        RECT 182.200 134.800 182.600 135.200 ;
        RECT 183.800 134.800 184.200 135.200 ;
        RECT 187.000 134.800 187.400 135.200 ;
        RECT 189.400 134.800 189.800 135.200 ;
        RECT 180.600 132.200 180.900 134.800 ;
        RECT 183.000 133.800 183.400 134.200 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 183.000 133.200 183.300 133.800 ;
        RECT 183.000 132.800 183.400 133.200 ;
        RECT 180.600 131.800 181.000 132.200 ;
        RECT 184.600 131.800 185.000 132.200 ;
        RECT 184.600 131.200 184.900 131.800 ;
        RECT 186.200 131.200 186.500 133.800 ;
        RECT 184.600 130.800 185.000 131.200 ;
        RECT 186.200 130.800 186.600 131.200 ;
        RECT 183.800 129.100 184.200 129.200 ;
        RECT 184.600 129.100 185.000 129.200 ;
        RECT 178.200 127.800 178.600 128.200 ;
        RECT 178.200 125.900 178.600 126.300 ;
        RECT 178.200 125.200 178.500 125.900 ;
        RECT 181.400 125.800 181.800 126.200 ;
        RECT 178.200 124.800 178.600 125.200 ;
        RECT 178.200 123.800 178.600 124.200 ;
        RECT 178.200 119.200 178.500 123.800 ;
        RECT 181.400 122.200 181.700 125.800 ;
        RECT 182.200 123.100 182.600 128.900 ;
        RECT 183.800 128.800 185.000 129.100 ;
        RECT 186.200 128.800 186.600 129.200 ;
        RECT 186.200 126.200 186.500 128.800 ;
        RECT 185.400 125.800 185.800 126.200 ;
        RECT 186.200 125.800 186.600 126.200 ;
        RECT 185.400 125.200 185.700 125.800 ;
        RECT 185.400 124.800 185.800 125.200 ;
        RECT 181.400 121.800 181.800 122.200 ;
        RECT 183.000 121.800 183.400 122.200 ;
        RECT 178.200 118.800 178.600 119.200 ;
        RECT 171.800 117.100 172.200 117.200 ;
        RECT 172.600 117.100 173.000 117.200 ;
        RECT 171.800 116.800 173.000 117.100 ;
        RECT 173.400 116.800 173.800 117.200 ;
        RECT 171.800 115.800 172.200 116.200 ;
        RECT 171.800 115.200 172.100 115.800 ;
        RECT 171.800 114.800 172.200 115.200 ;
        RECT 170.200 113.800 170.600 114.200 ;
        RECT 171.000 114.100 171.400 114.200 ;
        RECT 171.800 114.100 172.200 114.200 ;
        RECT 171.000 113.800 172.200 114.100 ;
        RECT 170.200 112.100 170.600 112.200 ;
        RECT 171.000 112.100 171.400 112.200 ;
        RECT 170.200 111.800 171.400 112.100 ;
        RECT 171.000 109.800 171.400 110.200 ;
        RECT 171.000 108.200 171.300 109.800 ;
        RECT 171.000 107.800 171.400 108.200 ;
        RECT 168.600 105.800 169.700 106.100 ;
        RECT 171.000 106.800 171.400 107.200 ;
        RECT 172.600 106.800 173.000 107.200 ;
        RECT 171.000 105.200 171.300 106.800 ;
        RECT 172.600 105.200 172.900 106.800 ;
        RECT 169.400 105.100 169.800 105.200 ;
        RECT 170.200 105.100 170.600 105.200 ;
        RECT 169.400 104.800 170.600 105.100 ;
        RECT 171.000 104.800 171.400 105.200 ;
        RECT 172.600 104.800 173.000 105.200 ;
        RECT 162.200 103.800 162.600 104.200 ;
        RECT 165.400 103.800 165.800 104.200 ;
        RECT 167.000 103.800 167.400 104.200 ;
        RECT 170.200 100.200 170.500 104.800 ;
        RECT 171.000 103.100 171.400 103.200 ;
        RECT 171.800 103.100 172.200 103.200 ;
        RECT 171.000 102.800 172.200 103.100 ;
        RECT 170.200 99.800 170.600 100.200 ;
        RECT 173.400 99.200 173.700 116.800 ;
        RECT 174.200 116.100 174.600 116.200 ;
        RECT 175.000 116.100 175.400 116.200 ;
        RECT 174.200 115.800 175.400 116.100 ;
        RECT 177.400 115.800 177.800 116.200 ;
        RECT 177.400 115.200 177.700 115.800 ;
        RECT 175.800 114.800 176.200 115.200 ;
        RECT 176.600 114.800 177.000 115.200 ;
        RECT 177.400 114.800 177.800 115.200 ;
        RECT 181.400 114.800 181.800 115.200 ;
        RECT 182.200 114.800 182.600 115.200 ;
        RECT 175.800 114.200 176.100 114.800 ;
        RECT 175.800 113.800 176.200 114.200 ;
        RECT 175.800 112.200 176.100 113.800 ;
        RECT 175.800 111.800 176.200 112.200 ;
        RECT 176.600 102.200 176.900 114.800 ;
        RECT 181.400 112.200 181.700 114.800 ;
        RECT 182.200 114.200 182.500 114.800 ;
        RECT 182.200 113.800 182.600 114.200 ;
        RECT 181.400 111.800 181.800 112.200 ;
        RECT 182.200 110.800 182.600 111.200 ;
        RECT 177.400 105.100 177.800 105.200 ;
        RECT 178.200 105.100 178.600 105.200 ;
        RECT 177.400 104.800 178.600 105.100 ;
        RECT 179.000 103.100 179.400 108.900 ;
        RECT 182.200 107.200 182.500 110.800 ;
        RECT 182.200 106.800 182.600 107.200 ;
        RECT 181.400 105.800 181.800 106.200 ;
        RECT 181.400 103.200 181.700 105.800 ;
        RECT 181.400 102.800 181.800 103.200 ;
        RECT 176.600 101.800 177.000 102.200 ;
        RECT 181.400 99.800 181.800 100.200 ;
        RECT 173.400 98.800 173.800 99.200 ;
        RECT 179.000 99.100 179.400 99.200 ;
        RECT 179.800 99.100 180.200 99.200 ;
        RECT 179.000 98.800 180.200 99.100 ;
        RECT 163.000 92.100 163.400 97.900 ;
        RECT 164.600 94.800 165.000 95.200 ;
        RECT 164.600 89.200 164.900 94.800 ;
        RECT 167.800 92.100 168.200 97.900 ;
        RECT 169.400 93.100 169.800 95.900 ;
        RECT 170.200 93.100 170.600 95.900 ;
        RECT 171.800 92.100 172.200 97.900 ;
        RECT 173.400 95.800 173.800 96.200 ;
        RECT 173.400 95.200 173.700 95.800 ;
        RECT 173.400 94.800 173.800 95.200 ;
        RECT 175.000 95.100 175.400 95.200 ;
        RECT 175.800 95.100 176.200 95.200 ;
        RECT 175.000 94.800 176.200 95.100 ;
        RECT 166.200 89.800 166.600 90.200 ;
        RECT 164.600 88.800 165.000 89.200 ;
        RECT 165.400 88.800 165.800 89.200 ;
        RECT 165.400 88.200 165.700 88.800 ;
        RECT 165.400 87.800 165.800 88.200 ;
        RECT 165.400 87.200 165.700 87.800 ;
        RECT 163.800 86.800 164.200 87.200 ;
        RECT 165.400 86.800 165.800 87.200 ;
        RECT 163.800 86.200 164.100 86.800 ;
        RECT 163.800 85.800 164.200 86.200 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 161.400 84.800 161.800 85.200 ;
        RECT 163.800 82.800 164.200 83.200 ;
        RECT 163.000 81.800 163.400 82.200 ;
        RECT 163.000 81.200 163.300 81.800 ;
        RECT 163.000 80.800 163.400 81.200 ;
        RECT 156.600 79.800 157.000 80.200 ;
        RECT 163.800 79.200 164.100 82.800 ;
        RECT 163.800 78.800 164.200 79.200 ;
        RECT 151.800 74.800 152.200 75.200 ;
        RECT 153.400 75.000 153.800 75.100 ;
        RECT 154.200 75.000 154.600 75.100 ;
        RECT 153.400 74.700 154.600 75.000 ;
        RECT 155.000 72.100 155.400 77.900 ;
        RECT 164.600 77.200 164.900 85.800 ;
        RECT 166.200 77.200 166.500 89.800 ;
        RECT 170.200 89.100 170.600 89.200 ;
        RECT 171.000 89.100 171.400 89.200 ;
        RECT 170.200 88.800 171.400 89.100 ;
        RECT 167.800 87.100 168.200 87.200 ;
        RECT 168.600 87.100 169.000 87.200 ;
        RECT 167.800 86.800 169.000 87.100 ;
        RECT 169.400 86.800 169.800 87.200 ;
        RECT 170.200 87.100 170.600 87.200 ;
        RECT 170.200 86.800 171.300 87.100 ;
        RECT 167.000 85.800 167.400 86.200 ;
        RECT 167.000 85.200 167.300 85.800 ;
        RECT 169.400 85.200 169.700 86.800 ;
        RECT 171.000 86.200 171.300 86.800 ;
        RECT 170.200 85.800 170.600 86.200 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 167.000 84.800 167.400 85.200 ;
        RECT 169.400 84.800 169.800 85.200 ;
        RECT 167.000 78.200 167.300 84.800 ;
        RECT 170.200 78.200 170.500 85.800 ;
        RECT 173.400 83.100 173.800 88.900 ;
        RECT 175.800 87.200 176.100 94.800 ;
        RECT 176.600 92.100 177.000 97.900 ;
        RECT 179.800 92.800 180.200 93.200 ;
        RECT 179.800 92.200 180.100 92.800 ;
        RECT 179.800 91.800 180.200 92.200 ;
        RECT 177.400 90.800 177.800 91.200 ;
        RECT 175.800 86.800 176.200 87.200 ;
        RECT 175.800 86.100 176.200 86.200 ;
        RECT 176.600 86.100 177.000 86.200 ;
        RECT 175.800 85.800 177.000 86.100 ;
        RECT 167.000 77.800 167.400 78.200 ;
        RECT 170.200 77.800 170.600 78.200 ;
        RECT 157.400 77.100 157.800 77.200 ;
        RECT 158.200 77.100 158.600 77.200 ;
        RECT 157.400 76.800 158.600 77.100 ;
        RECT 164.600 76.800 165.000 77.200 ;
        RECT 166.200 76.800 166.600 77.200 ;
        RECT 169.400 76.800 169.800 77.200 ;
        RECT 156.600 73.100 157.000 75.900 ;
        RECT 166.200 75.200 166.500 76.800 ;
        RECT 169.400 76.200 169.700 76.800 ;
        RECT 167.800 75.800 168.200 76.200 ;
        RECT 169.400 75.800 169.800 76.200 ;
        RECT 167.800 75.200 168.100 75.800 ;
        RECT 160.600 75.100 161.000 75.200 ;
        RECT 161.400 75.100 161.800 75.200 ;
        RECT 160.600 74.800 161.800 75.100 ;
        RECT 162.200 74.800 162.600 75.200 ;
        RECT 166.200 74.800 166.600 75.200 ;
        RECT 167.800 74.800 168.200 75.200 ;
        RECT 157.400 73.800 157.800 74.200 ;
        RECT 160.600 74.100 161.000 74.200 ;
        RECT 161.400 74.100 161.800 74.200 ;
        RECT 160.600 73.800 161.800 74.100 ;
        RECT 157.400 72.200 157.700 73.800 ;
        RECT 162.200 73.200 162.500 74.800 ;
        RECT 170.200 74.200 170.500 77.800 ;
        RECT 171.000 74.800 171.400 75.200 ;
        RECT 171.000 74.200 171.300 74.800 ;
        RECT 166.200 74.100 166.600 74.200 ;
        RECT 167.000 74.100 167.400 74.200 ;
        RECT 166.200 73.800 167.400 74.100 ;
        RECT 170.200 73.800 170.600 74.200 ;
        RECT 171.000 73.800 171.400 74.200 ;
        RECT 162.200 72.800 162.600 73.200 ;
        RECT 157.400 71.800 157.800 72.200 ;
        RECT 162.200 72.100 162.500 72.800 ;
        RECT 161.400 71.800 162.500 72.100 ;
        RECT 159.800 69.800 160.200 70.200 ;
        RECT 159.800 69.200 160.100 69.800 ;
        RECT 151.000 65.100 151.400 67.900 ;
        RECT 151.800 67.800 152.200 68.200 ;
        RECT 151.800 67.200 152.100 67.800 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 152.600 63.100 153.000 68.900 ;
        RECT 155.800 66.800 156.200 67.200 ;
        RECT 155.800 66.200 156.100 66.800 ;
        RECT 155.800 65.800 156.200 66.200 ;
        RECT 153.400 64.800 153.800 65.200 ;
        RECT 148.600 61.800 149.000 62.200 ;
        RECT 148.600 61.200 148.900 61.800 ;
        RECT 153.400 61.200 153.700 64.800 ;
        RECT 157.400 63.100 157.800 68.900 ;
        RECT 159.800 68.800 160.200 69.200 ;
        RECT 161.400 64.200 161.700 71.800 ;
        RECT 165.400 70.800 165.800 71.200 ;
        RECT 162.200 67.100 162.600 67.200 ;
        RECT 163.000 67.100 163.400 67.200 ;
        RECT 162.200 66.800 163.400 67.100 ;
        RECT 165.400 66.200 165.700 70.800 ;
        RECT 166.200 67.200 166.500 73.800 ;
        RECT 171.800 73.100 172.200 75.900 ;
        RECT 172.600 73.800 173.000 74.200 ;
        RECT 167.000 70.800 167.400 71.200 ;
        RECT 167.000 67.200 167.300 70.800 ;
        RECT 172.600 69.200 172.900 73.800 ;
        RECT 173.400 72.100 173.800 77.900 ;
        RECT 174.200 75.800 174.600 76.200 ;
        RECT 174.200 75.100 174.500 75.800 ;
        RECT 174.200 74.700 174.600 75.100 ;
        RECT 177.400 72.200 177.700 90.800 ;
        RECT 178.200 83.100 178.600 88.900 ;
        RECT 179.800 85.100 180.200 87.900 ;
        RECT 180.600 86.800 181.000 87.200 ;
        RECT 180.600 86.200 180.900 86.800 ;
        RECT 180.600 85.800 181.000 86.200 ;
        RECT 177.400 71.800 177.800 72.200 ;
        RECT 178.200 72.100 178.600 77.900 ;
        RECT 179.000 76.800 179.400 77.200 ;
        RECT 172.600 68.800 173.000 69.200 ;
        RECT 174.200 68.800 174.600 69.200 ;
        RECT 167.800 68.100 168.200 68.200 ;
        RECT 167.800 67.800 168.900 68.100 ;
        RECT 168.600 67.200 168.900 67.800 ;
        RECT 169.400 67.800 169.800 68.200 ;
        RECT 171.800 68.100 172.200 68.200 ;
        RECT 172.600 68.100 173.000 68.200 ;
        RECT 171.800 67.800 173.000 68.100 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 167.000 66.800 167.400 67.200 ;
        RECT 168.600 66.800 169.000 67.200 ;
        RECT 169.400 66.200 169.700 67.800 ;
        RECT 170.200 66.800 170.600 67.200 ;
        RECT 173.400 66.800 173.800 67.200 ;
        RECT 170.200 66.200 170.500 66.800 ;
        RECT 173.400 66.200 173.700 66.800 ;
        RECT 164.600 65.800 165.000 66.200 ;
        RECT 165.400 65.800 165.800 66.200 ;
        RECT 167.800 65.800 168.200 66.200 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 171.000 65.800 171.400 66.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 164.600 65.200 164.900 65.800 ;
        RECT 167.800 65.200 168.100 65.800 ;
        RECT 162.200 65.100 162.600 65.200 ;
        RECT 163.000 65.100 163.400 65.200 ;
        RECT 162.200 64.800 163.400 65.100 ;
        RECT 164.600 64.800 165.000 65.200 ;
        RECT 167.800 64.800 168.200 65.200 ;
        RECT 161.400 63.800 161.800 64.200 ;
        RECT 148.600 60.800 149.000 61.200 ;
        RECT 153.400 60.800 153.800 61.200 ;
        RECT 153.400 57.200 153.700 60.800 ;
        RECT 161.400 59.800 161.800 60.200 ;
        RECT 153.400 56.800 153.800 57.200 ;
        RECT 155.800 56.800 156.200 57.200 ;
        RECT 153.400 55.200 153.700 56.800 ;
        RECT 155.800 56.200 156.100 56.800 ;
        RECT 155.800 55.800 156.200 56.200 ;
        RECT 149.400 54.800 149.800 55.200 ;
        RECT 150.200 54.800 150.600 55.200 ;
        RECT 152.600 54.800 153.000 55.200 ;
        RECT 153.400 54.800 153.800 55.200 ;
        RECT 155.000 54.800 155.400 55.200 ;
        RECT 149.400 54.200 149.700 54.800 ;
        RECT 150.200 54.200 150.500 54.800 ;
        RECT 152.600 54.200 152.900 54.800 ;
        RECT 155.000 54.200 155.300 54.800 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 150.200 53.800 150.600 54.200 ;
        RECT 152.600 53.800 153.000 54.200 ;
        RECT 155.000 53.800 155.400 54.200 ;
        RECT 157.400 53.800 157.800 54.200 ;
        RECT 149.400 49.200 149.700 53.800 ;
        RECT 152.600 51.800 153.000 52.200 ;
        RECT 152.600 49.200 152.900 51.800 ;
        RECT 155.800 49.800 156.200 50.200 ;
        RECT 149.400 48.800 149.800 49.200 ;
        RECT 152.600 48.800 153.000 49.200 ;
        RECT 151.800 47.800 152.200 48.200 ;
        RECT 151.800 46.200 152.100 47.800 ;
        RECT 155.800 47.200 156.100 49.800 ;
        RECT 156.600 48.800 157.000 49.200 ;
        RECT 154.200 46.800 154.600 47.200 ;
        RECT 155.800 46.800 156.200 47.200 ;
        RECT 154.200 46.200 154.500 46.800 ;
        RECT 155.800 46.200 156.100 46.800 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 154.200 45.800 154.600 46.200 ;
        RECT 155.000 45.800 155.400 46.200 ;
        RECT 155.800 45.800 156.200 46.200 ;
        RECT 155.000 42.200 155.300 45.800 ;
        RECT 155.000 41.800 155.400 42.200 ;
        RECT 147.000 35.800 147.400 36.200 ;
        RECT 148.600 35.800 149.000 36.200 ;
        RECT 148.600 35.200 148.900 35.800 ;
        RECT 145.400 34.800 145.800 35.200 ;
        RECT 147.800 34.800 148.200 35.200 ;
        RECT 148.600 34.800 149.000 35.200 ;
        RECT 145.400 34.200 145.700 34.800 ;
        RECT 145.400 33.800 145.800 34.200 ;
        RECT 147.000 33.800 147.400 34.200 ;
        RECT 145.400 31.800 145.800 32.200 ;
        RECT 144.600 26.800 145.000 27.200 ;
        RECT 143.800 25.800 144.200 26.200 ;
        RECT 139.800 24.800 140.200 25.200 ;
        RECT 142.200 24.800 142.600 25.200 ;
        RECT 138.200 16.800 138.600 17.200 ;
        RECT 136.600 13.800 137.000 14.200 ;
        RECT 136.600 11.200 136.900 13.800 ;
        RECT 137.400 13.100 137.800 15.900 ;
        RECT 138.200 14.200 138.500 16.800 ;
        RECT 139.800 16.200 140.100 24.800 ;
        RECT 143.800 24.200 144.100 25.800 ;
        RECT 143.800 23.800 144.200 24.200 ;
        RECT 139.000 16.100 139.400 16.200 ;
        RECT 139.800 16.100 140.200 16.200 ;
        RECT 139.000 15.800 140.200 16.100 ;
        RECT 141.400 15.800 141.800 16.200 ;
        RECT 143.000 16.100 143.400 16.200 ;
        RECT 143.800 16.100 144.200 16.200 ;
        RECT 143.000 15.800 144.200 16.100 ;
        RECT 139.800 15.200 140.100 15.800 ;
        RECT 139.800 14.800 140.200 15.200 ;
        RECT 138.200 13.800 138.600 14.200 ;
        RECT 139.800 14.100 140.200 14.200 ;
        RECT 140.600 14.100 141.000 14.200 ;
        RECT 139.800 13.800 141.000 14.100 ;
        RECT 133.400 10.800 133.800 11.200 ;
        RECT 136.600 10.800 137.000 11.200 ;
        RECT 139.000 9.800 139.400 10.200 ;
        RECT 139.000 9.200 139.300 9.800 ;
        RECT 132.600 7.800 133.000 8.200 ;
        RECT 133.400 6.800 133.800 7.200 ;
        RECT 133.400 6.200 133.700 6.800 ;
        RECT 133.400 5.800 133.800 6.200 ;
        RECT 136.600 3.100 137.000 8.900 ;
        RECT 139.000 8.800 139.400 9.200 ;
        RECT 139.800 7.100 140.200 7.200 ;
        RECT 140.600 7.100 141.000 7.200 ;
        RECT 139.800 6.800 141.000 7.100 ;
        RECT 141.400 6.200 141.700 15.800 ;
        RECT 142.200 15.100 142.600 15.200 ;
        RECT 143.000 15.100 143.400 15.200 ;
        RECT 142.200 14.800 143.400 15.100 ;
        RECT 144.600 14.200 144.900 26.800 ;
        RECT 145.400 26.200 145.700 31.800 ;
        RECT 147.000 29.200 147.300 33.800 ;
        RECT 147.800 31.200 148.100 34.800 ;
        RECT 151.000 31.800 151.400 32.200 ;
        RECT 153.400 32.100 153.800 37.900 ;
        RECT 155.800 37.800 156.200 38.200 ;
        RECT 147.800 30.800 148.200 31.200 ;
        RECT 147.000 28.800 147.400 29.200 ;
        RECT 151.000 27.200 151.300 31.800 ;
        RECT 153.400 30.800 153.800 31.200 ;
        RECT 151.800 29.800 152.200 30.200 ;
        RECT 146.200 26.800 146.600 27.200 ;
        RECT 151.000 26.800 151.400 27.200 ;
        RECT 146.200 26.200 146.500 26.800 ;
        RECT 151.800 26.200 152.100 29.800 ;
        RECT 153.400 29.200 153.700 30.800 ;
        RECT 153.400 28.800 153.800 29.200 ;
        RECT 155.000 26.800 155.400 27.200 ;
        RECT 155.000 26.200 155.300 26.800 ;
        RECT 155.800 26.200 156.100 37.800 ;
        RECT 156.600 34.200 156.900 48.800 ;
        RECT 157.400 48.200 157.700 53.800 ;
        RECT 158.200 53.100 158.600 55.900 ;
        RECT 159.000 53.800 159.400 54.200 ;
        RECT 158.200 51.800 158.600 52.200 ;
        RECT 158.200 49.200 158.500 51.800 ;
        RECT 159.000 49.200 159.300 53.800 ;
        RECT 159.800 52.100 160.200 57.900 ;
        RECT 160.600 55.800 161.000 56.200 ;
        RECT 160.600 55.100 160.900 55.800 ;
        RECT 160.600 54.700 161.000 55.100 ;
        RECT 158.200 48.800 158.600 49.200 ;
        RECT 159.000 48.800 159.400 49.200 ;
        RECT 157.400 47.800 157.800 48.200 ;
        RECT 159.000 46.800 159.400 47.200 ;
        RECT 159.800 47.100 160.200 47.200 ;
        RECT 160.600 47.100 161.000 47.200 ;
        RECT 159.800 46.800 161.000 47.100 ;
        RECT 157.400 45.800 157.800 46.200 ;
        RECT 157.400 45.200 157.700 45.800 ;
        RECT 157.400 44.800 157.800 45.200 ;
        RECT 157.400 34.700 157.800 35.100 ;
        RECT 157.400 34.200 157.700 34.700 ;
        RECT 156.600 33.800 157.000 34.200 ;
        RECT 157.400 33.800 157.800 34.200 ;
        RECT 157.400 32.800 157.800 33.200 ;
        RECT 145.400 25.800 145.800 26.200 ;
        RECT 146.200 25.800 146.600 26.200 ;
        RECT 148.600 25.800 149.000 26.200 ;
        RECT 151.800 25.800 152.200 26.200 ;
        RECT 152.600 25.800 153.000 26.200 ;
        RECT 155.000 25.800 155.400 26.200 ;
        RECT 155.800 25.800 156.200 26.200 ;
        RECT 156.600 25.800 157.000 26.200 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 146.200 16.200 146.500 18.800 ;
        RECT 146.200 15.800 146.600 16.200 ;
        RECT 143.000 13.800 143.400 14.200 ;
        RECT 144.600 13.800 145.000 14.200 ;
        RECT 145.400 13.800 145.800 14.200 ;
        RECT 147.800 14.100 148.200 14.200 ;
        RECT 148.600 14.100 148.900 25.800 ;
        RECT 151.000 15.100 151.400 15.200 ;
        RECT 151.800 15.100 152.200 15.200 ;
        RECT 151.000 14.800 152.200 15.100 ;
        RECT 147.800 13.800 148.900 14.100 ;
        RECT 149.400 13.800 149.800 14.200 ;
        RECT 143.000 9.200 143.300 13.800 ;
        RECT 143.800 12.100 144.200 12.200 ;
        RECT 144.600 12.100 145.000 12.200 ;
        RECT 143.800 11.800 145.000 12.100 ;
        RECT 145.400 10.200 145.700 13.800 ;
        RECT 146.200 11.800 146.600 12.200 ;
        RECT 145.400 9.800 145.800 10.200 ;
        RECT 143.000 8.800 143.400 9.200 ;
        RECT 143.000 7.800 143.400 8.200 ;
        RECT 143.000 7.200 143.300 7.800 ;
        RECT 143.000 6.800 143.400 7.200 ;
        RECT 143.800 6.800 144.200 7.200 ;
        RECT 143.800 6.200 144.100 6.800 ;
        RECT 139.800 5.800 140.200 6.200 ;
        RECT 141.400 5.800 141.800 6.200 ;
        RECT 143.800 5.800 144.200 6.200 ;
        RECT 139.800 5.200 140.100 5.800 ;
        RECT 141.400 5.200 141.700 5.800 ;
        RECT 146.200 5.200 146.500 11.800 ;
        RECT 147.800 9.200 148.100 13.800 ;
        RECT 149.400 13.200 149.700 13.800 ;
        RECT 149.400 12.800 149.800 13.200 ;
        RECT 152.600 10.200 152.900 25.800 ;
        RECT 154.200 22.800 154.600 23.200 ;
        RECT 154.200 15.200 154.500 22.800 ;
        RECT 156.600 20.200 156.900 25.800 ;
        RECT 156.600 19.800 157.000 20.200 ;
        RECT 156.600 16.200 156.900 19.800 ;
        RECT 156.600 15.800 157.000 16.200 ;
        RECT 156.600 15.200 156.900 15.800 ;
        RECT 153.400 14.800 153.800 15.200 ;
        RECT 154.200 14.800 154.600 15.200 ;
        RECT 155.000 14.800 155.400 15.200 ;
        RECT 156.600 14.800 157.000 15.200 ;
        RECT 152.600 9.800 153.000 10.200 ;
        RECT 153.400 9.200 153.700 14.800 ;
        RECT 155.000 14.200 155.300 14.800 ;
        RECT 155.000 13.800 155.400 14.200 ;
        RECT 147.800 8.800 148.200 9.200 ;
        RECT 147.000 6.800 147.400 7.200 ;
        RECT 147.000 6.200 147.300 6.800 ;
        RECT 147.000 5.800 147.400 6.200 ;
        RECT 139.800 4.800 140.200 5.200 ;
        RECT 141.400 4.800 141.800 5.200 ;
        RECT 146.200 4.800 146.600 5.200 ;
        RECT 150.200 3.100 150.600 8.900 ;
        RECT 153.400 8.800 153.800 9.200 ;
        RECT 152.600 6.100 153.000 6.200 ;
        RECT 153.400 6.100 153.800 6.200 ;
        RECT 152.600 5.800 153.800 6.100 ;
        RECT 155.000 3.100 155.400 8.900 ;
        RECT 155.800 6.800 156.200 7.200 ;
        RECT 155.800 6.200 156.100 6.800 ;
        RECT 155.800 5.800 156.200 6.200 ;
        RECT 156.600 5.100 157.000 7.900 ;
        RECT 157.400 7.200 157.700 32.800 ;
        RECT 158.200 32.100 158.600 37.900 ;
        RECT 159.000 29.200 159.300 46.800 ;
        RECT 159.800 46.100 160.200 46.200 ;
        RECT 160.600 46.100 161.000 46.200 ;
        RECT 159.800 45.800 161.000 46.100 ;
        RECT 161.400 39.200 161.700 59.800 ;
        RECT 164.600 52.100 165.000 57.900 ;
        RECT 167.000 51.800 167.400 52.200 ;
        RECT 167.800 51.800 168.200 52.200 ;
        RECT 170.200 52.100 170.600 57.900 ;
        RECT 162.200 49.100 162.600 49.200 ;
        RECT 163.000 49.100 163.400 49.200 ;
        RECT 162.200 48.800 163.400 49.100 ;
        RECT 167.000 48.200 167.300 51.800 ;
        RECT 167.800 50.200 168.100 51.800 ;
        RECT 168.600 50.800 169.000 51.200 ;
        RECT 167.800 49.800 168.200 50.200 ;
        RECT 168.600 49.200 168.900 50.800 ;
        RECT 168.600 48.800 169.000 49.200 ;
        RECT 167.000 47.800 167.400 48.200 ;
        RECT 165.400 43.800 165.800 44.200 ;
        RECT 165.400 42.200 165.700 43.800 ;
        RECT 169.400 42.800 169.800 43.200 ;
        RECT 165.400 41.800 165.800 42.200 ;
        RECT 161.400 38.800 161.800 39.200 ;
        RECT 159.800 33.100 160.200 35.900 ;
        RECT 165.400 35.200 165.700 41.800 ;
        RECT 166.200 36.100 166.600 36.200 ;
        RECT 167.000 36.100 167.400 36.200 ;
        RECT 166.200 35.800 167.400 36.100 ;
        RECT 165.400 34.800 165.800 35.200 ;
        RECT 162.200 33.800 162.600 34.200 ;
        RECT 161.400 31.800 161.800 32.200 ;
        RECT 161.400 30.200 161.700 31.800 ;
        RECT 161.400 29.800 161.800 30.200 ;
        RECT 162.200 29.200 162.500 33.800 ;
        RECT 158.200 29.100 158.600 29.200 ;
        RECT 159.000 29.100 159.400 29.200 ;
        RECT 158.200 28.800 159.400 29.100 ;
        RECT 162.200 28.800 162.600 29.200 ;
        RECT 164.600 28.800 165.000 29.200 ;
        RECT 164.600 27.200 164.900 28.800 ;
        RECT 159.000 26.800 159.400 27.200 ;
        RECT 163.800 26.800 164.200 27.200 ;
        RECT 164.600 26.800 165.000 27.200 ;
        RECT 159.000 26.200 159.300 26.800 ;
        RECT 163.800 26.200 164.100 26.800 ;
        RECT 166.200 26.200 166.500 35.800 ;
        RECT 169.400 35.200 169.700 42.800 ;
        RECT 171.000 39.200 171.300 65.800 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 173.400 52.200 173.700 54.800 ;
        RECT 174.200 54.200 174.500 68.800 ;
        RECT 175.000 65.100 175.400 67.900 ;
        RECT 176.600 63.100 177.000 68.900 ;
        RECT 177.400 68.200 177.700 71.800 ;
        RECT 177.400 67.800 177.800 68.200 ;
        RECT 179.000 66.200 179.300 76.800 ;
        RECT 181.400 76.200 181.700 99.800 ;
        RECT 182.200 92.100 182.600 97.900 ;
        RECT 183.000 95.200 183.300 121.800 ;
        RECT 187.000 120.200 187.300 134.800 ;
        RECT 189.400 134.200 189.700 134.800 ;
        RECT 188.600 133.800 189.000 134.200 ;
        RECT 189.400 133.800 189.800 134.200 ;
        RECT 188.600 133.200 188.900 133.800 ;
        RECT 188.600 132.800 189.000 133.200 ;
        RECT 188.600 130.200 188.900 132.800 ;
        RECT 188.600 129.800 189.000 130.200 ;
        RECT 189.400 126.800 189.800 127.200 ;
        RECT 189.400 126.200 189.700 126.800 ;
        RECT 190.200 126.200 190.500 150.800 ;
        RECT 195.000 148.800 195.400 149.200 ;
        RECT 192.600 147.800 193.000 148.200 ;
        RECT 192.600 146.200 192.900 147.800 ;
        RECT 195.000 146.200 195.300 148.800 ;
        RECT 195.800 146.800 196.200 147.200 ;
        RECT 191.000 146.100 191.400 146.200 ;
        RECT 191.800 146.100 192.200 146.200 ;
        RECT 191.000 145.800 192.200 146.100 ;
        RECT 192.600 145.800 193.000 146.200 ;
        RECT 195.000 145.800 195.400 146.200 ;
        RECT 195.800 145.100 196.100 146.800 ;
        RECT 195.000 144.800 196.100 145.100 ;
        RECT 193.400 141.800 193.800 142.200 ;
        RECT 193.400 141.200 193.700 141.800 ;
        RECT 193.400 140.800 193.800 141.200 ;
        RECT 192.600 139.800 193.000 140.200 ;
        RECT 191.000 136.800 191.400 137.200 ;
        RECT 191.000 135.200 191.300 136.800 ;
        RECT 191.000 134.800 191.400 135.200 ;
        RECT 191.000 130.800 191.400 131.200 ;
        RECT 191.000 129.200 191.300 130.800 ;
        RECT 191.000 128.800 191.400 129.200 ;
        RECT 191.000 127.800 191.400 128.200 ;
        RECT 191.000 127.200 191.300 127.800 ;
        RECT 192.600 127.200 192.900 139.800 ;
        RECT 194.200 137.800 194.600 138.200 ;
        RECT 194.200 135.200 194.500 137.800 ;
        RECT 193.400 134.800 193.800 135.200 ;
        RECT 194.200 134.800 194.600 135.200 ;
        RECT 193.400 129.200 193.700 134.800 ;
        RECT 195.000 134.200 195.300 144.800 ;
        RECT 195.800 135.800 196.200 136.200 ;
        RECT 195.800 135.200 196.100 135.800 ;
        RECT 195.800 134.800 196.200 135.200 ;
        RECT 194.200 134.100 194.600 134.200 ;
        RECT 195.000 134.100 195.400 134.200 ;
        RECT 194.200 133.800 195.400 134.100 ;
        RECT 193.400 128.800 193.800 129.200 ;
        RECT 191.000 126.800 191.400 127.200 ;
        RECT 192.600 126.800 193.000 127.200 ;
        RECT 195.000 126.800 195.400 127.200 ;
        RECT 188.600 125.800 189.000 126.200 ;
        RECT 189.400 125.800 189.800 126.200 ;
        RECT 190.200 125.800 190.600 126.200 ;
        RECT 191.000 125.800 191.400 126.200 ;
        RECT 183.800 119.800 184.200 120.200 ;
        RECT 187.000 119.800 187.400 120.200 ;
        RECT 183.800 115.200 184.100 119.800 ;
        RECT 187.000 116.800 187.400 117.200 ;
        RECT 187.000 116.200 187.300 116.800 ;
        RECT 185.400 116.100 185.800 116.200 ;
        RECT 186.200 116.100 186.600 116.200 ;
        RECT 185.400 115.800 186.600 116.100 ;
        RECT 187.000 115.800 187.400 116.200 ;
        RECT 187.800 115.800 188.200 116.200 ;
        RECT 183.800 114.800 184.200 115.200 ;
        RECT 184.600 113.800 185.000 114.200 ;
        RECT 183.800 103.100 184.200 108.900 ;
        RECT 184.600 99.200 184.900 113.800 ;
        RECT 186.200 111.800 186.600 112.200 ;
        RECT 185.400 105.100 185.800 107.900 ;
        RECT 186.200 105.200 186.500 111.800 ;
        RECT 187.800 109.200 188.100 115.800 ;
        RECT 188.600 114.200 188.900 125.800 ;
        RECT 190.200 118.200 190.500 125.800 ;
        RECT 190.200 117.800 190.600 118.200 ;
        RECT 188.600 113.800 189.000 114.200 ;
        RECT 187.800 108.800 188.200 109.200 ;
        RECT 188.600 109.100 188.900 113.800 ;
        RECT 189.400 111.800 189.800 112.200 ;
        RECT 189.400 110.200 189.700 111.800 ;
        RECT 189.400 109.800 189.800 110.200 ;
        RECT 189.400 109.100 189.800 109.200 ;
        RECT 188.600 108.800 189.800 109.100 ;
        RECT 187.800 106.200 188.100 108.800 ;
        RECT 188.600 106.800 189.000 107.200 ;
        RECT 187.800 105.800 188.200 106.200 ;
        RECT 186.200 104.800 186.600 105.200 ;
        RECT 188.600 102.200 188.900 106.800 ;
        RECT 187.800 101.800 188.200 102.200 ;
        RECT 188.600 101.800 189.000 102.200 ;
        RECT 184.600 98.800 185.000 99.200 ;
        RECT 183.000 94.800 183.400 95.200 ;
        RECT 186.200 94.700 186.600 95.100 ;
        RECT 186.200 94.200 186.500 94.700 ;
        RECT 186.200 93.800 186.600 94.200 ;
        RECT 183.800 92.800 184.200 93.200 ;
        RECT 183.800 86.200 184.100 92.800 ;
        RECT 185.400 91.800 185.800 92.200 ;
        RECT 187.000 92.100 187.400 97.900 ;
        RECT 187.800 96.200 188.100 101.800 ;
        RECT 187.800 95.800 188.200 96.200 ;
        RECT 188.600 93.100 189.000 95.900 ;
        RECT 189.400 93.800 189.800 94.200 ;
        RECT 189.400 93.200 189.700 93.800 ;
        RECT 189.400 92.800 189.800 93.200 ;
        RECT 185.400 86.200 185.700 91.800 ;
        RECT 188.600 87.800 189.000 88.200 ;
        RECT 188.600 86.200 188.900 87.800 ;
        RECT 190.200 87.200 190.500 117.800 ;
        RECT 191.000 117.200 191.300 125.800 ;
        RECT 191.000 116.800 191.400 117.200 ;
        RECT 191.000 115.200 191.300 116.800 ;
        RECT 191.000 114.800 191.400 115.200 ;
        RECT 191.000 114.100 191.400 114.200 ;
        RECT 191.800 114.100 192.200 114.200 ;
        RECT 191.000 113.800 192.200 114.100 ;
        RECT 191.800 103.100 192.200 108.900 ;
        RECT 191.000 97.800 191.400 98.200 ;
        RECT 191.000 96.200 191.300 97.800 ;
        RECT 191.000 95.800 191.400 96.200 ;
        RECT 191.000 94.800 191.400 95.200 ;
        RECT 191.000 94.200 191.300 94.800 ;
        RECT 191.000 93.800 191.400 94.200 ;
        RECT 190.200 86.800 190.600 87.200 ;
        RECT 191.800 86.800 192.200 87.200 ;
        RECT 182.200 85.800 182.600 86.200 ;
        RECT 183.800 85.800 184.200 86.200 ;
        RECT 184.600 85.800 185.000 86.200 ;
        RECT 185.400 85.800 185.800 86.200 ;
        RECT 186.200 85.800 186.600 86.200 ;
        RECT 188.600 85.800 189.000 86.200 ;
        RECT 189.400 86.100 189.800 86.200 ;
        RECT 190.200 86.100 190.600 86.200 ;
        RECT 189.400 85.800 190.600 86.100 ;
        RECT 191.000 85.800 191.400 86.200 ;
        RECT 182.200 85.200 182.500 85.800 ;
        RECT 182.200 84.800 182.600 85.200 ;
        RECT 183.000 78.800 183.400 79.200 ;
        RECT 181.400 75.800 181.800 76.200 ;
        RECT 183.000 75.200 183.300 78.800 ;
        RECT 184.600 76.200 184.900 85.800 ;
        RECT 186.200 85.200 186.500 85.800 ;
        RECT 191.000 85.200 191.300 85.800 ;
        RECT 186.200 84.800 186.600 85.200 ;
        RECT 191.000 84.800 191.400 85.200 ;
        RECT 189.400 83.800 189.800 84.200 ;
        RECT 187.800 81.800 188.200 82.200 ;
        RECT 187.800 76.200 188.100 81.800 ;
        RECT 184.600 75.800 185.000 76.200 ;
        RECT 187.800 75.800 188.200 76.200 ;
        RECT 189.400 75.200 189.700 83.800 ;
        RECT 183.000 74.800 183.400 75.200 ;
        RECT 183.800 75.100 184.200 75.200 ;
        RECT 184.600 75.100 185.000 75.200 ;
        RECT 183.800 74.800 185.000 75.100 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 187.800 74.800 188.200 75.200 ;
        RECT 188.600 74.800 189.000 75.200 ;
        RECT 189.400 74.800 189.800 75.200 ;
        RECT 190.200 74.800 190.600 75.200 ;
        RECT 180.600 73.800 181.000 74.200 ;
        RECT 183.800 74.100 184.200 74.200 ;
        RECT 183.800 73.800 184.900 74.100 ;
        RECT 180.600 72.200 180.900 73.800 ;
        RECT 181.400 72.800 181.800 73.200 ;
        RECT 181.400 72.200 181.700 72.800 ;
        RECT 180.600 71.800 181.000 72.200 ;
        RECT 181.400 71.800 181.800 72.200 ;
        RECT 183.800 71.800 184.200 72.200 ;
        RECT 183.800 69.200 184.100 71.800 ;
        RECT 184.600 69.200 184.900 73.800 ;
        RECT 185.400 70.200 185.700 74.800 ;
        RECT 187.800 74.200 188.100 74.800 ;
        RECT 188.600 74.200 188.900 74.800 ;
        RECT 190.200 74.200 190.500 74.800 ;
        RECT 187.800 73.800 188.200 74.200 ;
        RECT 188.600 73.800 189.000 74.200 ;
        RECT 190.200 73.800 190.600 74.200 ;
        RECT 191.000 71.800 191.400 72.200 ;
        RECT 191.000 71.200 191.300 71.800 ;
        RECT 191.000 70.800 191.400 71.200 ;
        RECT 185.400 69.800 185.800 70.200 ;
        RECT 179.000 65.800 179.400 66.200 ;
        RECT 181.400 63.100 181.800 68.900 ;
        RECT 183.800 68.800 184.200 69.200 ;
        RECT 184.600 68.800 185.000 69.200 ;
        RECT 186.200 68.800 186.600 69.200 ;
        RECT 186.200 67.200 186.500 68.800 ;
        RECT 188.600 68.100 189.000 68.200 ;
        RECT 189.400 68.100 189.800 68.200 ;
        RECT 188.600 67.800 189.800 68.100 ;
        RECT 186.200 66.800 186.600 67.200 ;
        RECT 191.800 66.200 192.100 86.800 ;
        RECT 192.600 85.200 192.900 126.800 ;
        RECT 195.000 126.200 195.300 126.800 ;
        RECT 195.000 125.800 195.400 126.200 ;
        RECT 195.800 117.200 196.100 134.800 ;
        RECT 195.800 116.800 196.200 117.200 ;
        RECT 195.800 115.800 196.200 116.200 ;
        RECT 195.800 115.200 196.100 115.800 ;
        RECT 193.400 114.800 193.800 115.200 ;
        RECT 195.800 115.100 196.200 115.200 ;
        RECT 196.600 115.100 196.900 154.800 ;
        RECT 198.200 154.200 198.500 159.800 ;
        RECT 201.400 159.200 201.700 165.800 ;
        RECT 201.400 158.800 201.800 159.200 ;
        RECT 201.400 155.800 201.800 156.200 ;
        RECT 202.200 155.800 202.600 156.200 ;
        RECT 203.000 155.800 203.400 156.200 ;
        RECT 199.000 154.800 199.400 155.200 ;
        RECT 198.200 153.800 198.600 154.200 ;
        RECT 199.000 152.200 199.300 154.800 ;
        RECT 201.400 154.200 201.700 155.800 ;
        RECT 202.200 155.200 202.500 155.800 ;
        RECT 202.200 154.800 202.600 155.200 ;
        RECT 201.400 153.800 201.800 154.200 ;
        RECT 203.000 152.200 203.300 155.800 ;
        RECT 199.000 151.800 199.400 152.200 ;
        RECT 203.000 151.800 203.400 152.200 ;
        RECT 199.000 147.100 199.400 147.200 ;
        RECT 199.800 147.100 200.200 147.200 ;
        RECT 199.000 146.800 200.200 147.100 ;
        RECT 202.200 147.100 202.600 147.200 ;
        RECT 203.000 147.100 203.400 147.200 ;
        RECT 202.200 146.800 203.400 147.100 ;
        RECT 203.800 146.200 204.100 173.800 ;
        RECT 207.800 173.200 208.100 174.800 ;
        RECT 208.600 174.200 208.900 193.800 ;
        RECT 210.200 192.100 210.600 197.900 ;
        RECT 213.400 196.100 213.800 196.200 ;
        RECT 214.200 196.100 214.600 196.200 ;
        RECT 211.800 193.100 212.200 195.900 ;
        RECT 213.400 195.800 214.600 196.100 ;
        RECT 215.000 195.800 215.400 196.200 ;
        RECT 213.400 195.100 213.800 195.200 ;
        RECT 213.400 194.800 214.500 195.100 ;
        RECT 212.600 194.100 213.000 194.200 ;
        RECT 213.400 194.100 213.800 194.200 ;
        RECT 212.600 193.800 213.800 194.100 ;
        RECT 213.400 191.800 213.800 192.200 ;
        RECT 211.800 189.800 212.200 190.200 ;
        RECT 211.000 183.100 211.400 188.900 ;
        RECT 211.800 187.200 212.100 189.800 ;
        RECT 211.800 186.800 212.200 187.200 ;
        RECT 211.800 179.200 212.100 186.800 ;
        RECT 212.600 185.100 213.000 187.900 ;
        RECT 213.400 187.200 213.700 191.800 ;
        RECT 213.400 186.800 213.800 187.200 ;
        RECT 214.200 183.200 214.500 194.800 ;
        RECT 215.000 189.200 215.300 195.800 ;
        RECT 215.800 194.200 216.100 213.800 ;
        RECT 218.200 198.200 218.500 221.800 ;
        RECT 219.000 213.800 219.400 214.200 ;
        RECT 219.000 212.200 219.300 213.800 ;
        RECT 219.000 211.800 219.400 212.200 ;
        RECT 219.000 206.200 219.300 211.800 ;
        RECT 219.800 210.200 220.100 231.800 ;
        RECT 220.600 226.200 220.900 231.800 ;
        RECT 221.400 228.200 221.700 231.800 ;
        RECT 221.400 227.800 221.800 228.200 ;
        RECT 225.400 227.200 225.700 232.800 ;
        RECT 229.400 232.100 229.800 237.900 ;
        RECT 232.600 233.100 233.000 235.900 ;
        RECT 233.400 234.800 233.800 235.200 ;
        RECT 233.400 234.200 233.700 234.800 ;
        RECT 233.400 233.800 233.800 234.200 ;
        RECT 231.800 232.100 232.200 232.200 ;
        RECT 232.600 232.100 233.000 232.200 ;
        RECT 234.200 232.100 234.600 237.900 ;
        RECT 235.800 235.100 236.200 235.200 ;
        RECT 236.600 235.100 237.000 235.200 ;
        RECT 235.800 234.800 237.000 235.100 ;
        RECT 239.000 232.100 239.400 237.900 ;
        RECT 249.400 235.800 249.800 236.200 ;
        RECT 249.400 235.200 249.700 235.800 ;
        RECT 246.200 235.100 246.600 235.200 ;
        RECT 247.000 235.100 247.400 235.200 ;
        RECT 246.200 234.800 247.400 235.100 ;
        RECT 249.400 234.800 249.800 235.200 ;
        RECT 246.200 233.800 246.600 234.200 ;
        RECT 251.000 233.800 251.400 234.200 ;
        RECT 246.200 233.200 246.500 233.800 ;
        RECT 246.200 232.800 246.600 233.200 ;
        RECT 240.600 232.100 241.000 232.200 ;
        RECT 241.400 232.100 241.800 232.200 ;
        RECT 231.800 231.800 233.000 232.100 ;
        RECT 240.600 231.800 241.800 232.100 ;
        RECT 244.600 232.100 245.000 232.200 ;
        RECT 245.400 232.100 245.800 232.200 ;
        RECT 244.600 231.800 245.800 232.100 ;
        RECT 248.600 231.800 249.000 232.200 ;
        RECT 221.400 227.100 221.800 227.200 ;
        RECT 222.200 227.100 222.600 227.200 ;
        RECT 221.400 226.800 222.600 227.100 ;
        RECT 223.800 226.800 224.200 227.200 ;
        RECT 225.400 226.800 225.800 227.200 ;
        RECT 228.600 226.800 229.000 227.200 ;
        RECT 230.200 226.800 230.600 227.200 ;
        RECT 223.800 226.200 224.100 226.800 ;
        RECT 220.600 225.800 221.000 226.200 ;
        RECT 223.800 225.800 224.200 226.200 ;
        RECT 224.600 225.800 225.000 226.200 ;
        RECT 224.600 223.200 224.900 225.800 ;
        RECT 224.600 222.800 225.000 223.200 ;
        RECT 225.400 222.200 225.700 226.800 ;
        RECT 228.600 226.200 228.900 226.800 ;
        RECT 230.200 226.200 230.500 226.800 ;
        RECT 226.200 225.800 226.600 226.200 ;
        RECT 228.600 225.800 229.000 226.200 ;
        RECT 230.200 225.800 230.600 226.200 ;
        RECT 226.200 225.200 226.500 225.800 ;
        RECT 226.200 224.800 226.600 225.200 ;
        RECT 227.800 225.100 228.200 225.200 ;
        RECT 228.600 225.100 229.000 225.200 ;
        RECT 227.800 224.800 229.000 225.100 ;
        RECT 233.400 223.100 233.800 228.900 ;
        RECT 235.800 226.100 236.200 226.200 ;
        RECT 236.600 226.100 237.000 226.200 ;
        RECT 235.800 225.800 237.000 226.100 ;
        RECT 238.200 223.100 238.600 228.900 ;
        RECT 239.000 226.800 239.400 227.200 ;
        RECT 239.000 226.200 239.300 226.800 ;
        RECT 239.000 225.800 239.400 226.200 ;
        RECT 225.400 221.800 225.800 222.200 ;
        RECT 235.000 221.800 235.400 222.200 ;
        RECT 223.800 219.800 224.200 220.200 ;
        RECT 221.400 216.800 221.800 217.200 ;
        RECT 221.400 216.200 221.700 216.800 ;
        RECT 221.400 215.800 221.800 216.200 ;
        RECT 220.600 215.100 221.000 215.200 ;
        RECT 221.400 215.100 221.800 215.200 ;
        RECT 220.600 214.800 221.800 215.100 ;
        RECT 221.400 214.100 221.800 214.200 ;
        RECT 222.200 214.100 222.600 214.200 ;
        RECT 221.400 213.800 222.600 214.100 ;
        RECT 223.000 213.100 223.400 215.900 ;
        RECT 223.800 214.200 224.100 219.800 ;
        RECT 234.200 218.800 234.600 219.200 ;
        RECT 223.800 213.800 224.200 214.200 ;
        RECT 224.600 212.100 225.000 217.900 ;
        RECT 225.400 215.800 225.800 216.200 ;
        RECT 225.400 215.100 225.700 215.800 ;
        RECT 225.400 214.700 225.800 215.100 ;
        RECT 229.400 212.100 229.800 217.900 ;
        RECT 232.600 215.800 233.000 216.200 ;
        RECT 231.000 212.100 231.400 212.200 ;
        RECT 231.800 212.100 232.200 212.200 ;
        RECT 231.000 211.800 232.200 212.100 ;
        RECT 232.600 211.100 232.900 215.800 ;
        RECT 234.200 215.200 234.500 218.800 ;
        RECT 235.000 215.200 235.300 221.800 ;
        RECT 236.600 216.100 237.000 216.200 ;
        RECT 237.400 216.100 237.800 216.200 ;
        RECT 236.600 215.800 237.800 216.100 ;
        RECT 234.200 214.800 234.600 215.200 ;
        RECT 235.000 214.800 235.400 215.200 ;
        RECT 231.800 210.800 232.900 211.100 ;
        RECT 233.400 213.800 233.800 214.200 ;
        RECT 219.800 209.800 220.200 210.200 ;
        RECT 226.200 209.800 226.600 210.200 ;
        RECT 225.400 208.800 225.800 209.200 ;
        RECT 219.800 206.800 220.200 207.200 ;
        RECT 223.800 206.800 224.200 207.200 ;
        RECT 219.000 205.800 219.400 206.200 ;
        RECT 218.200 197.800 218.600 198.200 ;
        RECT 216.600 195.800 217.000 196.200 ;
        RECT 218.200 196.100 218.600 196.200 ;
        RECT 219.000 196.100 219.400 196.200 ;
        RECT 218.200 195.800 219.400 196.100 ;
        RECT 216.600 195.200 216.900 195.800 ;
        RECT 216.600 194.800 217.000 195.200 ;
        RECT 219.000 194.800 219.400 195.200 ;
        RECT 219.000 194.200 219.300 194.800 ;
        RECT 215.800 193.800 216.200 194.200 ;
        RECT 219.000 193.800 219.400 194.200 ;
        RECT 219.800 190.200 220.100 206.800 ;
        RECT 223.800 206.200 224.100 206.800 ;
        RECT 225.400 206.200 225.700 208.800 ;
        RECT 226.200 206.200 226.500 209.800 ;
        RECT 231.800 209.200 232.100 210.800 ;
        RECT 228.600 208.800 229.000 209.200 ;
        RECT 231.800 208.800 232.200 209.200 ;
        RECT 232.600 208.800 233.000 209.200 ;
        RECT 228.600 206.200 228.900 208.800 ;
        RECT 232.600 207.200 232.900 208.800 ;
        RECT 229.400 207.100 229.800 207.200 ;
        RECT 230.200 207.100 230.600 207.200 ;
        RECT 229.400 206.800 230.600 207.100 ;
        RECT 232.600 206.800 233.000 207.200 ;
        RECT 233.400 206.200 233.700 213.800 ;
        RECT 220.600 206.100 221.000 206.200 ;
        RECT 221.400 206.100 221.800 206.200 ;
        RECT 220.600 205.800 221.800 206.100 ;
        RECT 223.800 205.800 224.200 206.200 ;
        RECT 224.600 205.800 225.000 206.200 ;
        RECT 225.400 205.800 225.800 206.200 ;
        RECT 226.200 205.800 226.600 206.200 ;
        RECT 228.600 205.800 229.000 206.200 ;
        RECT 233.400 205.800 233.800 206.200 ;
        RECT 222.200 201.800 222.600 202.200 ;
        RECT 222.200 200.200 222.500 201.800 ;
        RECT 222.200 199.800 222.600 200.200 ;
        RECT 224.600 199.200 224.900 205.800 ;
        RECT 234.200 205.200 234.500 214.800 ;
        RECT 235.000 214.200 235.300 214.800 ;
        RECT 235.000 213.800 235.400 214.200 ;
        RECT 235.800 213.800 236.200 214.200 ;
        RECT 235.800 210.200 236.100 213.800 ;
        RECT 235.800 209.800 236.200 210.200 ;
        RECT 231.000 205.100 231.400 205.200 ;
        RECT 231.800 205.100 232.200 205.200 ;
        RECT 231.000 204.800 232.200 205.100 ;
        RECT 234.200 204.800 234.600 205.200 ;
        RECT 235.000 203.100 235.400 208.900 ;
        RECT 239.000 208.200 239.300 225.800 ;
        RECT 239.800 225.100 240.200 227.900 ;
        RECT 243.000 223.100 243.400 228.900 ;
        RECT 243.800 226.800 244.200 227.200 ;
        RECT 243.800 226.200 244.100 226.800 ;
        RECT 243.800 226.100 244.200 226.200 ;
        RECT 243.800 225.800 244.900 226.100 ;
        RECT 240.600 222.100 241.000 222.200 ;
        RECT 241.400 222.100 241.800 222.200 ;
        RECT 240.600 221.800 241.800 222.100 ;
        RECT 242.200 221.800 242.600 222.200 ;
        RECT 239.800 220.800 240.200 221.200 ;
        RECT 239.800 219.200 240.100 220.800 ;
        RECT 239.800 218.800 240.200 219.200 ;
        RECT 239.800 215.800 240.200 216.200 ;
        RECT 239.800 215.200 240.100 215.800 ;
        RECT 239.800 214.800 240.200 215.200 ;
        RECT 240.600 214.800 241.000 215.200 ;
        RECT 240.600 214.200 240.900 214.800 ;
        RECT 240.600 214.100 241.000 214.200 ;
        RECT 241.400 214.100 241.800 214.200 ;
        RECT 240.600 213.800 241.800 214.100 ;
        RECT 240.600 212.100 241.000 212.200 ;
        RECT 241.400 212.100 241.800 212.200 ;
        RECT 240.600 211.800 241.800 212.100 ;
        RECT 240.600 209.200 240.900 211.800 ;
        RECT 239.000 207.800 239.400 208.200 ;
        RECT 235.800 206.100 236.200 206.200 ;
        RECT 236.600 206.100 237.000 206.200 ;
        RECT 235.800 205.800 237.000 206.100 ;
        RECT 239.800 203.100 240.200 208.900 ;
        RECT 240.600 208.800 241.000 209.200 ;
        RECT 242.200 208.200 242.500 221.800 ;
        RECT 243.800 212.100 244.200 217.900 ;
        RECT 244.600 215.200 244.900 225.800 ;
        RECT 247.000 225.900 247.400 226.300 ;
        RECT 247.000 225.200 247.300 225.900 ;
        RECT 247.000 224.800 247.400 225.200 ;
        RECT 247.800 223.100 248.200 228.900 ;
        RECT 248.600 219.200 248.900 231.800 ;
        RECT 249.400 225.100 249.800 227.900 ;
        RECT 248.600 218.800 249.000 219.200 ;
        RECT 245.400 215.800 245.800 216.200 ;
        RECT 244.600 214.800 245.000 215.200 ;
        RECT 244.600 211.800 245.000 212.200 ;
        RECT 244.600 208.200 244.900 211.800 ;
        RECT 241.400 205.100 241.800 207.900 ;
        RECT 242.200 207.800 242.600 208.200 ;
        RECT 244.600 207.800 245.000 208.200 ;
        RECT 242.200 207.200 242.500 207.800 ;
        RECT 242.200 206.800 242.600 207.200 ;
        RECT 243.800 204.800 244.200 205.200 ;
        RECT 227.000 201.800 227.400 202.200 ;
        RECT 243.000 201.800 243.400 202.200 ;
        RECT 224.600 198.800 225.000 199.200 ;
        RECT 221.400 197.800 221.800 198.200 ;
        RECT 220.600 196.800 221.000 197.200 ;
        RECT 220.600 194.200 220.900 196.800 ;
        RECT 220.600 193.800 221.000 194.200 ;
        RECT 219.800 189.800 220.200 190.200 ;
        RECT 215.000 188.800 215.400 189.200 ;
        RECT 219.800 186.800 220.200 187.200 ;
        RECT 215.000 186.100 215.400 186.200 ;
        RECT 215.800 186.100 216.200 186.200 ;
        RECT 215.000 185.800 216.200 186.100 ;
        RECT 216.600 186.100 217.000 186.200 ;
        RECT 217.400 186.100 217.800 186.200 ;
        RECT 216.600 185.800 217.800 186.100 ;
        RECT 215.000 184.800 215.400 185.200 ;
        RECT 215.000 183.200 215.300 184.800 ;
        RECT 214.200 182.800 214.600 183.200 ;
        RECT 215.000 182.800 215.400 183.200 ;
        RECT 217.400 181.800 217.800 182.200 ;
        RECT 217.400 181.200 217.700 181.800 ;
        RECT 217.400 180.800 217.800 181.200 ;
        RECT 211.800 178.800 212.200 179.200 ;
        RECT 211.000 175.800 211.400 176.200 ;
        RECT 209.400 174.800 209.800 175.200 ;
        RECT 210.200 174.800 210.600 175.200 ;
        RECT 208.600 173.800 209.000 174.200 ;
        RECT 207.800 172.800 208.200 173.200 ;
        RECT 209.400 172.200 209.700 174.800 ;
        RECT 210.200 174.200 210.500 174.800 ;
        RECT 210.200 173.800 210.600 174.200 ;
        RECT 205.400 171.800 205.800 172.200 ;
        RECT 209.400 171.800 209.800 172.200 ;
        RECT 205.400 169.200 205.700 171.800 ;
        RECT 208.600 170.800 209.000 171.200 ;
        RECT 205.400 168.800 205.800 169.200 ;
        RECT 206.200 168.100 206.600 168.200 ;
        RECT 207.000 168.100 207.400 168.200 ;
        RECT 206.200 167.800 207.400 168.100 ;
        RECT 208.600 167.200 208.900 170.800 ;
        RECT 211.000 169.200 211.300 175.800 ;
        RECT 211.800 171.800 212.200 172.200 ;
        RECT 214.200 172.100 214.600 177.900 ;
        RECT 215.000 175.100 215.400 175.200 ;
        RECT 215.800 175.100 216.200 175.200 ;
        RECT 215.000 174.800 216.200 175.100 ;
        RECT 218.200 172.800 218.600 173.200 ;
        RECT 211.800 171.200 212.100 171.800 ;
        RECT 211.800 170.800 212.200 171.200 ;
        RECT 211.000 168.800 211.400 169.200 ;
        RECT 214.200 168.100 214.600 168.200 ;
        RECT 215.000 168.100 215.400 168.200 ;
        RECT 214.200 167.800 215.400 168.100 ;
        RECT 208.600 166.800 209.000 167.200 ;
        RECT 211.800 166.800 212.200 167.200 ;
        RECT 216.600 166.800 217.000 167.200 ;
        RECT 208.600 166.200 208.900 166.800 ;
        RECT 211.800 166.200 212.100 166.800 ;
        RECT 204.600 165.800 205.000 166.200 ;
        RECT 205.400 166.100 205.800 166.200 ;
        RECT 206.200 166.100 206.600 166.200 ;
        RECT 205.400 165.800 206.600 166.100 ;
        RECT 208.600 165.800 209.000 166.200 ;
        RECT 209.400 165.800 209.800 166.200 ;
        RECT 211.800 165.800 212.200 166.200 ;
        RECT 215.800 165.800 216.200 166.200 ;
        RECT 204.600 164.200 204.900 165.800 ;
        RECT 209.400 165.200 209.700 165.800 ;
        RECT 215.800 165.200 216.100 165.800 ;
        RECT 209.400 164.800 209.800 165.200 ;
        RECT 211.000 164.800 211.400 165.200 ;
        RECT 213.400 164.800 213.800 165.200 ;
        RECT 215.800 164.800 216.200 165.200 ;
        RECT 211.000 164.200 211.300 164.800 ;
        RECT 204.600 163.800 205.000 164.200 ;
        RECT 211.000 163.800 211.400 164.200 ;
        RECT 204.600 158.800 205.000 159.200 ;
        RECT 204.600 154.200 204.900 158.800 ;
        RECT 213.400 158.200 213.700 164.800 ;
        RECT 216.600 160.200 216.900 166.800 ;
        RECT 218.200 166.200 218.500 172.800 ;
        RECT 219.000 172.100 219.400 177.900 ;
        RECT 219.800 176.200 220.100 186.800 ;
        RECT 220.600 186.200 220.900 193.800 ;
        RECT 221.400 186.200 221.700 197.800 ;
        RECT 222.200 195.800 222.600 196.200 ;
        RECT 220.600 185.800 221.000 186.200 ;
        RECT 221.400 185.800 221.800 186.200 ;
        RECT 219.800 175.800 220.200 176.200 ;
        RECT 220.600 173.100 221.000 175.900 ;
        RECT 222.200 175.200 222.500 195.800 ;
        RECT 223.800 192.100 224.200 197.900 ;
        RECT 224.600 196.800 225.000 197.200 ;
        RECT 224.600 195.200 224.900 196.800 ;
        RECT 227.000 196.200 227.300 201.800 ;
        RECT 227.000 195.800 227.400 196.200 ;
        RECT 224.600 194.800 225.000 195.200 ;
        RECT 226.200 195.100 226.600 195.200 ;
        RECT 227.000 195.100 227.400 195.200 ;
        RECT 226.200 194.800 227.400 195.100 ;
        RECT 225.400 193.800 225.800 194.200 ;
        RECT 225.400 187.200 225.700 193.800 ;
        RECT 228.600 192.100 229.000 197.900 ;
        RECT 231.000 197.800 231.400 198.200 ;
        RECT 229.400 193.800 229.800 194.200 ;
        RECT 229.400 188.200 229.700 193.800 ;
        RECT 230.200 193.100 230.600 195.900 ;
        RECT 231.000 194.200 231.300 197.800 ;
        RECT 232.600 196.100 233.000 196.200 ;
        RECT 233.400 196.100 233.800 196.200 ;
        RECT 232.600 195.800 233.800 196.100 ;
        RECT 231.800 194.800 232.200 195.200 ;
        RECT 233.400 194.800 233.800 195.200 ;
        RECT 231.000 193.800 231.400 194.200 ;
        RECT 231.800 191.200 232.100 194.800 ;
        RECT 233.400 194.200 233.700 194.800 ;
        RECT 233.400 193.800 233.800 194.200 ;
        RECT 233.400 192.100 233.800 192.200 ;
        RECT 234.200 192.100 234.600 192.200 ;
        RECT 236.600 192.100 237.000 197.900 ;
        RECT 238.200 195.100 238.600 195.200 ;
        RECT 239.000 195.100 239.400 195.200 ;
        RECT 238.200 194.800 239.400 195.100 ;
        RECT 240.600 192.800 241.000 193.200 ;
        RECT 233.400 191.800 234.600 192.100 ;
        RECT 231.800 190.800 232.200 191.200 ;
        RECT 229.400 187.800 229.800 188.200 ;
        RECT 225.400 186.800 225.800 187.200 ;
        RECT 228.600 186.800 229.000 187.200 ;
        RECT 230.200 186.800 230.600 187.200 ;
        RECT 228.600 186.200 228.900 186.800 ;
        RECT 223.800 185.800 224.200 186.200 ;
        RECT 224.600 185.800 225.000 186.200 ;
        RECT 226.200 185.800 226.600 186.200 ;
        RECT 228.600 185.800 229.000 186.200 ;
        RECT 223.800 181.200 224.100 185.800 ;
        RECT 224.600 185.200 224.900 185.800 ;
        RECT 226.200 185.200 226.500 185.800 ;
        RECT 224.600 184.800 225.000 185.200 ;
        RECT 226.200 184.800 226.600 185.200 ;
        RECT 227.800 185.100 228.200 185.200 ;
        RECT 228.600 185.100 229.000 185.200 ;
        RECT 227.800 184.800 229.000 185.100 ;
        RECT 223.800 180.800 224.200 181.200 ;
        RECT 226.200 180.200 226.500 184.800 ;
        RECT 230.200 183.200 230.500 186.800 ;
        RECT 231.000 185.100 231.400 187.900 ;
        RECT 230.200 182.800 230.600 183.200 ;
        RECT 232.600 183.100 233.000 188.900 ;
        RECT 233.400 188.800 233.800 189.200 ;
        RECT 233.400 188.200 233.700 188.800 ;
        RECT 233.400 187.800 233.800 188.200 ;
        RECT 233.400 186.800 233.800 187.200 ;
        RECT 233.400 186.300 233.700 186.800 ;
        RECT 233.400 185.900 233.800 186.300 ;
        RECT 237.400 183.100 237.800 188.900 ;
        RECT 240.600 187.200 240.900 192.800 ;
        RECT 241.400 192.100 241.800 197.900 ;
        RECT 243.000 197.200 243.300 201.800 ;
        RECT 243.800 201.200 244.100 204.800 ;
        RECT 243.800 200.800 244.200 201.200 ;
        RECT 243.000 196.800 243.400 197.200 ;
        RECT 243.800 196.100 244.200 196.200 ;
        RECT 244.600 196.100 245.000 196.200 ;
        RECT 243.000 193.100 243.400 195.900 ;
        RECT 243.800 195.800 245.000 196.100 ;
        RECT 245.400 195.200 245.700 215.800 ;
        RECT 247.800 214.700 248.200 215.100 ;
        RECT 247.000 213.800 247.400 214.200 ;
        RECT 246.200 208.800 246.600 209.200 ;
        RECT 246.200 208.200 246.500 208.800 ;
        RECT 246.200 207.800 246.600 208.200 ;
        RECT 247.000 206.200 247.300 213.800 ;
        RECT 247.800 211.100 248.100 214.700 ;
        RECT 248.600 212.100 249.000 217.900 ;
        RECT 249.400 213.800 249.800 214.200 ;
        RECT 247.800 210.800 248.900 211.100 ;
        RECT 248.600 209.200 248.900 210.800 ;
        RECT 249.400 210.200 249.700 213.800 ;
        RECT 250.200 213.100 250.600 215.900 ;
        RECT 249.400 209.800 249.800 210.200 ;
        RECT 248.600 208.800 249.000 209.200 ;
        RECT 248.600 208.100 249.000 208.200 ;
        RECT 249.400 208.100 249.800 208.200 ;
        RECT 248.600 207.800 249.800 208.100 ;
        RECT 247.800 206.800 248.200 207.200 ;
        RECT 247.000 205.800 247.400 206.200 ;
        RECT 247.000 205.200 247.300 205.800 ;
        RECT 247.000 204.800 247.400 205.200 ;
        RECT 247.000 202.800 247.400 203.200 ;
        RECT 247.000 195.200 247.300 202.800 ;
        RECT 245.400 194.800 245.800 195.200 ;
        RECT 247.000 194.800 247.400 195.200 ;
        RECT 243.800 191.800 244.200 192.200 ;
        RECT 240.600 186.800 241.000 187.200 ;
        RECT 239.000 183.100 239.400 183.200 ;
        RECT 239.800 183.100 240.200 183.200 ;
        RECT 239.000 182.800 240.200 183.100 ;
        RECT 226.200 179.800 226.600 180.200 ;
        RECT 225.400 175.800 225.800 176.200 ;
        RECT 225.400 175.200 225.700 175.800 ;
        RECT 230.200 175.200 230.500 182.800 ;
        RECT 232.600 181.800 233.000 182.200 ;
        RECT 231.000 180.800 231.400 181.200 ;
        RECT 222.200 174.800 222.600 175.200 ;
        RECT 224.600 174.800 225.000 175.200 ;
        RECT 225.400 174.800 225.800 175.200 ;
        RECT 226.200 174.800 226.600 175.200 ;
        RECT 227.000 174.800 227.400 175.200 ;
        RECT 230.200 174.800 230.600 175.200 ;
        RECT 221.400 173.800 221.800 174.200 ;
        RECT 221.400 173.200 221.700 173.800 ;
        RECT 224.600 173.200 224.900 174.800 ;
        RECT 226.200 174.200 226.500 174.800 ;
        RECT 226.200 173.800 226.600 174.200 ;
        RECT 221.400 172.800 221.800 173.200 ;
        RECT 224.600 172.800 225.000 173.200 ;
        RECT 227.000 172.200 227.300 174.800 ;
        RECT 231.000 174.200 231.300 180.800 ;
        RECT 231.800 174.800 232.200 175.200 ;
        RECT 231.000 173.800 231.400 174.200 ;
        RECT 227.800 173.100 228.200 173.200 ;
        RECT 228.600 173.100 229.000 173.200 ;
        RECT 227.800 172.800 229.000 173.100 ;
        RECT 227.000 171.800 227.400 172.200 ;
        RECT 231.800 169.200 232.100 174.800 ;
        RECT 217.400 165.800 217.800 166.200 ;
        RECT 218.200 165.800 218.600 166.200 ;
        RECT 217.400 164.200 217.700 165.800 ;
        RECT 217.400 163.800 217.800 164.200 ;
        RECT 219.800 163.100 220.200 168.900 ;
        RECT 221.400 167.800 221.800 168.200 ;
        RECT 221.400 166.200 221.700 167.800 ;
        RECT 221.400 165.800 221.800 166.200 ;
        RECT 224.600 163.100 225.000 168.900 ;
        RECT 231.800 168.800 232.200 169.200 ;
        RECT 225.400 166.800 225.800 167.200 ;
        RECT 225.400 166.200 225.700 166.800 ;
        RECT 225.400 165.800 225.800 166.200 ;
        RECT 226.200 165.100 226.600 167.900 ;
        RECT 227.800 161.800 228.200 162.200 ;
        RECT 216.600 159.800 217.000 160.200 ;
        RECT 214.200 159.100 214.600 159.200 ;
        RECT 215.000 159.100 215.400 159.200 ;
        RECT 214.200 158.800 215.400 159.100 ;
        RECT 207.000 157.800 207.400 158.200 ;
        RECT 207.000 157.200 207.300 157.800 ;
        RECT 205.400 157.100 205.800 157.200 ;
        RECT 206.200 157.100 206.600 157.200 ;
        RECT 205.400 156.800 206.600 157.100 ;
        RECT 207.000 156.800 207.400 157.200 ;
        RECT 204.600 153.800 205.000 154.200 ;
        RECT 207.800 152.100 208.200 157.900 ;
        RECT 209.400 155.100 209.800 155.200 ;
        RECT 210.200 155.100 210.600 155.200 ;
        RECT 209.400 154.800 210.600 155.100 ;
        RECT 212.600 152.100 213.000 157.900 ;
        RECT 213.400 157.800 213.800 158.200 ;
        RECT 216.600 157.200 216.900 159.800 ;
        RECT 216.600 156.800 217.000 157.200 ;
        RECT 213.400 154.800 213.800 155.200 ;
        RECT 213.400 154.200 213.700 154.800 ;
        RECT 213.400 153.800 213.800 154.200 ;
        RECT 214.200 153.100 214.600 155.900 ;
        RECT 217.400 152.100 217.800 157.900 ;
        RECT 220.600 155.800 221.000 156.200 ;
        RECT 220.600 155.200 220.900 155.800 ;
        RECT 220.600 154.800 221.000 155.200 ;
        RECT 222.200 152.100 222.600 157.900 ;
        RECT 223.000 154.800 223.400 155.200 ;
        RECT 223.000 154.200 223.300 154.800 ;
        RECT 223.000 153.800 223.400 154.200 ;
        RECT 223.800 153.100 224.200 155.900 ;
        RECT 227.800 155.200 228.100 161.800 ;
        RECT 231.800 156.800 232.200 157.200 ;
        RECT 227.800 154.800 228.200 155.200 ;
        RECT 231.800 154.200 232.100 156.800 ;
        RECT 232.600 156.200 232.900 181.800 ;
        RECT 240.600 179.200 240.900 186.800 ;
        RECT 233.400 178.800 233.800 179.200 ;
        RECT 240.600 178.800 241.000 179.200 ;
        RECT 233.400 167.200 233.700 178.800 ;
        RECT 237.400 176.800 237.800 177.200 ;
        RECT 237.400 176.200 237.700 176.800 ;
        RECT 234.200 175.800 234.600 176.200 ;
        RECT 237.400 175.800 237.800 176.200 ;
        RECT 234.200 175.200 234.500 175.800 ;
        RECT 234.200 174.800 234.600 175.200 ;
        RECT 235.000 174.800 235.400 175.200 ;
        RECT 235.000 174.200 235.300 174.800 ;
        RECT 235.000 173.800 235.400 174.200 ;
        RECT 235.800 173.800 236.200 174.200 ;
        RECT 235.800 169.200 236.100 173.800 ;
        RECT 236.600 171.800 237.000 172.200 ;
        RECT 236.600 171.200 236.900 171.800 ;
        RECT 236.600 170.800 237.000 171.200 ;
        RECT 237.400 170.200 237.700 175.800 ;
        RECT 238.200 172.100 238.600 172.200 ;
        RECT 239.000 172.100 239.400 172.200 ;
        RECT 240.600 172.100 241.000 177.900 ;
        RECT 242.200 174.800 242.600 175.200 ;
        RECT 238.200 171.800 239.400 172.100 ;
        RECT 237.400 169.800 237.800 170.200 ;
        RECT 234.200 169.100 234.600 169.200 ;
        RECT 235.000 169.100 235.400 169.200 ;
        RECT 234.200 168.800 235.400 169.100 ;
        RECT 235.800 168.800 236.200 169.200 ;
        RECT 233.400 166.800 233.800 167.200 ;
        RECT 236.600 163.100 237.000 168.900 ;
        RECT 237.400 167.800 237.800 168.200 ;
        RECT 240.600 167.800 241.000 168.200 ;
        RECT 237.400 167.200 237.700 167.800 ;
        RECT 237.400 166.800 237.800 167.200 ;
        RECT 240.600 166.300 240.900 167.800 ;
        RECT 240.600 165.900 241.000 166.300 ;
        RECT 241.400 163.100 241.800 168.900 ;
        RECT 242.200 167.200 242.500 174.800 ;
        RECT 242.200 166.800 242.600 167.200 ;
        RECT 236.600 161.800 237.000 162.200 ;
        RECT 236.600 157.200 236.900 161.800 ;
        RECT 236.600 156.800 237.000 157.200 ;
        RECT 232.600 155.800 233.000 156.200 ;
        RECT 234.200 156.100 234.600 156.200 ;
        RECT 235.000 156.100 235.400 156.200 ;
        RECT 234.200 155.800 235.400 156.100 ;
        RECT 232.600 155.200 232.900 155.800 ;
        RECT 232.600 154.800 233.000 155.200 ;
        RECT 235.000 154.800 235.400 155.200 ;
        RECT 231.800 153.800 232.200 154.200 ;
        RECT 230.200 151.800 230.600 152.200 ;
        RECT 208.600 148.800 209.000 149.200 ;
        RECT 219.800 149.100 220.200 149.200 ;
        RECT 220.600 149.100 221.000 149.200 ;
        RECT 205.400 148.100 205.800 148.200 ;
        RECT 206.200 148.100 206.600 148.200 ;
        RECT 205.400 147.800 206.600 148.100 ;
        RECT 208.600 147.200 208.900 148.800 ;
        RECT 207.000 146.800 207.400 147.200 ;
        RECT 208.600 146.800 209.000 147.200 ;
        RECT 207.000 146.200 207.300 146.800 ;
        RECT 197.400 145.800 197.800 146.200 ;
        RECT 201.400 145.800 201.800 146.200 ;
        RECT 203.800 145.800 204.200 146.200 ;
        RECT 204.600 145.800 205.000 146.200 ;
        RECT 207.000 145.800 207.400 146.200 ;
        RECT 197.400 145.200 197.700 145.800 ;
        RECT 197.400 144.800 197.800 145.200 ;
        RECT 199.000 145.100 199.400 145.200 ;
        RECT 199.800 145.100 200.200 145.200 ;
        RECT 199.000 144.800 200.200 145.100 ;
        RECT 197.400 139.200 197.700 144.800 ;
        RECT 197.400 138.800 197.800 139.200 ;
        RECT 201.400 137.200 201.700 145.800 ;
        RECT 203.800 143.200 204.100 145.800 ;
        RECT 204.600 145.200 204.900 145.800 ;
        RECT 204.600 144.800 205.000 145.200 ;
        RECT 203.800 142.800 204.200 143.200 ;
        RECT 211.000 143.100 211.400 148.900 ;
        RECT 213.400 146.100 213.800 146.200 ;
        RECT 214.200 146.100 214.600 146.200 ;
        RECT 213.400 145.800 214.600 146.100 ;
        RECT 215.800 143.100 216.200 148.900 ;
        RECT 219.800 148.800 221.000 149.100 ;
        RECT 223.000 148.800 223.400 149.200 ;
        RECT 227.800 149.100 228.200 149.200 ;
        RECT 228.600 149.100 229.000 149.200 ;
        RECT 227.800 148.800 229.000 149.100 ;
        RECT 216.600 146.800 217.000 147.200 ;
        RECT 216.600 145.200 216.900 146.800 ;
        RECT 216.600 144.800 217.000 145.200 ;
        RECT 217.400 145.100 217.800 147.900 ;
        RECT 219.000 147.800 219.400 148.200 ;
        RECT 219.000 146.200 219.300 147.800 ;
        RECT 223.000 147.200 223.300 148.800 ;
        RECT 221.400 146.800 221.800 147.200 ;
        RECT 223.000 146.800 223.400 147.200 ;
        RECT 227.800 147.100 228.200 147.200 ;
        RECT 228.600 147.100 229.000 147.200 ;
        RECT 227.800 146.800 229.000 147.100 ;
        RECT 221.400 146.200 221.700 146.800 ;
        RECT 223.000 146.200 223.300 146.800 ;
        RECT 230.200 146.200 230.500 151.800 ;
        RECT 219.000 145.800 219.400 146.200 ;
        RECT 221.400 145.800 221.800 146.200 ;
        RECT 222.200 145.800 222.600 146.200 ;
        RECT 223.000 145.800 223.400 146.200 ;
        RECT 224.600 145.800 225.000 146.200 ;
        RECT 227.800 146.100 228.200 146.200 ;
        RECT 228.600 146.100 229.000 146.200 ;
        RECT 227.800 145.800 229.000 146.100 ;
        RECT 230.200 145.800 230.600 146.200 ;
        RECT 222.200 145.200 222.500 145.800 ;
        RECT 224.600 145.200 224.900 145.800 ;
        RECT 219.000 144.800 219.400 145.200 ;
        RECT 222.200 144.800 222.600 145.200 ;
        RECT 224.600 144.800 225.000 145.200 ;
        RECT 227.000 145.100 227.400 145.200 ;
        RECT 227.800 145.100 228.200 145.200 ;
        RECT 227.000 144.800 228.200 145.100 ;
        RECT 201.400 136.800 201.800 137.200 ;
        RECT 197.400 136.100 197.800 136.200 ;
        RECT 198.200 136.100 198.600 136.200 ;
        RECT 197.400 135.800 198.600 136.100 ;
        RECT 198.200 134.800 198.600 135.200 ;
        RECT 198.200 134.200 198.500 134.800 ;
        RECT 201.400 134.200 201.700 136.800 ;
        RECT 198.200 133.800 198.600 134.200 ;
        RECT 201.400 133.800 201.800 134.200 ;
        RECT 200.600 129.100 201.000 129.200 ;
        RECT 201.400 129.100 201.800 129.200 ;
        RECT 200.600 128.800 201.800 129.100 ;
        RECT 197.400 127.800 197.800 128.200 ;
        RECT 197.400 126.200 197.700 127.800 ;
        RECT 197.400 125.800 197.800 126.200 ;
        RECT 198.200 125.800 198.600 126.200 ;
        RECT 198.200 121.200 198.500 125.800 ;
        RECT 202.200 123.800 202.600 124.200 ;
        RECT 202.200 122.200 202.500 123.800 ;
        RECT 203.000 123.100 203.400 128.900 ;
        RECT 202.200 121.800 202.600 122.200 ;
        RECT 203.800 121.200 204.100 142.800 ;
        RECT 213.400 140.800 213.800 141.200 ;
        RECT 215.800 140.800 216.200 141.200 ;
        RECT 204.600 132.100 205.000 137.900 ;
        RECT 207.000 135.100 207.400 135.200 ;
        RECT 207.800 135.100 208.200 135.200 ;
        RECT 207.000 134.800 208.200 135.100 ;
        RECT 207.000 133.800 207.400 134.200 ;
        RECT 206.200 130.800 206.600 131.200 ;
        RECT 198.200 120.800 198.600 121.200 ;
        RECT 203.800 120.800 204.200 121.200 ;
        RECT 195.800 114.800 196.900 115.100 ;
        RECT 193.400 113.200 193.700 114.800 ;
        RECT 195.000 114.100 195.400 114.200 ;
        RECT 195.800 114.100 196.200 114.200 ;
        RECT 195.000 113.800 196.200 114.100 ;
        RECT 193.400 112.800 193.800 113.200 ;
        RECT 197.400 112.800 197.800 113.200 ;
        RECT 197.400 111.200 197.700 112.800 ;
        RECT 199.000 112.100 199.400 112.200 ;
        RECT 199.800 112.100 200.200 112.200 ;
        RECT 202.200 112.100 202.600 117.900 ;
        RECT 203.800 114.800 204.200 115.200 ;
        RECT 203.800 114.200 204.100 114.800 ;
        RECT 206.200 114.200 206.500 130.800 ;
        RECT 207.000 128.200 207.300 133.800 ;
        RECT 209.400 132.100 209.800 137.900 ;
        RECT 211.800 136.800 212.200 137.200 ;
        RECT 210.200 135.800 210.600 136.200 ;
        RECT 210.200 134.200 210.500 135.800 ;
        RECT 210.200 133.800 210.600 134.200 ;
        RECT 211.000 133.100 211.400 135.900 ;
        RECT 211.800 134.200 212.100 136.800 ;
        RECT 213.400 136.200 213.700 140.800 ;
        RECT 213.400 135.800 213.800 136.200 ;
        RECT 215.800 135.200 216.100 140.800 ;
        RECT 219.000 137.200 219.300 144.800 ;
        RECT 216.600 137.100 217.000 137.200 ;
        RECT 217.400 137.100 217.800 137.200 ;
        RECT 216.600 136.800 217.800 137.100 ;
        RECT 219.000 136.800 219.400 137.200 ;
        RECT 214.200 135.100 214.600 135.200 ;
        RECT 215.000 135.100 215.400 135.200 ;
        RECT 214.200 134.800 215.400 135.100 ;
        RECT 215.800 134.800 216.200 135.200 ;
        RECT 211.800 133.800 212.200 134.200 ;
        RECT 215.000 133.800 215.400 134.200 ;
        RECT 216.600 134.100 217.000 134.200 ;
        RECT 217.400 134.100 217.800 134.200 ;
        RECT 216.600 133.800 217.800 134.100 ;
        RECT 215.000 129.200 215.300 133.800 ;
        RECT 219.800 132.100 220.200 137.900 ;
        RECT 222.200 135.100 222.600 135.200 ;
        RECT 223.000 135.100 223.400 135.200 ;
        RECT 222.200 134.800 223.400 135.100 ;
        RECT 224.600 132.100 225.000 137.900 ;
        RECT 225.400 133.800 225.800 134.200 ;
        RECT 225.400 131.200 225.700 133.800 ;
        RECT 226.200 133.100 226.600 135.900 ;
        RECT 227.000 131.800 227.400 132.200 ;
        RECT 229.400 132.100 229.800 137.900 ;
        RECT 230.200 136.200 230.500 145.800 ;
        RECT 231.000 143.100 231.400 148.900 ;
        RECT 231.800 146.800 232.200 147.200 ;
        RECT 231.800 146.200 232.100 146.800 ;
        RECT 231.800 145.800 232.200 146.200 ;
        RECT 230.200 135.800 230.600 136.200 ;
        RECT 230.200 135.200 230.500 135.800 ;
        RECT 230.200 134.800 230.600 135.200 ;
        RECT 225.400 130.800 225.800 131.200 ;
        RECT 227.000 130.200 227.300 131.800 ;
        RECT 216.600 129.800 217.000 130.200 ;
        RECT 227.000 129.800 227.400 130.200 ;
        RECT 207.000 127.800 207.400 128.200 ;
        RECT 207.000 126.800 207.400 127.200 ;
        RECT 207.000 126.300 207.300 126.800 ;
        RECT 207.000 125.900 207.400 126.300 ;
        RECT 207.800 123.100 208.200 128.900 ;
        RECT 210.200 128.800 210.600 129.200 ;
        RECT 215.000 128.800 215.400 129.200 ;
        RECT 208.600 126.800 209.000 127.200 ;
        RECT 203.800 113.800 204.200 114.200 ;
        RECT 206.200 113.800 206.600 114.200 ;
        RECT 207.000 112.100 207.400 117.900 ;
        RECT 208.600 117.200 208.900 126.800 ;
        RECT 209.400 125.100 209.800 127.900 ;
        RECT 210.200 127.200 210.500 128.800 ;
        RECT 215.000 127.200 215.300 128.800 ;
        RECT 210.200 126.800 210.600 127.200 ;
        RECT 211.800 126.800 212.200 127.200 ;
        RECT 215.000 126.800 215.400 127.200 ;
        RECT 211.800 126.200 212.100 126.800 ;
        RECT 216.600 126.200 216.900 129.800 ;
        RECT 225.400 128.800 225.800 129.200 ;
        RECT 217.400 128.100 217.800 128.200 ;
        RECT 218.200 128.100 218.600 128.200 ;
        RECT 217.400 127.800 218.600 128.100 ;
        RECT 225.400 127.200 225.700 128.800 ;
        RECT 222.200 126.800 222.600 127.200 ;
        RECT 224.600 126.800 225.000 127.200 ;
        RECT 225.400 127.100 225.800 127.200 ;
        RECT 226.200 127.100 226.600 127.200 ;
        RECT 225.400 126.800 226.600 127.100 ;
        RECT 222.200 126.200 222.500 126.800 ;
        RECT 224.600 126.200 224.900 126.800 ;
        RECT 211.800 125.800 212.200 126.200 ;
        RECT 214.200 125.800 214.600 126.200 ;
        RECT 215.800 125.800 216.200 126.200 ;
        RECT 216.600 125.800 217.000 126.200 ;
        RECT 219.000 126.100 219.400 126.200 ;
        RECT 219.800 126.100 220.200 126.200 ;
        RECT 219.000 125.800 220.200 126.100 ;
        RECT 222.200 125.800 222.600 126.200 ;
        RECT 224.600 125.800 225.000 126.200 ;
        RECT 226.200 125.800 226.600 126.200 ;
        RECT 214.200 125.200 214.500 125.800 ;
        RECT 211.800 125.100 212.200 125.200 ;
        RECT 212.600 125.100 213.000 125.200 ;
        RECT 211.800 124.800 213.000 125.100 ;
        RECT 214.200 124.800 214.600 125.200 ;
        RECT 215.800 124.200 216.100 125.800 ;
        RECT 219.800 125.100 220.200 125.200 ;
        RECT 220.600 125.100 221.000 125.200 ;
        RECT 219.800 124.800 221.000 125.100 ;
        RECT 224.600 124.800 225.000 125.200 ;
        RECT 224.600 124.200 224.900 124.800 ;
        RECT 226.200 124.200 226.500 125.800 ;
        RECT 215.800 123.800 216.200 124.200 ;
        RECT 224.600 123.800 225.000 124.200 ;
        RECT 226.200 123.800 226.600 124.200 ;
        RECT 228.600 123.100 229.000 128.900 ;
        RECT 231.800 125.800 232.200 126.200 ;
        RECT 231.800 125.200 232.100 125.800 ;
        RECT 231.800 124.800 232.200 125.200 ;
        RECT 230.200 120.800 230.600 121.200 ;
        RECT 224.600 119.800 225.000 120.200 ;
        RECT 208.600 116.800 209.000 117.200 ;
        RECT 210.200 116.800 210.600 117.200 ;
        RECT 208.600 113.100 209.000 115.900 ;
        RECT 209.400 113.100 209.800 115.900 ;
        RECT 210.200 114.200 210.500 116.800 ;
        RECT 210.200 113.800 210.600 114.200 ;
        RECT 211.000 112.100 211.400 117.900 ;
        RECT 212.600 115.800 213.000 116.200 ;
        RECT 212.600 115.200 212.900 115.800 ;
        RECT 212.600 114.800 213.000 115.200 ;
        RECT 215.000 113.800 215.400 114.200 ;
        RECT 199.000 111.800 200.200 112.100 ;
        RECT 197.400 110.800 197.800 111.200 ;
        RECT 209.400 110.800 209.800 111.200 ;
        RECT 194.200 109.800 194.600 110.200 ;
        RECT 194.200 106.200 194.500 109.800 ;
        RECT 194.200 105.800 194.600 106.200 ;
        RECT 196.600 103.100 197.000 108.900 ;
        RECT 197.400 107.200 197.700 110.800 ;
        RECT 203.000 108.800 203.400 109.200 ;
        RECT 197.400 106.800 197.800 107.200 ;
        RECT 198.200 105.100 198.600 107.900 ;
        RECT 200.600 107.800 202.500 108.100 ;
        RECT 199.800 107.100 200.200 107.200 ;
        RECT 200.600 107.100 200.900 107.800 ;
        RECT 202.200 107.200 202.500 107.800 ;
        RECT 199.800 106.800 200.900 107.100 ;
        RECT 201.400 106.800 201.800 107.200 ;
        RECT 202.200 106.800 202.600 107.200 ;
        RECT 201.400 106.200 201.700 106.800 ;
        RECT 203.000 106.200 203.300 108.800 ;
        RECT 209.400 107.200 209.700 110.800 ;
        RECT 209.400 106.800 209.800 107.200 ;
        RECT 210.200 106.800 210.600 107.200 ;
        RECT 211.800 106.800 212.200 107.200 ;
        RECT 199.000 106.100 199.400 106.200 ;
        RECT 199.800 106.100 200.200 106.200 ;
        RECT 199.000 105.800 200.200 106.100 ;
        RECT 200.600 105.800 201.000 106.200 ;
        RECT 201.400 105.800 201.800 106.200 ;
        RECT 203.000 105.800 203.400 106.200 ;
        RECT 205.400 105.800 205.800 106.200 ;
        RECT 207.800 105.800 208.200 106.200 ;
        RECT 208.600 105.800 209.000 106.200 ;
        RECT 193.400 97.800 193.800 98.200 ;
        RECT 193.400 95.200 193.700 97.800 ;
        RECT 193.400 94.800 193.800 95.200 ;
        RECT 194.200 93.800 194.600 94.200 ;
        RECT 195.800 93.800 196.200 94.200 ;
        RECT 194.200 87.200 194.500 93.800 ;
        RECT 195.000 91.800 195.400 92.200 ;
        RECT 195.000 87.200 195.300 91.800 ;
        RECT 195.800 89.200 196.100 93.800 ;
        RECT 197.400 92.100 197.800 97.900 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 198.200 91.200 198.500 94.800 ;
        RECT 198.200 90.800 198.600 91.200 ;
        RECT 195.800 88.800 196.200 89.200 ;
        RECT 196.600 88.800 197.000 89.200 ;
        RECT 194.200 86.800 194.600 87.200 ;
        RECT 195.000 86.800 195.400 87.200 ;
        RECT 196.600 85.200 196.900 88.800 ;
        RECT 197.400 86.800 197.800 87.200 ;
        RECT 197.400 86.200 197.700 86.800 ;
        RECT 197.400 85.800 197.800 86.200 ;
        RECT 192.600 84.800 193.000 85.200 ;
        RECT 196.600 84.800 197.000 85.200 ;
        RECT 199.000 84.800 199.400 85.200 ;
        RECT 192.600 81.800 193.000 82.200 ;
        RECT 192.600 75.200 192.900 81.800 ;
        RECT 199.000 81.200 199.300 84.800 ;
        RECT 194.200 80.800 194.600 81.200 ;
        RECT 197.400 80.800 197.800 81.200 ;
        RECT 199.000 80.800 199.400 81.200 ;
        RECT 193.400 77.800 193.800 78.200 ;
        RECT 192.600 74.800 193.000 75.200 ;
        RECT 193.400 74.200 193.700 77.800 ;
        RECT 194.200 75.200 194.500 80.800 ;
        RECT 195.000 76.800 195.400 77.200 ;
        RECT 195.000 76.200 195.300 76.800 ;
        RECT 197.400 76.200 197.700 80.800 ;
        RECT 195.000 75.800 195.400 76.200 ;
        RECT 197.400 75.800 197.800 76.200 ;
        RECT 194.200 74.800 194.600 75.200 ;
        RECT 197.400 74.800 197.800 75.200 ;
        RECT 199.800 75.100 200.100 105.800 ;
        RECT 200.600 104.200 200.900 105.800 ;
        RECT 200.600 103.800 201.000 104.200 ;
        RECT 205.400 103.200 205.700 105.800 ;
        RECT 207.800 105.200 208.100 105.800 ;
        RECT 207.800 104.800 208.200 105.200 ;
        RECT 208.600 104.200 208.900 105.800 ;
        RECT 208.600 103.800 209.000 104.200 ;
        RECT 205.400 102.800 205.800 103.200 ;
        RECT 209.400 102.200 209.700 106.800 ;
        RECT 210.200 106.200 210.500 106.800 ;
        RECT 211.800 106.200 212.100 106.800 ;
        RECT 210.200 105.800 210.600 106.200 ;
        RECT 211.800 105.800 212.200 106.200 ;
        RECT 209.400 101.800 209.800 102.200 ;
        RECT 207.800 100.800 208.200 101.200 ;
        RECT 200.600 95.100 201.000 95.200 ;
        RECT 200.600 94.800 201.800 95.100 ;
        RECT 201.400 94.700 201.800 94.800 ;
        RECT 202.200 92.100 202.600 97.900 ;
        RECT 205.400 96.800 205.800 97.200 ;
        RECT 203.800 93.100 204.200 95.900 ;
        RECT 204.600 95.800 205.000 96.200 ;
        RECT 204.600 95.200 204.900 95.800 ;
        RECT 204.600 94.800 205.000 95.200 ;
        RECT 203.800 91.800 204.200 92.200 ;
        RECT 202.200 87.100 202.600 87.200 ;
        RECT 203.000 87.100 203.400 87.200 ;
        RECT 202.200 86.800 203.400 87.100 ;
        RECT 203.000 85.800 203.400 86.200 ;
        RECT 201.400 85.100 201.800 85.200 ;
        RECT 202.200 85.100 202.600 85.200 ;
        RECT 201.400 84.800 202.600 85.100 ;
        RECT 203.000 81.200 203.300 85.800 ;
        RECT 203.000 80.800 203.400 81.200 ;
        RECT 200.600 79.100 201.000 79.200 ;
        RECT 201.400 79.100 201.800 79.200 ;
        RECT 200.600 78.800 201.800 79.100 ;
        RECT 201.400 76.100 201.800 76.200 ;
        RECT 202.200 76.100 202.600 76.200 ;
        RECT 201.400 75.800 202.600 76.100 ;
        RECT 203.800 75.200 204.100 91.800 ;
        RECT 204.600 88.800 205.000 89.200 ;
        RECT 204.600 86.200 204.900 88.800 ;
        RECT 205.400 88.100 205.700 96.800 ;
        RECT 206.200 95.800 206.600 96.200 ;
        RECT 206.200 94.200 206.500 95.800 ;
        RECT 207.800 95.200 208.100 100.800 ;
        RECT 210.200 100.200 210.500 105.800 ;
        RECT 211.000 105.100 211.400 105.200 ;
        RECT 211.800 105.100 212.200 105.200 ;
        RECT 212.600 105.100 213.000 107.900 ;
        RECT 211.000 104.800 212.200 105.100 ;
        RECT 211.000 102.800 211.400 103.200 ;
        RECT 214.200 103.100 214.600 108.900 ;
        RECT 215.000 108.200 215.300 113.800 ;
        RECT 215.800 112.100 216.200 117.900 ;
        RECT 219.800 116.800 220.200 117.200 ;
        RECT 219.800 116.200 220.100 116.800 ;
        RECT 219.800 115.800 220.200 116.200 ;
        RECT 221.400 115.800 221.800 116.200 ;
        RECT 219.800 115.100 220.200 115.200 ;
        RECT 220.600 115.100 221.000 115.200 ;
        RECT 219.800 114.800 221.000 115.100 ;
        RECT 219.000 114.100 219.400 114.200 ;
        RECT 219.800 114.100 220.200 114.200 ;
        RECT 219.000 113.800 220.200 114.100 ;
        RECT 218.200 111.800 218.600 112.200 ;
        RECT 215.000 107.800 215.400 108.200 ;
        RECT 218.200 107.200 218.500 111.800 ;
        RECT 219.000 111.200 219.300 113.800 ;
        RECT 221.400 113.100 221.700 115.800 ;
        RECT 224.600 115.200 224.900 119.800 ;
        RECT 225.400 116.800 225.800 117.200 ;
        RECT 225.400 115.200 225.700 116.800 ;
        RECT 230.200 115.200 230.500 120.800 ;
        RECT 231.000 115.800 231.400 116.200 ;
        RECT 231.000 115.200 231.300 115.800 ;
        RECT 232.600 115.200 232.900 154.800 ;
        RECT 235.000 154.200 235.300 154.800 ;
        RECT 236.600 154.200 236.900 156.800 ;
        RECT 235.000 153.800 235.400 154.200 ;
        RECT 236.600 153.800 237.000 154.200 ;
        RECT 239.800 152.100 240.200 157.900 ;
        RECT 234.200 145.800 234.600 146.200 ;
        RECT 234.200 145.200 234.500 145.800 ;
        RECT 234.200 144.800 234.600 145.200 ;
        RECT 235.800 143.100 236.200 148.900 ;
        RECT 237.400 145.100 237.800 147.900 ;
        RECT 238.200 146.800 238.600 147.200 ;
        RECT 239.000 146.800 239.400 147.200 ;
        RECT 240.600 146.800 241.000 147.200 ;
        RECT 238.200 143.200 238.500 146.800 ;
        RECT 239.000 146.200 239.300 146.800 ;
        RECT 240.600 146.200 240.900 146.800 ;
        RECT 239.000 145.800 239.400 146.200 ;
        RECT 240.600 145.800 241.000 146.200 ;
        RECT 239.800 145.100 240.200 145.200 ;
        RECT 240.600 145.100 241.000 145.200 ;
        RECT 241.400 145.100 241.800 147.900 ;
        RECT 239.800 144.800 241.000 145.100 ;
        RECT 239.800 143.800 240.200 144.200 ;
        RECT 238.200 142.800 238.600 143.200 ;
        RECT 233.400 134.700 233.800 135.100 ;
        RECT 233.400 134.200 233.700 134.700 ;
        RECT 233.400 133.800 233.800 134.200 ;
        RECT 234.200 132.100 234.600 137.900 ;
        RECT 235.800 133.100 236.200 135.900 ;
        RECT 236.600 135.800 237.000 136.200 ;
        RECT 238.200 135.800 238.600 136.200 ;
        RECT 234.200 130.800 234.600 131.200 ;
        RECT 233.400 123.100 233.800 128.900 ;
        RECT 234.200 127.200 234.500 130.800 ;
        RECT 235.800 129.800 236.200 130.200 ;
        RECT 234.200 126.800 234.600 127.200 ;
        RECT 235.000 125.100 235.400 127.900 ;
        RECT 235.800 127.200 236.100 129.800 ;
        RECT 236.600 129.200 236.900 135.800 ;
        RECT 238.200 135.200 238.500 135.800 ;
        RECT 237.400 134.800 237.800 135.200 ;
        RECT 238.200 134.800 238.600 135.200 ;
        RECT 237.400 134.200 237.700 134.800 ;
        RECT 237.400 133.800 237.800 134.200 ;
        RECT 236.600 128.800 237.000 129.200 ;
        RECT 235.800 126.800 236.200 127.200 ;
        RECT 238.200 127.100 238.500 134.800 ;
        RECT 237.400 126.800 238.500 127.100 ;
        RECT 239.000 126.800 239.400 127.200 ;
        RECT 237.400 125.200 237.700 126.800 ;
        RECT 238.200 125.800 238.600 126.200 ;
        RECT 238.200 125.200 238.500 125.800 ;
        RECT 239.000 125.200 239.300 126.800 ;
        RECT 237.400 124.800 237.800 125.200 ;
        RECT 238.200 124.800 238.600 125.200 ;
        RECT 239.000 124.800 239.400 125.200 ;
        RECT 235.000 119.800 235.400 120.200 ;
        RECT 235.000 115.200 235.300 119.800 ;
        RECT 239.000 119.200 239.300 124.800 ;
        RECT 239.000 118.800 239.400 119.200 ;
        RECT 238.200 117.800 238.600 118.200 ;
        RECT 239.000 118.100 239.400 118.200 ;
        RECT 239.800 118.100 240.100 143.800 ;
        RECT 240.600 142.800 241.000 143.200 ;
        RECT 240.600 139.200 240.900 142.800 ;
        RECT 242.200 142.100 242.500 166.800 ;
        RECT 243.000 165.100 243.400 167.900 ;
        RECT 243.000 154.800 243.400 155.200 ;
        RECT 243.000 154.200 243.300 154.800 ;
        RECT 243.000 153.800 243.400 154.200 ;
        RECT 243.800 149.200 244.100 191.800 ;
        RECT 245.400 182.200 245.700 194.800 ;
        RECT 246.200 193.800 246.600 194.200 ;
        RECT 246.200 193.200 246.500 193.800 ;
        RECT 246.200 192.800 246.600 193.200 ;
        RECT 247.000 188.200 247.300 194.800 ;
        RECT 247.000 187.800 247.400 188.200 ;
        RECT 247.800 182.200 248.100 206.800 ;
        RECT 248.600 205.800 249.000 206.200 ;
        RECT 248.600 199.200 248.900 205.800 ;
        RECT 248.600 198.800 249.000 199.200 ;
        RECT 248.600 198.200 248.900 198.800 ;
        RECT 248.600 197.800 249.000 198.200 ;
        RECT 250.200 187.800 250.600 188.200 ;
        RECT 250.200 186.200 250.500 187.800 ;
        RECT 250.200 185.800 250.600 186.200 ;
        RECT 245.400 181.800 245.800 182.200 ;
        RECT 247.800 181.800 248.200 182.200 ;
        RECT 248.600 181.800 249.000 182.200 ;
        RECT 248.600 178.100 248.900 181.800 ;
        RECT 244.600 175.800 245.000 176.200 ;
        RECT 244.600 175.100 244.900 175.800 ;
        RECT 244.600 174.700 245.000 175.100 ;
        RECT 245.400 172.100 245.800 177.900 ;
        RECT 248.600 177.800 249.700 178.100 ;
        RECT 248.600 176.800 249.000 177.200 ;
        RECT 248.600 176.200 248.900 176.800 ;
        RECT 247.000 173.100 247.400 175.900 ;
        RECT 248.600 175.800 249.000 176.200 ;
        RECT 247.800 175.100 248.200 175.200 ;
        RECT 248.600 175.100 249.000 175.200 ;
        RECT 247.800 174.800 249.000 175.100 ;
        RECT 247.800 173.800 248.200 174.200 ;
        RECT 247.800 173.200 248.100 173.800 ;
        RECT 249.400 173.200 249.700 177.800 ;
        RECT 250.200 175.800 250.600 176.200 ;
        RECT 250.200 175.200 250.500 175.800 ;
        RECT 250.200 174.800 250.600 175.200 ;
        RECT 247.800 172.800 248.200 173.200 ;
        RECT 249.400 172.800 249.800 173.200 ;
        RECT 246.200 170.800 246.600 171.200 ;
        RECT 246.200 167.100 246.500 170.800 ;
        RECT 248.600 169.800 249.000 170.200 ;
        RECT 247.000 168.800 247.400 169.200 ;
        RECT 247.000 168.200 247.300 168.800 ;
        RECT 247.000 167.800 247.400 168.200 ;
        RECT 246.200 166.800 247.300 167.100 ;
        RECT 246.200 165.800 246.600 166.200 ;
        RECT 244.600 161.800 245.000 162.200 ;
        RECT 244.600 161.200 244.900 161.800 ;
        RECT 244.600 160.800 245.000 161.200 ;
        RECT 246.200 158.200 246.500 165.800 ;
        RECT 247.000 165.200 247.300 166.800 ;
        RECT 248.600 166.200 248.900 169.800 ;
        RECT 249.400 167.200 249.700 172.800 ;
        RECT 249.400 166.800 249.800 167.200 ;
        RECT 248.600 165.800 249.000 166.200 ;
        RECT 247.000 164.800 247.400 165.200 ;
        RECT 244.600 152.100 245.000 157.900 ;
        RECT 246.200 157.800 246.600 158.200 ;
        RECT 249.400 157.200 249.700 166.800 ;
        RECT 249.400 156.800 249.800 157.200 ;
        RECT 245.400 153.800 245.800 154.200 ;
        RECT 243.000 143.100 243.400 148.900 ;
        RECT 243.800 148.800 244.200 149.200 ;
        RECT 243.800 146.800 244.200 147.200 ;
        RECT 244.600 146.800 245.000 147.200 ;
        RECT 242.200 141.800 243.300 142.100 ;
        RECT 240.600 138.800 241.000 139.200 ;
        RECT 242.200 134.800 242.600 135.200 ;
        RECT 241.400 129.800 241.800 130.200 ;
        RECT 241.400 129.200 241.700 129.800 ;
        RECT 241.400 128.800 241.800 129.200 ;
        RECT 240.600 128.100 241.000 128.200 ;
        RECT 240.600 127.800 241.700 128.100 ;
        RECT 240.600 126.800 241.000 127.200 ;
        RECT 240.600 126.200 240.900 126.800 ;
        RECT 240.600 125.800 241.000 126.200 ;
        RECT 239.000 117.800 240.100 118.100 ;
        RECT 241.400 121.800 241.800 122.200 ;
        RECT 238.200 116.200 238.500 117.800 ;
        RECT 239.800 116.800 240.200 117.200 ;
        RECT 239.800 116.200 240.100 116.800 ;
        RECT 238.200 115.800 238.600 116.200 ;
        RECT 239.800 115.800 240.200 116.200 ;
        RECT 222.200 114.800 222.600 115.200 ;
        RECT 224.600 114.800 225.000 115.200 ;
        RECT 225.400 114.800 225.800 115.200 ;
        RECT 226.200 114.800 226.600 115.200 ;
        RECT 228.600 114.800 229.000 115.200 ;
        RECT 230.200 114.800 230.600 115.200 ;
        RECT 231.000 114.800 231.400 115.200 ;
        RECT 232.600 114.800 233.000 115.200 ;
        RECT 233.400 115.100 233.800 115.200 ;
        RECT 234.200 115.100 234.600 115.200 ;
        RECT 233.400 114.800 234.600 115.100 ;
        RECT 235.000 114.800 235.400 115.200 ;
        RECT 222.200 114.200 222.500 114.800 ;
        RECT 222.200 113.800 222.600 114.200 ;
        RECT 221.400 112.800 222.500 113.100 ;
        RECT 219.000 110.800 219.400 111.200 ;
        RECT 222.200 109.200 222.500 112.800 ;
        RECT 215.000 106.800 215.400 107.200 ;
        RECT 218.200 106.800 218.600 107.200 ;
        RECT 215.000 106.300 215.300 106.800 ;
        RECT 215.000 105.900 215.400 106.300 ;
        RECT 215.000 104.800 215.400 105.200 ;
        RECT 210.200 99.800 210.600 100.200 ;
        RECT 211.000 99.200 211.300 102.800 ;
        RECT 214.200 99.800 214.600 100.200 ;
        RECT 210.200 98.800 210.600 99.200 ;
        RECT 211.000 98.800 211.400 99.200 ;
        RECT 210.200 95.200 210.500 98.800 ;
        RECT 214.200 96.200 214.500 99.800 ;
        RECT 215.000 99.200 215.300 104.800 ;
        RECT 219.000 103.100 219.400 108.900 ;
        RECT 222.200 108.800 222.600 109.200 ;
        RECT 223.800 106.800 224.200 107.200 ;
        RECT 225.400 106.800 225.800 107.200 ;
        RECT 223.800 106.200 224.100 106.800 ;
        RECT 225.400 106.200 225.700 106.800 ;
        RECT 219.800 105.800 220.200 106.200 ;
        RECT 223.800 105.800 224.200 106.200 ;
        RECT 224.600 105.800 225.000 106.200 ;
        RECT 225.400 105.800 225.800 106.200 ;
        RECT 219.800 104.200 220.100 105.800 ;
        RECT 222.200 104.800 222.600 105.200 ;
        RECT 219.800 103.800 220.200 104.200 ;
        RECT 215.800 101.800 216.200 102.200 ;
        RECT 215.000 98.800 215.400 99.200 ;
        RECT 214.200 95.800 214.600 96.200 ;
        RECT 215.800 95.200 216.100 101.800 ;
        RECT 207.800 94.800 208.200 95.200 ;
        RECT 209.400 94.800 209.800 95.200 ;
        RECT 210.200 94.800 210.600 95.200 ;
        RECT 212.600 95.100 213.000 95.200 ;
        RECT 213.400 95.100 213.800 95.200 ;
        RECT 212.600 94.800 213.800 95.100 ;
        RECT 215.800 94.800 216.200 95.200 ;
        RECT 206.200 93.800 206.600 94.200 ;
        RECT 207.800 89.200 208.100 94.800 ;
        RECT 208.600 93.800 209.000 94.200 ;
        RECT 208.600 91.200 208.900 93.800 ;
        RECT 208.600 90.800 209.000 91.200 ;
        RECT 205.400 87.800 206.500 88.100 ;
        RECT 205.400 86.800 205.800 87.200 ;
        RECT 204.600 85.800 205.000 86.200 ;
        RECT 204.600 75.800 205.000 76.200 ;
        RECT 204.600 75.200 204.900 75.800 ;
        RECT 199.800 74.800 200.900 75.100 ;
        RECT 203.800 74.800 204.200 75.200 ;
        RECT 204.600 74.800 205.000 75.200 ;
        RECT 193.400 73.800 193.800 74.200 ;
        RECT 193.400 72.800 193.800 73.200 ;
        RECT 193.400 69.200 193.700 72.800 ;
        RECT 197.400 69.200 197.700 74.800 ;
        RECT 199.000 73.800 199.400 74.200 ;
        RECT 199.800 73.800 200.200 74.200 ;
        RECT 199.000 72.200 199.300 73.800 ;
        RECT 199.800 73.200 200.100 73.800 ;
        RECT 199.800 72.800 200.200 73.200 ;
        RECT 199.000 71.800 199.400 72.200 ;
        RECT 193.400 68.800 193.800 69.200 ;
        RECT 197.400 68.800 197.800 69.200 ;
        RECT 192.600 67.800 193.000 68.200 ;
        RECT 192.600 67.200 192.900 67.800 ;
        RECT 192.600 66.800 193.000 67.200 ;
        RECT 193.400 67.100 193.800 67.200 ;
        RECT 194.200 67.100 194.600 67.200 ;
        RECT 193.400 66.800 194.600 67.100 ;
        RECT 199.000 66.800 199.400 67.200 ;
        RECT 199.000 66.200 199.300 66.800 ;
        RECT 200.600 66.200 200.900 74.800 ;
        RECT 201.400 74.100 201.800 74.200 ;
        RECT 202.200 74.100 202.600 74.200 ;
        RECT 201.400 73.800 202.600 74.100 ;
        RECT 204.600 73.800 205.000 74.200 ;
        RECT 202.200 68.800 202.600 69.200 ;
        RECT 202.200 67.200 202.500 68.800 ;
        RECT 203.000 68.100 203.400 68.200 ;
        RECT 203.800 68.100 204.200 68.200 ;
        RECT 203.000 67.800 204.200 68.100 ;
        RECT 204.600 67.200 204.900 73.800 ;
        RECT 205.400 67.200 205.700 86.800 ;
        RECT 206.200 74.200 206.500 87.800 ;
        RECT 207.000 83.100 207.400 88.900 ;
        RECT 207.800 88.800 208.200 89.200 ;
        RECT 208.600 87.200 208.900 90.800 ;
        RECT 208.600 86.800 209.000 87.200 ;
        RECT 209.400 84.200 209.700 94.800 ;
        RECT 215.800 94.200 216.100 94.800 ;
        RECT 215.800 93.800 216.200 94.200 ;
        RECT 216.600 91.800 217.000 92.200 ;
        RECT 219.000 92.100 219.400 97.900 ;
        RECT 219.800 95.200 220.100 103.800 ;
        RECT 220.600 102.100 221.000 102.200 ;
        RECT 221.400 102.100 221.800 102.200 ;
        RECT 220.600 101.800 221.800 102.100 ;
        RECT 221.400 100.800 221.800 101.200 ;
        RECT 220.600 95.800 221.000 96.200 ;
        RECT 219.800 94.800 220.200 95.200 ;
        RECT 210.200 85.800 210.600 86.200 ;
        RECT 210.200 85.200 210.500 85.800 ;
        RECT 210.200 84.800 210.600 85.200 ;
        RECT 209.400 83.800 209.800 84.200 ;
        RECT 210.200 83.800 210.600 84.200 ;
        RECT 207.000 75.800 207.400 76.200 ;
        RECT 207.000 75.200 207.300 75.800 ;
        RECT 207.000 74.800 207.400 75.200 ;
        RECT 207.800 74.800 208.200 75.200 ;
        RECT 208.600 74.800 209.000 75.200 ;
        RECT 206.200 73.800 206.600 74.200 ;
        RECT 202.200 66.800 202.600 67.200 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 204.600 66.800 205.000 67.200 ;
        RECT 205.400 66.800 205.800 67.200 ;
        RECT 187.000 66.100 187.400 66.200 ;
        RECT 187.800 66.100 188.200 66.200 ;
        RECT 187.000 65.800 188.200 66.100 ;
        RECT 190.200 65.800 190.600 66.200 ;
        RECT 191.000 65.800 191.400 66.200 ;
        RECT 191.800 65.800 192.200 66.200 ;
        RECT 194.200 66.100 194.600 66.200 ;
        RECT 195.000 66.100 195.400 66.200 ;
        RECT 194.200 65.800 195.400 66.100 ;
        RECT 195.800 65.800 196.200 66.200 ;
        RECT 199.000 65.800 199.400 66.200 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 200.600 65.800 201.000 66.200 ;
        RECT 183.800 65.100 184.200 65.200 ;
        RECT 184.600 65.100 185.000 65.200 ;
        RECT 183.800 64.800 185.000 65.100 ;
        RECT 190.200 59.200 190.500 65.800 ;
        RECT 191.000 65.200 191.300 65.800 ;
        RECT 191.000 64.800 191.400 65.200 ;
        RECT 195.800 65.100 196.100 65.800 ;
        RECT 195.000 64.800 196.100 65.100 ;
        RECT 199.800 65.200 200.100 65.800 ;
        RECT 199.800 64.800 200.200 65.200 ;
        RECT 195.000 59.200 195.300 64.800 ;
        RECT 188.600 58.800 189.000 59.200 ;
        RECT 190.200 58.800 190.600 59.200 ;
        RECT 195.000 58.800 195.400 59.200 ;
        RECT 174.200 53.800 174.600 54.200 ;
        RECT 173.400 51.800 173.800 52.200 ;
        RECT 175.000 52.100 175.400 57.900 ;
        RECT 175.800 57.800 176.200 58.200 ;
        RECT 175.800 54.200 176.100 57.800 ;
        RECT 175.800 53.800 176.200 54.200 ;
        RECT 175.800 49.200 176.100 53.800 ;
        RECT 176.600 53.100 177.000 55.900 ;
        RECT 177.400 53.100 177.800 55.900 ;
        RECT 179.000 52.100 179.400 57.900 ;
        RECT 182.200 54.800 182.600 55.200 ;
        RECT 182.200 54.200 182.500 54.800 ;
        RECT 180.600 53.800 181.000 54.200 ;
        RECT 182.200 53.800 182.600 54.200 ;
        RECT 175.800 48.800 176.200 49.200 ;
        RECT 180.600 47.200 180.900 53.800 ;
        RECT 183.800 52.100 184.200 57.900 ;
        RECT 187.000 54.800 187.400 55.200 ;
        RECT 187.000 54.200 187.300 54.800 ;
        RECT 188.600 54.200 188.900 58.800 ;
        RECT 203.000 56.200 203.300 66.800 ;
        RECT 205.400 65.800 205.800 66.200 ;
        RECT 206.200 65.800 206.600 66.200 ;
        RECT 204.600 58.800 205.000 59.200 ;
        RECT 189.400 55.800 189.800 56.200 ;
        RECT 203.000 55.800 203.400 56.200 ;
        RECT 204.600 56.100 204.900 58.800 ;
        RECT 205.400 57.200 205.700 65.800 ;
        RECT 206.200 59.200 206.500 65.800 ;
        RECT 206.200 58.800 206.600 59.200 ;
        RECT 207.800 58.200 208.100 74.800 ;
        RECT 208.600 72.200 208.900 74.800 ;
        RECT 208.600 71.800 209.000 72.200 ;
        RECT 209.400 71.800 209.800 72.200 ;
        RECT 209.400 70.200 209.700 71.800 ;
        RECT 209.400 69.800 209.800 70.200 ;
        RECT 209.400 67.800 209.800 68.200 ;
        RECT 209.400 66.200 209.700 67.800 ;
        RECT 209.400 65.800 209.800 66.200 ;
        RECT 207.800 57.800 208.200 58.200 ;
        RECT 205.400 56.800 205.800 57.200 ;
        RECT 204.600 55.800 205.700 56.100 ;
        RECT 189.400 55.200 189.700 55.800 ;
        RECT 203.000 55.200 203.300 55.800 ;
        RECT 189.400 54.800 189.800 55.200 ;
        RECT 191.800 54.800 192.200 55.200 ;
        RECT 195.800 54.800 196.200 55.200 ;
        RECT 196.600 54.800 197.000 55.200 ;
        RECT 198.200 55.100 198.600 55.200 ;
        RECT 199.000 55.100 199.400 55.200 ;
        RECT 198.200 54.800 199.400 55.100 ;
        RECT 201.400 54.800 201.800 55.200 ;
        RECT 203.000 54.800 203.400 55.200 ;
        RECT 187.000 53.800 187.400 54.200 ;
        RECT 187.800 53.800 188.200 54.200 ;
        RECT 188.600 53.800 189.000 54.200 ;
        RECT 190.200 54.100 190.600 54.200 ;
        RECT 191.000 54.100 191.400 54.200 ;
        RECT 190.200 53.800 191.400 54.100 ;
        RECT 187.000 53.100 187.400 53.200 ;
        RECT 187.800 53.100 188.100 53.800 ;
        RECT 191.800 53.200 192.100 54.800 ;
        RECT 195.800 54.200 196.100 54.800 ;
        RECT 192.600 53.800 193.000 54.200 ;
        RECT 195.800 53.800 196.200 54.200 ;
        RECT 187.000 52.800 188.100 53.100 ;
        RECT 190.200 52.800 190.600 53.200 ;
        RECT 191.800 52.800 192.200 53.200 ;
        RECT 186.200 52.100 186.600 52.200 ;
        RECT 187.000 52.100 187.400 52.200 ;
        RECT 186.200 51.800 187.400 52.100 ;
        RECT 190.200 49.200 190.500 52.800 ;
        RECT 191.800 52.200 192.100 52.800 ;
        RECT 191.800 51.800 192.200 52.200 ;
        RECT 192.600 49.200 192.900 53.800 ;
        RECT 196.600 52.200 196.900 54.800 ;
        RECT 201.400 54.200 201.700 54.800 ;
        RECT 197.400 53.800 197.800 54.200 ;
        RECT 201.400 53.800 201.800 54.200 ;
        RECT 197.400 53.200 197.700 53.800 ;
        RECT 197.400 52.800 197.800 53.200 ;
        RECT 196.600 51.800 197.000 52.200 ;
        RECT 200.600 51.800 201.000 52.200 ;
        RECT 196.600 51.200 196.900 51.800 ;
        RECT 196.600 50.800 197.000 51.200 ;
        RECT 190.200 48.800 190.600 49.200 ;
        RECT 192.600 48.800 193.000 49.200 ;
        RECT 180.600 47.100 181.000 47.200 ;
        RECT 181.400 47.100 181.800 47.200 ;
        RECT 180.600 46.800 181.800 47.100 ;
        RECT 187.000 46.100 187.400 46.200 ;
        RECT 187.800 46.100 188.200 46.200 ;
        RECT 187.000 45.800 188.200 46.100 ;
        RECT 188.600 45.800 189.000 46.200 ;
        RECT 191.000 45.800 191.400 46.200 ;
        RECT 188.600 45.200 188.900 45.800 ;
        RECT 179.800 44.800 180.200 45.200 ;
        RECT 188.600 44.800 189.000 45.200 ;
        RECT 178.200 42.800 178.600 43.200 ;
        RECT 178.200 42.200 178.500 42.800 ;
        RECT 172.600 41.800 173.000 42.200 ;
        RECT 178.200 41.800 178.600 42.200 ;
        RECT 171.000 38.800 171.400 39.200 ;
        RECT 167.000 34.800 167.400 35.200 ;
        RECT 168.600 34.800 169.000 35.200 ;
        RECT 169.400 34.800 169.800 35.200 ;
        RECT 170.200 34.800 170.600 35.200 ;
        RECT 167.000 34.200 167.300 34.800 ;
        RECT 168.600 34.200 168.900 34.800 ;
        RECT 167.000 33.800 167.400 34.200 ;
        RECT 168.600 33.800 169.000 34.200 ;
        RECT 167.000 32.200 167.300 33.800 ;
        RECT 169.400 33.200 169.700 34.800 ;
        RECT 170.200 34.200 170.500 34.800 ;
        RECT 170.200 33.800 170.600 34.200 ;
        RECT 171.800 33.800 172.200 34.200 ;
        RECT 169.400 32.800 169.800 33.200 ;
        RECT 167.000 31.800 167.400 32.200 ;
        RECT 167.800 31.800 168.200 32.200 ;
        RECT 171.000 31.800 171.400 32.200 ;
        RECT 167.000 29.800 167.400 30.200 ;
        RECT 167.000 29.200 167.300 29.800 ;
        RECT 167.000 28.800 167.400 29.200 ;
        RECT 167.000 28.200 167.300 28.800 ;
        RECT 167.000 27.800 167.400 28.200 ;
        RECT 167.800 26.200 168.100 31.800 ;
        RECT 169.400 27.800 169.800 28.200 ;
        RECT 169.400 27.200 169.700 27.800 ;
        RECT 171.000 27.200 171.300 31.800 ;
        RECT 171.800 29.200 172.100 33.800 ;
        RECT 171.800 28.800 172.200 29.200 ;
        RECT 169.400 26.800 169.800 27.200 ;
        RECT 171.000 26.800 171.400 27.200 ;
        RECT 159.000 25.800 159.400 26.200 ;
        RECT 161.400 25.800 161.800 26.200 ;
        RECT 163.000 26.100 163.400 26.200 ;
        RECT 163.800 26.100 164.200 26.200 ;
        RECT 163.000 25.800 164.200 26.100 ;
        RECT 166.200 25.800 166.600 26.200 ;
        RECT 167.800 25.800 168.200 26.200 ;
        RECT 169.400 26.100 169.800 26.200 ;
        RECT 170.200 26.100 170.600 26.200 ;
        RECT 169.400 25.800 170.600 26.100 ;
        RECT 161.400 25.200 161.700 25.800 ;
        RECT 161.400 24.800 161.800 25.200 ;
        RECT 165.400 23.800 165.800 24.200 ;
        RECT 158.200 21.800 158.600 22.200 ;
        RECT 158.200 17.200 158.500 21.800 ;
        RECT 159.000 18.100 159.400 18.200 ;
        RECT 159.800 18.100 160.200 18.200 ;
        RECT 159.000 17.800 160.200 18.100 ;
        RECT 158.200 16.800 158.600 17.200 ;
        RECT 159.800 16.800 160.200 17.200 ;
        RECT 158.200 15.100 158.600 15.200 ;
        RECT 159.000 15.100 159.400 15.200 ;
        RECT 158.200 14.800 159.400 15.100 ;
        RECT 159.800 14.200 160.100 16.800 ;
        RECT 159.800 13.800 160.200 14.200 ;
        RECT 159.800 8.200 160.100 13.800 ;
        RECT 160.600 13.100 161.000 15.900 ;
        RECT 161.400 13.800 161.800 14.200 ;
        RECT 159.800 7.800 160.200 8.200 ;
        RECT 161.400 7.200 161.700 13.800 ;
        RECT 162.200 12.100 162.600 17.900 ;
        RECT 163.000 17.800 163.400 18.200 ;
        RECT 163.000 15.100 163.300 17.800 ;
        RECT 164.600 16.800 165.000 17.200 ;
        RECT 163.000 14.700 163.400 15.100 ;
        RECT 163.800 10.800 164.200 11.200 ;
        RECT 163.800 7.200 164.100 10.800 ;
        RECT 164.600 7.200 164.900 16.800 ;
        RECT 157.400 6.800 157.800 7.200 ;
        RECT 161.400 6.800 161.800 7.200 ;
        RECT 163.800 6.800 164.200 7.200 ;
        RECT 164.600 6.800 165.000 7.200 ;
        RECT 157.400 6.200 157.700 6.800 ;
        RECT 165.400 6.200 165.700 23.800 ;
        RECT 170.200 20.800 170.600 21.200 ;
        RECT 167.000 12.100 167.400 17.900 ;
        RECT 169.400 16.800 169.800 17.200 ;
        RECT 169.400 14.200 169.700 16.800 ;
        RECT 170.200 16.200 170.500 20.800 ;
        RECT 170.200 15.800 170.600 16.200 ;
        RECT 171.000 14.200 171.300 26.800 ;
        RECT 172.600 23.200 172.900 41.800 ;
        RECT 179.800 39.200 180.100 44.800 ;
        RECT 186.200 41.800 186.600 42.200 ;
        RECT 186.200 39.200 186.500 41.800 ;
        RECT 179.800 38.800 180.200 39.200 ;
        RECT 186.200 38.800 186.600 39.200 ;
        RECT 182.200 36.800 182.600 37.200 ;
        RECT 187.000 37.100 187.400 37.200 ;
        RECT 187.800 37.100 188.200 37.200 ;
        RECT 187.000 36.800 188.200 37.100 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 176.600 35.100 177.000 35.200 ;
        RECT 177.400 35.100 177.800 35.200 ;
        RECT 176.600 34.800 177.800 35.100 ;
        RECT 178.200 34.800 178.600 35.200 ;
        RECT 172.600 22.800 173.000 23.200 ;
        RECT 171.800 18.800 172.200 19.200 ;
        RECT 171.800 14.200 172.100 18.800 ;
        RECT 172.600 18.200 172.900 22.800 ;
        RECT 173.400 19.200 173.700 34.800 ;
        RECT 177.400 34.200 177.700 34.800 ;
        RECT 177.400 33.800 177.800 34.200 ;
        RECT 175.800 31.800 176.200 32.200 ;
        RECT 175.800 31.200 176.100 31.800 ;
        RECT 175.800 30.800 176.200 31.200 ;
        RECT 178.200 29.200 178.500 34.800 ;
        RECT 182.200 34.200 182.500 36.800 ;
        RECT 183.800 35.800 184.200 36.200 ;
        RECT 186.200 36.100 186.600 36.200 ;
        RECT 187.000 36.100 187.400 36.200 ;
        RECT 186.200 35.800 187.400 36.100 ;
        RECT 183.800 35.200 184.100 35.800 ;
        RECT 183.800 34.800 184.200 35.200 ;
        RECT 185.400 35.100 185.800 35.200 ;
        RECT 186.200 35.100 186.600 35.200 ;
        RECT 185.400 34.800 186.600 35.100 ;
        RECT 182.200 33.800 182.600 34.200 ;
        RECT 174.200 23.100 174.600 28.900 ;
        RECT 178.200 28.800 178.600 29.200 ;
        RECT 177.400 27.800 177.800 28.200 ;
        RECT 176.600 26.800 177.000 27.200 ;
        RECT 174.200 20.800 174.600 21.200 ;
        RECT 173.400 18.800 173.800 19.200 ;
        RECT 172.600 17.800 173.000 18.200 ;
        RECT 174.200 15.200 174.500 20.800 ;
        RECT 175.000 19.100 175.400 19.200 ;
        RECT 175.800 19.100 176.200 19.200 ;
        RECT 175.000 18.800 176.200 19.100 ;
        RECT 172.600 15.100 173.000 15.200 ;
        RECT 173.400 15.100 173.800 15.200 ;
        RECT 172.600 14.800 173.800 15.100 ;
        RECT 174.200 14.800 174.600 15.200 ;
        RECT 169.400 13.800 169.800 14.200 ;
        RECT 171.000 13.800 171.400 14.200 ;
        RECT 171.800 13.800 172.200 14.200 ;
        RECT 174.200 14.100 174.600 14.200 ;
        RECT 175.000 14.100 175.400 14.200 ;
        RECT 174.200 13.800 175.400 14.100 ;
        RECT 167.800 8.800 168.200 9.200 ;
        RECT 169.400 9.100 169.800 9.200 ;
        RECT 170.200 9.100 170.600 9.200 ;
        RECT 169.400 8.800 170.600 9.100 ;
        RECT 167.800 7.200 168.100 8.800 ;
        RECT 167.000 6.800 167.400 7.200 ;
        RECT 167.800 6.800 168.200 7.200 ;
        RECT 167.000 6.200 167.300 6.800 ;
        RECT 157.400 5.800 157.800 6.200 ;
        RECT 165.400 5.800 165.800 6.200 ;
        RECT 167.000 5.800 167.400 6.200 ;
        RECT 169.400 5.800 169.800 6.200 ;
        RECT 169.400 5.200 169.700 5.800 ;
        RECT 169.400 4.800 169.800 5.200 ;
        RECT 172.600 3.100 173.000 8.900 ;
        RECT 176.600 8.200 176.900 26.800 ;
        RECT 177.400 26.200 177.700 27.800 ;
        RECT 177.400 25.800 177.800 26.200 ;
        RECT 179.000 23.100 179.400 28.900 ;
        RECT 181.400 28.800 181.800 29.200 ;
        RECT 180.600 25.100 181.000 27.900 ;
        RECT 181.400 27.200 181.700 28.800 ;
        RECT 181.400 26.800 181.800 27.200 ;
        RECT 183.000 25.800 183.400 26.200 ;
        RECT 183.000 25.200 183.300 25.800 ;
        RECT 182.200 25.100 182.600 25.200 ;
        RECT 183.000 25.100 183.400 25.200 ;
        RECT 182.200 24.800 183.400 25.100 ;
        RECT 183.800 22.200 184.100 34.800 ;
        RECT 187.000 34.100 187.400 34.200 ;
        RECT 186.200 33.800 187.400 34.100 ;
        RECT 186.200 32.200 186.500 33.800 ;
        RECT 186.200 31.800 186.600 32.200 ;
        RECT 190.200 32.100 190.600 37.900 ;
        RECT 186.200 28.200 186.500 31.800 ;
        RECT 187.000 29.100 187.400 29.200 ;
        RECT 187.800 29.100 188.200 29.200 ;
        RECT 187.000 28.800 188.200 29.100 ;
        RECT 186.200 27.800 186.600 28.200 ;
        RECT 186.200 27.200 186.500 27.800 ;
        RECT 186.200 26.800 186.600 27.200 ;
        RECT 184.600 26.100 185.000 26.200 ;
        RECT 185.400 26.100 185.800 26.200 ;
        RECT 184.600 25.800 185.800 26.100 ;
        RECT 185.400 25.100 185.800 25.200 ;
        RECT 186.200 25.100 186.600 25.200 ;
        RECT 185.400 24.800 186.600 25.100 ;
        RECT 189.400 23.100 189.800 28.900 ;
        RECT 190.200 25.800 190.600 26.200 ;
        RECT 183.800 21.800 184.200 22.200 ;
        RECT 190.200 22.100 190.500 25.800 ;
        RECT 191.000 23.200 191.300 45.800 ;
        RECT 195.000 43.100 195.400 48.900 ;
        RECT 195.800 46.800 196.200 47.200 ;
        RECT 199.000 46.800 199.400 47.200 ;
        RECT 195.800 46.200 196.100 46.800 ;
        RECT 199.000 46.300 199.300 46.800 ;
        RECT 195.800 45.800 196.200 46.200 ;
        RECT 199.000 45.900 199.400 46.300 ;
        RECT 191.800 38.800 192.200 39.200 ;
        RECT 191.800 35.200 192.100 38.800 ;
        RECT 193.400 35.800 193.800 36.200 ;
        RECT 193.400 35.200 193.700 35.800 ;
        RECT 191.800 34.800 192.200 35.200 ;
        RECT 193.400 34.800 193.800 35.200 ;
        RECT 191.000 22.800 191.400 23.200 ;
        RECT 189.400 21.800 190.500 22.100 ;
        RECT 178.200 12.100 178.600 17.900 ;
        RECT 179.800 15.100 180.200 15.200 ;
        RECT 180.600 15.100 181.000 15.200 ;
        RECT 179.800 14.800 181.000 15.100 ;
        RECT 183.000 12.100 183.400 17.900 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 183.800 14.200 184.100 14.800 ;
        RECT 183.800 13.800 184.200 14.200 ;
        RECT 184.600 13.100 185.000 15.900 ;
        RECT 186.200 15.800 186.600 16.200 ;
        RECT 187.800 16.100 188.200 16.200 ;
        RECT 188.600 16.100 189.000 16.200 ;
        RECT 187.800 15.800 189.000 16.100 ;
        RECT 186.200 15.200 186.500 15.800 ;
        RECT 186.200 14.800 186.600 15.200 ;
        RECT 185.400 14.100 185.800 14.200 ;
        RECT 186.200 14.100 186.600 14.200 ;
        RECT 185.400 13.800 186.600 14.100 ;
        RECT 176.600 7.800 177.000 8.200 ;
        RECT 175.800 6.800 176.200 7.200 ;
        RECT 175.800 6.200 176.100 6.800 ;
        RECT 175.800 5.800 176.200 6.200 ;
        RECT 177.400 3.100 177.800 8.900 ;
        RECT 181.400 8.800 181.800 9.200 ;
        RECT 185.400 9.100 185.700 13.800 ;
        RECT 187.800 12.800 188.200 13.200 ;
        RECT 187.800 12.200 188.100 12.800 ;
        RECT 187.800 11.800 188.200 12.200 ;
        RECT 184.600 8.800 185.700 9.100 ;
        RECT 178.200 7.800 178.600 8.200 ;
        RECT 178.200 7.200 178.500 7.800 ;
        RECT 178.200 6.800 178.600 7.200 ;
        RECT 179.000 5.100 179.400 7.900 ;
        RECT 181.400 7.200 181.700 8.800 ;
        RECT 184.600 7.200 184.900 8.800 ;
        RECT 180.600 6.800 181.000 7.200 ;
        RECT 181.400 6.800 181.800 7.200 ;
        RECT 183.800 6.800 184.200 7.200 ;
        RECT 184.600 6.800 185.000 7.200 ;
        RECT 180.600 5.200 180.900 6.800 ;
        RECT 183.800 6.200 184.100 6.800 ;
        RECT 183.800 5.800 184.200 6.200 ;
        RECT 179.800 5.100 180.200 5.200 ;
        RECT 180.600 5.100 181.000 5.200 ;
        RECT 179.800 4.800 181.000 5.100 ;
        RECT 183.800 4.800 184.200 5.200 ;
        RECT 185.400 5.100 185.800 7.900 ;
        RECT 183.800 4.200 184.100 4.800 ;
        RECT 183.800 3.800 184.200 4.200 ;
        RECT 187.000 3.100 187.400 8.900 ;
        RECT 189.400 8.200 189.700 21.800 ;
        RECT 190.200 16.800 190.600 17.200 ;
        RECT 190.200 14.200 190.500 16.800 ;
        RECT 190.200 13.800 190.600 14.200 ;
        RECT 191.000 13.100 191.400 15.900 ;
        RECT 191.800 15.200 192.100 34.800 ;
        RECT 195.000 32.100 195.400 37.900 ;
        RECT 195.800 31.100 196.100 45.800 ;
        RECT 199.000 44.800 199.400 45.200 ;
        RECT 199.000 39.200 199.300 44.800 ;
        RECT 199.800 43.100 200.200 48.900 ;
        RECT 200.600 46.200 200.900 51.800 ;
        RECT 204.600 50.800 205.000 51.200 ;
        RECT 200.600 45.800 201.000 46.200 ;
        RECT 201.400 45.100 201.800 47.900 ;
        RECT 203.000 46.800 203.400 47.200 ;
        RECT 203.000 46.200 203.300 46.800 ;
        RECT 204.600 46.200 204.900 50.800 ;
        RECT 205.400 49.200 205.700 55.800 ;
        RECT 207.800 53.800 208.200 54.200 ;
        RECT 205.400 48.800 205.800 49.200 ;
        RECT 207.000 48.800 207.400 49.200 ;
        RECT 207.000 46.200 207.300 48.800 ;
        RECT 207.800 47.200 208.100 53.800 ;
        RECT 208.600 49.100 209.000 49.200 ;
        RECT 209.400 49.100 209.800 49.200 ;
        RECT 208.600 48.800 209.800 49.100 ;
        RECT 207.800 46.800 208.200 47.200 ;
        RECT 203.000 45.800 203.400 46.200 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 207.000 45.800 207.400 46.200 ;
        RECT 207.800 45.800 208.200 46.200 ;
        RECT 207.800 44.200 208.100 45.800 ;
        RECT 207.800 43.800 208.200 44.200 ;
        RECT 199.000 38.800 199.400 39.200 ;
        RECT 207.000 38.800 207.400 39.200 ;
        RECT 197.400 37.800 197.800 38.200 ;
        RECT 196.600 33.100 197.000 35.900 ;
        RECT 197.400 35.200 197.700 37.800 ;
        RECT 197.400 34.800 197.800 35.200 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 200.600 34.800 201.000 35.200 ;
        RECT 195.000 30.800 196.100 31.100 ;
        RECT 196.600 30.800 197.000 31.200 ;
        RECT 192.600 25.800 193.000 26.200 ;
        RECT 193.400 25.800 193.800 26.200 ;
        RECT 192.600 25.200 192.900 25.800 ;
        RECT 192.600 24.800 193.000 25.200 ;
        RECT 191.800 14.800 192.200 15.200 ;
        RECT 191.800 14.200 192.100 14.800 ;
        RECT 191.800 13.800 192.200 14.200 ;
        RECT 192.600 12.100 193.000 17.900 ;
        RECT 193.400 9.200 193.700 25.800 ;
        RECT 194.200 23.100 194.600 28.900 ;
        RECT 195.000 27.200 195.300 30.800 ;
        RECT 195.000 26.800 195.400 27.200 ;
        RECT 195.800 25.100 196.200 27.900 ;
        RECT 196.600 26.200 196.900 30.800 ;
        RECT 198.200 29.200 198.500 34.800 ;
        RECT 198.200 28.800 198.600 29.200 ;
        RECT 200.600 29.100 200.900 34.800 ;
        RECT 204.600 32.800 205.000 33.200 ;
        RECT 202.200 32.100 202.600 32.200 ;
        RECT 203.000 32.100 203.400 32.200 ;
        RECT 202.200 31.800 203.400 32.100 ;
        RECT 204.600 29.200 204.900 32.800 ;
        RECT 205.400 31.800 205.800 32.200 ;
        RECT 206.200 32.100 206.600 37.900 ;
        RECT 207.000 35.200 207.300 38.800 ;
        RECT 207.000 34.800 207.400 35.200 ;
        RECT 208.600 34.800 209.000 35.200 ;
        RECT 200.600 28.800 201.700 29.100 ;
        RECT 204.600 28.800 205.000 29.200 ;
        RECT 196.600 25.800 197.000 26.200 ;
        RECT 197.400 25.800 197.800 26.200 ;
        RECT 199.800 26.100 200.200 26.200 ;
        RECT 200.600 26.100 201.000 26.200 ;
        RECT 199.800 25.800 201.000 26.100 ;
        RECT 197.400 25.200 197.700 25.800 ;
        RECT 197.400 24.800 197.800 25.200 ;
        RECT 194.200 14.800 194.600 15.200 ;
        RECT 194.200 13.200 194.500 14.800 ;
        RECT 195.000 13.800 195.400 14.200 ;
        RECT 194.200 12.800 194.600 13.200 ;
        RECT 193.400 9.100 193.800 9.200 ;
        RECT 194.200 9.100 194.600 9.200 ;
        RECT 189.400 7.800 189.800 8.200 ;
        RECT 189.400 7.200 189.700 7.800 ;
        RECT 189.400 6.800 189.800 7.200 ;
        RECT 187.800 5.900 188.200 6.300 ;
        RECT 187.800 5.200 188.100 5.900 ;
        RECT 187.800 4.800 188.200 5.200 ;
        RECT 191.800 3.100 192.200 8.900 ;
        RECT 193.400 8.800 194.600 9.100 ;
        RECT 195.000 7.200 195.300 13.800 ;
        RECT 197.400 12.100 197.800 17.900 ;
        RECT 199.000 17.100 199.400 17.200 ;
        RECT 199.800 17.100 200.200 17.200 ;
        RECT 199.000 16.800 200.200 17.100 ;
        RECT 201.400 14.200 201.700 28.800 ;
        RECT 205.400 27.200 205.700 31.800 ;
        RECT 208.600 29.200 208.900 34.800 ;
        RECT 208.600 28.800 209.000 29.200 ;
        RECT 210.200 27.200 210.500 83.800 ;
        RECT 211.800 83.100 212.200 88.900 ;
        RECT 212.600 87.800 213.000 88.200 ;
        RECT 212.600 87.200 212.900 87.800 ;
        RECT 212.600 86.800 213.000 87.200 ;
        RECT 213.400 85.100 213.800 87.900 ;
        RECT 214.200 86.800 214.600 87.200 ;
        RECT 216.600 87.100 216.900 91.800 ;
        RECT 220.600 89.200 220.900 95.800 ;
        RECT 220.600 88.800 221.000 89.200 ;
        RECT 217.400 87.100 217.800 87.200 ;
        RECT 216.600 86.800 217.800 87.100 ;
        RECT 219.000 87.100 219.400 87.200 ;
        RECT 219.800 87.100 220.200 87.200 ;
        RECT 219.000 86.800 220.200 87.100 ;
        RECT 214.200 86.200 214.500 86.800 ;
        RECT 217.400 86.200 217.700 86.800 ;
        RECT 221.400 86.200 221.700 100.800 ;
        RECT 222.200 95.200 222.500 104.800 ;
        RECT 224.600 104.200 224.900 105.800 ;
        RECT 224.600 103.800 225.000 104.200 ;
        RECT 226.200 103.200 226.500 114.800 ;
        RECT 228.600 114.200 228.900 114.800 ;
        RECT 228.600 113.800 229.000 114.200 ;
        RECT 227.000 111.800 227.400 112.200 ;
        RECT 227.000 109.200 227.300 111.800 ;
        RECT 227.000 108.800 227.400 109.200 ;
        RECT 228.600 108.800 229.000 109.200 ;
        RECT 227.800 106.800 228.200 107.200 ;
        RECT 227.800 106.200 228.100 106.800 ;
        RECT 227.800 105.800 228.200 106.200 ;
        RECT 227.000 104.800 227.400 105.200 ;
        RECT 227.000 104.200 227.300 104.800 ;
        RECT 227.000 103.800 227.400 104.200 ;
        RECT 226.200 102.800 226.600 103.200 ;
        RECT 222.200 94.800 222.600 95.200 ;
        RECT 223.000 94.700 223.400 95.100 ;
        RECT 223.000 94.200 223.300 94.700 ;
        RECT 223.000 93.800 223.400 94.200 ;
        RECT 222.200 91.800 222.600 92.200 ;
        RECT 223.800 92.100 224.200 97.900 ;
        RECT 226.200 96.100 226.600 96.200 ;
        RECT 227.000 96.100 227.400 96.200 ;
        RECT 225.400 93.100 225.800 95.900 ;
        RECT 226.200 95.800 227.400 96.100 ;
        RECT 228.600 95.200 228.900 108.800 ;
        RECT 229.400 105.800 229.800 106.200 ;
        RECT 229.400 105.200 229.700 105.800 ;
        RECT 229.400 104.800 229.800 105.200 ;
        RECT 230.200 101.200 230.500 114.800 ;
        RECT 231.800 113.800 232.200 114.200 ;
        RECT 231.800 113.200 232.100 113.800 ;
        RECT 231.800 112.800 232.200 113.200 ;
        RECT 231.800 106.800 232.200 107.200 ;
        RECT 231.800 106.200 232.100 106.800 ;
        RECT 231.800 105.800 232.200 106.200 ;
        RECT 230.200 100.800 230.600 101.200 ;
        RECT 232.600 96.200 232.900 114.800 ;
        RECT 238.200 114.200 238.500 115.800 ;
        RECT 237.400 113.800 237.800 114.200 ;
        RECT 238.200 113.800 238.600 114.200 ;
        RECT 237.400 113.200 237.700 113.800 ;
        RECT 237.400 112.800 237.800 113.200 ;
        RECT 240.600 113.100 241.000 115.900 ;
        RECT 241.400 115.200 241.700 121.800 ;
        RECT 242.200 120.200 242.500 134.800 ;
        RECT 243.000 123.200 243.300 141.800 ;
        RECT 243.800 139.200 244.100 146.800 ;
        RECT 244.600 146.200 244.900 146.800 ;
        RECT 244.600 145.800 245.000 146.200 ;
        RECT 243.800 138.800 244.200 139.200 ;
        RECT 243.800 131.800 244.200 132.200 ;
        RECT 243.800 131.200 244.100 131.800 ;
        RECT 243.800 130.800 244.200 131.200 ;
        RECT 243.000 122.800 243.400 123.200 ;
        RECT 243.800 123.100 244.200 128.900 ;
        RECT 245.400 127.200 245.700 153.800 ;
        RECT 246.200 153.100 246.600 155.900 ;
        RECT 247.800 155.100 248.200 155.200 ;
        RECT 248.600 155.100 249.000 155.200 ;
        RECT 247.800 154.800 249.000 155.100 ;
        RECT 248.600 153.800 249.000 154.200 ;
        RECT 247.000 152.800 247.400 153.200 ;
        RECT 247.000 129.200 247.300 152.800 ;
        RECT 247.800 151.800 248.200 152.200 ;
        RECT 247.800 150.200 248.100 151.800 ;
        RECT 247.800 149.800 248.200 150.200 ;
        RECT 247.800 143.100 248.200 148.900 ;
        RECT 248.600 132.200 248.900 153.800 ;
        RECT 250.200 151.800 250.600 152.200 ;
        RECT 250.200 151.200 250.500 151.800 ;
        RECT 250.200 150.800 250.600 151.200 ;
        RECT 250.200 148.800 250.600 149.200 ;
        RECT 250.200 148.200 250.500 148.800 ;
        RECT 250.200 147.800 250.600 148.200 ;
        RECT 249.400 133.800 249.800 134.200 ;
        RECT 248.600 131.800 249.000 132.200 ;
        RECT 247.000 128.800 247.400 129.200 ;
        RECT 245.400 126.800 245.800 127.200 ;
        RECT 244.600 126.100 245.000 126.200 ;
        RECT 245.400 126.100 245.800 126.200 ;
        RECT 244.600 125.800 245.800 126.100 ;
        RECT 245.400 122.800 245.800 123.200 ;
        RECT 248.600 123.100 249.000 128.900 ;
        RECT 249.400 127.200 249.700 133.800 ;
        RECT 249.400 126.800 249.800 127.200 ;
        RECT 250.200 125.100 250.600 127.900 ;
        RECT 242.200 119.800 242.600 120.200 ;
        RECT 241.400 114.800 241.800 115.200 ;
        RECT 241.400 113.800 241.800 114.200 ;
        RECT 241.400 113.200 241.700 113.800 ;
        RECT 241.400 112.800 241.800 113.200 ;
        RECT 236.600 111.800 237.000 112.200 ;
        RECT 236.600 109.200 236.900 111.800 ;
        RECT 237.400 109.200 237.700 112.800 ;
        RECT 242.200 112.100 242.600 117.900 ;
        RECT 243.000 115.800 243.400 116.200 ;
        RECT 243.000 115.100 243.300 115.800 ;
        RECT 243.000 114.700 243.400 115.100 ;
        RECT 241.400 110.800 241.800 111.200 ;
        RECT 241.400 109.200 241.700 110.800 ;
        RECT 236.600 108.800 237.000 109.200 ;
        RECT 237.400 108.800 237.800 109.200 ;
        RECT 241.400 108.800 241.800 109.200 ;
        RECT 243.800 108.800 244.200 109.200 ;
        RECT 243.800 107.200 244.100 108.800 ;
        RECT 239.000 106.800 239.400 107.200 ;
        RECT 243.800 106.800 244.200 107.200 ;
        RECT 239.000 106.200 239.300 106.800 ;
        RECT 235.800 105.800 236.200 106.200 ;
        RECT 239.000 105.800 239.400 106.200 ;
        RECT 240.600 105.800 241.000 106.200 ;
        RECT 243.000 106.100 243.400 106.200 ;
        RECT 243.800 106.100 244.200 106.200 ;
        RECT 243.000 105.800 244.200 106.100 ;
        RECT 244.600 105.800 245.000 106.200 ;
        RECT 231.800 95.800 232.200 96.200 ;
        RECT 232.600 95.800 233.000 96.200 ;
        RECT 226.200 94.800 226.600 95.200 ;
        RECT 228.600 94.800 229.000 95.200 ;
        RECT 230.200 95.100 230.600 95.200 ;
        RECT 231.000 95.100 231.400 95.200 ;
        RECT 230.200 94.800 231.400 95.100 ;
        RECT 226.200 94.200 226.500 94.800 ;
        RECT 226.200 93.800 226.600 94.200 ;
        RECT 222.200 86.200 222.500 91.800 ;
        RECT 226.200 88.800 226.600 89.200 ;
        RECT 226.200 87.200 226.500 88.800 ;
        RECT 226.200 86.800 226.600 87.200 ;
        RECT 214.200 85.800 214.600 86.200 ;
        RECT 215.000 85.800 215.400 86.200 ;
        RECT 217.400 85.800 217.800 86.200 ;
        RECT 218.200 86.100 218.600 86.200 ;
        RECT 219.000 86.100 219.400 86.200 ;
        RECT 218.200 85.800 219.400 86.100 ;
        RECT 221.400 85.800 221.800 86.200 ;
        RECT 222.200 85.800 222.600 86.200 ;
        RECT 227.800 85.800 228.200 86.200 ;
        RECT 214.200 80.800 214.600 81.200 ;
        RECT 212.600 79.800 213.000 80.200 ;
        RECT 211.000 77.800 211.400 78.200 ;
        RECT 211.000 72.200 211.300 77.800 ;
        RECT 211.800 74.800 212.200 75.200 ;
        RECT 211.800 74.200 212.100 74.800 ;
        RECT 212.600 74.200 212.900 79.800 ;
        RECT 214.200 76.200 214.500 80.800 ;
        RECT 215.000 78.200 215.300 85.800 ;
        RECT 219.800 85.100 220.200 85.200 ;
        RECT 220.600 85.100 221.000 85.200 ;
        RECT 219.800 84.800 221.000 85.100 ;
        RECT 219.800 82.200 220.100 84.800 ;
        RECT 219.800 81.800 220.200 82.200 ;
        RECT 215.000 77.800 215.400 78.200 ;
        RECT 216.600 76.800 217.000 77.200 ;
        RECT 216.600 76.200 216.900 76.800 ;
        RECT 214.200 75.800 214.600 76.200 ;
        RECT 215.000 76.100 215.400 76.200 ;
        RECT 215.800 76.100 216.200 76.200 ;
        RECT 215.000 75.800 216.200 76.100 ;
        RECT 216.600 75.800 217.000 76.200 ;
        RECT 219.000 76.100 219.400 76.200 ;
        RECT 219.800 76.100 220.200 76.200 ;
        RECT 219.000 75.800 220.200 76.100 ;
        RECT 211.800 73.800 212.200 74.200 ;
        RECT 212.600 73.800 213.000 74.200 ;
        RECT 211.000 71.800 211.400 72.200 ;
        RECT 211.000 69.200 211.300 71.800 ;
        RECT 212.600 70.200 212.900 73.800 ;
        RECT 213.400 71.800 213.800 72.200 ;
        RECT 212.600 69.800 213.000 70.200 ;
        RECT 211.000 68.800 211.400 69.200 ;
        RECT 213.400 67.200 213.700 71.800 ;
        RECT 211.800 67.100 212.200 67.200 ;
        RECT 212.600 67.100 213.000 67.200 ;
        RECT 211.800 66.800 213.000 67.100 ;
        RECT 213.400 66.800 213.800 67.200 ;
        RECT 213.400 65.800 213.800 66.200 ;
        RECT 213.400 63.200 213.700 65.800 ;
        RECT 213.400 63.100 213.800 63.200 ;
        RECT 214.200 63.100 214.500 75.800 ;
        RECT 215.000 74.800 215.400 75.200 ;
        RECT 219.800 75.100 220.200 75.200 ;
        RECT 219.000 74.800 220.200 75.100 ;
        RECT 215.000 74.200 215.300 74.800 ;
        RECT 215.000 73.800 215.400 74.200 ;
        RECT 217.400 73.800 217.800 74.200 ;
        RECT 217.400 72.200 217.700 73.800 ;
        RECT 217.400 71.800 217.800 72.200 ;
        RECT 215.800 69.800 216.200 70.200 ;
        RECT 215.800 69.200 216.100 69.800 ;
        RECT 215.800 68.800 216.200 69.200 ;
        RECT 215.000 66.800 215.400 67.200 ;
        RECT 215.000 66.200 215.300 66.800 ;
        RECT 215.000 65.800 215.400 66.200 ;
        RECT 215.000 64.800 215.400 65.200 ;
        RECT 215.000 64.200 215.300 64.800 ;
        RECT 215.000 63.800 215.400 64.200 ;
        RECT 218.200 63.100 218.600 68.900 ;
        RECT 213.400 62.800 214.500 63.100 ;
        RECT 213.400 55.100 213.800 55.200 ;
        RECT 214.200 55.100 214.600 55.200 ;
        RECT 213.400 54.800 214.600 55.100 ;
        RECT 215.000 51.800 215.400 52.200 ;
        RECT 217.400 52.100 217.800 57.900 ;
        RECT 218.200 54.800 218.600 55.200 ;
        RECT 218.200 54.200 218.500 54.800 ;
        RECT 218.200 53.800 218.600 54.200 ;
        RECT 215.000 51.200 215.300 51.800 ;
        RECT 215.000 50.800 215.400 51.200 ;
        RECT 211.000 43.100 211.400 48.900 ;
        RECT 211.800 46.800 212.200 47.200 ;
        RECT 211.800 46.200 212.100 46.800 ;
        RECT 214.200 46.200 214.600 46.300 ;
        RECT 215.000 46.200 215.400 46.300 ;
        RECT 211.800 45.800 212.200 46.200 ;
        RECT 214.200 45.900 215.400 46.200 ;
        RECT 215.800 43.100 216.200 48.900 ;
        RECT 218.200 48.800 218.600 49.200 ;
        RECT 217.400 45.100 217.800 47.900 ;
        RECT 218.200 47.200 218.500 48.800 ;
        RECT 218.200 46.800 218.600 47.200 ;
        RECT 211.000 32.100 211.400 37.900 ;
        RECT 213.400 36.800 213.800 37.200 ;
        RECT 213.400 36.200 213.700 36.800 ;
        RECT 212.600 33.100 213.000 35.900 ;
        RECT 213.400 35.800 213.800 36.200 ;
        RECT 211.800 27.800 212.200 28.200 ;
        RECT 211.800 27.200 212.100 27.800 ;
        RECT 205.400 26.800 205.800 27.200 ;
        RECT 207.800 26.800 208.200 27.200 ;
        RECT 210.200 26.800 210.600 27.200 ;
        RECT 211.800 27.100 212.200 27.200 ;
        RECT 212.600 27.100 213.000 27.200 ;
        RECT 211.800 26.800 213.000 27.100 ;
        RECT 205.400 26.200 205.700 26.800 ;
        RECT 205.400 25.800 205.800 26.200 ;
        RECT 207.800 25.200 208.100 26.800 ;
        RECT 210.200 26.200 210.500 26.800 ;
        RECT 209.400 25.800 209.800 26.200 ;
        RECT 210.200 25.800 210.600 26.200 ;
        RECT 212.600 26.100 213.000 26.200 ;
        RECT 213.400 26.100 213.700 35.800 ;
        RECT 215.000 34.800 215.400 35.200 ;
        RECT 215.800 34.800 216.200 35.200 ;
        RECT 216.600 35.100 217.000 35.200 ;
        RECT 217.400 35.100 217.800 35.200 ;
        RECT 216.600 34.800 218.500 35.100 ;
        RECT 215.000 34.200 215.300 34.800 ;
        RECT 215.800 34.200 216.100 34.800 ;
        RECT 215.000 33.800 215.400 34.200 ;
        RECT 215.800 33.800 216.200 34.200 ;
        RECT 212.600 25.800 213.700 26.100 ;
        RECT 214.200 31.800 214.600 32.200 ;
        RECT 207.800 24.800 208.200 25.200 ;
        RECT 204.600 21.800 205.000 22.200 ;
        RECT 204.600 15.200 204.900 21.800 ;
        RECT 206.200 17.800 206.600 18.200 ;
        RECT 206.200 15.200 206.500 17.800 ;
        RECT 209.400 15.200 209.700 25.800 ;
        RECT 214.200 25.200 214.500 31.800 ;
        RECT 218.200 29.200 218.500 34.800 ;
        RECT 219.000 34.200 219.300 74.800 ;
        RECT 219.800 73.800 220.200 74.200 ;
        RECT 220.600 73.800 221.000 74.200 ;
        RECT 219.800 73.200 220.100 73.800 ;
        RECT 219.800 72.800 220.200 73.200 ;
        RECT 220.600 69.200 220.900 73.800 ;
        RECT 220.600 68.800 221.000 69.200 ;
        RECT 220.600 66.800 221.000 67.200 ;
        RECT 220.600 66.200 220.900 66.800 ;
        RECT 220.600 65.800 221.000 66.200 ;
        RECT 221.400 60.200 221.700 85.800 ;
        RECT 227.800 85.200 228.100 85.800 ;
        RECT 228.600 85.200 228.900 94.800 ;
        RECT 231.800 94.200 232.100 95.800 ;
        RECT 232.600 95.200 232.900 95.800 ;
        RECT 232.600 94.800 233.000 95.200 ;
        RECT 229.400 93.800 229.800 94.200 ;
        RECT 231.800 93.800 232.200 94.200 ;
        RECT 234.200 93.800 234.600 94.200 ;
        RECT 229.400 91.200 229.700 93.800 ;
        RECT 234.200 92.200 234.500 93.800 ;
        RECT 235.000 93.100 235.400 95.900 ;
        RECT 235.800 94.200 236.100 105.800 ;
        RECT 240.600 105.200 240.900 105.800 ;
        RECT 240.600 104.800 241.000 105.200 ;
        RECT 235.800 93.800 236.200 94.200 ;
        RECT 234.200 91.800 234.600 92.200 ;
        RECT 229.400 90.800 229.800 91.200 ;
        RECT 231.000 90.800 231.400 91.200 ;
        RECT 230.200 89.800 230.600 90.200 ;
        RECT 230.200 86.200 230.500 89.800 ;
        RECT 231.000 87.200 231.300 90.800 ;
        RECT 231.000 86.800 231.400 87.200 ;
        RECT 230.200 85.800 230.600 86.200 ;
        RECT 227.800 84.800 228.200 85.200 ;
        RECT 228.600 84.800 229.000 85.200 ;
        RECT 230.200 84.800 230.600 85.200 ;
        RECT 231.800 85.100 232.200 87.900 ;
        RECT 232.600 87.800 233.000 88.200 ;
        RECT 232.600 87.200 232.900 87.800 ;
        RECT 232.600 86.800 233.000 87.200 ;
        RECT 230.200 84.200 230.500 84.800 ;
        RECT 230.200 83.800 230.600 84.200 ;
        RECT 232.600 84.100 232.900 86.800 ;
        RECT 231.800 83.800 232.900 84.100 ;
        RECT 224.600 82.800 225.000 83.200 ;
        RECT 223.800 81.800 224.200 82.200 ;
        RECT 223.800 75.200 224.100 81.800 ;
        RECT 224.600 75.200 224.900 82.800 ;
        RECT 225.400 76.800 225.800 77.200 ;
        RECT 225.400 75.200 225.700 76.800 ;
        RECT 223.800 74.800 224.200 75.200 ;
        RECT 224.600 74.800 225.000 75.200 ;
        RECT 225.400 74.800 225.800 75.200 ;
        RECT 227.800 72.100 228.200 77.900 ;
        RECT 230.200 77.800 230.600 78.200 ;
        RECT 229.400 74.800 229.800 75.200 ;
        RECT 229.400 74.200 229.700 74.800 ;
        RECT 229.400 73.800 229.800 74.200 ;
        RECT 223.000 63.100 223.400 68.900 ;
        RECT 226.200 68.800 226.600 69.200 ;
        RECT 223.800 67.800 224.200 68.200 ;
        RECT 223.800 67.200 224.100 67.800 ;
        RECT 223.800 66.800 224.200 67.200 ;
        RECT 224.600 65.100 225.000 67.900 ;
        RECT 225.400 67.800 225.800 68.200 ;
        RECT 225.400 67.200 225.700 67.800 ;
        RECT 225.400 66.800 225.800 67.200 ;
        RECT 226.200 66.200 226.500 68.800 ;
        RECT 229.400 68.100 229.800 68.200 ;
        RECT 228.600 67.800 229.800 68.100 ;
        RECT 228.600 66.200 228.900 67.800 ;
        RECT 230.200 67.200 230.500 77.800 ;
        RECT 231.800 73.200 232.100 83.800 ;
        RECT 233.400 83.100 233.800 88.900 ;
        RECT 234.200 85.900 234.600 86.300 ;
        RECT 234.200 85.200 234.500 85.900 ;
        RECT 234.200 84.800 234.600 85.200 ;
        RECT 231.800 72.800 232.200 73.200 ;
        RECT 231.800 68.200 232.100 72.800 ;
        RECT 232.600 72.100 233.000 77.900 ;
        RECT 234.200 73.100 234.600 75.900 ;
        RECT 235.000 74.100 235.400 74.200 ;
        RECT 235.800 74.100 236.100 93.800 ;
        RECT 236.600 92.100 237.000 97.900 ;
        RECT 237.400 95.800 237.800 96.200 ;
        RECT 237.400 95.100 237.700 95.800 ;
        RECT 237.400 94.700 237.800 95.100 ;
        RECT 240.600 90.200 240.900 104.800 ;
        RECT 241.400 92.100 241.800 97.900 ;
        RECT 244.600 96.200 244.900 105.800 ;
        RECT 242.200 95.800 242.600 96.200 ;
        RECT 243.800 96.100 244.200 96.200 ;
        RECT 244.600 96.100 245.000 96.200 ;
        RECT 243.800 95.800 245.000 96.100 ;
        RECT 240.600 89.800 241.000 90.200 ;
        RECT 239.800 89.100 240.200 89.200 ;
        RECT 240.600 89.100 241.000 89.200 ;
        RECT 238.200 83.100 238.600 88.900 ;
        RECT 239.800 88.800 241.000 89.100 ;
        RECT 241.400 87.800 241.800 88.200 ;
        RECT 241.400 87.200 241.700 87.800 ;
        RECT 241.400 86.800 241.800 87.200 ;
        RECT 242.200 86.200 242.500 95.800 ;
        RECT 243.000 92.100 243.400 92.200 ;
        RECT 243.800 92.100 244.200 92.200 ;
        RECT 243.000 91.800 244.200 92.100 ;
        RECT 244.600 91.800 245.000 92.200 ;
        RECT 242.200 85.800 242.600 86.200 ;
        RECT 243.000 86.100 243.400 86.200 ;
        RECT 243.800 86.100 244.200 86.200 ;
        RECT 243.000 85.800 244.200 86.100 ;
        RECT 235.000 73.800 236.100 74.100 ;
        RECT 242.200 74.200 242.500 85.800 ;
        RECT 243.800 85.100 244.200 85.200 ;
        RECT 244.600 85.100 244.900 91.800 ;
        RECT 245.400 89.200 245.700 122.800 ;
        RECT 248.600 118.100 249.000 118.200 ;
        RECT 249.400 118.100 249.800 118.200 ;
        RECT 247.000 112.100 247.400 117.900 ;
        RECT 248.600 117.800 249.800 118.100 ;
        RECT 249.400 109.100 249.800 109.200 ;
        RECT 250.200 109.100 250.600 109.200 ;
        RECT 249.400 108.800 250.600 109.100 ;
        RECT 248.600 102.800 249.000 103.200 ;
        RECT 248.600 99.200 248.900 102.800 ;
        RECT 248.600 98.800 249.000 99.200 ;
        RECT 251.000 95.200 251.300 233.800 ;
        RECT 251.800 200.800 252.200 201.200 ;
        RECT 251.800 156.200 252.100 200.800 ;
        RECT 251.800 155.800 252.200 156.200 ;
        RECT 246.200 95.100 246.600 95.200 ;
        RECT 247.000 95.100 247.400 95.200 ;
        RECT 246.200 94.800 247.400 95.100 ;
        RECT 247.800 94.800 248.200 95.200 ;
        RECT 251.000 94.800 251.400 95.200 ;
        RECT 247.800 94.200 248.100 94.800 ;
        RECT 246.200 94.100 246.600 94.200 ;
        RECT 247.000 94.100 247.400 94.200 ;
        RECT 246.200 93.800 247.400 94.100 ;
        RECT 247.800 93.800 248.200 94.200 ;
        RECT 251.000 89.200 251.300 94.800 ;
        RECT 245.400 88.800 245.800 89.200 ;
        RECT 251.000 88.800 251.400 89.200 ;
        RECT 243.800 84.800 244.900 85.100 ;
        RECT 247.000 87.800 247.400 88.200 ;
        RECT 247.000 75.200 247.300 87.800 ;
        RECT 250.200 87.100 250.600 87.200 ;
        RECT 251.000 87.100 251.400 87.200 ;
        RECT 250.200 86.800 251.400 87.100 ;
        RECT 247.800 76.100 248.200 76.200 ;
        RECT 248.600 76.100 249.000 76.200 ;
        RECT 247.800 75.800 249.000 76.100 ;
        RECT 251.800 75.200 252.100 155.800 ;
        RECT 243.800 75.100 244.200 75.200 ;
        RECT 244.600 75.100 245.000 75.200 ;
        RECT 243.800 74.800 245.000 75.100 ;
        RECT 246.200 74.800 246.600 75.200 ;
        RECT 247.000 74.800 247.400 75.200 ;
        RECT 251.800 74.800 252.200 75.200 ;
        RECT 246.200 74.200 246.500 74.800 ;
        RECT 247.000 74.200 247.300 74.800 ;
        RECT 242.200 73.800 242.600 74.200 ;
        RECT 246.200 73.800 246.600 74.200 ;
        RECT 247.000 73.800 247.400 74.200 ;
        RECT 249.400 74.100 249.800 74.200 ;
        RECT 250.200 74.100 250.600 74.200 ;
        RECT 249.400 73.800 250.600 74.100 ;
        RECT 242.200 72.800 242.600 73.200 ;
        RECT 240.600 71.800 241.000 72.200 ;
        RECT 232.600 69.100 233.000 69.200 ;
        RECT 233.400 69.100 233.800 69.200 ;
        RECT 232.600 68.800 233.800 69.100 ;
        RECT 231.800 67.800 232.200 68.200 ;
        RECT 230.200 66.800 230.600 67.200 ;
        RECT 226.200 65.800 226.600 66.200 ;
        RECT 228.600 65.800 229.000 66.200 ;
        RECT 229.400 65.800 229.800 66.200 ;
        RECT 226.200 61.800 226.600 62.200 ;
        RECT 221.400 59.800 221.800 60.200 ;
        RECT 221.400 54.700 221.800 55.100 ;
        RECT 221.400 54.200 221.700 54.700 ;
        RECT 221.400 53.800 221.800 54.200 ;
        RECT 222.200 52.100 222.600 57.900 ;
        RECT 223.800 53.100 224.200 55.900 ;
        RECT 226.200 54.200 226.500 61.800 ;
        RECT 227.800 59.800 228.200 60.200 ;
        RECT 227.800 59.200 228.100 59.800 ;
        RECT 228.600 59.200 228.900 65.800 ;
        RECT 229.400 65.200 229.700 65.800 ;
        RECT 229.400 64.800 229.800 65.200 ;
        RECT 227.800 58.800 228.200 59.200 ;
        RECT 228.600 58.800 229.000 59.200 ;
        RECT 228.600 57.800 229.000 58.200 ;
        RECT 227.800 56.800 228.200 57.200 ;
        RECT 227.000 54.800 227.400 55.200 ;
        RECT 227.000 54.200 227.300 54.800 ;
        RECT 224.600 54.100 225.000 54.200 ;
        RECT 225.400 54.100 225.800 54.200 ;
        RECT 224.600 53.800 225.800 54.100 ;
        RECT 226.200 53.800 226.600 54.200 ;
        RECT 227.000 53.800 227.400 54.200 ;
        RECT 224.600 52.800 225.000 53.200 ;
        RECT 223.800 50.800 224.200 51.200 ;
        RECT 223.800 48.200 224.100 50.800 ;
        RECT 224.600 49.200 224.900 52.800 ;
        RECT 224.600 48.800 225.000 49.200 ;
        RECT 220.600 47.800 221.000 48.200 ;
        RECT 223.000 47.800 223.400 48.200 ;
        RECT 223.800 47.800 224.200 48.200 ;
        RECT 219.800 46.800 220.200 47.200 ;
        RECT 219.800 46.200 220.100 46.800 ;
        RECT 219.800 45.800 220.200 46.200 ;
        RECT 219.800 44.800 220.200 45.200 ;
        RECT 219.800 44.200 220.100 44.800 ;
        RECT 219.800 43.800 220.200 44.200 ;
        RECT 219.800 34.800 220.200 35.200 ;
        RECT 219.000 33.800 219.400 34.200 ;
        RECT 218.200 28.800 218.600 29.200 ;
        RECT 215.000 27.100 215.400 27.200 ;
        RECT 215.800 27.100 216.200 27.200 ;
        RECT 215.000 26.800 216.200 27.100 ;
        RECT 215.000 25.800 215.400 26.200 ;
        RECT 216.600 26.100 217.000 26.200 ;
        RECT 217.400 26.100 217.800 26.200 ;
        RECT 216.600 25.800 217.800 26.100 ;
        RECT 215.000 25.200 215.300 25.800 ;
        RECT 214.200 24.800 214.600 25.200 ;
        RECT 215.000 24.800 215.400 25.200 ;
        RECT 211.800 22.800 212.200 23.200 ;
        RECT 211.800 19.200 212.100 22.800 ;
        RECT 211.800 18.800 212.200 19.200 ;
        RECT 210.200 15.800 210.600 16.200 ;
        RECT 213.400 15.800 213.800 16.200 ;
        RECT 218.200 15.800 218.600 16.200 ;
        RECT 210.200 15.200 210.500 15.800 ;
        RECT 213.400 15.200 213.700 15.800 ;
        RECT 218.200 15.200 218.500 15.800 ;
        RECT 204.600 14.800 205.000 15.200 ;
        RECT 205.400 14.800 205.800 15.200 ;
        RECT 206.200 14.800 206.600 15.200 ;
        RECT 209.400 14.800 209.800 15.200 ;
        RECT 210.200 14.800 210.600 15.200 ;
        RECT 211.000 14.800 211.400 15.200 ;
        RECT 213.400 14.800 213.800 15.200 ;
        RECT 215.000 15.100 215.400 15.200 ;
        RECT 215.800 15.100 216.200 15.200 ;
        RECT 215.000 14.800 216.200 15.100 ;
        RECT 218.200 14.800 218.600 15.200 ;
        RECT 201.400 13.800 201.800 14.200 ;
        RECT 205.400 13.200 205.700 14.800 ;
        RECT 207.000 14.100 207.400 14.200 ;
        RECT 207.800 14.100 208.200 14.200 ;
        RECT 207.000 13.800 208.200 14.100 ;
        RECT 200.600 12.800 201.000 13.200 ;
        RECT 205.400 12.800 205.800 13.200 ;
        RECT 200.600 7.200 200.900 12.800 ;
        RECT 205.400 10.200 205.700 12.800 ;
        RECT 205.400 9.800 205.800 10.200 ;
        RECT 209.400 9.200 209.700 14.800 ;
        RECT 211.000 13.200 211.300 14.800 ;
        RECT 219.800 14.200 220.100 34.800 ;
        RECT 220.600 34.200 220.900 47.800 ;
        RECT 223.000 47.200 223.300 47.800 ;
        RECT 223.000 46.800 223.400 47.200 ;
        RECT 226.200 47.100 226.500 53.800 ;
        RECT 227.000 48.200 227.300 53.800 ;
        RECT 227.800 49.200 228.100 56.800 ;
        RECT 227.800 48.800 228.200 49.200 ;
        RECT 227.000 47.800 227.400 48.200 ;
        RECT 225.400 46.800 226.500 47.100 ;
        RECT 227.800 46.800 228.200 47.200 ;
        RECT 225.400 46.200 225.700 46.800 ;
        RECT 222.200 45.800 222.600 46.200 ;
        RECT 225.400 45.800 225.800 46.200 ;
        RECT 226.200 45.800 226.600 46.200 ;
        RECT 227.000 45.800 227.400 46.200 ;
        RECT 222.200 44.200 222.500 45.800 ;
        RECT 226.200 45.200 226.500 45.800 ;
        RECT 226.200 44.800 226.600 45.200 ;
        RECT 222.200 43.800 222.600 44.200 ;
        RECT 223.800 36.800 224.200 37.200 ;
        RECT 223.800 36.200 224.100 36.800 ;
        RECT 221.400 35.800 221.800 36.200 ;
        RECT 223.800 35.800 224.200 36.200 ;
        RECT 221.400 35.200 221.700 35.800 ;
        RECT 221.400 34.800 221.800 35.200 ;
        RECT 227.000 34.200 227.300 45.800 ;
        RECT 220.600 33.800 221.000 34.200 ;
        RECT 226.200 33.800 226.600 34.200 ;
        RECT 227.000 33.800 227.400 34.200 ;
        RECT 223.000 31.800 223.400 32.200 ;
        RECT 220.600 23.100 221.000 28.900 ;
        RECT 223.000 27.200 223.300 31.800 ;
        RECT 226.200 29.200 226.500 33.800 ;
        RECT 223.000 26.800 223.400 27.200 ;
        RECT 222.200 25.800 222.600 26.200 ;
        RECT 223.800 25.800 224.200 26.200 ;
        RECT 221.400 19.800 221.800 20.200 ;
        RECT 221.400 15.200 221.700 19.800 ;
        RECT 221.400 14.800 221.800 15.200 ;
        RECT 214.200 14.100 214.600 14.200 ;
        RECT 215.000 14.100 215.400 14.200 ;
        RECT 214.200 13.800 215.400 14.100 ;
        RECT 216.600 13.800 217.000 14.200 ;
        RECT 219.800 13.800 220.200 14.200 ;
        RECT 220.600 14.100 221.000 14.200 ;
        RECT 221.400 14.100 221.800 14.200 ;
        RECT 220.600 13.800 221.800 14.100 ;
        RECT 211.000 12.800 211.400 13.200 ;
        RECT 211.000 9.800 211.400 10.200 ;
        RECT 211.000 9.200 211.300 9.800 ;
        RECT 195.000 6.800 195.400 7.200 ;
        RECT 197.400 7.100 197.800 7.200 ;
        RECT 198.200 7.100 198.600 7.200 ;
        RECT 197.400 6.800 198.600 7.100 ;
        RECT 200.600 6.800 201.000 7.200 ;
        RECT 195.800 5.800 196.200 6.200 ;
        RECT 195.800 3.200 196.100 5.800 ;
        RECT 198.200 4.800 198.600 5.200 ;
        RECT 202.200 5.100 202.600 7.900 ;
        RECT 198.200 3.200 198.500 4.800 ;
        RECT 195.800 2.800 196.200 3.200 ;
        RECT 198.200 2.800 198.600 3.200 ;
        RECT 203.800 3.100 204.200 8.900 ;
        RECT 206.200 7.800 206.600 8.200 ;
        RECT 206.200 7.200 206.500 7.800 ;
        RECT 204.600 6.800 205.000 7.200 ;
        RECT 206.200 6.800 206.600 7.200 ;
        RECT 204.600 6.300 204.900 6.800 ;
        RECT 204.600 5.900 205.000 6.300 ;
        RECT 208.600 3.100 209.000 8.900 ;
        RECT 209.400 8.800 209.800 9.200 ;
        RECT 211.000 8.800 211.400 9.200 ;
        RECT 211.800 5.100 212.200 7.900 ;
        RECT 213.400 3.100 213.800 8.900 ;
        RECT 215.800 7.800 216.200 8.200 ;
        RECT 215.800 7.200 216.100 7.800 ;
        RECT 215.800 6.800 216.200 7.200 ;
        RECT 216.600 6.200 216.900 13.800 ;
        RECT 219.800 9.100 220.100 13.800 ;
        RECT 220.600 9.100 221.000 9.200 ;
        RECT 216.600 5.800 217.000 6.200 ;
        RECT 218.200 3.100 218.600 8.900 ;
        RECT 219.800 8.800 221.000 9.100 ;
        RECT 221.400 7.200 221.700 13.800 ;
        RECT 222.200 8.200 222.500 25.800 ;
        RECT 223.800 25.200 224.100 25.800 ;
        RECT 223.800 24.800 224.200 25.200 ;
        RECT 225.400 23.100 225.800 28.900 ;
        RECT 226.200 28.800 226.600 29.200 ;
        RECT 227.000 25.100 227.400 27.900 ;
        RECT 227.800 27.200 228.100 46.800 ;
        RECT 228.600 29.200 228.900 57.800 ;
        RECT 229.400 38.100 229.700 64.800 ;
        RECT 230.200 60.200 230.500 66.800 ;
        RECT 231.800 64.800 232.200 65.200 ;
        RECT 231.000 61.800 231.400 62.200 ;
        RECT 230.200 59.800 230.600 60.200 ;
        RECT 230.200 52.100 230.600 57.900 ;
        RECT 231.000 56.200 231.300 61.800 ;
        RECT 231.800 61.200 232.100 64.800 ;
        RECT 235.000 63.100 235.400 68.900 ;
        RECT 235.800 67.800 236.200 68.200 ;
        RECT 239.000 67.800 239.400 68.200 ;
        RECT 235.800 67.200 236.100 67.800 ;
        RECT 235.800 66.800 236.200 67.200 ;
        RECT 239.000 66.300 239.300 67.800 ;
        RECT 239.000 65.900 239.400 66.300 ;
        RECT 239.800 63.100 240.200 68.900 ;
        RECT 240.600 67.200 240.900 71.800 ;
        RECT 242.200 69.200 242.500 72.800 ;
        RECT 245.400 71.800 245.800 72.200 ;
        RECT 242.200 68.800 242.600 69.200 ;
        RECT 240.600 66.800 241.000 67.200 ;
        RECT 241.400 65.100 241.800 67.900 ;
        RECT 242.200 65.100 242.600 67.900 ;
        RECT 243.800 63.100 244.200 68.900 ;
        RECT 245.400 68.200 245.700 71.800 ;
        RECT 245.400 67.800 245.800 68.200 ;
        RECT 245.400 66.800 245.800 67.200 ;
        RECT 245.400 66.200 245.700 66.800 ;
        RECT 245.400 65.800 245.800 66.200 ;
        RECT 246.200 62.200 246.500 73.800 ;
        RECT 247.800 71.800 248.200 72.200 ;
        RECT 246.200 61.800 246.600 62.200 ;
        RECT 231.800 60.800 232.200 61.200 ;
        RECT 239.000 60.800 239.400 61.200 ;
        RECT 232.600 56.800 233.000 57.200 ;
        RECT 231.000 55.800 231.400 56.200 ;
        RECT 231.000 55.100 231.400 55.200 ;
        RECT 231.800 55.100 232.200 55.200 ;
        RECT 231.000 54.800 232.200 55.100 ;
        RECT 231.000 45.800 231.400 46.200 ;
        RECT 229.400 37.800 230.500 38.100 ;
        RECT 229.400 36.800 229.800 37.200 ;
        RECT 229.400 35.200 229.700 36.800 ;
        RECT 230.200 35.200 230.500 37.800 ;
        RECT 229.400 34.800 229.800 35.200 ;
        RECT 230.200 34.800 230.600 35.200 ;
        RECT 231.000 33.200 231.300 45.800 ;
        RECT 232.600 35.200 232.900 56.800 ;
        RECT 233.400 55.100 233.800 55.200 ;
        RECT 233.400 54.800 234.600 55.100 ;
        RECT 234.200 54.700 234.600 54.800 ;
        RECT 234.200 51.800 234.600 52.200 ;
        RECT 235.000 52.100 235.400 57.900 ;
        RECT 237.400 56.800 237.800 57.200 ;
        RECT 237.400 56.200 237.700 56.800 ;
        RECT 235.800 53.800 236.200 54.200 ;
        RECT 234.200 47.100 234.500 51.800 ;
        RECT 235.800 47.200 236.100 53.800 ;
        RECT 236.600 53.100 237.000 55.900 ;
        RECT 237.400 55.800 237.800 56.200 ;
        RECT 239.000 55.200 239.300 60.800 ;
        RECT 239.800 59.100 240.200 59.200 ;
        RECT 240.600 59.100 241.000 59.200 ;
        RECT 247.800 59.100 248.100 71.800 ;
        RECT 251.000 69.800 251.400 70.200 ;
        RECT 251.000 69.200 251.300 69.800 ;
        RECT 248.600 63.100 249.000 68.900 ;
        RECT 251.000 68.800 251.400 69.200 ;
        RECT 239.800 58.800 241.000 59.100 ;
        RECT 247.000 58.800 248.100 59.100 ;
        RECT 237.400 55.100 237.800 55.200 ;
        RECT 238.200 55.100 238.600 55.200 ;
        RECT 237.400 54.800 238.600 55.100 ;
        RECT 239.000 54.800 239.400 55.200 ;
        RECT 239.800 54.100 240.200 54.200 ;
        RECT 240.600 54.100 241.000 54.200 ;
        RECT 239.800 53.800 241.000 54.100 ;
        RECT 243.000 52.100 243.400 57.900 ;
        RECT 247.000 55.100 247.300 58.800 ;
        RECT 247.000 54.700 247.400 55.100 ;
        RECT 246.200 53.800 246.600 54.200 ;
        RECT 240.600 48.800 241.000 49.200 ;
        RECT 240.600 47.200 240.900 48.800 ;
        RECT 234.200 46.800 235.300 47.100 ;
        RECT 235.000 46.200 235.300 46.800 ;
        RECT 235.800 46.800 236.200 47.200 ;
        RECT 238.200 47.100 238.600 47.200 ;
        RECT 239.000 47.100 239.400 47.200 ;
        RECT 238.200 46.800 239.400 47.100 ;
        RECT 240.600 46.800 241.000 47.200 ;
        RECT 233.400 46.100 233.800 46.200 ;
        RECT 234.200 46.100 234.600 46.200 ;
        RECT 233.400 45.800 234.600 46.100 ;
        RECT 235.000 45.800 235.400 46.200 ;
        RECT 235.800 35.200 236.100 46.800 ;
        RECT 236.600 46.100 237.000 46.200 ;
        RECT 237.400 46.100 237.800 46.200 ;
        RECT 236.600 45.800 237.800 46.100 ;
        RECT 239.000 45.800 239.400 46.200 ;
        RECT 239.000 45.200 239.300 45.800 ;
        RECT 239.000 44.800 239.400 45.200 ;
        RECT 241.400 45.100 241.800 47.900 ;
        RECT 242.200 46.800 242.600 47.200 ;
        RECT 242.200 42.100 242.500 46.800 ;
        RECT 243.000 43.100 243.400 48.900 ;
        RECT 243.800 46.800 244.200 47.200 ;
        RECT 243.800 46.300 244.100 46.800 ;
        RECT 243.800 45.900 244.200 46.300 ;
        RECT 242.200 41.800 243.300 42.100 ;
        RECT 241.400 36.800 241.800 37.200 ;
        RECT 237.400 35.800 237.800 36.200 ;
        RECT 239.800 36.100 240.200 36.200 ;
        RECT 240.600 36.100 241.000 36.200 ;
        RECT 239.800 35.800 241.000 36.100 ;
        RECT 237.400 35.200 237.700 35.800 ;
        RECT 232.600 34.800 233.000 35.200 ;
        RECT 235.800 34.800 236.200 35.200 ;
        RECT 237.400 34.800 237.800 35.200 ;
        RECT 239.800 34.800 240.200 35.200 ;
        RECT 232.600 34.200 232.900 34.800 ;
        RECT 239.800 34.200 240.100 34.800 ;
        RECT 232.600 33.800 233.000 34.200 ;
        RECT 234.200 34.100 234.600 34.200 ;
        RECT 235.000 34.100 235.400 34.200 ;
        RECT 234.200 33.800 235.400 34.100 ;
        RECT 236.600 33.800 237.000 34.200 ;
        RECT 239.800 33.800 240.200 34.200 ;
        RECT 231.000 32.800 231.400 33.200 ;
        RECT 231.000 29.200 231.300 32.800 ;
        RECT 234.200 31.800 234.600 32.200 ;
        RECT 228.600 28.800 229.000 29.200 ;
        RECT 229.400 29.100 229.800 29.200 ;
        RECT 230.200 29.100 230.600 29.200 ;
        RECT 229.400 28.800 230.600 29.100 ;
        RECT 231.000 28.800 231.400 29.200 ;
        RECT 227.800 26.800 228.200 27.200 ;
        RECT 229.400 24.800 229.800 25.200 ;
        RECT 229.400 24.200 229.700 24.800 ;
        RECT 229.400 23.800 229.800 24.200 ;
        RECT 232.600 23.100 233.000 28.900 ;
        RECT 234.200 26.200 234.500 31.800 ;
        RECT 236.600 27.200 236.900 33.800 ;
        RECT 239.000 29.100 239.400 29.200 ;
        RECT 239.800 29.100 240.200 29.200 ;
        RECT 235.800 26.800 236.200 27.200 ;
        RECT 236.600 26.800 237.000 27.200 ;
        RECT 235.800 26.200 236.100 26.800 ;
        RECT 234.200 25.800 234.600 26.200 ;
        RECT 235.800 25.800 236.200 26.200 ;
        RECT 223.800 19.800 224.200 20.200 ;
        RECT 223.800 16.200 224.100 19.800 ;
        RECT 236.600 19.200 236.900 26.800 ;
        RECT 237.400 23.100 237.800 28.900 ;
        RECT 239.000 28.800 240.200 29.100 ;
        RECT 239.000 25.100 239.400 27.900 ;
        RECT 236.600 18.800 237.000 19.200 ;
        RECT 225.400 16.800 225.800 17.200 ;
        RECT 225.400 16.200 225.700 16.800 ;
        RECT 223.800 15.800 224.200 16.200 ;
        RECT 225.400 15.800 225.800 16.200 ;
        RECT 223.800 14.800 224.200 15.200 ;
        RECT 223.800 14.200 224.100 14.800 ;
        RECT 225.400 14.200 225.700 15.800 ;
        RECT 223.800 13.800 224.200 14.200 ;
        RECT 225.400 13.800 225.800 14.200 ;
        RECT 227.000 12.800 227.400 13.200 ;
        RECT 227.000 9.200 227.300 12.800 ;
        RECT 228.600 12.100 229.000 17.900 ;
        RECT 231.000 15.100 231.400 15.200 ;
        RECT 231.800 15.100 232.200 15.200 ;
        RECT 231.000 14.800 232.200 15.100 ;
        RECT 233.400 12.100 233.800 17.900 ;
        RECT 240.600 16.200 240.900 35.800 ;
        RECT 241.400 34.200 241.700 36.800 ;
        RECT 241.400 33.800 241.800 34.200 ;
        RECT 242.200 33.100 242.600 35.900 ;
        RECT 243.000 34.200 243.300 41.800 ;
        RECT 243.000 33.800 243.400 34.200 ;
        RECT 243.000 33.200 243.300 33.800 ;
        RECT 243.000 32.800 243.400 33.200 ;
        RECT 243.800 32.100 244.200 37.900 ;
        RECT 244.600 35.800 245.000 36.200 ;
        RECT 244.600 35.100 244.900 35.800 ;
        RECT 244.600 34.700 245.000 35.100 ;
        RECT 242.200 23.100 242.600 28.900 ;
        RECT 246.200 28.200 246.500 53.800 ;
        RECT 247.800 52.100 248.200 57.900 ;
        RECT 249.400 53.100 249.800 55.900 ;
        RECT 249.400 49.100 249.800 49.200 ;
        RECT 250.200 49.100 250.600 49.200 ;
        RECT 247.800 43.100 248.200 48.900 ;
        RECT 249.400 48.800 250.600 49.100 ;
        RECT 251.800 44.200 252.100 74.800 ;
        RECT 251.800 43.800 252.200 44.200 ;
        RECT 248.600 32.100 249.000 37.900 ;
        RECT 250.200 37.100 250.600 37.200 ;
        RECT 251.000 37.100 251.400 37.200 ;
        RECT 250.200 36.800 251.400 37.100 ;
        RECT 251.000 35.800 251.400 36.200 ;
        RECT 250.200 29.800 250.600 30.200 ;
        RECT 246.200 27.800 246.600 28.200 ;
        RECT 243.800 25.800 244.200 26.200 ;
        RECT 244.600 26.100 245.000 26.200 ;
        RECT 245.400 26.100 245.800 26.200 ;
        RECT 244.600 25.800 245.800 26.100 ;
        RECT 243.800 19.200 244.100 25.800 ;
        RECT 247.000 23.100 247.400 28.900 ;
        RECT 248.600 25.100 249.000 27.900 ;
        RECT 249.400 27.800 249.800 28.200 ;
        RECT 249.400 27.200 249.700 27.800 ;
        RECT 249.400 26.800 249.800 27.200 ;
        RECT 250.200 26.200 250.500 29.800 ;
        RECT 250.200 25.800 250.600 26.200 ;
        RECT 251.000 19.200 251.300 35.800 ;
        RECT 251.800 30.200 252.100 43.800 ;
        RECT 251.800 29.800 252.200 30.200 ;
        RECT 251.800 28.800 252.200 29.200 ;
        RECT 251.800 28.200 252.100 28.800 ;
        RECT 251.800 27.800 252.200 28.200 ;
        RECT 251.800 25.800 252.200 26.200 ;
        RECT 251.800 25.200 252.100 25.800 ;
        RECT 251.800 24.800 252.200 25.200 ;
        RECT 251.800 23.800 252.200 24.200 ;
        RECT 243.800 18.800 244.200 19.200 ;
        RECT 251.000 18.800 251.400 19.200 ;
        RECT 234.200 14.800 234.600 15.200 ;
        RECT 234.200 14.200 234.500 14.800 ;
        RECT 234.200 13.800 234.600 14.200 ;
        RECT 235.000 13.100 235.400 15.900 ;
        RECT 240.600 15.800 241.000 16.200 ;
        RECT 249.400 16.100 249.800 16.200 ;
        RECT 250.200 16.100 250.600 16.200 ;
        RECT 249.400 15.800 250.600 16.100 ;
        RECT 235.800 14.800 236.200 15.200 ;
        RECT 235.800 14.200 236.100 14.800 ;
        RECT 251.800 14.200 252.100 23.800 ;
        RECT 235.800 13.800 236.200 14.200 ;
        RECT 242.200 14.100 242.600 14.200 ;
        RECT 243.000 14.100 243.400 14.200 ;
        RECT 242.200 13.800 243.400 14.100 ;
        RECT 251.800 13.800 252.200 14.200 ;
        RECT 227.000 8.800 227.400 9.200 ;
        RECT 222.200 7.800 222.600 8.200 ;
        RECT 221.400 6.800 221.800 7.200 ;
        RECT 223.800 7.100 224.200 7.200 ;
        RECT 224.600 7.100 225.000 7.200 ;
        RECT 223.800 6.800 225.000 7.100 ;
        RECT 221.400 6.100 221.800 6.200 ;
        RECT 222.200 6.100 222.600 6.200 ;
        RECT 221.400 5.800 222.600 6.100 ;
        RECT 224.600 5.800 225.000 6.200 ;
        RECT 224.600 5.200 224.900 5.800 ;
        RECT 224.600 4.800 225.000 5.200 ;
        RECT 229.400 3.100 229.800 8.900 ;
        RECT 232.600 6.800 233.000 7.200 ;
        RECT 232.600 6.200 232.900 6.800 ;
        RECT 232.600 5.800 233.000 6.200 ;
        RECT 234.200 3.100 234.600 8.900 ;
        RECT 235.000 7.800 235.400 8.200 ;
        RECT 235.000 7.200 235.300 7.800 ;
        RECT 235.000 6.800 235.400 7.200 ;
        RECT 235.800 5.100 236.200 7.900 ;
        RECT 242.200 7.200 242.500 13.800 ;
        RECT 243.800 9.100 244.200 9.200 ;
        RECT 244.600 9.100 245.000 9.200 ;
        RECT 243.800 8.800 245.000 9.100 ;
        RECT 247.800 9.100 248.200 9.200 ;
        RECT 248.600 9.100 249.000 9.200 ;
        RECT 247.800 8.800 249.000 9.100 ;
        RECT 242.200 6.800 242.600 7.200 ;
        RECT 243.000 7.100 243.400 7.200 ;
        RECT 243.800 7.100 244.200 7.200 ;
        RECT 243.000 6.800 244.200 7.100 ;
      LAYER via2 ;
        RECT 5.400 233.800 5.800 234.200 ;
        RECT 1.400 221.800 1.800 222.200 ;
        RECT 19.000 225.800 19.400 226.200 ;
        RECT 1.400 218.800 1.800 219.200 ;
        RECT 1.400 208.800 1.800 209.200 ;
        RECT 1.400 186.800 1.800 187.200 ;
        RECT 12.600 205.800 13.000 206.200 ;
        RECT 17.400 205.800 17.800 206.200 ;
        RECT 7.800 185.800 8.200 186.200 ;
        RECT 3.000 184.800 3.400 185.200 ;
        RECT 1.400 177.800 1.800 178.200 ;
        RECT 14.200 175.800 14.600 176.200 ;
        RECT 11.800 174.800 12.200 175.200 ;
        RECT 18.200 175.800 18.600 176.200 ;
        RECT 14.200 173.800 14.600 174.200 ;
        RECT 11.800 165.800 12.200 166.200 ;
        RECT 5.400 154.800 5.800 155.200 ;
        RECT 55.800 236.800 56.200 237.200 ;
        RECT 55.800 233.800 56.200 234.200 ;
        RECT 41.400 224.800 41.800 225.200 ;
        RECT 31.800 195.800 32.200 196.200 ;
        RECT 22.200 173.800 22.600 174.200 ;
        RECT 19.800 165.800 20.200 166.200 ;
        RECT 29.400 174.800 29.800 175.200 ;
        RECT 33.400 185.800 33.800 186.200 ;
        RECT 30.200 167.800 30.600 168.200 ;
        RECT 75.000 234.800 75.400 235.200 ;
        RECT 75.800 233.800 76.200 234.200 ;
        RECT 65.400 195.800 65.800 196.200 ;
        RECT 22.200 154.800 22.600 155.200 ;
        RECT 11.000 153.800 11.400 154.200 ;
        RECT 3.800 138.800 4.200 139.200 ;
        RECT 12.600 146.800 13.000 147.200 ;
        RECT 15.000 145.800 15.400 146.200 ;
        RECT 20.600 145.800 21.000 146.200 ;
        RECT 8.600 134.800 9.000 135.200 ;
        RECT 16.600 134.800 17.000 135.200 ;
        RECT 15.000 133.800 15.400 134.200 ;
        RECT 11.000 124.800 11.400 125.200 ;
        RECT 17.400 125.800 17.800 126.200 ;
        RECT 11.800 114.800 12.200 115.200 ;
        RECT 26.200 153.800 26.600 154.200 ;
        RECT 27.800 145.800 28.200 146.200 ;
        RECT 25.400 141.800 25.800 142.200 ;
        RECT 43.000 164.800 43.400 165.200 ;
        RECT 69.400 215.800 69.800 216.200 ;
        RECT 72.600 214.800 73.000 215.200 ;
        RECT 69.400 205.800 69.800 206.200 ;
        RECT 71.800 213.800 72.200 214.200 ;
        RECT 112.600 235.800 113.000 236.200 ;
        RECT 86.200 224.800 86.600 225.200 ;
        RECT 70.200 194.800 70.600 195.200 ;
        RECT 95.800 225.800 96.200 226.200 ;
        RECT 92.600 214.800 93.000 215.200 ;
        RECT 91.000 211.800 91.400 212.200 ;
        RECT 80.600 194.800 81.000 195.200 ;
        RECT 69.400 182.800 69.800 183.200 ;
        RECT 59.000 177.800 59.400 178.200 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 63.000 168.800 63.400 169.200 ;
        RECT 99.000 211.800 99.400 212.200 ;
        RECT 107.800 226.800 108.200 227.200 ;
        RECT 101.400 195.800 101.800 196.200 ;
        RECT 95.800 194.800 96.200 195.200 ;
        RECT 93.400 191.800 93.800 192.200 ;
        RECT 100.600 194.800 101.000 195.200 ;
        RECT 80.600 185.800 81.000 186.200 ;
        RECT 86.200 186.800 86.600 187.200 ;
        RECT 87.800 184.800 88.200 185.200 ;
        RECT 64.600 165.800 65.000 166.200 ;
        RECT 70.200 165.800 70.600 166.200 ;
        RECT 43.800 145.800 44.200 146.200 ;
        RECT 47.800 145.800 48.200 146.200 ;
        RECT 65.400 155.800 65.800 156.200 ;
        RECT 45.400 138.800 45.800 139.200 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 23.000 116.800 23.400 117.200 ;
        RECT 7.800 94.800 8.200 95.200 ;
        RECT 20.600 95.800 21.000 96.200 ;
        RECT 8.600 84.800 9.000 85.200 ;
        RECT 1.400 66.800 1.800 67.200 ;
        RECT 5.400 65.800 5.800 66.200 ;
        RECT 20.600 88.800 21.000 89.200 ;
        RECT 19.800 83.800 20.200 84.200 ;
        RECT 28.600 115.800 29.000 116.200 ;
        RECT 38.200 114.800 38.600 115.200 ;
        RECT 26.200 95.800 26.600 96.200 ;
        RECT 24.600 93.800 25.000 94.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 24.600 74.800 25.000 75.200 ;
        RECT 19.000 73.800 19.400 74.200 ;
        RECT 25.400 73.800 25.800 74.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.000 44.800 15.400 45.200 ;
        RECT 1.400 26.800 1.800 27.200 ;
        RECT 11.000 24.800 11.400 25.200 ;
        RECT 43.800 115.800 44.200 116.200 ;
        RECT 43.800 114.800 44.200 115.200 ;
        RECT 48.600 116.800 49.000 117.200 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 63.800 133.800 64.200 134.200 ;
        RECT 65.400 126.800 65.800 127.200 ;
        RECT 62.200 124.800 62.600 125.200 ;
        RECT 48.600 106.800 49.000 107.200 ;
        RECT 59.000 115.800 59.400 116.200 ;
        RECT 59.000 114.800 59.400 115.200 ;
        RECT 38.200 85.800 38.600 86.200 ;
        RECT 33.400 75.800 33.800 76.200 ;
        RECT 128.600 235.800 129.000 236.200 ;
        RECT 128.600 233.800 129.000 234.200 ;
        RECT 118.200 225.800 118.600 226.200 ;
        RECT 157.400 234.800 157.800 235.200 ;
        RECT 139.800 224.800 140.200 225.200 ;
        RECT 131.000 213.800 131.400 214.200 ;
        RECT 107.000 185.800 107.400 186.200 ;
        RECT 162.200 227.800 162.600 228.200 ;
        RECT 146.200 211.800 146.600 212.200 ;
        RECT 127.800 205.800 128.200 206.200 ;
        RECT 118.200 191.800 118.600 192.200 ;
        RECT 111.000 186.800 111.400 187.200 ;
        RECT 115.000 184.800 115.400 185.200 ;
        RECT 105.400 176.800 105.800 177.200 ;
        RECT 116.600 175.800 117.000 176.200 ;
        RECT 108.600 165.800 109.000 166.200 ;
        RECT 116.600 165.800 117.000 166.200 ;
        RECT 75.800 145.800 76.200 146.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 84.600 134.800 85.000 135.200 ;
        RECT 75.000 115.800 75.400 116.200 ;
        RECT 73.400 104.800 73.800 105.200 ;
        RECT 102.200 153.800 102.600 154.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 65.400 85.800 65.800 86.200 ;
        RECT 28.600 53.800 29.000 54.200 ;
        RECT 58.200 66.800 58.600 67.200 ;
        RECT 78.200 94.800 78.600 95.200 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 63.000 65.800 63.400 66.200 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 35.800 46.800 36.200 47.200 ;
        RECT 36.600 43.800 37.000 44.200 ;
        RECT 47.000 54.800 47.400 55.200 ;
        RECT 15.000 14.800 15.400 15.200 ;
        RECT 19.800 13.800 20.200 14.200 ;
        RECT 39.800 34.800 40.200 35.200 ;
        RECT 44.600 34.800 45.000 35.200 ;
        RECT 40.600 33.800 41.000 34.200 ;
        RECT 41.400 22.800 41.800 23.200 ;
        RECT 43.800 18.800 44.200 19.200 ;
        RECT 62.200 53.800 62.600 54.200 ;
        RECT 63.800 53.800 64.200 54.200 ;
        RECT 60.600 52.800 61.000 53.200 ;
        RECT 85.400 84.800 85.800 85.200 ;
        RECT 107.800 153.800 108.200 154.200 ;
        RECT 108.600 151.800 109.000 152.200 ;
        RECT 118.200 154.800 118.600 155.200 ;
        RECT 106.200 134.800 106.600 135.200 ;
        RECT 114.200 135.800 114.600 136.200 ;
        RECT 140.600 194.800 141.000 195.200 ;
        RECT 147.000 194.800 147.400 195.200 ;
        RECT 131.800 173.800 132.200 174.200 ;
        RECT 149.400 193.800 149.800 194.200 ;
        RECT 147.800 188.800 148.200 189.200 ;
        RECT 152.600 186.800 153.000 187.200 ;
        RECT 160.600 196.800 161.000 197.200 ;
        RECT 145.400 174.800 145.800 175.200 ;
        RECT 133.400 154.800 133.800 155.200 ;
        RECT 126.200 153.800 126.600 154.200 ;
        RECT 107.000 115.800 107.400 116.200 ;
        RECT 155.000 175.800 155.400 176.200 ;
        RECT 182.200 228.800 182.600 229.200 ;
        RECT 180.600 214.800 181.000 215.200 ;
        RECT 199.000 233.800 199.400 234.200 ;
        RECT 195.000 208.800 195.400 209.200 ;
        RECT 190.200 206.800 190.600 207.200 ;
        RECT 194.200 205.800 194.600 206.200 ;
        RECT 193.400 194.800 193.800 195.200 ;
        RECT 178.200 182.800 178.600 183.200 ;
        RECT 194.200 191.800 194.600 192.200 ;
        RECT 221.400 235.800 221.800 236.200 ;
        RECT 227.000 234.800 227.400 235.200 ;
        RECT 203.800 191.800 204.200 192.200 ;
        RECT 160.600 165.800 161.000 166.200 ;
        RECT 144.600 155.800 145.000 156.200 ;
        RECT 148.600 155.800 149.000 156.200 ;
        RECT 159.000 155.800 159.400 156.200 ;
        RECT 147.000 153.800 147.400 154.200 ;
        RECT 111.800 104.800 112.200 105.200 ;
        RECT 107.000 94.700 107.400 95.100 ;
        RECT 96.600 86.800 97.000 87.200 ;
        RECT 92.600 73.800 93.000 74.200 ;
        RECT 90.200 66.800 90.600 67.200 ;
        RECT 93.400 66.800 93.800 67.200 ;
        RECT 82.200 65.800 82.600 66.200 ;
        RECT 91.000 65.800 91.400 66.200 ;
        RECT 85.400 58.800 85.800 59.200 ;
        RECT 71.800 54.700 72.200 55.100 ;
        RECT 80.600 54.800 81.000 55.200 ;
        RECT 91.800 54.800 92.200 55.200 ;
        RECT 95.800 54.800 96.200 55.200 ;
        RECT 71.000 48.800 71.400 49.200 ;
        RECT 73.400 46.800 73.800 47.200 ;
        RECT 72.600 45.800 73.000 46.200 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 59.000 26.800 59.400 27.200 ;
        RECT 43.800 6.800 44.200 7.200 ;
        RECT 58.200 25.800 58.600 26.200 ;
        RECT 60.600 24.800 61.000 25.200 ;
        RECT 73.400 25.800 73.800 26.200 ;
        RECT 79.000 26.800 79.400 27.200 ;
        RECT 92.600 48.800 93.000 49.200 ;
        RECT 88.600 46.800 89.000 47.200 ;
        RECT 91.000 45.800 91.400 46.200 ;
        RECT 103.800 74.800 104.200 75.200 ;
        RECT 107.800 73.800 108.200 74.200 ;
        RECT 99.800 56.800 100.200 57.200 ;
        RECT 89.400 32.800 89.800 33.200 ;
        RECT 107.000 67.800 107.400 68.200 ;
        RECT 131.800 104.800 132.200 105.200 ;
        RECT 123.800 94.000 124.200 94.400 ;
        RECT 115.800 74.800 116.200 75.200 ;
        RECT 116.600 67.800 117.000 68.200 ;
        RECT 119.800 73.800 120.200 74.200 ;
        RECT 119.800 68.800 120.200 69.200 ;
        RECT 113.400 64.800 113.800 65.200 ;
        RECT 155.800 147.800 156.200 148.200 ;
        RECT 147.800 133.800 148.200 134.200 ;
        RECT 143.800 115.800 144.200 116.200 ;
        RECT 134.200 93.800 134.600 94.200 ;
        RECT 129.400 74.800 129.800 75.200 ;
        RECT 107.800 45.800 108.200 46.200 ;
        RECT 97.400 28.800 97.800 29.200 ;
        RECT 83.000 13.800 83.400 14.200 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 84.600 6.800 85.000 7.200 ;
        RECT 84.600 4.800 85.000 5.200 ;
        RECT 117.400 55.800 117.800 56.200 ;
        RECT 120.600 52.800 121.000 53.200 ;
        RECT 113.400 25.800 113.800 26.200 ;
        RECT 140.600 83.800 141.000 84.200 ;
        RECT 147.800 113.800 148.200 114.200 ;
        RECT 149.400 111.800 149.800 112.200 ;
        RECT 168.600 166.800 169.000 167.200 ;
        RECT 178.200 168.800 178.600 169.200 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 178.200 153.800 178.600 154.200 ;
        RECT 169.400 134.800 169.800 135.200 ;
        RECT 172.600 133.800 173.000 134.200 ;
        RECT 139.000 74.800 139.400 75.200 ;
        RECT 135.800 66.800 136.200 67.200 ;
        RECT 143.000 65.800 143.400 66.200 ;
        RECT 128.600 54.800 129.000 55.200 ;
        RECT 142.200 53.800 142.600 54.200 ;
        RECT 131.000 36.800 131.400 37.200 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 127.800 31.800 128.200 32.200 ;
        RECT 107.000 5.800 107.400 6.200 ;
        RECT 104.600 4.800 105.000 5.200 ;
        RECT 129.400 16.800 129.800 17.200 ;
        RECT 127.000 6.800 127.400 7.200 ;
        RECT 148.600 76.800 149.000 77.200 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 158.200 85.800 158.600 86.200 ;
        RECT 179.800 146.800 180.200 147.200 ;
        RECT 179.800 134.800 180.200 135.200 ;
        RECT 172.600 116.800 173.000 117.200 ;
        RECT 171.800 113.800 172.200 114.200 ;
        RECT 171.000 111.800 171.400 112.200 ;
        RECT 171.800 102.800 172.200 103.200 ;
        RECT 175.000 115.800 175.400 116.200 ;
        RECT 179.800 98.800 180.200 99.200 ;
        RECT 168.600 86.800 169.000 87.200 ;
        RECT 158.200 76.800 158.600 77.200 ;
        RECT 161.400 73.800 161.800 74.200 ;
        RECT 167.000 73.800 167.400 74.200 ;
        RECT 172.600 67.800 173.000 68.200 ;
        RECT 163.000 64.800 163.400 65.200 ;
        RECT 140.600 13.800 141.000 14.200 ;
        RECT 140.600 6.800 141.000 7.200 ;
        RECT 143.000 14.800 143.400 15.200 ;
        RECT 151.800 14.800 152.200 15.200 ;
        RECT 144.600 11.800 145.000 12.200 ;
        RECT 160.600 45.800 161.000 46.200 ;
        RECT 163.000 48.800 163.400 49.200 ;
        RECT 159.000 28.800 159.400 29.200 ;
        RECT 203.000 146.800 203.400 147.200 ;
        RECT 214.200 195.800 214.600 196.200 ;
        RECT 213.400 193.800 213.800 194.200 ;
        RECT 232.600 231.800 233.000 232.200 ;
        RECT 236.600 234.800 237.000 235.200 ;
        RECT 245.400 231.800 245.800 232.200 ;
        RECT 222.200 226.800 222.600 227.200 ;
        RECT 230.200 206.800 230.600 207.200 ;
        RECT 241.400 221.800 241.800 222.200 ;
        RECT 241.400 213.800 241.800 214.200 ;
        RECT 217.400 185.800 217.800 186.200 ;
        RECT 207.000 167.800 207.400 168.200 ;
        RECT 215.000 167.800 215.400 168.200 ;
        RECT 206.200 165.800 206.600 166.200 ;
        RECT 244.600 195.800 245.000 196.200 ;
        RECT 228.600 172.800 229.000 173.200 ;
        RECT 206.200 156.800 206.600 157.200 ;
        RECT 239.000 171.800 239.400 172.200 ;
        RECT 235.000 168.800 235.400 169.200 ;
        RECT 206.200 147.800 206.600 148.200 ;
        RECT 220.600 148.800 221.000 149.200 ;
        RECT 228.600 146.800 229.000 147.200 ;
        RECT 228.600 145.800 229.000 146.200 ;
        RECT 227.800 144.800 228.200 145.200 ;
        RECT 201.400 128.800 201.800 129.200 ;
        RECT 195.800 113.800 196.200 114.200 ;
        RECT 217.400 133.800 217.800 134.200 ;
        RECT 218.200 127.800 218.600 128.200 ;
        RECT 226.200 126.800 226.600 127.200 ;
        RECT 219.800 125.800 220.200 126.200 ;
        RECT 212.600 124.800 213.000 125.200 ;
        RECT 199.800 105.800 200.200 106.200 ;
        RECT 203.000 86.800 203.400 87.200 ;
        RECT 202.200 84.800 202.600 85.200 ;
        RECT 201.400 78.800 201.800 79.200 ;
        RECT 202.200 75.800 202.600 76.200 ;
        RECT 220.600 114.800 221.000 115.200 ;
        RECT 219.800 113.800 220.200 114.200 ;
        RECT 234.200 114.800 234.600 115.200 ;
        RECT 213.400 94.800 213.800 95.200 ;
        RECT 203.800 67.800 204.200 68.200 ;
        RECT 187.000 51.800 187.400 52.200 ;
        RECT 181.400 46.800 181.800 47.200 ;
        RECT 159.800 17.800 160.200 18.200 ;
        RECT 187.000 35.800 187.400 36.200 ;
        RECT 187.800 28.800 188.200 29.200 ;
        RECT 186.200 24.800 186.600 25.200 ;
        RECT 186.200 13.800 186.600 14.200 ;
        RECT 180.600 4.800 181.000 5.200 ;
        RECT 209.400 48.800 209.800 49.200 ;
        RECT 200.600 25.800 201.000 26.200 ;
        RECT 217.400 86.800 217.800 87.200 ;
        RECT 219.800 86.800 220.200 87.200 ;
        RECT 227.000 95.800 227.400 96.200 ;
        RECT 243.800 105.800 244.200 106.200 ;
        RECT 231.000 94.800 231.400 95.200 ;
        RECT 219.000 85.800 219.400 86.200 ;
        RECT 215.800 75.800 216.200 76.200 ;
        RECT 212.600 26.800 213.000 27.200 ;
        RECT 217.400 34.800 217.800 35.200 ;
        RECT 229.400 67.800 229.800 68.200 ;
        RECT 247.000 93.800 247.400 94.200 ;
        RECT 248.600 75.800 249.000 76.200 ;
        RECT 244.600 74.800 245.000 75.200 ;
        RECT 233.400 68.800 233.800 69.200 ;
        RECT 225.400 53.800 225.800 54.200 ;
        RECT 215.800 26.800 216.200 27.200 ;
        RECT 207.800 13.800 208.200 14.200 ;
        RECT 221.400 13.800 221.800 14.200 ;
        RECT 231.800 54.800 232.200 55.200 ;
        RECT 240.600 53.800 241.000 54.200 ;
        RECT 237.400 45.800 237.800 46.200 ;
        RECT 240.600 35.800 241.000 36.200 ;
        RECT 243.800 6.800 244.200 7.200 ;
      LAYER metal3 ;
        RECT 74.200 237.800 74.600 238.200 ;
        RECT 85.400 238.100 85.800 238.200 ;
        RECT 112.600 238.100 113.000 238.200 ;
        RECT 85.400 237.800 113.000 238.100 ;
        RECT 55.800 237.100 56.200 237.200 ;
        RECT 57.400 237.100 57.800 237.200 ;
        RECT 55.800 236.800 57.800 237.100 ;
        RECT 63.800 237.100 64.200 237.200 ;
        RECT 74.200 237.100 74.500 237.800 ;
        RECT 63.800 236.800 74.500 237.100 ;
        RECT 104.600 237.100 105.000 237.200 ;
        RECT 111.000 237.100 111.400 237.200 ;
        RECT 104.600 236.800 111.400 237.100 ;
        RECT 191.800 236.800 192.200 237.200 ;
        RECT 7.000 236.100 7.400 236.200 ;
        RECT 8.600 236.100 9.000 236.200 ;
        RECT 7.000 235.800 9.000 236.100 ;
        RECT 29.400 236.100 29.800 236.200 ;
        RECT 31.000 236.100 31.400 236.200 ;
        RECT 29.400 235.800 31.400 236.100 ;
        RECT 36.600 235.800 37.000 236.200 ;
        RECT 55.800 236.100 56.200 236.200 ;
        RECT 59.000 236.100 59.400 236.200 ;
        RECT 110.200 236.100 110.600 236.200 ;
        RECT 55.800 235.800 110.600 236.100 ;
        RECT 112.600 236.100 113.000 236.200 ;
        RECT 121.400 236.100 121.800 236.200 ;
        RECT 112.600 235.800 121.800 236.100 ;
        RECT 128.600 236.100 129.000 236.200 ;
        RECT 130.200 236.100 130.600 236.200 ;
        RECT 128.600 235.800 130.600 236.100 ;
        RECT 132.600 236.100 133.000 236.200 ;
        RECT 134.200 236.100 134.600 236.200 ;
        RECT 132.600 235.800 134.600 236.100 ;
        RECT 184.600 236.100 185.000 236.200 ;
        RECT 191.800 236.100 192.100 236.800 ;
        RECT 184.600 235.800 192.100 236.100 ;
        RECT 199.000 236.100 199.400 236.200 ;
        RECT 208.600 236.100 209.000 236.200 ;
        RECT 199.000 235.800 209.000 236.100 ;
        RECT 209.400 236.100 209.800 236.200 ;
        RECT 221.400 236.100 221.800 236.200 ;
        RECT 238.200 236.100 238.600 236.200 ;
        RECT 209.400 235.800 238.600 236.100 ;
        RECT 9.400 235.100 9.800 235.200 ;
        RECT 16.600 235.100 17.000 235.200 ;
        RECT 9.400 234.800 17.000 235.100 ;
        RECT 19.000 235.100 19.400 235.200 ;
        RECT 28.600 235.100 29.000 235.200 ;
        RECT 19.000 234.800 29.000 235.100 ;
        RECT 31.800 235.100 32.200 235.200 ;
        RECT 36.600 235.100 36.900 235.800 ;
        RECT 31.800 234.800 36.900 235.100 ;
        RECT 51.000 235.100 51.400 235.200 ;
        RECT 55.800 235.100 56.200 235.200 ;
        RECT 51.000 234.800 56.200 235.100 ;
        RECT 59.800 234.800 60.200 235.200 ;
        RECT 71.800 235.100 72.200 235.200 ;
        RECT 75.000 235.100 75.400 235.200 ;
        RECT 127.800 235.100 128.200 235.200 ;
        RECT 71.800 234.800 128.200 235.100 ;
        RECT 147.800 235.100 148.200 235.200 ;
        RECT 151.000 235.100 151.400 235.200 ;
        RECT 147.800 234.800 151.400 235.100 ;
        RECT 156.600 235.100 157.000 235.200 ;
        RECT 157.400 235.100 157.800 235.200 ;
        RECT 159.800 235.100 160.200 235.200 ;
        RECT 156.600 234.800 160.200 235.100 ;
        RECT 170.200 234.800 170.600 235.200 ;
        RECT 183.000 235.100 183.400 235.200 ;
        RECT 191.000 235.100 191.400 235.200 ;
        RECT 183.000 234.800 191.400 235.100 ;
        RECT 193.400 235.100 193.800 235.200 ;
        RECT 204.600 235.100 205.000 235.200 ;
        RECT 193.400 234.800 205.000 235.100 ;
        RECT 207.000 235.100 207.400 235.200 ;
        RECT 209.400 235.100 209.800 235.200 ;
        RECT 207.000 234.800 209.800 235.100 ;
        RECT 223.800 234.800 224.200 235.200 ;
        RECT 227.000 235.100 227.400 235.200 ;
        RECT 231.000 235.100 231.400 235.200 ;
        RECT 227.000 234.800 231.400 235.100 ;
        RECT 233.400 234.800 233.800 235.200 ;
        RECT 235.800 235.100 236.200 235.200 ;
        RECT 236.600 235.100 237.000 235.200 ;
        RECT 235.800 234.800 237.000 235.100 ;
        RECT 241.400 235.100 241.800 235.200 ;
        RECT 246.200 235.100 246.600 235.200 ;
        RECT 249.400 235.100 249.800 235.200 ;
        RECT 241.400 234.800 249.800 235.100 ;
        RECT 2.200 234.100 2.600 234.200 ;
        RECT 4.600 234.100 5.000 234.200 ;
        RECT 5.400 234.100 5.800 234.200 ;
        RECT 27.800 234.100 28.200 234.200 ;
        RECT 2.200 233.800 5.800 234.100 ;
        RECT 22.200 233.800 28.200 234.100 ;
        RECT 45.400 234.100 45.800 234.200 ;
        RECT 55.800 234.100 56.200 234.200 ;
        RECT 58.200 234.100 58.600 234.200 ;
        RECT 45.400 233.800 58.600 234.100 ;
        RECT 59.800 234.100 60.100 234.800 ;
        RECT 75.800 234.100 76.200 234.200 ;
        RECT 76.600 234.100 77.000 234.200 ;
        RECT 91.000 234.100 91.400 234.200 ;
        RECT 59.800 233.800 77.000 234.100 ;
        RECT 83.800 233.800 91.400 234.100 ;
        RECT 97.400 234.100 97.800 234.200 ;
        RECT 110.200 234.100 110.600 234.200 ;
        RECT 119.000 234.100 119.400 234.200 ;
        RECT 97.400 233.800 100.900 234.100 ;
        RECT 110.200 233.800 119.400 234.100 ;
        RECT 119.800 234.100 120.200 234.200 ;
        RECT 128.600 234.100 129.000 234.200 ;
        RECT 119.800 233.800 129.000 234.100 ;
        RECT 147.000 234.100 147.400 234.200 ;
        RECT 156.600 234.100 157.000 234.200 ;
        RECT 147.000 233.800 157.000 234.100 ;
        RECT 159.000 234.100 159.400 234.200 ;
        RECT 167.800 234.100 168.200 234.200 ;
        RECT 159.000 233.800 168.200 234.100 ;
        RECT 170.200 234.100 170.500 234.800 ;
        RECT 223.800 234.200 224.100 234.800 ;
        RECT 188.600 234.100 189.000 234.200 ;
        RECT 199.000 234.100 199.400 234.200 ;
        RECT 214.200 234.100 214.600 234.200 ;
        RECT 170.200 233.800 214.600 234.100 ;
        RECT 220.600 234.100 221.000 234.200 ;
        RECT 221.400 234.100 221.800 234.200 ;
        RECT 220.600 233.800 221.800 234.100 ;
        RECT 223.800 233.800 224.200 234.200 ;
        RECT 230.200 234.100 230.600 234.200 ;
        RECT 233.400 234.100 233.700 234.800 ;
        RECT 230.200 233.800 233.700 234.100 ;
        RECT 246.200 233.800 246.600 234.200 ;
        RECT 22.200 233.200 22.500 233.800 ;
        RECT 83.800 233.200 84.100 233.800 ;
        RECT 100.600 233.200 100.900 233.800 ;
        RECT 246.200 233.200 246.500 233.800 ;
        RECT 6.200 233.100 6.600 233.200 ;
        RECT 17.400 233.100 17.800 233.200 ;
        RECT 22.200 233.100 22.600 233.200 ;
        RECT 6.200 232.800 22.600 233.100 ;
        RECT 28.600 233.100 29.000 233.200 ;
        RECT 34.200 233.100 34.600 233.200 ;
        RECT 36.600 233.100 37.000 233.200 ;
        RECT 28.600 232.800 37.000 233.100 ;
        RECT 53.400 233.100 53.800 233.200 ;
        RECT 63.000 233.100 63.400 233.200 ;
        RECT 53.400 232.800 63.400 233.100 ;
        RECT 83.800 232.800 84.200 233.200 ;
        RECT 100.600 233.100 101.000 233.200 ;
        RECT 117.400 233.100 117.800 233.200 ;
        RECT 124.600 233.100 125.000 233.200 ;
        RECT 100.600 232.800 125.000 233.100 ;
        RECT 178.200 233.100 178.600 233.200 ;
        RECT 199.000 233.100 199.400 233.200 ;
        RECT 178.200 232.800 199.400 233.100 ;
        RECT 210.200 233.100 210.600 233.200 ;
        RECT 225.400 233.100 225.800 233.200 ;
        RECT 210.200 232.800 225.800 233.100 ;
        RECT 246.200 232.800 246.600 233.200 ;
        RECT 33.400 232.100 33.800 232.200 ;
        RECT 42.200 232.100 42.600 232.200 ;
        RECT 64.600 232.100 65.000 232.200 ;
        RECT 33.400 231.800 65.000 232.100 ;
        RECT 70.200 232.100 70.600 232.200 ;
        RECT 91.800 232.100 92.200 232.200 ;
        RECT 70.200 231.800 92.200 232.100 ;
        RECT 97.400 232.100 97.800 232.200 ;
        RECT 119.000 232.100 119.400 232.200 ;
        RECT 97.400 231.800 119.400 232.100 ;
        RECT 130.200 232.100 130.600 232.200 ;
        RECT 205.400 232.100 205.800 232.200 ;
        RECT 220.600 232.100 221.000 232.200 ;
        RECT 130.200 231.800 176.100 232.100 ;
        RECT 205.400 231.800 221.000 232.100 ;
        RECT 232.600 232.100 233.000 232.200 ;
        RECT 233.400 232.100 233.800 232.200 ;
        RECT 232.600 231.800 233.800 232.100 ;
        RECT 239.000 232.100 239.400 232.200 ;
        RECT 240.600 232.100 241.000 232.200 ;
        RECT 239.000 231.800 241.000 232.100 ;
        RECT 244.600 232.100 245.000 232.200 ;
        RECT 245.400 232.100 245.800 232.200 ;
        RECT 244.600 231.800 245.800 232.100 ;
        RECT 75.800 231.100 76.200 231.200 ;
        RECT 76.600 231.100 77.000 231.200 ;
        RECT 75.800 230.800 77.000 231.100 ;
        RECT 80.600 231.100 81.000 231.200 ;
        RECT 85.400 231.100 85.800 231.200 ;
        RECT 80.600 230.800 85.800 231.100 ;
        RECT 108.600 231.100 109.000 231.200 ;
        RECT 123.000 231.100 123.400 231.200 ;
        RECT 108.600 230.800 123.400 231.100 ;
        RECT 126.200 231.100 126.600 231.200 ;
        RECT 144.600 231.100 145.000 231.200 ;
        RECT 126.200 230.800 145.000 231.100 ;
        RECT 148.600 231.100 149.000 231.200 ;
        RECT 175.000 231.100 175.400 231.200 ;
        RECT 148.600 230.800 175.400 231.100 ;
        RECT 175.800 231.100 176.100 231.800 ;
        RECT 181.400 231.100 181.800 231.200 ;
        RECT 175.800 230.800 181.800 231.100 ;
        RECT 191.000 231.100 191.400 231.200 ;
        RECT 195.800 231.100 196.200 231.200 ;
        RECT 191.000 230.800 196.200 231.100 ;
        RECT 82.200 230.100 82.600 230.200 ;
        RECT 97.400 230.100 97.800 230.200 ;
        RECT 82.200 229.800 97.800 230.100 ;
        RECT 134.200 230.100 134.600 230.200 ;
        RECT 135.800 230.100 136.200 230.200 ;
        RECT 134.200 229.800 136.200 230.100 ;
        RECT 136.600 230.100 137.000 230.200 ;
        RECT 147.000 230.100 147.400 230.200 ;
        RECT 150.200 230.100 150.600 230.200 ;
        RECT 136.600 229.800 150.600 230.100 ;
        RECT 161.400 230.100 161.800 230.200 ;
        RECT 187.800 230.100 188.200 230.200 ;
        RECT 161.400 229.800 188.200 230.100 ;
        RECT 22.200 229.100 22.600 229.200 ;
        RECT 31.000 229.100 31.400 229.200 ;
        RECT 33.400 229.100 33.800 229.200 ;
        RECT 22.200 228.800 33.800 229.100 ;
        RECT 42.200 229.100 42.600 229.200 ;
        RECT 51.000 229.100 51.400 229.200 ;
        RECT 55.000 229.100 55.400 229.200 ;
        RECT 42.200 228.800 55.400 229.100 ;
        RECT 87.000 229.100 87.400 229.200 ;
        RECT 109.400 229.100 109.800 229.200 ;
        RECT 115.000 229.100 115.400 229.200 ;
        RECT 120.600 229.100 121.000 229.200 ;
        RECT 131.800 229.100 132.200 229.200 ;
        RECT 138.200 229.100 138.600 229.200 ;
        RECT 87.000 228.800 138.600 229.100 ;
        RECT 153.400 229.100 153.800 229.200 ;
        RECT 182.200 229.100 182.600 229.200 ;
        RECT 186.200 229.100 186.600 229.200 ;
        RECT 153.400 228.800 186.600 229.100 ;
        RECT 190.200 229.100 190.600 229.200 ;
        RECT 190.200 228.800 204.100 229.100 ;
        RECT 203.800 228.200 204.100 228.800 ;
        RECT 67.800 228.100 68.200 228.200 ;
        RECT 75.800 228.100 76.200 228.200 ;
        RECT 85.400 228.100 85.800 228.200 ;
        RECT 67.800 227.800 85.800 228.100 ;
        RECT 90.200 228.100 90.600 228.200 ;
        RECT 91.000 228.100 91.400 228.200 ;
        RECT 90.200 227.800 91.400 228.100 ;
        RECT 94.200 228.100 94.600 228.200 ;
        RECT 97.400 228.100 97.800 228.200 ;
        RECT 110.200 228.100 110.600 228.200 ;
        RECT 94.200 227.800 110.600 228.100 ;
        RECT 127.000 228.100 127.400 228.200 ;
        RECT 128.600 228.100 129.000 228.200 ;
        RECT 141.400 228.100 141.800 228.200 ;
        RECT 127.000 227.800 141.800 228.100 ;
        RECT 142.200 228.100 142.600 228.200 ;
        RECT 162.200 228.100 162.600 228.200 ;
        RECT 142.200 227.800 162.600 228.100 ;
        RECT 171.800 228.100 172.200 228.200 ;
        RECT 190.200 228.100 190.600 228.200 ;
        RECT 201.400 228.100 201.800 228.200 ;
        RECT 171.800 227.800 201.800 228.100 ;
        RECT 203.800 228.100 204.200 228.200 ;
        RECT 219.000 228.100 219.400 228.200 ;
        RECT 203.800 227.800 219.400 228.100 ;
        RECT 221.400 228.100 221.800 228.200 ;
        RECT 235.800 228.100 236.200 228.200 ;
        RECT 221.400 227.800 236.200 228.100 ;
        RECT 11.000 227.100 11.400 227.200 ;
        RECT 35.800 227.100 36.200 227.200 ;
        RECT 11.000 226.800 36.200 227.100 ;
        RECT 56.600 227.100 57.000 227.200 ;
        RECT 62.200 227.100 62.600 227.200 ;
        RECT 56.600 226.800 62.600 227.100 ;
        RECT 79.000 226.800 79.400 227.200 ;
        RECT 91.000 227.100 91.400 227.200 ;
        RECT 100.600 227.100 101.000 227.200 ;
        RECT 91.000 226.800 101.000 227.100 ;
        RECT 103.000 226.800 103.400 227.200 ;
        RECT 105.400 227.100 105.800 227.200 ;
        RECT 107.800 227.100 108.200 227.200 ;
        RECT 122.200 227.100 122.600 227.200 ;
        RECT 147.800 227.100 148.200 227.200 ;
        RECT 105.400 226.800 108.200 227.100 ;
        RECT 119.800 226.800 148.200 227.100 ;
        RECT 154.200 227.100 154.600 227.200 ;
        RECT 155.000 227.100 155.400 227.200 ;
        RECT 154.200 226.800 155.400 227.100 ;
        RECT 183.000 226.800 183.400 227.200 ;
        RECT 192.600 226.800 193.000 227.200 ;
        RECT 195.000 227.100 195.400 227.200 ;
        RECT 222.200 227.100 222.600 227.200 ;
        RECT 195.000 226.800 222.600 227.100 ;
        RECT 223.800 227.100 224.200 227.200 ;
        RECT 230.200 227.100 230.600 227.200 ;
        RECT 223.800 226.800 230.600 227.100 ;
        RECT 243.800 226.800 244.200 227.200 ;
        RECT 19.000 226.100 19.400 226.200 ;
        RECT 20.600 226.100 21.000 226.200 ;
        RECT 39.000 226.100 39.400 226.200 ;
        RECT 19.000 225.800 21.000 226.100 ;
        RECT 35.000 225.800 39.400 226.100 ;
        RECT 40.600 226.100 41.000 226.200 ;
        RECT 40.600 225.800 45.700 226.100 ;
        RECT 35.000 225.200 35.300 225.800 ;
        RECT 45.400 225.200 45.700 225.800 ;
        RECT 59.800 225.800 60.200 226.200 ;
        RECT 63.000 226.100 63.400 226.200 ;
        RECT 74.200 226.100 74.600 226.200 ;
        RECT 79.000 226.100 79.300 226.800 ;
        RECT 63.000 225.800 79.300 226.100 ;
        RECT 81.400 226.100 81.800 226.200 ;
        RECT 86.200 226.100 86.600 226.200 ;
        RECT 81.400 225.800 86.600 226.100 ;
        RECT 87.800 225.800 88.200 226.200 ;
        RECT 95.800 226.100 96.200 226.200 ;
        RECT 101.400 226.100 101.800 226.200 ;
        RECT 95.800 225.800 101.800 226.100 ;
        RECT 103.000 226.100 103.300 226.800 ;
        RECT 119.800 226.200 120.100 226.800 ;
        RECT 108.600 226.100 109.000 226.200 ;
        RECT 103.000 225.800 109.000 226.100 ;
        RECT 118.200 226.100 118.600 226.200 ;
        RECT 119.800 226.100 120.200 226.200 ;
        RECT 118.200 225.800 120.200 226.100 ;
        RECT 124.600 226.100 125.000 226.200 ;
        RECT 138.200 226.100 138.600 226.200 ;
        RECT 143.000 226.100 143.400 226.200 ;
        RECT 144.600 226.100 145.000 226.200 ;
        RECT 124.600 225.800 145.000 226.100 ;
        RECT 146.200 226.100 146.600 226.200 ;
        RECT 164.600 226.100 165.000 226.200 ;
        RECT 183.000 226.100 183.300 226.800 ;
        RECT 146.200 225.800 183.300 226.100 ;
        RECT 189.400 226.100 189.800 226.200 ;
        RECT 192.600 226.100 192.900 226.800 ;
        RECT 189.400 225.800 192.900 226.100 ;
        RECT 196.600 226.100 197.000 226.200 ;
        RECT 197.400 226.100 197.800 226.200 ;
        RECT 199.800 226.100 200.200 226.200 ;
        RECT 196.600 225.800 200.200 226.100 ;
        RECT 215.000 226.100 215.400 226.200 ;
        RECT 215.800 226.100 216.200 226.200 ;
        RECT 215.000 225.800 216.200 226.100 ;
        RECT 226.200 225.800 226.600 226.200 ;
        RECT 228.600 226.100 229.000 226.200 ;
        RECT 235.800 226.100 236.200 226.200 ;
        RECT 228.600 225.800 236.200 226.100 ;
        RECT 239.000 226.100 239.400 226.200 ;
        RECT 243.800 226.100 244.100 226.800 ;
        RECT 239.000 225.800 244.100 226.100 ;
        RECT 247.000 225.800 247.400 226.200 ;
        RECT 59.800 225.200 60.100 225.800 ;
        RECT 19.800 225.100 20.200 225.200 ;
        RECT 25.400 225.100 25.800 225.200 ;
        RECT 19.800 224.800 25.800 225.100 ;
        RECT 35.000 224.800 35.400 225.200 ;
        RECT 38.200 225.100 38.600 225.200 ;
        RECT 41.400 225.100 41.800 225.200 ;
        RECT 43.800 225.100 44.200 225.200 ;
        RECT 38.200 224.800 44.200 225.100 ;
        RECT 45.400 224.800 45.800 225.200 ;
        RECT 59.800 224.800 60.200 225.200 ;
        RECT 86.200 225.100 86.600 225.200 ;
        RECT 87.800 225.100 88.100 225.800 ;
        RECT 226.200 225.200 226.500 225.800 ;
        RECT 247.000 225.200 247.300 225.800 ;
        RECT 86.200 224.800 88.100 225.100 ;
        RECT 107.800 225.100 108.200 225.200 ;
        RECT 110.200 225.100 110.600 225.200 ;
        RECT 111.000 225.100 111.400 225.200 ;
        RECT 132.600 225.100 133.000 225.200 ;
        RECT 107.800 224.800 133.000 225.100 ;
        RECT 135.000 225.100 135.400 225.200 ;
        RECT 139.800 225.100 140.200 225.200 ;
        RECT 135.000 224.800 140.200 225.100 ;
        RECT 140.600 225.100 141.000 225.200 ;
        RECT 158.200 225.100 158.600 225.200 ;
        RECT 175.800 225.100 176.200 225.200 ;
        RECT 140.600 224.800 176.200 225.100 ;
        RECT 182.200 224.800 182.600 225.200 ;
        RECT 183.000 225.100 183.400 225.200 ;
        RECT 204.600 225.100 205.000 225.200 ;
        RECT 183.000 224.800 205.000 225.100 ;
        RECT 214.200 225.100 214.600 225.200 ;
        RECT 215.800 225.100 216.200 225.200 ;
        RECT 214.200 224.800 216.200 225.100 ;
        RECT 226.200 225.100 226.600 225.200 ;
        RECT 227.800 225.100 228.200 225.200 ;
        RECT 228.600 225.100 229.000 225.200 ;
        RECT 226.200 224.800 229.000 225.100 ;
        RECT 247.000 224.800 247.400 225.200 ;
        RECT 8.600 224.100 9.000 224.200 ;
        RECT 16.600 224.100 17.000 224.200 ;
        RECT 28.600 224.100 29.000 224.200 ;
        RECT 37.400 224.100 37.800 224.200 ;
        RECT 8.600 223.800 37.800 224.100 ;
        RECT 59.000 224.100 59.400 224.200 ;
        RECT 105.400 224.100 105.800 224.200 ;
        RECT 59.000 223.800 105.800 224.100 ;
        RECT 107.000 224.100 107.400 224.200 ;
        RECT 112.600 224.100 113.000 224.200 ;
        RECT 107.000 223.800 113.000 224.100 ;
        RECT 116.600 224.100 117.000 224.200 ;
        RECT 136.600 224.100 137.000 224.200 ;
        RECT 140.600 224.100 140.900 224.800 ;
        RECT 182.200 224.200 182.500 224.800 ;
        RECT 116.600 223.800 140.900 224.100 ;
        RECT 148.600 224.100 149.000 224.200 ;
        RECT 160.600 224.100 161.000 224.200 ;
        RECT 163.000 224.100 163.400 224.200 ;
        RECT 148.600 223.800 163.400 224.100 ;
        RECT 182.200 223.800 182.600 224.200 ;
        RECT 185.400 224.100 185.800 224.200 ;
        RECT 197.400 224.100 197.800 224.200 ;
        RECT 185.400 223.800 197.800 224.100 ;
        RECT 199.800 224.100 200.200 224.200 ;
        RECT 244.600 224.100 245.000 224.200 ;
        RECT 199.800 223.800 245.000 224.100 ;
        RECT 13.400 223.100 13.800 223.200 ;
        RECT 87.000 223.100 87.400 223.200 ;
        RECT 13.400 222.800 87.400 223.100 ;
        RECT 90.200 223.100 90.600 223.200 ;
        RECT 120.600 223.100 121.000 223.200 ;
        RECT 90.200 222.800 121.000 223.100 ;
        RECT 127.800 223.100 128.200 223.200 ;
        RECT 134.200 223.100 134.600 223.200 ;
        RECT 127.800 222.800 134.600 223.100 ;
        RECT 155.800 223.100 156.200 223.200 ;
        RECT 183.000 223.100 183.400 223.200 ;
        RECT 155.800 222.800 183.400 223.100 ;
        RECT 224.600 223.100 225.000 223.200 ;
        RECT 235.000 223.100 235.400 223.200 ;
        RECT 224.600 222.800 235.400 223.100 ;
        RECT 1.400 222.100 1.800 222.200 ;
        RECT 25.400 222.100 25.800 222.200 ;
        RECT 1.400 221.800 25.800 222.100 ;
        RECT 32.600 222.100 33.000 222.200 ;
        RECT 57.400 222.100 57.800 222.200 ;
        RECT 32.600 221.800 57.800 222.100 ;
        RECT 63.800 222.100 64.200 222.200 ;
        RECT 89.400 222.100 89.800 222.200 ;
        RECT 63.800 221.800 89.800 222.100 ;
        RECT 115.000 222.100 115.400 222.200 ;
        RECT 115.800 222.100 116.200 222.200 ;
        RECT 115.000 221.800 116.200 222.100 ;
        RECT 119.000 222.100 119.400 222.200 ;
        RECT 121.400 222.100 121.800 222.200 ;
        RECT 119.000 221.800 121.800 222.100 ;
        RECT 156.600 222.100 157.000 222.200 ;
        RECT 159.800 222.100 160.200 222.200 ;
        RECT 178.200 222.100 178.600 222.200 ;
        RECT 195.800 222.100 196.200 222.200 ;
        RECT 199.000 222.100 199.400 222.200 ;
        RECT 156.600 221.800 199.400 222.100 ;
        RECT 209.400 222.100 209.800 222.200 ;
        RECT 214.200 222.100 214.600 222.200 ;
        RECT 216.600 222.100 217.000 222.200 ;
        RECT 209.400 221.800 217.000 222.100 ;
        RECT 225.400 222.100 225.800 222.200 ;
        RECT 235.000 222.100 235.400 222.200 ;
        RECT 225.400 221.800 235.400 222.100 ;
        RECT 241.400 222.100 241.800 222.200 ;
        RECT 242.200 222.100 242.600 222.200 ;
        RECT 241.400 221.800 242.600 222.100 ;
        RECT 7.000 221.100 7.400 221.200 ;
        RECT 19.000 221.100 19.400 221.200 ;
        RECT 7.000 220.800 19.400 221.100 ;
        RECT 67.000 221.100 67.400 221.200 ;
        RECT 68.600 221.100 69.000 221.200 ;
        RECT 67.000 220.800 69.000 221.100 ;
        RECT 103.800 221.100 104.200 221.200 ;
        RECT 116.600 221.100 117.000 221.200 ;
        RECT 103.800 220.800 117.000 221.100 ;
        RECT 213.400 221.100 213.800 221.200 ;
        RECT 239.800 221.100 240.200 221.200 ;
        RECT 213.400 220.800 240.200 221.100 ;
        RECT 61.400 220.100 61.800 220.200 ;
        RECT 63.800 220.100 64.200 220.200 ;
        RECT 61.400 219.800 64.200 220.100 ;
        RECT 66.200 220.100 66.600 220.200 ;
        RECT 69.400 220.100 69.800 220.200 ;
        RECT 66.200 219.800 69.800 220.100 ;
        RECT 87.000 220.100 87.400 220.200 ;
        RECT 91.000 220.100 91.400 220.200 ;
        RECT 106.200 220.100 106.600 220.200 ;
        RECT 87.000 219.800 106.600 220.100 ;
        RECT 215.800 220.100 216.200 220.200 ;
        RECT 223.800 220.100 224.200 220.200 ;
        RECT 215.800 219.800 224.200 220.100 ;
        RECT 1.400 219.100 1.800 219.200 ;
        RECT 15.000 219.100 15.400 219.200 ;
        RECT 96.600 219.100 97.000 219.200 ;
        RECT 1.400 218.800 97.000 219.100 ;
        RECT 159.800 219.100 160.200 219.200 ;
        RECT 211.800 219.100 212.200 219.200 ;
        RECT 234.200 219.100 234.600 219.200 ;
        RECT 159.800 218.800 234.600 219.100 ;
        RECT 245.400 219.100 245.800 219.200 ;
        RECT 248.600 219.100 249.000 219.200 ;
        RECT 245.400 218.800 249.000 219.100 ;
        RECT 70.200 217.800 70.600 218.200 ;
        RECT 99.800 218.100 100.200 218.200 ;
        RECT 106.200 218.100 106.600 218.200 ;
        RECT 99.800 217.800 106.600 218.100 ;
        RECT 124.600 218.100 125.000 218.200 ;
        RECT 136.600 218.100 137.000 218.200 ;
        RECT 124.600 217.800 137.000 218.100 ;
        RECT 148.600 218.100 149.000 218.200 ;
        RECT 182.200 218.100 182.600 218.200 ;
        RECT 148.600 217.800 182.600 218.100 ;
        RECT 190.200 218.100 190.600 218.200 ;
        RECT 191.800 218.100 192.200 218.200 ;
        RECT 190.200 217.800 192.200 218.100 ;
        RECT 197.400 218.100 197.800 218.200 ;
        RECT 210.200 218.100 210.600 218.200 ;
        RECT 197.400 217.800 210.600 218.100 ;
        RECT 8.600 217.100 9.000 217.200 ;
        RECT 11.000 217.100 11.400 217.200 ;
        RECT 14.200 217.100 14.600 217.200 ;
        RECT 16.600 217.100 17.000 217.200 ;
        RECT 8.600 216.800 17.000 217.100 ;
        RECT 34.200 217.100 34.600 217.200 ;
        RECT 35.000 217.100 35.400 217.200 ;
        RECT 34.200 216.800 35.400 217.100 ;
        RECT 65.400 217.100 65.800 217.200 ;
        RECT 70.200 217.100 70.500 217.800 ;
        RECT 65.400 216.800 70.500 217.100 ;
        RECT 91.800 216.800 92.200 217.200 ;
        RECT 100.600 217.100 101.000 217.200 ;
        RECT 163.000 217.100 163.400 217.200 ;
        RECT 165.400 217.100 165.800 217.200 ;
        RECT 212.600 217.100 213.000 217.200 ;
        RECT 217.400 217.100 217.800 217.200 ;
        RECT 100.600 216.800 217.800 217.100 ;
        RECT 221.400 216.800 221.800 217.200 ;
        RECT 7.000 216.100 7.400 216.200 ;
        RECT 11.800 216.100 12.200 216.200 ;
        RECT 7.000 215.800 12.200 216.100 ;
        RECT 28.600 216.100 29.000 216.200 ;
        RECT 31.800 216.100 32.200 216.200 ;
        RECT 35.800 216.100 36.200 216.200 ;
        RECT 28.600 215.800 36.200 216.100 ;
        RECT 43.800 216.100 44.200 216.200 ;
        RECT 62.200 216.100 62.600 216.200 ;
        RECT 43.800 215.800 62.600 216.100 ;
        RECT 64.600 216.100 65.000 216.200 ;
        RECT 69.400 216.100 69.800 216.200 ;
        RECT 64.600 215.800 69.800 216.100 ;
        RECT 84.600 216.100 85.000 216.200 ;
        RECT 91.800 216.100 92.100 216.800 ;
        RECT 84.600 215.800 92.100 216.100 ;
        RECT 94.200 216.100 94.600 216.200 ;
        RECT 157.400 216.100 157.800 216.200 ;
        RECT 159.000 216.100 159.400 216.200 ;
        RECT 94.200 215.800 159.400 216.100 ;
        RECT 205.400 216.100 205.800 216.200 ;
        RECT 221.400 216.100 221.700 216.800 ;
        RECT 225.400 216.100 225.800 216.200 ;
        RECT 205.400 215.800 208.100 216.100 ;
        RECT 221.400 215.800 225.800 216.100 ;
        RECT 236.600 216.100 237.000 216.200 ;
        RECT 237.400 216.100 237.800 216.200 ;
        RECT 239.800 216.100 240.200 216.200 ;
        RECT 245.400 216.100 245.800 216.200 ;
        RECT 236.600 215.800 245.800 216.100 ;
        RECT 207.800 215.200 208.100 215.800 ;
        RECT 10.200 215.100 10.600 215.200 ;
        RECT 11.000 215.100 11.400 215.200 ;
        RECT 13.400 215.100 13.800 215.200 ;
        RECT 10.200 214.800 13.800 215.100 ;
        RECT 20.600 215.100 21.000 215.200 ;
        RECT 70.200 215.100 70.600 215.200 ;
        RECT 20.600 214.800 70.600 215.100 ;
        RECT 72.600 215.100 73.000 215.200 ;
        RECT 76.600 215.100 77.000 215.200 ;
        RECT 90.200 215.100 90.600 215.200 ;
        RECT 91.000 215.100 91.400 215.200 ;
        RECT 72.600 214.800 91.400 215.100 ;
        RECT 92.600 215.100 93.000 215.200 ;
        RECT 95.800 215.100 96.200 215.200 ;
        RECT 100.600 215.100 101.000 215.200 ;
        RECT 92.600 214.800 101.000 215.100 ;
        RECT 105.400 214.800 105.800 215.200 ;
        RECT 122.200 215.100 122.600 215.200 ;
        RECT 125.400 215.100 125.800 215.200 ;
        RECT 122.200 214.800 125.800 215.100 ;
        RECT 130.200 215.100 130.600 215.200 ;
        RECT 131.000 215.100 131.400 215.200 ;
        RECT 133.400 215.100 133.800 215.200 ;
        RECT 130.200 214.800 133.800 215.100 ;
        RECT 147.000 215.100 147.400 215.200 ;
        RECT 150.200 215.100 150.600 215.200 ;
        RECT 147.000 214.800 150.600 215.100 ;
        RECT 153.400 215.100 153.800 215.200 ;
        RECT 166.200 215.100 166.600 215.200 ;
        RECT 168.600 215.100 169.000 215.200 ;
        RECT 153.400 214.800 169.000 215.100 ;
        RECT 180.600 215.100 181.000 215.200 ;
        RECT 185.400 215.100 185.800 215.200 ;
        RECT 199.800 215.100 200.200 215.200 ;
        RECT 180.600 214.800 200.200 215.100 ;
        RECT 207.800 214.800 208.200 215.200 ;
        RECT 217.400 215.100 217.800 215.200 ;
        RECT 220.600 215.100 221.000 215.200 ;
        RECT 217.400 214.800 221.000 215.100 ;
        RECT 235.000 215.100 235.400 215.200 ;
        RECT 240.600 215.100 241.000 215.200 ;
        RECT 235.000 214.800 241.000 215.100 ;
        RECT 30.200 214.100 30.600 214.200 ;
        RECT 34.200 214.100 34.600 214.200 ;
        RECT 30.200 213.800 34.600 214.100 ;
        RECT 40.600 214.100 41.000 214.200 ;
        RECT 71.800 214.100 72.200 214.200 ;
        RECT 77.400 214.100 77.800 214.200 ;
        RECT 40.600 213.800 77.800 214.100 ;
        RECT 91.000 214.100 91.400 214.200 ;
        RECT 105.400 214.100 105.700 214.800 ;
        RECT 91.000 213.800 105.700 214.100 ;
        RECT 106.200 214.100 106.600 214.200 ;
        RECT 108.600 214.100 109.000 214.200 ;
        RECT 106.200 213.800 109.000 214.100 ;
        RECT 119.000 214.100 119.400 214.200 ;
        RECT 131.000 214.100 131.400 214.200 ;
        RECT 119.000 213.800 131.400 214.100 ;
        RECT 132.600 214.100 133.000 214.200 ;
        RECT 138.200 214.100 138.600 214.200 ;
        RECT 132.600 213.800 138.600 214.100 ;
        RECT 143.800 214.100 144.200 214.200 ;
        RECT 145.400 214.100 145.800 214.200 ;
        RECT 143.800 213.800 145.800 214.100 ;
        RECT 164.600 214.100 165.000 214.200 ;
        RECT 170.200 214.100 170.600 214.200 ;
        RECT 164.600 213.800 170.600 214.100 ;
        RECT 181.400 214.100 181.800 214.200 ;
        RECT 187.800 214.100 188.200 214.200 ;
        RECT 181.400 213.800 188.200 214.100 ;
        RECT 204.600 214.100 205.000 214.200 ;
        RECT 215.800 214.100 216.200 214.200 ;
        RECT 221.400 214.100 221.800 214.200 ;
        RECT 204.600 213.800 221.800 214.100 ;
        RECT 241.400 214.100 241.800 214.200 ;
        RECT 247.000 214.100 247.400 214.200 ;
        RECT 241.400 213.800 247.400 214.100 ;
        RECT 21.400 213.100 21.800 213.200 ;
        RECT 43.800 213.100 44.200 213.200 ;
        RECT 52.600 213.100 53.000 213.200 ;
        RECT 21.400 212.800 53.000 213.100 ;
        RECT 74.200 213.100 74.600 213.200 ;
        RECT 75.000 213.100 75.400 213.200 ;
        RECT 74.200 212.800 75.400 213.100 ;
        RECT 107.800 213.100 108.200 213.200 ;
        RECT 115.000 213.100 115.400 213.200 ;
        RECT 107.800 212.800 115.400 213.100 ;
        RECT 107.800 212.200 108.100 212.800 ;
        RECT 20.600 212.100 21.000 212.200 ;
        RECT 23.800 212.100 24.200 212.200 ;
        RECT 20.600 211.800 24.200 212.100 ;
        RECT 32.600 212.100 33.000 212.200 ;
        RECT 41.400 212.100 41.800 212.200 ;
        RECT 32.600 211.800 41.800 212.100 ;
        RECT 74.200 212.100 74.600 212.200 ;
        RECT 75.800 212.100 76.200 212.200 ;
        RECT 74.200 211.800 76.200 212.100 ;
        RECT 91.000 212.100 91.400 212.200 ;
        RECT 94.200 212.100 94.600 212.200 ;
        RECT 91.000 211.800 94.600 212.100 ;
        RECT 96.600 212.100 97.000 212.200 ;
        RECT 99.000 212.100 99.400 212.200 ;
        RECT 96.600 211.800 99.400 212.100 ;
        RECT 107.800 211.800 108.200 212.200 ;
        RECT 124.600 212.100 125.000 212.200 ;
        RECT 135.000 212.100 135.400 212.200 ;
        RECT 143.800 212.100 144.200 212.200 ;
        RECT 124.600 211.800 144.200 212.100 ;
        RECT 145.400 212.100 145.800 212.200 ;
        RECT 146.200 212.100 146.600 212.200 ;
        RECT 145.400 211.800 146.600 212.100 ;
        RECT 167.000 212.100 167.400 212.200 ;
        RECT 219.000 212.100 219.400 212.200 ;
        RECT 231.000 212.100 231.400 212.200 ;
        RECT 167.000 211.800 176.900 212.100 ;
        RECT 219.000 211.800 231.400 212.100 ;
        RECT 240.600 212.100 241.000 212.200 ;
        RECT 244.600 212.100 245.000 212.200 ;
        RECT 240.600 211.800 245.000 212.100 ;
        RECT 176.600 211.200 176.900 211.800 ;
        RECT 10.200 211.100 10.600 211.200 ;
        RECT 15.800 211.100 16.200 211.200 ;
        RECT 40.600 211.100 41.000 211.200 ;
        RECT 10.200 210.800 41.000 211.100 ;
        RECT 54.200 211.100 54.600 211.200 ;
        RECT 66.200 211.100 66.600 211.200 ;
        RECT 54.200 210.800 66.600 211.100 ;
        RECT 72.600 211.100 73.000 211.200 ;
        RECT 76.600 211.100 77.000 211.200 ;
        RECT 72.600 210.800 77.000 211.100 ;
        RECT 79.000 211.100 79.400 211.200 ;
        RECT 94.200 211.100 94.600 211.200 ;
        RECT 79.000 210.800 94.600 211.100 ;
        RECT 113.400 211.100 113.800 211.200 ;
        RECT 117.400 211.100 117.800 211.200 ;
        RECT 113.400 210.800 117.800 211.100 ;
        RECT 131.000 211.100 131.400 211.200 ;
        RECT 143.000 211.100 143.400 211.200 ;
        RECT 148.600 211.100 149.000 211.200 ;
        RECT 156.600 211.100 157.000 211.200 ;
        RECT 162.200 211.100 162.600 211.200 ;
        RECT 165.400 211.100 165.800 211.200 ;
        RECT 131.000 210.800 165.800 211.100 ;
        RECT 176.600 210.800 177.000 211.200 ;
        RECT 24.600 210.100 25.000 210.200 ;
        RECT 58.200 210.100 58.600 210.200 ;
        RECT 24.600 209.800 58.600 210.100 ;
        RECT 103.000 210.100 103.400 210.200 ;
        RECT 107.800 210.100 108.200 210.200 ;
        RECT 103.000 209.800 108.200 210.100 ;
        RECT 135.000 210.100 135.400 210.200 ;
        RECT 141.400 210.100 141.800 210.200 ;
        RECT 135.000 209.800 141.800 210.100 ;
        RECT 160.600 210.100 161.000 210.200 ;
        RECT 191.000 210.100 191.400 210.200 ;
        RECT 219.800 210.100 220.200 210.200 ;
        RECT 226.200 210.100 226.600 210.200 ;
        RECT 235.800 210.100 236.200 210.200 ;
        RECT 160.600 209.800 200.900 210.100 ;
        RECT 219.800 209.800 236.200 210.100 ;
        RECT 249.400 209.800 249.800 210.200 ;
        RECT 1.400 209.100 1.800 209.200 ;
        RECT 27.800 209.100 28.200 209.200 ;
        RECT 54.200 209.100 54.600 209.200 ;
        RECT 1.400 208.800 15.300 209.100 ;
        RECT 27.800 208.800 54.600 209.100 ;
        RECT 57.400 209.100 57.800 209.200 ;
        RECT 73.400 209.100 73.800 209.200 ;
        RECT 123.000 209.100 123.400 209.200 ;
        RECT 169.400 209.100 169.800 209.200 ;
        RECT 57.400 208.800 169.800 209.100 ;
        RECT 191.000 209.100 191.400 209.200 ;
        RECT 193.400 209.100 193.800 209.200 ;
        RECT 195.000 209.100 195.400 209.200 ;
        RECT 195.800 209.100 196.200 209.200 ;
        RECT 191.000 208.800 193.800 209.100 ;
        RECT 194.200 208.800 196.200 209.100 ;
        RECT 200.600 209.100 200.900 209.800 ;
        RECT 249.400 209.200 249.700 209.800 ;
        RECT 225.400 209.100 225.800 209.200 ;
        RECT 200.600 208.800 225.800 209.100 ;
        RECT 228.600 209.100 229.000 209.200 ;
        RECT 240.600 209.100 241.000 209.200 ;
        RECT 228.600 208.800 241.000 209.100 ;
        RECT 246.200 208.800 246.600 209.200 ;
        RECT 249.400 208.800 249.800 209.200 ;
        RECT 15.000 208.200 15.300 208.800 ;
        RECT 8.600 207.800 9.000 208.200 ;
        RECT 15.000 207.800 15.400 208.200 ;
        RECT 35.800 208.100 36.200 208.200 ;
        RECT 27.800 207.800 36.200 208.100 ;
        RECT 65.400 208.100 65.800 208.200 ;
        RECT 75.000 208.100 75.400 208.200 ;
        RECT 65.400 207.800 75.400 208.100 ;
        RECT 77.400 208.100 77.800 208.200 ;
        RECT 88.600 208.100 89.000 208.200 ;
        RECT 90.200 208.100 90.600 208.200 ;
        RECT 77.400 207.800 90.600 208.100 ;
        RECT 97.400 208.100 97.800 208.200 ;
        RECT 100.600 208.100 101.000 208.200 ;
        RECT 103.000 208.100 103.400 208.200 ;
        RECT 97.400 207.800 103.400 208.100 ;
        RECT 115.800 208.100 116.200 208.200 ;
        RECT 123.800 208.100 124.200 208.200 ;
        RECT 115.800 207.800 124.200 208.100 ;
        RECT 136.600 207.800 137.000 208.200 ;
        RECT 144.600 208.100 145.000 208.200 ;
        RECT 145.400 208.100 145.800 208.200 ;
        RECT 144.600 207.800 145.800 208.100 ;
        RECT 159.800 208.100 160.200 208.200 ;
        RECT 161.400 208.100 161.800 208.200 ;
        RECT 159.800 207.800 161.800 208.100 ;
        RECT 170.200 208.100 170.600 208.200 ;
        RECT 176.600 208.100 177.000 208.200 ;
        RECT 179.800 208.100 180.200 208.200 ;
        RECT 170.200 207.800 180.200 208.100 ;
        RECT 188.600 208.100 189.000 208.200 ;
        RECT 195.000 208.100 195.400 208.200 ;
        RECT 202.200 208.100 202.600 208.200 ;
        RECT 242.200 208.100 242.600 208.200 ;
        RECT 188.600 207.800 202.600 208.100 ;
        RECT 203.000 207.800 242.600 208.100 ;
        RECT 246.200 208.100 246.500 208.800 ;
        RECT 248.600 208.100 249.000 208.200 ;
        RECT 246.200 207.800 249.000 208.100 ;
        RECT 8.600 207.200 8.900 207.800 ;
        RECT 8.600 206.800 9.000 207.200 ;
        RECT 15.000 207.100 15.300 207.800 ;
        RECT 27.800 207.200 28.100 207.800 ;
        RECT 22.200 207.100 22.600 207.200 ;
        RECT 15.000 206.800 22.600 207.100 ;
        RECT 27.800 206.800 28.200 207.200 ;
        RECT 29.400 207.100 29.800 207.200 ;
        RECT 62.200 207.100 62.600 207.200 ;
        RECT 123.800 207.100 124.200 207.200 ;
        RECT 29.400 206.800 124.200 207.100 ;
        RECT 136.600 207.100 136.900 207.800 ;
        RECT 149.400 207.100 149.800 207.200 ;
        RECT 136.600 206.800 149.800 207.100 ;
        RECT 154.200 207.100 154.600 207.200 ;
        RECT 159.000 207.100 159.400 207.200 ;
        RECT 154.200 206.800 159.400 207.100 ;
        RECT 163.800 207.100 164.200 207.200 ;
        RECT 167.000 207.100 167.400 207.200 ;
        RECT 163.800 206.800 167.400 207.100 ;
        RECT 167.800 207.100 168.200 207.200 ;
        RECT 173.400 207.100 173.800 207.200 ;
        RECT 167.800 206.800 173.800 207.100 ;
        RECT 187.000 207.100 187.400 207.200 ;
        RECT 190.200 207.100 190.600 207.200 ;
        RECT 187.000 206.800 190.600 207.100 ;
        RECT 191.800 207.100 192.200 207.200 ;
        RECT 203.000 207.100 203.300 207.800 ;
        RECT 223.800 207.100 224.200 207.200 ;
        RECT 230.200 207.100 230.600 207.200 ;
        RECT 232.600 207.100 233.000 207.200 ;
        RECT 191.800 206.800 203.300 207.100 ;
        RECT 211.800 206.800 213.700 207.100 ;
        RECT 223.800 206.800 233.000 207.100 ;
        RECT 6.200 206.100 6.600 206.200 ;
        RECT 12.600 206.100 13.000 206.200 ;
        RECT 6.200 205.800 13.000 206.100 ;
        RECT 17.400 206.100 17.800 206.200 ;
        RECT 19.000 206.100 19.400 206.200 ;
        RECT 17.400 205.800 19.400 206.100 ;
        RECT 27.800 206.100 28.200 206.200 ;
        RECT 29.400 206.100 29.700 206.800 ;
        RECT 211.800 206.200 212.100 206.800 ;
        RECT 213.400 206.200 213.700 206.800 ;
        RECT 27.800 205.800 29.700 206.100 ;
        RECT 37.400 206.100 37.800 206.200 ;
        RECT 49.400 206.100 49.800 206.200 ;
        RECT 51.000 206.100 51.400 206.200 ;
        RECT 37.400 205.800 40.900 206.100 ;
        RECT 49.400 205.800 51.400 206.100 ;
        RECT 59.000 206.100 59.400 206.200 ;
        RECT 60.600 206.100 61.000 206.200 ;
        RECT 63.000 206.100 63.400 206.200 ;
        RECT 59.000 205.800 63.400 206.100 ;
        RECT 67.000 206.100 67.400 206.200 ;
        RECT 69.400 206.100 69.800 206.200 ;
        RECT 73.400 206.100 73.800 206.200 ;
        RECT 67.000 205.800 69.800 206.100 ;
        RECT 71.800 205.800 73.800 206.100 ;
        RECT 97.400 206.100 97.800 206.200 ;
        RECT 101.400 206.100 101.800 206.200 ;
        RECT 97.400 205.800 101.800 206.100 ;
        RECT 102.200 206.100 102.600 206.200 ;
        RECT 104.600 206.100 105.000 206.200 ;
        RECT 102.200 205.800 105.000 206.100 ;
        RECT 105.400 206.100 105.800 206.200 ;
        RECT 112.600 206.100 113.000 206.200 ;
        RECT 105.400 205.800 113.000 206.100 ;
        RECT 127.800 206.100 128.200 206.200 ;
        RECT 128.600 206.100 129.000 206.200 ;
        RECT 138.200 206.100 138.600 206.200 ;
        RECT 127.800 205.800 138.600 206.100 ;
        RECT 139.800 206.100 140.200 206.200 ;
        RECT 142.200 206.100 142.600 206.200 ;
        RECT 139.800 205.800 142.600 206.100 ;
        RECT 147.800 206.100 148.200 206.200 ;
        RECT 194.200 206.100 194.600 206.200 ;
        RECT 197.400 206.100 197.800 206.200 ;
        RECT 147.800 205.800 197.800 206.100 ;
        RECT 199.000 206.100 199.400 206.200 ;
        RECT 199.800 206.100 200.200 206.200 ;
        RECT 199.000 205.800 200.200 206.100 ;
        RECT 211.800 205.800 212.200 206.200 ;
        RECT 213.400 205.800 213.800 206.200 ;
        RECT 219.000 206.100 219.400 206.200 ;
        RECT 220.600 206.100 221.000 206.200 ;
        RECT 219.000 205.800 221.000 206.100 ;
        RECT 233.400 206.100 233.800 206.200 ;
        RECT 235.800 206.100 236.200 206.200 ;
        RECT 248.600 206.100 249.000 206.200 ;
        RECT 233.400 205.800 236.200 206.100 ;
        RECT 247.000 205.800 249.000 206.100 ;
        RECT 40.600 205.200 40.900 205.800 ;
        RECT 71.800 205.200 72.100 205.800 ;
        RECT 98.200 205.200 98.500 205.800 ;
        RECT 112.600 205.200 112.900 205.800 ;
        RECT 247.000 205.200 247.300 205.800 ;
        RECT 11.000 205.100 11.400 205.200 ;
        RECT 13.400 205.100 13.800 205.200 ;
        RECT 11.000 204.800 13.800 205.100 ;
        RECT 32.600 205.100 33.000 205.200 ;
        RECT 39.000 205.100 39.400 205.200 ;
        RECT 32.600 204.800 39.400 205.100 ;
        RECT 40.600 204.800 41.000 205.200 ;
        RECT 44.600 205.100 45.000 205.200 ;
        RECT 59.000 205.100 59.400 205.200 ;
        RECT 44.600 204.800 59.400 205.100 ;
        RECT 71.800 204.800 72.200 205.200 ;
        RECT 98.200 204.800 98.600 205.200 ;
        RECT 112.600 204.800 113.000 205.200 ;
        RECT 121.400 205.100 121.800 205.200 ;
        RECT 133.400 205.100 133.800 205.200 ;
        RECT 121.400 204.800 133.800 205.100 ;
        RECT 169.400 205.100 169.800 205.200 ;
        RECT 180.600 205.100 181.000 205.200 ;
        RECT 169.400 204.800 181.000 205.100 ;
        RECT 192.600 205.100 193.000 205.200 ;
        RECT 193.400 205.100 193.800 205.200 ;
        RECT 192.600 204.800 193.800 205.100 ;
        RECT 196.600 205.100 197.000 205.200 ;
        RECT 208.600 205.100 209.000 205.200 ;
        RECT 196.600 204.800 209.000 205.100 ;
        RECT 231.000 205.100 231.400 205.200 ;
        RECT 234.200 205.100 234.600 205.200 ;
        RECT 231.000 204.800 234.600 205.100 ;
        RECT 247.000 204.800 247.400 205.200 ;
        RECT 13.400 204.200 13.700 204.800 ;
        RECT 13.400 203.800 13.800 204.200 ;
        RECT 55.800 204.100 56.200 204.200 ;
        RECT 63.000 204.100 63.400 204.200 ;
        RECT 55.800 203.800 63.400 204.100 ;
        RECT 79.800 204.100 80.200 204.200 ;
        RECT 82.200 204.100 82.600 204.200 ;
        RECT 79.800 203.800 82.600 204.100 ;
        RECT 89.400 204.100 89.800 204.200 ;
        RECT 102.200 204.100 102.600 204.200 ;
        RECT 89.400 203.800 102.600 204.100 ;
        RECT 104.600 204.100 105.000 204.200 ;
        RECT 166.200 204.100 166.600 204.200 ;
        RECT 168.600 204.100 169.000 204.200 ;
        RECT 205.400 204.100 205.800 204.200 ;
        RECT 104.600 203.800 205.800 204.100 ;
        RECT 95.000 203.100 95.400 203.200 ;
        RECT 103.000 203.100 103.400 203.200 ;
        RECT 95.000 202.800 103.400 203.100 ;
        RECT 113.400 203.100 113.800 203.200 ;
        RECT 115.800 203.100 116.200 203.200 ;
        RECT 113.400 202.800 116.200 203.100 ;
        RECT 130.200 203.100 130.600 203.200 ;
        RECT 187.800 203.100 188.200 203.200 ;
        RECT 130.200 202.800 188.200 203.100 ;
        RECT 244.600 203.100 245.000 203.200 ;
        RECT 247.000 203.100 247.400 203.200 ;
        RECT 244.600 202.800 247.400 203.100 ;
        RECT 34.200 202.100 34.600 202.200 ;
        RECT 50.200 202.100 50.600 202.200 ;
        RECT 34.200 201.800 50.600 202.100 ;
        RECT 59.000 202.100 59.400 202.200 ;
        RECT 64.600 202.100 65.000 202.200 ;
        RECT 70.200 202.100 70.600 202.200 ;
        RECT 59.000 201.800 70.600 202.100 ;
        RECT 112.600 202.100 113.000 202.200 ;
        RECT 143.800 202.100 144.200 202.200 ;
        RECT 147.800 202.100 148.200 202.200 ;
        RECT 112.600 201.800 148.200 202.100 ;
        RECT 60.600 201.100 61.000 201.200 ;
        RECT 112.600 201.100 113.000 201.200 ;
        RECT 60.600 200.800 113.000 201.100 ;
        RECT 115.000 201.100 115.400 201.200 ;
        RECT 136.600 201.100 137.000 201.200 ;
        RECT 115.000 200.800 137.000 201.100 ;
        RECT 156.600 201.100 157.000 201.200 ;
        RECT 161.400 201.100 161.800 201.200 ;
        RECT 156.600 200.800 161.800 201.100 ;
        RECT 172.600 201.100 173.000 201.200 ;
        RECT 243.800 201.100 244.200 201.200 ;
        RECT 251.800 201.100 252.200 201.200 ;
        RECT 172.600 200.800 252.200 201.100 ;
        RECT 76.600 200.100 77.000 200.200 ;
        RECT 127.000 200.100 127.400 200.200 ;
        RECT 76.600 199.800 127.400 200.100 ;
        RECT 132.600 200.100 133.000 200.200 ;
        RECT 144.600 200.100 145.000 200.200 ;
        RECT 132.600 199.800 145.000 200.100 ;
        RECT 195.000 200.100 195.400 200.200 ;
        RECT 222.200 200.100 222.600 200.200 ;
        RECT 195.000 199.800 222.600 200.100 ;
        RECT 19.000 199.100 19.400 199.200 ;
        RECT 23.000 199.100 23.400 199.200 ;
        RECT 19.000 198.800 23.400 199.100 ;
        RECT 27.000 199.100 27.400 199.200 ;
        RECT 44.600 199.100 45.000 199.200 ;
        RECT 74.200 199.100 74.600 199.200 ;
        RECT 75.000 199.100 75.400 199.200 ;
        RECT 27.000 198.800 75.400 199.100 ;
        RECT 97.400 199.100 97.800 199.200 ;
        RECT 160.600 199.100 161.000 199.200 ;
        RECT 97.400 198.800 161.000 199.100 ;
        RECT 222.200 199.100 222.600 199.200 ;
        RECT 224.600 199.100 225.000 199.200 ;
        RECT 222.200 198.800 225.000 199.100 ;
        RECT 50.200 198.100 50.600 198.200 ;
        RECT 55.800 198.100 56.200 198.200 ;
        RECT 50.200 197.800 56.200 198.100 ;
        RECT 126.200 197.800 126.600 198.200 ;
        RECT 127.000 198.100 127.400 198.200 ;
        RECT 139.800 198.100 140.200 198.200 ;
        RECT 140.600 198.100 141.000 198.200 ;
        RECT 127.000 197.800 141.000 198.100 ;
        RECT 141.400 198.100 141.800 198.200 ;
        RECT 163.000 198.100 163.400 198.200 ;
        RECT 141.400 197.800 163.400 198.100 ;
        RECT 166.200 198.100 166.600 198.200 ;
        RECT 166.200 197.800 173.700 198.100 ;
        RECT 126.200 197.200 126.500 197.800 ;
        RECT 173.400 197.200 173.700 197.800 ;
        RECT 186.200 197.800 186.600 198.200 ;
        RECT 218.200 198.100 218.600 198.200 ;
        RECT 221.400 198.100 221.800 198.200 ;
        RECT 218.200 197.800 221.800 198.100 ;
        RECT 231.000 198.100 231.400 198.200 ;
        RECT 236.600 198.100 237.000 198.200 ;
        RECT 248.600 198.100 249.000 198.200 ;
        RECT 231.000 197.800 249.000 198.100 ;
        RECT 186.200 197.200 186.500 197.800 ;
        RECT 6.200 197.100 6.600 197.200 ;
        RECT 10.200 197.100 10.600 197.200 ;
        RECT 6.200 196.800 10.600 197.100 ;
        RECT 27.000 197.100 27.400 197.200 ;
        RECT 40.600 197.100 41.000 197.200 ;
        RECT 46.200 197.100 46.600 197.200 ;
        RECT 27.000 196.800 46.600 197.100 ;
        RECT 67.800 196.800 68.200 197.200 ;
        RECT 126.200 196.800 126.600 197.200 ;
        RECT 135.000 197.100 135.400 197.200 ;
        RECT 160.600 197.100 161.000 197.200 ;
        RECT 169.400 197.100 169.800 197.200 ;
        RECT 135.000 196.800 169.800 197.100 ;
        RECT 173.400 196.800 173.800 197.200 ;
        RECT 186.200 196.800 186.600 197.200 ;
        RECT 209.400 197.100 209.800 197.200 ;
        RECT 224.600 197.100 225.000 197.200 ;
        RECT 209.400 196.800 225.000 197.100 ;
        RECT 243.000 197.100 243.400 197.200 ;
        RECT 251.800 197.100 252.200 197.200 ;
        RECT 243.000 196.800 252.200 197.100 ;
        RECT 31.800 196.100 32.200 196.200 ;
        RECT 35.000 196.100 35.400 196.200 ;
        RECT 31.000 195.800 35.400 196.100 ;
        RECT 51.000 196.100 51.400 196.200 ;
        RECT 52.600 196.100 53.000 196.200 ;
        RECT 51.000 195.800 53.000 196.100 ;
        RECT 64.600 196.100 65.000 196.200 ;
        RECT 65.400 196.100 65.800 196.200 ;
        RECT 64.600 195.800 65.800 196.100 ;
        RECT 67.800 196.100 68.100 196.800 ;
        RECT 68.600 196.100 69.000 196.200 ;
        RECT 67.800 195.800 69.000 196.100 ;
        RECT 71.000 196.100 71.400 196.200 ;
        RECT 95.800 196.100 96.200 196.200 ;
        RECT 71.000 195.800 96.200 196.100 ;
        RECT 96.600 196.100 97.000 196.200 ;
        RECT 101.400 196.100 101.800 196.200 ;
        RECT 96.600 195.800 101.800 196.100 ;
        RECT 120.600 195.800 121.000 196.200 ;
        RECT 132.600 196.100 133.000 196.200 ;
        RECT 165.400 196.100 165.800 196.200 ;
        RECT 181.400 196.100 181.800 196.200 ;
        RECT 132.600 195.800 181.800 196.100 ;
        RECT 199.800 196.100 200.200 196.200 ;
        RECT 207.800 196.100 208.200 196.200 ;
        RECT 199.800 195.800 208.200 196.100 ;
        RECT 208.600 196.100 209.000 196.200 ;
        RECT 214.200 196.100 214.600 196.200 ;
        RECT 208.600 195.800 214.600 196.100 ;
        RECT 216.600 196.100 217.000 196.200 ;
        RECT 218.200 196.100 218.600 196.200 ;
        RECT 219.800 196.100 220.200 196.200 ;
        RECT 216.600 195.800 220.200 196.100 ;
        RECT 222.200 196.100 222.600 196.200 ;
        RECT 227.000 196.100 227.400 196.200 ;
        RECT 222.200 195.800 227.400 196.100 ;
        RECT 232.600 195.800 233.000 196.200 ;
        RECT 242.200 196.100 242.600 196.200 ;
        RECT 244.600 196.100 245.000 196.200 ;
        RECT 242.200 195.800 245.000 196.100 ;
        RECT 8.600 195.100 9.000 195.200 ;
        RECT 28.600 195.100 29.000 195.200 ;
        RECT 31.000 195.100 31.400 195.200 ;
        RECT 8.600 194.800 12.900 195.100 ;
        RECT 28.600 194.800 31.400 195.100 ;
        RECT 41.400 195.100 41.800 195.200 ;
        RECT 41.400 194.800 45.700 195.100 ;
        RECT 12.600 194.200 12.900 194.800 ;
        RECT 45.400 194.200 45.700 194.800 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 58.200 195.100 58.600 195.200 ;
        RECT 60.600 195.100 61.000 195.200 ;
        RECT 58.200 194.800 61.000 195.100 ;
        RECT 62.200 195.100 62.600 195.200 ;
        RECT 63.000 195.100 63.400 195.200 ;
        RECT 62.200 194.800 63.400 195.100 ;
        RECT 68.600 194.800 69.000 195.200 ;
        RECT 70.200 194.800 70.600 195.200 ;
        RECT 79.800 195.100 80.200 195.200 ;
        RECT 80.600 195.100 81.000 195.200 ;
        RECT 79.800 194.800 81.000 195.100 ;
        RECT 95.000 195.100 95.400 195.200 ;
        RECT 95.800 195.100 96.200 195.200 ;
        RECT 95.000 194.800 96.200 195.100 ;
        RECT 100.600 195.100 101.000 195.200 ;
        RECT 107.800 195.100 108.200 195.200 ;
        RECT 100.600 194.800 108.200 195.100 ;
        RECT 111.000 195.100 111.400 195.200 ;
        RECT 120.600 195.100 120.900 195.800 ;
        RECT 232.600 195.200 232.900 195.800 ;
        RECT 131.800 195.100 132.200 195.200 ;
        RECT 111.000 194.800 120.900 195.100 ;
        RECT 130.200 194.800 132.200 195.100 ;
        RECT 140.600 194.800 141.000 195.200 ;
        RECT 143.000 195.100 143.400 195.200 ;
        RECT 143.800 195.100 144.200 195.200 ;
        RECT 143.000 194.800 144.200 195.100 ;
        RECT 147.000 195.100 147.400 195.200 ;
        RECT 157.400 195.100 157.800 195.200 ;
        RECT 147.000 194.800 157.800 195.100 ;
        RECT 171.000 195.100 171.400 195.200 ;
        RECT 172.600 195.100 173.000 195.200 ;
        RECT 171.000 194.800 173.000 195.100 ;
        RECT 193.400 195.100 193.800 195.200 ;
        RECT 195.800 195.100 196.200 195.200 ;
        RECT 193.400 194.800 196.200 195.100 ;
        RECT 200.600 195.100 201.000 195.200 ;
        RECT 215.800 195.100 216.200 195.200 ;
        RECT 200.600 194.800 216.200 195.100 ;
        RECT 219.000 195.100 219.400 195.200 ;
        RECT 226.200 195.100 226.600 195.200 ;
        RECT 219.000 194.800 226.600 195.100 ;
        RECT 232.600 194.800 233.000 195.200 ;
        RECT 233.400 195.100 233.800 195.200 ;
        RECT 238.200 195.100 238.600 195.200 ;
        RECT 233.400 194.800 238.600 195.100 ;
        RECT 51.800 194.200 52.100 194.800 ;
        RECT 60.600 194.200 60.900 194.800 ;
        RECT 68.600 194.200 68.900 194.800 ;
        RECT 70.200 194.200 70.500 194.800 ;
        RECT 130.200 194.200 130.500 194.800 ;
        RECT 140.600 194.200 140.900 194.800 ;
        RECT 200.600 194.200 200.900 194.800 ;
        RECT 12.600 193.800 13.000 194.200 ;
        RECT 43.000 194.100 43.400 194.200 ;
        RECT 31.800 193.800 43.400 194.100 ;
        RECT 45.400 193.800 45.800 194.200 ;
        RECT 51.800 193.800 52.200 194.200 ;
        RECT 60.600 193.800 61.000 194.200 ;
        RECT 64.600 194.100 65.000 194.200 ;
        RECT 65.400 194.100 65.800 194.200 ;
        RECT 64.600 193.800 65.800 194.100 ;
        RECT 68.600 193.800 69.000 194.200 ;
        RECT 70.200 193.800 70.600 194.200 ;
        RECT 72.600 193.800 73.000 194.200 ;
        RECT 77.400 194.100 77.800 194.200 ;
        RECT 79.800 194.100 80.200 194.200 ;
        RECT 106.200 194.100 106.600 194.200 ;
        RECT 77.400 193.800 80.200 194.100 ;
        RECT 89.400 193.800 106.600 194.100 ;
        RECT 115.000 194.100 115.400 194.200 ;
        RECT 127.800 194.100 128.200 194.200 ;
        RECT 115.000 193.800 128.200 194.100 ;
        RECT 130.200 193.800 130.600 194.200 ;
        RECT 137.400 193.800 137.800 194.200 ;
        RECT 140.600 194.100 141.000 194.200 ;
        RECT 143.800 194.100 144.200 194.200 ;
        RECT 140.600 193.800 144.200 194.100 ;
        RECT 144.600 193.800 145.000 194.200 ;
        RECT 149.400 194.100 149.800 194.200 ;
        RECT 152.600 194.100 153.000 194.200 ;
        RECT 149.400 193.800 153.000 194.100 ;
        RECT 200.600 193.800 201.000 194.200 ;
        RECT 208.600 194.100 209.000 194.200 ;
        RECT 213.400 194.100 213.800 194.200 ;
        RECT 215.800 194.100 216.200 194.200 ;
        RECT 225.400 194.100 225.800 194.200 ;
        RECT 208.600 193.800 225.800 194.100 ;
        RECT 244.600 194.100 245.000 194.200 ;
        RECT 246.200 194.100 246.600 194.200 ;
        RECT 244.600 193.800 246.600 194.100 ;
        RECT 31.800 193.200 32.100 193.800 ;
        RECT 31.800 192.800 32.200 193.200 ;
        RECT 61.400 193.100 61.800 193.200 ;
        RECT 63.800 193.100 64.200 193.200 ;
        RECT 72.600 193.100 72.900 193.800 ;
        RECT 61.400 192.800 72.900 193.100 ;
        RECT 89.400 193.200 89.700 193.800 ;
        RECT 137.400 193.200 137.700 193.800 ;
        RECT 144.600 193.200 144.900 193.800 ;
        RECT 246.200 193.200 246.500 193.800 ;
        RECT 89.400 192.800 89.800 193.200 ;
        RECT 95.000 193.100 95.400 193.200 ;
        RECT 96.600 193.100 97.000 193.200 ;
        RECT 95.000 192.800 97.000 193.100 ;
        RECT 117.400 193.100 117.800 193.200 ;
        RECT 125.400 193.100 125.800 193.200 ;
        RECT 117.400 192.800 125.800 193.100 ;
        RECT 137.400 192.800 137.800 193.200 ;
        RECT 144.600 192.800 145.000 193.200 ;
        RECT 147.800 193.100 148.200 193.200 ;
        RECT 158.200 193.100 158.600 193.200 ;
        RECT 147.800 192.800 158.600 193.100 ;
        RECT 191.000 193.100 191.400 193.200 ;
        RECT 191.800 193.100 192.200 193.200 ;
        RECT 191.000 192.800 192.200 193.100 ;
        RECT 246.200 192.800 246.600 193.200 ;
        RECT 21.400 191.800 21.800 192.200 ;
        RECT 67.800 192.100 68.200 192.200 ;
        RECT 93.400 192.100 93.800 192.200 ;
        RECT 67.800 191.800 93.800 192.100 ;
        RECT 115.800 192.100 116.200 192.200 ;
        RECT 118.200 192.100 118.600 192.200 ;
        RECT 141.400 192.100 141.800 192.200 ;
        RECT 115.800 191.800 141.800 192.100 ;
        RECT 143.800 192.100 144.200 192.200 ;
        RECT 187.800 192.100 188.200 192.200 ;
        RECT 143.800 191.800 188.200 192.100 ;
        RECT 188.600 192.100 189.000 192.200 ;
        RECT 194.200 192.100 194.600 192.200 ;
        RECT 188.600 191.800 194.600 192.100 ;
        RECT 197.400 192.100 197.800 192.200 ;
        RECT 203.800 192.100 204.200 192.200 ;
        RECT 213.400 192.100 213.800 192.200 ;
        RECT 197.400 191.800 213.800 192.100 ;
        RECT 218.200 192.100 218.600 192.200 ;
        RECT 233.400 192.100 233.800 192.200 ;
        RECT 218.200 191.800 233.800 192.100 ;
        RECT 21.400 191.200 21.700 191.800 ;
        RECT 21.400 190.800 21.800 191.200 ;
        RECT 129.400 191.100 129.800 191.200 ;
        RECT 153.400 191.100 153.800 191.200 ;
        RECT 129.400 190.800 153.800 191.100 ;
        RECT 187.000 191.100 187.400 191.200 ;
        RECT 190.200 191.100 190.600 191.200 ;
        RECT 187.000 190.800 190.600 191.100 ;
        RECT 210.200 191.100 210.600 191.200 ;
        RECT 231.800 191.100 232.200 191.200 ;
        RECT 210.200 190.800 232.200 191.100 ;
        RECT 80.600 190.100 81.000 190.200 ;
        RECT 90.200 190.100 90.600 190.200 ;
        RECT 95.800 190.100 96.200 190.200 ;
        RECT 80.600 189.800 96.200 190.100 ;
        RECT 123.800 190.100 124.200 190.200 ;
        RECT 144.600 190.100 145.000 190.200 ;
        RECT 123.800 189.800 145.000 190.100 ;
        RECT 211.800 190.100 212.200 190.200 ;
        RECT 219.800 190.100 220.200 190.200 ;
        RECT 211.800 189.800 220.200 190.100 ;
        RECT 34.200 188.800 34.600 189.200 ;
        RECT 40.600 189.100 41.000 189.200 ;
        RECT 47.000 189.100 47.400 189.200 ;
        RECT 48.600 189.100 49.000 189.200 ;
        RECT 40.600 188.800 49.000 189.100 ;
        RECT 54.200 189.100 54.600 189.200 ;
        RECT 71.800 189.100 72.200 189.200 ;
        RECT 54.200 188.800 72.200 189.100 ;
        RECT 87.800 189.100 88.200 189.200 ;
        RECT 92.600 189.100 93.000 189.200 ;
        RECT 87.800 188.800 93.000 189.100 ;
        RECT 130.200 189.100 130.600 189.200 ;
        RECT 131.000 189.100 131.400 189.200 ;
        RECT 130.200 188.800 131.400 189.100 ;
        RECT 131.800 189.100 132.200 189.200 ;
        RECT 147.800 189.100 148.200 189.200 ;
        RECT 131.800 188.800 148.200 189.100 ;
        RECT 148.600 189.100 149.000 189.200 ;
        RECT 151.800 189.100 152.200 189.200 ;
        RECT 160.600 189.100 161.000 189.200 ;
        RECT 165.400 189.100 165.800 189.200 ;
        RECT 148.600 188.800 152.900 189.100 ;
        RECT 160.600 188.800 165.800 189.100 ;
        RECT 179.000 189.100 179.400 189.200 ;
        RECT 186.200 189.100 186.600 189.200 ;
        RECT 189.400 189.100 189.800 189.200 ;
        RECT 179.000 188.800 189.800 189.100 ;
        RECT 199.800 189.100 200.200 189.200 ;
        RECT 203.000 189.100 203.400 189.200 ;
        RECT 199.800 188.800 203.400 189.100 ;
        RECT 233.400 188.800 233.800 189.200 ;
        RECT 34.200 188.100 34.500 188.800 ;
        RECT 43.800 188.100 44.200 188.200 ;
        RECT 51.000 188.100 51.400 188.200 ;
        RECT 34.200 187.800 51.400 188.100 ;
        RECT 55.800 188.100 56.200 188.200 ;
        RECT 63.000 188.100 63.400 188.200 ;
        RECT 55.800 187.800 63.400 188.100 ;
        RECT 65.400 188.100 65.800 188.200 ;
        RECT 81.400 188.100 81.800 188.200 ;
        RECT 91.000 188.100 91.400 188.200 ;
        RECT 65.400 187.800 91.400 188.100 ;
        RECT 95.800 188.100 96.200 188.200 ;
        RECT 117.400 188.100 117.800 188.200 ;
        RECT 95.800 187.800 117.800 188.100 ;
        RECT 125.400 188.100 125.800 188.200 ;
        RECT 155.000 188.100 155.400 188.200 ;
        RECT 125.400 187.800 155.400 188.100 ;
        RECT 174.200 187.800 174.600 188.200 ;
        RECT 186.200 188.100 186.600 188.200 ;
        RECT 187.000 188.100 187.400 188.200 ;
        RECT 186.200 187.800 187.400 188.100 ;
        RECT 229.400 188.100 229.800 188.200 ;
        RECT 233.400 188.100 233.700 188.800 ;
        RECT 229.400 187.800 233.700 188.100 ;
        RECT 247.000 188.100 247.400 188.200 ;
        RECT 250.200 188.100 250.600 188.200 ;
        RECT 247.000 187.800 250.600 188.100 ;
        RECT 1.400 187.100 1.800 187.200 ;
        RECT 11.000 187.100 11.400 187.200 ;
        RECT 1.400 186.800 11.400 187.100 ;
        RECT 20.600 187.100 21.000 187.200 ;
        RECT 22.200 187.100 22.600 187.200 ;
        RECT 29.400 187.100 29.800 187.200 ;
        RECT 33.400 187.100 33.800 187.200 ;
        RECT 39.000 187.100 39.400 187.200 ;
        RECT 20.600 186.800 39.400 187.100 ;
        RECT 45.400 186.800 45.800 187.200 ;
        RECT 60.600 187.100 61.000 187.200 ;
        RECT 67.000 187.100 67.400 187.200 ;
        RECT 60.600 186.800 67.400 187.100 ;
        RECT 67.800 186.800 68.200 187.200 ;
        RECT 73.400 187.100 73.800 187.200 ;
        RECT 74.200 187.100 74.600 187.200 ;
        RECT 73.400 186.800 74.600 187.100 ;
        RECT 84.600 187.100 85.000 187.200 ;
        RECT 86.200 187.100 86.600 187.200 ;
        RECT 96.600 187.100 97.000 187.200 ;
        RECT 84.600 186.800 97.000 187.100 ;
        RECT 99.800 187.100 100.200 187.200 ;
        RECT 111.000 187.100 111.400 187.200 ;
        RECT 99.800 186.800 111.400 187.100 ;
        RECT 116.600 187.100 117.000 187.200 ;
        RECT 117.400 187.100 117.800 187.200 ;
        RECT 116.600 186.800 117.800 187.100 ;
        RECT 126.200 186.800 126.600 187.200 ;
        RECT 127.000 187.100 127.400 187.200 ;
        RECT 139.800 187.100 140.200 187.200 ;
        RECT 127.000 186.800 140.200 187.100 ;
        RECT 143.000 187.100 143.400 187.200 ;
        RECT 144.600 187.100 145.000 187.200 ;
        RECT 148.600 187.100 149.000 187.200 ;
        RECT 143.000 186.800 149.000 187.100 ;
        RECT 149.400 187.100 149.800 187.200 ;
        RECT 152.600 187.100 153.000 187.200 ;
        RECT 149.400 186.800 153.000 187.100 ;
        RECT 154.200 186.800 154.600 187.200 ;
        RECT 158.200 187.100 158.600 187.200 ;
        RECT 162.200 187.100 162.600 187.200 ;
        RECT 174.200 187.100 174.500 187.800 ;
        RECT 175.000 187.100 175.400 187.200 ;
        RECT 179.800 187.100 180.200 187.200 ;
        RECT 158.200 186.800 180.200 187.100 ;
        RECT 183.000 187.100 183.400 187.200 ;
        RECT 195.800 187.100 196.200 187.200 ;
        RECT 207.000 187.100 207.400 187.200 ;
        RECT 183.000 186.800 196.200 187.100 ;
        RECT 198.200 186.800 207.400 187.100 ;
        RECT 233.400 186.800 233.800 187.200 ;
        RECT 7.800 186.100 8.200 186.200 ;
        RECT 9.400 186.100 9.800 186.200 ;
        RECT 7.800 185.800 9.800 186.100 ;
        RECT 11.800 186.100 12.200 186.200 ;
        RECT 14.200 186.100 14.600 186.200 ;
        RECT 19.000 186.100 19.400 186.200 ;
        RECT 11.800 185.800 19.400 186.100 ;
        RECT 23.800 186.100 24.200 186.200 ;
        RECT 33.400 186.100 33.800 186.200 ;
        RECT 35.000 186.100 35.400 186.200 ;
        RECT 23.800 185.800 32.100 186.100 ;
        RECT 33.400 185.800 35.400 186.100 ;
        RECT 43.000 186.100 43.400 186.200 ;
        RECT 45.400 186.100 45.700 186.800 ;
        RECT 43.000 185.800 45.700 186.100 ;
        RECT 47.000 186.100 47.400 186.200 ;
        RECT 57.400 186.100 57.800 186.200 ;
        RECT 67.800 186.100 68.100 186.800 ;
        RECT 47.000 185.800 57.800 186.100 ;
        RECT 63.800 185.800 68.100 186.100 ;
        RECT 71.800 185.800 72.200 186.200 ;
        RECT 80.600 186.100 81.000 186.200 ;
        RECT 87.800 186.100 88.200 186.200 ;
        RECT 80.600 185.800 88.200 186.100 ;
        RECT 107.000 186.100 107.400 186.200 ;
        RECT 114.200 186.100 114.600 186.200 ;
        RECT 107.000 185.800 114.600 186.100 ;
        RECT 119.800 186.100 120.200 186.200 ;
        RECT 126.200 186.100 126.500 186.800 ;
        RECT 154.200 186.200 154.500 186.800 ;
        RECT 198.200 186.200 198.500 186.800 ;
        RECT 119.800 185.800 126.500 186.100 ;
        RECT 131.000 185.800 131.400 186.200 ;
        RECT 141.400 186.100 141.800 186.200 ;
        RECT 150.200 186.100 150.600 186.200 ;
        RECT 141.400 185.800 150.600 186.100 ;
        RECT 154.200 185.800 154.600 186.200 ;
        RECT 161.400 185.800 161.800 186.200 ;
        RECT 165.400 186.100 165.800 186.200 ;
        RECT 169.400 186.100 169.800 186.200 ;
        RECT 165.400 185.800 169.800 186.100 ;
        RECT 184.600 186.100 185.000 186.200 ;
        RECT 185.400 186.100 185.800 186.200 ;
        RECT 184.600 185.800 185.800 186.100 ;
        RECT 187.800 186.100 188.200 186.200 ;
        RECT 188.600 186.100 189.000 186.200 ;
        RECT 187.800 185.800 189.000 186.100 ;
        RECT 198.200 185.800 198.600 186.200 ;
        RECT 199.800 185.800 200.200 186.200 ;
        RECT 209.400 186.100 209.800 186.200 ;
        RECT 215.000 186.100 215.400 186.200 ;
        RECT 209.400 185.800 215.400 186.100 ;
        RECT 217.400 186.100 217.800 186.200 ;
        RECT 218.200 186.100 218.600 186.200 ;
        RECT 217.400 185.800 218.600 186.100 ;
        RECT 228.600 186.100 229.000 186.200 ;
        RECT 233.400 186.100 233.700 186.800 ;
        RECT 228.600 185.800 233.700 186.100 ;
        RECT 31.800 185.200 32.100 185.800 ;
        RECT 57.400 185.200 57.700 185.800 ;
        RECT 63.800 185.200 64.100 185.800 ;
        RECT 71.800 185.200 72.100 185.800 ;
        RECT 131.000 185.200 131.300 185.800 ;
        RECT 3.000 185.100 3.400 185.200 ;
        RECT 4.600 185.100 5.000 185.200 ;
        RECT 29.400 185.100 29.800 185.200 ;
        RECT 3.000 184.800 5.000 185.100 ;
        RECT 13.400 184.800 29.800 185.100 ;
        RECT 31.800 184.800 32.200 185.200 ;
        RECT 43.800 185.100 44.200 185.200 ;
        RECT 53.400 185.100 53.800 185.200 ;
        RECT 43.800 184.800 53.800 185.100 ;
        RECT 57.400 184.800 57.800 185.200 ;
        RECT 63.800 184.800 64.200 185.200 ;
        RECT 66.200 185.100 66.600 185.200 ;
        RECT 67.000 185.100 67.400 185.200 ;
        RECT 66.200 184.800 67.400 185.100 ;
        RECT 71.800 184.800 72.200 185.200 ;
        RECT 87.800 185.100 88.200 185.200 ;
        RECT 89.400 185.100 89.800 185.200 ;
        RECT 87.800 184.800 89.800 185.100 ;
        RECT 115.000 185.100 115.400 185.200 ;
        RECT 118.200 185.100 118.600 185.200 ;
        RECT 115.000 184.800 118.600 185.100 ;
        RECT 131.000 184.800 131.400 185.200 ;
        RECT 132.600 184.800 133.000 185.200 ;
        RECT 146.200 185.100 146.600 185.200 ;
        RECT 156.600 185.100 157.000 185.200 ;
        RECT 146.200 184.800 157.000 185.100 ;
        RECT 157.400 185.100 157.800 185.200 ;
        RECT 158.200 185.100 158.600 185.200 ;
        RECT 157.400 184.800 158.600 185.100 ;
        RECT 161.400 185.100 161.700 185.800 ;
        RECT 164.600 185.100 165.000 185.200 ;
        RECT 161.400 184.800 165.000 185.100 ;
        RECT 171.000 185.100 171.400 185.200 ;
        RECT 199.800 185.100 200.100 185.800 ;
        RECT 171.000 184.800 200.100 185.100 ;
        RECT 218.200 185.100 218.600 185.200 ;
        RECT 224.600 185.100 225.000 185.200 ;
        RECT 218.200 184.800 225.000 185.100 ;
        RECT 226.200 185.100 226.600 185.200 ;
        RECT 227.800 185.100 228.200 185.200 ;
        RECT 241.400 185.100 241.800 185.200 ;
        RECT 226.200 184.800 241.800 185.100 ;
        RECT 13.400 184.200 13.700 184.800 ;
        RECT 132.600 184.200 132.900 184.800 ;
        RECT 13.400 183.800 13.800 184.200 ;
        RECT 15.800 184.100 16.200 184.200 ;
        RECT 38.200 184.100 38.600 184.200 ;
        RECT 15.800 183.800 38.600 184.100 ;
        RECT 53.400 184.100 53.800 184.200 ;
        RECT 62.200 184.100 62.600 184.200 ;
        RECT 53.400 183.800 62.600 184.100 ;
        RECT 66.200 184.100 66.600 184.200 ;
        RECT 107.000 184.100 107.400 184.200 ;
        RECT 66.200 183.800 107.400 184.100 ;
        RECT 132.600 183.800 133.000 184.200 ;
        RECT 139.000 184.100 139.400 184.200 ;
        RECT 147.000 184.100 147.400 184.200 ;
        RECT 139.000 183.800 147.400 184.100 ;
        RECT 147.800 184.100 148.200 184.200 ;
        RECT 160.600 184.100 161.000 184.200 ;
        RECT 147.800 183.800 161.000 184.100 ;
        RECT 181.400 184.100 181.800 184.200 ;
        RECT 183.000 184.100 183.400 184.200 ;
        RECT 183.800 184.100 184.200 184.200 ;
        RECT 181.400 183.800 184.200 184.100 ;
        RECT 185.400 184.100 185.800 184.200 ;
        RECT 186.200 184.100 186.600 184.200 ;
        RECT 185.400 183.800 186.600 184.100 ;
        RECT 189.400 184.100 189.800 184.200 ;
        RECT 199.800 184.100 200.200 184.200 ;
        RECT 189.400 183.800 200.200 184.100 ;
        RECT 57.400 183.100 57.800 183.200 ;
        RECT 69.400 183.100 69.800 183.200 ;
        RECT 57.400 182.800 69.800 183.100 ;
        RECT 79.800 183.100 80.200 183.200 ;
        RECT 103.800 183.100 104.200 183.200 ;
        RECT 79.800 182.800 104.200 183.100 ;
        RECT 147.800 183.100 148.200 183.200 ;
        RECT 178.200 183.100 178.600 183.200 ;
        RECT 147.800 182.800 178.600 183.100 ;
        RECT 181.400 183.100 181.800 183.200 ;
        RECT 214.200 183.100 214.600 183.200 ;
        RECT 215.000 183.100 215.400 183.200 ;
        RECT 181.400 182.800 215.400 183.100 ;
        RECT 230.200 183.100 230.600 183.200 ;
        RECT 239.000 183.100 239.400 183.200 ;
        RECT 230.200 182.800 239.400 183.100 ;
        RECT 42.200 182.100 42.600 182.200 ;
        RECT 44.600 182.100 45.000 182.200 ;
        RECT 85.400 182.100 85.800 182.200 ;
        RECT 42.200 181.800 85.800 182.100 ;
        RECT 87.000 182.100 87.400 182.200 ;
        RECT 92.600 182.100 93.000 182.200 ;
        RECT 95.000 182.100 95.400 182.200 ;
        RECT 162.200 182.100 162.600 182.200 ;
        RECT 232.600 182.100 233.000 182.200 ;
        RECT 87.000 181.800 233.000 182.100 ;
        RECT 239.800 182.100 240.200 182.200 ;
        RECT 245.400 182.100 245.800 182.200 ;
        RECT 239.800 181.800 245.800 182.100 ;
        RECT 247.800 182.100 248.200 182.200 ;
        RECT 248.600 182.100 249.000 182.200 ;
        RECT 247.800 181.800 249.000 182.100 ;
        RECT 50.200 181.100 50.600 181.200 ;
        RECT 105.400 181.100 105.800 181.200 ;
        RECT 143.000 181.100 143.400 181.200 ;
        RECT 50.200 180.800 143.400 181.100 ;
        RECT 174.200 181.100 174.600 181.200 ;
        RECT 177.400 181.100 177.800 181.200 ;
        RECT 174.200 180.800 177.800 181.100 ;
        RECT 181.400 181.100 181.800 181.200 ;
        RECT 184.600 181.100 185.000 181.200 ;
        RECT 181.400 180.800 185.000 181.100 ;
        RECT 199.000 181.100 199.400 181.200 ;
        RECT 217.400 181.100 217.800 181.200 ;
        RECT 199.000 180.800 217.800 181.100 ;
        RECT 223.800 181.100 224.200 181.200 ;
        RECT 231.000 181.100 231.400 181.200 ;
        RECT 223.800 180.800 231.400 181.100 ;
        RECT 9.400 180.100 9.800 180.200 ;
        RECT 44.600 180.100 45.000 180.200 ;
        RECT 9.400 179.800 45.000 180.100 ;
        RECT 66.200 180.100 66.600 180.200 ;
        RECT 138.200 180.100 138.600 180.200 ;
        RECT 66.200 179.800 138.600 180.100 ;
        RECT 155.000 180.100 155.400 180.200 ;
        RECT 223.000 180.100 223.400 180.200 ;
        RECT 226.200 180.100 226.600 180.200 ;
        RECT 155.000 179.800 226.600 180.100 ;
        RECT 25.400 179.100 25.800 179.200 ;
        RECT 30.200 179.100 30.600 179.200 ;
        RECT 51.000 179.100 51.400 179.200 ;
        RECT 25.400 178.800 29.700 179.100 ;
        RECT 30.200 178.800 51.400 179.100 ;
        RECT 51.800 179.100 52.200 179.200 ;
        RECT 59.000 179.100 59.400 179.200 ;
        RECT 51.800 178.800 59.400 179.100 ;
        RECT 112.600 179.100 113.000 179.200 ;
        RECT 135.000 179.100 135.400 179.200 ;
        RECT 112.600 178.800 135.400 179.100 ;
        RECT 151.800 179.100 152.200 179.200 ;
        RECT 155.800 179.100 156.200 179.200 ;
        RECT 159.000 179.100 159.400 179.200 ;
        RECT 151.800 178.800 159.400 179.100 ;
        RECT 171.800 179.100 172.200 179.200 ;
        RECT 210.200 179.100 210.600 179.200 ;
        RECT 171.800 178.800 210.600 179.100 ;
        RECT 211.800 179.100 212.200 179.200 ;
        RECT 233.400 179.100 233.800 179.200 ;
        RECT 240.600 179.100 241.000 179.200 ;
        RECT 211.800 178.800 241.000 179.100 ;
        RECT 1.400 178.100 1.800 178.200 ;
        RECT 15.000 178.100 15.400 178.200 ;
        RECT 24.600 178.100 25.000 178.200 ;
        RECT 1.400 177.800 25.000 178.100 ;
        RECT 29.400 178.100 29.700 178.800 ;
        RECT 48.600 178.100 49.000 178.200 ;
        RECT 29.400 177.800 49.000 178.100 ;
        RECT 59.000 178.100 59.400 178.200 ;
        RECT 63.800 178.100 64.200 178.200 ;
        RECT 59.000 177.800 64.200 178.100 ;
        RECT 91.800 178.100 92.200 178.200 ;
        RECT 121.400 178.100 121.800 178.200 ;
        RECT 91.800 177.800 121.800 178.100 ;
        RECT 174.200 177.800 174.600 178.200 ;
        RECT 175.800 178.100 176.200 178.200 ;
        RECT 182.200 178.100 182.600 178.200 ;
        RECT 185.400 178.100 185.800 178.200 ;
        RECT 175.800 177.800 185.800 178.100 ;
        RECT 8.600 177.100 9.000 177.200 ;
        RECT 17.400 177.100 17.800 177.200 ;
        RECT 24.600 177.100 25.000 177.200 ;
        RECT 8.600 176.800 25.000 177.100 ;
        RECT 31.000 177.100 31.400 177.200 ;
        RECT 31.800 177.100 32.200 177.200 ;
        RECT 31.000 176.800 32.200 177.100 ;
        RECT 52.600 176.800 53.000 177.200 ;
        RECT 63.000 176.800 63.400 177.200 ;
        RECT 103.000 177.100 103.400 177.200 ;
        RECT 105.400 177.100 105.800 177.200 ;
        RECT 114.200 177.100 114.600 177.200 ;
        RECT 103.000 176.800 114.600 177.100 ;
        RECT 119.800 177.100 120.200 177.200 ;
        RECT 171.800 177.100 172.200 177.200 ;
        RECT 119.800 176.800 172.200 177.100 ;
        RECT 174.200 177.100 174.500 177.800 ;
        RECT 180.600 177.100 181.000 177.200 ;
        RECT 174.200 176.800 181.000 177.100 ;
        RECT 210.200 177.100 210.600 177.200 ;
        RECT 237.400 177.100 237.800 177.200 ;
        RECT 210.200 176.800 237.800 177.100 ;
        RECT 248.600 176.800 249.000 177.200 ;
        RECT 7.000 175.800 7.400 176.200 ;
        RECT 14.200 176.100 14.600 176.200 ;
        RECT 16.600 176.100 17.000 176.200 ;
        RECT 14.200 175.800 17.000 176.100 ;
        RECT 18.200 176.100 18.600 176.200 ;
        RECT 19.000 176.100 19.400 176.200 ;
        RECT 18.200 175.800 19.400 176.100 ;
        RECT 23.000 176.100 23.400 176.200 ;
        RECT 27.000 176.100 27.400 176.200 ;
        RECT 32.600 176.100 33.000 176.200 ;
        RECT 23.000 175.800 33.000 176.100 ;
        RECT 39.800 175.800 40.200 176.200 ;
        RECT 51.000 176.100 51.400 176.200 ;
        RECT 52.600 176.100 52.900 176.800 ;
        RECT 51.000 175.800 52.900 176.100 ;
        RECT 63.000 176.100 63.300 176.800 ;
        RECT 70.200 176.100 70.600 176.200 ;
        RECT 63.000 175.800 70.600 176.100 ;
        RECT 72.600 176.100 73.000 176.200 ;
        RECT 98.200 176.100 98.600 176.200 ;
        RECT 72.600 175.800 98.600 176.100 ;
        RECT 101.400 175.800 101.800 176.200 ;
        RECT 116.600 176.100 117.000 176.200 ;
        RECT 118.200 176.100 118.600 176.200 ;
        RECT 116.600 175.800 118.600 176.100 ;
        RECT 126.200 175.800 126.600 176.200 ;
        RECT 129.400 175.800 129.800 176.200 ;
        RECT 135.000 176.100 135.400 176.200 ;
        RECT 147.800 176.100 148.200 176.200 ;
        RECT 135.000 175.800 148.200 176.100 ;
        RECT 149.400 176.100 149.800 176.200 ;
        RECT 150.200 176.100 150.600 176.200 ;
        RECT 155.000 176.100 155.400 176.200 ;
        RECT 159.800 176.100 160.200 176.200 ;
        RECT 166.200 176.100 166.600 176.200 ;
        RECT 149.400 175.800 150.600 176.100 ;
        RECT 154.200 175.800 159.300 176.100 ;
        RECT 159.800 175.800 166.600 176.100 ;
        RECT 168.600 176.100 169.000 176.200 ;
        RECT 175.800 176.100 176.200 176.200 ;
        RECT 168.600 175.800 176.200 176.100 ;
        RECT 206.200 176.100 206.600 176.200 ;
        RECT 219.800 176.100 220.200 176.200 ;
        RECT 206.200 175.800 220.200 176.100 ;
        RECT 225.400 175.800 225.800 176.200 ;
        RECT 234.200 176.100 234.600 176.200 ;
        RECT 237.400 176.100 237.800 176.200 ;
        RECT 234.200 175.800 237.800 176.100 ;
        RECT 244.600 176.100 245.000 176.200 ;
        RECT 248.600 176.100 248.900 176.800 ;
        RECT 251.000 176.100 251.400 176.200 ;
        RECT 244.600 175.800 248.900 176.100 ;
        RECT 250.200 175.800 251.400 176.100 ;
        RECT 7.000 175.100 7.300 175.800 ;
        RECT 11.800 175.100 12.200 175.200 ;
        RECT 7.000 174.800 12.200 175.100 ;
        RECT 14.200 175.100 14.600 175.200 ;
        RECT 18.200 175.100 18.600 175.200 ;
        RECT 21.400 175.100 21.800 175.200 ;
        RECT 14.200 174.800 21.800 175.100 ;
        RECT 29.400 175.100 29.800 175.200 ;
        RECT 39.800 175.100 40.100 175.800 ;
        RECT 101.400 175.200 101.700 175.800 ;
        RECT 126.200 175.200 126.500 175.800 ;
        RECT 46.200 175.100 46.600 175.200 ;
        RECT 47.000 175.100 47.400 175.200 ;
        RECT 29.400 174.800 36.900 175.100 ;
        RECT 39.800 174.800 44.100 175.100 ;
        RECT 46.200 174.800 47.400 175.100 ;
        RECT 52.600 175.100 53.000 175.200 ;
        RECT 54.200 175.100 54.600 175.200 ;
        RECT 52.600 174.800 54.600 175.100 ;
        RECT 63.800 174.800 64.200 175.200 ;
        RECT 86.200 175.100 86.600 175.200 ;
        RECT 78.200 174.800 86.600 175.100 ;
        RECT 95.800 175.100 96.200 175.200 ;
        RECT 96.600 175.100 97.000 175.200 ;
        RECT 95.800 174.800 97.000 175.100 ;
        RECT 101.400 174.800 101.800 175.200 ;
        RECT 115.800 175.100 116.200 175.200 ;
        RECT 110.200 174.800 116.200 175.100 ;
        RECT 126.200 174.800 126.600 175.200 ;
        RECT 129.400 175.100 129.700 175.800 ;
        RECT 133.400 175.100 133.800 175.200 ;
        RECT 129.400 174.800 133.800 175.100 ;
        RECT 145.400 175.100 145.800 175.200 ;
        RECT 148.600 175.100 149.000 175.200 ;
        RECT 145.400 174.800 149.000 175.100 ;
        RECT 150.200 175.100 150.500 175.800 ;
        RECT 153.400 175.100 153.800 175.200 ;
        RECT 150.200 174.800 153.800 175.100 ;
        RECT 155.000 175.100 155.400 175.200 ;
        RECT 156.600 175.100 157.000 175.200 ;
        RECT 155.000 174.800 157.000 175.100 ;
        RECT 159.000 175.100 159.300 175.800 ;
        RECT 160.600 175.100 161.000 175.200 ;
        RECT 159.000 174.800 161.000 175.100 ;
        RECT 168.600 175.100 168.900 175.800 ;
        RECT 225.400 175.200 225.700 175.800 ;
        RECT 250.200 175.200 250.500 175.800 ;
        RECT 170.200 175.100 170.600 175.200 ;
        RECT 168.600 174.800 170.600 175.100 ;
        RECT 171.800 175.100 172.200 175.200 ;
        RECT 173.400 175.100 173.800 175.200 ;
        RECT 171.800 174.800 173.800 175.100 ;
        RECT 175.000 175.100 175.400 175.200 ;
        RECT 175.800 175.100 176.200 175.200 ;
        RECT 175.000 174.800 176.200 175.100 ;
        RECT 183.800 175.100 184.200 175.200 ;
        RECT 191.800 175.100 192.200 175.200 ;
        RECT 183.800 174.800 192.200 175.100 ;
        RECT 196.600 175.100 197.000 175.200 ;
        RECT 203.800 175.100 204.200 175.200 ;
        RECT 215.000 175.100 215.400 175.200 ;
        RECT 196.600 174.800 204.200 175.100 ;
        RECT 210.200 174.800 215.400 175.100 ;
        RECT 216.600 175.100 217.000 175.200 ;
        RECT 225.400 175.100 225.800 175.200 ;
        RECT 216.600 174.800 225.800 175.100 ;
        RECT 235.000 174.800 235.400 175.200 ;
        RECT 247.800 174.800 248.200 175.200 ;
        RECT 250.200 174.800 250.600 175.200 ;
        RECT 36.600 174.200 36.900 174.800 ;
        RECT 43.800 174.200 44.100 174.800 ;
        RECT 63.800 174.200 64.100 174.800 ;
        RECT 78.200 174.200 78.500 174.800 ;
        RECT 110.200 174.700 110.600 174.800 ;
        RECT 210.200 174.200 210.500 174.800 ;
        RECT 235.000 174.200 235.300 174.800 ;
        RECT 247.800 174.200 248.100 174.800 ;
        RECT 10.200 174.100 10.600 174.200 ;
        RECT 14.200 174.100 14.600 174.200 ;
        RECT 22.200 174.100 22.600 174.200 ;
        RECT 26.200 174.100 26.600 174.200 ;
        RECT 10.200 173.800 14.600 174.100 ;
        RECT 21.400 173.800 26.600 174.100 ;
        RECT 36.600 173.800 37.000 174.200 ;
        RECT 43.800 173.800 44.200 174.200 ;
        RECT 54.200 173.800 56.900 174.100 ;
        RECT 63.800 173.800 64.200 174.200 ;
        RECT 78.200 173.800 78.600 174.200 ;
        RECT 79.000 174.100 79.400 174.200 ;
        RECT 97.400 174.100 97.800 174.200 ;
        RECT 79.000 173.800 97.800 174.100 ;
        RECT 102.200 174.100 102.600 174.200 ;
        RECT 103.800 174.100 104.200 174.200 ;
        RECT 123.000 174.100 123.400 174.200 ;
        RECT 102.200 173.800 123.400 174.100 ;
        RECT 127.800 174.100 128.200 174.200 ;
        RECT 130.200 174.100 130.600 174.200 ;
        RECT 127.800 173.800 130.600 174.100 ;
        RECT 131.800 173.800 132.200 174.200 ;
        RECT 137.400 174.100 137.800 174.200 ;
        RECT 143.800 174.100 144.200 174.200 ;
        RECT 137.400 173.800 144.200 174.100 ;
        RECT 148.600 174.100 149.000 174.200 ;
        RECT 155.800 174.100 156.200 174.200 ;
        RECT 148.600 173.800 156.200 174.100 ;
        RECT 170.200 174.100 170.600 174.200 ;
        RECT 171.000 174.100 171.400 174.200 ;
        RECT 170.200 173.800 171.400 174.100 ;
        RECT 195.800 174.100 196.200 174.200 ;
        RECT 198.200 174.100 198.600 174.200 ;
        RECT 195.800 173.800 198.600 174.100 ;
        RECT 200.600 174.100 201.000 174.200 ;
        RECT 203.800 174.100 204.200 174.200 ;
        RECT 200.600 173.800 204.200 174.100 ;
        RECT 204.600 174.100 205.000 174.200 ;
        RECT 206.200 174.100 206.600 174.200 ;
        RECT 204.600 173.800 206.600 174.100 ;
        RECT 210.200 173.800 210.600 174.200 ;
        RECT 211.000 174.100 211.400 174.200 ;
        RECT 226.200 174.100 226.600 174.200 ;
        RECT 211.000 173.800 226.600 174.100 ;
        RECT 235.000 173.800 235.400 174.200 ;
        RECT 247.800 173.800 248.200 174.200 ;
        RECT 54.200 173.200 54.500 173.800 ;
        RECT 56.600 173.200 56.900 173.800 ;
        RECT 131.800 173.200 132.100 173.800 ;
        RECT 12.600 173.100 13.000 173.200 ;
        RECT 18.200 173.100 18.600 173.200 ;
        RECT 20.600 173.100 21.000 173.200 ;
        RECT 35.000 173.100 35.400 173.200 ;
        RECT 12.600 172.800 35.400 173.100 ;
        RECT 54.200 172.800 54.600 173.200 ;
        RECT 56.600 172.800 57.000 173.200 ;
        RECT 77.400 173.100 77.800 173.200 ;
        RECT 88.600 173.100 89.000 173.200 ;
        RECT 77.400 172.800 89.000 173.100 ;
        RECT 94.200 173.100 94.600 173.200 ;
        RECT 98.200 173.100 98.600 173.200 ;
        RECT 94.200 172.800 98.600 173.100 ;
        RECT 131.000 172.800 131.400 173.200 ;
        RECT 131.800 172.800 132.200 173.200 ;
        RECT 142.200 173.100 142.600 173.200 ;
        RECT 165.400 173.100 165.800 173.200 ;
        RECT 142.200 172.800 165.800 173.100 ;
        RECT 167.000 173.100 167.400 173.200 ;
        RECT 169.400 173.100 169.800 173.200 ;
        RECT 167.000 172.800 169.800 173.100 ;
        RECT 207.800 173.100 208.200 173.200 ;
        RECT 221.400 173.100 221.800 173.200 ;
        RECT 207.800 172.800 221.800 173.100 ;
        RECT 224.600 173.100 225.000 173.200 ;
        RECT 228.600 173.100 229.000 173.200 ;
        RECT 224.600 172.800 229.000 173.100 ;
        RECT 247.800 173.100 248.200 173.200 ;
        RECT 249.400 173.100 249.800 173.200 ;
        RECT 247.800 172.800 249.800 173.100 ;
        RECT 131.000 172.200 131.300 172.800 ;
        RECT 59.800 172.100 60.200 172.200 ;
        RECT 60.600 172.100 61.000 172.200 ;
        RECT 63.000 172.100 63.400 172.200 ;
        RECT 59.800 171.800 63.400 172.100 ;
        RECT 68.600 172.100 69.000 172.200 ;
        RECT 79.000 172.100 79.400 172.200 ;
        RECT 68.600 171.800 79.400 172.100 ;
        RECT 83.800 172.100 84.200 172.200 ;
        RECT 87.000 172.100 87.400 172.200 ;
        RECT 83.800 171.800 87.400 172.100 ;
        RECT 97.400 172.100 97.800 172.200 ;
        RECT 123.800 172.100 124.200 172.200 ;
        RECT 97.400 171.800 124.200 172.100 ;
        RECT 131.000 171.800 131.400 172.200 ;
        RECT 139.800 172.100 140.200 172.200 ;
        RECT 133.400 171.800 140.200 172.100 ;
        RECT 209.400 172.100 209.800 172.200 ;
        RECT 211.000 172.100 211.400 172.200 ;
        RECT 209.400 171.800 211.400 172.100 ;
        RECT 227.000 172.100 227.400 172.200 ;
        RECT 239.000 172.100 239.400 172.200 ;
        RECT 240.600 172.100 241.000 172.200 ;
        RECT 227.000 171.800 241.000 172.100 ;
        RECT 23.800 171.100 24.200 171.200 ;
        RECT 37.400 171.100 37.800 171.200 ;
        RECT 23.800 170.800 37.800 171.100 ;
        RECT 51.000 171.100 51.400 171.200 ;
        RECT 84.600 171.100 85.000 171.200 ;
        RECT 51.000 170.800 85.000 171.100 ;
        RECT 103.800 171.100 104.200 171.200 ;
        RECT 114.200 171.100 114.600 171.200 ;
        RECT 119.000 171.100 119.400 171.200 ;
        RECT 123.000 171.100 123.400 171.200 ;
        RECT 129.400 171.100 129.800 171.200 ;
        RECT 133.400 171.100 133.700 171.800 ;
        RECT 103.800 170.800 129.800 171.100 ;
        RECT 131.800 170.800 133.700 171.100 ;
        RECT 134.200 171.100 134.600 171.200 ;
        RECT 147.800 171.100 148.200 171.200 ;
        RECT 192.600 171.100 193.000 171.200 ;
        RECT 134.200 170.800 193.000 171.100 ;
        RECT 208.600 171.100 209.000 171.200 ;
        RECT 211.800 171.100 212.200 171.200 ;
        RECT 208.600 170.800 212.200 171.100 ;
        RECT 236.600 171.100 237.000 171.200 ;
        RECT 246.200 171.100 246.600 171.200 ;
        RECT 236.600 170.800 246.600 171.100 ;
        RECT 52.600 170.100 53.000 170.200 ;
        RECT 70.200 170.100 70.600 170.200 ;
        RECT 52.600 169.800 70.600 170.100 ;
        RECT 87.000 170.100 87.400 170.200 ;
        RECT 95.000 170.100 95.400 170.200 ;
        RECT 87.000 169.800 95.400 170.100 ;
        RECT 102.200 170.100 102.600 170.200 ;
        RECT 103.800 170.100 104.200 170.200 ;
        RECT 102.200 169.800 104.200 170.100 ;
        RECT 122.200 170.100 122.600 170.200 ;
        RECT 131.800 170.100 132.100 170.800 ;
        RECT 122.200 169.800 132.100 170.100 ;
        RECT 132.600 169.800 133.000 170.200 ;
        RECT 165.400 170.100 165.800 170.200 ;
        RECT 172.600 170.100 173.000 170.200 ;
        RECT 187.000 170.100 187.400 170.200 ;
        RECT 165.400 169.800 187.400 170.100 ;
        RECT 192.600 170.100 193.000 170.200 ;
        RECT 195.000 170.100 195.400 170.200 ;
        RECT 192.600 169.800 195.400 170.100 ;
        RECT 237.400 170.100 237.800 170.200 ;
        RECT 243.800 170.100 244.200 170.200 ;
        RECT 248.600 170.100 249.000 170.200 ;
        RECT 237.400 169.800 249.000 170.100 ;
        RECT 11.800 169.100 12.200 169.200 ;
        RECT 20.600 169.100 21.000 169.200 ;
        RECT 11.800 168.800 21.000 169.100 ;
        RECT 23.000 168.800 23.400 169.200 ;
        RECT 35.000 169.100 35.400 169.200 ;
        RECT 45.400 169.100 45.800 169.200 ;
        RECT 35.000 168.800 45.800 169.100 ;
        RECT 55.800 168.800 56.200 169.200 ;
        RECT 63.000 169.100 63.400 169.200 ;
        RECT 67.800 169.100 68.200 169.200 ;
        RECT 73.400 169.100 73.800 169.200 ;
        RECT 63.000 168.800 73.800 169.100 ;
        RECT 95.800 169.100 96.200 169.200 ;
        RECT 108.600 169.100 109.000 169.200 ;
        RECT 119.000 169.100 119.400 169.200 ;
        RECT 95.800 168.800 109.000 169.100 ;
        RECT 113.400 168.800 119.400 169.100 ;
        RECT 124.600 169.100 125.000 169.200 ;
        RECT 132.600 169.100 132.900 169.800 ;
        RECT 124.600 168.800 132.900 169.100 ;
        RECT 164.600 169.100 165.000 169.200 ;
        RECT 178.200 169.100 178.600 169.200 ;
        RECT 164.600 168.800 178.600 169.100 ;
        RECT 182.200 169.100 182.600 169.200 ;
        RECT 205.400 169.100 205.800 169.200 ;
        RECT 182.200 168.800 205.800 169.100 ;
        RECT 231.800 169.100 232.200 169.200 ;
        RECT 235.000 169.100 235.400 169.200 ;
        RECT 235.800 169.100 236.200 169.200 ;
        RECT 231.800 168.800 236.200 169.100 ;
        RECT 247.000 168.800 247.400 169.200 ;
        RECT 23.000 168.100 23.300 168.800 ;
        RECT 24.600 168.100 25.000 168.200 ;
        RECT 23.000 167.800 25.000 168.100 ;
        RECT 30.200 168.100 30.600 168.200 ;
        RECT 35.800 168.100 36.200 168.200 ;
        RECT 30.200 167.800 36.200 168.100 ;
        RECT 41.400 168.100 41.800 168.200 ;
        RECT 55.800 168.100 56.100 168.800 ;
        RECT 113.400 168.200 113.700 168.800 ;
        RECT 41.400 167.800 56.100 168.100 ;
        RECT 63.800 168.100 64.200 168.200 ;
        RECT 75.800 168.100 76.200 168.200 ;
        RECT 78.200 168.100 78.600 168.200 ;
        RECT 63.800 167.800 78.600 168.100 ;
        RECT 87.800 168.100 88.200 168.200 ;
        RECT 97.400 168.100 97.800 168.200 ;
        RECT 100.600 168.100 101.000 168.200 ;
        RECT 87.800 167.800 101.000 168.100 ;
        RECT 113.400 167.800 113.800 168.200 ;
        RECT 128.600 168.100 129.000 168.200 ;
        RECT 131.000 168.100 131.400 168.200 ;
        RECT 128.600 167.800 131.400 168.100 ;
        RECT 142.200 167.800 142.600 168.200 ;
        RECT 174.200 168.100 174.600 168.200 ;
        RECT 183.000 168.100 183.400 168.200 ;
        RECT 174.200 167.800 183.400 168.100 ;
        RECT 187.000 168.100 187.400 168.200 ;
        RECT 192.600 168.100 193.000 168.200 ;
        RECT 187.000 167.800 193.000 168.100 ;
        RECT 193.400 168.100 193.800 168.200 ;
        RECT 207.000 168.100 207.400 168.200 ;
        RECT 193.400 167.800 207.400 168.100 ;
        RECT 215.000 168.100 215.400 168.200 ;
        RECT 221.400 168.100 221.800 168.200 ;
        RECT 215.000 167.800 221.800 168.100 ;
        RECT 240.600 168.100 241.000 168.200 ;
        RECT 247.000 168.100 247.300 168.800 ;
        RECT 240.600 167.800 247.300 168.100 ;
        RECT 15.000 167.100 15.400 167.200 ;
        RECT 19.000 167.100 19.400 167.200 ;
        RECT 15.000 166.800 19.400 167.100 ;
        RECT 25.400 167.100 25.800 167.200 ;
        RECT 31.800 167.100 32.200 167.200 ;
        RECT 25.400 166.800 32.200 167.100 ;
        RECT 33.400 167.100 33.800 167.200 ;
        RECT 39.000 167.100 39.400 167.200 ;
        RECT 40.600 167.100 41.000 167.200 ;
        RECT 33.400 166.800 41.000 167.100 ;
        RECT 45.400 167.100 45.800 167.200 ;
        RECT 49.400 167.100 49.800 167.200 ;
        RECT 45.400 166.800 49.800 167.100 ;
        RECT 51.800 167.100 52.200 167.200 ;
        RECT 85.400 167.100 85.800 167.200 ;
        RECT 51.800 166.800 85.800 167.100 ;
        RECT 92.600 167.100 93.000 167.200 ;
        RECT 94.200 167.100 94.600 167.200 ;
        RECT 123.800 167.100 124.200 167.200 ;
        RECT 92.600 166.800 124.200 167.100 ;
        RECT 129.400 167.100 129.800 167.200 ;
        RECT 142.200 167.100 142.500 167.800 ;
        RECT 129.400 166.800 142.500 167.100 ;
        RECT 167.800 167.100 168.200 167.200 ;
        RECT 168.600 167.100 169.000 167.200 ;
        RECT 167.800 166.800 169.000 167.100 ;
        RECT 171.000 167.100 171.400 167.200 ;
        RECT 222.200 167.100 222.600 167.200 ;
        RECT 237.400 167.100 237.800 167.200 ;
        RECT 171.000 166.800 222.600 167.100 ;
        RECT 225.400 166.800 237.800 167.100 ;
        RECT 225.400 166.200 225.700 166.800 ;
        RECT 11.800 166.100 12.200 166.200 ;
        RECT 17.400 166.100 17.800 166.200 ;
        RECT 11.800 165.800 17.800 166.100 ;
        RECT 19.000 166.100 19.400 166.200 ;
        RECT 19.800 166.100 20.200 166.200 ;
        RECT 19.000 165.800 20.200 166.100 ;
        RECT 35.000 166.100 35.400 166.200 ;
        RECT 64.600 166.100 65.000 166.200 ;
        RECT 66.200 166.100 66.600 166.200 ;
        RECT 35.000 165.800 47.300 166.100 ;
        RECT 64.600 165.800 66.600 166.100 ;
        RECT 69.400 166.100 69.800 166.200 ;
        RECT 70.200 166.100 70.600 166.200 ;
        RECT 69.400 165.800 70.600 166.100 ;
        RECT 71.000 166.100 71.400 166.200 ;
        RECT 74.200 166.100 74.600 166.200 ;
        RECT 79.800 166.100 80.200 166.200 ;
        RECT 71.000 165.800 80.200 166.100 ;
        RECT 93.400 166.100 93.800 166.200 ;
        RECT 101.400 166.100 101.800 166.200 ;
        RECT 93.400 165.800 101.800 166.100 ;
        RECT 108.600 166.100 109.000 166.200 ;
        RECT 116.600 166.100 117.000 166.200 ;
        RECT 108.600 165.800 117.000 166.100 ;
        RECT 122.200 166.100 122.600 166.200 ;
        RECT 124.600 166.100 125.000 166.200 ;
        RECT 122.200 165.800 125.000 166.100 ;
        RECT 126.200 166.100 126.600 166.200 ;
        RECT 127.800 166.100 128.200 166.200 ;
        RECT 126.200 165.800 128.200 166.100 ;
        RECT 144.600 166.100 145.000 166.200 ;
        RECT 149.400 166.100 149.800 166.200 ;
        RECT 144.600 165.800 149.800 166.100 ;
        RECT 155.800 165.800 156.200 166.200 ;
        RECT 159.800 166.100 160.200 166.200 ;
        RECT 160.600 166.100 161.000 166.200 ;
        RECT 159.800 165.800 161.000 166.100 ;
        RECT 170.200 166.100 170.600 166.200 ;
        RECT 173.400 166.100 173.800 166.200 ;
        RECT 175.000 166.100 175.400 166.200 ;
        RECT 177.400 166.100 177.800 166.200 ;
        RECT 170.200 165.800 174.500 166.100 ;
        RECT 175.000 165.800 177.800 166.100 ;
        RECT 179.800 166.100 180.200 166.200 ;
        RECT 192.600 166.100 193.000 166.200 ;
        RECT 195.800 166.100 196.200 166.200 ;
        RECT 179.800 165.800 196.200 166.100 ;
        RECT 206.200 166.100 206.600 166.200 ;
        RECT 208.600 166.100 209.000 166.200 ;
        RECT 206.200 165.800 209.000 166.100 ;
        RECT 209.400 166.100 209.800 166.200 ;
        RECT 211.800 166.100 212.200 166.200 ;
        RECT 217.400 166.100 217.800 166.200 ;
        RECT 209.400 165.800 217.800 166.100 ;
        RECT 218.200 166.100 218.600 166.200 ;
        RECT 225.400 166.100 225.800 166.200 ;
        RECT 218.200 165.800 225.800 166.100 ;
        RECT 47.000 165.200 47.300 165.800 ;
        RECT 155.800 165.200 156.100 165.800 ;
        RECT 4.600 165.100 5.000 165.200 ;
        RECT 31.800 165.100 32.200 165.200 ;
        RECT 34.200 165.100 34.600 165.200 ;
        RECT 4.600 164.800 34.600 165.100 ;
        RECT 42.200 165.100 42.600 165.200 ;
        RECT 43.000 165.100 43.400 165.200 ;
        RECT 44.600 165.100 45.000 165.200 ;
        RECT 42.200 164.800 45.000 165.100 ;
        RECT 47.000 164.800 47.400 165.200 ;
        RECT 56.600 165.100 57.000 165.200 ;
        RECT 79.000 165.100 79.400 165.200 ;
        RECT 81.400 165.100 81.800 165.200 ;
        RECT 56.600 164.800 64.100 165.100 ;
        RECT 79.000 164.800 81.800 165.100 ;
        RECT 83.800 165.100 84.200 165.200 ;
        RECT 84.600 165.100 85.000 165.200 ;
        RECT 83.800 164.800 85.000 165.100 ;
        RECT 95.800 165.100 96.200 165.200 ;
        RECT 118.200 165.100 118.600 165.200 ;
        RECT 138.200 165.100 138.600 165.200 ;
        RECT 95.800 164.800 118.600 165.100 ;
        RECT 128.600 164.800 138.600 165.100 ;
        RECT 142.200 165.100 142.600 165.200 ;
        RECT 155.000 165.100 155.400 165.200 ;
        RECT 142.200 164.800 155.400 165.100 ;
        RECT 155.800 164.800 156.200 165.200 ;
        RECT 160.600 165.100 161.000 165.200 ;
        RECT 161.400 165.100 161.800 165.200 ;
        RECT 160.600 164.800 161.800 165.100 ;
        RECT 162.200 164.800 162.600 165.200 ;
        RECT 165.400 165.100 165.800 165.200 ;
        RECT 167.800 165.100 168.200 165.200 ;
        RECT 165.400 164.800 168.200 165.100 ;
        RECT 175.000 165.100 175.400 165.200 ;
        RECT 175.800 165.100 176.200 165.200 ;
        RECT 175.000 164.800 176.200 165.100 ;
        RECT 176.600 165.100 177.000 165.200 ;
        RECT 187.000 165.100 187.400 165.200 ;
        RECT 176.600 164.800 187.400 165.100 ;
        RECT 211.000 164.800 211.400 165.200 ;
        RECT 213.400 165.100 213.800 165.200 ;
        RECT 215.800 165.100 216.200 165.200 ;
        RECT 213.400 164.800 216.200 165.100 ;
        RECT 63.800 164.200 64.100 164.800 ;
        RECT 128.600 164.200 128.900 164.800 ;
        RECT 18.200 164.100 18.600 164.200 ;
        RECT 37.400 164.100 37.800 164.200 ;
        RECT 43.800 164.100 44.200 164.200 ;
        RECT 18.200 163.800 19.300 164.100 ;
        RECT 37.400 163.800 44.200 164.100 ;
        RECT 44.600 164.100 45.000 164.200 ;
        RECT 46.200 164.100 46.600 164.200 ;
        RECT 44.600 163.800 46.600 164.100 ;
        RECT 51.000 164.100 51.400 164.200 ;
        RECT 58.200 164.100 58.600 164.200 ;
        RECT 51.000 163.800 58.600 164.100 ;
        RECT 63.800 163.800 64.200 164.200 ;
        RECT 84.600 163.800 85.000 164.200 ;
        RECT 87.800 164.100 88.200 164.200 ;
        RECT 89.400 164.100 89.800 164.200 ;
        RECT 99.000 164.100 99.400 164.200 ;
        RECT 103.000 164.100 103.400 164.200 ;
        RECT 116.600 164.100 117.000 164.200 ;
        RECT 87.800 163.800 117.000 164.100 ;
        RECT 128.600 163.800 129.000 164.200 ;
        RECT 162.200 164.100 162.500 164.800 ;
        RECT 211.000 164.200 211.300 164.800 ;
        RECT 180.600 164.100 181.000 164.200 ;
        RECT 162.200 163.800 181.000 164.100 ;
        RECT 184.600 164.100 185.000 164.200 ;
        RECT 204.600 164.100 205.000 164.200 ;
        RECT 184.600 163.800 205.000 164.100 ;
        RECT 211.000 163.800 211.400 164.200 ;
        RECT 19.000 163.200 19.300 163.800 ;
        RECT 19.000 162.800 19.400 163.200 ;
        RECT 36.600 163.100 37.000 163.200 ;
        RECT 51.800 163.100 52.200 163.200 ;
        RECT 36.600 162.800 52.200 163.100 ;
        RECT 84.600 163.100 84.900 163.800 ;
        RECT 130.200 163.100 130.600 163.200 ;
        RECT 84.600 162.800 130.600 163.100 ;
        RECT 131.000 163.100 131.400 163.200 ;
        RECT 143.000 163.100 143.400 163.200 ;
        RECT 195.800 163.100 196.200 163.200 ;
        RECT 131.000 162.800 196.200 163.100 ;
        RECT 39.000 162.100 39.400 162.200 ;
        RECT 47.800 162.100 48.200 162.200 ;
        RECT 39.000 161.800 48.200 162.100 ;
        RECT 51.800 162.100 52.200 162.200 ;
        RECT 54.200 162.100 54.600 162.200 ;
        RECT 58.200 162.100 58.600 162.200 ;
        RECT 51.800 161.800 58.600 162.100 ;
        RECT 123.800 162.100 124.200 162.200 ;
        RECT 154.200 162.100 154.600 162.200 ;
        RECT 123.800 161.800 154.600 162.100 ;
        RECT 159.800 162.100 160.200 162.200 ;
        RECT 171.800 162.100 172.200 162.200 ;
        RECT 159.800 161.800 172.200 162.100 ;
        RECT 236.600 162.100 237.000 162.200 ;
        RECT 237.400 162.100 237.800 162.200 ;
        RECT 236.600 161.800 237.800 162.100 ;
        RECT 39.800 160.800 40.200 161.200 ;
        RECT 66.200 161.100 66.600 161.200 ;
        RECT 87.800 161.100 88.200 161.200 ;
        RECT 114.200 161.100 114.600 161.200 ;
        RECT 117.400 161.100 117.800 161.200 ;
        RECT 66.200 160.800 117.800 161.100 ;
        RECT 152.600 161.100 153.000 161.200 ;
        RECT 157.400 161.100 157.800 161.200 ;
        RECT 152.600 160.800 157.800 161.100 ;
        RECT 172.600 161.100 173.000 161.200 ;
        RECT 198.200 161.100 198.600 161.200 ;
        RECT 172.600 160.800 198.600 161.100 ;
        RECT 242.200 161.100 242.600 161.200 ;
        RECT 244.600 161.100 245.000 161.200 ;
        RECT 242.200 160.800 245.000 161.100 ;
        RECT 39.800 160.200 40.100 160.800 ;
        RECT 39.800 159.800 40.200 160.200 ;
        RECT 64.600 160.100 65.000 160.200 ;
        RECT 71.800 160.100 72.200 160.200 ;
        RECT 112.600 160.100 113.000 160.200 ;
        RECT 132.600 160.100 133.000 160.200 ;
        RECT 64.600 159.800 133.000 160.100 ;
        RECT 198.200 160.100 198.600 160.200 ;
        RECT 216.600 160.100 217.000 160.200 ;
        RECT 198.200 159.800 217.000 160.100 ;
        RECT 27.800 158.800 28.200 159.200 ;
        RECT 76.600 159.100 77.000 159.200 ;
        RECT 79.000 159.100 79.400 159.200 ;
        RECT 76.600 158.800 79.400 159.100 ;
        RECT 117.400 159.100 117.800 159.200 ;
        RECT 129.400 159.100 129.800 159.200 ;
        RECT 117.400 158.800 129.800 159.100 ;
        RECT 132.600 159.100 133.000 159.200 ;
        RECT 133.400 159.100 133.800 159.200 ;
        RECT 132.600 158.800 133.800 159.100 ;
        RECT 135.800 159.100 136.200 159.200 ;
        RECT 184.600 159.100 185.000 159.200 ;
        RECT 135.800 158.800 185.000 159.100 ;
        RECT 201.400 159.100 201.800 159.200 ;
        RECT 204.600 159.100 205.000 159.200 ;
        RECT 214.200 159.100 214.600 159.200 ;
        RECT 201.400 158.800 214.600 159.100 ;
        RECT 27.800 158.200 28.100 158.800 ;
        RECT 27.800 157.800 28.200 158.200 ;
        RECT 43.000 158.100 43.400 158.200 ;
        RECT 68.600 158.100 69.000 158.200 ;
        RECT 43.000 157.800 69.000 158.100 ;
        RECT 81.400 157.800 81.800 158.200 ;
        RECT 118.200 158.100 118.600 158.200 ;
        RECT 189.400 158.100 189.800 158.200 ;
        RECT 207.000 158.100 207.400 158.200 ;
        RECT 118.200 157.800 154.500 158.100 ;
        RECT 189.400 157.800 207.400 158.100 ;
        RECT 209.400 158.100 209.800 158.200 ;
        RECT 213.400 158.100 213.800 158.200 ;
        RECT 209.400 157.800 213.800 158.100 ;
        RECT 216.600 158.100 217.000 158.200 ;
        RECT 246.200 158.100 246.600 158.200 ;
        RECT 216.600 157.800 246.600 158.100 ;
        RECT 81.400 157.200 81.700 157.800 ;
        RECT 45.400 157.100 45.800 157.200 ;
        RECT 52.600 157.100 53.000 157.200 ;
        RECT 45.400 156.800 53.000 157.100 ;
        RECT 59.800 157.100 60.200 157.200 ;
        RECT 66.200 157.100 66.600 157.200 ;
        RECT 59.800 156.800 66.600 157.100 ;
        RECT 81.400 156.800 81.800 157.200 ;
        RECT 103.000 157.100 103.400 157.200 ;
        RECT 126.200 157.100 126.600 157.200 ;
        RECT 103.000 156.800 126.600 157.100 ;
        RECT 154.200 157.100 154.500 157.800 ;
        RECT 171.800 157.100 172.200 157.200 ;
        RECT 173.400 157.100 173.800 157.200 ;
        RECT 175.800 157.100 176.200 157.200 ;
        RECT 206.200 157.100 206.600 157.200 ;
        RECT 154.200 156.800 176.200 157.100 ;
        RECT 192.600 156.800 206.600 157.100 ;
        RECT 216.600 157.100 217.000 157.200 ;
        RECT 231.800 157.100 232.200 157.200 ;
        RECT 249.400 157.100 249.800 157.200 ;
        RECT 216.600 156.800 249.800 157.100 ;
        RECT 192.600 156.200 192.900 156.800 ;
        RECT 10.200 156.100 10.600 156.200 ;
        RECT 11.000 156.100 11.400 156.200 ;
        RECT 14.200 156.100 14.600 156.200 ;
        RECT 10.200 155.800 14.600 156.100 ;
        RECT 19.800 156.100 20.200 156.200 ;
        RECT 29.400 156.100 29.800 156.200 ;
        RECT 65.400 156.100 65.800 156.200 ;
        RECT 67.000 156.100 67.400 156.200 ;
        RECT 19.800 155.800 64.100 156.100 ;
        RECT 65.400 155.800 67.400 156.100 ;
        RECT 67.800 156.100 68.200 156.200 ;
        RECT 75.800 156.100 76.200 156.200 ;
        RECT 67.800 155.800 76.200 156.100 ;
        RECT 78.200 156.100 78.600 156.200 ;
        RECT 87.000 156.100 87.400 156.200 ;
        RECT 78.200 155.800 87.400 156.100 ;
        RECT 114.200 156.100 114.600 156.200 ;
        RECT 124.600 156.100 125.000 156.200 ;
        RECT 127.800 156.100 128.200 156.200 ;
        RECT 114.200 155.800 128.200 156.100 ;
        RECT 130.200 155.800 130.600 156.200 ;
        RECT 142.200 156.100 142.600 156.200 ;
        RECT 143.800 156.100 144.200 156.200 ;
        RECT 144.600 156.100 145.000 156.200 ;
        RECT 142.200 155.800 145.000 156.100 ;
        RECT 147.800 156.100 148.200 156.200 ;
        RECT 148.600 156.100 149.000 156.200 ;
        RECT 147.800 155.800 149.000 156.100 ;
        RECT 155.800 156.100 156.200 156.200 ;
        RECT 159.000 156.100 159.400 156.200 ;
        RECT 160.600 156.100 161.000 156.200 ;
        RECT 155.800 155.800 161.000 156.100 ;
        RECT 163.800 155.800 164.200 156.200 ;
        RECT 175.000 156.100 175.400 156.200 ;
        RECT 182.200 156.100 182.600 156.200 ;
        RECT 192.600 156.100 193.000 156.200 ;
        RECT 175.000 155.800 181.700 156.100 ;
        RECT 182.200 155.800 193.000 156.100 ;
        RECT 195.800 156.100 196.200 156.200 ;
        RECT 202.200 156.100 202.600 156.200 ;
        RECT 220.600 156.100 221.000 156.200 ;
        RECT 195.800 155.800 197.700 156.100 ;
        RECT 202.200 155.800 221.000 156.100 ;
        RECT 232.600 156.100 233.000 156.200 ;
        RECT 234.200 156.100 234.600 156.200 ;
        RECT 232.600 155.800 234.600 156.100 ;
        RECT 5.400 155.100 5.800 155.200 ;
        RECT 12.600 155.100 13.000 155.200 ;
        RECT 5.400 154.800 13.000 155.100 ;
        RECT 16.600 155.100 17.000 155.200 ;
        RECT 18.200 155.100 18.600 155.200 ;
        RECT 16.600 154.800 18.600 155.100 ;
        RECT 20.600 154.800 21.000 155.200 ;
        RECT 22.200 155.100 22.600 155.200 ;
        RECT 23.800 155.100 24.200 155.200 ;
        RECT 22.200 154.800 24.200 155.100 ;
        RECT 35.800 155.100 36.200 155.200 ;
        RECT 36.600 155.100 37.000 155.200 ;
        RECT 35.800 154.800 37.000 155.100 ;
        RECT 38.200 155.100 38.600 155.200 ;
        RECT 47.800 155.100 48.200 155.200 ;
        RECT 48.600 155.100 49.000 155.200 ;
        RECT 38.200 154.800 46.500 155.100 ;
        RECT 47.800 154.800 49.000 155.100 ;
        RECT 63.000 154.800 63.400 155.200 ;
        RECT 63.800 155.100 64.100 155.800 ;
        RECT 77.400 155.100 77.800 155.200 ;
        RECT 63.800 154.800 77.800 155.100 ;
        RECT 79.000 155.100 79.400 155.200 ;
        RECT 81.400 155.100 81.800 155.200 ;
        RECT 79.000 154.800 81.800 155.100 ;
        RECT 93.400 155.100 93.800 155.200 ;
        RECT 99.800 155.100 100.200 155.200 ;
        RECT 105.400 155.100 105.800 155.200 ;
        RECT 93.400 154.800 105.800 155.100 ;
        RECT 111.800 155.100 112.200 155.200 ;
        RECT 115.000 155.100 115.400 155.200 ;
        RECT 111.800 154.800 115.400 155.100 ;
        RECT 118.200 155.100 118.600 155.200 ;
        RECT 123.800 155.100 124.200 155.200 ;
        RECT 130.200 155.100 130.500 155.800 ;
        RECT 163.800 155.200 164.100 155.800 ;
        RECT 118.200 154.800 123.300 155.100 ;
        RECT 123.800 154.800 130.500 155.100 ;
        RECT 133.400 155.100 133.800 155.200 ;
        RECT 145.400 155.100 145.800 155.200 ;
        RECT 133.400 154.800 145.800 155.100 ;
        RECT 163.800 154.800 164.200 155.200 ;
        RECT 167.000 155.100 167.400 155.200 ;
        RECT 177.400 155.100 177.800 155.200 ;
        RECT 167.000 154.800 177.800 155.100 ;
        RECT 181.400 155.100 181.700 155.800 ;
        RECT 187.800 155.100 188.200 155.200 ;
        RECT 181.400 154.800 188.200 155.100 ;
        RECT 194.200 155.100 194.600 155.200 ;
        RECT 196.600 155.100 197.000 155.200 ;
        RECT 194.200 154.800 197.000 155.100 ;
        RECT 197.400 155.100 197.700 155.800 ;
        RECT 209.400 155.100 209.800 155.200 ;
        RECT 197.400 154.800 209.800 155.100 ;
        RECT 213.400 155.100 213.800 155.200 ;
        RECT 223.000 155.100 223.400 155.200 ;
        RECT 227.800 155.100 228.200 155.200 ;
        RECT 213.400 154.800 228.200 155.100 ;
        RECT 235.000 155.100 235.400 155.200 ;
        RECT 247.800 155.100 248.200 155.200 ;
        RECT 248.600 155.100 249.000 155.200 ;
        RECT 235.000 154.800 243.300 155.100 ;
        RECT 247.800 154.800 249.000 155.100 ;
        RECT 20.600 154.200 20.900 154.800 ;
        RECT 46.200 154.200 46.500 154.800 ;
        RECT 11.000 154.100 11.400 154.200 ;
        RECT 15.800 154.100 16.200 154.200 ;
        RECT 11.000 153.800 16.200 154.100 ;
        RECT 20.600 153.800 21.000 154.200 ;
        RECT 26.200 154.100 26.600 154.200 ;
        RECT 42.200 154.100 42.600 154.200 ;
        RECT 26.200 153.800 42.600 154.100 ;
        RECT 46.200 153.800 46.600 154.200 ;
        RECT 54.200 154.100 54.600 154.200 ;
        RECT 63.000 154.100 63.300 154.800 ;
        RECT 54.200 153.800 63.300 154.100 ;
        RECT 68.600 154.100 69.000 154.200 ;
        RECT 84.600 154.100 85.000 154.200 ;
        RECT 68.600 153.800 85.000 154.100 ;
        RECT 85.400 154.100 85.800 154.200 ;
        RECT 94.200 154.100 94.600 154.200 ;
        RECT 96.600 154.100 97.000 154.200 ;
        RECT 85.400 153.800 97.000 154.100 ;
        RECT 102.200 154.100 102.600 154.200 ;
        RECT 103.800 154.100 104.200 154.200 ;
        RECT 105.400 154.100 105.800 154.200 ;
        RECT 102.200 153.800 105.800 154.100 ;
        RECT 107.800 154.100 108.200 154.200 ;
        RECT 109.400 154.100 109.800 154.200 ;
        RECT 122.200 154.100 122.600 154.200 ;
        RECT 107.800 153.800 122.600 154.100 ;
        RECT 123.000 154.100 123.300 154.800 ;
        RECT 243.000 154.200 243.300 154.800 ;
        RECT 126.200 154.100 126.600 154.200 ;
        RECT 123.000 153.800 126.600 154.100 ;
        RECT 143.000 154.100 143.400 154.200 ;
        RECT 147.000 154.100 147.400 154.200 ;
        RECT 147.800 154.100 148.200 154.200 ;
        RECT 143.000 153.800 148.200 154.100 ;
        RECT 157.400 154.100 157.800 154.200 ;
        RECT 166.200 154.100 166.600 154.200 ;
        RECT 157.400 153.800 166.600 154.100 ;
        RECT 171.800 154.100 172.200 154.200 ;
        RECT 173.400 154.100 173.800 154.200 ;
        RECT 178.200 154.100 178.600 154.200 ;
        RECT 179.000 154.100 179.400 154.200 ;
        RECT 183.000 154.100 183.400 154.200 ;
        RECT 171.800 153.800 173.800 154.100 ;
        RECT 177.400 153.800 183.400 154.100 ;
        RECT 243.000 153.800 243.400 154.200 ;
        RECT 22.200 153.100 22.600 153.200 ;
        RECT 30.200 153.100 30.600 153.200 ;
        RECT 22.200 152.800 30.600 153.100 ;
        RECT 34.200 153.100 34.600 153.200 ;
        RECT 56.600 153.100 57.000 153.200 ;
        RECT 68.600 153.100 69.000 153.200 ;
        RECT 34.200 152.800 69.000 153.100 ;
        RECT 153.400 153.100 153.800 153.200 ;
        RECT 170.200 153.100 170.600 153.200 ;
        RECT 175.000 153.100 175.400 153.200 ;
        RECT 153.400 152.800 175.400 153.100 ;
        RECT 17.400 152.100 17.800 152.200 ;
        RECT 42.200 152.100 42.600 152.200 ;
        RECT 17.400 151.800 42.600 152.100 ;
        RECT 76.600 152.100 77.000 152.200 ;
        RECT 80.600 152.100 81.000 152.200 ;
        RECT 76.600 151.800 81.000 152.100 ;
        RECT 99.800 152.100 100.200 152.200 ;
        RECT 107.000 152.100 107.400 152.200 ;
        RECT 99.800 151.800 107.400 152.100 ;
        RECT 108.600 152.100 109.000 152.200 ;
        RECT 124.600 152.100 125.000 152.200 ;
        RECT 108.600 151.800 125.000 152.100 ;
        RECT 198.200 152.100 198.600 152.200 ;
        RECT 199.000 152.100 199.400 152.200 ;
        RECT 203.000 152.100 203.400 152.200 ;
        RECT 198.200 151.800 203.400 152.100 ;
        RECT 35.000 151.100 35.400 151.200 ;
        RECT 47.000 151.100 47.400 151.200 ;
        RECT 35.000 150.800 47.400 151.100 ;
        RECT 55.800 151.100 56.200 151.200 ;
        RECT 74.200 151.100 74.600 151.200 ;
        RECT 55.800 150.800 74.600 151.100 ;
        RECT 111.000 151.100 111.400 151.200 ;
        RECT 123.000 151.100 123.400 151.200 ;
        RECT 135.800 151.100 136.200 151.200 ;
        RECT 111.000 150.800 121.700 151.100 ;
        RECT 123.000 150.800 136.200 151.100 ;
        RECT 139.800 151.100 140.200 151.200 ;
        RECT 163.000 151.100 163.400 151.200 ;
        RECT 139.800 150.800 163.400 151.100 ;
        RECT 186.200 151.100 186.600 151.200 ;
        RECT 190.200 151.100 190.600 151.200 ;
        RECT 186.200 150.800 190.600 151.100 ;
        RECT 250.200 150.800 250.600 151.200 ;
        RECT 121.400 150.200 121.700 150.800 ;
        RECT 250.200 150.200 250.500 150.800 ;
        RECT 105.400 150.100 105.800 150.200 ;
        RECT 116.600 150.100 117.000 150.200 ;
        RECT 118.200 150.100 118.600 150.200 ;
        RECT 105.400 149.800 118.600 150.100 ;
        RECT 121.400 150.100 121.800 150.200 ;
        RECT 131.000 150.100 131.400 150.200 ;
        RECT 121.400 149.800 131.400 150.100 ;
        RECT 168.600 150.100 169.000 150.200 ;
        RECT 178.200 150.100 178.600 150.200 ;
        RECT 168.600 149.800 178.600 150.100 ;
        RECT 241.400 150.100 241.800 150.200 ;
        RECT 247.800 150.100 248.200 150.200 ;
        RECT 241.400 149.800 248.200 150.100 ;
        RECT 250.200 149.800 250.600 150.200 ;
        RECT 32.600 149.100 33.000 149.200 ;
        RECT 35.800 149.100 36.200 149.200 ;
        RECT 32.600 148.800 36.200 149.100 ;
        RECT 67.000 149.100 67.400 149.200 ;
        RECT 67.800 149.100 68.200 149.200 ;
        RECT 67.000 148.800 68.200 149.100 ;
        RECT 73.400 148.800 73.800 149.200 ;
        RECT 77.400 149.100 77.800 149.200 ;
        RECT 91.000 149.100 91.400 149.200 ;
        RECT 77.400 148.800 91.400 149.100 ;
        RECT 107.000 149.100 107.400 149.200 ;
        RECT 132.600 149.100 133.000 149.200 ;
        RECT 107.000 148.800 133.000 149.100 ;
        RECT 138.200 149.100 138.600 149.200 ;
        RECT 152.600 149.100 153.000 149.200 ;
        RECT 138.200 148.800 153.000 149.100 ;
        RECT 161.400 149.100 161.800 149.200 ;
        RECT 166.200 149.100 166.600 149.200 ;
        RECT 170.200 149.100 170.600 149.200 ;
        RECT 161.400 148.800 170.600 149.100 ;
        RECT 195.000 149.100 195.400 149.200 ;
        RECT 220.600 149.100 221.000 149.200 ;
        RECT 195.000 148.800 221.000 149.100 ;
        RECT 223.000 149.100 223.400 149.200 ;
        RECT 227.800 149.100 228.200 149.200 ;
        RECT 223.000 148.800 228.200 149.100 ;
        RECT 243.000 149.100 243.400 149.200 ;
        RECT 243.800 149.100 244.200 149.200 ;
        RECT 243.000 148.800 244.200 149.100 ;
        RECT 73.400 148.200 73.700 148.800 ;
        RECT 79.800 148.200 80.100 148.800 ;
        RECT 40.600 148.100 41.000 148.200 ;
        RECT 48.600 148.100 49.000 148.200 ;
        RECT 54.200 148.100 54.600 148.200 ;
        RECT 58.200 148.100 58.600 148.200 ;
        RECT 40.600 147.800 58.600 148.100 ;
        RECT 73.400 147.800 73.800 148.200 ;
        RECT 79.800 147.800 80.200 148.200 ;
        RECT 89.400 148.100 89.800 148.200 ;
        RECT 108.600 148.100 109.000 148.200 ;
        RECT 123.000 148.100 123.400 148.200 ;
        RECT 89.400 147.800 123.400 148.100 ;
        RECT 135.000 148.100 135.400 148.200 ;
        RECT 136.600 148.100 137.000 148.200 ;
        RECT 149.400 148.100 149.800 148.200 ;
        RECT 135.000 147.800 149.800 148.100 ;
        RECT 155.800 148.100 156.200 148.200 ;
        RECT 172.600 148.100 173.000 148.200 ;
        RECT 174.200 148.100 174.600 148.200 ;
        RECT 155.800 147.800 174.600 148.100 ;
        RECT 192.600 148.100 193.000 148.200 ;
        RECT 206.200 148.100 206.600 148.200 ;
        RECT 192.600 147.800 206.600 148.100 ;
        RECT 219.000 148.100 219.400 148.200 ;
        RECT 221.400 148.100 221.800 148.200 ;
        RECT 250.200 148.100 250.600 148.200 ;
        RECT 219.000 147.800 250.600 148.100 ;
        RECT 3.800 147.100 4.200 147.200 ;
        RECT 12.600 147.100 13.000 147.200 ;
        RECT 3.800 146.800 13.000 147.100 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 25.400 147.100 25.800 147.200 ;
        RECT 14.200 146.800 25.800 147.100 ;
        RECT 34.200 147.100 34.600 147.200 ;
        RECT 35.800 147.100 36.200 147.200 ;
        RECT 34.200 146.800 36.200 147.100 ;
        RECT 37.400 146.800 37.800 147.200 ;
        RECT 44.600 147.100 45.000 147.200 ;
        RECT 56.600 147.100 57.000 147.200 ;
        RECT 44.600 146.800 57.000 147.100 ;
        RECT 69.400 147.100 69.800 147.200 ;
        RECT 75.000 147.100 75.400 147.200 ;
        RECT 69.400 146.800 75.400 147.100 ;
        RECT 95.000 147.100 95.400 147.200 ;
        RECT 100.600 147.100 101.000 147.200 ;
        RECT 95.000 146.800 101.000 147.100 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 129.400 147.100 129.800 147.200 ;
        RECT 135.800 147.100 136.200 147.200 ;
        RECT 129.400 146.800 136.200 147.100 ;
        RECT 143.000 147.100 143.400 147.200 ;
        RECT 148.600 147.100 149.000 147.200 ;
        RECT 143.000 146.800 149.000 147.100 ;
        RECT 159.000 147.100 159.400 147.200 ;
        RECT 164.600 147.100 165.000 147.200 ;
        RECT 159.000 146.800 165.000 147.100 ;
        RECT 167.800 147.100 168.200 147.200 ;
        RECT 179.800 147.100 180.200 147.200 ;
        RECT 167.800 146.800 180.200 147.100 ;
        RECT 199.000 147.100 199.400 147.200 ;
        RECT 202.200 147.100 202.600 147.200 ;
        RECT 199.000 146.800 202.600 147.100 ;
        RECT 203.000 147.100 203.400 147.200 ;
        RECT 207.000 147.100 207.400 147.200 ;
        RECT 208.600 147.100 209.000 147.200 ;
        RECT 203.000 146.800 209.000 147.100 ;
        RECT 221.400 147.100 221.800 147.200 ;
        RECT 223.000 147.100 223.400 147.200 ;
        RECT 221.400 146.800 223.400 147.100 ;
        RECT 228.600 147.100 229.000 147.200 ;
        RECT 238.200 147.100 238.600 147.200 ;
        RECT 228.600 146.800 238.600 147.100 ;
        RECT 239.000 146.800 239.400 147.200 ;
        RECT 244.600 146.800 245.000 147.200 ;
        RECT 37.400 146.200 37.700 146.800 ;
        RECT 11.800 146.100 12.200 146.200 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 15.000 146.100 15.400 146.200 ;
        RECT 11.800 145.800 15.400 146.100 ;
        RECT 20.600 146.100 21.000 146.200 ;
        RECT 27.800 146.100 28.200 146.200 ;
        RECT 20.600 145.800 28.200 146.100 ;
        RECT 32.600 146.100 33.000 146.200 ;
        RECT 34.200 146.100 34.600 146.200 ;
        RECT 32.600 145.800 34.600 146.100 ;
        RECT 37.400 145.800 37.800 146.200 ;
        RECT 43.000 146.100 43.400 146.200 ;
        RECT 43.800 146.100 44.200 146.200 ;
        RECT 43.000 145.800 44.200 146.100 ;
        RECT 47.800 146.100 48.200 146.200 ;
        RECT 51.800 146.100 52.200 146.200 ;
        RECT 75.800 146.100 76.200 146.200 ;
        RECT 84.600 146.100 85.000 146.200 ;
        RECT 47.800 145.800 52.200 146.100 ;
        RECT 75.000 145.800 85.000 146.100 ;
        RECT 86.200 146.100 86.600 146.200 ;
        RECT 95.800 146.100 96.200 146.200 ;
        RECT 99.000 146.100 99.400 146.200 ;
        RECT 86.200 145.800 99.400 146.100 ;
        RECT 102.200 146.100 102.600 146.200 ;
        RECT 110.200 146.100 110.500 146.800 ;
        RECT 102.200 145.800 110.500 146.100 ;
        RECT 125.400 146.100 125.800 146.200 ;
        RECT 151.000 146.100 151.400 146.200 ;
        RECT 170.200 146.100 170.600 146.200 ;
        RECT 179.000 146.100 179.400 146.200 ;
        RECT 125.400 145.800 170.600 146.100 ;
        RECT 172.600 145.800 179.400 146.100 ;
        RECT 183.800 146.100 184.200 146.200 ;
        RECT 190.200 146.100 190.600 146.200 ;
        RECT 191.000 146.100 191.400 146.200 ;
        RECT 183.800 145.800 191.400 146.100 ;
        RECT 201.400 146.100 201.800 146.200 ;
        RECT 213.400 146.100 213.800 146.200 ;
        RECT 214.200 146.100 214.600 146.200 ;
        RECT 201.400 145.800 204.900 146.100 ;
        RECT 213.400 145.800 214.600 146.100 ;
        RECT 222.200 145.800 222.600 146.200 ;
        RECT 224.600 146.100 225.000 146.200 ;
        RECT 228.600 146.100 229.000 146.200 ;
        RECT 229.400 146.100 229.800 146.200 ;
        RECT 224.600 145.800 229.800 146.100 ;
        RECT 230.200 146.100 230.600 146.200 ;
        RECT 231.800 146.100 232.200 146.200 ;
        RECT 230.200 145.800 232.200 146.100 ;
        RECT 238.200 146.100 238.600 146.200 ;
        RECT 239.000 146.100 239.300 146.800 ;
        RECT 238.200 145.800 239.300 146.100 ;
        RECT 240.600 146.100 241.000 146.200 ;
        RECT 244.600 146.100 244.900 146.800 ;
        RECT 240.600 145.800 244.900 146.100 ;
        RECT 147.000 145.200 147.300 145.800 ;
        RECT 172.600 145.200 172.900 145.800 ;
        RECT 204.600 145.200 204.900 145.800 ;
        RECT 222.200 145.200 222.500 145.800 ;
        RECT 47.000 145.100 47.400 145.200 ;
        RECT 47.800 145.100 48.200 145.200 ;
        RECT 47.000 144.800 48.200 145.100 ;
        RECT 67.800 145.100 68.200 145.200 ;
        RECT 83.800 145.100 84.200 145.200 ;
        RECT 67.800 144.800 84.200 145.100 ;
        RECT 121.400 145.100 121.800 145.200 ;
        RECT 130.200 145.100 130.600 145.200 ;
        RECT 121.400 144.800 130.600 145.100 ;
        RECT 147.000 144.800 147.400 145.200 ;
        RECT 147.800 145.100 148.200 145.200 ;
        RECT 152.600 145.100 153.000 145.200 ;
        RECT 147.800 144.800 153.000 145.100 ;
        RECT 155.800 145.100 156.200 145.200 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 171.000 145.100 171.400 145.200 ;
        RECT 155.800 144.800 171.400 145.100 ;
        RECT 172.600 144.800 173.000 145.200 ;
        RECT 197.400 145.100 197.800 145.200 ;
        RECT 199.000 145.100 199.400 145.200 ;
        RECT 197.400 144.800 199.400 145.100 ;
        RECT 204.600 144.800 205.000 145.200 ;
        RECT 216.600 145.100 217.000 145.200 ;
        RECT 219.000 145.100 219.400 145.200 ;
        RECT 216.600 144.800 219.400 145.100 ;
        RECT 222.200 144.800 222.600 145.200 ;
        RECT 227.800 145.100 228.200 145.200 ;
        RECT 234.200 145.100 234.600 145.200 ;
        RECT 227.000 144.800 234.600 145.100 ;
        RECT 235.800 145.100 236.200 145.200 ;
        RECT 239.800 145.100 240.200 145.200 ;
        RECT 235.800 144.800 240.200 145.100 ;
        RECT 5.400 144.100 5.800 144.200 ;
        RECT 16.600 144.100 17.000 144.200 ;
        RECT 5.400 143.800 17.000 144.100 ;
        RECT 26.200 144.100 26.600 144.200 ;
        RECT 28.600 144.100 29.000 144.200 ;
        RECT 87.800 144.100 88.200 144.200 ;
        RECT 26.200 143.800 88.200 144.100 ;
        RECT 95.000 144.100 95.400 144.200 ;
        RECT 97.400 144.100 97.800 144.200 ;
        RECT 95.000 143.800 97.800 144.100 ;
        RECT 239.000 144.100 239.400 144.200 ;
        RECT 239.800 144.100 240.200 144.200 ;
        RECT 239.000 143.800 240.200 144.100 ;
        RECT 21.400 143.100 21.800 143.200 ;
        RECT 101.400 143.100 101.800 143.200 ;
        RECT 117.400 143.100 117.800 143.200 ;
        RECT 203.800 143.100 204.200 143.200 ;
        RECT 21.400 142.800 204.200 143.100 ;
        RECT 238.200 143.100 238.600 143.200 ;
        RECT 239.000 143.100 239.400 143.200 ;
        RECT 240.600 143.100 241.000 143.200 ;
        RECT 238.200 142.800 241.000 143.100 ;
        RECT 25.400 142.100 25.800 142.200 ;
        RECT 30.200 142.100 30.600 142.200 ;
        RECT 37.400 142.100 37.800 142.200 ;
        RECT 25.400 141.800 37.800 142.100 ;
        RECT 75.000 142.100 75.400 142.200 ;
        RECT 76.600 142.100 77.000 142.200 ;
        RECT 75.000 141.800 77.000 142.100 ;
        RECT 93.400 142.100 93.800 142.200 ;
        RECT 116.600 142.100 117.000 142.200 ;
        RECT 93.400 141.800 117.000 142.100 ;
        RECT 143.000 142.100 143.400 142.200 ;
        RECT 147.800 142.100 148.200 142.200 ;
        RECT 155.000 142.100 155.400 142.200 ;
        RECT 143.000 141.800 155.400 142.100 ;
        RECT 158.200 142.100 158.600 142.200 ;
        RECT 184.600 142.100 185.000 142.200 ;
        RECT 158.200 141.800 185.000 142.100 ;
        RECT 36.600 141.100 37.000 141.200 ;
        RECT 43.000 141.100 43.400 141.200 ;
        RECT 36.600 140.800 43.400 141.100 ;
        RECT 51.000 141.100 51.400 141.200 ;
        RECT 66.200 141.100 66.600 141.200 ;
        RECT 51.000 140.800 66.600 141.100 ;
        RECT 88.600 141.100 89.000 141.200 ;
        RECT 94.200 141.100 94.600 141.200 ;
        RECT 88.600 140.800 94.600 141.100 ;
        RECT 127.000 141.100 127.400 141.200 ;
        RECT 146.200 141.100 146.600 141.200 ;
        RECT 127.000 140.800 146.600 141.100 ;
        RECT 183.800 141.100 184.200 141.200 ;
        RECT 193.400 141.100 193.800 141.200 ;
        RECT 183.800 140.800 193.800 141.100 ;
        RECT 212.600 141.100 213.000 141.200 ;
        RECT 213.400 141.100 213.800 141.200 ;
        RECT 215.800 141.100 216.200 141.200 ;
        RECT 212.600 140.800 216.200 141.100 ;
        RECT 10.200 140.100 10.600 140.200 ;
        RECT 23.000 140.100 23.400 140.200 ;
        RECT 10.200 139.800 23.400 140.100 ;
        RECT 51.800 140.100 52.200 140.200 ;
        RECT 65.400 140.100 65.800 140.200 ;
        RECT 72.600 140.100 73.000 140.200 ;
        RECT 51.800 139.800 73.000 140.100 ;
        RECT 73.400 140.100 73.800 140.200 ;
        RECT 75.800 140.100 76.200 140.200 ;
        RECT 73.400 139.800 76.200 140.100 ;
        RECT 78.200 140.100 78.600 140.200 ;
        RECT 111.800 140.100 112.200 140.200 ;
        RECT 78.200 139.800 112.200 140.100 ;
        RECT 187.800 140.100 188.200 140.200 ;
        RECT 192.600 140.100 193.000 140.200 ;
        RECT 187.800 139.800 193.000 140.100 ;
        RECT 3.800 139.100 4.200 139.200 ;
        RECT 12.600 139.100 13.000 139.200 ;
        RECT 27.000 139.100 27.400 139.200 ;
        RECT 45.400 139.100 45.800 139.200 ;
        RECT 67.800 139.100 68.200 139.200 ;
        RECT 3.800 138.800 27.400 139.100 ;
        RECT 44.600 138.800 68.200 139.100 ;
        RECT 85.400 139.100 85.800 139.200 ;
        RECT 93.400 139.100 93.800 139.200 ;
        RECT 85.400 138.800 93.800 139.100 ;
        RECT 107.000 139.100 107.400 139.200 ;
        RECT 111.000 139.100 111.400 139.200 ;
        RECT 155.800 139.100 156.200 139.200 ;
        RECT 107.000 138.800 156.200 139.100 ;
        RECT 156.600 139.100 157.000 139.200 ;
        RECT 197.400 139.100 197.800 139.200 ;
        RECT 156.600 138.800 197.800 139.100 ;
        RECT 15.000 138.100 15.400 138.200 ;
        RECT 17.400 138.100 17.800 138.200 ;
        RECT 59.800 138.100 60.200 138.200 ;
        RECT 15.000 137.800 60.200 138.100 ;
        RECT 63.000 138.100 63.400 138.200 ;
        RECT 71.800 138.100 72.200 138.200 ;
        RECT 101.400 138.100 101.800 138.200 ;
        RECT 63.000 137.800 101.800 138.100 ;
        RECT 120.600 138.100 121.000 138.200 ;
        RECT 133.400 138.100 133.800 138.200 ;
        RECT 120.600 137.800 133.800 138.100 ;
        RECT 155.000 138.100 155.400 138.200 ;
        RECT 194.200 138.100 194.600 138.200 ;
        RECT 155.000 137.800 194.600 138.100 ;
        RECT 48.600 137.100 49.000 137.200 ;
        RECT 24.600 136.800 49.000 137.100 ;
        RECT 64.600 137.100 65.000 137.200 ;
        RECT 70.200 137.100 70.600 137.200 ;
        RECT 64.600 136.800 70.600 137.100 ;
        RECT 73.400 136.800 73.800 137.200 ;
        RECT 86.200 137.100 86.600 137.200 ;
        RECT 109.400 137.100 109.800 137.200 ;
        RECT 131.000 137.100 131.400 137.200 ;
        RECT 86.200 136.800 131.400 137.100 ;
        RECT 167.800 136.800 168.200 137.200 ;
        RECT 184.600 136.800 185.000 137.200 ;
        RECT 191.000 137.100 191.400 137.200 ;
        RECT 211.800 137.100 212.200 137.200 ;
        RECT 216.600 137.100 217.000 137.200 ;
        RECT 191.000 136.800 217.000 137.100 ;
        RECT 24.600 136.200 24.900 136.800 ;
        RECT 16.600 136.100 17.000 136.200 ;
        RECT 16.600 135.800 20.100 136.100 ;
        RECT 24.600 135.800 25.000 136.200 ;
        RECT 27.000 136.100 27.400 136.200 ;
        RECT 64.600 136.100 65.000 136.200 ;
        RECT 27.000 135.800 65.000 136.100 ;
        RECT 73.400 136.100 73.700 136.800 ;
        RECT 85.400 136.100 85.800 136.200 ;
        RECT 73.400 135.800 85.800 136.100 ;
        RECT 86.200 136.100 86.600 136.200 ;
        RECT 87.800 136.100 88.200 136.200 ;
        RECT 89.400 136.100 89.800 136.200 ;
        RECT 86.200 135.800 89.800 136.100 ;
        RECT 93.400 135.800 93.800 136.200 ;
        RECT 100.600 136.100 101.000 136.200 ;
        RECT 114.200 136.100 114.600 136.200 ;
        RECT 115.800 136.100 116.200 136.200 ;
        RECT 100.600 135.800 116.200 136.100 ;
        RECT 119.800 136.100 120.200 136.200 ;
        RECT 123.800 136.100 124.200 136.200 ;
        RECT 119.800 135.800 124.200 136.100 ;
        RECT 135.800 136.100 136.200 136.200 ;
        RECT 139.000 136.100 139.400 136.200 ;
        RECT 135.800 135.800 139.400 136.100 ;
        RECT 146.200 136.100 146.600 136.200 ;
        RECT 147.800 136.100 148.200 136.200 ;
        RECT 165.400 136.100 165.800 136.200 ;
        RECT 146.200 135.800 165.800 136.100 ;
        RECT 167.800 136.100 168.100 136.800 ;
        RECT 176.600 136.100 177.000 136.200 ;
        RECT 167.800 135.800 177.000 136.100 ;
        RECT 182.200 136.100 182.600 136.200 ;
        RECT 184.600 136.100 184.900 136.800 ;
        RECT 182.200 135.800 184.900 136.100 ;
        RECT 195.800 136.100 196.200 136.200 ;
        RECT 197.400 136.100 197.800 136.200 ;
        RECT 195.800 135.800 197.800 136.100 ;
        RECT 210.200 136.100 210.600 136.200 ;
        RECT 230.200 136.100 230.600 136.200 ;
        RECT 210.200 135.800 230.600 136.100 ;
        RECT 231.800 136.100 232.200 136.200 ;
        RECT 238.200 136.100 238.600 136.200 ;
        RECT 231.800 135.800 238.600 136.100 ;
        RECT 19.800 135.200 20.100 135.800 ;
        RECT 8.600 135.100 9.000 135.200 ;
        RECT 16.600 135.100 17.000 135.200 ;
        RECT 8.600 134.800 17.000 135.100 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 41.400 135.100 41.800 135.200 ;
        RECT 40.600 134.800 41.800 135.100 ;
        RECT 43.000 135.100 43.400 135.200 ;
        RECT 45.400 135.100 45.800 135.200 ;
        RECT 43.000 134.800 45.800 135.100 ;
        RECT 46.200 135.100 46.600 135.200 ;
        RECT 47.000 135.100 47.400 135.200 ;
        RECT 46.200 134.800 47.400 135.100 ;
        RECT 51.800 135.100 52.200 135.200 ;
        RECT 63.000 135.100 63.400 135.200 ;
        RECT 51.800 134.800 63.400 135.100 ;
        RECT 79.800 135.100 80.200 135.200 ;
        RECT 81.400 135.100 81.800 135.200 ;
        RECT 84.600 135.100 85.000 135.200 ;
        RECT 85.400 135.100 85.800 135.200 ;
        RECT 79.800 134.800 85.800 135.100 ;
        RECT 88.600 135.100 89.000 135.200 ;
        RECT 93.400 135.100 93.700 135.800 ;
        RECT 123.800 135.200 124.100 135.800 ;
        RECT 88.600 134.800 93.700 135.100 ;
        RECT 95.800 135.100 96.200 135.200 ;
        RECT 104.600 135.100 105.000 135.200 ;
        RECT 95.800 134.800 105.000 135.100 ;
        RECT 106.200 135.100 106.600 135.200 ;
        RECT 113.400 135.100 113.800 135.200 ;
        RECT 106.200 134.800 113.800 135.100 ;
        RECT 123.800 135.100 124.200 135.200 ;
        RECT 125.400 135.100 125.800 135.200 ;
        RECT 123.800 134.800 125.800 135.100 ;
        RECT 150.200 135.100 150.600 135.200 ;
        RECT 153.400 135.100 153.800 135.200 ;
        RECT 150.200 134.800 153.800 135.100 ;
        RECT 156.600 135.100 157.000 135.200 ;
        RECT 157.400 135.100 157.800 135.200 ;
        RECT 156.600 134.800 157.800 135.100 ;
        RECT 164.600 135.100 165.000 135.200 ;
        RECT 169.400 135.100 169.800 135.200 ;
        RECT 164.600 134.800 169.800 135.100 ;
        RECT 171.800 135.100 172.200 135.200 ;
        RECT 174.200 135.100 174.600 135.200 ;
        RECT 171.800 134.800 174.600 135.100 ;
        RECT 179.800 135.100 180.200 135.200 ;
        RECT 189.400 135.100 189.800 135.200 ;
        RECT 179.800 134.800 189.800 135.100 ;
        RECT 198.200 135.100 198.600 135.200 ;
        RECT 207.000 135.100 207.400 135.200 ;
        RECT 198.200 134.800 207.400 135.100 ;
        RECT 214.200 135.100 214.600 135.200 ;
        RECT 222.200 135.100 222.600 135.200 ;
        RECT 214.200 134.800 222.600 135.100 ;
        RECT 233.400 134.800 237.700 135.100 ;
        RECT 233.400 134.200 233.700 134.800 ;
        RECT 237.400 134.200 237.700 134.800 ;
        RECT 15.000 134.100 15.400 134.200 ;
        RECT 15.800 134.100 16.200 134.200 ;
        RECT 26.200 134.100 26.600 134.200 ;
        RECT 28.600 134.100 29.000 134.200 ;
        RECT 15.000 133.800 29.000 134.100 ;
        RECT 40.600 134.100 41.000 134.200 ;
        RECT 52.600 134.100 53.000 134.200 ;
        RECT 40.600 133.800 53.000 134.100 ;
        RECT 58.200 134.100 58.600 134.200 ;
        RECT 63.800 134.100 64.200 134.200 ;
        RECT 58.200 133.800 64.200 134.100 ;
        RECT 75.800 134.100 76.200 134.200 ;
        RECT 79.000 134.100 79.400 134.200 ;
        RECT 75.800 133.800 79.400 134.100 ;
        RECT 80.600 134.100 81.000 134.200 ;
        RECT 103.000 134.100 103.400 134.200 ;
        RECT 80.600 133.800 103.400 134.100 ;
        RECT 116.600 134.100 117.000 134.200 ;
        RECT 126.200 134.100 126.600 134.200 ;
        RECT 116.600 133.800 126.600 134.100 ;
        RECT 147.800 134.100 148.200 134.200 ;
        RECT 148.600 134.100 149.000 134.200 ;
        RECT 147.800 133.800 149.000 134.100 ;
        RECT 151.800 134.100 152.200 134.200 ;
        RECT 155.000 134.100 155.400 134.200 ;
        RECT 151.800 133.800 155.400 134.100 ;
        RECT 159.000 134.100 159.400 134.200 ;
        RECT 172.600 134.100 173.000 134.200 ;
        RECT 159.000 133.800 173.000 134.100 ;
        RECT 175.800 134.100 176.200 134.200 ;
        RECT 187.800 134.100 188.200 134.200 ;
        RECT 194.200 134.100 194.600 134.200 ;
        RECT 175.800 133.800 188.200 134.100 ;
        RECT 188.600 133.800 194.600 134.100 ;
        RECT 215.000 134.100 215.400 134.200 ;
        RECT 217.400 134.100 217.800 134.200 ;
        RECT 215.000 133.800 217.800 134.100 ;
        RECT 233.400 133.800 233.800 134.200 ;
        RECT 237.400 133.800 237.800 134.200 ;
        RECT 188.600 133.200 188.900 133.800 ;
        RECT 13.400 133.100 13.800 133.200 ;
        RECT 19.000 133.100 19.400 133.200 ;
        RECT 13.400 132.800 19.400 133.100 ;
        RECT 21.400 133.100 21.800 133.200 ;
        RECT 25.400 133.100 25.800 133.200 ;
        RECT 27.800 133.100 28.200 133.200 ;
        RECT 21.400 132.800 28.200 133.100 ;
        RECT 43.000 133.100 43.400 133.200 ;
        RECT 51.000 133.100 51.400 133.200 ;
        RECT 43.000 132.800 51.400 133.100 ;
        RECT 54.200 133.100 54.600 133.200 ;
        RECT 60.600 133.100 61.000 133.200 ;
        RECT 74.200 133.100 74.600 133.200 ;
        RECT 54.200 132.800 74.600 133.100 ;
        RECT 84.600 133.100 85.000 133.200 ;
        RECT 88.600 133.100 89.000 133.200 ;
        RECT 84.600 132.800 89.000 133.100 ;
        RECT 130.200 133.100 130.600 133.200 ;
        RECT 137.400 133.100 137.800 133.200 ;
        RECT 183.000 133.100 183.400 133.200 ;
        RECT 187.000 133.100 187.400 133.200 ;
        RECT 130.200 132.800 187.400 133.100 ;
        RECT 188.600 132.800 189.000 133.200 ;
        RECT 14.200 132.100 14.600 132.200 ;
        RECT 31.800 132.100 32.200 132.200 ;
        RECT 14.200 131.800 32.200 132.100 ;
        RECT 39.000 132.100 39.400 132.200 ;
        RECT 45.400 132.100 45.800 132.200 ;
        RECT 83.800 132.100 84.200 132.200 ;
        RECT 39.000 131.800 84.200 132.100 ;
        RECT 90.200 132.100 90.600 132.200 ;
        RECT 97.400 132.100 97.800 132.200 ;
        RECT 99.000 132.100 99.400 132.200 ;
        RECT 90.200 131.800 99.400 132.100 ;
        RECT 113.400 132.100 113.800 132.200 ;
        RECT 122.200 132.100 122.600 132.200 ;
        RECT 127.000 132.100 127.400 132.200 ;
        RECT 113.400 131.800 127.400 132.100 ;
        RECT 131.800 132.100 132.200 132.200 ;
        RECT 140.600 132.100 141.000 132.200 ;
        RECT 180.600 132.100 181.000 132.200 ;
        RECT 186.200 132.100 186.600 132.200 ;
        RECT 131.800 131.800 186.600 132.100 ;
        RECT 228.600 132.100 229.000 132.200 ;
        RECT 248.600 132.100 249.000 132.200 ;
        RECT 228.600 131.800 249.000 132.100 ;
        RECT 37.400 131.100 37.800 131.200 ;
        RECT 44.600 131.100 45.000 131.200 ;
        RECT 37.400 130.800 45.000 131.100 ;
        RECT 52.600 131.100 53.000 131.200 ;
        RECT 59.800 131.100 60.200 131.200 ;
        RECT 52.600 130.800 60.200 131.100 ;
        RECT 79.800 131.100 80.200 131.200 ;
        RECT 82.200 131.100 82.600 131.200 ;
        RECT 79.800 130.800 82.600 131.100 ;
        RECT 124.600 131.100 125.000 131.200 ;
        RECT 133.400 131.100 133.800 131.200 ;
        RECT 124.600 130.800 133.800 131.100 ;
        RECT 135.000 131.100 135.400 131.200 ;
        RECT 138.200 131.100 138.600 131.200 ;
        RECT 151.800 131.100 152.200 131.200 ;
        RECT 156.600 131.100 157.000 131.200 ;
        RECT 135.000 130.800 157.000 131.100 ;
        RECT 169.400 131.100 169.800 131.200 ;
        RECT 184.600 131.100 185.000 131.200 ;
        RECT 169.400 130.800 185.000 131.100 ;
        RECT 186.200 131.100 186.600 131.200 ;
        RECT 191.000 131.100 191.400 131.200 ;
        RECT 186.200 130.800 191.400 131.100 ;
        RECT 206.200 131.100 206.600 131.200 ;
        RECT 225.400 131.100 225.800 131.200 ;
        RECT 234.200 131.100 234.600 131.200 ;
        RECT 243.800 131.100 244.200 131.200 ;
        RECT 206.200 130.800 244.200 131.100 ;
        RECT 32.600 130.100 33.000 130.200 ;
        RECT 47.000 130.100 47.400 130.200 ;
        RECT 32.600 129.800 47.400 130.100 ;
        RECT 53.400 130.100 53.800 130.200 ;
        RECT 68.600 130.100 69.000 130.200 ;
        RECT 82.200 130.100 82.600 130.200 ;
        RECT 53.400 129.800 82.600 130.100 ;
        RECT 115.800 130.100 116.200 130.200 ;
        RECT 131.000 130.100 131.400 130.200 ;
        RECT 115.800 129.800 131.400 130.100 ;
        RECT 145.400 130.100 145.800 130.200 ;
        RECT 157.400 130.100 157.800 130.200 ;
        RECT 164.600 130.100 165.000 130.200 ;
        RECT 175.000 130.100 175.400 130.200 ;
        RECT 188.600 130.100 189.000 130.200 ;
        RECT 145.400 129.800 189.000 130.100 ;
        RECT 216.600 130.100 217.000 130.200 ;
        RECT 227.000 130.100 227.400 130.200 ;
        RECT 235.800 130.100 236.200 130.200 ;
        RECT 216.600 129.800 236.200 130.100 ;
        RECT 241.400 129.800 241.800 130.200 ;
        RECT 19.000 129.100 19.400 129.200 ;
        RECT 39.000 129.100 39.400 129.200 ;
        RECT 19.000 128.800 39.400 129.100 ;
        RECT 43.800 128.800 44.200 129.200 ;
        RECT 45.400 128.800 45.800 129.200 ;
        RECT 58.200 129.100 58.600 129.200 ;
        RECT 71.000 129.100 71.400 129.200 ;
        RECT 87.000 129.100 87.400 129.200 ;
        RECT 58.200 128.800 62.500 129.100 ;
        RECT 71.000 128.800 87.400 129.100 ;
        RECT 89.400 129.100 89.800 129.200 ;
        RECT 91.000 129.100 91.400 129.200 ;
        RECT 89.400 128.800 91.400 129.100 ;
        RECT 93.400 129.100 93.800 129.200 ;
        RECT 119.800 129.100 120.200 129.200 ;
        RECT 128.600 129.100 129.000 129.200 ;
        RECT 93.400 128.800 129.000 129.100 ;
        RECT 138.200 129.100 138.600 129.200 ;
        RECT 139.800 129.100 140.200 129.200 ;
        RECT 154.200 129.100 154.600 129.200 ;
        RECT 138.200 128.800 154.600 129.100 ;
        RECT 165.400 129.100 165.800 129.200 ;
        RECT 167.000 129.100 167.400 129.200 ;
        RECT 165.400 128.800 167.400 129.100 ;
        RECT 175.000 129.100 175.400 129.200 ;
        RECT 183.800 129.100 184.200 129.200 ;
        RECT 186.200 129.100 186.600 129.200 ;
        RECT 175.000 128.800 186.600 129.100 ;
        RECT 193.400 129.100 193.800 129.200 ;
        RECT 201.400 129.100 201.800 129.200 ;
        RECT 210.200 129.100 210.600 129.200 ;
        RECT 193.400 128.800 210.600 129.100 ;
        RECT 215.000 129.100 215.400 129.200 ;
        RECT 225.400 129.100 225.800 129.200 ;
        RECT 215.000 128.800 225.800 129.100 ;
        RECT 241.400 129.100 241.700 129.800 ;
        RECT 247.000 129.100 247.400 129.200 ;
        RECT 241.400 128.800 247.400 129.100 ;
        RECT 9.400 128.100 9.800 128.200 ;
        RECT 11.800 128.100 12.200 128.200 ;
        RECT 28.600 128.100 29.000 128.200 ;
        RECT 9.400 127.800 29.000 128.100 ;
        RECT 43.800 128.100 44.100 128.800 ;
        RECT 45.400 128.100 45.700 128.800 ;
        RECT 43.800 127.800 45.700 128.100 ;
        RECT 62.200 128.200 62.500 128.800 ;
        RECT 62.200 127.800 62.600 128.200 ;
        RECT 69.400 128.100 69.800 128.200 ;
        RECT 84.600 128.100 85.000 128.200 ;
        RECT 69.400 127.800 85.000 128.100 ;
        RECT 86.200 128.100 86.600 128.200 ;
        RECT 101.400 128.100 101.800 128.200 ;
        RECT 86.200 127.800 101.800 128.100 ;
        RECT 102.200 128.100 102.600 128.200 ;
        RECT 119.000 128.100 119.400 128.200 ;
        RECT 102.200 127.800 119.400 128.100 ;
        RECT 142.200 128.100 142.600 128.200 ;
        RECT 147.000 128.100 147.400 128.200 ;
        RECT 142.200 127.800 147.400 128.100 ;
        RECT 150.200 128.100 150.600 128.200 ;
        RECT 159.800 128.100 160.200 128.200 ;
        RECT 150.200 127.800 160.200 128.100 ;
        RECT 174.200 128.100 174.600 128.200 ;
        RECT 181.400 128.100 181.800 128.200 ;
        RECT 174.200 127.800 181.800 128.100 ;
        RECT 191.000 128.100 191.400 128.200 ;
        RECT 195.000 128.100 195.400 128.200 ;
        RECT 191.000 127.800 195.400 128.100 ;
        RECT 197.400 128.100 197.800 128.200 ;
        RECT 218.200 128.100 218.600 128.200 ;
        RECT 197.400 127.800 218.600 128.100 ;
        RECT 240.600 128.100 241.000 128.200 ;
        RECT 241.400 128.100 241.800 128.200 ;
        RECT 240.600 127.800 241.800 128.100 ;
        RECT 5.400 127.100 5.800 127.200 ;
        RECT 17.400 127.100 17.800 127.200 ;
        RECT 22.200 127.100 22.600 127.200 ;
        RECT 5.400 126.800 12.900 127.100 ;
        RECT 17.400 126.800 22.600 127.100 ;
        RECT 23.800 127.100 24.200 127.200 ;
        RECT 29.400 127.100 29.800 127.200 ;
        RECT 23.800 126.800 29.800 127.100 ;
        RECT 42.200 126.800 42.600 127.200 ;
        RECT 49.400 127.100 49.800 127.200 ;
        RECT 65.400 127.100 65.800 127.200 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 69.400 127.100 69.800 127.200 ;
        RECT 49.400 126.800 69.800 127.100 ;
        RECT 78.200 127.100 78.600 127.200 ;
        RECT 82.200 127.100 82.600 127.200 ;
        RECT 78.200 126.800 82.600 127.100 ;
        RECT 94.200 126.800 94.600 127.200 ;
        RECT 97.400 126.800 97.800 127.200 ;
        RECT 101.400 127.100 101.800 127.200 ;
        RECT 102.200 127.100 102.600 127.200 ;
        RECT 101.400 126.800 102.600 127.100 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 114.200 127.100 114.600 127.200 ;
        RECT 115.000 127.100 115.400 127.200 ;
        RECT 114.200 126.800 115.400 127.100 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 136.600 127.100 137.000 127.200 ;
        RECT 141.400 127.100 141.800 127.200 ;
        RECT 136.600 126.800 141.800 127.100 ;
        RECT 143.800 127.100 144.200 127.200 ;
        RECT 161.400 127.100 161.800 127.200 ;
        RECT 173.400 127.100 173.800 127.200 ;
        RECT 143.800 126.800 173.800 127.100 ;
        RECT 189.400 127.100 189.800 127.200 ;
        RECT 195.000 127.100 195.400 127.200 ;
        RECT 189.400 126.800 195.400 127.100 ;
        RECT 207.000 126.800 207.400 127.200 ;
        RECT 220.600 127.100 221.000 127.200 ;
        RECT 224.600 127.100 225.000 127.200 ;
        RECT 220.600 126.800 225.000 127.100 ;
        RECT 226.200 127.100 226.600 127.200 ;
        RECT 239.000 127.100 239.400 127.200 ;
        RECT 226.200 126.800 239.400 127.100 ;
        RECT 245.400 127.100 245.800 127.200 ;
        RECT 247.000 127.100 247.400 127.200 ;
        RECT 245.400 126.800 247.400 127.100 ;
        RECT 12.600 126.200 12.900 126.800 ;
        RECT 12.600 125.800 13.000 126.200 ;
        RECT 16.600 126.100 17.000 126.200 ;
        RECT 17.400 126.100 17.800 126.200 ;
        RECT 16.600 125.800 17.800 126.100 ;
        RECT 18.200 125.800 18.600 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 30.200 125.800 36.200 126.100 ;
        RECT 38.200 125.800 38.600 126.200 ;
        RECT 42.200 126.100 42.500 126.800 ;
        RECT 94.200 126.200 94.500 126.800 ;
        RECT 97.400 126.200 97.700 126.800 ;
        RECT 44.600 126.100 45.000 126.200 ;
        RECT 48.600 126.100 49.000 126.200 ;
        RECT 42.200 125.800 49.000 126.100 ;
        RECT 58.200 126.100 58.600 126.200 ;
        RECT 68.600 126.100 69.000 126.200 ;
        RECT 58.200 125.800 69.000 126.100 ;
        RECT 77.400 126.100 77.800 126.200 ;
        RECT 78.200 126.100 78.600 126.200 ;
        RECT 77.400 125.800 78.600 126.100 ;
        RECT 82.200 126.100 82.600 126.200 ;
        RECT 83.000 126.100 83.400 126.200 ;
        RECT 92.600 126.100 93.000 126.200 ;
        RECT 82.200 125.800 93.000 126.100 ;
        RECT 94.200 125.800 94.600 126.200 ;
        RECT 97.400 125.800 97.800 126.200 ;
        RECT 100.600 126.100 101.000 126.200 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 100.600 125.800 105.000 126.100 ;
        RECT 108.600 126.100 108.900 126.800 ;
        RECT 110.200 126.100 110.600 126.200 ;
        RECT 108.600 125.800 110.600 126.100 ;
        RECT 118.200 126.100 118.600 126.200 ;
        RECT 123.800 126.100 124.100 126.800 ;
        RECT 118.200 125.800 124.100 126.100 ;
        RECT 155.800 126.100 156.200 126.300 ;
        RECT 161.400 126.100 161.800 126.200 ;
        RECT 155.800 125.800 161.800 126.100 ;
        RECT 165.400 126.100 165.800 126.200 ;
        RECT 175.800 126.100 176.200 126.200 ;
        RECT 165.400 125.800 176.200 126.100 ;
        RECT 185.400 125.800 185.800 126.200 ;
        RECT 191.000 126.100 191.400 126.200 ;
        RECT 199.000 126.100 199.400 126.200 ;
        RECT 191.000 125.800 199.400 126.100 ;
        RECT 207.000 126.100 207.300 126.800 ;
        RECT 211.800 126.100 212.200 126.200 ;
        RECT 207.000 125.800 212.200 126.100 ;
        RECT 219.800 126.100 220.200 126.200 ;
        RECT 222.200 126.100 222.600 126.200 ;
        RECT 226.200 126.100 226.600 126.200 ;
        RECT 239.000 126.100 239.400 126.200 ;
        RECT 219.800 125.800 226.600 126.100 ;
        RECT 238.200 125.800 239.400 126.100 ;
        RECT 240.600 126.100 241.000 126.200 ;
        RECT 244.600 126.100 245.000 126.200 ;
        RECT 240.600 125.800 245.000 126.100 ;
        RECT 4.600 125.100 5.000 125.200 ;
        RECT 11.000 125.100 11.400 125.200 ;
        RECT 14.200 125.100 14.600 125.200 ;
        RECT 4.600 124.800 14.600 125.100 ;
        RECT 18.200 125.100 18.500 125.800 ;
        RECT 30.200 125.200 30.500 125.800 ;
        RECT 38.200 125.200 38.500 125.800 ;
        RECT 185.400 125.200 185.700 125.800 ;
        RECT 238.200 125.200 238.500 125.800 ;
        RECT 19.800 125.100 20.200 125.200 ;
        RECT 18.200 124.800 20.200 125.100 ;
        RECT 30.200 124.800 30.600 125.200 ;
        RECT 33.400 125.100 33.800 125.200 ;
        RECT 35.000 125.100 35.400 125.200 ;
        RECT 33.400 124.800 35.400 125.100 ;
        RECT 38.200 124.800 38.600 125.200 ;
        RECT 46.200 125.100 46.600 125.200 ;
        RECT 55.800 125.100 56.200 125.200 ;
        RECT 46.200 124.800 56.200 125.100 ;
        RECT 62.200 125.100 62.600 125.200 ;
        RECT 63.800 125.100 64.200 125.200 ;
        RECT 62.200 124.800 64.200 125.100 ;
        RECT 64.600 125.100 65.000 125.200 ;
        RECT 65.400 125.100 65.800 125.200 ;
        RECT 71.000 125.100 71.400 125.200 ;
        RECT 64.600 124.800 71.400 125.100 ;
        RECT 72.600 125.100 73.000 125.200 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 86.200 125.100 86.600 125.200 ;
        RECT 72.600 124.800 86.600 125.100 ;
        RECT 92.600 125.100 93.000 125.200 ;
        RECT 111.000 125.100 111.400 125.200 ;
        RECT 92.600 124.800 111.400 125.100 ;
        RECT 115.000 125.100 115.400 125.200 ;
        RECT 117.400 125.100 117.800 125.200 ;
        RECT 115.000 124.800 117.800 125.100 ;
        RECT 127.800 125.100 128.200 125.200 ;
        RECT 160.600 125.100 161.000 125.200 ;
        RECT 163.800 125.100 164.200 125.200 ;
        RECT 166.200 125.100 166.600 125.200 ;
        RECT 127.800 124.800 166.600 125.100 ;
        RECT 172.600 125.100 173.000 125.200 ;
        RECT 178.200 125.100 178.600 125.200 ;
        RECT 172.600 124.800 178.600 125.100 ;
        RECT 185.400 124.800 185.800 125.200 ;
        RECT 211.800 125.100 212.200 125.200 ;
        RECT 212.600 125.100 213.000 125.200 ;
        RECT 214.200 125.100 214.600 125.200 ;
        RECT 211.800 124.800 214.600 125.100 ;
        RECT 219.800 125.100 220.200 125.200 ;
        RECT 220.600 125.100 221.000 125.200 ;
        RECT 231.800 125.100 232.200 125.200 ;
        RECT 219.800 124.800 221.000 125.100 ;
        RECT 224.600 124.800 232.200 125.100 ;
        RECT 238.200 124.800 238.600 125.200 ;
        RECT 239.000 125.100 239.400 125.200 ;
        RECT 248.600 125.100 249.000 125.200 ;
        RECT 239.000 124.800 249.000 125.100 ;
        RECT 224.600 124.200 224.900 124.800 ;
        RECT 10.200 124.100 10.600 124.200 ;
        RECT 31.800 124.100 32.200 124.200 ;
        RECT 10.200 123.800 32.200 124.100 ;
        RECT 35.800 124.100 36.200 124.200 ;
        RECT 43.000 124.100 43.400 124.200 ;
        RECT 47.000 124.100 47.400 124.200 ;
        RECT 139.800 124.100 140.200 124.200 ;
        RECT 35.800 123.800 140.200 124.100 ;
        RECT 153.400 124.100 153.800 124.200 ;
        RECT 166.200 124.100 166.600 124.200 ;
        RECT 153.400 123.800 166.600 124.100 ;
        RECT 168.600 124.100 169.000 124.200 ;
        RECT 178.200 124.100 178.600 124.200 ;
        RECT 168.600 123.800 178.600 124.100 ;
        RECT 192.600 124.100 193.000 124.200 ;
        RECT 215.000 124.100 215.400 124.200 ;
        RECT 215.800 124.100 216.200 124.200 ;
        RECT 192.600 123.800 216.200 124.100 ;
        RECT 224.600 123.800 225.000 124.200 ;
        RECT 46.200 123.100 46.600 123.200 ;
        RECT 49.400 123.100 49.800 123.200 ;
        RECT 46.200 122.800 49.800 123.100 ;
        RECT 71.000 123.100 71.400 123.200 ;
        RECT 89.400 123.100 89.800 123.200 ;
        RECT 71.000 122.800 89.800 123.100 ;
        RECT 95.000 123.100 95.400 123.200 ;
        RECT 100.600 123.100 101.000 123.200 ;
        RECT 95.000 122.800 101.000 123.100 ;
        RECT 103.000 123.100 103.400 123.200 ;
        RECT 171.000 123.100 171.400 123.200 ;
        RECT 173.400 123.100 173.800 123.200 ;
        RECT 179.800 123.100 180.200 123.200 ;
        RECT 103.000 122.800 180.200 123.100 ;
        RECT 243.000 123.100 243.400 123.200 ;
        RECT 245.400 123.100 245.800 123.200 ;
        RECT 243.000 122.800 245.800 123.100 ;
        RECT 12.600 122.100 13.000 122.200 ;
        RECT 13.400 122.100 13.800 122.200 ;
        RECT 67.000 122.100 67.400 122.200 ;
        RECT 12.600 121.800 67.400 122.100 ;
        RECT 74.200 122.100 74.600 122.200 ;
        RECT 87.800 122.100 88.200 122.200 ;
        RECT 103.800 122.100 104.200 122.200 ;
        RECT 74.200 121.800 104.200 122.100 ;
        RECT 105.400 122.100 105.800 122.200 ;
        RECT 110.200 122.100 110.600 122.200 ;
        RECT 105.400 121.800 110.600 122.100 ;
        RECT 115.800 122.100 116.200 122.200 ;
        RECT 141.400 122.100 141.800 122.200 ;
        RECT 143.800 122.100 144.200 122.200 ;
        RECT 115.800 121.800 144.200 122.100 ;
        RECT 181.400 122.100 181.800 122.200 ;
        RECT 183.000 122.100 183.400 122.200 ;
        RECT 202.200 122.100 202.600 122.200 ;
        RECT 181.400 121.800 202.600 122.100 ;
        RECT 25.400 121.100 25.800 121.200 ;
        RECT 34.200 121.100 34.600 121.200 ;
        RECT 25.400 120.800 34.600 121.100 ;
        RECT 67.000 121.100 67.400 121.200 ;
        RECT 115.800 121.100 116.200 121.200 ;
        RECT 67.000 120.800 116.200 121.100 ;
        RECT 121.400 121.100 121.800 121.200 ;
        RECT 139.000 121.100 139.400 121.200 ;
        RECT 121.400 120.800 139.400 121.100 ;
        RECT 191.800 121.100 192.200 121.200 ;
        RECT 195.800 121.100 196.200 121.200 ;
        RECT 198.200 121.100 198.600 121.200 ;
        RECT 191.800 120.800 198.600 121.100 ;
        RECT 203.800 121.100 204.200 121.200 ;
        RECT 230.200 121.100 230.600 121.200 ;
        RECT 203.800 120.800 230.600 121.100 ;
        RECT 63.800 119.800 64.200 120.200 ;
        RECT 66.200 120.100 66.600 120.200 ;
        RECT 71.800 120.100 72.200 120.200 ;
        RECT 66.200 119.800 72.200 120.100 ;
        RECT 79.800 120.100 80.200 120.200 ;
        RECT 80.600 120.100 81.000 120.200 ;
        RECT 79.800 119.800 81.000 120.100 ;
        RECT 90.200 120.100 90.600 120.200 ;
        RECT 95.000 120.100 95.400 120.200 ;
        RECT 90.200 119.800 95.400 120.100 ;
        RECT 101.400 120.100 101.800 120.200 ;
        RECT 115.800 120.100 116.200 120.200 ;
        RECT 101.400 119.800 116.200 120.100 ;
        RECT 183.800 120.100 184.200 120.200 ;
        RECT 187.000 120.100 187.400 120.200 ;
        RECT 224.600 120.100 225.000 120.200 ;
        RECT 235.000 120.100 235.400 120.200 ;
        RECT 242.200 120.100 242.600 120.200 ;
        RECT 246.200 120.100 246.600 120.200 ;
        RECT 183.800 119.800 246.600 120.100 ;
        RECT 63.800 119.200 64.100 119.800 ;
        RECT 18.200 119.100 18.600 119.200 ;
        RECT 21.400 119.100 21.800 119.200 ;
        RECT 18.200 118.800 21.800 119.100 ;
        RECT 63.800 118.800 64.200 119.200 ;
        RECT 69.400 119.100 69.800 119.200 ;
        RECT 79.000 119.100 79.400 119.200 ;
        RECT 94.200 119.100 94.600 119.200 ;
        RECT 69.400 118.800 94.600 119.100 ;
        RECT 107.000 119.100 107.400 119.200 ;
        RECT 114.200 119.100 114.600 119.200 ;
        RECT 107.000 118.800 114.600 119.100 ;
        RECT 139.800 119.100 140.200 119.200 ;
        RECT 232.600 119.100 233.000 119.200 ;
        RECT 239.000 119.100 239.400 119.200 ;
        RECT 139.800 118.800 239.400 119.100 ;
        RECT 74.200 118.100 74.600 118.200 ;
        RECT 81.400 118.100 81.800 118.200 ;
        RECT 109.400 118.100 109.800 118.200 ;
        RECT 115.000 118.100 115.400 118.200 ;
        RECT 74.200 117.800 81.800 118.100 ;
        RECT 104.600 117.800 115.400 118.100 ;
        RECT 115.800 118.100 116.200 118.200 ;
        RECT 190.200 118.100 190.600 118.200 ;
        RECT 115.800 117.800 190.600 118.100 ;
        RECT 225.400 117.800 225.800 118.200 ;
        RECT 238.200 118.100 238.600 118.200 ;
        RECT 248.600 118.100 249.000 118.200 ;
        RECT 238.200 117.800 249.000 118.100 ;
        RECT 104.600 117.200 104.900 117.800 ;
        RECT 225.400 117.200 225.700 117.800 ;
        RECT 9.400 117.100 9.800 117.200 ;
        RECT 12.600 117.100 13.000 117.200 ;
        RECT 21.400 117.100 21.800 117.200 ;
        RECT 9.400 116.800 21.800 117.100 ;
        RECT 23.000 117.100 23.400 117.200 ;
        RECT 23.800 117.100 24.200 117.200 ;
        RECT 23.000 116.800 24.200 117.100 ;
        RECT 48.600 117.100 49.000 117.200 ;
        RECT 62.200 117.100 62.600 117.200 ;
        RECT 48.600 116.800 62.600 117.100 ;
        RECT 64.600 116.800 65.000 117.200 ;
        RECT 79.800 117.100 80.200 117.200 ;
        RECT 88.600 117.100 89.000 117.200 ;
        RECT 93.400 117.100 93.800 117.200 ;
        RECT 104.600 117.100 105.000 117.200 ;
        RECT 79.800 116.800 105.000 117.100 ;
        RECT 106.200 117.100 106.600 117.200 ;
        RECT 115.000 117.100 115.400 117.200 ;
        RECT 146.200 117.100 146.600 117.200 ;
        RECT 106.200 116.800 146.600 117.100 ;
        RECT 158.200 116.800 158.600 117.200 ;
        RECT 164.600 117.100 165.000 117.200 ;
        RECT 172.600 117.100 173.000 117.200 ;
        RECT 164.600 116.800 173.000 117.100 ;
        RECT 173.400 117.100 173.800 117.200 ;
        RECT 187.000 117.100 187.400 117.200 ;
        RECT 191.000 117.100 191.400 117.200 ;
        RECT 173.400 116.800 191.400 117.100 ;
        RECT 195.800 116.800 196.200 117.200 ;
        RECT 208.600 117.100 209.000 117.200 ;
        RECT 210.200 117.100 210.600 117.200 ;
        RECT 208.600 116.800 210.600 117.100 ;
        RECT 219.800 116.800 220.200 117.200 ;
        RECT 225.400 116.800 225.800 117.200 ;
        RECT 239.800 116.800 240.200 117.200 ;
        RECT 7.800 116.100 8.200 116.200 ;
        RECT 22.200 116.100 22.600 116.200 ;
        RECT 7.800 115.800 22.600 116.100 ;
        RECT 28.600 116.100 29.000 116.200 ;
        RECT 31.800 116.100 32.200 116.200 ;
        RECT 28.600 115.800 32.200 116.100 ;
        RECT 43.800 116.100 44.200 116.200 ;
        RECT 45.400 116.100 45.800 116.200 ;
        RECT 43.800 115.800 45.800 116.100 ;
        RECT 53.400 116.100 53.800 116.200 ;
        RECT 59.000 116.100 59.400 116.200 ;
        RECT 53.400 115.800 59.400 116.100 ;
        RECT 64.600 116.100 64.900 116.800 ;
        RECT 68.600 116.100 69.000 116.200 ;
        RECT 64.600 115.800 69.000 116.100 ;
        RECT 75.000 116.100 75.400 116.200 ;
        RECT 87.000 116.100 87.400 116.200 ;
        RECT 75.000 115.800 87.400 116.100 ;
        RECT 95.000 116.100 95.400 116.200 ;
        RECT 97.400 116.100 97.800 116.200 ;
        RECT 95.000 115.800 97.800 116.100 ;
        RECT 107.000 116.100 107.400 116.200 ;
        RECT 108.600 116.100 109.000 116.200 ;
        RECT 107.000 115.800 109.000 116.100 ;
        RECT 130.200 116.100 130.600 116.200 ;
        RECT 137.400 116.100 137.800 116.200 ;
        RECT 139.800 116.100 140.200 116.200 ;
        RECT 130.200 115.800 140.200 116.100 ;
        RECT 143.800 116.100 144.200 116.200 ;
        RECT 146.200 116.100 146.600 116.200 ;
        RECT 143.800 115.800 146.600 116.100 ;
        RECT 154.200 116.100 154.600 116.200 ;
        RECT 158.200 116.100 158.500 116.800 ;
        RECT 195.800 116.200 196.100 116.800 ;
        RECT 154.200 115.800 158.500 116.100 ;
        RECT 171.800 116.100 172.200 116.200 ;
        RECT 175.000 116.100 175.400 116.200 ;
        RECT 175.800 116.100 176.200 116.200 ;
        RECT 171.800 115.800 176.200 116.100 ;
        RECT 177.400 115.800 177.800 116.200 ;
        RECT 185.400 116.100 185.800 116.200 ;
        RECT 187.800 116.100 188.200 116.200 ;
        RECT 185.400 115.800 188.200 116.100 ;
        RECT 195.800 115.800 196.200 116.200 ;
        RECT 212.600 116.100 213.000 116.200 ;
        RECT 219.800 116.100 220.100 116.800 ;
        RECT 239.800 116.200 240.100 116.800 ;
        RECT 212.600 115.800 220.100 116.100 ;
        RECT 231.000 116.100 231.400 116.200 ;
        RECT 238.200 116.100 238.600 116.200 ;
        RECT 231.000 115.800 238.600 116.100 ;
        RECT 239.800 115.800 240.200 116.200 ;
        RECT 243.000 115.800 243.400 116.200 ;
        RECT 171.800 115.200 172.100 115.800 ;
        RECT 11.800 115.100 12.200 115.200 ;
        RECT 16.600 115.100 17.000 115.200 ;
        RECT 11.800 114.800 17.000 115.100 ;
        RECT 30.200 114.800 30.600 115.200 ;
        RECT 38.200 115.100 38.600 115.200 ;
        RECT 43.800 115.100 44.200 115.200 ;
        RECT 38.200 114.800 44.200 115.100 ;
        RECT 57.400 114.800 57.800 115.200 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 60.600 115.100 61.000 115.200 ;
        RECT 59.000 114.800 61.000 115.100 ;
        RECT 67.000 115.100 67.400 115.200 ;
        RECT 67.000 114.800 68.100 115.100 ;
        RECT 11.000 114.100 11.400 114.200 ;
        RECT 11.800 114.100 12.200 114.200 ;
        RECT 14.200 114.100 14.600 114.200 ;
        RECT 30.200 114.100 30.500 114.800 ;
        RECT 11.000 113.800 30.500 114.100 ;
        RECT 46.200 114.100 46.600 114.200 ;
        RECT 57.400 114.100 57.700 114.800 ;
        RECT 46.200 113.800 57.700 114.100 ;
        RECT 67.800 114.200 68.100 114.800 ;
        RECT 78.200 114.800 78.600 115.200 ;
        RECT 80.600 115.100 81.000 115.200 ;
        RECT 81.400 115.100 81.800 115.200 ;
        RECT 83.000 115.100 83.400 115.200 ;
        RECT 80.600 114.800 83.400 115.100 ;
        RECT 94.200 115.100 94.600 115.200 ;
        RECT 95.800 115.100 96.200 115.200 ;
        RECT 96.600 115.100 97.000 115.200 ;
        RECT 94.200 114.800 97.000 115.100 ;
        RECT 99.000 115.100 99.400 115.200 ;
        RECT 102.200 115.100 102.600 115.200 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 113.400 115.100 113.800 115.200 ;
        RECT 99.000 114.800 105.000 115.100 ;
        RECT 107.800 114.800 113.800 115.100 ;
        RECT 118.200 115.100 118.600 115.200 ;
        RECT 123.000 115.100 123.400 115.200 ;
        RECT 118.200 114.800 123.400 115.100 ;
        RECT 156.600 115.100 157.000 115.200 ;
        RECT 162.200 115.100 162.600 115.200 ;
        RECT 156.600 114.800 162.600 115.100 ;
        RECT 171.800 114.800 172.200 115.200 ;
        RECT 175.800 115.100 176.200 115.200 ;
        RECT 177.400 115.100 177.700 115.800 ;
        RECT 243.000 115.200 243.300 115.800 ;
        RECT 175.800 114.800 177.700 115.100 ;
        RECT 182.200 114.800 182.600 115.200 ;
        RECT 193.400 115.100 193.800 115.200 ;
        RECT 195.800 115.100 196.200 115.200 ;
        RECT 197.400 115.100 197.800 115.200 ;
        RECT 193.400 114.800 197.800 115.100 ;
        RECT 220.600 115.100 221.000 115.200 ;
        RECT 232.600 115.100 233.000 115.200 ;
        RECT 220.600 114.800 233.000 115.100 ;
        RECT 234.200 115.100 234.600 115.200 ;
        RECT 241.400 115.100 241.800 115.200 ;
        RECT 234.200 114.800 241.800 115.100 ;
        RECT 243.000 114.800 243.400 115.200 ;
        RECT 78.200 114.200 78.500 114.800 ;
        RECT 107.800 114.200 108.100 114.800 ;
        RECT 67.800 113.800 68.200 114.200 ;
        RECT 71.000 114.100 71.400 114.200 ;
        RECT 74.200 114.100 74.600 114.200 ;
        RECT 71.000 113.800 74.600 114.100 ;
        RECT 78.200 113.800 78.600 114.200 ;
        RECT 96.600 114.100 97.000 114.200 ;
        RECT 104.600 114.100 105.000 114.200 ;
        RECT 96.600 113.800 105.000 114.100 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 135.800 114.100 136.200 114.200 ;
        RECT 136.600 114.100 137.000 114.200 ;
        RECT 135.800 113.800 137.000 114.100 ;
        RECT 147.800 114.100 148.200 114.200 ;
        RECT 159.800 114.100 160.200 114.200 ;
        RECT 170.200 114.100 170.600 114.200 ;
        RECT 171.800 114.100 172.200 114.200 ;
        RECT 182.200 114.100 182.500 114.800 ;
        RECT 191.000 114.100 191.400 114.200 ;
        RECT 147.800 113.800 191.400 114.100 ;
        RECT 195.800 114.100 196.200 114.200 ;
        RECT 203.800 114.100 204.200 114.200 ;
        RECT 195.800 113.800 204.200 114.100 ;
        RECT 219.800 114.100 220.200 114.200 ;
        RECT 222.200 114.100 222.600 114.200 ;
        RECT 219.800 113.800 222.600 114.100 ;
        RECT 228.600 114.100 229.000 114.200 ;
        RECT 231.800 114.100 232.200 114.200 ;
        RECT 228.600 113.800 232.200 114.100 ;
        RECT 237.400 114.100 237.800 114.200 ;
        RECT 237.400 113.800 241.700 114.100 ;
        RECT 241.400 113.200 241.700 113.800 ;
        RECT 7.000 113.100 7.400 113.200 ;
        RECT 17.400 113.100 17.800 113.200 ;
        RECT 34.200 113.100 34.600 113.200 ;
        RECT 7.000 112.800 34.600 113.100 ;
        RECT 43.800 113.100 44.200 113.200 ;
        RECT 44.600 113.100 45.000 113.200 ;
        RECT 46.200 113.100 46.600 113.200 ;
        RECT 88.600 113.100 89.000 113.200 ;
        RECT 99.800 113.100 100.200 113.200 ;
        RECT 43.800 112.800 83.300 113.100 ;
        RECT 88.600 112.800 100.200 113.100 ;
        RECT 103.800 113.100 104.200 113.200 ;
        RECT 104.600 113.100 105.000 113.200 ;
        RECT 115.000 113.100 115.400 113.200 ;
        RECT 103.800 112.800 115.400 113.100 ;
        RECT 118.200 113.100 118.600 113.200 ;
        RECT 120.600 113.100 121.000 113.200 ;
        RECT 118.200 112.800 121.000 113.100 ;
        RECT 134.200 113.100 134.600 113.200 ;
        RECT 193.400 113.100 193.800 113.200 ;
        RECT 134.200 112.800 193.800 113.100 ;
        RECT 197.400 113.100 197.800 113.200 ;
        RECT 230.200 113.100 230.600 113.200 ;
        RECT 237.400 113.100 237.800 113.200 ;
        RECT 197.400 112.800 237.800 113.100 ;
        RECT 241.400 112.800 241.800 113.200 ;
        RECT 66.200 112.100 66.600 112.200 ;
        RECT 72.600 112.100 73.000 112.200 ;
        RECT 82.200 112.100 82.600 112.200 ;
        RECT 66.200 111.800 82.600 112.100 ;
        RECT 83.000 112.100 83.300 112.800 ;
        RECT 100.600 112.100 101.000 112.200 ;
        RECT 83.000 111.800 101.000 112.100 ;
        RECT 103.800 112.100 104.200 112.200 ;
        RECT 105.400 112.100 105.800 112.200 ;
        RECT 103.800 111.800 105.800 112.100 ;
        RECT 107.800 112.100 108.200 112.200 ;
        RECT 127.800 112.100 128.200 112.200 ;
        RECT 107.800 111.800 128.200 112.100 ;
        RECT 129.400 112.100 129.800 112.200 ;
        RECT 142.200 112.100 142.600 112.200 ;
        RECT 129.400 111.800 142.600 112.100 ;
        RECT 149.400 112.100 149.800 112.200 ;
        RECT 153.400 112.100 153.800 112.200 ;
        RECT 149.400 111.800 153.800 112.100 ;
        RECT 155.000 112.100 155.400 112.200 ;
        RECT 157.400 112.100 157.800 112.200 ;
        RECT 155.000 111.800 157.800 112.100 ;
        RECT 160.600 112.100 161.000 112.200 ;
        RECT 161.400 112.100 161.800 112.200 ;
        RECT 160.600 111.800 161.800 112.100 ;
        RECT 164.600 112.100 165.000 112.200 ;
        RECT 167.000 112.100 167.400 112.200 ;
        RECT 164.600 111.800 167.400 112.100 ;
        RECT 171.000 112.100 171.400 112.200 ;
        RECT 175.800 112.100 176.200 112.200 ;
        RECT 171.000 111.800 176.200 112.100 ;
        RECT 181.400 112.100 181.800 112.200 ;
        RECT 199.000 112.100 199.400 112.200 ;
        RECT 181.400 111.800 199.400 112.100 ;
        RECT 241.400 111.800 241.800 112.200 ;
        RECT 241.400 111.200 241.700 111.800 ;
        RECT 39.800 111.100 40.200 111.200 ;
        RECT 49.400 111.100 49.800 111.200 ;
        RECT 67.000 111.100 67.400 111.200 ;
        RECT 71.000 111.100 71.400 111.200 ;
        RECT 39.800 110.800 71.400 111.100 ;
        RECT 103.800 111.100 104.200 111.200 ;
        RECT 111.000 111.100 111.400 111.200 ;
        RECT 114.200 111.100 114.600 111.200 ;
        RECT 103.800 110.800 114.600 111.100 ;
        RECT 119.800 111.100 120.200 111.200 ;
        RECT 122.200 111.100 122.600 111.200 ;
        RECT 119.800 110.800 122.600 111.100 ;
        RECT 135.800 111.100 136.200 111.200 ;
        RECT 139.800 111.100 140.200 111.200 ;
        RECT 135.800 110.800 140.200 111.100 ;
        RECT 148.600 111.100 149.000 111.200 ;
        RECT 165.400 111.100 165.800 111.200 ;
        RECT 170.200 111.100 170.600 111.200 ;
        RECT 148.600 110.800 170.600 111.100 ;
        RECT 182.200 111.100 182.600 111.200 ;
        RECT 197.400 111.100 197.800 111.200 ;
        RECT 182.200 110.800 197.800 111.100 ;
        RECT 209.400 111.100 209.800 111.200 ;
        RECT 219.000 111.100 219.400 111.200 ;
        RECT 209.400 110.800 219.400 111.100 ;
        RECT 241.400 110.800 241.800 111.200 ;
        RECT 71.800 110.100 72.200 110.200 ;
        RECT 79.000 110.100 79.400 110.200 ;
        RECT 71.800 109.800 79.400 110.100 ;
        RECT 82.200 110.100 82.600 110.200 ;
        RECT 87.000 110.100 87.400 110.200 ;
        RECT 82.200 109.800 87.400 110.100 ;
        RECT 105.400 110.100 105.800 110.200 ;
        RECT 107.800 110.100 108.200 110.200 ;
        RECT 118.200 110.100 118.600 110.200 ;
        RECT 105.400 109.800 118.600 110.100 ;
        RECT 119.000 110.100 119.400 110.200 ;
        RECT 123.000 110.100 123.400 110.200 ;
        RECT 119.000 109.800 123.400 110.100 ;
        RECT 128.600 110.100 129.000 110.200 ;
        RECT 133.400 110.100 133.800 110.200 ;
        RECT 128.600 109.800 133.800 110.100 ;
        RECT 135.000 110.100 135.400 110.200 ;
        RECT 163.800 110.100 164.200 110.200 ;
        RECT 168.600 110.100 169.000 110.200 ;
        RECT 135.000 109.800 169.000 110.100 ;
        RECT 169.400 110.100 169.800 110.200 ;
        RECT 171.000 110.100 171.400 110.200 ;
        RECT 169.400 109.800 171.400 110.100 ;
        RECT 189.400 110.100 189.800 110.200 ;
        RECT 194.200 110.100 194.600 110.200 ;
        RECT 189.400 109.800 194.600 110.100 ;
        RECT 249.400 109.800 249.800 110.200 ;
        RECT 249.400 109.200 249.700 109.800 ;
        RECT 1.400 109.100 1.800 109.200 ;
        RECT 18.200 109.100 18.600 109.200 ;
        RECT 1.400 108.800 18.600 109.100 ;
        RECT 23.000 109.100 23.400 109.200 ;
        RECT 27.800 109.100 28.200 109.200 ;
        RECT 36.600 109.100 37.000 109.200 ;
        RECT 23.000 108.800 37.000 109.100 ;
        RECT 54.200 109.100 54.600 109.200 ;
        RECT 59.000 109.100 59.400 109.200 ;
        RECT 54.200 108.800 59.400 109.100 ;
        RECT 60.600 109.100 61.000 109.200 ;
        RECT 83.000 109.100 83.400 109.200 ;
        RECT 60.600 108.800 83.400 109.100 ;
        RECT 84.600 109.100 85.000 109.200 ;
        RECT 92.600 109.100 93.000 109.200 ;
        RECT 84.600 108.800 93.000 109.100 ;
        RECT 115.000 109.100 115.400 109.200 ;
        RECT 187.800 109.100 188.200 109.200 ;
        RECT 198.200 109.100 198.600 109.200 ;
        RECT 115.000 108.800 198.600 109.100 ;
        RECT 203.000 109.100 203.400 109.200 ;
        RECT 227.000 109.100 227.400 109.200 ;
        RECT 203.000 108.800 227.400 109.100 ;
        RECT 228.600 109.100 229.000 109.200 ;
        RECT 229.400 109.100 229.800 109.200 ;
        RECT 228.600 108.800 229.800 109.100 ;
        RECT 236.600 109.100 237.000 109.200 ;
        RECT 241.400 109.100 241.800 109.200 ;
        RECT 243.800 109.100 244.200 109.200 ;
        RECT 244.600 109.100 245.000 109.200 ;
        RECT 236.600 108.800 245.000 109.100 ;
        RECT 249.400 108.800 249.800 109.200 ;
        RECT 12.600 106.800 13.000 107.200 ;
        RECT 13.400 107.100 13.800 107.200 ;
        RECT 23.000 107.100 23.400 107.200 ;
        RECT 13.400 106.800 23.400 107.100 ;
        RECT 27.000 107.100 27.400 107.200 ;
        RECT 30.200 107.100 30.600 107.200 ;
        RECT 27.000 106.800 30.600 107.100 ;
        RECT 42.200 107.100 42.600 107.200 ;
        RECT 48.600 107.100 49.000 107.200 ;
        RECT 50.200 107.100 50.600 107.200 ;
        RECT 42.200 106.800 50.600 107.100 ;
        RECT 55.000 107.100 55.400 107.200 ;
        RECT 64.600 107.100 65.000 107.200 ;
        RECT 55.000 106.800 65.000 107.100 ;
        RECT 84.600 107.100 85.000 107.200 ;
        RECT 95.000 107.100 95.400 107.200 ;
        RECT 97.400 107.100 97.800 107.200 ;
        RECT 134.200 107.100 134.600 107.200 ;
        RECT 183.000 107.100 183.400 107.200 ;
        RECT 210.200 107.100 210.600 107.200 ;
        RECT 84.600 106.800 210.600 107.100 ;
        RECT 215.000 106.800 215.400 107.200 ;
        RECT 218.200 107.100 218.600 107.200 ;
        RECT 223.800 107.100 224.200 107.200 ;
        RECT 225.400 107.100 225.800 107.200 ;
        RECT 218.200 106.800 225.800 107.100 ;
        RECT 227.800 107.100 228.200 107.200 ;
        RECT 237.400 107.100 237.800 107.200 ;
        RECT 239.000 107.100 239.400 107.200 ;
        RECT 227.800 106.800 239.400 107.100 ;
        RECT 243.800 106.800 244.200 107.200 ;
        RECT 12.600 106.200 12.900 106.800 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 19.000 106.100 19.400 106.300 ;
        RECT 24.600 106.100 25.000 106.200 ;
        RECT 19.000 105.800 25.000 106.100 ;
        RECT 43.800 106.100 44.200 106.200 ;
        RECT 63.800 106.100 64.200 106.200 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 43.800 105.800 69.000 106.100 ;
        RECT 72.600 106.100 73.000 106.200 ;
        RECT 79.000 106.100 79.400 106.200 ;
        RECT 72.600 105.800 79.400 106.100 ;
        RECT 86.200 106.100 86.600 106.200 ;
        RECT 91.800 106.100 92.200 106.200 ;
        RECT 103.800 106.100 104.200 106.200 ;
        RECT 86.200 105.800 104.200 106.100 ;
        RECT 105.400 106.100 105.800 106.200 ;
        RECT 108.600 106.100 109.000 106.200 ;
        RECT 123.800 106.100 124.200 106.200 ;
        RECT 105.400 105.800 124.200 106.100 ;
        RECT 132.600 106.100 133.000 106.200 ;
        RECT 196.600 106.100 197.000 106.200 ;
        RECT 199.800 106.100 200.200 106.200 ;
        RECT 132.600 105.800 200.200 106.100 ;
        RECT 200.600 106.100 201.000 106.200 ;
        RECT 201.400 106.100 201.800 106.200 ;
        RECT 200.600 105.800 201.800 106.100 ;
        RECT 207.800 105.800 208.200 106.200 ;
        RECT 211.800 106.100 212.200 106.200 ;
        RECT 215.000 106.100 215.300 106.800 ;
        RECT 243.800 106.200 244.100 106.800 ;
        RECT 211.800 105.800 215.300 106.100 ;
        RECT 219.800 106.100 220.200 106.200 ;
        RECT 231.800 106.100 232.200 106.200 ;
        RECT 235.800 106.100 236.200 106.200 ;
        RECT 219.800 105.800 236.200 106.100 ;
        RECT 240.600 106.100 241.000 106.200 ;
        RECT 243.800 106.100 244.200 106.200 ;
        RECT 240.600 105.800 244.200 106.100 ;
        RECT 244.600 106.100 245.000 106.200 ;
        RECT 247.800 106.100 248.200 106.200 ;
        RECT 244.600 105.800 248.200 106.100 ;
        RECT 207.800 105.200 208.100 105.800 ;
        RECT 60.600 105.100 61.000 105.200 ;
        RECT 66.200 105.100 66.600 105.200 ;
        RECT 60.600 104.800 66.600 105.100 ;
        RECT 70.200 105.100 70.600 105.200 ;
        RECT 72.600 105.100 73.000 105.200 ;
        RECT 73.400 105.100 73.800 105.200 ;
        RECT 70.200 104.800 73.800 105.100 ;
        RECT 97.400 105.100 97.800 105.200 ;
        RECT 98.200 105.100 98.600 105.200 ;
        RECT 97.400 104.800 98.600 105.100 ;
        RECT 100.600 105.100 101.000 105.200 ;
        RECT 103.000 105.100 103.400 105.200 ;
        RECT 107.000 105.100 107.400 105.200 ;
        RECT 100.600 104.800 107.400 105.100 ;
        RECT 109.400 105.100 109.800 105.200 ;
        RECT 110.200 105.100 110.600 105.200 ;
        RECT 109.400 104.800 110.600 105.100 ;
        RECT 111.800 105.100 112.200 105.200 ;
        RECT 123.800 105.100 124.200 105.200 ;
        RECT 127.000 105.100 127.400 105.200 ;
        RECT 111.800 104.800 127.400 105.100 ;
        RECT 131.000 105.100 131.400 105.200 ;
        RECT 131.800 105.100 132.200 105.200 ;
        RECT 131.000 104.800 132.200 105.100 ;
        RECT 133.400 105.100 133.800 105.200 ;
        RECT 136.600 105.100 137.000 105.200 ;
        RECT 133.400 104.800 137.000 105.100 ;
        RECT 142.200 105.100 142.600 105.200 ;
        RECT 143.800 105.100 144.200 105.200 ;
        RECT 142.200 104.800 144.200 105.100 ;
        RECT 155.800 105.100 156.200 105.200 ;
        RECT 159.000 105.100 159.400 105.200 ;
        RECT 155.800 104.800 159.400 105.100 ;
        RECT 162.200 104.800 162.600 105.200 ;
        RECT 165.400 105.100 165.800 105.200 ;
        RECT 169.400 105.100 169.800 105.200 ;
        RECT 165.400 104.800 169.800 105.100 ;
        RECT 171.000 105.100 171.400 105.200 ;
        RECT 172.600 105.100 173.000 105.200 ;
        RECT 171.000 104.800 173.000 105.100 ;
        RECT 177.400 105.100 177.800 105.200 ;
        RECT 191.000 105.100 191.400 105.200 ;
        RECT 177.400 104.800 191.400 105.100 ;
        RECT 207.800 104.800 208.200 105.200 ;
        RECT 211.000 105.100 211.400 105.200 ;
        RECT 215.000 105.100 215.400 105.200 ;
        RECT 211.000 104.800 215.400 105.100 ;
        RECT 215.800 105.100 216.200 105.200 ;
        RECT 229.400 105.100 229.800 105.200 ;
        RECT 230.200 105.100 230.600 105.200 ;
        RECT 215.800 104.800 227.300 105.100 ;
        RECT 229.400 104.800 230.600 105.100 ;
        RECT 23.000 104.100 23.400 104.200 ;
        RECT 24.600 104.100 25.000 104.200 ;
        RECT 27.000 104.100 27.400 104.200 ;
        RECT 55.800 104.100 56.200 104.200 ;
        RECT 23.000 103.800 56.200 104.100 ;
        RECT 101.400 104.100 101.800 104.200 ;
        RECT 106.200 104.100 106.600 104.200 ;
        RECT 120.600 104.100 121.000 104.200 ;
        RECT 101.400 103.800 121.000 104.100 ;
        RECT 134.200 104.100 134.600 104.200 ;
        RECT 135.000 104.100 135.400 104.200 ;
        RECT 134.200 103.800 135.400 104.100 ;
        RECT 140.600 104.100 141.000 104.200 ;
        RECT 157.400 104.100 157.800 104.200 ;
        RECT 140.600 103.800 157.800 104.100 ;
        RECT 162.200 104.100 162.500 104.800 ;
        RECT 227.000 104.200 227.300 104.800 ;
        RECT 165.400 104.100 165.800 104.200 ;
        RECT 162.200 103.800 165.800 104.100 ;
        RECT 167.000 104.100 167.400 104.200 ;
        RECT 200.600 104.100 201.000 104.200 ;
        RECT 167.000 103.800 201.000 104.100 ;
        RECT 207.800 104.100 208.200 104.200 ;
        RECT 208.600 104.100 209.000 104.200 ;
        RECT 218.200 104.100 218.600 104.200 ;
        RECT 207.800 103.800 218.600 104.100 ;
        RECT 219.800 104.100 220.200 104.200 ;
        RECT 222.200 104.100 222.600 104.200 ;
        RECT 224.600 104.100 225.000 104.200 ;
        RECT 219.800 103.800 225.000 104.100 ;
        RECT 227.000 103.800 227.400 104.200 ;
        RECT 230.200 104.100 230.600 104.200 ;
        RECT 231.800 104.100 232.200 104.200 ;
        RECT 230.200 103.800 232.200 104.100 ;
        RECT 22.200 103.100 22.600 103.200 ;
        RECT 59.000 103.100 59.400 103.200 ;
        RECT 67.800 103.100 68.200 103.200 ;
        RECT 22.200 102.800 68.200 103.100 ;
        RECT 89.400 103.100 89.800 103.200 ;
        RECT 118.200 103.100 118.600 103.200 ;
        RECT 89.400 102.800 118.600 103.100 ;
        RECT 119.000 103.100 119.400 103.200 ;
        RECT 129.400 103.100 129.800 103.200 ;
        RECT 119.000 102.800 129.800 103.100 ;
        RECT 147.000 103.100 147.400 103.200 ;
        RECT 155.800 103.100 156.200 103.200 ;
        RECT 156.600 103.100 157.000 103.200 ;
        RECT 171.800 103.100 172.200 103.200 ;
        RECT 181.400 103.100 181.800 103.200 ;
        RECT 147.000 102.800 157.000 103.100 ;
        RECT 171.000 102.800 181.800 103.100 ;
        RECT 205.400 103.100 205.800 103.200 ;
        RECT 211.000 103.100 211.400 103.200 ;
        RECT 205.400 102.800 211.400 103.100 ;
        RECT 226.200 103.100 226.600 103.200 ;
        RECT 248.600 103.100 249.000 103.200 ;
        RECT 226.200 102.800 249.000 103.100 ;
        RECT 39.000 102.100 39.400 102.200 ;
        RECT 41.400 102.100 41.800 102.200 ;
        RECT 61.400 102.100 61.800 102.200 ;
        RECT 39.000 101.800 61.800 102.100 ;
        RECT 75.800 102.100 76.200 102.200 ;
        RECT 106.200 102.100 106.600 102.200 ;
        RECT 75.800 101.800 106.600 102.100 ;
        RECT 107.800 102.100 108.200 102.200 ;
        RECT 112.600 102.100 113.000 102.200 ;
        RECT 115.000 102.100 115.400 102.200 ;
        RECT 107.800 101.800 115.400 102.100 ;
        RECT 122.200 102.100 122.600 102.200 ;
        RECT 176.600 102.100 177.000 102.200 ;
        RECT 184.600 102.100 185.000 102.200 ;
        RECT 122.200 101.800 185.000 102.100 ;
        RECT 188.600 102.100 189.000 102.200 ;
        RECT 209.400 102.100 209.800 102.200 ;
        RECT 212.600 102.100 213.000 102.200 ;
        RECT 188.600 101.800 213.000 102.100 ;
        RECT 215.800 102.100 216.200 102.200 ;
        RECT 220.600 102.100 221.000 102.200 ;
        RECT 215.800 101.800 221.000 102.100 ;
        RECT 89.400 101.100 89.800 101.200 ;
        RECT 95.000 101.100 95.400 101.200 ;
        RECT 89.400 100.800 95.400 101.100 ;
        RECT 114.200 101.100 114.600 101.200 ;
        RECT 130.200 101.100 130.600 101.200 ;
        RECT 114.200 100.800 130.600 101.100 ;
        RECT 155.000 101.100 155.400 101.200 ;
        RECT 159.800 101.100 160.200 101.200 ;
        RECT 155.000 100.800 160.200 101.100 ;
        RECT 207.800 101.100 208.200 101.200 ;
        RECT 209.400 101.100 209.800 101.200 ;
        RECT 207.800 100.800 209.800 101.100 ;
        RECT 221.400 101.100 221.800 101.200 ;
        RECT 230.200 101.100 230.600 101.200 ;
        RECT 221.400 100.800 230.600 101.100 ;
        RECT 82.200 100.100 82.600 100.200 ;
        RECT 83.800 100.100 84.200 100.200 ;
        RECT 82.200 99.800 84.200 100.100 ;
        RECT 90.200 100.100 90.600 100.200 ;
        RECT 93.400 100.100 93.800 100.200 ;
        RECT 90.200 99.800 93.800 100.100 ;
        RECT 95.000 100.100 95.400 100.200 ;
        RECT 95.800 100.100 96.200 100.200 ;
        RECT 95.000 99.800 96.200 100.100 ;
        RECT 96.600 100.100 97.000 100.200 ;
        RECT 111.000 100.100 111.400 100.200 ;
        RECT 96.600 99.800 111.400 100.100 ;
        RECT 116.600 100.100 117.000 100.200 ;
        RECT 125.400 100.100 125.800 100.200 ;
        RECT 116.600 99.800 125.800 100.100 ;
        RECT 170.200 100.100 170.600 100.200 ;
        RECT 181.400 100.100 181.800 100.200 ;
        RECT 170.200 99.800 181.800 100.100 ;
        RECT 210.200 100.100 210.600 100.200 ;
        RECT 214.200 100.100 214.600 100.200 ;
        RECT 215.800 100.100 216.200 100.200 ;
        RECT 210.200 99.800 216.200 100.100 ;
        RECT 47.000 99.100 47.400 99.200 ;
        RECT 80.600 99.100 81.000 99.200 ;
        RECT 47.000 98.800 81.000 99.100 ;
        RECT 83.800 99.100 84.200 99.200 ;
        RECT 87.000 99.100 87.400 99.200 ;
        RECT 99.800 99.100 100.200 99.200 ;
        RECT 113.400 99.100 113.800 99.200 ;
        RECT 83.800 98.800 113.800 99.100 ;
        RECT 118.200 99.100 118.600 99.200 ;
        RECT 121.400 99.100 121.800 99.200 ;
        RECT 138.200 99.100 138.600 99.200 ;
        RECT 173.400 99.100 173.800 99.200 ;
        RECT 118.200 98.800 173.800 99.100 ;
        RECT 179.800 99.100 180.200 99.200 ;
        RECT 184.600 99.100 185.000 99.200 ;
        RECT 210.200 99.100 210.600 99.200 ;
        RECT 179.800 98.800 210.600 99.100 ;
        RECT 2.200 98.100 2.600 98.200 ;
        RECT 42.200 98.100 42.600 98.200 ;
        RECT 98.200 98.100 98.600 98.200 ;
        RECT 2.200 97.800 98.600 98.100 ;
        RECT 127.000 98.100 127.400 98.200 ;
        RECT 191.000 98.100 191.400 98.200 ;
        RECT 193.400 98.100 193.800 98.200 ;
        RECT 195.800 98.100 196.200 98.200 ;
        RECT 127.000 97.800 196.200 98.100 ;
        RECT 23.000 97.100 23.400 97.200 ;
        RECT 27.800 97.100 28.200 97.200 ;
        RECT 23.000 96.800 28.200 97.100 ;
        RECT 30.200 97.100 30.600 97.200 ;
        RECT 34.200 97.100 34.600 97.200 ;
        RECT 45.400 97.100 45.800 97.200 ;
        RECT 30.200 96.800 45.800 97.100 ;
        RECT 55.000 97.100 55.400 97.200 ;
        RECT 67.800 97.100 68.200 97.200 ;
        RECT 70.200 97.100 70.600 97.200 ;
        RECT 96.600 97.100 97.000 97.200 ;
        RECT 55.000 96.800 66.500 97.100 ;
        RECT 67.800 96.800 97.000 97.100 ;
        RECT 99.800 97.100 100.200 97.200 ;
        RECT 111.800 97.100 112.200 97.200 ;
        RECT 119.000 97.100 119.400 97.200 ;
        RECT 99.800 96.800 119.400 97.100 ;
        RECT 156.600 97.100 157.000 97.200 ;
        RECT 178.200 97.100 178.600 97.200 ;
        RECT 156.600 96.800 178.600 97.100 ;
        RECT 187.000 97.100 187.400 97.200 ;
        RECT 205.400 97.100 205.800 97.200 ;
        RECT 187.000 96.800 205.800 97.100 ;
        RECT 20.600 96.100 21.000 96.200 ;
        RECT 22.200 96.100 22.600 96.200 ;
        RECT 20.600 95.800 22.600 96.100 ;
        RECT 26.200 96.100 26.600 96.200 ;
        RECT 27.800 96.100 28.200 96.200 ;
        RECT 29.400 96.100 29.800 96.200 ;
        RECT 33.400 96.100 33.800 96.200 ;
        RECT 26.200 95.800 29.800 96.100 ;
        RECT 31.800 95.800 33.800 96.100 ;
        RECT 60.600 96.100 61.000 96.200 ;
        RECT 62.200 96.100 62.600 96.200 ;
        RECT 65.400 96.100 65.800 96.200 ;
        RECT 60.600 95.800 65.800 96.100 ;
        RECT 66.200 96.100 66.500 96.800 ;
        RECT 68.600 96.100 69.000 96.200 ;
        RECT 66.200 95.800 69.000 96.100 ;
        RECT 90.200 96.100 90.600 96.200 ;
        RECT 95.800 96.100 96.200 96.200 ;
        RECT 103.000 96.100 103.400 96.200 ;
        RECT 111.800 96.100 112.200 96.200 ;
        RECT 90.200 95.800 112.200 96.100 ;
        RECT 117.400 96.100 117.800 96.200 ;
        RECT 132.600 96.100 133.000 96.200 ;
        RECT 135.000 96.100 135.400 96.200 ;
        RECT 117.400 95.800 135.400 96.100 ;
        RECT 157.400 96.100 157.800 96.200 ;
        RECT 172.600 96.100 173.000 96.200 ;
        RECT 157.400 95.800 173.000 96.100 ;
        RECT 173.400 96.100 173.800 96.200 ;
        RECT 187.800 96.100 188.200 96.200 ;
        RECT 173.400 95.800 188.200 96.100 ;
        RECT 204.600 95.800 205.000 96.200 ;
        RECT 220.600 96.100 221.000 96.200 ;
        RECT 227.000 96.100 227.400 96.200 ;
        RECT 220.600 95.800 227.400 96.100 ;
        RECT 231.800 96.100 232.200 96.200 ;
        RECT 237.400 96.100 237.800 96.200 ;
        RECT 231.800 95.800 237.800 96.100 ;
        RECT 242.200 96.100 242.600 96.200 ;
        RECT 243.000 96.100 243.400 96.200 ;
        RECT 243.800 96.100 244.200 96.200 ;
        RECT 242.200 95.800 244.200 96.100 ;
        RECT 31.800 95.200 32.100 95.800 ;
        RECT 157.400 95.200 157.700 95.800 ;
        RECT 3.000 94.800 3.400 95.200 ;
        RECT 7.800 95.100 8.200 95.200 ;
        RECT 19.800 95.100 20.200 95.200 ;
        RECT 7.800 94.800 20.200 95.100 ;
        RECT 31.800 94.800 32.200 95.200 ;
        RECT 52.600 94.800 53.000 95.200 ;
        RECT 60.600 95.100 61.000 95.200 ;
        RECT 67.800 95.100 68.200 95.200 ;
        RECT 60.600 94.800 68.200 95.100 ;
        RECT 69.400 95.100 69.800 95.200 ;
        RECT 71.800 95.100 72.200 95.200 ;
        RECT 69.400 94.800 72.200 95.100 ;
        RECT 74.200 95.100 74.600 95.200 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 74.200 94.800 78.600 95.100 ;
        RECT 85.400 95.100 85.800 95.200 ;
        RECT 95.800 95.100 96.200 95.200 ;
        RECT 85.400 94.800 96.200 95.100 ;
        RECT 96.600 95.100 97.000 95.200 ;
        RECT 101.400 95.100 101.800 95.200 ;
        RECT 96.600 94.800 101.800 95.100 ;
        RECT 102.200 95.100 102.600 95.200 ;
        RECT 119.800 95.100 120.200 95.200 ;
        RECT 120.600 95.100 121.000 95.200 ;
        RECT 102.200 94.800 107.400 95.100 ;
        RECT 119.800 94.800 121.000 95.100 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 175.000 95.100 175.400 95.200 ;
        RECT 183.000 95.100 183.400 95.200 ;
        RECT 191.000 95.100 191.400 95.200 ;
        RECT 175.000 94.800 183.400 95.100 ;
        RECT 186.200 94.800 191.400 95.100 ;
        RECT 200.600 95.100 201.000 95.200 ;
        RECT 204.600 95.100 204.900 95.800 ;
        RECT 200.600 94.800 204.900 95.100 ;
        RECT 213.400 95.100 213.800 95.200 ;
        RECT 215.800 95.100 216.200 95.200 ;
        RECT 213.400 94.800 216.200 95.100 ;
        RECT 222.200 95.100 222.600 95.200 ;
        RECT 231.000 95.100 231.400 95.200 ;
        RECT 232.600 95.100 233.000 95.200 ;
        RECT 222.200 94.800 233.000 95.100 ;
        RECT 235.000 95.100 235.400 95.200 ;
        RECT 243.000 95.100 243.400 95.200 ;
        RECT 246.200 95.100 246.600 95.200 ;
        RECT 235.000 94.800 246.600 95.100 ;
        RECT 3.000 94.100 3.300 94.800 ;
        RECT 11.000 94.100 11.400 94.200 ;
        RECT 3.000 93.800 11.400 94.100 ;
        RECT 12.600 94.100 13.000 94.200 ;
        RECT 16.600 94.100 17.000 94.200 ;
        RECT 18.200 94.100 18.600 94.200 ;
        RECT 12.600 93.800 18.600 94.100 ;
        RECT 24.600 94.100 25.000 94.200 ;
        RECT 30.200 94.100 30.600 94.200 ;
        RECT 24.600 93.800 30.600 94.100 ;
        RECT 31.000 94.100 31.400 94.200 ;
        RECT 35.000 94.100 35.400 94.200 ;
        RECT 31.000 93.800 35.400 94.100 ;
        RECT 38.200 94.100 38.600 94.200 ;
        RECT 52.600 94.100 52.900 94.800 ;
        RECT 107.000 94.700 107.400 94.800 ;
        RECT 98.200 94.100 98.600 94.200 ;
        RECT 101.400 94.100 101.800 94.200 ;
        RECT 38.200 93.800 76.100 94.100 ;
        RECT 98.200 93.800 101.800 94.100 ;
        RECT 102.200 94.100 102.600 94.200 ;
        RECT 103.000 94.100 103.400 94.200 ;
        RECT 102.200 93.800 103.400 94.100 ;
        RECT 112.600 94.100 113.000 94.200 ;
        RECT 115.000 94.100 115.400 94.200 ;
        RECT 112.600 93.800 115.400 94.100 ;
        RECT 123.800 94.100 124.200 94.400 ;
        RECT 186.200 94.200 186.500 94.800 ;
        RECT 134.200 94.100 134.600 94.200 ;
        RECT 139.000 94.100 139.400 94.200 ;
        RECT 123.800 93.800 139.400 94.100 ;
        RECT 139.800 93.800 140.200 94.200 ;
        RECT 141.400 94.100 141.800 94.200 ;
        RECT 155.800 94.100 156.200 94.200 ;
        RECT 175.000 94.100 175.400 94.200 ;
        RECT 141.400 93.800 175.400 94.100 ;
        RECT 186.200 93.800 186.600 94.200 ;
        RECT 195.800 94.100 196.200 94.200 ;
        RECT 206.200 94.100 206.600 94.200 ;
        RECT 195.800 93.800 206.600 94.100 ;
        RECT 223.000 94.100 223.400 94.200 ;
        RECT 226.200 94.100 226.600 94.200 ;
        RECT 223.000 93.800 226.600 94.100 ;
        RECT 233.400 94.100 233.800 94.200 ;
        RECT 247.000 94.100 247.400 94.200 ;
        RECT 247.800 94.100 248.200 94.200 ;
        RECT 233.400 93.800 248.200 94.100 ;
        RECT 75.800 93.200 76.100 93.800 ;
        RECT 0.600 93.100 1.000 93.200 ;
        RECT 7.800 93.100 8.200 93.200 ;
        RECT 0.600 92.800 8.200 93.100 ;
        RECT 15.000 93.100 15.400 93.200 ;
        RECT 46.200 93.100 46.600 93.200 ;
        RECT 15.000 92.800 46.600 93.100 ;
        RECT 75.800 92.800 76.200 93.200 ;
        RECT 87.800 93.100 88.200 93.200 ;
        RECT 107.800 93.100 108.200 93.200 ;
        RECT 87.800 92.800 108.200 93.100 ;
        RECT 117.400 93.100 117.800 93.200 ;
        RECT 125.400 93.100 125.800 93.200 ;
        RECT 117.400 92.800 125.800 93.100 ;
        RECT 128.600 93.100 129.000 93.200 ;
        RECT 131.800 93.100 132.200 93.200 ;
        RECT 128.600 92.800 132.200 93.100 ;
        RECT 137.400 93.100 137.800 93.200 ;
        RECT 139.800 93.100 140.100 93.800 ;
        RECT 137.400 92.800 140.100 93.100 ;
        RECT 143.000 93.100 143.400 93.200 ;
        RECT 179.800 93.100 180.200 93.200 ;
        RECT 183.800 93.100 184.200 93.200 ;
        RECT 189.400 93.100 189.800 93.200 ;
        RECT 143.000 92.800 174.500 93.100 ;
        RECT 179.800 92.800 189.800 93.100 ;
        RECT 38.200 92.100 38.600 92.200 ;
        RECT 40.600 92.100 41.000 92.200 ;
        RECT 38.200 91.800 41.000 92.100 ;
        RECT 43.000 92.100 43.400 92.200 ;
        RECT 49.400 92.100 49.800 92.200 ;
        RECT 43.000 91.800 49.800 92.100 ;
        RECT 80.600 92.100 81.000 92.200 ;
        RECT 84.600 92.100 85.000 92.200 ;
        RECT 80.600 91.800 85.000 92.100 ;
        RECT 93.400 92.100 93.800 92.200 ;
        RECT 96.600 92.100 97.000 92.200 ;
        RECT 93.400 91.800 97.000 92.100 ;
        RECT 106.200 92.100 106.600 92.200 ;
        RECT 122.200 92.100 122.600 92.200 ;
        RECT 106.200 91.800 122.600 92.100 ;
        RECT 126.200 92.100 126.600 92.200 ;
        RECT 146.200 92.100 146.600 92.200 ;
        RECT 126.200 91.800 146.600 92.100 ;
        RECT 174.200 92.100 174.500 92.800 ;
        RECT 183.800 92.100 184.200 92.200 ;
        RECT 185.400 92.100 185.800 92.200 ;
        RECT 174.200 91.800 185.800 92.100 ;
        RECT 186.200 92.100 186.600 92.200 ;
        RECT 203.800 92.100 204.200 92.200 ;
        RECT 186.200 91.800 204.200 92.100 ;
        RECT 222.200 92.100 222.600 92.200 ;
        RECT 234.200 92.100 234.600 92.200 ;
        RECT 243.000 92.100 243.400 92.200 ;
        RECT 222.200 91.800 243.400 92.100 ;
        RECT 45.400 91.100 45.800 91.200 ;
        RECT 64.600 91.100 65.000 91.200 ;
        RECT 45.400 90.800 65.000 91.100 ;
        RECT 102.200 91.100 102.600 91.200 ;
        RECT 114.200 91.100 114.600 91.200 ;
        RECT 102.200 90.800 114.600 91.100 ;
        RECT 116.600 91.100 117.000 91.200 ;
        RECT 132.600 91.100 133.000 91.200 ;
        RECT 116.600 90.800 133.000 91.100 ;
        RECT 133.400 91.100 133.800 91.200 ;
        RECT 147.000 91.100 147.400 91.200 ;
        RECT 133.400 90.800 147.400 91.100 ;
        RECT 159.000 91.100 159.400 91.200 ;
        RECT 159.800 91.100 160.200 91.200 ;
        RECT 159.000 90.800 160.200 91.100 ;
        RECT 177.400 91.100 177.800 91.200 ;
        RECT 198.200 91.100 198.600 91.200 ;
        RECT 177.400 90.800 198.600 91.100 ;
        RECT 208.600 91.100 209.000 91.200 ;
        RECT 229.400 91.100 229.800 91.200 ;
        RECT 231.000 91.100 231.400 91.200 ;
        RECT 208.600 90.800 231.400 91.100 ;
        RECT 87.000 90.100 87.400 90.200 ;
        RECT 96.600 90.100 97.000 90.200 ;
        RECT 87.000 89.800 97.000 90.100 ;
        RECT 115.800 90.100 116.200 90.200 ;
        RECT 117.400 90.100 117.800 90.200 ;
        RECT 115.800 89.800 117.800 90.100 ;
        RECT 120.600 90.100 121.000 90.200 ;
        RECT 127.800 90.100 128.200 90.200 ;
        RECT 120.600 89.800 128.200 90.100 ;
        RECT 129.400 90.100 129.800 90.200 ;
        RECT 132.600 90.100 133.000 90.200 ;
        RECT 143.000 90.100 143.400 90.200 ;
        RECT 129.400 89.800 143.400 90.100 ;
        RECT 146.200 90.100 146.600 90.200 ;
        RECT 166.200 90.100 166.600 90.200 ;
        RECT 146.200 89.800 166.600 90.100 ;
        RECT 230.200 90.100 230.600 90.200 ;
        RECT 240.600 90.100 241.000 90.200 ;
        RECT 230.200 89.800 241.000 90.100 ;
        RECT 20.600 89.100 21.000 89.200 ;
        RECT 23.800 89.100 24.200 89.200 ;
        RECT 20.600 88.800 24.200 89.100 ;
        RECT 41.400 89.100 41.800 89.200 ;
        RECT 60.600 89.100 61.000 89.200 ;
        RECT 64.600 89.100 65.000 89.200 ;
        RECT 41.400 88.800 45.700 89.100 ;
        RECT 60.600 88.800 65.000 89.100 ;
        RECT 81.400 89.100 81.800 89.200 ;
        RECT 87.800 89.100 88.200 89.200 ;
        RECT 81.400 88.800 88.200 89.100 ;
        RECT 94.200 89.100 94.600 89.200 ;
        RECT 97.400 89.100 97.800 89.200 ;
        RECT 103.000 89.100 103.400 89.200 ;
        RECT 94.200 88.800 103.400 89.100 ;
        RECT 111.000 89.100 111.400 89.200 ;
        RECT 116.600 89.100 117.000 89.200 ;
        RECT 111.000 88.800 117.000 89.100 ;
        RECT 122.200 89.100 122.600 89.200 ;
        RECT 123.000 89.100 123.400 89.200 ;
        RECT 135.800 89.100 136.200 89.200 ;
        RECT 158.200 89.100 158.600 89.200 ;
        RECT 122.200 88.800 158.600 89.100 ;
        RECT 159.800 89.100 160.200 89.200 ;
        RECT 164.600 89.100 165.000 89.200 ;
        RECT 159.800 88.800 165.000 89.100 ;
        RECT 165.400 89.100 165.800 89.200 ;
        RECT 170.200 89.100 170.600 89.200 ;
        RECT 165.400 88.800 170.600 89.100 ;
        RECT 175.000 89.100 175.400 89.200 ;
        RECT 196.600 89.100 197.000 89.200 ;
        RECT 207.800 89.100 208.200 89.200 ;
        RECT 175.000 88.800 208.200 89.100 ;
        RECT 226.200 89.100 226.600 89.200 ;
        RECT 239.800 89.100 240.200 89.200 ;
        RECT 226.200 88.800 240.200 89.100 ;
        RECT 251.000 88.800 251.400 89.200 ;
        RECT 45.400 88.200 45.700 88.800 ;
        RECT 251.000 88.200 251.300 88.800 ;
        RECT 6.200 88.100 6.600 88.200 ;
        RECT 11.000 88.100 11.400 88.200 ;
        RECT 23.000 88.100 23.400 88.200 ;
        RECT 35.000 88.100 35.400 88.200 ;
        RECT 6.200 87.800 35.400 88.100 ;
        RECT 45.400 87.800 45.800 88.200 ;
        RECT 55.000 87.800 55.400 88.200 ;
        RECT 55.800 88.100 56.200 88.200 ;
        RECT 58.200 88.100 58.600 88.200 ;
        RECT 90.200 88.100 90.600 88.200 ;
        RECT 55.800 87.800 90.600 88.100 ;
        RECT 103.000 88.100 103.400 88.200 ;
        RECT 115.000 88.100 115.400 88.200 ;
        RECT 125.400 88.100 125.800 88.200 ;
        RECT 127.000 88.100 127.400 88.200 ;
        RECT 127.800 88.100 128.200 88.200 ;
        RECT 103.000 87.800 128.200 88.100 ;
        RECT 129.400 88.100 129.800 88.200 ;
        RECT 141.400 88.100 141.800 88.200 ;
        RECT 129.400 87.800 141.800 88.100 ;
        RECT 148.600 88.100 149.000 88.200 ;
        RECT 151.800 88.100 152.200 88.200 ;
        RECT 148.600 87.800 152.200 88.100 ;
        RECT 159.000 88.100 159.400 88.200 ;
        RECT 159.800 88.100 160.200 88.200 ;
        RECT 159.000 87.800 160.200 88.100 ;
        RECT 188.600 88.100 189.000 88.200 ;
        RECT 212.600 88.100 213.000 88.200 ;
        RECT 232.600 88.100 233.000 88.200 ;
        RECT 188.600 87.800 209.700 88.100 ;
        RECT 212.600 87.800 233.000 88.100 ;
        RECT 241.400 88.100 241.800 88.200 ;
        RECT 247.000 88.100 247.400 88.200 ;
        RECT 241.400 87.800 247.400 88.100 ;
        RECT 251.000 87.800 251.400 88.200 ;
        RECT 29.400 87.100 29.800 87.200 ;
        RECT 44.600 87.100 45.000 87.200 ;
        RECT 55.000 87.100 55.300 87.800 ;
        RECT 71.000 87.100 71.400 87.200 ;
        RECT 85.400 87.100 85.800 87.200 ;
        RECT 87.800 87.100 88.200 87.200 ;
        RECT 29.400 86.800 71.400 87.100 ;
        RECT 73.400 86.800 75.300 87.100 ;
        RECT 85.400 86.800 88.200 87.100 ;
        RECT 95.800 87.100 96.200 87.200 ;
        RECT 96.600 87.100 97.000 87.200 ;
        RECT 95.800 86.800 97.000 87.100 ;
        RECT 114.200 87.100 114.600 87.200 ;
        RECT 119.800 87.100 120.200 87.200 ;
        RECT 114.200 86.800 120.200 87.100 ;
        RECT 120.600 86.800 121.000 87.200 ;
        RECT 124.600 87.100 125.000 87.200 ;
        RECT 129.400 87.100 129.800 87.200 ;
        RECT 131.000 87.100 131.400 87.200 ;
        RECT 124.600 86.800 131.400 87.100 ;
        RECT 134.200 86.800 134.600 87.200 ;
        RECT 140.600 87.100 141.000 87.200 ;
        RECT 150.200 87.100 150.600 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 140.600 86.800 160.200 87.100 ;
        RECT 163.800 87.100 164.200 87.200 ;
        RECT 165.400 87.100 165.800 87.200 ;
        RECT 163.800 86.800 165.800 87.100 ;
        RECT 168.600 87.100 169.000 87.200 ;
        RECT 170.200 87.100 170.600 87.200 ;
        RECT 168.600 86.800 170.600 87.100 ;
        RECT 171.000 87.100 171.400 87.200 ;
        RECT 180.600 87.100 181.000 87.200 ;
        RECT 171.000 86.800 181.000 87.100 ;
        RECT 190.200 87.100 190.600 87.200 ;
        RECT 191.800 87.100 192.200 87.200 ;
        RECT 190.200 86.800 192.200 87.100 ;
        RECT 194.200 87.100 194.600 87.200 ;
        RECT 203.000 87.100 203.400 87.200 ;
        RECT 205.400 87.100 205.800 87.200 ;
        RECT 208.600 87.100 209.000 87.200 ;
        RECT 194.200 86.800 209.000 87.100 ;
        RECT 209.400 87.100 209.700 87.800 ;
        RECT 241.400 87.200 241.700 87.800 ;
        RECT 214.200 87.100 214.600 87.200 ;
        RECT 209.400 86.800 214.600 87.100 ;
        RECT 217.400 87.100 217.800 87.200 ;
        RECT 219.800 87.100 220.200 87.200 ;
        RECT 217.400 86.800 220.200 87.100 ;
        RECT 241.400 86.800 241.800 87.200 ;
        RECT 247.000 87.100 247.400 87.200 ;
        RECT 250.200 87.100 250.600 87.200 ;
        RECT 247.000 86.800 250.600 87.100 ;
        RECT 73.400 86.200 73.700 86.800 ;
        RECT 75.000 86.200 75.300 86.800 ;
        RECT 33.400 85.800 33.800 86.200 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 35.800 86.100 36.200 86.200 ;
        RECT 38.200 86.100 38.600 86.200 ;
        RECT 35.800 85.800 38.600 86.100 ;
        RECT 40.600 86.100 41.000 86.200 ;
        RECT 60.600 86.100 61.000 86.200 ;
        RECT 40.600 85.800 61.000 86.100 ;
        RECT 64.600 86.100 65.000 86.200 ;
        RECT 65.400 86.100 65.800 86.200 ;
        RECT 64.600 85.800 65.800 86.100 ;
        RECT 73.400 85.800 73.800 86.200 ;
        RECT 75.000 86.100 75.400 86.200 ;
        RECT 80.600 86.100 81.000 86.200 ;
        RECT 75.000 85.800 81.000 86.100 ;
        RECT 88.600 86.100 89.000 86.200 ;
        RECT 91.000 86.100 91.400 86.200 ;
        RECT 88.600 85.800 91.400 86.100 ;
        RECT 92.600 86.100 93.000 86.200 ;
        RECT 94.200 86.100 94.600 86.200 ;
        RECT 95.800 86.100 96.200 86.200 ;
        RECT 92.600 85.800 96.200 86.100 ;
        RECT 115.800 86.100 116.200 86.200 ;
        RECT 118.200 86.100 118.600 86.200 ;
        RECT 115.800 85.800 118.600 86.100 ;
        RECT 120.600 86.100 120.900 86.800 ;
        RECT 123.800 86.100 124.200 86.200 ;
        RECT 120.600 85.800 124.200 86.100 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 128.600 86.100 129.000 86.200 ;
        RECT 125.400 85.800 129.000 86.100 ;
        RECT 131.800 86.100 132.200 86.200 ;
        RECT 134.200 86.100 134.500 86.800 ;
        RECT 144.600 86.100 145.000 86.200 ;
        RECT 131.800 85.800 145.000 86.100 ;
        RECT 146.200 86.100 146.600 86.300 ;
        RECT 153.400 86.100 153.800 86.200 ;
        RECT 146.200 85.800 153.800 86.100 ;
        RECT 158.200 86.100 158.600 86.200 ;
        RECT 170.200 86.100 170.600 86.200 ;
        RECT 158.200 85.800 170.600 86.100 ;
        RECT 171.000 86.100 171.400 86.200 ;
        RECT 175.800 86.100 176.200 86.200 ;
        RECT 188.600 86.100 189.000 86.200 ;
        RECT 189.400 86.100 189.800 86.200 ;
        RECT 197.400 86.100 197.800 86.200 ;
        RECT 204.600 86.100 205.000 86.200 ;
        RECT 171.000 85.800 176.200 86.100 ;
        RECT 182.200 85.800 186.500 86.100 ;
        RECT 188.600 85.800 189.800 86.100 ;
        RECT 191.000 85.800 205.000 86.100 ;
        RECT 219.000 86.100 219.400 86.200 ;
        RECT 221.400 86.100 221.800 86.200 ;
        RECT 219.000 85.800 221.800 86.100 ;
        RECT 227.800 86.100 228.200 86.200 ;
        RECT 230.200 86.100 230.600 86.200 ;
        RECT 227.800 85.800 230.600 86.100 ;
        RECT 231.000 86.100 231.400 86.200 ;
        RECT 243.000 86.100 243.400 86.200 ;
        RECT 231.000 85.800 243.400 86.100 ;
        RECT 33.400 85.200 33.700 85.800 ;
        RECT 34.200 85.200 34.500 85.800 ;
        RECT 125.400 85.200 125.700 85.800 ;
        RECT 182.200 85.200 182.500 85.800 ;
        RECT 186.200 85.200 186.500 85.800 ;
        RECT 191.000 85.200 191.300 85.800 ;
        RECT 2.200 85.100 2.600 85.200 ;
        RECT 8.600 85.100 9.000 85.200 ;
        RECT 2.200 84.800 9.000 85.100 ;
        RECT 33.400 84.800 33.800 85.200 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 57.400 85.100 57.800 85.200 ;
        RECT 70.200 85.100 70.600 85.200 ;
        RECT 57.400 84.800 70.600 85.100 ;
        RECT 85.400 85.100 85.800 85.200 ;
        RECT 89.400 85.100 89.800 85.200 ;
        RECT 85.400 84.800 89.800 85.100 ;
        RECT 91.800 85.100 92.200 85.200 ;
        RECT 101.400 85.100 101.800 85.200 ;
        RECT 91.800 84.800 101.800 85.100 ;
        RECT 104.600 85.100 105.000 85.200 ;
        RECT 107.800 85.100 108.200 85.200 ;
        RECT 104.600 84.800 108.200 85.100 ;
        RECT 110.200 85.100 110.600 85.200 ;
        RECT 116.600 85.100 117.000 85.200 ;
        RECT 110.200 84.800 117.000 85.100 ;
        RECT 119.800 85.100 120.200 85.200 ;
        RECT 121.400 85.100 121.800 85.200 ;
        RECT 119.800 84.800 121.800 85.100 ;
        RECT 125.400 84.800 125.800 85.200 ;
        RECT 127.000 85.100 127.400 85.200 ;
        RECT 135.000 85.100 135.400 85.200 ;
        RECT 127.000 84.800 135.400 85.100 ;
        RECT 150.200 85.100 150.600 85.200 ;
        RECT 152.600 85.100 153.000 85.200 ;
        RECT 155.800 85.100 156.200 85.200 ;
        RECT 156.600 85.100 157.000 85.200 ;
        RECT 150.200 84.800 157.000 85.100 ;
        RECT 161.400 85.100 161.800 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 161.400 84.800 162.600 85.100 ;
        RECT 167.000 85.100 167.400 85.200 ;
        RECT 169.400 85.100 169.800 85.200 ;
        RECT 167.000 84.800 169.800 85.100 ;
        RECT 182.200 84.800 182.600 85.200 ;
        RECT 186.200 84.800 186.600 85.200 ;
        RECT 191.000 84.800 191.400 85.200 ;
        RECT 192.600 84.800 193.000 85.200 ;
        RECT 202.200 85.100 202.600 85.200 ;
        RECT 210.200 85.100 210.600 85.200 ;
        RECT 201.400 84.800 210.600 85.100 ;
        RECT 219.800 85.100 220.200 85.200 ;
        RECT 228.600 85.100 229.000 85.200 ;
        RECT 234.200 85.100 234.600 85.200 ;
        RECT 219.800 84.800 229.000 85.100 ;
        RECT 230.200 84.800 234.600 85.100 ;
        RECT 192.600 84.200 192.900 84.800 ;
        RECT 230.200 84.200 230.500 84.800 ;
        RECT 19.800 84.100 20.200 84.200 ;
        RECT 23.000 84.100 23.400 84.200 ;
        RECT 32.600 84.100 33.000 84.200 ;
        RECT 19.800 83.800 33.000 84.100 ;
        RECT 44.600 84.100 45.000 84.200 ;
        RECT 69.400 84.100 69.800 84.200 ;
        RECT 44.600 83.800 69.800 84.100 ;
        RECT 70.200 84.100 70.600 84.200 ;
        RECT 86.200 84.100 86.600 84.200 ;
        RECT 70.200 83.800 86.600 84.100 ;
        RECT 96.600 84.100 97.000 84.200 ;
        RECT 104.600 84.100 105.000 84.200 ;
        RECT 117.400 84.100 117.800 84.200 ;
        RECT 96.600 83.800 117.800 84.100 ;
        RECT 139.800 84.100 140.200 84.200 ;
        RECT 140.600 84.100 141.000 84.200 ;
        RECT 139.800 83.800 141.000 84.100 ;
        RECT 178.200 84.100 178.600 84.200 ;
        RECT 189.400 84.100 189.800 84.200 ;
        RECT 178.200 83.800 189.800 84.100 ;
        RECT 192.600 83.800 193.000 84.200 ;
        RECT 208.600 84.100 209.000 84.200 ;
        RECT 209.400 84.100 209.800 84.200 ;
        RECT 208.600 83.800 209.800 84.100 ;
        RECT 210.200 84.100 210.600 84.200 ;
        RECT 220.600 84.100 221.000 84.200 ;
        RECT 210.200 83.800 221.000 84.100 ;
        RECT 230.200 83.800 230.600 84.200 ;
        RECT 17.400 83.100 17.800 83.200 ;
        RECT 38.200 83.100 38.600 83.200 ;
        RECT 70.200 83.100 70.600 83.200 ;
        RECT 17.400 82.800 70.600 83.100 ;
        RECT 71.800 83.100 72.200 83.200 ;
        RECT 79.000 83.100 79.400 83.200 ;
        RECT 82.200 83.100 82.600 83.200 ;
        RECT 96.600 83.100 96.900 83.800 ;
        RECT 71.800 82.800 96.900 83.100 ;
        RECT 120.600 83.100 121.000 83.200 ;
        RECT 163.800 83.100 164.200 83.200 ;
        RECT 207.800 83.100 208.200 83.200 ;
        RECT 224.600 83.100 225.000 83.200 ;
        RECT 120.600 82.800 225.000 83.100 ;
        RECT 27.800 82.100 28.200 82.200 ;
        RECT 88.600 82.100 89.000 82.200 ;
        RECT 27.800 81.800 89.000 82.100 ;
        RECT 91.000 82.100 91.400 82.200 ;
        RECT 95.000 82.100 95.400 82.200 ;
        RECT 91.000 81.800 95.400 82.100 ;
        RECT 159.800 82.100 160.200 82.200 ;
        RECT 219.800 82.100 220.200 82.200 ;
        RECT 159.800 81.800 220.200 82.100 ;
        RECT 51.000 81.100 51.400 81.200 ;
        RECT 59.800 81.100 60.200 81.200 ;
        RECT 92.600 81.100 93.000 81.200 ;
        RECT 51.000 80.800 93.000 81.100 ;
        RECT 118.200 81.100 118.600 81.200 ;
        RECT 133.400 81.100 133.800 81.200 ;
        RECT 118.200 80.800 133.800 81.100 ;
        RECT 163.000 81.100 163.400 81.200 ;
        RECT 175.000 81.100 175.400 81.200 ;
        RECT 163.000 80.800 175.400 81.100 ;
        RECT 175.800 81.100 176.200 81.200 ;
        RECT 194.200 81.100 194.600 81.200 ;
        RECT 197.400 81.100 197.800 81.200 ;
        RECT 175.800 80.800 197.800 81.100 ;
        RECT 199.000 81.100 199.400 81.200 ;
        RECT 203.000 81.100 203.400 81.200 ;
        RECT 211.000 81.100 211.400 81.200 ;
        RECT 214.200 81.100 214.600 81.200 ;
        RECT 199.000 80.800 214.600 81.100 ;
        RECT 53.400 80.100 53.800 80.200 ;
        RECT 58.200 80.100 58.600 80.200 ;
        RECT 53.400 79.800 58.600 80.100 ;
        RECT 72.600 80.100 73.000 80.200 ;
        RECT 79.800 80.100 80.200 80.200 ;
        RECT 95.000 80.100 95.400 80.200 ;
        RECT 72.600 79.800 95.400 80.100 ;
        RECT 113.400 80.100 113.800 80.200 ;
        RECT 142.200 80.100 142.600 80.200 ;
        RECT 113.400 79.800 142.600 80.100 ;
        RECT 156.600 80.100 157.000 80.200 ;
        RECT 212.600 80.100 213.000 80.200 ;
        RECT 156.600 79.800 213.000 80.100 ;
        RECT 36.600 79.100 37.000 79.200 ;
        RECT 52.600 79.100 53.000 79.200 ;
        RECT 36.600 78.800 53.000 79.100 ;
        RECT 102.200 79.100 102.600 79.200 ;
        RECT 131.800 79.100 132.200 79.200 ;
        RECT 137.400 79.100 137.800 79.200 ;
        RECT 102.200 78.800 137.800 79.100 ;
        RECT 183.000 79.100 183.400 79.200 ;
        RECT 201.400 79.100 201.800 79.200 ;
        RECT 183.000 78.800 201.800 79.100 ;
        RECT 63.000 78.100 63.400 78.200 ;
        RECT 87.800 78.100 88.200 78.200 ;
        RECT 63.000 77.800 88.200 78.100 ;
        RECT 88.600 78.100 89.000 78.200 ;
        RECT 91.000 78.100 91.400 78.200 ;
        RECT 88.600 77.800 91.400 78.100 ;
        RECT 98.200 78.100 98.600 78.200 ;
        RECT 102.200 78.100 102.600 78.200 ;
        RECT 116.600 78.100 117.000 78.200 ;
        RECT 98.200 77.800 117.000 78.100 ;
        RECT 119.800 78.100 120.200 78.200 ;
        RECT 136.600 78.100 137.000 78.200 ;
        RECT 119.800 77.800 137.000 78.100 ;
        RECT 143.800 78.100 144.200 78.200 ;
        RECT 167.000 78.100 167.400 78.200 ;
        RECT 167.800 78.100 168.200 78.200 ;
        RECT 143.800 77.800 168.200 78.100 ;
        RECT 170.200 78.100 170.600 78.200 ;
        RECT 193.400 78.100 193.800 78.200 ;
        RECT 211.000 78.100 211.400 78.200 ;
        RECT 170.200 77.800 211.400 78.100 ;
        RECT 215.000 78.100 215.400 78.200 ;
        RECT 230.200 78.100 230.600 78.200 ;
        RECT 215.000 77.800 230.600 78.100 ;
        RECT 14.200 77.100 14.600 77.200 ;
        RECT 19.800 77.100 20.200 77.200 ;
        RECT 14.200 76.800 20.200 77.100 ;
        RECT 34.200 77.100 34.600 77.200 ;
        RECT 43.000 77.100 43.400 77.200 ;
        RECT 45.400 77.100 45.800 77.200 ;
        RECT 34.200 76.800 45.800 77.100 ;
        RECT 49.400 77.100 49.800 77.200 ;
        RECT 55.800 77.100 56.200 77.200 ;
        RECT 49.400 76.800 56.200 77.100 ;
        RECT 74.200 77.100 74.600 77.200 ;
        RECT 81.400 77.100 81.800 77.200 ;
        RECT 74.200 76.800 81.800 77.100 ;
        RECT 91.000 77.100 91.400 77.200 ;
        RECT 94.200 77.100 94.600 77.200 ;
        RECT 91.000 76.800 94.600 77.100 ;
        RECT 103.800 77.100 104.200 77.200 ;
        RECT 110.200 77.100 110.600 77.200 ;
        RECT 103.800 76.800 110.600 77.100 ;
        RECT 130.200 77.100 130.600 77.200 ;
        RECT 131.000 77.100 131.400 77.200 ;
        RECT 130.200 76.800 131.400 77.100 ;
        RECT 131.800 77.100 132.200 77.200 ;
        RECT 148.600 77.100 149.000 77.200 ;
        RECT 158.200 77.100 158.600 77.200 ;
        RECT 131.800 76.800 158.600 77.100 ;
        RECT 164.600 77.100 165.000 77.200 ;
        RECT 165.400 77.100 165.800 77.200 ;
        RECT 164.600 76.800 165.800 77.100 ;
        RECT 166.200 77.100 166.600 77.200 ;
        RECT 169.400 77.100 169.800 77.200 ;
        RECT 166.200 76.800 169.800 77.100 ;
        RECT 179.000 77.100 179.400 77.200 ;
        RECT 197.400 77.100 197.800 77.200 ;
        RECT 216.600 77.100 217.000 77.200 ;
        RECT 179.000 76.800 195.300 77.100 ;
        RECT 197.400 76.800 217.000 77.100 ;
        RECT 195.000 76.200 195.300 76.800 ;
        RECT 11.800 75.800 12.200 76.200 ;
        RECT 19.000 75.800 19.400 76.200 ;
        RECT 30.200 76.100 30.600 76.200 ;
        RECT 31.000 76.100 31.400 76.200 ;
        RECT 32.600 76.100 33.000 76.200 ;
        RECT 33.400 76.100 33.800 76.200 ;
        RECT 30.200 75.800 33.800 76.100 ;
        RECT 76.600 76.100 77.000 76.200 ;
        RECT 91.800 76.100 92.200 76.200 ;
        RECT 92.600 76.100 93.000 76.200 ;
        RECT 76.600 75.800 93.000 76.100 ;
        RECT 103.000 76.100 103.400 76.200 ;
        RECT 104.600 76.100 105.000 76.200 ;
        RECT 108.600 76.100 109.000 76.200 ;
        RECT 103.000 75.800 109.000 76.100 ;
        RECT 109.400 76.100 109.800 76.200 ;
        RECT 110.200 76.100 110.600 76.200 ;
        RECT 109.400 75.800 110.600 76.100 ;
        RECT 117.400 75.800 117.800 76.200 ;
        RECT 127.800 76.100 128.200 76.200 ;
        RECT 133.400 76.100 133.800 76.200 ;
        RECT 127.800 75.800 133.800 76.100 ;
        RECT 136.600 75.800 137.000 76.200 ;
        RECT 167.800 76.100 168.200 76.200 ;
        RECT 174.200 76.100 174.600 76.200 ;
        RECT 167.800 75.800 174.600 76.100 ;
        RECT 183.800 76.100 184.200 76.200 ;
        RECT 184.600 76.100 185.000 76.200 ;
        RECT 183.800 75.800 185.000 76.100 ;
        RECT 187.800 76.100 188.200 76.200 ;
        RECT 194.200 76.100 194.600 76.200 ;
        RECT 187.800 75.800 194.600 76.100 ;
        RECT 195.000 75.800 195.400 76.200 ;
        RECT 202.200 76.100 202.600 76.200 ;
        RECT 202.200 75.800 204.900 76.100 ;
        RECT 11.800 75.200 12.100 75.800 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 13.400 75.100 13.800 75.200 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 13.400 74.800 17.000 75.100 ;
        RECT 19.000 75.100 19.300 75.800 ;
        RECT 21.400 75.100 21.800 75.200 ;
        RECT 19.000 74.800 21.800 75.100 ;
        RECT 24.600 75.100 25.000 75.200 ;
        RECT 29.400 75.100 29.800 75.200 ;
        RECT 24.600 74.800 29.800 75.100 ;
        RECT 32.600 75.100 33.000 75.200 ;
        RECT 53.400 75.100 53.800 75.200 ;
        RECT 61.400 75.100 61.800 75.200 ;
        RECT 32.600 74.800 37.700 75.100 ;
        RECT 53.400 74.800 61.800 75.100 ;
        RECT 64.600 75.100 65.000 75.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 64.600 74.800 67.400 75.100 ;
        RECT 72.600 75.100 73.000 75.200 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 98.200 75.100 98.600 75.200 ;
        RECT 72.600 74.800 98.600 75.100 ;
        RECT 103.000 75.100 103.400 75.200 ;
        RECT 103.800 75.100 104.200 75.200 ;
        RECT 103.000 74.800 104.200 75.100 ;
        RECT 107.800 74.800 108.200 75.200 ;
        RECT 115.800 75.100 116.200 75.200 ;
        RECT 116.600 75.100 117.000 75.200 ;
        RECT 115.800 74.800 117.000 75.100 ;
        RECT 117.400 75.100 117.700 75.800 ;
        RECT 136.600 75.200 136.900 75.800 ;
        RECT 204.600 75.200 204.900 75.800 ;
        RECT 207.000 75.800 207.400 76.200 ;
        RECT 215.800 76.100 216.200 76.200 ;
        RECT 219.000 76.100 219.400 76.200 ;
        RECT 215.800 75.800 219.400 76.100 ;
        RECT 248.600 76.100 249.000 76.200 ;
        RECT 249.400 76.100 249.800 76.200 ;
        RECT 248.600 75.800 249.800 76.100 ;
        RECT 207.000 75.200 207.300 75.800 ;
        RECT 122.200 75.100 122.600 75.200 ;
        RECT 117.400 74.800 122.600 75.100 ;
        RECT 129.400 75.100 129.800 75.200 ;
        RECT 131.000 75.100 131.400 75.200 ;
        RECT 129.400 74.800 131.400 75.100 ;
        RECT 131.800 75.100 132.200 75.200 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 131.800 74.800 135.300 75.100 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 139.000 75.100 139.400 75.200 ;
        RECT 140.600 75.100 141.000 75.200 ;
        RECT 160.600 75.100 161.000 75.200 ;
        RECT 162.200 75.100 162.600 75.200 ;
        RECT 169.400 75.100 169.800 75.200 ;
        RECT 138.200 74.800 141.000 75.100 ;
        RECT 153.400 74.800 161.700 75.100 ;
        RECT 162.200 74.800 169.800 75.100 ;
        RECT 171.000 74.800 171.400 75.200 ;
        RECT 183.800 75.100 184.200 75.200 ;
        RECT 184.600 75.100 185.000 75.200 ;
        RECT 183.800 74.800 185.000 75.100 ;
        RECT 187.800 75.100 188.200 75.200 ;
        RECT 195.000 75.100 195.400 75.200 ;
        RECT 197.400 75.100 197.800 75.200 ;
        RECT 187.800 74.800 190.500 75.100 ;
        RECT 195.000 74.800 197.800 75.100 ;
        RECT 204.600 74.800 205.000 75.200 ;
        RECT 207.000 74.800 207.400 75.200 ;
        RECT 215.000 75.100 215.400 75.200 ;
        RECT 225.400 75.100 225.800 75.200 ;
        RECT 215.000 74.800 225.800 75.100 ;
        RECT 244.600 75.100 245.000 75.200 ;
        RECT 246.200 75.100 246.600 75.200 ;
        RECT 244.600 74.800 246.600 75.100 ;
        RECT 37.400 74.200 37.700 74.800 ;
        RECT 107.800 74.200 108.100 74.800 ;
        RECT 153.400 74.700 153.800 74.800 ;
        RECT 5.400 74.100 5.800 74.200 ;
        RECT 12.600 74.100 13.000 74.200 ;
        RECT 19.000 74.100 19.400 74.200 ;
        RECT 23.800 74.100 24.200 74.200 ;
        RECT 5.400 73.800 24.200 74.100 ;
        RECT 25.400 74.100 25.800 74.200 ;
        RECT 27.000 74.100 27.400 74.200 ;
        RECT 31.000 74.100 31.400 74.200 ;
        RECT 25.400 73.800 31.400 74.100 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 44.600 73.800 45.000 74.200 ;
        RECT 52.600 74.100 53.000 74.200 ;
        RECT 54.200 74.100 54.600 74.200 ;
        RECT 52.600 73.800 54.600 74.100 ;
        RECT 63.000 74.100 63.400 74.200 ;
        RECT 89.400 74.100 89.800 74.200 ;
        RECT 92.600 74.100 93.000 74.200 ;
        RECT 94.200 74.100 94.600 74.200 ;
        RECT 95.000 74.100 95.400 74.200 ;
        RECT 63.000 73.800 85.700 74.100 ;
        RECT 89.400 73.800 95.400 74.100 ;
        RECT 104.600 74.100 105.000 74.200 ;
        RECT 106.200 74.100 106.600 74.200 ;
        RECT 104.600 73.800 106.600 74.100 ;
        RECT 107.800 74.100 108.200 74.200 ;
        RECT 117.400 74.100 117.800 74.200 ;
        RECT 107.800 73.800 117.800 74.100 ;
        RECT 119.800 74.100 120.200 74.200 ;
        RECT 151.800 74.100 152.200 74.200 ;
        RECT 119.800 73.800 152.200 74.100 ;
        RECT 160.600 74.100 161.000 74.200 ;
        RECT 161.400 74.100 161.800 74.200 ;
        RECT 160.600 73.800 161.800 74.100 ;
        RECT 167.000 74.100 167.400 74.200 ;
        RECT 170.200 74.100 170.600 74.200 ;
        RECT 167.000 73.800 170.600 74.100 ;
        RECT 171.000 74.100 171.300 74.800 ;
        RECT 190.200 74.200 190.500 74.800 ;
        RECT 180.600 74.100 181.000 74.200 ;
        RECT 188.600 74.100 189.000 74.200 ;
        RECT 171.000 73.800 189.000 74.100 ;
        RECT 190.200 73.800 190.600 74.200 ;
        RECT 200.600 74.100 201.000 74.200 ;
        RECT 201.400 74.100 201.800 74.200 ;
        RECT 200.600 73.800 201.800 74.100 ;
        RECT 204.600 74.100 205.000 74.200 ;
        RECT 205.400 74.100 205.800 74.200 ;
        RECT 204.600 73.800 205.800 74.100 ;
        RECT 211.800 74.100 212.200 74.200 ;
        RECT 215.000 74.100 215.300 74.800 ;
        RECT 229.400 74.100 229.800 74.200 ;
        RECT 211.800 73.800 215.300 74.100 ;
        RECT 219.800 73.800 229.800 74.100 ;
        RECT 239.800 74.100 240.200 74.200 ;
        RECT 242.200 74.100 242.600 74.200 ;
        RECT 239.800 73.800 242.600 74.100 ;
        RECT 247.000 74.100 247.400 74.200 ;
        RECT 249.400 74.100 249.800 74.200 ;
        RECT 247.000 73.800 249.800 74.100 ;
        RECT 44.600 73.200 44.900 73.800 ;
        RECT 85.400 73.200 85.700 73.800 ;
        RECT 219.800 73.200 220.100 73.800 ;
        RECT 44.600 72.800 45.000 73.200 ;
        RECT 71.800 73.100 72.200 73.200 ;
        RECT 77.400 73.100 77.800 73.200 ;
        RECT 71.800 72.800 77.800 73.100 ;
        RECT 85.400 73.100 85.800 73.200 ;
        RECT 103.800 73.100 104.200 73.200 ;
        RECT 115.000 73.100 115.400 73.200 ;
        RECT 115.800 73.100 116.200 73.200 ;
        RECT 85.400 72.800 116.200 73.100 ;
        RECT 116.600 73.100 117.000 73.200 ;
        RECT 124.600 73.100 125.000 73.200 ;
        RECT 116.600 72.800 125.000 73.100 ;
        RECT 129.400 73.100 129.800 73.200 ;
        RECT 130.200 73.100 130.600 73.200 ;
        RECT 129.400 72.800 130.600 73.100 ;
        RECT 169.400 73.100 169.800 73.200 ;
        RECT 193.400 73.100 193.800 73.200 ;
        RECT 199.800 73.100 200.200 73.200 ;
        RECT 169.400 72.800 181.700 73.100 ;
        RECT 193.400 72.800 200.200 73.100 ;
        RECT 219.800 72.800 220.200 73.200 ;
        RECT 44.600 72.100 45.000 72.200 ;
        RECT 46.200 72.100 46.600 72.200 ;
        RECT 44.600 71.800 46.600 72.100 ;
        RECT 50.200 72.100 50.600 72.200 ;
        RECT 68.600 72.100 69.000 72.200 ;
        RECT 50.200 71.800 69.000 72.100 ;
        RECT 77.400 72.100 77.700 72.800 ;
        RECT 181.400 72.200 181.700 72.800 ;
        RECT 86.200 72.100 86.600 72.200 ;
        RECT 77.400 71.800 86.600 72.100 ;
        RECT 90.200 72.100 90.600 72.200 ;
        RECT 102.200 72.100 102.600 72.200 ;
        RECT 90.200 71.800 102.600 72.100 ;
        RECT 111.800 72.100 112.200 72.200 ;
        RECT 113.400 72.100 113.800 72.200 ;
        RECT 123.000 72.100 123.400 72.200 ;
        RECT 111.800 71.800 123.400 72.100 ;
        RECT 127.800 72.100 128.200 72.200 ;
        RECT 139.000 72.100 139.400 72.200 ;
        RECT 143.800 72.100 144.200 72.200 ;
        RECT 127.800 71.800 144.200 72.100 ;
        RECT 157.400 72.100 157.800 72.200 ;
        RECT 177.400 72.100 177.800 72.200 ;
        RECT 157.400 71.800 177.800 72.100 ;
        RECT 181.400 71.800 181.800 72.200 ;
        RECT 183.800 72.100 184.200 72.200 ;
        RECT 199.000 72.100 199.400 72.200 ;
        RECT 208.600 72.100 209.000 72.200 ;
        RECT 183.800 71.800 209.000 72.100 ;
        RECT 211.000 72.100 211.400 72.200 ;
        RECT 217.400 72.100 217.800 72.200 ;
        RECT 211.000 71.800 217.800 72.100 ;
        RECT 45.400 71.100 45.800 71.200 ;
        RECT 53.400 71.100 53.800 71.200 ;
        RECT 75.800 71.100 76.200 71.200 ;
        RECT 45.400 70.800 76.200 71.100 ;
        RECT 83.000 71.100 83.400 71.200 ;
        RECT 97.400 71.100 97.800 71.200 ;
        RECT 83.000 70.800 97.800 71.100 ;
        RECT 100.600 71.100 101.000 71.200 ;
        RECT 115.800 71.100 116.200 71.200 ;
        RECT 100.600 70.800 116.200 71.100 ;
        RECT 116.600 71.100 117.000 71.200 ;
        RECT 129.400 71.100 129.800 71.200 ;
        RECT 116.600 70.800 129.800 71.100 ;
        RECT 132.600 71.100 133.000 71.200 ;
        RECT 141.400 71.100 141.800 71.200 ;
        RECT 132.600 70.800 141.800 71.100 ;
        RECT 142.200 71.100 142.600 71.200 ;
        RECT 162.200 71.100 162.600 71.200 ;
        RECT 165.400 71.100 165.800 71.200 ;
        RECT 142.200 70.800 165.800 71.100 ;
        RECT 167.000 71.100 167.400 71.200 ;
        RECT 191.000 71.100 191.400 71.200 ;
        RECT 167.000 70.800 191.400 71.100 ;
        RECT 17.400 70.100 17.800 70.200 ;
        RECT 19.800 70.100 20.200 70.200 ;
        RECT 34.200 70.100 34.600 70.200 ;
        RECT 17.400 69.800 34.600 70.100 ;
        RECT 71.000 70.100 71.400 70.200 ;
        RECT 89.400 70.100 89.800 70.200 ;
        RECT 92.600 70.100 93.000 70.200 ;
        RECT 94.200 70.100 94.600 70.200 ;
        RECT 71.000 69.800 89.800 70.100 ;
        RECT 90.200 69.800 94.600 70.100 ;
        RECT 105.400 70.100 105.800 70.200 ;
        RECT 106.200 70.100 106.600 70.200 ;
        RECT 143.800 70.100 144.200 70.200 ;
        RECT 105.400 69.800 144.200 70.100 ;
        RECT 159.800 70.100 160.200 70.200 ;
        RECT 185.400 70.100 185.800 70.200 ;
        RECT 159.800 69.800 185.800 70.100 ;
        RECT 203.800 70.100 204.200 70.200 ;
        RECT 209.400 70.100 209.800 70.200 ;
        RECT 203.800 69.800 209.800 70.100 ;
        RECT 212.600 70.100 213.000 70.200 ;
        RECT 215.800 70.100 216.200 70.200 ;
        RECT 212.600 69.800 216.200 70.100 ;
        RECT 251.000 69.800 251.400 70.200 ;
        RECT 10.200 69.100 10.600 69.200 ;
        RECT 21.400 69.100 21.800 69.200 ;
        RECT 10.200 68.800 21.800 69.100 ;
        RECT 29.400 69.100 29.800 69.200 ;
        RECT 63.000 69.100 63.400 69.200 ;
        RECT 67.000 69.100 67.400 69.200 ;
        RECT 29.400 68.800 67.400 69.100 ;
        RECT 68.600 69.100 69.000 69.200 ;
        RECT 90.200 69.100 90.500 69.800 ;
        RECT 251.000 69.200 251.300 69.800 ;
        RECT 68.600 68.800 90.500 69.100 ;
        RECT 91.000 69.100 91.400 69.200 ;
        RECT 95.800 69.100 96.200 69.200 ;
        RECT 115.000 69.100 115.400 69.200 ;
        RECT 91.000 68.800 92.900 69.100 ;
        RECT 95.800 68.800 115.400 69.100 ;
        RECT 115.800 69.100 116.200 69.200 ;
        RECT 118.200 69.100 118.600 69.200 ;
        RECT 115.800 68.800 118.600 69.100 ;
        RECT 119.800 69.100 120.200 69.200 ;
        RECT 123.800 69.100 124.200 69.200 ;
        RECT 128.600 69.100 129.000 69.200 ;
        RECT 172.600 69.100 173.000 69.200 ;
        RECT 174.200 69.100 174.600 69.200 ;
        RECT 119.800 68.800 129.000 69.100 ;
        RECT 151.800 68.800 174.600 69.100 ;
        RECT 186.200 69.100 186.600 69.200 ;
        RECT 202.200 69.100 202.600 69.200 ;
        RECT 220.600 69.100 221.000 69.200 ;
        RECT 186.200 68.800 193.700 69.100 ;
        RECT 202.200 68.800 221.000 69.100 ;
        RECT 226.200 69.100 226.600 69.200 ;
        RECT 233.400 69.100 233.800 69.200 ;
        RECT 242.200 69.100 242.600 69.200 ;
        RECT 226.200 68.800 242.600 69.100 ;
        RECT 251.000 68.800 251.400 69.200 ;
        RECT 4.600 68.100 5.000 68.200 ;
        RECT 5.400 68.100 5.800 68.200 ;
        RECT 4.600 67.800 5.800 68.100 ;
        RECT 21.400 67.800 21.800 68.200 ;
        RECT 31.800 68.100 32.200 68.200 ;
        RECT 35.800 68.100 36.200 68.200 ;
        RECT 31.800 67.800 36.200 68.100 ;
        RECT 39.800 68.100 40.200 68.200 ;
        RECT 51.800 68.100 52.200 68.200 ;
        RECT 39.800 67.800 52.200 68.100 ;
        RECT 55.800 68.100 56.200 68.200 ;
        RECT 58.200 68.100 58.600 68.200 ;
        RECT 76.600 68.100 77.000 68.200 ;
        RECT 55.800 67.800 77.000 68.100 ;
        RECT 77.400 68.100 77.800 68.200 ;
        RECT 83.000 68.100 83.400 68.200 ;
        RECT 77.400 67.800 83.400 68.100 ;
        RECT 83.800 68.100 84.200 68.200 ;
        RECT 87.800 68.100 88.200 68.200 ;
        RECT 91.800 68.100 92.200 68.200 ;
        RECT 83.800 67.800 92.200 68.100 ;
        RECT 92.600 68.100 92.900 68.800 ;
        RECT 151.800 68.200 152.100 68.800 ;
        RECT 100.600 68.100 101.000 68.200 ;
        RECT 92.600 67.800 101.000 68.100 ;
        RECT 104.600 67.800 105.000 68.200 ;
        RECT 106.200 68.100 106.600 68.200 ;
        RECT 107.000 68.100 107.400 68.200 ;
        RECT 106.200 67.800 107.400 68.100 ;
        RECT 114.200 68.100 114.600 68.200 ;
        RECT 116.600 68.100 117.000 68.200 ;
        RECT 114.200 67.800 117.000 68.100 ;
        RECT 127.800 68.100 128.200 68.200 ;
        RECT 133.400 68.100 133.800 68.200 ;
        RECT 127.800 67.800 133.800 68.100 ;
        RECT 151.800 67.800 152.200 68.200 ;
        RECT 167.800 68.100 168.200 68.200 ;
        RECT 168.600 68.100 169.000 68.200 ;
        RECT 167.800 67.800 169.000 68.100 ;
        RECT 169.400 68.100 169.800 68.200 ;
        RECT 172.600 68.100 173.000 68.200 ;
        RECT 169.400 67.800 173.000 68.100 ;
        RECT 188.600 68.100 189.000 68.200 ;
        RECT 192.600 68.100 193.000 68.200 ;
        RECT 188.600 67.800 193.000 68.100 ;
        RECT 193.400 68.100 193.700 68.800 ;
        RECT 203.800 68.100 204.200 68.200 ;
        RECT 193.400 67.800 204.200 68.100 ;
        RECT 209.400 68.100 209.800 68.200 ;
        RECT 216.600 68.100 217.000 68.200 ;
        RECT 209.400 67.800 217.000 68.100 ;
        RECT 223.800 67.800 224.200 68.200 ;
        RECT 224.600 68.100 225.000 68.200 ;
        RECT 225.400 68.100 225.800 68.200 ;
        RECT 224.600 67.800 225.800 68.100 ;
        RECT 228.600 68.100 229.000 68.200 ;
        RECT 229.400 68.100 229.800 68.200 ;
        RECT 228.600 67.800 229.800 68.100 ;
        RECT 231.000 68.100 231.400 68.200 ;
        RECT 231.800 68.100 232.200 68.200 ;
        RECT 231.000 67.800 232.200 68.100 ;
        RECT 239.000 68.100 239.400 68.200 ;
        RECT 245.400 68.100 245.800 68.200 ;
        RECT 239.000 67.800 245.800 68.100 ;
        RECT 1.400 67.100 1.800 67.200 ;
        RECT 6.200 67.100 6.600 67.200 ;
        RECT 9.400 67.100 9.800 67.200 ;
        RECT 1.400 66.800 9.800 67.100 ;
        RECT 15.000 67.100 15.400 67.200 ;
        RECT 21.400 67.100 21.700 67.800 ;
        RECT 15.000 66.800 21.700 67.100 ;
        RECT 29.400 66.800 29.800 67.200 ;
        RECT 32.600 67.100 33.000 67.200 ;
        RECT 33.400 67.100 33.800 67.200 ;
        RECT 32.600 66.800 33.800 67.100 ;
        RECT 35.000 66.800 35.400 67.200 ;
        RECT 41.400 67.100 41.800 67.200 ;
        RECT 45.400 67.100 45.800 67.200 ;
        RECT 41.400 66.800 45.800 67.100 ;
        RECT 46.200 67.100 46.600 67.200 ;
        RECT 48.600 67.100 49.000 67.200 ;
        RECT 46.200 66.800 49.000 67.100 ;
        RECT 51.000 67.100 51.400 67.200 ;
        RECT 53.400 67.100 53.800 67.200 ;
        RECT 51.000 66.800 53.800 67.100 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 58.200 66.800 58.600 67.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 65.400 67.100 65.800 67.200 ;
        RECT 64.600 66.800 65.800 67.100 ;
        RECT 67.800 67.100 68.200 67.200 ;
        RECT 70.200 67.100 70.600 67.200 ;
        RECT 67.800 66.800 70.600 67.100 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 75.800 67.100 76.200 67.200 ;
        RECT 90.200 67.100 90.600 67.200 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 75.800 66.800 94.600 67.100 ;
        RECT 104.600 67.100 104.900 67.800 ;
        RECT 122.200 67.100 122.600 67.200 ;
        RECT 104.600 66.800 122.600 67.100 ;
        RECT 125.400 67.100 125.800 67.200 ;
        RECT 130.200 67.100 130.600 67.200 ;
        RECT 125.400 66.800 130.600 67.100 ;
        RECT 135.800 67.100 136.200 67.200 ;
        RECT 137.400 67.100 137.800 67.200 ;
        RECT 135.800 66.800 137.800 67.100 ;
        RECT 144.600 67.100 145.000 67.200 ;
        RECT 151.800 67.100 152.100 67.800 ;
        RECT 144.600 66.800 152.100 67.100 ;
        RECT 155.800 67.100 156.200 67.200 ;
        RECT 162.200 67.100 162.600 67.200 ;
        RECT 155.800 66.800 162.600 67.100 ;
        RECT 170.200 66.800 170.600 67.200 ;
        RECT 173.400 66.800 173.800 67.200 ;
        RECT 192.600 67.100 193.000 67.200 ;
        RECT 193.400 67.100 193.800 67.200 ;
        RECT 192.600 66.800 193.800 67.100 ;
        RECT 199.000 66.800 199.400 67.200 ;
        RECT 203.000 67.100 203.400 67.200 ;
        RECT 211.800 67.100 212.200 67.200 ;
        RECT 212.600 67.100 213.000 67.200 ;
        RECT 203.000 66.800 213.000 67.100 ;
        RECT 213.400 67.100 213.800 67.200 ;
        RECT 214.200 67.100 214.600 67.200 ;
        RECT 213.400 66.800 214.600 67.100 ;
        RECT 215.000 67.100 215.400 67.200 ;
        RECT 220.600 67.100 221.000 67.200 ;
        RECT 215.000 66.800 221.000 67.100 ;
        RECT 223.800 67.100 224.100 67.800 ;
        RECT 235.800 67.100 236.200 67.200 ;
        RECT 223.800 66.800 236.200 67.100 ;
        RECT 245.400 66.800 245.800 67.200 ;
        RECT 29.400 66.200 29.700 66.800 ;
        RECT 35.000 66.200 35.300 66.800 ;
        RECT 2.200 66.100 2.600 66.200 ;
        RECT 4.600 66.100 5.000 66.200 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 27.800 66.100 28.200 66.200 ;
        RECT 2.200 65.800 5.800 66.100 ;
        RECT 7.800 65.800 28.200 66.100 ;
        RECT 29.400 65.800 29.800 66.200 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 37.400 65.800 38.600 66.100 ;
        RECT 39.800 66.100 40.200 66.200 ;
        RECT 40.600 66.100 41.000 66.200 ;
        RECT 45.400 66.100 45.800 66.200 ;
        RECT 39.800 65.800 41.000 66.100 ;
        RECT 41.400 65.800 45.800 66.100 ;
        RECT 47.000 66.100 47.400 66.200 ;
        RECT 55.000 66.100 55.300 66.800 ;
        RECT 47.000 65.800 55.300 66.100 ;
        RECT 58.200 66.200 58.500 66.800 ;
        RECT 75.000 66.200 75.300 66.800 ;
        RECT 170.200 66.200 170.500 66.800 ;
        RECT 173.400 66.200 173.700 66.800 ;
        RECT 199.000 66.200 199.300 66.800 ;
        RECT 245.400 66.200 245.700 66.800 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 68.600 66.100 69.000 66.200 ;
        RECT 63.000 65.800 69.000 66.100 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 73.400 65.800 74.600 66.100 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 75.800 65.800 77.000 66.100 ;
        RECT 79.000 66.100 79.400 66.200 ;
        RECT 79.800 66.100 80.200 66.200 ;
        RECT 79.000 65.800 80.200 66.100 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 82.200 66.100 82.600 66.200 ;
        RECT 81.400 65.800 82.600 66.100 ;
        RECT 84.600 66.100 85.000 66.200 ;
        RECT 91.000 66.100 91.400 66.200 ;
        RECT 109.400 66.100 109.800 66.200 ;
        RECT 111.800 66.100 112.200 66.200 ;
        RECT 84.600 65.800 91.400 66.100 ;
        RECT 107.000 65.800 109.800 66.100 ;
        RECT 110.200 65.800 112.200 66.100 ;
        RECT 114.200 66.100 114.600 66.200 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 132.600 66.100 133.000 66.200 ;
        RECT 114.200 65.800 133.000 66.100 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 143.000 66.100 143.400 66.200 ;
        RECT 135.800 65.800 143.400 66.100 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 175.000 66.100 175.400 66.200 ;
        RECT 187.000 66.100 187.400 66.200 ;
        RECT 175.000 65.800 187.400 66.100 ;
        RECT 191.000 65.800 191.400 66.200 ;
        RECT 194.200 66.100 194.600 66.200 ;
        RECT 195.000 66.100 195.400 66.200 ;
        RECT 194.200 65.800 195.400 66.100 ;
        RECT 199.000 65.800 199.400 66.200 ;
        RECT 205.400 66.100 205.800 66.200 ;
        RECT 206.200 66.100 206.600 66.200 ;
        RECT 205.400 65.800 229.700 66.100 ;
        RECT 245.400 65.800 245.800 66.200 ;
        RECT 7.800 65.200 8.100 65.800 ;
        RECT 41.400 65.200 41.700 65.800 ;
        RECT 107.000 65.200 107.300 65.800 ;
        RECT 110.200 65.200 110.500 65.800 ;
        RECT 191.000 65.200 191.300 65.800 ;
        RECT 229.400 65.200 229.700 65.800 ;
        RECT 7.800 64.800 8.200 65.200 ;
        RECT 29.400 65.100 29.800 65.200 ;
        RECT 31.000 65.100 31.400 65.200 ;
        RECT 29.400 64.800 31.400 65.100 ;
        RECT 41.400 64.800 41.800 65.200 ;
        RECT 51.800 64.800 52.200 65.200 ;
        RECT 57.400 64.800 57.800 65.200 ;
        RECT 58.200 65.100 58.600 65.200 ;
        RECT 79.000 65.100 79.400 65.200 ;
        RECT 58.200 64.800 79.400 65.100 ;
        RECT 86.200 65.100 86.600 65.200 ;
        RECT 93.400 65.100 93.800 65.200 ;
        RECT 86.200 64.800 93.800 65.100 ;
        RECT 107.000 64.800 107.400 65.200 ;
        RECT 107.800 64.800 108.200 65.200 ;
        RECT 110.200 64.800 110.600 65.200 ;
        RECT 113.400 65.100 113.800 65.200 ;
        RECT 116.600 65.100 117.000 65.200 ;
        RECT 113.400 64.800 117.000 65.100 ;
        RECT 118.200 65.100 118.600 65.200 ;
        RECT 120.600 65.100 121.000 65.200 ;
        RECT 118.200 64.800 121.000 65.100 ;
        RECT 141.400 65.100 141.800 65.200 ;
        RECT 153.400 65.100 153.800 65.200 ;
        RECT 141.400 64.800 153.800 65.100 ;
        RECT 161.400 65.100 161.800 65.200 ;
        RECT 163.000 65.100 163.400 65.200 ;
        RECT 164.600 65.100 165.000 65.200 ;
        RECT 161.400 64.800 165.000 65.100 ;
        RECT 167.800 65.100 168.200 65.200 ;
        RECT 183.800 65.100 184.200 65.200 ;
        RECT 167.800 64.800 184.200 65.100 ;
        RECT 191.000 65.100 191.400 65.200 ;
        RECT 199.800 65.100 200.200 65.200 ;
        RECT 191.000 64.800 200.200 65.100 ;
        RECT 214.200 65.100 214.600 65.200 ;
        RECT 214.200 64.800 215.300 65.100 ;
        RECT 229.400 64.800 229.800 65.200 ;
        RECT 51.800 64.100 52.100 64.800 ;
        RECT 55.800 64.100 56.200 64.200 ;
        RECT 51.800 63.800 56.200 64.100 ;
        RECT 57.400 64.100 57.700 64.800 ;
        RECT 107.800 64.200 108.100 64.800 ;
        RECT 215.000 64.200 215.300 64.800 ;
        RECT 59.000 64.100 59.400 64.200 ;
        RECT 57.400 63.800 59.400 64.100 ;
        RECT 59.800 64.100 60.200 64.200 ;
        RECT 60.600 64.100 61.000 64.200 ;
        RECT 59.800 63.800 61.000 64.100 ;
        RECT 63.800 64.100 64.200 64.200 ;
        RECT 79.000 64.100 79.400 64.200 ;
        RECT 101.400 64.100 101.800 64.200 ;
        RECT 63.800 63.800 79.400 64.100 ;
        RECT 79.800 63.800 101.800 64.100 ;
        RECT 107.800 63.800 108.200 64.200 ;
        RECT 115.800 64.100 116.200 64.200 ;
        RECT 123.000 64.100 123.400 64.200 ;
        RECT 115.800 63.800 123.400 64.100 ;
        RECT 127.000 64.100 127.400 64.200 ;
        RECT 139.800 64.100 140.200 64.200 ;
        RECT 127.000 63.800 140.200 64.100 ;
        RECT 143.000 64.100 143.400 64.200 ;
        RECT 161.400 64.100 161.800 64.200 ;
        RECT 143.000 63.800 161.800 64.100 ;
        RECT 215.000 63.800 215.400 64.200 ;
        RECT 34.200 63.100 34.600 63.200 ;
        RECT 79.800 63.100 80.100 63.800 ;
        RECT 34.200 62.800 80.100 63.100 ;
        RECT 87.800 62.800 88.200 63.200 ;
        RECT 129.400 63.100 129.800 63.200 ;
        RECT 213.400 63.100 213.800 63.200 ;
        RECT 129.400 62.800 213.800 63.100 ;
        RECT 52.600 62.100 53.000 62.200 ;
        RECT 87.800 62.100 88.100 62.800 ;
        RECT 88.600 62.100 89.000 62.200 ;
        RECT 226.200 62.100 226.600 62.200 ;
        RECT 246.200 62.100 246.600 62.200 ;
        RECT 52.600 61.800 246.600 62.100 ;
        RECT 50.200 61.100 50.600 61.200 ;
        RECT 59.000 61.100 59.400 61.200 ;
        RECT 50.200 60.800 59.400 61.100 ;
        RECT 63.800 61.100 64.200 61.200 ;
        RECT 66.200 61.100 66.600 61.200 ;
        RECT 91.000 61.100 91.400 61.200 ;
        RECT 63.800 60.800 91.400 61.100 ;
        RECT 91.800 61.100 92.200 61.200 ;
        RECT 120.600 61.100 121.000 61.200 ;
        RECT 91.800 60.800 121.000 61.100 ;
        RECT 139.000 61.100 139.400 61.200 ;
        RECT 146.200 61.100 146.600 61.200 ;
        RECT 148.600 61.100 149.000 61.200 ;
        RECT 139.000 60.800 149.000 61.100 ;
        RECT 153.400 61.100 153.800 61.200 ;
        RECT 231.800 61.100 232.200 61.200 ;
        RECT 238.200 61.100 238.600 61.200 ;
        RECT 239.000 61.100 239.400 61.200 ;
        RECT 153.400 60.800 239.400 61.100 ;
        RECT 51.800 60.100 52.200 60.200 ;
        RECT 87.800 60.100 88.200 60.200 ;
        RECT 51.800 59.800 88.200 60.100 ;
        RECT 101.400 60.100 101.800 60.200 ;
        RECT 125.400 60.100 125.800 60.200 ;
        RECT 129.400 60.100 129.800 60.200 ;
        RECT 101.400 59.800 129.800 60.100 ;
        RECT 161.400 60.100 161.800 60.200 ;
        RECT 221.400 60.100 221.800 60.200 ;
        RECT 161.400 59.800 221.800 60.100 ;
        RECT 227.800 60.100 228.200 60.200 ;
        RECT 230.200 60.100 230.600 60.200 ;
        RECT 227.800 59.800 230.600 60.100 ;
        RECT 16.600 59.100 17.000 59.200 ;
        RECT 27.000 59.100 27.400 59.200 ;
        RECT 29.400 59.100 29.800 59.200 ;
        RECT 68.600 59.100 69.000 59.200 ;
        RECT 16.600 58.800 69.000 59.100 ;
        RECT 78.200 59.100 78.600 59.200 ;
        RECT 85.400 59.100 85.800 59.200 ;
        RECT 78.200 58.800 85.800 59.100 ;
        RECT 94.200 59.100 94.600 59.200 ;
        RECT 115.000 59.100 115.400 59.200 ;
        RECT 94.200 58.800 115.400 59.100 ;
        RECT 137.400 59.100 137.800 59.200 ;
        RECT 188.600 59.100 189.000 59.200 ;
        RECT 137.400 58.800 189.000 59.100 ;
        RECT 190.200 59.100 190.600 59.200 ;
        RECT 204.600 59.100 205.000 59.200 ;
        RECT 190.200 58.800 205.000 59.100 ;
        RECT 228.600 59.100 229.000 59.200 ;
        RECT 239.800 59.100 240.200 59.200 ;
        RECT 228.600 58.800 240.200 59.100 ;
        RECT 0.600 58.100 1.000 58.200 ;
        RECT 9.400 58.100 9.800 58.200 ;
        RECT 14.200 58.100 14.600 58.200 ;
        RECT 0.600 57.800 14.600 58.100 ;
        RECT 43.000 58.100 43.400 58.200 ;
        RECT 51.800 58.100 52.200 58.200 ;
        RECT 43.000 57.800 52.200 58.100 ;
        RECT 61.400 58.100 61.800 58.200 ;
        RECT 80.600 58.100 81.000 58.200 ;
        RECT 61.400 57.800 81.000 58.100 ;
        RECT 108.600 58.100 109.000 58.200 ;
        RECT 115.000 58.100 115.400 58.200 ;
        RECT 108.600 57.800 115.400 58.100 ;
        RECT 175.800 58.100 176.200 58.200 ;
        RECT 207.800 58.100 208.200 58.200 ;
        RECT 175.800 57.800 208.200 58.100 ;
        RECT 228.600 58.100 229.000 58.200 ;
        RECT 230.200 58.100 230.600 58.200 ;
        RECT 228.600 57.800 230.600 58.100 ;
        RECT 232.600 57.800 233.000 58.200 ;
        RECT 232.600 57.200 232.900 57.800 ;
        RECT 2.200 56.800 2.600 57.200 ;
        RECT 44.600 56.800 45.000 57.200 ;
        RECT 55.000 57.100 55.400 57.200 ;
        RECT 72.600 57.100 73.000 57.200 ;
        RECT 55.000 56.800 73.000 57.100 ;
        RECT 81.400 57.100 81.800 57.200 ;
        RECT 99.800 57.100 100.200 57.200 ;
        RECT 108.600 57.100 109.000 57.200 ;
        RECT 81.400 56.800 109.000 57.100 ;
        RECT 110.200 57.100 110.600 57.200 ;
        RECT 112.600 57.100 113.000 57.200 ;
        RECT 110.200 56.800 113.000 57.100 ;
        RECT 114.200 57.100 114.600 57.200 ;
        RECT 120.600 57.100 121.000 57.200 ;
        RECT 137.400 57.100 137.800 57.200 ;
        RECT 114.200 56.800 137.800 57.100 ;
        RECT 153.400 57.100 153.800 57.200 ;
        RECT 155.800 57.100 156.200 57.200 ;
        RECT 153.400 56.800 156.200 57.100 ;
        RECT 205.400 57.100 205.800 57.200 ;
        RECT 227.800 57.100 228.200 57.200 ;
        RECT 205.400 56.800 228.200 57.100 ;
        RECT 232.600 56.800 233.000 57.200 ;
        RECT 237.400 56.800 237.800 57.200 ;
        RECT 2.200 56.200 2.500 56.800 ;
        RECT 44.600 56.200 44.900 56.800 ;
        RECT 2.200 56.100 2.600 56.200 ;
        RECT 4.600 56.100 5.000 56.200 ;
        RECT 2.200 55.800 5.000 56.100 ;
        RECT 8.600 55.800 9.000 56.200 ;
        RECT 44.600 55.800 45.000 56.200 ;
        RECT 45.400 56.100 45.800 56.200 ;
        RECT 46.200 56.100 46.600 56.200 ;
        RECT 45.400 55.800 46.600 56.100 ;
        RECT 57.400 56.100 57.800 56.200 ;
        RECT 62.200 56.100 62.600 56.200 ;
        RECT 57.400 55.800 62.600 56.100 ;
        RECT 63.800 56.100 64.200 56.200 ;
        RECT 66.200 56.100 66.600 56.200 ;
        RECT 63.800 55.800 66.600 56.100 ;
        RECT 67.800 56.100 68.200 56.200 ;
        RECT 74.200 56.100 74.600 56.200 ;
        RECT 77.400 56.100 77.800 56.200 ;
        RECT 67.800 55.800 77.800 56.100 ;
        RECT 87.000 56.100 87.400 56.200 ;
        RECT 91.800 56.100 92.200 56.200 ;
        RECT 87.000 55.800 92.200 56.100 ;
        RECT 105.400 55.800 105.800 56.200 ;
        RECT 111.800 56.100 112.200 56.200 ;
        RECT 117.400 56.100 117.800 56.200 ;
        RECT 118.200 56.100 118.600 56.200 ;
        RECT 111.800 55.800 118.600 56.100 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 160.600 55.800 161.000 56.200 ;
        RECT 189.400 56.100 189.800 56.200 ;
        RECT 203.000 56.100 203.400 56.200 ;
        RECT 189.400 55.800 203.400 56.100 ;
        RECT 231.000 56.100 231.400 56.200 ;
        RECT 237.400 56.100 237.700 56.800 ;
        RECT 231.000 55.800 237.700 56.100 ;
        RECT 8.600 55.100 8.900 55.800 ;
        RECT 3.800 54.800 8.900 55.100 ;
        RECT 25.400 55.100 25.800 55.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 25.400 54.800 41.000 55.100 ;
        RECT 46.200 55.100 46.600 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 46.200 54.800 47.400 55.100 ;
        RECT 51.000 55.100 51.400 55.200 ;
        RECT 61.400 55.100 61.800 55.200 ;
        RECT 51.000 54.800 61.800 55.100 ;
        RECT 66.200 55.100 66.600 55.200 ;
        RECT 80.600 55.100 81.000 55.200 ;
        RECT 83.000 55.100 83.400 55.200 ;
        RECT 66.200 54.800 72.200 55.100 ;
        RECT 79.800 54.800 83.400 55.100 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 87.800 55.100 88.200 55.200 ;
        RECT 91.800 55.100 92.200 55.200 ;
        RECT 95.800 55.100 96.200 55.200 ;
        RECT 87.800 54.800 88.900 55.100 ;
        RECT 91.800 54.800 96.200 55.100 ;
        RECT 105.400 55.100 105.700 55.800 ;
        RECT 110.200 55.100 110.600 55.200 ;
        RECT 105.400 54.800 110.600 55.100 ;
        RECT 128.600 55.100 129.000 55.200 ;
        RECT 133.400 55.100 133.700 55.800 ;
        RECT 128.600 54.800 133.700 55.100 ;
        RECT 140.600 55.100 141.000 55.200 ;
        RECT 152.600 55.100 153.000 55.200 ;
        RECT 140.600 54.800 153.000 55.100 ;
        RECT 155.000 55.100 155.400 55.200 ;
        RECT 160.600 55.100 160.900 55.800 ;
        RECT 155.000 54.800 160.900 55.100 ;
        RECT 167.800 55.100 168.200 55.200 ;
        RECT 198.200 55.100 198.600 55.200 ;
        RECT 201.400 55.100 201.800 55.200 ;
        RECT 167.800 54.800 201.800 55.100 ;
        RECT 213.400 55.100 213.800 55.200 ;
        RECT 231.800 55.100 232.200 55.200 ;
        RECT 213.400 54.800 232.200 55.100 ;
        RECT 233.400 55.100 233.800 55.200 ;
        RECT 237.400 55.100 237.800 55.200 ;
        RECT 233.400 54.800 237.800 55.100 ;
        RECT 3.800 54.200 4.100 54.800 ;
        RECT 71.800 54.700 72.200 54.800 ;
        RECT 86.200 54.200 86.500 54.800 ;
        RECT 88.600 54.200 88.900 54.800 ;
        RECT 218.200 54.200 218.500 54.800 ;
        RECT 3.800 53.800 4.200 54.200 ;
        RECT 4.600 54.100 5.000 54.200 ;
        RECT 5.400 54.100 5.800 54.200 ;
        RECT 4.600 53.800 5.800 54.100 ;
        RECT 19.000 54.100 19.400 54.200 ;
        RECT 28.600 54.100 29.000 54.200 ;
        RECT 19.000 53.800 29.000 54.100 ;
        RECT 32.600 54.100 33.000 54.200 ;
        RECT 36.600 54.100 37.000 54.200 ;
        RECT 32.600 53.800 37.000 54.100 ;
        RECT 46.200 54.100 46.600 54.200 ;
        RECT 56.600 54.100 57.000 54.200 ;
        RECT 46.200 53.800 57.000 54.100 ;
        RECT 61.400 54.100 61.800 54.200 ;
        RECT 62.200 54.100 62.600 54.200 ;
        RECT 61.400 53.800 62.600 54.100 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 63.000 53.800 64.200 54.100 ;
        RECT 86.200 53.800 86.600 54.200 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 92.600 54.100 93.000 54.200 ;
        RECT 107.000 54.100 107.400 54.200 ;
        RECT 129.400 54.100 129.800 54.200 ;
        RECT 92.600 53.800 129.800 54.100 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 143.800 54.100 144.200 54.200 ;
        RECT 142.200 53.800 144.200 54.100 ;
        RECT 145.400 54.100 145.800 54.200 ;
        RECT 149.400 54.100 149.800 54.200 ;
        RECT 145.400 53.800 149.800 54.100 ;
        RECT 150.200 54.100 150.600 54.200 ;
        RECT 151.800 54.100 152.200 54.200 ;
        RECT 175.800 54.100 176.200 54.200 ;
        RECT 150.200 53.800 176.200 54.100 ;
        RECT 182.200 54.100 182.600 54.200 ;
        RECT 187.000 54.100 187.400 54.200 ;
        RECT 182.200 53.800 187.400 54.100 ;
        RECT 187.800 54.100 188.200 54.200 ;
        RECT 190.200 54.100 190.600 54.200 ;
        RECT 192.600 54.100 193.000 54.200 ;
        RECT 195.800 54.100 196.200 54.200 ;
        RECT 197.400 54.100 197.800 54.200 ;
        RECT 187.800 53.800 191.300 54.100 ;
        RECT 192.600 53.800 197.800 54.100 ;
        RECT 218.200 53.800 218.600 54.200 ;
        RECT 221.400 54.100 221.800 54.200 ;
        RECT 225.400 54.100 225.800 54.200 ;
        RECT 221.400 53.800 225.800 54.100 ;
        RECT 227.000 54.100 227.400 54.200 ;
        RECT 235.800 54.100 236.200 54.200 ;
        RECT 240.600 54.100 241.000 54.200 ;
        RECT 242.200 54.100 242.600 54.200 ;
        RECT 227.000 53.800 242.600 54.100 ;
        RECT 3.800 53.100 4.200 53.200 ;
        RECT 7.000 53.100 7.400 53.200 ;
        RECT 3.800 52.800 7.400 53.100 ;
        RECT 27.800 53.100 28.200 53.200 ;
        RECT 46.200 53.100 46.600 53.200 ;
        RECT 27.800 52.800 46.600 53.100 ;
        RECT 58.200 52.800 58.600 53.200 ;
        RECT 60.600 53.100 61.000 53.200 ;
        RECT 73.400 53.100 73.800 53.200 ;
        RECT 60.600 52.800 73.800 53.100 ;
        RECT 85.400 53.100 85.800 53.200 ;
        RECT 93.400 53.100 93.800 53.200 ;
        RECT 85.400 52.800 93.800 53.100 ;
        RECT 103.000 53.100 103.400 53.200 ;
        RECT 109.400 53.100 109.800 53.200 ;
        RECT 103.000 52.800 109.800 53.100 ;
        RECT 118.200 53.100 118.600 53.200 ;
        RECT 119.000 53.100 119.400 53.200 ;
        RECT 118.200 52.800 119.400 53.100 ;
        RECT 119.800 53.100 120.200 53.200 ;
        RECT 120.600 53.100 121.000 53.200 ;
        RECT 119.800 52.800 121.000 53.100 ;
        RECT 123.800 53.100 124.200 53.200 ;
        RECT 146.200 53.100 146.600 53.200 ;
        RECT 123.800 52.800 146.600 53.100 ;
        RECT 190.200 53.100 190.600 53.200 ;
        RECT 200.600 53.100 201.000 53.200 ;
        RECT 190.200 52.800 201.000 53.100 ;
        RECT 42.200 52.100 42.600 52.200 ;
        RECT 58.200 52.100 58.500 52.800 ;
        RECT 42.200 51.800 58.500 52.100 ;
        RECT 97.400 52.100 97.800 52.200 ;
        RECT 119.800 52.100 120.200 52.200 ;
        RECT 97.400 51.800 120.200 52.100 ;
        RECT 136.600 52.100 137.000 52.200 ;
        RECT 152.600 52.100 153.000 52.200 ;
        RECT 136.600 51.800 153.000 52.100 ;
        RECT 158.200 52.100 158.600 52.200 ;
        RECT 173.400 52.100 173.800 52.200 ;
        RECT 158.200 51.800 173.800 52.100 ;
        RECT 187.000 52.100 187.400 52.200 ;
        RECT 191.800 52.100 192.200 52.200 ;
        RECT 187.000 51.800 192.200 52.100 ;
        RECT 196.600 52.100 197.000 52.200 ;
        RECT 234.200 52.100 234.600 52.200 ;
        RECT 243.000 52.100 243.400 52.200 ;
        RECT 196.600 51.800 243.400 52.100 ;
        RECT 15.000 51.100 15.400 51.200 ;
        RECT 92.600 51.100 93.000 51.200 ;
        RECT 15.000 50.800 93.000 51.100 ;
        RECT 107.800 51.100 108.200 51.200 ;
        RECT 113.400 51.100 113.800 51.200 ;
        RECT 119.000 51.100 119.400 51.200 ;
        RECT 130.200 51.100 130.600 51.200 ;
        RECT 135.800 51.100 136.200 51.200 ;
        RECT 140.600 51.100 141.000 51.200 ;
        RECT 107.800 50.800 141.000 51.100 ;
        RECT 143.800 51.100 144.200 51.200 ;
        RECT 168.600 51.100 169.000 51.200 ;
        RECT 183.800 51.100 184.200 51.200 ;
        RECT 196.600 51.100 197.000 51.200 ;
        RECT 143.800 50.800 197.000 51.100 ;
        RECT 204.600 51.100 205.000 51.200 ;
        RECT 215.000 51.100 215.400 51.200 ;
        RECT 223.800 51.100 224.200 51.200 ;
        RECT 204.600 50.800 224.200 51.100 ;
        RECT 9.400 50.100 9.800 50.200 ;
        RECT 11.800 50.100 12.200 50.200 ;
        RECT 9.400 49.800 12.200 50.100 ;
        RECT 28.600 50.100 29.000 50.200 ;
        RECT 31.000 50.100 31.400 50.200 ;
        RECT 28.600 49.800 31.400 50.100 ;
        RECT 37.400 50.100 37.800 50.200 ;
        RECT 48.600 50.100 49.000 50.200 ;
        RECT 37.400 49.800 49.000 50.100 ;
        RECT 58.200 50.100 58.600 50.200 ;
        RECT 60.600 50.100 61.000 50.200 ;
        RECT 58.200 49.800 61.000 50.100 ;
        RECT 114.200 50.100 114.600 50.200 ;
        RECT 138.200 50.100 138.600 50.200 ;
        RECT 114.200 49.800 138.600 50.100 ;
        RECT 155.800 50.100 156.200 50.200 ;
        RECT 167.800 50.100 168.200 50.200 ;
        RECT 155.800 49.800 168.200 50.100 ;
        RECT 10.200 49.100 10.600 49.200 ;
        RECT 23.800 49.100 24.200 49.200 ;
        RECT 43.800 49.100 44.200 49.200 ;
        RECT 10.200 48.800 44.200 49.100 ;
        RECT 45.400 49.100 45.800 49.200 ;
        RECT 69.400 49.100 69.800 49.200 ;
        RECT 45.400 48.800 69.800 49.100 ;
        RECT 71.000 49.100 71.400 49.200 ;
        RECT 75.800 49.100 76.200 49.200 ;
        RECT 79.000 49.100 79.400 49.200 ;
        RECT 71.000 48.800 79.400 49.100 ;
        RECT 92.600 49.100 93.000 49.200 ;
        RECT 101.400 49.100 101.800 49.200 ;
        RECT 92.600 48.800 101.800 49.100 ;
        RECT 112.600 48.800 113.000 49.200 ;
        RECT 156.600 49.100 157.000 49.200 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 163.000 49.100 163.400 49.200 ;
        RECT 184.600 49.100 185.000 49.200 ;
        RECT 156.600 48.800 159.400 49.100 ;
        RECT 162.200 48.800 185.000 49.100 ;
        RECT 207.000 49.100 207.400 49.200 ;
        RECT 209.400 49.100 209.800 49.200 ;
        RECT 218.200 49.100 218.600 49.200 ;
        RECT 207.000 48.800 218.600 49.100 ;
        RECT 234.200 49.100 234.600 49.200 ;
        RECT 240.600 49.100 241.000 49.200 ;
        RECT 249.400 49.100 249.800 49.200 ;
        RECT 234.200 48.800 249.800 49.100 ;
        RECT 11.800 48.100 12.200 48.200 ;
        RECT 15.000 48.100 15.400 48.200 ;
        RECT 30.200 48.100 30.600 48.200 ;
        RECT 71.000 48.100 71.400 48.200 ;
        RECT 11.800 47.800 71.400 48.100 ;
        RECT 99.800 47.800 100.200 48.200 ;
        RECT 112.600 48.100 112.900 48.800 ;
        RECT 122.200 48.100 122.600 48.200 ;
        RECT 127.800 48.100 128.200 48.200 ;
        RECT 112.600 47.800 128.200 48.100 ;
        RECT 151.800 48.100 152.200 48.200 ;
        RECT 157.400 48.100 157.800 48.200 ;
        RECT 167.000 48.100 167.400 48.200 ;
        RECT 151.800 47.800 167.400 48.100 ;
        RECT 220.600 48.100 221.000 48.200 ;
        RECT 223.000 48.100 223.400 48.200 ;
        RECT 227.000 48.100 227.400 48.200 ;
        RECT 220.600 47.800 227.400 48.100 ;
        RECT 29.400 47.100 29.800 47.200 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 29.400 46.800 30.600 47.100 ;
        RECT 35.800 47.100 36.200 47.200 ;
        RECT 46.200 47.100 46.600 47.200 ;
        RECT 35.800 46.800 46.600 47.100 ;
        RECT 53.400 47.100 53.800 47.200 ;
        RECT 64.600 47.100 65.000 47.200 ;
        RECT 73.400 47.100 73.800 47.200 ;
        RECT 53.400 46.800 62.500 47.100 ;
        RECT 64.600 46.800 73.800 47.100 ;
        RECT 79.800 47.100 80.200 47.200 ;
        RECT 88.600 47.100 89.000 47.200 ;
        RECT 79.800 46.800 89.000 47.100 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 98.200 46.800 98.600 47.200 ;
        RECT 99.800 47.100 100.100 47.800 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 118.200 47.100 118.600 47.200 ;
        RECT 99.800 46.800 118.600 47.100 ;
        RECT 121.400 47.100 121.800 47.200 ;
        RECT 130.200 47.100 130.600 47.200 ;
        RECT 121.400 46.800 130.600 47.100 ;
        RECT 154.200 46.800 154.600 47.200 ;
        RECT 159.000 47.100 159.400 47.200 ;
        RECT 159.800 47.100 160.200 47.200 ;
        RECT 159.000 46.800 160.200 47.100 ;
        RECT 181.400 47.100 181.800 47.200 ;
        RECT 195.800 47.100 196.200 47.200 ;
        RECT 181.400 46.800 196.200 47.100 ;
        RECT 199.000 46.800 199.400 47.200 ;
        RECT 207.800 47.100 208.200 47.200 ;
        RECT 211.800 47.100 212.200 47.200 ;
        RECT 207.800 46.800 212.200 47.100 ;
        RECT 217.400 47.100 217.800 47.200 ;
        RECT 227.800 47.100 228.200 47.200 ;
        RECT 217.400 46.800 228.200 47.100 ;
        RECT 238.200 47.100 238.600 47.200 ;
        RECT 243.800 47.100 244.200 47.200 ;
        RECT 238.200 46.800 244.200 47.100 ;
        RECT 62.200 46.200 62.500 46.800 ;
        RECT 91.000 46.200 91.300 46.800 ;
        RECT 11.800 46.100 12.200 46.200 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 15.000 46.100 15.400 46.200 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 34.200 46.100 34.600 46.200 ;
        RECT 11.800 45.800 34.600 46.100 ;
        RECT 62.200 45.800 62.600 46.200 ;
        RECT 72.600 46.100 73.000 46.200 ;
        RECT 74.200 46.100 74.600 46.200 ;
        RECT 84.600 46.100 85.000 46.200 ;
        RECT 72.600 45.800 85.000 46.100 ;
        RECT 87.800 46.100 88.200 46.200 ;
        RECT 91.000 46.100 91.400 46.200 ;
        RECT 87.800 45.800 91.400 46.100 ;
        RECT 98.200 46.100 98.500 46.800 ;
        RECT 103.800 46.100 104.200 46.200 ;
        RECT 98.200 45.800 104.200 46.100 ;
        RECT 104.600 46.100 105.000 46.200 ;
        RECT 107.800 46.100 108.200 46.200 ;
        RECT 111.000 46.100 111.400 46.200 ;
        RECT 104.600 45.800 111.400 46.100 ;
        RECT 119.800 46.100 120.200 46.200 ;
        RECT 122.200 46.100 122.600 46.200 ;
        RECT 119.800 45.800 122.600 46.100 ;
        RECT 154.200 46.100 154.500 46.800 ;
        RECT 155.800 46.100 156.200 46.200 ;
        RECT 154.200 45.800 156.200 46.100 ;
        RECT 157.400 46.100 157.800 46.200 ;
        RECT 159.800 46.100 160.200 46.200 ;
        RECT 160.600 46.100 161.000 46.200 ;
        RECT 157.400 45.800 161.000 46.100 ;
        RECT 186.200 46.100 186.600 46.200 ;
        RECT 187.000 46.100 187.400 46.200 ;
        RECT 187.800 46.100 188.200 46.200 ;
        RECT 186.200 45.800 188.200 46.100 ;
        RECT 199.000 46.100 199.300 46.800 ;
        RECT 200.600 46.100 201.000 46.200 ;
        RECT 199.000 45.800 201.000 46.100 ;
        RECT 203.000 46.100 203.400 46.200 ;
        RECT 211.800 46.100 212.100 46.800 ;
        RECT 203.000 45.800 212.100 46.100 ;
        RECT 214.200 46.100 214.600 46.300 ;
        RECT 219.800 46.100 220.200 46.200 ;
        RECT 214.200 45.800 220.200 46.100 ;
        RECT 225.400 46.100 225.800 46.200 ;
        RECT 233.400 46.100 233.800 46.200 ;
        RECT 234.200 46.100 234.600 46.200 ;
        RECT 225.400 45.800 226.500 46.100 ;
        RECT 233.400 45.800 234.600 46.100 ;
        RECT 237.400 46.100 237.800 46.200 ;
        RECT 239.000 46.100 239.400 46.200 ;
        RECT 237.400 45.800 239.400 46.100 ;
        RECT 226.200 45.200 226.500 45.800 ;
        RECT 239.000 45.200 239.300 45.800 ;
        RECT 15.000 45.100 15.400 45.200 ;
        RECT 18.200 45.100 18.600 45.200 ;
        RECT 14.200 44.800 18.600 45.100 ;
        RECT 32.600 45.100 33.000 45.200 ;
        RECT 40.600 45.100 41.000 45.200 ;
        RECT 32.600 44.800 41.000 45.100 ;
        RECT 45.400 44.800 45.800 45.200 ;
        RECT 58.200 44.800 58.600 45.200 ;
        RECT 59.800 45.100 60.200 45.200 ;
        RECT 77.400 45.100 77.800 45.200 ;
        RECT 59.800 44.800 77.800 45.100 ;
        RECT 84.600 45.100 85.000 45.200 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 84.600 44.800 85.800 45.100 ;
        RECT 93.400 45.100 93.800 45.200 ;
        RECT 120.600 45.100 121.000 45.200 ;
        RECT 93.400 44.800 121.000 45.100 ;
        RECT 179.800 45.100 180.200 45.200 ;
        RECT 188.600 45.100 189.000 45.200 ;
        RECT 179.800 44.800 189.000 45.100 ;
        RECT 195.000 45.100 195.400 45.200 ;
        RECT 199.000 45.100 199.400 45.200 ;
        RECT 195.000 44.800 199.400 45.100 ;
        RECT 226.200 44.800 226.600 45.200 ;
        RECT 239.000 44.800 239.400 45.200 ;
        RECT 2.200 44.100 2.600 44.200 ;
        RECT 36.600 44.100 37.000 44.200 ;
        RECT 45.400 44.100 45.700 44.800 ;
        RECT 2.200 43.800 45.700 44.100 ;
        RECT 58.200 44.200 58.500 44.800 ;
        RECT 58.200 43.800 58.600 44.200 ;
        RECT 60.600 44.100 61.000 44.200 ;
        RECT 82.200 44.100 82.600 44.200 ;
        RECT 103.000 44.100 103.400 44.200 ;
        RECT 60.600 43.800 103.400 44.100 ;
        RECT 111.000 44.100 111.400 44.200 ;
        RECT 134.200 44.100 134.600 44.200 ;
        RECT 111.000 43.800 134.600 44.100 ;
        RECT 165.400 44.100 165.800 44.200 ;
        RECT 185.400 44.100 185.800 44.200 ;
        RECT 207.800 44.100 208.200 44.200 ;
        RECT 165.400 43.800 208.200 44.100 ;
        RECT 219.800 44.100 220.200 44.200 ;
        RECT 222.200 44.100 222.600 44.200 ;
        RECT 251.800 44.100 252.200 44.200 ;
        RECT 219.800 43.800 252.200 44.100 ;
        RECT 12.600 43.100 13.000 43.200 ;
        RECT 52.600 43.100 53.000 43.200 ;
        RECT 12.600 42.800 53.000 43.100 ;
        RECT 95.000 43.100 95.400 43.200 ;
        RECT 118.200 43.100 118.600 43.200 ;
        RECT 167.000 43.100 167.400 43.200 ;
        RECT 169.400 43.100 169.800 43.200 ;
        RECT 95.000 42.800 169.800 43.100 ;
        RECT 178.200 43.100 178.600 43.200 ;
        RECT 189.400 43.100 189.800 43.200 ;
        RECT 178.200 42.800 189.800 43.100 ;
        RECT 55.000 42.100 55.400 42.200 ;
        RECT 97.400 42.100 97.800 42.200 ;
        RECT 55.000 41.800 97.800 42.100 ;
        RECT 120.600 42.100 121.000 42.200 ;
        RECT 135.800 42.100 136.200 42.200 ;
        RECT 155.000 42.100 155.400 42.200 ;
        RECT 178.200 42.100 178.500 42.800 ;
        RECT 120.600 41.800 178.500 42.100 ;
        RECT 86.200 41.100 86.600 41.200 ;
        RECT 88.600 41.100 89.000 41.200 ;
        RECT 90.200 41.100 90.600 41.200 ;
        RECT 86.200 40.800 90.600 41.100 ;
        RECT 120.600 41.100 121.000 41.200 ;
        RECT 146.200 41.100 146.600 41.200 ;
        RECT 120.600 40.800 146.600 41.100 ;
        RECT 86.200 40.100 86.600 40.200 ;
        RECT 122.200 40.100 122.600 40.200 ;
        RECT 86.200 39.800 122.600 40.100 ;
        RECT 15.800 39.100 16.200 39.200 ;
        RECT 18.200 39.100 18.600 39.200 ;
        RECT 27.000 39.100 27.400 39.200 ;
        RECT 15.800 38.800 27.400 39.100 ;
        RECT 95.800 39.100 96.200 39.200 ;
        RECT 141.400 39.100 141.800 39.200 ;
        RECT 143.800 39.100 144.200 39.200 ;
        RECT 95.800 38.800 144.200 39.100 ;
        RECT 186.200 39.100 186.600 39.200 ;
        RECT 191.800 39.100 192.200 39.200 ;
        RECT 207.000 39.100 207.400 39.200 ;
        RECT 186.200 38.800 207.400 39.100 ;
        RECT 72.600 38.100 73.000 38.200 ;
        RECT 88.600 38.100 89.000 38.200 ;
        RECT 98.200 38.100 98.600 38.200 ;
        RECT 111.000 38.100 111.400 38.200 ;
        RECT 72.600 37.800 111.400 38.100 ;
        RECT 134.200 38.100 134.600 38.200 ;
        RECT 155.800 38.100 156.200 38.200 ;
        RECT 134.200 37.800 156.200 38.100 ;
        RECT 164.600 38.100 165.000 38.200 ;
        RECT 191.800 38.100 192.200 38.200 ;
        RECT 197.400 38.100 197.800 38.200 ;
        RECT 164.600 37.800 197.800 38.100 ;
        RECT 5.400 37.100 5.800 37.200 ;
        RECT 15.000 37.100 15.400 37.200 ;
        RECT 35.000 37.100 35.400 37.200 ;
        RECT 5.400 36.800 35.400 37.100 ;
        RECT 37.400 37.100 37.800 37.200 ;
        RECT 39.000 37.100 39.400 37.200 ;
        RECT 37.400 36.800 39.400 37.100 ;
        RECT 51.800 37.100 52.200 37.200 ;
        RECT 55.000 37.100 55.400 37.200 ;
        RECT 51.800 36.800 55.400 37.100 ;
        RECT 85.400 37.100 85.800 37.200 ;
        RECT 91.800 37.100 92.200 37.200 ;
        RECT 96.600 37.100 97.000 37.200 ;
        RECT 85.400 36.800 97.000 37.100 ;
        RECT 110.200 37.100 110.600 37.200 ;
        RECT 119.000 37.100 119.400 37.200 ;
        RECT 121.400 37.100 121.800 37.200 ;
        RECT 110.200 36.800 121.800 37.100 ;
        RECT 128.600 37.100 129.000 37.200 ;
        RECT 131.000 37.100 131.400 37.200 ;
        RECT 139.800 37.100 140.200 37.200 ;
        RECT 128.600 36.800 140.200 37.100 ;
        RECT 166.200 36.800 166.600 37.200 ;
        RECT 182.200 37.100 182.600 37.200 ;
        RECT 187.000 37.100 187.400 37.200 ;
        RECT 182.200 36.800 187.400 37.100 ;
        RECT 213.400 36.800 213.800 37.200 ;
        RECT 223.800 36.800 224.200 37.200 ;
        RECT 229.400 37.100 229.800 37.200 ;
        RECT 241.400 37.100 241.800 37.200 ;
        RECT 250.200 37.100 250.600 37.200 ;
        RECT 229.400 36.800 250.600 37.100 ;
        RECT 166.200 36.200 166.500 36.800 ;
        RECT 10.200 36.100 10.600 36.200 ;
        RECT 41.400 36.100 41.800 36.200 ;
        RECT 10.200 35.800 41.800 36.100 ;
        RECT 43.000 36.100 43.400 36.200 ;
        RECT 47.800 36.100 48.200 36.200 ;
        RECT 50.200 36.100 50.600 36.200 ;
        RECT 43.000 35.800 50.600 36.100 ;
        RECT 55.800 36.100 56.200 36.200 ;
        RECT 67.000 36.100 67.400 36.200 ;
        RECT 87.000 36.100 87.400 36.200 ;
        RECT 55.800 35.800 87.400 36.100 ;
        RECT 107.800 36.100 108.200 36.200 ;
        RECT 113.400 36.100 113.800 36.200 ;
        RECT 107.800 35.800 113.800 36.100 ;
        RECT 114.200 36.100 114.600 36.200 ;
        RECT 147.000 36.100 147.400 36.200 ;
        RECT 148.600 36.100 149.000 36.200 ;
        RECT 164.600 36.100 165.000 36.200 ;
        RECT 114.200 35.800 165.000 36.100 ;
        RECT 166.200 35.800 166.600 36.200 ;
        RECT 187.000 36.100 187.400 36.200 ;
        RECT 193.400 36.100 193.800 36.200 ;
        RECT 186.200 35.800 193.800 36.100 ;
        RECT 198.200 36.100 198.600 36.200 ;
        RECT 213.400 36.100 213.700 36.800 ;
        RECT 198.200 35.800 213.700 36.100 ;
        RECT 221.400 36.100 221.800 36.200 ;
        RECT 223.000 36.100 223.400 36.200 ;
        RECT 223.800 36.100 224.100 36.800 ;
        RECT 221.400 35.800 224.100 36.100 ;
        RECT 237.400 36.100 237.800 36.200 ;
        RECT 239.800 36.100 240.200 36.200 ;
        RECT 240.600 36.100 241.000 36.200 ;
        RECT 237.400 35.800 241.000 36.100 ;
        RECT 244.600 35.800 245.000 36.200 ;
        RECT 250.200 36.100 250.600 36.200 ;
        RECT 251.000 36.100 251.400 36.200 ;
        RECT 250.200 35.800 251.400 36.100 ;
        RECT 11.000 35.100 11.400 35.200 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 15.000 35.100 15.400 35.200 ;
        RECT 11.000 34.800 13.000 35.100 ;
        RECT 14.200 34.800 15.400 35.100 ;
        RECT 19.800 35.100 20.200 35.200 ;
        RECT 25.400 35.100 25.800 35.200 ;
        RECT 29.400 35.100 29.800 35.200 ;
        RECT 19.800 34.800 29.800 35.100 ;
        RECT 39.000 35.100 39.400 35.200 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 39.000 34.800 40.200 35.100 ;
        RECT 41.400 35.100 41.800 35.200 ;
        RECT 44.600 35.100 45.000 35.200 ;
        RECT 51.000 35.100 51.400 35.200 ;
        RECT 41.400 34.800 51.400 35.100 ;
        RECT 51.800 35.100 52.200 35.200 ;
        RECT 52.600 35.100 53.000 35.200 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 51.800 34.800 61.000 35.100 ;
        RECT 67.000 35.100 67.400 35.200 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 67.000 34.800 68.200 35.100 ;
        RECT 69.400 35.100 69.800 35.200 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 69.400 34.800 70.600 35.100 ;
        RECT 82.200 35.100 82.600 35.200 ;
        RECT 88.600 35.100 89.000 35.200 ;
        RECT 82.200 34.800 89.000 35.100 ;
        RECT 92.600 35.100 93.000 35.200 ;
        RECT 93.400 35.100 93.800 35.200 ;
        RECT 92.600 34.800 93.800 35.100 ;
        RECT 97.400 35.100 97.800 35.200 ;
        RECT 105.400 35.100 105.800 35.200 ;
        RECT 108.600 35.100 109.000 35.200 ;
        RECT 97.400 34.800 109.000 35.100 ;
        RECT 130.200 35.100 130.600 35.200 ;
        RECT 165.400 35.100 165.800 35.200 ;
        RECT 130.200 34.800 165.800 35.100 ;
        RECT 167.000 35.100 167.400 35.200 ;
        RECT 176.600 35.100 177.000 35.200 ;
        RECT 167.000 34.800 177.000 35.100 ;
        RECT 181.400 35.100 181.800 35.200 ;
        RECT 183.800 35.100 184.200 35.200 ;
        RECT 185.400 35.100 185.800 35.200 ;
        RECT 181.400 34.800 185.800 35.100 ;
        RECT 215.000 35.100 215.400 35.200 ;
        RECT 217.400 35.100 217.800 35.200 ;
        RECT 215.000 34.800 217.800 35.100 ;
        RECT 239.800 35.100 240.200 35.200 ;
        RECT 244.600 35.100 244.900 35.800 ;
        RECT 239.800 34.800 244.900 35.100 ;
        RECT 14.200 34.200 14.500 34.800 ;
        RECT 14.200 33.800 14.600 34.200 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 23.000 34.100 23.400 34.200 ;
        RECT 17.400 33.800 23.400 34.100 ;
        RECT 38.200 34.100 38.600 34.200 ;
        RECT 40.600 34.100 41.000 34.200 ;
        RECT 38.200 33.800 41.000 34.100 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 54.200 34.100 54.600 34.200 ;
        RECT 56.600 34.100 57.000 34.200 ;
        RECT 54.200 33.800 57.000 34.100 ;
        RECT 76.600 34.100 77.000 34.200 ;
        RECT 76.600 33.800 87.300 34.100 ;
        RECT 3.800 33.100 4.200 33.200 ;
        RECT 21.400 33.100 21.800 33.200 ;
        RECT 3.800 32.800 21.800 33.100 ;
        RECT 24.600 33.100 25.000 33.200 ;
        RECT 52.600 33.100 52.900 33.800 ;
        RECT 87.000 33.200 87.300 33.800 ;
        RECT 96.600 33.800 97.000 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 107.800 34.100 108.200 34.200 ;
        RECT 131.800 34.100 132.200 34.200 ;
        RECT 104.600 33.800 132.200 34.100 ;
        RECT 136.600 34.100 137.000 34.200 ;
        RECT 141.400 34.100 141.800 34.200 ;
        RECT 136.600 33.800 141.800 34.100 ;
        RECT 145.400 34.100 145.800 34.200 ;
        RECT 147.000 34.100 147.400 34.200 ;
        RECT 145.400 33.800 147.400 34.100 ;
        RECT 157.400 34.100 157.800 34.200 ;
        RECT 162.200 34.100 162.600 34.200 ;
        RECT 157.400 33.800 162.600 34.100 ;
        RECT 168.600 34.100 169.000 34.200 ;
        RECT 170.200 34.100 170.600 34.200 ;
        RECT 171.800 34.100 172.200 34.200 ;
        RECT 168.600 33.800 172.200 34.100 ;
        RECT 177.400 34.100 177.800 34.200 ;
        RECT 215.800 34.100 216.200 34.200 ;
        RECT 219.800 34.100 220.200 34.200 ;
        RECT 177.400 33.800 220.200 34.100 ;
        RECT 232.600 34.100 233.000 34.200 ;
        RECT 234.200 34.100 234.600 34.200 ;
        RECT 232.600 33.800 234.600 34.100 ;
        RECT 236.600 34.100 237.000 34.200 ;
        RECT 236.600 33.800 243.300 34.100 ;
        RECT 24.600 32.800 52.900 33.100 ;
        RECT 55.000 33.100 55.400 33.200 ;
        RECT 56.600 33.100 57.000 33.200 ;
        RECT 55.000 32.800 57.000 33.100 ;
        RECT 83.000 33.100 83.400 33.200 ;
        RECT 84.600 33.100 85.000 33.200 ;
        RECT 83.000 32.800 85.000 33.100 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 89.400 33.100 89.800 33.200 ;
        RECT 91.800 33.100 92.200 33.200 ;
        RECT 88.600 32.800 92.200 33.100 ;
        RECT 96.600 33.100 96.900 33.800 ;
        RECT 243.000 33.200 243.300 33.800 ;
        RECT 105.400 33.100 105.800 33.200 ;
        RECT 111.800 33.100 112.200 33.200 ;
        RECT 96.600 32.800 112.200 33.100 ;
        RECT 169.400 33.100 169.800 33.200 ;
        RECT 204.600 33.100 205.000 33.200 ;
        RECT 208.600 33.100 209.000 33.200 ;
        RECT 169.400 32.800 209.000 33.100 ;
        RECT 243.000 32.800 243.400 33.200 ;
        RECT 32.600 32.100 33.000 32.200 ;
        RECT 33.400 32.100 33.800 32.200 ;
        RECT 32.600 31.800 33.800 32.100 ;
        RECT 63.800 32.100 64.200 32.200 ;
        RECT 96.600 32.100 97.000 32.200 ;
        RECT 63.800 31.800 97.000 32.100 ;
        RECT 101.400 32.100 101.800 32.200 ;
        RECT 127.800 32.100 128.200 32.200 ;
        RECT 145.400 32.100 145.800 32.200 ;
        RECT 167.000 32.100 167.400 32.200 ;
        RECT 101.400 31.800 128.200 32.100 ;
        RECT 128.600 31.800 167.400 32.100 ;
        RECT 171.000 32.100 171.400 32.200 ;
        RECT 186.200 32.100 186.600 32.200 ;
        RECT 171.000 31.800 186.600 32.100 ;
        RECT 202.200 32.100 202.600 32.200 ;
        RECT 205.400 32.100 205.800 32.200 ;
        RECT 202.200 31.800 205.800 32.100 ;
        RECT 20.600 31.100 21.000 31.200 ;
        RECT 31.000 31.100 31.400 31.200 ;
        RECT 20.600 30.800 31.400 31.100 ;
        RECT 68.600 31.100 69.000 31.200 ;
        RECT 73.400 31.100 73.800 31.200 ;
        RECT 68.600 30.800 73.800 31.100 ;
        RECT 100.600 31.100 101.000 31.200 ;
        RECT 128.600 31.100 128.900 31.800 ;
        RECT 100.600 30.800 128.900 31.100 ;
        RECT 147.800 31.100 148.200 31.200 ;
        RECT 153.400 31.100 153.800 31.200 ;
        RECT 147.800 30.800 153.800 31.100 ;
        RECT 157.400 31.100 157.800 31.200 ;
        RECT 175.800 31.100 176.200 31.200 ;
        RECT 196.600 31.100 197.000 31.200 ;
        RECT 157.400 30.800 197.000 31.100 ;
        RECT 2.200 30.100 2.600 30.200 ;
        RECT 4.600 30.100 5.000 30.200 ;
        RECT 10.200 30.100 10.600 30.200 ;
        RECT 2.200 29.800 10.600 30.100 ;
        RECT 30.200 29.800 30.600 30.200 ;
        RECT 31.000 30.100 31.400 30.200 ;
        RECT 38.200 30.100 38.600 30.200 ;
        RECT 31.000 29.800 38.600 30.100 ;
        RECT 61.400 30.100 61.800 30.200 ;
        RECT 85.400 30.100 85.800 30.200 ;
        RECT 61.400 29.800 85.800 30.100 ;
        RECT 140.600 30.100 141.000 30.200 ;
        RECT 141.400 30.100 141.800 30.200 ;
        RECT 140.600 29.800 141.800 30.100 ;
        RECT 151.800 30.100 152.200 30.200 ;
        RECT 161.400 30.100 161.800 30.200 ;
        RECT 151.800 29.800 161.800 30.100 ;
        RECT 167.000 30.100 167.400 30.200 ;
        RECT 186.200 30.100 186.600 30.200 ;
        RECT 167.000 29.800 186.600 30.100 ;
        RECT 250.200 30.100 250.600 30.200 ;
        RECT 251.800 30.100 252.200 30.200 ;
        RECT 250.200 29.800 252.200 30.100 ;
        RECT 6.200 29.100 6.600 29.200 ;
        RECT 19.800 29.100 20.200 29.200 ;
        RECT 6.200 28.800 20.200 29.100 ;
        RECT 30.200 29.100 30.500 29.800 ;
        RECT 50.200 29.100 50.600 29.200 ;
        RECT 30.200 28.800 50.600 29.100 ;
        RECT 79.800 29.100 80.200 29.200 ;
        RECT 82.200 29.100 82.600 29.200 ;
        RECT 79.800 28.800 82.600 29.100 ;
        RECT 83.800 29.100 84.200 29.200 ;
        RECT 85.400 29.100 85.700 29.800 ;
        RECT 83.800 28.800 85.700 29.100 ;
        RECT 97.400 29.100 97.800 29.200 ;
        RECT 106.200 29.100 106.600 29.200 ;
        RECT 97.400 28.800 106.600 29.100 ;
        RECT 114.200 28.800 114.600 29.200 ;
        RECT 126.200 29.100 126.600 29.200 ;
        RECT 131.800 29.100 132.200 29.200 ;
        RECT 140.600 29.100 141.000 29.200 ;
        RECT 159.000 29.100 159.400 29.200 ;
        RECT 164.600 29.100 165.000 29.200 ;
        RECT 126.200 28.800 141.000 29.100 ;
        RECT 158.200 28.800 165.000 29.100 ;
        RECT 178.200 29.100 178.600 29.200 ;
        RECT 181.400 29.100 181.800 29.200 ;
        RECT 187.800 29.100 188.200 29.200 ;
        RECT 178.200 28.800 188.200 29.100 ;
        RECT 226.200 29.100 226.600 29.200 ;
        RECT 229.400 29.100 229.800 29.200 ;
        RECT 226.200 28.800 229.800 29.100 ;
        RECT 231.000 29.100 231.400 29.200 ;
        RECT 239.000 29.100 239.400 29.200 ;
        RECT 231.000 28.800 239.400 29.100 ;
        RECT 248.600 29.100 249.000 29.200 ;
        RECT 248.600 28.800 252.100 29.100 ;
        RECT 11.000 28.100 11.400 28.200 ;
        RECT 11.800 28.100 12.200 28.200 ;
        RECT 11.000 27.800 12.200 28.100 ;
        RECT 48.600 28.100 49.000 28.200 ;
        RECT 66.200 28.100 66.600 28.200 ;
        RECT 48.600 27.800 66.600 28.100 ;
        RECT 70.200 28.100 70.600 28.200 ;
        RECT 75.800 28.100 76.200 28.200 ;
        RECT 100.600 28.100 101.000 28.200 ;
        RECT 70.200 27.800 101.000 28.100 ;
        RECT 110.200 27.800 110.600 28.200 ;
        RECT 111.000 27.800 111.400 28.200 ;
        RECT 114.200 28.100 114.500 28.800 ;
        RECT 251.800 28.200 252.100 28.800 ;
        RECT 119.800 28.100 120.200 28.200 ;
        RECT 114.200 27.800 120.200 28.100 ;
        RECT 131.800 28.100 132.200 28.200 ;
        RECT 167.000 28.100 167.400 28.200 ;
        RECT 131.800 27.800 167.400 28.100 ;
        RECT 169.400 28.100 169.800 28.200 ;
        RECT 177.400 28.100 177.800 28.200 ;
        RECT 169.400 27.800 177.800 28.100 ;
        RECT 186.200 28.100 186.600 28.200 ;
        RECT 211.800 28.100 212.200 28.200 ;
        RECT 186.200 27.800 212.200 28.100 ;
        RECT 249.400 27.800 249.800 28.200 ;
        RECT 251.800 27.800 252.200 28.200 ;
        RECT 110.200 27.200 110.500 27.800 ;
        RECT 1.400 27.100 1.800 27.200 ;
        RECT 7.800 27.100 8.200 27.200 ;
        RECT 1.400 26.800 8.200 27.100 ;
        RECT 47.000 27.100 47.400 27.200 ;
        RECT 59.000 27.100 59.400 27.200 ;
        RECT 47.000 26.800 59.400 27.100 ;
        RECT 65.400 27.100 65.800 27.200 ;
        RECT 79.000 27.100 79.400 27.200 ;
        RECT 65.400 26.800 79.400 27.100 ;
        RECT 80.600 26.800 81.000 27.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 99.800 26.800 100.200 27.200 ;
        RECT 103.000 27.100 103.400 27.200 ;
        RECT 108.600 27.100 109.000 27.200 ;
        RECT 103.000 26.800 109.000 27.100 ;
        RECT 110.200 26.800 110.600 27.200 ;
        RECT 111.000 27.100 111.300 27.800 ;
        RECT 127.000 27.100 127.400 27.200 ;
        RECT 111.000 26.800 127.400 27.100 ;
        RECT 127.800 27.100 128.200 27.200 ;
        RECT 128.600 27.100 129.000 27.200 ;
        RECT 127.800 26.800 129.000 27.100 ;
        RECT 129.400 27.100 129.800 27.200 ;
        RECT 135.000 27.100 135.400 27.200 ;
        RECT 129.400 26.800 135.400 27.100 ;
        RECT 141.400 27.100 141.800 27.200 ;
        RECT 142.200 27.100 142.600 27.200 ;
        RECT 141.400 26.800 142.600 27.100 ;
        RECT 143.000 27.100 143.400 27.200 ;
        RECT 146.200 27.100 146.600 27.200 ;
        RECT 143.000 26.800 146.600 27.100 ;
        RECT 151.000 27.100 151.400 27.200 ;
        RECT 155.000 27.100 155.400 27.200 ;
        RECT 159.000 27.100 159.400 27.200 ;
        RECT 151.000 26.800 159.400 27.100 ;
        RECT 163.800 27.100 164.200 27.200 ;
        RECT 207.800 27.100 208.200 27.200 ;
        RECT 210.200 27.100 210.600 27.200 ;
        RECT 163.800 26.800 210.600 27.100 ;
        RECT 212.600 27.100 213.000 27.200 ;
        RECT 215.800 27.100 216.200 27.200 ;
        RECT 212.600 26.800 216.200 27.100 ;
        RECT 216.600 26.800 217.000 27.200 ;
        RECT 223.000 27.100 223.400 27.200 ;
        RECT 235.800 27.100 236.200 27.200 ;
        RECT 223.000 26.800 236.200 27.100 ;
        RECT 236.600 27.100 237.000 27.200 ;
        RECT 249.400 27.100 249.700 27.800 ;
        RECT 236.600 26.800 249.700 27.100 ;
        RECT 7.800 26.100 8.200 26.200 ;
        RECT 10.200 26.100 10.600 26.200 ;
        RECT 7.800 25.800 10.600 26.100 ;
        RECT 36.600 26.100 37.000 26.300 ;
        RECT 80.600 26.200 80.900 26.800 ;
        RECT 42.200 26.100 42.600 26.200 ;
        RECT 36.600 25.800 42.600 26.100 ;
        RECT 50.200 26.100 50.600 26.200 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 73.400 26.100 73.800 26.200 ;
        RECT 76.600 26.100 77.000 26.200 ;
        RECT 50.200 25.800 52.900 26.100 ;
        RECT 58.200 25.800 60.100 26.100 ;
        RECT 71.000 25.800 77.000 26.100 ;
        RECT 78.200 26.100 78.600 26.200 ;
        RECT 80.600 26.100 81.000 26.200 ;
        RECT 78.200 25.800 81.000 26.100 ;
        RECT 83.800 26.100 84.100 26.800 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 83.800 25.800 89.800 26.100 ;
        RECT 95.800 26.100 96.200 26.200 ;
        RECT 99.800 26.100 100.100 26.800 ;
        RECT 95.800 25.800 100.100 26.100 ;
        RECT 107.800 26.100 108.200 26.200 ;
        RECT 110.200 26.100 110.600 26.200 ;
        RECT 107.800 25.800 110.600 26.100 ;
        RECT 113.400 26.100 113.800 26.200 ;
        RECT 115.000 26.100 115.400 26.200 ;
        RECT 113.400 25.800 115.400 26.100 ;
        RECT 128.600 26.100 128.900 26.800 ;
        RECT 216.600 26.200 216.900 26.800 ;
        RECT 130.200 26.100 130.600 26.200 ;
        RECT 156.600 26.100 157.000 26.200 ;
        RECT 128.600 25.800 157.000 26.100 ;
        RECT 160.600 26.100 161.000 26.200 ;
        RECT 161.400 26.100 161.800 26.200 ;
        RECT 163.000 26.100 163.400 26.200 ;
        RECT 160.600 25.800 163.400 26.100 ;
        RECT 166.200 26.100 166.600 26.200 ;
        RECT 169.400 26.100 169.800 26.200 ;
        RECT 166.200 25.800 169.800 26.100 ;
        RECT 183.000 26.100 183.400 26.200 ;
        RECT 184.600 26.100 185.000 26.200 ;
        RECT 183.000 25.800 185.000 26.100 ;
        RECT 193.400 26.100 193.800 26.200 ;
        RECT 200.600 26.100 201.000 26.200 ;
        RECT 205.400 26.100 205.800 26.200 ;
        RECT 193.400 25.800 197.700 26.100 ;
        RECT 200.600 25.800 205.800 26.100 ;
        RECT 209.400 26.100 209.800 26.200 ;
        RECT 216.600 26.100 217.000 26.200 ;
        RECT 209.400 25.800 217.000 26.100 ;
        RECT 234.200 26.100 234.600 26.200 ;
        RECT 244.600 26.100 245.000 26.200 ;
        RECT 234.200 25.800 245.000 26.100 ;
        RECT 251.800 25.800 252.200 26.200 ;
        RECT 52.600 25.200 52.900 25.800 ;
        RECT 59.800 25.200 60.100 25.800 ;
        RECT 197.400 25.200 197.700 25.800 ;
        RECT 251.800 25.200 252.100 25.800 ;
        RECT 11.000 25.100 11.400 25.200 ;
        RECT 14.200 25.100 14.600 25.200 ;
        RECT 10.200 24.800 14.600 25.100 ;
        RECT 52.600 24.800 53.000 25.200 ;
        RECT 59.800 25.100 60.200 25.200 ;
        RECT 60.600 25.100 61.000 25.200 ;
        RECT 59.800 24.800 61.000 25.100 ;
        RECT 139.800 25.100 140.200 25.200 ;
        RECT 182.200 25.100 182.600 25.200 ;
        RECT 186.200 25.100 186.600 25.200 ;
        RECT 192.600 25.100 193.000 25.200 ;
        RECT 139.800 24.800 182.600 25.100 ;
        RECT 185.400 24.800 193.000 25.100 ;
        RECT 197.400 24.800 197.800 25.200 ;
        RECT 215.000 25.100 215.400 25.200 ;
        RECT 223.800 25.100 224.200 25.200 ;
        RECT 215.000 24.800 224.200 25.100 ;
        RECT 251.800 24.800 252.200 25.200 ;
        RECT 55.000 24.100 55.400 24.200 ;
        RECT 60.600 24.100 61.000 24.200 ;
        RECT 55.000 23.800 61.000 24.100 ;
        RECT 116.600 24.100 117.000 24.200 ;
        RECT 125.400 24.100 125.800 24.200 ;
        RECT 143.000 24.100 143.400 24.200 ;
        RECT 116.600 23.800 143.400 24.100 ;
        RECT 143.800 24.100 144.200 24.200 ;
        RECT 165.400 24.100 165.800 24.200 ;
        RECT 143.800 23.800 165.800 24.100 ;
        RECT 196.600 24.100 197.000 24.200 ;
        RECT 229.400 24.100 229.800 24.200 ;
        RECT 196.600 23.800 229.800 24.100 ;
        RECT 240.600 24.100 241.000 24.200 ;
        RECT 251.800 24.100 252.200 24.200 ;
        RECT 240.600 23.800 252.200 24.100 ;
        RECT 41.400 23.100 41.800 23.200 ;
        RECT 61.400 23.100 61.800 23.200 ;
        RECT 41.400 22.800 61.800 23.100 ;
        RECT 64.600 23.100 65.000 23.200 ;
        RECT 107.800 23.100 108.200 23.200 ;
        RECT 154.200 23.100 154.600 23.200 ;
        RECT 172.600 23.100 173.000 23.200 ;
        RECT 64.600 22.800 173.000 23.100 ;
        RECT 191.000 23.100 191.400 23.200 ;
        RECT 211.800 23.100 212.200 23.200 ;
        RECT 191.000 22.800 212.200 23.100 ;
        RECT 17.400 21.800 17.800 22.200 ;
        RECT 47.000 22.100 47.400 22.200 ;
        RECT 87.800 22.100 88.200 22.200 ;
        RECT 47.000 21.800 88.200 22.100 ;
        RECT 126.200 22.100 126.600 22.200 ;
        RECT 129.400 22.100 129.800 22.200 ;
        RECT 126.200 21.800 129.800 22.100 ;
        RECT 137.400 22.100 137.800 22.200 ;
        RECT 183.800 22.100 184.200 22.200 ;
        RECT 137.400 21.800 184.200 22.100 ;
        RECT 17.400 21.200 17.700 21.800 ;
        RECT 17.400 20.800 17.800 21.200 ;
        RECT 70.200 21.100 70.600 21.200 ;
        RECT 71.000 21.100 71.400 21.200 ;
        RECT 95.000 21.100 95.400 21.200 ;
        RECT 70.200 20.800 95.400 21.100 ;
        RECT 159.800 21.100 160.200 21.200 ;
        RECT 170.200 21.100 170.600 21.200 ;
        RECT 174.200 21.100 174.600 21.200 ;
        RECT 159.800 20.800 174.600 21.100 ;
        RECT 88.600 19.800 89.000 20.200 ;
        RECT 156.600 20.100 157.000 20.200 ;
        RECT 221.400 20.100 221.800 20.200 ;
        RECT 223.800 20.100 224.200 20.200 ;
        RECT 156.600 19.800 224.200 20.100 ;
        RECT 88.600 19.200 88.900 19.800 ;
        RECT 43.000 19.100 43.400 19.200 ;
        RECT 43.800 19.100 44.200 19.200 ;
        RECT 43.000 18.800 44.200 19.100 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 111.800 19.100 112.200 19.200 ;
        RECT 112.600 19.100 113.000 19.200 ;
        RECT 111.800 18.800 113.000 19.100 ;
        RECT 138.200 19.100 138.600 19.200 ;
        RECT 143.800 19.100 144.200 19.200 ;
        RECT 146.200 19.100 146.600 19.200 ;
        RECT 138.200 18.800 146.600 19.100 ;
        RECT 171.800 19.100 172.200 19.200 ;
        RECT 173.400 19.100 173.800 19.200 ;
        RECT 175.000 19.100 175.400 19.200 ;
        RECT 171.800 18.800 175.400 19.100 ;
        RECT 48.600 18.100 49.000 18.200 ;
        RECT 64.600 18.100 65.000 18.200 ;
        RECT 48.600 17.800 65.000 18.100 ;
        RECT 107.000 18.100 107.400 18.200 ;
        RECT 128.600 18.100 129.000 18.200 ;
        RECT 159.800 18.100 160.200 18.200 ;
        RECT 163.000 18.100 163.400 18.200 ;
        RECT 107.000 17.800 129.000 18.100 ;
        RECT 159.000 17.800 163.400 18.100 ;
        RECT 172.600 18.100 173.000 18.200 ;
        RECT 206.200 18.100 206.600 18.200 ;
        RECT 215.000 18.100 215.400 18.200 ;
        RECT 172.600 17.800 215.400 18.100 ;
        RECT 10.200 17.100 10.600 17.200 ;
        RECT 15.800 17.100 16.200 17.200 ;
        RECT 10.200 16.800 16.200 17.100 ;
        RECT 26.200 17.100 26.600 17.200 ;
        RECT 33.400 17.100 33.800 17.200 ;
        RECT 53.400 17.100 53.800 17.200 ;
        RECT 26.200 16.800 53.800 17.100 ;
        RECT 62.200 17.100 62.600 17.200 ;
        RECT 64.600 17.100 65.000 17.200 ;
        RECT 97.400 17.100 97.800 17.200 ;
        RECT 62.200 16.800 97.800 17.100 ;
        RECT 108.600 17.100 109.000 17.200 ;
        RECT 113.400 17.100 113.800 17.200 ;
        RECT 108.600 16.800 113.800 17.100 ;
        RECT 129.400 17.100 129.800 17.200 ;
        RECT 138.200 17.100 138.600 17.200 ;
        RECT 129.400 16.800 138.600 17.100 ;
        RECT 158.200 17.100 158.600 17.200 ;
        RECT 159.800 17.100 160.200 17.200 ;
        RECT 164.600 17.100 165.000 17.200 ;
        RECT 158.200 16.800 165.000 17.100 ;
        RECT 190.200 17.100 190.600 17.200 ;
        RECT 199.000 17.100 199.400 17.200 ;
        RECT 190.200 16.800 199.400 17.100 ;
        RECT 7.000 16.100 7.400 16.200 ;
        RECT 12.600 16.100 13.000 16.200 ;
        RECT 7.000 15.800 13.000 16.100 ;
        RECT 15.000 16.100 15.400 16.200 ;
        RECT 17.400 16.100 17.800 16.200 ;
        RECT 15.000 15.800 17.800 16.100 ;
        RECT 26.200 15.800 26.600 16.200 ;
        RECT 65.400 15.800 65.800 16.200 ;
        RECT 80.600 16.100 81.000 16.200 ;
        RECT 99.800 16.100 100.200 16.200 ;
        RECT 80.600 15.800 100.200 16.100 ;
        RECT 103.000 16.100 103.400 16.200 ;
        RECT 103.800 16.100 104.200 16.200 ;
        RECT 103.000 15.800 104.200 16.100 ;
        RECT 109.400 16.100 109.800 16.200 ;
        RECT 110.200 16.100 110.600 16.200 ;
        RECT 112.600 16.100 113.000 16.200 ;
        RECT 139.000 16.100 139.400 16.200 ;
        RECT 109.400 15.800 139.400 16.100 ;
        RECT 141.400 16.100 141.800 16.200 ;
        RECT 143.000 16.100 143.400 16.200 ;
        RECT 141.400 15.800 143.400 16.100 ;
        RECT 146.200 16.100 146.600 16.200 ;
        RECT 186.200 16.100 186.600 16.200 ;
        RECT 187.800 16.100 188.200 16.200 ;
        RECT 146.200 15.800 188.200 16.100 ;
        RECT 210.200 15.800 210.600 16.200 ;
        RECT 213.400 16.100 213.800 16.200 ;
        RECT 225.400 16.100 225.800 16.200 ;
        RECT 213.400 15.800 225.800 16.100 ;
        RECT 240.600 16.100 241.000 16.200 ;
        RECT 249.400 16.100 249.800 16.200 ;
        RECT 240.600 15.800 249.800 16.100 ;
        RECT 0.600 15.100 1.000 15.200 ;
        RECT 10.200 15.100 10.600 15.200 ;
        RECT 11.000 15.100 11.400 15.200 ;
        RECT 0.600 14.800 11.400 15.100 ;
        RECT 11.800 15.100 12.200 15.200 ;
        RECT 15.000 15.100 15.400 15.200 ;
        RECT 19.000 15.100 19.400 15.200 ;
        RECT 11.800 14.800 19.400 15.100 ;
        RECT 20.600 15.100 21.000 15.200 ;
        RECT 26.200 15.100 26.500 15.800 ;
        RECT 20.600 14.800 26.500 15.100 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 61.400 15.100 61.800 15.200 ;
        RECT 65.400 15.100 65.700 15.800 ;
        RECT 61.400 14.800 65.700 15.100 ;
        RECT 71.800 14.800 72.200 15.200 ;
        RECT 82.200 15.100 82.600 15.200 ;
        RECT 83.800 15.100 84.200 15.200 ;
        RECT 101.400 15.100 101.800 15.200 ;
        RECT 108.600 15.100 109.000 15.200 ;
        RECT 119.000 15.100 119.400 15.200 ;
        RECT 131.800 15.100 132.200 15.200 ;
        RECT 82.200 14.800 101.800 15.100 ;
        RECT 102.200 14.800 109.000 15.100 ;
        RECT 111.800 14.800 119.400 15.100 ;
        RECT 123.800 14.800 132.200 15.100 ;
        RECT 139.800 15.100 140.200 15.200 ;
        RECT 143.000 15.100 143.400 15.200 ;
        RECT 139.800 14.800 143.400 15.100 ;
        RECT 151.800 15.100 152.200 15.200 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 151.800 14.800 155.400 15.100 ;
        RECT 156.600 15.100 157.000 15.200 ;
        RECT 158.200 15.100 158.600 15.200 ;
        RECT 156.600 14.800 158.600 15.100 ;
        RECT 172.600 15.100 173.000 15.200 ;
        RECT 179.800 15.100 180.200 15.200 ;
        RECT 172.600 14.800 180.200 15.100 ;
        RECT 183.800 15.100 184.200 15.200 ;
        RECT 191.800 15.100 192.200 15.200 ;
        RECT 183.800 14.800 192.200 15.100 ;
        RECT 204.600 15.100 205.000 15.200 ;
        RECT 210.200 15.100 210.500 15.800 ;
        RECT 204.600 14.800 210.500 15.100 ;
        RECT 215.000 15.100 215.400 15.200 ;
        RECT 215.800 15.100 216.200 15.200 ;
        RECT 218.200 15.100 218.600 15.200 ;
        RECT 215.000 14.800 218.600 15.100 ;
        RECT 223.800 15.100 224.200 15.200 ;
        RECT 231.000 15.100 231.400 15.200 ;
        RECT 223.800 14.800 231.400 15.100 ;
        RECT 234.200 14.800 234.600 15.200 ;
        RECT 235.800 14.800 236.200 15.200 ;
        RECT 14.200 14.100 14.600 14.200 ;
        RECT 15.000 14.100 15.400 14.200 ;
        RECT 14.200 13.800 15.400 14.100 ;
        RECT 19.800 14.100 20.200 14.200 ;
        RECT 21.400 14.100 21.800 14.200 ;
        RECT 19.800 13.800 21.800 14.100 ;
        RECT 59.800 14.100 60.100 14.800 ;
        RECT 71.800 14.100 72.100 14.800 ;
        RECT 102.200 14.200 102.500 14.800 ;
        RECT 111.800 14.200 112.100 14.800 ;
        RECT 123.800 14.200 124.100 14.800 ;
        RECT 59.800 13.800 72.100 14.100 ;
        RECT 74.200 14.100 74.600 14.200 ;
        RECT 83.000 14.100 83.400 14.200 ;
        RECT 74.200 13.800 83.400 14.100 ;
        RECT 102.200 13.800 102.600 14.200 ;
        RECT 111.800 13.800 112.200 14.200 ;
        RECT 112.600 14.100 113.000 14.200 ;
        RECT 113.400 14.100 113.800 14.200 ;
        RECT 112.600 13.800 113.800 14.100 ;
        RECT 123.800 13.800 124.200 14.200 ;
        RECT 134.200 14.100 134.600 14.200 ;
        RECT 140.600 14.100 141.000 14.200 ;
        RECT 134.200 13.800 141.000 14.100 ;
        RECT 143.000 14.100 143.400 14.200 ;
        RECT 144.600 14.100 145.000 14.200 ;
        RECT 143.000 13.800 145.000 14.100 ;
        RECT 155.000 14.100 155.400 14.200 ;
        RECT 169.400 14.100 169.800 14.200 ;
        RECT 155.000 13.800 169.800 14.100 ;
        RECT 171.000 14.100 171.400 14.200 ;
        RECT 174.200 14.100 174.600 14.200 ;
        RECT 171.000 13.800 174.600 14.100 ;
        RECT 186.200 14.100 186.600 14.200 ;
        RECT 195.000 14.100 195.400 14.200 ;
        RECT 207.800 14.100 208.200 14.200 ;
        RECT 214.200 14.100 214.600 14.200 ;
        RECT 221.400 14.100 221.800 14.200 ;
        RECT 186.200 13.800 221.800 14.100 ;
        RECT 234.200 14.100 234.500 14.800 ;
        RECT 235.800 14.100 236.100 14.800 ;
        RECT 234.200 13.800 236.100 14.100 ;
        RECT 7.000 13.100 7.400 13.200 ;
        RECT 24.600 13.100 25.000 13.200 ;
        RECT 34.200 13.100 34.600 13.200 ;
        RECT 7.000 12.800 34.600 13.100 ;
        RECT 69.400 13.100 69.800 13.200 ;
        RECT 78.200 13.100 78.600 13.200 ;
        RECT 69.400 12.800 78.600 13.100 ;
        RECT 100.600 13.100 101.000 13.200 ;
        RECT 124.600 13.100 125.000 13.200 ;
        RECT 100.600 12.800 125.000 13.100 ;
        RECT 127.800 13.100 128.200 13.200 ;
        RECT 149.400 13.100 149.800 13.200 ;
        RECT 194.200 13.100 194.600 13.200 ;
        RECT 127.800 12.800 149.800 13.100 ;
        RECT 187.800 12.800 194.600 13.100 ;
        RECT 200.600 13.100 201.000 13.200 ;
        RECT 205.400 13.100 205.800 13.200 ;
        RECT 200.600 12.800 205.800 13.100 ;
        RECT 211.000 13.100 211.400 13.200 ;
        RECT 227.000 13.100 227.400 13.200 ;
        RECT 211.000 12.800 227.400 13.100 ;
        RECT 187.800 12.200 188.100 12.800 ;
        RECT 23.000 12.100 23.400 12.200 ;
        RECT 31.800 12.100 32.200 12.200 ;
        RECT 35.800 12.100 36.200 12.200 ;
        RECT 23.000 11.800 36.200 12.100 ;
        RECT 56.600 12.100 57.000 12.200 ;
        RECT 65.400 12.100 65.800 12.200 ;
        RECT 71.000 12.100 71.400 12.200 ;
        RECT 56.600 11.800 71.400 12.100 ;
        RECT 75.000 12.100 75.400 12.200 ;
        RECT 91.000 12.100 91.400 12.200 ;
        RECT 100.600 12.100 101.000 12.200 ;
        RECT 75.000 11.800 101.000 12.100 ;
        RECT 103.800 12.100 104.200 12.200 ;
        RECT 120.600 12.100 121.000 12.200 ;
        RECT 103.800 11.800 121.000 12.100 ;
        RECT 122.200 12.100 122.600 12.200 ;
        RECT 132.600 12.100 133.000 12.200 ;
        RECT 122.200 11.800 133.000 12.100 ;
        RECT 139.800 12.100 140.200 12.200 ;
        RECT 144.600 12.100 145.000 12.200 ;
        RECT 139.800 11.800 145.000 12.100 ;
        RECT 187.800 11.800 188.200 12.200 ;
        RECT 119.800 11.100 120.200 11.200 ;
        RECT 133.400 11.100 133.800 11.200 ;
        RECT 119.800 10.800 133.800 11.100 ;
        RECT 136.600 11.100 137.000 11.200 ;
        RECT 163.800 11.100 164.200 11.200 ;
        RECT 136.600 10.800 164.200 11.100 ;
        RECT 17.400 10.100 17.800 10.200 ;
        RECT 27.000 10.100 27.400 10.200 ;
        RECT 44.600 10.100 45.000 10.200 ;
        RECT 17.400 9.800 45.000 10.100 ;
        RECT 101.400 10.100 101.800 10.200 ;
        RECT 128.600 10.100 129.000 10.200 ;
        RECT 137.400 10.100 137.800 10.200 ;
        RECT 101.400 9.800 137.800 10.100 ;
        RECT 139.000 10.100 139.400 10.200 ;
        RECT 145.400 10.100 145.800 10.200 ;
        RECT 152.600 10.100 153.000 10.200 ;
        RECT 139.000 9.800 153.000 10.100 ;
        RECT 205.400 10.100 205.800 10.200 ;
        RECT 211.000 10.100 211.400 10.200 ;
        RECT 205.400 9.800 211.400 10.100 ;
        RECT 29.400 9.100 29.800 9.200 ;
        RECT 33.400 9.100 33.800 9.200 ;
        RECT 41.400 9.100 41.800 9.200 ;
        RECT 29.400 8.800 41.800 9.100 ;
        RECT 43.000 9.100 43.400 9.200 ;
        RECT 69.400 9.100 69.800 9.200 ;
        RECT 43.000 8.800 69.800 9.100 ;
        RECT 71.000 9.100 71.400 9.200 ;
        RECT 81.400 9.100 81.800 9.200 ;
        RECT 87.000 9.100 87.400 9.200 ;
        RECT 107.000 9.100 107.400 9.200 ;
        RECT 127.000 9.100 127.400 9.200 ;
        RECT 129.400 9.100 129.800 9.200 ;
        RECT 143.000 9.100 143.400 9.200 ;
        RECT 71.000 8.800 87.400 9.100 ;
        RECT 89.400 8.800 143.400 9.100 ;
        RECT 153.400 9.100 153.800 9.200 ;
        RECT 167.800 9.100 168.200 9.200 ;
        RECT 169.400 9.100 169.800 9.200 ;
        RECT 153.400 8.800 169.800 9.100 ;
        RECT 181.400 9.100 181.800 9.200 ;
        RECT 193.400 9.100 193.800 9.200 ;
        RECT 181.400 8.800 193.800 9.100 ;
        RECT 209.400 9.100 209.800 9.200 ;
        RECT 243.800 9.100 244.200 9.200 ;
        RECT 209.400 8.800 244.200 9.100 ;
        RECT 246.200 9.100 246.600 9.200 ;
        RECT 247.800 9.100 248.200 9.200 ;
        RECT 246.200 8.800 248.200 9.100 ;
        RECT 89.400 8.200 89.700 8.800 ;
        RECT 21.400 8.100 21.800 8.200 ;
        RECT 27.800 8.100 28.200 8.200 ;
        RECT 31.800 8.100 32.200 8.200 ;
        RECT 35.800 8.100 36.200 8.200 ;
        RECT 21.400 7.800 36.200 8.100 ;
        RECT 58.200 7.800 58.600 8.200 ;
        RECT 73.400 7.800 73.800 8.200 ;
        RECT 89.400 7.800 89.800 8.200 ;
        RECT 95.800 8.100 96.200 8.200 ;
        RECT 107.800 8.100 108.200 8.200 ;
        RECT 95.800 7.800 108.200 8.100 ;
        RECT 143.000 8.100 143.400 8.200 ;
        RECT 159.800 8.100 160.200 8.200 ;
        RECT 143.000 7.800 160.200 8.100 ;
        RECT 178.200 8.100 178.600 8.200 ;
        RECT 189.400 8.100 189.800 8.200 ;
        RECT 206.200 8.100 206.600 8.200 ;
        RECT 215.800 8.100 216.200 8.200 ;
        RECT 222.200 8.100 222.600 8.200 ;
        RECT 235.000 8.100 235.400 8.200 ;
        RECT 178.200 7.800 235.400 8.100 ;
        RECT 11.800 7.100 12.200 7.200 ;
        RECT 14.200 7.100 14.600 7.200 ;
        RECT 32.600 7.100 33.000 7.200 ;
        RECT 43.800 7.100 44.200 7.200 ;
        RECT 11.800 6.800 44.200 7.100 ;
        RECT 45.400 7.100 45.800 7.200 ;
        RECT 55.800 7.100 56.200 7.200 ;
        RECT 45.400 6.800 56.200 7.100 ;
        RECT 58.200 7.100 58.500 7.800 ;
        RECT 73.400 7.100 73.700 7.800 ;
        RECT 58.200 6.800 73.700 7.100 ;
        RECT 75.800 7.100 76.200 7.200 ;
        RECT 84.600 7.100 85.000 7.200 ;
        RECT 75.800 6.800 85.000 7.100 ;
        RECT 86.200 7.100 86.600 7.200 ;
        RECT 111.000 7.100 111.400 7.200 ;
        RECT 118.200 7.100 118.600 7.200 ;
        RECT 127.000 7.100 127.400 7.200 ;
        RECT 86.200 6.800 111.400 7.100 ;
        RECT 114.200 6.800 116.100 7.100 ;
        RECT 118.200 6.800 127.400 7.100 ;
        RECT 133.400 7.100 133.800 7.200 ;
        RECT 140.600 7.100 141.000 7.200 ;
        RECT 133.400 6.800 141.000 7.100 ;
        RECT 143.800 6.800 144.200 7.200 ;
        RECT 161.400 7.100 161.800 7.200 ;
        RECT 155.800 6.800 161.800 7.100 ;
        RECT 167.000 7.100 167.400 7.200 ;
        RECT 175.800 7.100 176.200 7.200 ;
        RECT 167.000 6.800 176.200 7.100 ;
        RECT 180.600 7.100 181.000 7.200 ;
        RECT 183.800 7.100 184.200 7.200 ;
        RECT 196.600 7.100 197.000 7.200 ;
        RECT 180.600 6.800 197.000 7.100 ;
        RECT 197.400 7.100 197.800 7.200 ;
        RECT 204.600 7.100 205.000 7.200 ;
        RECT 197.400 6.800 205.000 7.100 ;
        RECT 223.800 7.100 224.200 7.200 ;
        RECT 232.600 7.100 233.000 7.200 ;
        RECT 223.800 6.800 233.000 7.100 ;
        RECT 235.000 7.100 235.300 7.800 ;
        RECT 242.200 7.100 242.600 7.200 ;
        RECT 235.000 6.800 242.600 7.100 ;
        RECT 243.800 7.100 244.200 7.200 ;
        RECT 247.000 7.100 247.400 7.200 ;
        RECT 243.800 6.800 247.400 7.100 ;
        RECT 14.200 6.100 14.600 6.200 ;
        RECT 17.400 6.100 17.800 6.200 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 14.200 5.800 19.400 6.100 ;
        RECT 19.800 6.100 20.200 6.200 ;
        RECT 43.000 6.100 43.400 6.200 ;
        RECT 46.200 6.100 46.600 6.200 ;
        RECT 19.800 5.800 46.600 6.100 ;
        RECT 67.800 6.100 68.200 6.200 ;
        RECT 68.600 6.100 69.000 6.200 ;
        RECT 67.800 5.800 69.000 6.100 ;
        RECT 69.400 6.100 69.800 6.200 ;
        RECT 87.000 6.100 87.400 6.200 ;
        RECT 69.400 5.800 87.400 6.100 ;
        RECT 96.600 6.100 97.000 6.300 ;
        RECT 114.200 6.200 114.500 6.800 ;
        RECT 115.800 6.200 116.100 6.800 ;
        RECT 143.800 6.200 144.100 6.800 ;
        RECT 155.800 6.200 156.100 6.800 ;
        RECT 157.400 6.200 157.700 6.800 ;
        RECT 103.800 6.100 104.200 6.200 ;
        RECT 96.600 5.800 104.200 6.100 ;
        RECT 107.000 6.100 107.400 6.200 ;
        RECT 108.600 6.100 109.000 6.200 ;
        RECT 107.000 5.800 109.000 6.100 ;
        RECT 110.200 6.100 110.600 6.200 ;
        RECT 114.200 6.100 114.600 6.200 ;
        RECT 110.200 5.800 114.600 6.100 ;
        RECT 115.800 5.800 116.200 6.200 ;
        RECT 126.200 6.100 126.600 6.200 ;
        RECT 128.600 6.100 129.000 6.200 ;
        RECT 126.200 5.800 129.000 6.100 ;
        RECT 139.800 6.100 140.200 6.200 ;
        RECT 140.600 6.100 141.000 6.200 ;
        RECT 139.800 5.800 141.000 6.100 ;
        RECT 143.800 5.800 144.200 6.200 ;
        RECT 147.000 6.100 147.400 6.200 ;
        RECT 152.600 6.100 153.000 6.200 ;
        RECT 147.000 5.800 153.000 6.100 ;
        RECT 155.800 5.800 156.200 6.200 ;
        RECT 157.400 5.800 157.800 6.200 ;
        RECT 165.400 6.100 165.800 6.200 ;
        RECT 169.400 6.100 169.800 6.200 ;
        RECT 221.400 6.100 221.800 6.200 ;
        RECT 224.600 6.100 225.000 6.200 ;
        RECT 165.400 5.800 225.000 6.100 ;
        RECT 16.600 5.100 17.000 5.200 ;
        RECT 20.600 5.100 21.000 5.200 ;
        RECT 16.600 4.800 21.000 5.100 ;
        RECT 31.000 5.100 31.400 5.200 ;
        RECT 35.800 5.100 36.200 5.200 ;
        RECT 31.000 4.800 36.200 5.100 ;
        RECT 84.600 5.100 85.000 5.200 ;
        RECT 86.200 5.100 86.600 5.200 ;
        RECT 84.600 4.800 86.600 5.100 ;
        RECT 104.600 5.100 105.000 5.200 ;
        RECT 106.200 5.100 106.600 5.200 ;
        RECT 141.400 5.100 141.800 5.200 ;
        RECT 180.600 5.100 181.000 5.200 ;
        RECT 187.800 5.100 188.200 5.200 ;
        RECT 104.600 4.800 181.000 5.100 ;
        RECT 183.800 4.800 188.200 5.100 ;
        RECT 183.800 4.200 184.100 4.800 ;
        RECT 183.800 3.800 184.200 4.200 ;
        RECT 111.000 3.100 111.400 3.200 ;
        RECT 195.800 3.100 196.200 3.200 ;
        RECT 198.200 3.100 198.600 3.200 ;
        RECT 111.000 2.800 198.600 3.100 ;
      LAYER via3 ;
        RECT 238.200 235.800 238.600 236.200 ;
        RECT 231.000 234.800 231.400 235.200 ;
        RECT 4.600 233.800 5.000 234.200 ;
        RECT 119.000 233.800 119.400 234.200 ;
        RECT 34.200 232.800 34.600 233.200 ;
        RECT 233.400 231.800 233.800 232.200 ;
        RECT 76.600 230.800 77.000 231.200 ;
        RECT 181.400 230.800 181.800 231.200 ;
        RECT 97.400 229.800 97.800 230.200 ;
        RECT 135.800 229.800 136.200 230.200 ;
        RECT 91.000 227.800 91.400 228.200 ;
        RECT 235.800 227.800 236.200 228.200 ;
        RECT 122.200 226.800 122.600 227.200 ;
        RECT 39.000 225.800 39.400 226.200 ;
        RECT 144.600 225.800 145.000 226.200 ;
        RECT 197.400 225.800 197.800 226.200 ;
        RECT 215.800 225.800 216.200 226.200 ;
        RECT 43.800 224.800 44.200 225.200 ;
        RECT 110.200 224.800 110.600 225.200 ;
        RECT 228.600 224.800 229.000 225.200 ;
        RECT 105.400 223.800 105.800 224.200 ;
        RECT 244.600 223.800 245.000 224.200 ;
        RECT 134.200 222.800 134.600 223.200 ;
        RECT 235.000 222.800 235.400 223.200 ;
        RECT 57.400 221.800 57.800 222.200 ;
        RECT 69.400 219.800 69.800 220.200 ;
        RECT 106.200 219.800 106.600 220.200 ;
        RECT 211.800 218.800 212.200 219.200 ;
        RECT 182.200 217.800 182.600 218.200 ;
        RECT 212.600 216.800 213.000 217.200 ;
        RECT 237.400 215.800 237.800 216.200 ;
        RECT 11.000 214.800 11.400 215.200 ;
        RECT 100.600 214.800 101.000 215.200 ;
        RECT 131.000 214.800 131.400 215.200 ;
        RECT 185.400 214.800 185.800 215.200 ;
        RECT 94.200 210.800 94.600 211.200 ;
        RECT 73.400 208.800 73.800 209.200 ;
        RECT 169.400 208.800 169.800 209.200 ;
        RECT 145.400 207.800 145.800 208.200 ;
        RECT 112.600 205.800 113.000 206.200 ;
        RECT 199.800 205.800 200.200 206.200 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 193.400 204.800 193.800 205.200 ;
        RECT 102.200 203.800 102.600 204.200 ;
        RECT 115.800 202.800 116.200 203.200 ;
        RECT 50.200 201.800 50.600 202.200 ;
        RECT 23.000 198.800 23.400 199.200 ;
        RECT 75.000 198.800 75.400 199.200 ;
        RECT 140.600 197.800 141.000 198.200 ;
        RECT 236.600 197.800 237.000 198.200 ;
        RECT 251.800 196.800 252.200 197.200 ;
        RECT 165.400 195.800 165.800 196.200 ;
        RECT 219.800 195.800 220.200 196.200 ;
        RECT 60.600 194.800 61.000 195.200 ;
        RECT 63.000 194.800 63.400 195.200 ;
        RECT 143.800 194.800 144.200 195.200 ;
        RECT 215.800 194.800 216.200 195.200 ;
        RECT 65.400 193.800 65.800 194.200 ;
        RECT 143.800 193.800 144.200 194.200 ;
        RECT 246.200 193.800 246.600 194.200 ;
        RECT 63.800 192.800 64.200 193.200 ;
        RECT 231.800 190.800 232.200 191.200 ;
        RECT 74.200 186.800 74.600 187.200 ;
        RECT 117.400 186.800 117.800 187.200 ;
        RECT 148.600 186.800 149.000 187.200 ;
        RECT 175.000 186.800 175.400 187.200 ;
        RECT 35.000 185.800 35.400 186.200 ;
        RECT 57.400 185.800 57.800 186.200 ;
        RECT 218.200 185.800 218.600 186.200 ;
        RECT 158.200 184.800 158.600 185.200 ;
        RECT 241.400 184.800 241.800 185.200 ;
        RECT 38.200 183.800 38.600 184.200 ;
        RECT 107.000 183.800 107.400 184.200 ;
        RECT 183.000 183.800 183.400 184.200 ;
        RECT 85.400 181.800 85.800 182.200 ;
        RECT 248.600 181.800 249.000 182.200 ;
        RECT 105.400 180.800 105.800 181.200 ;
        RECT 223.000 179.800 223.400 180.200 ;
        RECT 51.000 178.800 51.400 179.200 ;
        RECT 210.200 178.800 210.600 179.200 ;
        RECT 182.200 177.800 182.600 178.200 ;
        RECT 185.400 177.800 185.800 178.200 ;
        RECT 31.800 176.800 32.200 177.200 ;
        RECT 16.600 175.800 17.000 176.200 ;
        RECT 19.000 175.800 19.400 176.200 ;
        RECT 147.800 175.800 148.200 176.200 ;
        RECT 150.200 175.800 150.600 176.200 ;
        RECT 237.400 175.800 237.800 176.200 ;
        RECT 251.000 175.800 251.400 176.200 ;
        RECT 86.200 174.800 86.600 175.200 ;
        RECT 96.600 174.800 97.000 175.200 ;
        RECT 133.400 174.800 133.800 175.200 ;
        RECT 175.800 174.800 176.200 175.200 ;
        RECT 225.400 174.800 225.800 175.200 ;
        RECT 123.000 173.800 123.400 174.200 ;
        RECT 20.600 172.800 21.000 173.200 ;
        RECT 79.000 171.800 79.400 172.200 ;
        RECT 123.800 171.800 124.200 172.200 ;
        RECT 211.000 171.800 211.400 172.200 ;
        RECT 240.600 171.800 241.000 172.200 ;
        RECT 192.600 170.800 193.000 171.200 ;
        RECT 103.800 169.800 104.200 170.200 ;
        RECT 243.800 169.800 244.200 170.200 ;
        RECT 94.200 166.800 94.600 167.200 ;
        RECT 222.200 166.800 222.600 167.200 ;
        RECT 17.400 165.800 17.800 166.200 ;
        RECT 84.600 164.800 85.000 165.200 ;
        RECT 155.000 164.800 155.400 165.200 ;
        RECT 116.600 163.800 117.000 164.200 ;
        RECT 195.800 162.800 196.200 163.200 ;
        RECT 58.200 161.800 58.600 162.200 ;
        RECT 237.400 161.800 237.800 162.200 ;
        RECT 132.600 159.800 133.000 160.200 ;
        RECT 184.600 158.800 185.000 159.200 ;
        RECT 171.800 156.800 172.200 157.200 ;
        RECT 29.400 155.800 29.800 156.200 ;
        RECT 143.800 155.800 144.200 156.200 ;
        RECT 248.600 154.800 249.000 155.200 ;
        RECT 105.400 153.800 105.800 154.200 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 74.200 150.800 74.600 151.200 ;
        RECT 67.800 148.800 68.200 149.200 ;
        RECT 221.400 147.800 221.800 148.200 ;
        RECT 135.800 146.800 136.200 147.200 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 14.200 145.800 14.600 146.200 ;
        RECT 170.200 145.800 170.600 146.200 ;
        RECT 190.200 145.800 190.600 146.200 ;
        RECT 214.200 145.800 214.600 146.200 ;
        RECT 229.400 145.800 229.800 146.200 ;
        RECT 47.800 144.800 48.200 145.200 ;
        RECT 130.200 144.800 130.600 145.200 ;
        RECT 171.000 144.800 171.400 145.200 ;
        RECT 87.800 143.800 88.200 144.200 ;
        RECT 97.400 143.800 97.800 144.200 ;
        RECT 101.400 142.800 101.800 143.200 ;
        RECT 239.000 142.800 239.400 143.200 ;
        RECT 147.800 141.800 148.200 142.200 ;
        RECT 65.400 139.800 65.800 140.200 ;
        RECT 72.600 139.800 73.000 140.200 ;
        RECT 12.600 138.800 13.000 139.200 ;
        RECT 111.000 138.800 111.400 139.200 ;
        RECT 59.800 137.800 60.200 138.200 ;
        RECT 71.800 137.800 72.200 138.200 ;
        RECT 101.400 137.800 101.800 138.200 ;
        RECT 131.000 136.800 131.400 137.200 ;
        RECT 64.600 135.800 65.000 136.200 ;
        RECT 89.400 135.800 89.800 136.200 ;
        RECT 123.800 135.800 124.200 136.200 ;
        RECT 139.000 135.800 139.400 136.200 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 45.400 134.800 45.800 135.200 ;
        RECT 85.400 134.800 85.800 135.200 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 187.800 133.800 188.200 134.200 ;
        RECT 137.400 132.800 137.800 133.200 ;
        RECT 187.000 132.800 187.400 133.200 ;
        RECT 83.800 131.800 84.200 132.200 ;
        RECT 97.400 131.800 97.800 132.200 ;
        RECT 140.600 131.800 141.000 132.200 ;
        RECT 186.200 131.800 186.600 132.200 ;
        RECT 82.200 130.800 82.600 131.200 ;
        RECT 47.000 129.800 47.400 130.200 ;
        RECT 68.600 129.800 69.000 130.200 ;
        RECT 82.200 129.800 82.600 130.200 ;
        RECT 157.400 129.800 157.800 130.200 ;
        RECT 167.000 128.800 167.400 129.200 ;
        RECT 181.400 127.800 181.800 128.200 ;
        RECT 195.000 127.800 195.400 128.200 ;
        RECT 241.400 127.800 241.800 128.200 ;
        RECT 102.200 126.800 102.600 127.200 ;
        RECT 115.000 126.800 115.400 127.200 ;
        RECT 161.400 126.800 161.800 127.200 ;
        RECT 239.000 126.800 239.400 127.200 ;
        RECT 247.000 126.800 247.400 127.200 ;
        RECT 92.600 125.800 93.000 126.200 ;
        RECT 175.800 125.800 176.200 126.200 ;
        RECT 199.000 125.800 199.400 126.200 ;
        RECT 239.000 125.800 239.400 126.200 ;
        RECT 35.000 124.800 35.400 125.200 ;
        RECT 86.200 124.800 86.600 125.200 ;
        RECT 166.200 124.800 166.600 125.200 ;
        RECT 220.600 124.800 221.000 125.200 ;
        RECT 248.600 124.800 249.000 125.200 ;
        RECT 139.800 123.800 140.200 124.200 ;
        RECT 215.000 123.800 215.400 124.200 ;
        RECT 100.600 122.800 101.000 123.200 ;
        RECT 179.800 122.800 180.200 123.200 ;
        RECT 13.400 121.800 13.800 122.200 ;
        RECT 67.000 121.800 67.400 122.200 ;
        RECT 87.800 121.800 88.200 122.200 ;
        RECT 195.800 120.800 196.200 121.200 ;
        RECT 71.800 119.800 72.200 120.200 ;
        RECT 115.800 119.800 116.200 120.200 ;
        RECT 246.200 119.800 246.600 120.200 ;
        RECT 232.600 118.800 233.000 119.200 ;
        RECT 115.000 117.800 115.400 118.200 ;
        RECT 115.000 116.800 115.400 117.200 ;
        RECT 87.000 115.800 87.400 116.200 ;
        RECT 175.800 115.800 176.200 116.200 ;
        RECT 60.600 114.800 61.000 115.200 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 197.400 114.800 197.800 115.200 ;
        RECT 230.200 112.800 230.600 113.200 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 127.800 111.800 128.200 112.200 ;
        RECT 71.000 110.800 71.400 111.200 ;
        RECT 170.200 110.800 170.600 111.200 ;
        RECT 79.000 109.800 79.400 110.200 ;
        RECT 107.800 109.800 108.200 110.200 ;
        RECT 118.200 109.800 118.600 110.200 ;
        RECT 163.800 109.800 164.200 110.200 ;
        RECT 168.600 109.800 169.000 110.200 ;
        RECT 27.800 108.800 28.200 109.200 ;
        RECT 198.200 108.800 198.600 109.200 ;
        RECT 229.400 108.800 229.800 109.200 ;
        RECT 241.400 108.800 241.800 109.200 ;
        RECT 244.600 108.800 245.000 109.200 ;
        RECT 183.000 106.800 183.400 107.200 ;
        RECT 237.400 106.800 237.800 107.200 ;
        RECT 67.800 105.800 68.200 106.200 ;
        RECT 108.600 105.800 109.000 106.200 ;
        RECT 123.800 105.800 124.200 106.200 ;
        RECT 196.600 105.800 197.000 106.200 ;
        RECT 247.800 105.800 248.200 106.200 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 191.000 104.800 191.400 105.200 ;
        RECT 230.200 104.800 230.600 105.200 ;
        RECT 120.600 103.800 121.000 104.200 ;
        RECT 218.200 103.800 218.600 104.200 ;
        RECT 222.200 103.800 222.600 104.200 ;
        RECT 231.800 103.800 232.200 104.200 ;
        RECT 59.000 102.800 59.400 103.200 ;
        RECT 118.200 102.800 118.600 103.200 ;
        RECT 155.800 102.800 156.200 103.200 ;
        RECT 106.200 101.800 106.600 102.200 ;
        RECT 184.600 101.800 185.000 102.200 ;
        RECT 212.600 101.800 213.000 102.200 ;
        RECT 130.200 100.800 130.600 101.200 ;
        RECT 209.400 100.800 209.800 101.200 ;
        RECT 95.800 99.800 96.200 100.200 ;
        RECT 125.400 99.800 125.800 100.200 ;
        RECT 215.800 99.800 216.200 100.200 ;
        RECT 80.600 98.800 81.000 99.200 ;
        RECT 138.200 98.800 138.600 99.200 ;
        RECT 42.200 97.800 42.600 98.200 ;
        RECT 195.800 97.800 196.200 98.200 ;
        RECT 34.200 96.800 34.600 97.200 ;
        RECT 96.600 96.800 97.000 97.200 ;
        RECT 178.200 96.800 178.600 97.200 ;
        RECT 111.800 95.800 112.200 96.200 ;
        RECT 132.600 95.800 133.000 96.200 ;
        RECT 172.600 95.800 173.000 96.200 ;
        RECT 243.000 95.800 243.400 96.200 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 243.000 94.800 243.400 95.200 ;
        RECT 101.400 93.800 101.800 94.200 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 175.000 93.800 175.400 94.200 ;
        RECT 183.800 91.800 184.200 92.200 ;
        RECT 64.600 90.800 65.000 91.200 ;
        RECT 114.200 90.800 114.600 91.200 ;
        RECT 159.800 90.800 160.200 91.200 ;
        RECT 127.800 87.800 128.200 88.200 ;
        RECT 141.400 87.800 141.800 88.200 ;
        RECT 159.800 87.800 160.200 88.200 ;
        RECT 87.800 86.800 88.200 87.200 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 91.000 85.800 91.400 86.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 156.600 84.800 157.000 85.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 69.400 83.800 69.800 84.200 ;
        RECT 117.400 83.800 117.800 84.200 ;
        RECT 220.600 83.800 221.000 84.200 ;
        RECT 38.200 82.800 38.600 83.200 ;
        RECT 70.200 82.800 70.600 83.200 ;
        RECT 207.800 82.800 208.200 83.200 ;
        RECT 59.800 80.800 60.200 81.200 ;
        RECT 133.400 80.800 133.800 81.200 ;
        RECT 175.000 80.800 175.400 81.200 ;
        RECT 211.000 80.800 211.400 81.200 ;
        RECT 79.800 79.800 80.200 80.200 ;
        RECT 52.600 78.800 53.000 79.200 ;
        RECT 131.800 78.800 132.200 79.200 ;
        RECT 116.600 77.800 117.000 78.200 ;
        RECT 167.800 77.800 168.200 78.200 ;
        RECT 165.400 76.800 165.800 77.200 ;
        RECT 31.000 75.800 31.400 76.200 ;
        RECT 32.600 75.800 33.000 76.200 ;
        RECT 110.200 75.800 110.600 76.200 ;
        RECT 194.200 75.800 194.600 76.200 ;
        RECT 15.800 74.800 16.200 75.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 249.400 75.800 249.800 76.200 ;
        RECT 131.000 74.800 131.400 75.200 ;
        RECT 169.400 74.800 169.800 75.200 ;
        RECT 184.600 74.800 185.000 75.200 ;
        RECT 31.000 73.800 31.400 74.200 ;
        RECT 151.800 73.800 152.200 74.200 ;
        RECT 205.400 73.800 205.800 74.200 ;
        RECT 115.800 72.800 116.200 73.200 ;
        RECT 130.200 72.800 130.600 73.200 ;
        RECT 46.200 71.800 46.600 72.200 ;
        RECT 139.000 71.800 139.400 72.200 ;
        RECT 143.800 71.800 144.200 72.200 ;
        RECT 75.800 70.800 76.200 71.200 ;
        RECT 97.400 70.800 97.800 71.200 ;
        RECT 162.200 70.800 162.600 71.200 ;
        RECT 94.200 69.800 94.600 70.200 ;
        RECT 21.400 68.800 21.800 69.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 115.000 68.800 115.400 69.200 ;
        RECT 5.400 67.800 5.800 68.200 ;
        RECT 58.200 67.800 58.600 68.200 ;
        RECT 100.600 67.800 101.000 68.200 ;
        RECT 168.600 67.800 169.000 68.200 ;
        RECT 216.600 67.800 217.000 68.200 ;
        RECT 33.400 66.800 33.800 67.200 ;
        RECT 48.600 66.800 49.000 67.200 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 65.400 66.800 65.800 67.200 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 212.600 66.800 213.000 67.200 ;
        RECT 214.200 66.800 214.600 67.200 ;
        RECT 4.600 65.800 5.000 66.200 ;
        RECT 27.800 65.800 28.200 66.200 ;
        RECT 38.200 65.800 38.600 66.200 ;
        RECT 40.600 65.800 41.000 66.200 ;
        RECT 45.400 65.800 45.800 66.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 195.000 65.800 195.400 66.200 ;
        RECT 116.600 64.800 117.000 65.200 ;
        RECT 120.600 64.800 121.000 65.200 ;
        RECT 55.800 63.800 56.200 64.200 ;
        RECT 79.000 63.800 79.400 64.200 ;
        RECT 88.600 61.800 89.000 62.200 ;
        RECT 59.000 60.800 59.400 61.200 ;
        RECT 91.000 60.800 91.400 61.200 ;
        RECT 238.200 60.800 238.600 61.200 ;
        RECT 68.600 58.800 69.000 59.200 ;
        RECT 230.200 57.800 230.600 58.200 ;
        RECT 137.400 56.800 137.800 57.200 ;
        RECT 46.200 55.800 46.600 56.200 ;
        RECT 74.200 55.800 74.600 56.200 ;
        RECT 91.800 55.800 92.200 56.200 ;
        RECT 231.800 54.800 232.200 55.200 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 107.000 53.800 107.400 54.200 ;
        RECT 151.800 53.800 152.200 54.200 ;
        RECT 242.200 53.800 242.600 54.200 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 73.400 52.800 73.800 53.200 ;
        RECT 119.000 52.800 119.400 53.200 ;
        RECT 200.600 52.800 201.000 53.200 ;
        RECT 243.000 51.800 243.400 52.200 ;
        RECT 183.800 50.800 184.200 51.200 ;
        RECT 184.600 48.800 185.000 49.200 ;
        RECT 30.200 46.800 30.600 47.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 111.000 45.800 111.400 46.200 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 187.800 45.800 188.200 46.200 ;
        RECT 234.200 45.800 234.600 46.200 ;
        RECT 40.600 44.800 41.000 45.200 ;
        RECT 85.400 44.800 85.800 45.200 ;
        RECT 103.000 43.800 103.400 44.200 ;
        RECT 185.400 43.800 185.800 44.200 ;
        RECT 118.200 42.800 118.600 43.200 ;
        RECT 167.000 42.800 167.400 43.200 ;
        RECT 189.400 42.800 189.800 43.200 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 88.600 40.800 89.000 41.200 ;
        RECT 88.600 37.800 89.000 38.200 ;
        RECT 191.800 37.800 192.200 38.200 ;
        RECT 50.200 35.800 50.600 36.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 164.600 35.800 165.000 36.200 ;
        RECT 223.000 35.800 223.400 36.200 ;
        RECT 239.800 35.800 240.200 36.200 ;
        RECT 15.000 34.800 15.400 35.200 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 52.600 34.800 53.000 35.200 ;
        RECT 60.600 34.800 61.000 35.200 ;
        RECT 107.800 33.800 108.200 34.200 ;
        RECT 131.800 33.800 132.200 34.200 ;
        RECT 219.800 33.800 220.200 34.200 ;
        RECT 208.600 32.800 209.000 33.200 ;
        RECT 10.200 29.800 10.600 30.200 ;
        RECT 141.400 29.800 141.800 30.200 ;
        RECT 186.200 29.800 186.600 30.200 ;
        RECT 11.800 27.800 12.200 28.200 ;
        RECT 100.600 27.800 101.000 28.200 ;
        RECT 128.600 26.800 129.000 27.200 ;
        RECT 80.600 25.800 81.000 26.200 ;
        RECT 143.000 23.800 143.400 24.200 ;
        RECT 87.800 21.800 88.200 22.200 ;
        RECT 129.400 21.800 129.800 22.200 ;
        RECT 71.000 20.800 71.400 21.200 ;
        RECT 112.600 18.800 113.000 19.200 ;
        RECT 143.800 18.800 144.200 19.200 ;
        RECT 215.000 17.800 215.400 18.200 ;
        RECT 97.400 16.800 97.800 17.200 ;
        RECT 103.800 15.800 104.200 16.200 ;
        RECT 110.200 15.800 110.600 16.200 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 101.400 14.800 101.800 15.200 ;
        RECT 131.800 14.800 132.200 15.200 ;
        RECT 215.800 14.800 216.200 15.200 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 113.400 13.800 113.800 14.200 ;
        RECT 137.400 9.800 137.800 10.200 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 35.800 7.800 36.200 8.200 ;
        RECT 196.600 6.800 197.000 7.200 ;
        RECT 247.000 6.800 247.400 7.200 ;
        RECT 17.400 5.800 17.800 6.200 ;
        RECT 68.600 5.800 69.000 6.200 ;
        RECT 108.600 5.800 109.000 6.200 ;
        RECT 140.600 5.800 141.000 6.200 ;
      LAYER metal4 ;
        RECT 238.200 235.800 238.600 236.200 ;
        RECT 19.000 234.800 19.400 235.200 ;
        RECT 156.600 234.800 157.000 235.200 ;
        RECT 183.000 234.800 183.400 235.200 ;
        RECT 231.000 234.800 231.400 235.200 ;
        RECT 235.800 235.100 236.200 235.200 ;
        RECT 236.600 235.100 237.000 235.200 ;
        RECT 235.800 234.800 237.000 235.100 ;
        RECT 4.600 234.100 5.000 234.200 ;
        RECT 5.400 234.100 5.800 234.200 ;
        RECT 4.600 233.800 5.800 234.100 ;
        RECT 8.600 223.800 9.000 224.200 ;
        RECT 8.600 207.200 8.900 223.800 ;
        RECT 11.000 214.800 11.400 215.200 ;
        RECT 8.600 206.800 9.000 207.200 ;
        RECT 10.200 156.100 10.600 156.200 ;
        RECT 11.000 156.100 11.300 214.800 ;
        RECT 10.200 155.800 11.300 156.100 ;
        RECT 13.400 204.800 13.800 205.200 ;
        RECT 4.600 124.800 5.000 125.200 ;
        RECT 2.200 84.800 2.600 85.200 ;
        RECT 2.200 56.200 2.500 84.800 ;
        RECT 4.600 66.200 4.900 124.800 ;
        RECT 5.400 67.800 5.800 68.200 ;
        RECT 4.600 65.800 5.000 66.200 ;
        RECT 4.600 65.200 4.900 65.800 ;
        RECT 4.600 64.800 5.000 65.200 ;
        RECT 2.200 55.800 2.600 56.200 ;
        RECT 5.400 54.200 5.700 67.800 ;
        RECT 5.400 53.800 5.800 54.200 ;
        RECT 10.200 30.200 10.500 155.800 ;
        RECT 12.600 138.800 13.000 139.200 ;
        RECT 12.600 106.200 12.900 138.800 ;
        RECT 13.400 122.200 13.700 204.800 ;
        RECT 19.000 176.200 19.300 234.800 ;
        RECT 119.000 233.800 119.400 234.200 ;
        RECT 122.200 233.800 122.600 234.200 ;
        RECT 34.200 232.800 34.600 233.200 ;
        RECT 34.200 217.200 34.500 232.800 ;
        RECT 97.400 231.800 97.800 232.200 ;
        RECT 76.600 231.100 77.000 231.200 ;
        RECT 75.800 230.800 77.000 231.100 ;
        RECT 39.000 226.100 39.400 226.200 ;
        RECT 39.800 226.100 40.200 226.200 ;
        RECT 39.000 225.800 40.200 226.100 ;
        RECT 59.000 226.100 59.400 226.200 ;
        RECT 59.800 226.100 60.200 226.200 ;
        RECT 59.000 225.800 60.200 226.100 ;
        RECT 43.800 224.800 44.200 225.200 ;
        RECT 34.200 216.800 34.600 217.200 ;
        RECT 23.000 198.800 23.400 199.200 ;
        RECT 21.400 190.800 21.800 191.200 ;
        RECT 16.600 175.800 17.000 176.200 ;
        RECT 19.000 175.800 19.400 176.200 ;
        RECT 14.200 174.800 14.600 175.200 ;
        RECT 14.200 146.200 14.500 174.800 ;
        RECT 14.200 145.800 14.600 146.200 ;
        RECT 13.400 121.800 13.800 122.200 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 11.800 75.100 12.200 75.200 ;
        RECT 12.600 75.100 13.000 75.200 ;
        RECT 11.800 74.800 13.000 75.100 ;
        RECT 11.800 47.800 12.200 48.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 10.200 29.800 10.600 30.200 ;
        RECT 10.200 17.200 10.500 29.800 ;
        RECT 10.200 16.800 10.600 17.200 ;
        RECT 11.000 15.200 11.300 34.800 ;
        RECT 11.800 28.200 12.100 47.800 ;
        RECT 14.200 46.200 14.500 145.800 ;
        RECT 16.600 136.200 16.900 175.800 ;
        RECT 19.000 167.200 19.300 175.800 ;
        RECT 20.600 172.800 21.000 173.200 ;
        RECT 19.000 166.800 19.400 167.200 ;
        RECT 19.000 166.200 19.300 166.800 ;
        RECT 17.400 165.800 17.800 166.200 ;
        RECT 19.000 165.800 19.400 166.200 ;
        RECT 17.400 165.100 17.700 165.800 ;
        RECT 17.400 164.800 18.500 165.100 ;
        RECT 18.200 164.200 18.500 164.800 ;
        RECT 18.200 163.800 18.600 164.200 ;
        RECT 16.600 135.800 17.000 136.200 ;
        RECT 16.600 126.200 16.900 135.800 ;
        RECT 16.600 125.800 17.000 126.200 ;
        RECT 15.800 77.800 16.200 78.200 ;
        RECT 15.800 75.200 16.100 77.800 ;
        RECT 15.800 74.800 16.200 75.200 ;
        RECT 16.600 59.200 16.900 125.800 ;
        RECT 16.600 58.800 17.000 59.200 ;
        RECT 15.000 50.800 15.400 51.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 15.000 35.200 15.300 50.800 ;
        RECT 15.000 34.800 15.400 35.200 ;
        RECT 11.800 27.800 12.200 28.200 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 11.800 7.200 12.100 27.800 ;
        RECT 17.400 20.800 17.800 21.200 ;
        RECT 15.000 15.800 15.400 16.200 ;
        RECT 15.000 14.200 15.300 15.800 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 17.400 6.200 17.700 20.800 ;
        RECT 19.000 15.200 19.300 165.800 ;
        RECT 20.600 154.200 20.900 172.800 ;
        RECT 20.600 153.800 21.000 154.200 ;
        RECT 21.400 143.200 21.700 190.800 ;
        RECT 21.400 142.800 21.800 143.200 ;
        RECT 21.400 69.200 21.700 142.800 ;
        RECT 23.000 104.200 23.300 198.800 ;
        RECT 41.400 194.800 41.800 195.200 ;
        RECT 35.000 185.800 35.400 186.200 ;
        RECT 31.800 177.100 32.200 177.200 ;
        RECT 31.000 176.800 32.200 177.100 ;
        RECT 27.800 157.800 28.200 158.200 ;
        RECT 27.800 109.200 28.100 157.800 ;
        RECT 29.400 155.800 29.800 156.200 ;
        RECT 27.800 108.800 28.200 109.200 ;
        RECT 23.000 103.800 23.400 104.200 ;
        RECT 21.400 68.800 21.800 69.200 ;
        RECT 29.400 67.200 29.700 155.800 ;
        RECT 31.000 76.200 31.300 176.800 ;
        RECT 35.000 166.200 35.300 185.800 ;
        RECT 38.200 183.800 38.600 184.200 ;
        RECT 35.000 165.800 35.400 166.200 ;
        RECT 35.000 125.200 35.300 165.800 ;
        RECT 38.200 155.200 38.500 183.800 ;
        RECT 39.800 159.800 40.200 160.200 ;
        RECT 38.200 154.800 38.600 155.200 ;
        RECT 37.400 145.800 37.800 146.200 ;
        RECT 37.400 145.200 37.700 145.800 ;
        RECT 37.400 144.800 37.800 145.200 ;
        RECT 38.200 126.200 38.500 154.800 ;
        RECT 38.200 125.800 38.600 126.200 ;
        RECT 35.000 124.800 35.400 125.200 ;
        RECT 34.200 96.800 34.600 97.200 ;
        RECT 33.400 85.800 33.800 86.200 ;
        RECT 33.400 84.200 33.700 85.800 ;
        RECT 34.200 85.200 34.500 96.800 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 33.400 83.800 33.800 84.200 ;
        RECT 31.000 75.800 31.400 76.200 ;
        RECT 32.600 76.100 33.000 76.200 ;
        RECT 33.400 76.100 33.800 76.200 ;
        RECT 32.600 75.800 33.800 76.100 ;
        RECT 31.000 74.100 31.400 74.200 ;
        RECT 31.800 74.100 32.200 74.200 ;
        RECT 31.000 73.800 32.200 74.100 ;
        RECT 35.000 69.200 35.300 124.800 ;
        RECT 35.800 123.800 36.200 124.200 ;
        RECT 35.000 68.800 35.400 69.200 ;
        RECT 29.400 66.800 29.800 67.200 ;
        RECT 33.400 67.100 33.800 67.200 ;
        RECT 34.200 67.100 34.600 67.200 ;
        RECT 33.400 66.800 34.600 67.100 ;
        RECT 27.800 66.100 28.200 66.200 ;
        RECT 28.600 66.100 29.000 66.200 ;
        RECT 27.800 65.800 29.000 66.100 ;
        RECT 29.400 47.100 29.700 66.800 ;
        RECT 35.000 66.200 35.300 68.800 ;
        RECT 35.000 65.800 35.400 66.200 ;
        RECT 30.200 47.100 30.600 47.200 ;
        RECT 29.400 46.800 30.600 47.100 ;
        RECT 32.600 32.100 33.000 32.200 ;
        RECT 32.600 31.800 33.700 32.100 ;
        RECT 19.000 15.100 19.400 15.200 ;
        RECT 19.000 14.800 20.100 15.100 ;
        RECT 19.800 6.200 20.100 14.800 ;
        RECT 33.400 9.200 33.700 31.800 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 35.800 8.200 36.100 123.800 ;
        RECT 38.200 83.200 38.500 125.800 ;
        RECT 39.800 111.200 40.100 159.800 ;
        RECT 40.600 135.100 41.000 135.200 ;
        RECT 41.400 135.100 41.700 194.800 ;
        RECT 40.600 134.800 41.700 135.100 ;
        RECT 42.200 164.800 42.600 165.200 ;
        RECT 39.800 110.800 40.200 111.200 ;
        RECT 39.000 101.800 39.400 102.200 ;
        RECT 38.200 82.800 38.600 83.200 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 37.400 65.800 38.600 66.100 ;
        RECT 39.000 35.200 39.300 101.800 ;
        RECT 42.200 98.200 42.500 164.800 ;
        RECT 43.000 157.800 43.400 158.200 ;
        RECT 43.000 146.200 43.300 157.800 ;
        RECT 43.000 145.800 43.400 146.200 ;
        RECT 42.200 97.800 42.600 98.200 ;
        RECT 40.600 67.100 41.000 67.200 ;
        RECT 41.400 67.100 41.800 67.200 ;
        RECT 40.600 66.800 41.800 67.100 ;
        RECT 40.600 65.800 41.000 66.200 ;
        RECT 40.600 45.200 40.900 65.800 ;
        RECT 43.000 58.200 43.300 145.800 ;
        RECT 43.800 113.200 44.100 224.800 ;
        RECT 75.800 224.200 76.100 230.800 ;
        RECT 97.400 230.200 97.700 231.800 ;
        RECT 97.400 229.800 97.800 230.200 ;
        RECT 91.000 228.100 91.400 228.200 ;
        RECT 90.200 227.800 91.400 228.100 ;
        RECT 75.800 223.800 76.200 224.200 ;
        RECT 90.200 223.200 90.500 227.800 ;
        RECT 110.200 225.100 110.600 225.200 ;
        RECT 110.200 224.800 111.300 225.100 ;
        RECT 105.400 223.800 105.800 224.200 ;
        RECT 90.200 222.800 90.600 223.200 ;
        RECT 57.400 221.800 57.800 222.200 ;
        RECT 50.200 201.800 50.600 202.200 ;
        RECT 47.000 185.800 47.400 186.200 ;
        RECT 46.200 174.800 46.600 175.200 ;
        RECT 46.200 135.200 46.500 174.800 ;
        RECT 45.400 134.800 45.800 135.200 ;
        RECT 46.200 134.800 46.600 135.200 ;
        RECT 43.800 112.800 44.200 113.200 ;
        RECT 44.600 72.800 45.000 73.200 ;
        RECT 43.000 57.800 43.400 58.200 ;
        RECT 44.600 57.200 44.900 72.800 ;
        RECT 45.400 71.200 45.700 134.800 ;
        RECT 46.200 72.200 46.500 134.800 ;
        RECT 47.000 130.200 47.300 185.800 ;
        RECT 50.200 181.200 50.500 201.800 ;
        RECT 51.800 194.800 52.200 195.200 ;
        RECT 51.800 194.200 52.100 194.800 ;
        RECT 51.800 193.800 52.200 194.200 ;
        RECT 57.400 186.200 57.700 221.800 ;
        RECT 69.400 219.800 69.800 220.200 ;
        RECT 59.800 212.800 60.200 213.200 ;
        RECT 59.000 201.800 59.400 202.200 ;
        RECT 57.400 186.100 57.800 186.200 ;
        RECT 58.200 186.100 58.600 186.200 ;
        RECT 57.400 185.800 58.600 186.100 ;
        RECT 50.200 180.800 50.600 181.200 ;
        RECT 51.000 178.800 51.400 179.200 ;
        RECT 51.000 171.200 51.300 178.800 ;
        RECT 51.000 170.800 51.400 171.200 ;
        RECT 58.200 161.800 58.600 162.200 ;
        RECT 47.800 145.800 48.200 146.200 ;
        RECT 47.800 145.200 48.100 145.800 ;
        RECT 47.800 144.800 48.200 145.200 ;
        RECT 58.200 134.200 58.500 161.800 ;
        RECT 58.200 133.800 58.600 134.200 ;
        RECT 47.000 129.800 47.400 130.200 ;
        RECT 51.000 80.800 51.400 81.200 ;
        RECT 46.200 71.800 46.600 72.200 ;
        RECT 50.200 71.800 50.600 72.200 ;
        RECT 45.400 70.800 45.800 71.200 ;
        RECT 48.600 67.100 49.000 67.200 ;
        RECT 49.400 67.100 49.800 67.200 ;
        RECT 48.600 66.800 49.800 67.100 ;
        RECT 45.400 66.100 45.800 66.200 ;
        RECT 46.200 66.100 46.600 66.200 ;
        RECT 45.400 65.800 46.600 66.100 ;
        RECT 44.600 56.800 45.000 57.200 ;
        RECT 45.400 56.100 45.800 56.200 ;
        RECT 46.200 56.100 46.600 56.200 ;
        RECT 45.400 55.800 46.600 56.100 ;
        RECT 46.200 54.800 46.600 55.200 ;
        RECT 46.200 53.200 46.500 54.800 ;
        RECT 46.200 52.800 46.600 53.200 ;
        RECT 40.600 44.800 41.000 45.200 ;
        RECT 50.200 36.200 50.500 71.800 ;
        RECT 43.000 35.800 43.400 36.200 ;
        RECT 50.200 35.800 50.600 36.200 ;
        RECT 39.000 34.800 39.400 35.200 ;
        RECT 43.000 19.200 43.300 35.800 ;
        RECT 51.000 35.200 51.300 80.800 ;
        RECT 52.600 78.800 53.000 79.200 ;
        RECT 52.600 35.200 52.900 78.800 ;
        RECT 58.200 68.200 58.500 133.800 ;
        RECT 59.000 103.200 59.300 201.800 ;
        RECT 59.800 172.200 60.100 212.800 ;
        RECT 64.600 195.800 65.000 196.200 ;
        RECT 60.600 194.800 61.000 195.200 ;
        RECT 63.000 195.100 63.400 195.200 ;
        RECT 63.800 195.100 64.200 195.200 ;
        RECT 63.000 194.800 64.200 195.100 ;
        RECT 60.600 177.200 60.900 194.800 ;
        RECT 63.800 192.800 64.200 193.200 ;
        RECT 60.600 176.800 61.000 177.200 ;
        RECT 59.800 171.800 60.200 172.200 ;
        RECT 59.800 138.200 60.100 171.800 ;
        RECT 59.800 137.800 60.200 138.200 ;
        RECT 59.000 102.800 59.400 103.200 ;
        RECT 59.800 81.200 60.100 137.800 ;
        RECT 60.600 115.200 60.900 176.800 ;
        RECT 63.800 174.200 64.100 192.800 ;
        RECT 63.800 173.800 64.200 174.200 ;
        RECT 64.600 160.200 64.900 195.800 ;
        RECT 68.600 194.800 69.000 195.200 ;
        RECT 65.400 193.800 65.800 194.200 ;
        RECT 64.600 159.800 65.000 160.200 ;
        RECT 65.400 140.200 65.700 193.800 ;
        RECT 66.200 184.800 66.600 185.200 ;
        RECT 66.200 180.200 66.500 184.800 ;
        RECT 66.200 179.800 66.600 180.200 ;
        RECT 65.400 139.800 65.800 140.200 ;
        RECT 64.600 135.800 65.000 136.200 ;
        RECT 64.600 125.200 64.900 135.800 ;
        RECT 64.600 124.800 65.000 125.200 ;
        RECT 63.800 118.800 64.200 119.200 ;
        RECT 60.600 114.800 61.000 115.200 ;
        RECT 59.800 80.800 60.200 81.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 53.400 67.800 53.800 68.200 ;
        RECT 58.200 67.800 58.600 68.200 ;
        RECT 53.400 67.200 53.700 67.800 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 58.200 65.800 58.600 66.200 ;
        RECT 55.800 64.100 56.200 64.200 ;
        RECT 56.600 64.100 57.000 64.200 ;
        RECT 55.800 63.800 57.000 64.100 ;
        RECT 58.200 45.200 58.500 65.800 ;
        RECT 59.800 64.100 60.200 64.200 ;
        RECT 60.600 64.100 61.000 64.200 ;
        RECT 59.800 63.800 61.000 64.100 ;
        RECT 59.000 60.800 59.400 61.200 ;
        RECT 59.000 58.200 59.300 60.800 ;
        RECT 59.000 57.800 59.400 58.200 ;
        RECT 61.400 57.800 61.800 58.200 ;
        RECT 61.400 54.200 61.700 57.800 ;
        RECT 63.000 54.200 63.300 68.800 ;
        RECT 63.800 61.200 64.100 118.800 ;
        RECT 66.200 115.100 66.500 179.800 ;
        RECT 67.800 149.100 68.200 149.200 ;
        RECT 67.000 148.800 68.200 149.100 ;
        RECT 67.000 122.200 67.300 148.800 ;
        RECT 68.600 130.200 68.900 194.800 ;
        RECT 69.400 166.200 69.700 219.800 ;
        RECT 100.600 216.800 101.000 217.200 ;
        RECT 94.200 215.800 94.600 216.200 ;
        RECT 74.200 213.100 74.600 213.200 ;
        RECT 74.200 212.800 75.300 213.100 ;
        RECT 73.400 208.800 73.800 209.200 ;
        RECT 70.200 194.800 70.600 195.200 ;
        RECT 70.200 194.200 70.500 194.800 ;
        RECT 70.200 193.800 70.600 194.200 ;
        RECT 71.800 185.800 72.200 186.200 ;
        RECT 69.400 165.800 69.800 166.200 ;
        RECT 71.800 138.200 72.100 185.800 ;
        RECT 73.400 149.200 73.700 208.800 ;
        RECT 75.000 199.200 75.300 212.800 ;
        RECT 94.200 211.200 94.500 215.800 ;
        RECT 100.600 215.200 100.900 216.800 ;
        RECT 100.600 214.800 101.000 215.200 ;
        RECT 96.600 211.800 97.000 212.200 ;
        RECT 94.200 210.800 94.600 211.200 ;
        RECT 85.400 201.800 85.800 202.200 ;
        RECT 75.000 198.800 75.400 199.200 ;
        RECT 82.200 195.800 82.600 196.200 ;
        RECT 79.800 194.800 80.200 195.200 ;
        RECT 74.200 186.800 74.600 187.200 ;
        RECT 74.200 151.200 74.500 186.800 ;
        RECT 79.000 173.800 79.400 174.200 ;
        RECT 79.000 172.200 79.300 173.800 ;
        RECT 79.000 171.800 79.400 172.200 ;
        RECT 74.200 150.800 74.600 151.200 ;
        RECT 73.400 148.800 73.800 149.200 ;
        RECT 72.600 139.800 73.000 140.200 ;
        RECT 71.800 137.800 72.200 138.200 ;
        RECT 68.600 129.800 69.000 130.200 ;
        RECT 72.600 125.200 72.900 139.800 ;
        RECT 72.600 124.800 73.000 125.200 ;
        RECT 67.000 121.800 67.400 122.200 ;
        RECT 67.000 121.200 67.300 121.800 ;
        RECT 67.000 120.800 67.400 121.200 ;
        RECT 71.800 119.800 72.200 120.200 ;
        RECT 69.400 118.800 69.800 119.200 ;
        RECT 67.000 115.100 67.400 115.200 ;
        RECT 66.200 114.800 67.400 115.100 ;
        RECT 64.600 90.800 65.000 91.200 ;
        RECT 64.600 87.200 64.900 90.800 ;
        RECT 64.600 86.800 65.000 87.200 ;
        RECT 64.600 86.200 64.900 86.800 ;
        RECT 64.600 85.800 65.000 86.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 65.400 67.100 65.800 67.200 ;
        RECT 64.600 66.800 65.800 67.100 ;
        RECT 63.800 60.800 64.200 61.200 ;
        RECT 61.400 53.800 61.800 54.200 ;
        RECT 63.000 53.800 63.400 54.200 ;
        RECT 58.200 44.800 58.600 45.200 ;
        RECT 60.600 43.800 61.000 44.200 ;
        RECT 60.600 35.200 60.900 43.800 ;
        RECT 67.000 36.200 67.300 114.800 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 67.800 105.800 69.000 106.100 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 67.800 94.200 68.100 94.800 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 69.400 84.200 69.700 118.800 ;
        RECT 71.000 110.800 71.400 111.200 ;
        RECT 69.400 83.800 69.800 84.200 ;
        RECT 70.200 82.800 70.600 83.200 ;
        RECT 68.600 68.800 69.000 69.200 ;
        RECT 68.600 59.200 68.900 68.800 ;
        RECT 68.600 58.800 69.000 59.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 69.400 35.800 69.800 36.200 ;
        RECT 69.400 35.200 69.700 35.800 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 52.600 34.800 53.000 35.200 ;
        RECT 60.600 34.800 61.000 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 70.200 28.200 70.500 82.800 ;
        RECT 70.200 27.800 70.600 28.200 ;
        RECT 59.800 24.800 60.200 25.200 ;
        RECT 59.800 24.200 60.100 24.800 ;
        RECT 59.800 23.800 60.200 24.200 ;
        RECT 71.000 21.200 71.300 110.800 ;
        RECT 71.800 83.200 72.100 119.800 ;
        RECT 72.600 104.800 73.000 105.200 ;
        RECT 71.800 82.800 72.200 83.200 ;
        RECT 72.600 80.200 72.900 104.800 ;
        RECT 72.600 79.800 73.000 80.200 ;
        RECT 73.400 53.200 73.700 148.800 ;
        RECT 74.200 122.200 74.500 150.800 ;
        RECT 79.800 135.200 80.100 194.800 ;
        RECT 81.400 156.800 81.800 157.200 ;
        RECT 79.800 134.800 80.200 135.200 ;
        RECT 74.200 121.800 74.600 122.200 ;
        RECT 79.800 120.100 80.200 120.200 ;
        RECT 79.800 119.800 80.900 120.100 ;
        RECT 78.200 115.100 78.600 115.200 ;
        RECT 79.000 115.100 79.400 115.200 ;
        RECT 78.200 114.800 79.400 115.100 ;
        RECT 79.000 109.800 79.400 110.200 ;
        RECT 75.000 72.800 75.400 73.200 ;
        RECT 75.000 66.200 75.300 72.800 ;
        RECT 75.800 70.800 76.200 71.200 ;
        RECT 75.800 67.200 76.100 70.800 ;
        RECT 75.800 66.800 76.200 67.200 ;
        RECT 79.000 66.200 79.300 109.800 ;
        RECT 80.600 99.200 80.900 119.800 ;
        RECT 81.400 115.200 81.700 156.800 ;
        RECT 82.200 131.200 82.500 195.800 ;
        RECT 85.400 182.200 85.700 201.800 ;
        RECT 95.000 195.800 95.400 196.200 ;
        RECT 95.000 195.200 95.300 195.800 ;
        RECT 95.000 194.800 95.400 195.200 ;
        RECT 95.000 192.800 95.400 193.200 ;
        RECT 85.400 181.800 85.800 182.200 ;
        RECT 87.000 181.800 87.400 182.200 ;
        RECT 84.600 165.100 85.000 165.200 ;
        RECT 83.800 164.800 85.000 165.100 ;
        RECT 83.800 132.200 84.100 164.800 ;
        RECT 85.400 154.200 85.700 181.800 ;
        RECT 86.200 174.800 86.600 175.200 ;
        RECT 85.400 153.800 85.800 154.200 ;
        RECT 86.200 137.200 86.500 174.800 ;
        RECT 86.200 136.800 86.600 137.200 ;
        RECT 85.400 134.800 85.800 135.200 ;
        RECT 83.800 131.800 84.200 132.200 ;
        RECT 82.200 130.800 82.600 131.200 ;
        RECT 82.200 129.800 82.600 130.200 ;
        RECT 82.200 126.200 82.500 129.800 ;
        RECT 82.200 125.800 82.600 126.200 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 82.200 100.200 82.500 111.800 ;
        RECT 82.200 99.800 82.600 100.200 ;
        RECT 83.800 99.200 84.100 131.800 ;
        RECT 84.600 106.800 85.000 107.200 ;
        RECT 80.600 98.800 81.000 99.200 ;
        RECT 83.800 98.800 84.200 99.200 ;
        RECT 80.600 91.800 81.000 92.200 ;
        RECT 79.800 79.800 80.200 80.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 75.800 65.800 77.000 66.100 ;
        RECT 79.000 65.800 79.400 66.200 ;
        RECT 74.200 56.200 74.500 65.800 ;
        RECT 79.000 64.200 79.300 65.800 ;
        RECT 79.000 63.800 79.400 64.200 ;
        RECT 74.200 55.800 74.600 56.200 ;
        RECT 73.400 52.800 73.800 53.200 ;
        RECT 79.800 29.200 80.100 79.800 ;
        RECT 79.800 28.800 80.200 29.200 ;
        RECT 80.600 26.200 80.900 91.800 ;
        RECT 83.000 68.100 83.400 68.200 ;
        RECT 83.800 68.100 84.200 68.200 ;
        RECT 83.000 67.800 84.200 68.100 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 82.200 66.100 82.600 66.200 ;
        RECT 81.400 65.800 82.600 66.100 ;
        RECT 84.600 46.200 84.900 106.800 ;
        RECT 85.400 95.200 85.700 134.800 ;
        RECT 86.200 124.800 86.600 125.200 ;
        RECT 86.200 106.200 86.500 124.800 ;
        RECT 87.000 116.200 87.300 181.800 ;
        RECT 94.200 166.800 94.600 167.200 ;
        RECT 87.800 163.800 88.200 164.200 ;
        RECT 87.800 144.200 88.100 163.800 ;
        RECT 87.800 143.800 88.200 144.200 ;
        RECT 88.600 140.800 89.000 141.200 ;
        RECT 87.800 121.800 88.200 122.200 ;
        RECT 87.000 115.800 87.400 116.200 ;
        RECT 86.200 105.800 86.600 106.200 ;
        RECT 85.400 94.800 85.800 95.200 ;
        RECT 87.000 90.200 87.300 115.800 ;
        RECT 87.000 89.800 87.400 90.200 ;
        RECT 87.800 87.200 88.100 121.800 ;
        RECT 87.800 86.800 88.200 87.200 ;
        RECT 88.600 62.200 88.900 140.800 ;
        RECT 89.400 135.800 89.800 136.200 ;
        RECT 89.400 103.200 89.700 135.800 ;
        RECT 94.200 126.200 94.500 166.800 ;
        RECT 92.600 125.800 93.000 126.200 ;
        RECT 94.200 125.800 94.600 126.200 ;
        RECT 92.600 105.200 92.900 125.800 ;
        RECT 95.000 116.200 95.300 192.800 ;
        RECT 96.600 175.200 96.900 211.800 ;
        RECT 97.400 205.800 97.800 206.200 ;
        RECT 97.400 199.200 97.700 205.800 ;
        RECT 97.400 198.800 97.800 199.200 ;
        RECT 96.600 174.800 97.000 175.200 ;
        RECT 95.800 164.800 96.200 165.200 ;
        RECT 95.000 115.800 95.400 116.200 ;
        RECT 94.200 107.800 94.600 108.200 ;
        RECT 92.600 104.800 93.000 105.200 ;
        RECT 89.400 102.800 89.800 103.200 ;
        RECT 92.600 86.200 92.900 104.800 ;
        RECT 93.400 91.800 93.800 92.200 ;
        RECT 91.000 86.100 91.400 86.200 ;
        RECT 91.800 86.100 92.200 86.200 ;
        RECT 91.000 85.800 92.200 86.100 ;
        RECT 92.600 85.800 93.000 86.200 ;
        RECT 91.000 81.800 91.400 82.200 ;
        RECT 88.600 61.800 89.000 62.200 ;
        RECT 86.200 54.800 86.600 55.200 ;
        RECT 87.800 54.800 88.200 55.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 84.600 45.100 84.900 45.800 ;
        RECT 85.400 45.100 85.800 45.200 ;
        RECT 84.600 44.800 85.800 45.100 ;
        RECT 86.200 40.200 86.500 54.800 ;
        RECT 86.200 39.800 86.600 40.200 ;
        RECT 80.600 25.800 81.000 26.200 ;
        RECT 87.800 22.200 88.100 54.800 ;
        RECT 88.600 41.200 88.900 61.800 ;
        RECT 91.000 61.200 91.300 81.800 ;
        RECT 93.400 67.100 93.700 91.800 ;
        RECT 94.200 70.200 94.500 107.800 ;
        RECT 95.800 100.200 96.100 164.800 ;
        RECT 97.400 144.200 97.700 198.800 ;
        RECT 97.400 143.800 97.800 144.200 ;
        RECT 100.600 136.200 100.900 214.800 ;
        RECT 105.400 206.200 105.700 223.800 ;
        RECT 106.200 219.800 106.600 220.200 ;
        RECT 105.400 205.800 105.800 206.200 ;
        RECT 102.200 203.800 102.600 204.200 ;
        RECT 101.400 174.800 101.800 175.200 ;
        RECT 101.400 143.200 101.700 174.800 ;
        RECT 102.200 174.200 102.500 203.800 ;
        RECT 105.400 180.800 105.800 181.200 ;
        RECT 102.200 173.800 102.600 174.200 ;
        RECT 103.800 169.800 104.200 170.200 ;
        RECT 101.400 142.800 101.800 143.200 ;
        RECT 101.400 137.800 101.800 138.200 ;
        RECT 100.600 135.800 101.000 136.200 ;
        RECT 97.400 131.800 97.800 132.200 ;
        RECT 97.400 127.200 97.700 131.800 ;
        RECT 97.400 126.800 97.800 127.200 ;
        RECT 101.400 127.100 101.700 137.800 ;
        RECT 102.200 127.100 102.600 127.200 ;
        RECT 101.400 126.800 102.600 127.100 ;
        RECT 100.600 122.800 101.000 123.200 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 96.600 114.200 96.900 114.800 ;
        RECT 96.600 113.800 97.000 114.200 ;
        RECT 95.800 99.800 96.200 100.200 ;
        RECT 96.600 99.800 97.000 100.200 ;
        RECT 96.600 97.200 96.900 99.800 ;
        RECT 96.600 96.800 97.000 97.200 ;
        RECT 95.800 86.800 96.200 87.200 ;
        RECT 94.200 69.800 94.600 70.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 93.400 66.800 94.600 67.100 ;
        RECT 91.000 60.800 91.400 61.200 ;
        RECT 91.800 60.800 92.200 61.200 ;
        RECT 91.000 47.200 91.300 60.800 ;
        RECT 91.800 56.200 92.100 60.800 ;
        RECT 91.800 55.800 92.200 56.200 ;
        RECT 91.000 46.800 91.400 47.200 ;
        RECT 88.600 40.800 89.000 41.200 ;
        RECT 95.800 39.200 96.100 86.800 ;
        RECT 100.600 73.200 100.900 122.800 ;
        RECT 103.800 113.200 104.100 169.800 ;
        RECT 105.400 154.200 105.700 180.800 ;
        RECT 105.400 153.800 105.800 154.200 ;
        RECT 104.600 114.800 105.000 115.200 ;
        RECT 103.800 112.800 104.200 113.200 ;
        RECT 101.400 93.800 101.800 94.200 ;
        RECT 103.000 93.800 103.400 94.200 ;
        RECT 100.600 72.800 101.000 73.200 ;
        RECT 97.400 70.800 97.800 71.200 ;
        RECT 100.600 70.800 101.000 71.200 ;
        RECT 97.400 52.200 97.700 70.800 ;
        RECT 100.600 68.200 100.900 70.800 ;
        RECT 100.600 67.800 101.000 68.200 ;
        RECT 101.400 60.200 101.700 93.800 ;
        RECT 103.000 88.200 103.300 93.800 ;
        RECT 103.000 87.800 103.400 88.200 ;
        RECT 103.000 75.200 103.300 87.800 ;
        RECT 104.600 85.200 104.900 114.800 ;
        RECT 104.600 84.800 105.000 85.200 ;
        RECT 103.000 74.800 103.400 75.200 ;
        RECT 105.400 74.200 105.700 153.800 ;
        RECT 106.200 117.200 106.500 219.800 ;
        RECT 107.800 211.800 108.200 212.200 ;
        RECT 107.000 183.800 107.400 184.200 ;
        RECT 107.000 119.200 107.300 183.800 ;
        RECT 107.800 166.200 108.100 211.800 ;
        RECT 107.800 165.800 108.200 166.200 ;
        RECT 107.000 118.800 107.400 119.200 ;
        RECT 106.200 116.800 106.600 117.200 ;
        RECT 106.200 101.800 106.600 102.200 ;
        RECT 106.200 92.200 106.500 101.800 ;
        RECT 106.200 91.800 106.600 92.200 ;
        RECT 105.400 73.800 105.800 74.200 ;
        RECT 105.400 70.200 105.700 73.800 ;
        RECT 105.400 69.800 105.800 70.200 ;
        RECT 106.200 68.200 106.500 91.800 ;
        RECT 106.200 67.800 106.600 68.200 ;
        RECT 101.400 59.800 101.800 60.200 ;
        RECT 107.000 54.200 107.300 118.800 ;
        RECT 107.800 112.200 108.100 165.800 ;
        RECT 111.000 139.200 111.300 224.800 ;
        RECT 115.000 223.800 115.400 224.200 ;
        RECT 115.000 222.200 115.300 223.800 ;
        RECT 119.000 222.200 119.300 233.800 ;
        RECT 122.200 227.200 122.500 233.800 ;
        RECT 135.800 229.800 136.200 230.200 ;
        RECT 135.800 227.200 136.100 229.800 ;
        RECT 122.200 226.800 122.600 227.200 ;
        RECT 135.800 226.800 136.200 227.200 ;
        RECT 154.200 227.100 154.600 227.200 ;
        RECT 155.000 227.100 155.400 227.200 ;
        RECT 154.200 226.800 155.400 227.100 ;
        RECT 115.000 222.100 115.400 222.200 ;
        RECT 115.000 221.800 116.100 222.100 ;
        RECT 112.600 206.100 113.000 206.200 ;
        RECT 113.400 206.100 113.800 206.200 ;
        RECT 112.600 205.800 113.800 206.100 ;
        RECT 115.800 203.200 116.100 221.800 ;
        RECT 119.000 221.800 119.400 222.200 ;
        RECT 115.800 202.800 116.200 203.200 ;
        RECT 111.800 202.100 112.200 202.200 ;
        RECT 112.600 202.100 113.000 202.200 ;
        RECT 111.800 201.800 113.000 202.100 ;
        RECT 117.400 186.800 117.800 187.200 ;
        RECT 117.400 183.200 117.700 186.800 ;
        RECT 117.400 182.800 117.800 183.200 ;
        RECT 116.600 163.800 117.000 164.200 ;
        RECT 114.200 155.800 114.600 156.200 ;
        RECT 111.000 138.800 111.400 139.200 ;
        RECT 107.800 111.800 108.200 112.200 ;
        RECT 107.800 109.800 108.200 110.200 ;
        RECT 107.800 75.200 108.100 109.800 ;
        RECT 108.600 105.800 109.000 106.200 ;
        RECT 107.800 74.800 108.200 75.200 ;
        RECT 107.800 63.800 108.200 64.200 ;
        RECT 107.000 53.800 107.400 54.200 ;
        RECT 97.400 51.800 97.800 52.200 ;
        RECT 95.800 38.800 96.200 39.200 ;
        RECT 88.600 37.800 89.000 38.200 ;
        RECT 87.800 21.800 88.200 22.200 ;
        RECT 71.000 20.800 71.400 21.200 ;
        RECT 88.600 19.200 88.900 37.800 ;
        RECT 43.000 18.800 43.400 19.200 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 97.400 17.200 97.700 51.800 ;
        RECT 103.000 43.800 103.400 44.200 ;
        RECT 100.600 30.800 101.000 31.200 ;
        RECT 100.600 28.200 100.900 30.800 ;
        RECT 100.600 27.800 101.000 28.200 ;
        RECT 97.400 16.800 97.800 17.200 ;
        RECT 103.000 16.200 103.300 43.800 ;
        RECT 107.800 34.200 108.100 63.800 ;
        RECT 107.800 33.800 108.200 34.200 ;
        RECT 103.000 16.100 103.400 16.200 ;
        RECT 103.800 16.100 104.200 16.200 ;
        RECT 103.000 15.800 104.200 16.100 ;
        RECT 101.400 14.800 101.800 15.200 ;
        RECT 101.400 10.200 101.700 14.800 ;
        RECT 101.400 9.800 101.800 10.200 ;
        RECT 35.800 7.800 36.200 8.200 ;
        RECT 108.600 6.200 108.900 105.800 ;
        RECT 109.400 105.100 109.800 105.200 ;
        RECT 110.200 105.100 110.600 105.200 ;
        RECT 109.400 104.800 110.600 105.100 ;
        RECT 111.800 95.800 112.200 96.200 ;
        RECT 111.000 88.800 111.400 89.200 ;
        RECT 111.000 76.200 111.300 88.800 ;
        RECT 111.800 85.200 112.100 95.800 ;
        RECT 114.200 95.200 114.500 155.800 ;
        RECT 115.000 126.800 115.400 127.200 ;
        RECT 115.000 118.200 115.300 126.800 ;
        RECT 115.800 119.800 116.200 120.200 ;
        RECT 115.800 118.200 116.100 119.800 ;
        RECT 115.000 117.800 115.400 118.200 ;
        RECT 115.800 117.800 116.200 118.200 ;
        RECT 115.000 116.800 115.400 117.200 ;
        RECT 114.200 94.800 114.600 95.200 ;
        RECT 114.200 91.200 114.500 94.800 ;
        RECT 114.200 90.800 114.600 91.200 ;
        RECT 111.800 84.800 112.200 85.200 ;
        RECT 110.200 76.100 110.600 76.200 ;
        RECT 109.400 75.800 110.600 76.100 ;
        RECT 111.000 75.800 111.400 76.200 ;
        RECT 109.400 16.100 109.700 75.800 ;
        RECT 110.200 65.800 110.600 66.200 ;
        RECT 110.200 65.200 110.500 65.800 ;
        RECT 110.200 64.800 110.600 65.200 ;
        RECT 110.200 56.800 110.600 57.200 ;
        RECT 110.200 28.200 110.500 56.800 ;
        RECT 111.000 46.200 111.300 75.800 ;
        RECT 115.000 69.200 115.300 116.800 ;
        RECT 115.800 90.200 116.100 117.800 ;
        RECT 116.600 91.200 116.900 163.800 ;
        RECT 117.400 159.200 117.700 182.800 ;
        RECT 117.400 158.800 117.800 159.200 ;
        RECT 118.200 112.800 118.600 113.200 ;
        RECT 118.200 110.200 118.500 112.800 ;
        RECT 118.200 109.800 118.600 110.200 ;
        RECT 119.000 106.200 119.300 221.800 ;
        RECT 122.200 154.200 122.500 226.800 ;
        RECT 124.600 225.800 125.000 226.200 ;
        RECT 144.600 225.800 145.000 226.200 ;
        RECT 124.600 225.200 124.900 225.800 ;
        RECT 144.600 225.200 144.900 225.800 ;
        RECT 124.600 224.800 125.000 225.200 ;
        RECT 144.600 224.800 145.000 225.200 ;
        RECT 148.600 223.800 149.000 224.200 ;
        RECT 134.200 222.800 134.600 223.200 ;
        RECT 131.000 214.800 131.400 215.200 ;
        RECT 131.000 213.200 131.300 214.800 ;
        RECT 131.000 212.800 131.400 213.200 ;
        RECT 130.200 202.800 130.600 203.200 ;
        RECT 126.200 196.800 126.600 197.200 ;
        RECT 126.200 175.200 126.500 196.800 ;
        RECT 130.200 194.200 130.500 202.800 ;
        RECT 132.600 195.800 133.000 196.200 ;
        RECT 130.200 193.800 130.600 194.200 ;
        RECT 130.200 189.200 130.500 193.800 ;
        RECT 130.200 188.800 130.600 189.200 ;
        RECT 126.200 174.800 126.600 175.200 ;
        RECT 123.000 173.800 123.400 174.200 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 119.000 105.800 119.400 106.200 ;
        RECT 119.000 103.200 119.300 105.800 ;
        RECT 120.600 104.100 121.000 104.200 ;
        RECT 121.400 104.100 121.800 104.200 ;
        RECT 120.600 103.800 121.800 104.100 ;
        RECT 118.200 102.800 118.600 103.200 ;
        RECT 119.000 102.800 119.400 103.200 ;
        RECT 118.200 99.200 118.500 102.800 ;
        RECT 118.200 98.800 118.600 99.200 ;
        RECT 117.400 95.800 117.800 96.200 ;
        RECT 116.600 90.800 117.000 91.200 ;
        RECT 115.800 89.800 116.200 90.200 ;
        RECT 115.800 73.200 116.100 89.800 ;
        RECT 116.600 78.200 116.900 90.800 ;
        RECT 117.400 84.200 117.700 95.800 ;
        RECT 122.200 89.200 122.500 153.800 ;
        RECT 123.000 151.200 123.300 173.800 ;
        RECT 123.800 171.800 124.200 172.200 ;
        RECT 123.800 165.200 124.100 171.800 ;
        RECT 123.800 164.800 124.200 165.200 ;
        RECT 123.000 150.800 123.400 151.200 ;
        RECT 125.400 145.800 125.800 146.200 ;
        RECT 123.800 135.800 124.200 136.200 ;
        RECT 123.800 106.200 124.100 135.800 ;
        RECT 123.800 105.800 124.200 106.200 ;
        RECT 125.400 100.200 125.700 145.800 ;
        RECT 130.200 145.200 130.500 188.800 ;
        RECT 131.000 184.800 131.400 185.200 ;
        RECT 131.000 173.200 131.300 184.800 ;
        RECT 132.600 184.200 132.900 195.800 ;
        RECT 134.200 186.200 134.500 222.800 ;
        RECT 143.800 213.800 144.200 214.200 ;
        RECT 140.600 198.100 141.000 198.200 ;
        RECT 139.800 197.800 141.000 198.100 ;
        RECT 137.400 193.800 137.800 194.200 ;
        RECT 134.200 185.800 134.600 186.200 ;
        RECT 132.600 183.800 133.000 184.200 ;
        RECT 131.000 172.800 131.400 173.200 ;
        RECT 131.800 172.800 132.200 173.200 ;
        RECT 131.000 162.800 131.400 163.200 ;
        RECT 130.200 144.800 130.600 145.200 ;
        RECT 131.000 137.200 131.300 162.800 ;
        RECT 131.000 136.800 131.400 137.200 ;
        RECT 130.200 132.800 130.600 133.200 ;
        RECT 127.800 124.800 128.200 125.200 ;
        RECT 127.800 112.200 128.100 124.800 ;
        RECT 127.800 111.800 128.200 112.200 ;
        RECT 130.200 101.200 130.500 132.800 ;
        RECT 131.800 106.200 132.100 172.800 ;
        RECT 132.600 160.200 132.900 183.800 ;
        RECT 133.400 174.800 133.800 175.200 ;
        RECT 132.600 159.800 133.000 160.200 ;
        RECT 132.600 158.800 133.000 159.200 ;
        RECT 132.600 106.200 132.900 158.800 ;
        RECT 131.000 105.800 131.400 106.200 ;
        RECT 131.800 105.800 132.200 106.200 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 131.000 105.200 131.300 105.800 ;
        RECT 131.000 104.800 131.400 105.200 ;
        RECT 130.200 100.800 130.600 101.200 ;
        RECT 125.400 99.800 125.800 100.200 ;
        RECT 128.600 92.800 129.000 93.200 ;
        RECT 122.200 88.800 122.600 89.200 ;
        RECT 117.400 83.800 117.800 84.200 ;
        RECT 122.200 78.200 122.500 88.800 ;
        RECT 127.800 87.800 128.200 88.200 ;
        RECT 123.800 85.800 124.200 86.200 ;
        RECT 125.400 85.800 125.800 86.200 ;
        RECT 116.600 77.800 117.000 78.200 ;
        RECT 119.800 77.800 120.200 78.200 ;
        RECT 122.200 77.800 122.600 78.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 116.600 73.200 116.900 74.800 ;
        RECT 115.800 72.800 116.200 73.200 ;
        RECT 116.600 72.800 117.000 73.200 ;
        RECT 116.600 70.800 117.000 71.200 ;
        RECT 115.800 69.800 116.200 70.200 ;
        RECT 115.800 69.200 116.100 69.800 ;
        RECT 115.000 68.800 115.400 69.200 ;
        RECT 115.800 68.800 116.200 69.200 ;
        RECT 114.200 65.800 114.600 66.200 ;
        RECT 114.200 65.200 114.500 65.800 ;
        RECT 114.200 64.800 114.600 65.200 ;
        RECT 114.200 57.800 114.600 58.200 ;
        RECT 114.200 57.200 114.500 57.800 ;
        RECT 114.200 56.800 114.600 57.200 ;
        RECT 111.000 45.800 111.400 46.200 ;
        RECT 115.000 37.200 115.300 68.800 ;
        RECT 116.600 65.200 116.900 70.800 ;
        RECT 116.600 64.800 117.000 65.200 ;
        RECT 119.800 56.200 120.100 77.800 ;
        RECT 123.800 73.200 124.100 85.800 ;
        RECT 125.400 85.200 125.700 85.800 ;
        RECT 125.400 84.800 125.800 85.200 ;
        RECT 123.800 72.800 124.200 73.200 ;
        RECT 127.800 68.200 128.100 87.800 ;
        RECT 127.800 67.800 128.200 68.200 ;
        RECT 120.600 64.800 121.000 65.200 ;
        RECT 119.800 55.800 120.200 56.200 ;
        RECT 119.800 53.200 120.100 55.800 ;
        RECT 119.000 53.100 119.400 53.200 ;
        RECT 118.200 52.800 119.400 53.100 ;
        RECT 119.800 52.800 120.200 53.200 ;
        RECT 118.200 43.200 118.500 52.800 ;
        RECT 118.200 42.800 118.600 43.200 ;
        RECT 120.600 41.200 120.900 64.800 ;
        RECT 120.600 40.800 121.000 41.200 ;
        RECT 115.000 36.800 115.400 37.200 ;
        RECT 114.200 35.800 114.600 36.200 ;
        RECT 114.200 35.200 114.500 35.800 ;
        RECT 114.200 34.800 114.600 35.200 ;
        RECT 110.200 27.800 110.600 28.200 ;
        RECT 128.600 27.200 128.900 92.800 ;
        RECT 129.400 89.800 129.800 90.200 ;
        RECT 129.400 87.200 129.700 89.800 ;
        RECT 129.400 86.800 129.800 87.200 ;
        RECT 130.200 77.200 130.500 100.800 ;
        RECT 130.200 76.800 130.600 77.200 ;
        RECT 131.000 75.200 131.300 104.800 ;
        RECT 131.800 79.200 132.100 105.800 ;
        RECT 132.600 96.200 132.900 105.800 ;
        RECT 133.400 105.200 133.700 174.800 ;
        RECT 134.200 171.200 134.500 185.800 ;
        RECT 134.200 170.800 134.600 171.200 ;
        RECT 135.800 146.800 136.200 147.200 ;
        RECT 135.800 114.200 136.100 146.800 ;
        RECT 137.400 133.200 137.700 193.800 ;
        RECT 139.000 135.800 139.400 136.200 ;
        RECT 137.400 132.800 137.800 133.200 ;
        RECT 135.800 113.800 136.200 114.200 ;
        RECT 133.400 104.800 133.800 105.200 ;
        RECT 134.200 104.100 134.600 104.200 ;
        RECT 135.000 104.100 135.400 104.200 ;
        RECT 134.200 103.800 135.400 104.100 ;
        RECT 132.600 95.800 133.000 96.200 ;
        RECT 135.800 94.200 136.100 113.800 ;
        RECT 138.200 98.800 138.600 99.200 ;
        RECT 135.800 93.800 136.200 94.200 ;
        RECT 133.400 90.800 133.800 91.200 ;
        RECT 133.400 81.200 133.700 90.800 ;
        RECT 133.400 80.800 133.800 81.200 ;
        RECT 131.800 78.800 132.200 79.200 ;
        RECT 131.800 76.800 132.200 77.200 ;
        RECT 131.800 75.200 132.100 76.800 ;
        RECT 131.000 74.800 131.400 75.200 ;
        RECT 131.800 74.800 132.200 75.200 ;
        RECT 130.200 73.100 130.600 73.200 ;
        RECT 129.400 72.800 130.600 73.100 ;
        RECT 128.600 26.800 129.000 27.200 ;
        RECT 129.400 22.200 129.700 72.800 ;
        RECT 135.800 42.200 136.100 93.800 ;
        RECT 137.400 92.800 137.800 93.200 ;
        RECT 136.600 74.800 137.000 75.200 ;
        RECT 136.600 52.200 136.900 74.800 ;
        RECT 137.400 66.200 137.700 92.800 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 137.400 57.200 137.700 65.800 ;
        RECT 137.400 56.800 137.800 57.200 ;
        RECT 136.600 51.800 137.000 52.200 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 131.800 33.800 132.200 34.200 ;
        RECT 131.800 28.200 132.100 33.800 ;
        RECT 131.800 27.800 132.200 28.200 ;
        RECT 129.400 21.800 129.800 22.200 ;
        RECT 112.600 18.800 113.000 19.200 ;
        RECT 110.200 16.100 110.600 16.200 ;
        RECT 109.400 15.800 110.600 16.100 ;
        RECT 112.600 14.100 112.900 18.800 ;
        RECT 131.800 15.200 132.100 27.800 ;
        RECT 138.200 24.200 138.500 98.800 ;
        RECT 139.000 84.200 139.300 135.800 ;
        RECT 139.800 124.200 140.100 197.800 ;
        RECT 143.800 195.200 144.100 213.800 ;
        RECT 145.400 211.800 145.800 212.200 ;
        RECT 145.400 208.200 145.700 211.800 ;
        RECT 145.400 207.800 145.800 208.200 ;
        RECT 144.600 195.800 145.000 196.200 ;
        RECT 143.800 194.800 144.200 195.200 ;
        RECT 140.600 193.800 141.000 194.200 ;
        RECT 143.800 193.800 144.200 194.200 ;
        RECT 140.600 132.200 140.900 193.800 ;
        RECT 143.800 192.200 144.100 193.800 ;
        RECT 144.600 193.200 144.900 195.800 ;
        RECT 144.600 193.100 145.000 193.200 ;
        RECT 145.400 193.100 145.800 193.200 ;
        RECT 144.600 192.800 145.800 193.100 ;
        RECT 143.800 191.800 144.200 192.200 ;
        RECT 148.600 187.200 148.900 223.800 ;
        RECT 148.600 186.800 149.000 187.200 ;
        RECT 149.400 187.100 149.800 187.200 ;
        RECT 150.200 187.100 150.600 187.200 ;
        RECT 149.400 186.800 150.600 187.100 ;
        RECT 154.200 185.800 154.600 186.200 ;
        RECT 154.200 184.200 154.500 185.800 ;
        RECT 154.200 183.800 154.600 184.200 ;
        RECT 147.800 182.800 148.200 183.200 ;
        RECT 147.800 176.200 148.100 182.800 ;
        RECT 155.000 179.800 155.400 180.200 ;
        RECT 150.200 176.800 150.600 177.200 ;
        RECT 150.200 176.200 150.500 176.800 ;
        RECT 147.800 175.800 148.200 176.200 ;
        RECT 150.200 175.800 150.600 176.200 ;
        RECT 155.000 165.200 155.300 179.800 ;
        RECT 155.000 164.800 155.400 165.200 ;
        RECT 155.800 164.800 156.200 165.200 ;
        RECT 143.800 155.800 144.200 156.200 ;
        RECT 147.800 155.800 148.200 156.200 ;
        RECT 140.600 131.800 141.000 132.200 ;
        RECT 139.800 123.800 140.200 124.200 ;
        RECT 139.800 119.200 140.100 123.800 ;
        RECT 139.800 118.800 140.200 119.200 ;
        RECT 139.800 84.200 140.100 118.800 ;
        RECT 143.800 108.200 144.100 155.800 ;
        RECT 147.800 142.200 148.100 155.800 ;
        RECT 147.800 141.800 148.200 142.200 ;
        RECT 151.800 133.800 152.200 134.200 ;
        RECT 143.800 107.800 144.200 108.200 ;
        RECT 141.400 87.800 141.800 88.200 ;
        RECT 139.000 83.800 139.400 84.200 ;
        RECT 139.800 83.800 140.200 84.200 ;
        RECT 139.000 72.200 139.300 83.800 ;
        RECT 139.000 71.800 139.400 72.200 ;
        RECT 141.400 65.200 141.700 87.800 ;
        RECT 149.400 85.100 149.800 85.200 ;
        RECT 150.200 85.100 150.600 85.200 ;
        RECT 149.400 84.800 150.600 85.100 ;
        RECT 151.800 74.200 152.100 133.800 ;
        RECT 155.800 103.200 156.100 164.800 ;
        RECT 156.600 139.200 156.900 234.800 ;
        RECT 181.400 230.800 181.800 231.200 ;
        RECT 169.400 208.800 169.800 209.200 ;
        RECT 169.400 205.200 169.700 208.800 ;
        RECT 169.400 204.800 169.800 205.200 ;
        RECT 165.400 195.800 165.800 196.200 ;
        RECT 158.200 185.100 158.600 185.200 ;
        RECT 159.000 185.100 159.400 185.200 ;
        RECT 158.200 184.800 159.400 185.100 ;
        RECT 159.800 166.800 160.200 167.200 ;
        RECT 159.800 166.200 160.100 166.800 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 160.600 164.800 161.000 165.200 ;
        RECT 156.600 138.800 157.000 139.200 ;
        RECT 155.800 102.800 156.200 103.200 ;
        RECT 156.600 85.200 156.900 138.800 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 157.400 130.200 157.700 134.800 ;
        RECT 157.400 129.800 157.800 130.200 ;
        RECT 160.600 112.200 160.900 164.800 ;
        RECT 163.800 154.800 164.200 155.200 ;
        RECT 161.400 126.800 161.800 127.200 ;
        RECT 160.600 111.800 161.000 112.200 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 156.600 84.800 157.000 85.200 ;
        RECT 151.800 73.800 152.200 74.200 ;
        RECT 143.800 71.800 144.200 72.200 ;
        RECT 141.400 64.800 141.800 65.200 ;
        RECT 143.800 51.200 144.100 71.800 ;
        RECT 151.800 54.200 152.100 73.800 ;
        RECT 151.800 53.800 152.200 54.200 ;
        RECT 143.800 50.800 144.200 51.200 ;
        RECT 157.400 31.200 157.700 94.800 ;
        RECT 159.800 90.800 160.200 91.200 ;
        RECT 159.800 88.200 160.100 90.800 ;
        RECT 159.800 87.800 160.200 88.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 160.600 87.100 161.000 87.200 ;
        RECT 159.800 86.800 161.000 87.100 ;
        RECT 159.800 81.800 160.200 82.200 ;
        RECT 159.800 46.200 160.100 81.800 ;
        RECT 160.600 74.800 161.000 75.200 ;
        RECT 160.600 74.200 160.900 74.800 ;
        RECT 160.600 73.800 161.000 74.200 ;
        RECT 161.400 65.200 161.700 126.800 ;
        RECT 163.800 110.200 164.100 154.800 ;
        RECT 163.800 109.800 164.200 110.200 ;
        RECT 165.400 105.200 165.700 195.800 ;
        RECT 167.000 172.800 167.400 173.200 ;
        RECT 167.000 155.200 167.300 172.800 ;
        RECT 167.800 166.800 168.200 167.200 ;
        RECT 167.800 166.200 168.100 166.800 ;
        RECT 167.800 165.800 168.200 166.200 ;
        RECT 167.000 154.800 167.400 155.200 ;
        RECT 167.000 129.200 167.300 154.800 ;
        RECT 167.000 128.800 167.400 129.200 ;
        RECT 166.200 124.800 166.600 125.200 ;
        RECT 165.400 104.800 165.800 105.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 162.200 71.200 162.500 84.800 ;
        RECT 165.400 77.100 165.800 77.200 ;
        RECT 164.600 76.800 165.800 77.100 ;
        RECT 164.600 73.200 164.900 76.800 ;
        RECT 164.600 72.800 165.000 73.200 ;
        RECT 162.200 70.800 162.600 71.200 ;
        RECT 161.400 64.800 161.800 65.200 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 164.600 37.800 165.000 38.200 ;
        RECT 159.800 36.800 160.200 37.200 ;
        RECT 157.400 30.800 157.800 31.200 ;
        RECT 141.400 29.800 141.800 30.200 ;
        RECT 141.400 27.200 141.700 29.800 ;
        RECT 141.400 26.800 141.800 27.200 ;
        RECT 143.000 26.800 143.400 27.200 ;
        RECT 143.000 24.200 143.300 26.800 ;
        RECT 138.200 23.800 138.600 24.200 ;
        RECT 143.000 23.800 143.400 24.200 ;
        RECT 137.400 21.800 137.800 22.200 ;
        RECT 131.800 14.800 132.200 15.200 ;
        RECT 113.400 14.100 113.800 14.200 ;
        RECT 112.600 13.800 113.800 14.100 ;
        RECT 137.400 10.200 137.700 21.800 ;
        RECT 138.200 19.200 138.500 23.800 ;
        RECT 138.200 18.800 138.600 19.200 ;
        RECT 143.800 18.800 144.200 19.200 ;
        RECT 139.800 11.800 140.200 12.200 ;
        RECT 137.400 9.800 137.800 10.200 ;
        RECT 17.400 5.800 17.800 6.200 ;
        RECT 19.800 5.800 20.200 6.200 ;
        RECT 67.800 6.100 68.200 6.200 ;
        RECT 68.600 6.100 69.000 6.200 ;
        RECT 67.800 5.800 69.000 6.100 ;
        RECT 108.600 5.800 109.000 6.200 ;
        RECT 109.400 6.100 109.800 6.200 ;
        RECT 110.200 6.100 110.600 6.200 ;
        RECT 109.400 5.800 110.600 6.100 ;
        RECT 139.800 6.100 140.100 11.800 ;
        RECT 143.800 6.200 144.100 18.800 ;
        RECT 157.400 16.200 157.700 30.800 ;
        RECT 159.800 21.200 160.100 36.800 ;
        RECT 164.600 36.200 164.900 37.800 ;
        RECT 166.200 37.200 166.500 124.800 ;
        RECT 167.000 43.200 167.300 128.800 ;
        RECT 169.400 110.200 169.700 204.800 ;
        RECT 175.000 186.800 175.400 187.200 ;
        RECT 171.000 184.800 171.400 185.200 ;
        RECT 170.200 173.800 170.600 174.200 ;
        RECT 170.200 146.200 170.500 173.800 ;
        RECT 170.200 145.800 170.600 146.200 ;
        RECT 171.000 145.200 171.300 184.800 ;
        RECT 175.000 175.100 175.300 186.800 ;
        RECT 181.400 183.200 181.700 230.800 ;
        RECT 183.000 225.200 183.300 234.800 ;
        RECT 220.600 234.100 221.000 234.200 ;
        RECT 220.600 233.800 221.700 234.100 ;
        RECT 197.400 225.800 197.800 226.200 ;
        RECT 215.800 225.800 216.200 226.200 ;
        RECT 183.000 224.800 183.400 225.200 ;
        RECT 182.200 223.800 182.600 224.200 ;
        RECT 182.200 218.200 182.500 223.800 ;
        RECT 182.200 217.800 182.600 218.200 ;
        RECT 181.400 182.800 181.800 183.200 ;
        RECT 175.800 175.100 176.200 175.200 ;
        RECT 175.000 174.800 176.200 175.100 ;
        RECT 176.600 165.800 177.000 166.200 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 176.600 165.200 176.900 165.800 ;
        RECT 175.000 165.100 175.400 165.200 ;
        RECT 175.000 164.800 176.100 165.100 ;
        RECT 176.600 164.800 177.000 165.200 ;
        RECT 172.600 160.800 173.000 161.200 ;
        RECT 171.800 156.800 172.200 157.200 ;
        RECT 171.000 144.800 171.400 145.200 ;
        RECT 171.800 115.200 172.100 156.800 ;
        RECT 171.800 114.800 172.200 115.200 ;
        RECT 170.200 110.800 170.600 111.200 ;
        RECT 168.600 109.800 169.000 110.200 ;
        RECT 169.400 109.800 169.800 110.200 ;
        RECT 167.800 77.800 168.200 78.200 ;
        RECT 167.800 55.200 168.100 77.800 ;
        RECT 168.600 68.200 168.900 109.800 ;
        RECT 169.400 75.200 169.700 109.800 ;
        RECT 169.400 74.800 169.800 75.200 ;
        RECT 169.400 73.800 169.800 74.200 ;
        RECT 169.400 73.200 169.700 73.800 ;
        RECT 169.400 72.800 169.800 73.200 ;
        RECT 168.600 67.800 169.000 68.200 ;
        RECT 170.200 66.200 170.500 110.800 ;
        RECT 172.600 96.200 172.900 160.800 ;
        RECT 175.800 126.200 176.100 164.800 ;
        RECT 175.800 125.800 176.200 126.200 ;
        RECT 179.800 123.200 180.100 165.800 ;
        RECT 181.400 128.200 181.700 182.800 ;
        RECT 182.200 178.200 182.500 217.800 ;
        RECT 183.000 184.200 183.300 224.800 ;
        RECT 190.200 217.800 190.600 218.200 ;
        RECT 185.400 214.800 185.800 215.200 ;
        RECT 184.600 186.100 185.000 186.200 ;
        RECT 185.400 186.100 185.700 214.800 ;
        RECT 190.200 206.200 190.500 217.800 ;
        RECT 190.200 205.800 190.600 206.200 ;
        RECT 186.200 196.800 186.600 197.200 ;
        RECT 186.200 188.200 186.500 196.800 ;
        RECT 187.000 190.800 187.400 191.200 ;
        RECT 186.200 187.800 186.600 188.200 ;
        RECT 184.600 185.800 185.700 186.100 ;
        RECT 183.000 183.800 183.400 184.200 ;
        RECT 184.600 184.100 185.000 184.200 ;
        RECT 185.400 184.100 185.800 184.200 ;
        RECT 184.600 183.800 185.800 184.100 ;
        RECT 182.200 177.800 182.600 178.200 ;
        RECT 181.400 127.800 181.800 128.200 ;
        RECT 179.800 122.800 180.200 123.200 ;
        RECT 175.800 115.800 176.200 116.200 ;
        RECT 172.600 95.800 173.000 96.200 ;
        RECT 175.000 93.800 175.400 94.200 ;
        RECT 175.000 89.200 175.300 93.800 ;
        RECT 175.000 88.800 175.400 89.200 ;
        RECT 171.000 87.100 171.400 87.200 ;
        RECT 171.800 87.100 172.200 87.200 ;
        RECT 171.000 86.800 172.200 87.100 ;
        RECT 175.800 81.200 176.100 115.800 ;
        RECT 178.200 96.800 178.600 97.200 ;
        RECT 178.200 84.200 178.500 96.800 ;
        RECT 178.200 83.800 178.600 84.200 ;
        RECT 175.000 80.800 175.400 81.200 ;
        RECT 175.800 80.800 176.200 81.200 ;
        RECT 173.400 66.800 173.800 67.200 ;
        RECT 173.400 66.200 173.700 66.800 ;
        RECT 175.000 66.200 175.300 80.800 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 175.000 65.800 175.400 66.200 ;
        RECT 167.800 54.800 168.200 55.200 ;
        RECT 167.000 42.800 167.400 43.200 ;
        RECT 166.200 36.800 166.600 37.200 ;
        RECT 164.600 35.800 165.000 36.200 ;
        RECT 181.400 35.200 181.700 127.800 ;
        RECT 183.000 107.200 183.300 183.800 ;
        RECT 185.400 177.800 185.800 178.200 ;
        RECT 185.400 174.200 185.700 177.800 ;
        RECT 185.400 173.800 185.800 174.200 ;
        RECT 184.600 163.800 185.000 164.200 ;
        RECT 184.600 159.200 184.900 163.800 ;
        RECT 184.600 158.800 185.000 159.200 ;
        RECT 183.800 145.800 184.200 146.200 ;
        RECT 183.000 106.800 183.400 107.200 ;
        RECT 183.800 92.200 184.100 145.800 ;
        RECT 184.600 102.200 184.900 158.800 ;
        RECT 185.400 126.200 185.700 173.800 ;
        RECT 187.000 133.200 187.300 190.800 ;
        RECT 187.800 186.800 188.200 187.200 ;
        RECT 187.800 186.200 188.100 186.800 ;
        RECT 187.800 185.800 188.200 186.200 ;
        RECT 187.800 140.200 188.100 185.800 ;
        RECT 190.200 146.200 190.500 205.800 ;
        RECT 193.400 205.100 193.800 205.200 ;
        RECT 192.600 204.800 193.800 205.100 ;
        RECT 191.000 193.100 191.400 193.200 ;
        RECT 191.000 192.800 192.100 193.100 ;
        RECT 190.200 145.800 190.600 146.200 ;
        RECT 187.800 139.800 188.200 140.200 ;
        RECT 191.800 139.200 192.100 192.800 ;
        RECT 192.600 171.200 192.900 204.800 ;
        RECT 196.600 174.800 197.000 175.200 ;
        RECT 195.800 173.800 196.200 174.200 ;
        RECT 192.600 170.800 193.000 171.200 ;
        RECT 187.800 138.800 188.200 139.200 ;
        RECT 191.800 138.800 192.200 139.200 ;
        RECT 187.800 134.200 188.100 138.800 ;
        RECT 187.800 133.800 188.200 134.200 ;
        RECT 187.000 132.800 187.400 133.200 ;
        RECT 186.200 131.800 186.600 132.200 ;
        RECT 185.400 125.800 185.800 126.200 ;
        RECT 184.600 101.800 185.000 102.200 ;
        RECT 183.800 91.800 184.200 92.200 ;
        RECT 183.800 75.800 184.200 76.200 ;
        RECT 183.800 51.200 184.100 75.800 ;
        RECT 184.600 75.200 184.900 101.800 ;
        RECT 184.600 74.800 185.000 75.200 ;
        RECT 183.800 50.800 184.200 51.200 ;
        RECT 184.600 49.200 184.900 74.800 ;
        RECT 184.600 48.800 185.000 49.200 ;
        RECT 185.400 44.200 185.700 125.800 ;
        RECT 186.200 92.200 186.500 131.800 ;
        RECT 187.000 97.200 187.300 132.800 ;
        RECT 187.000 96.800 187.400 97.200 ;
        RECT 186.200 91.800 186.600 92.200 ;
        RECT 187.800 46.200 188.100 133.800 ;
        RECT 192.600 124.200 192.900 170.800 ;
        RECT 193.400 167.800 193.800 168.200 ;
        RECT 193.400 167.200 193.700 167.800 ;
        RECT 193.400 166.800 193.800 167.200 ;
        RECT 195.800 163.200 196.100 173.800 ;
        RECT 195.800 162.800 196.200 163.200 ;
        RECT 195.000 127.800 195.400 128.200 ;
        RECT 192.600 123.800 193.000 124.200 ;
        RECT 191.800 120.800 192.200 121.200 ;
        RECT 191.000 104.800 191.400 105.200 ;
        RECT 191.000 104.200 191.300 104.800 ;
        RECT 191.000 103.800 191.400 104.200 ;
        RECT 188.600 86.100 189.000 86.200 ;
        RECT 188.600 85.800 189.700 86.100 ;
        RECT 186.200 45.800 186.600 46.200 ;
        RECT 187.800 45.800 188.200 46.200 ;
        RECT 185.400 43.800 185.800 44.200 ;
        RECT 181.400 34.800 181.800 35.200 ;
        RECT 186.200 30.200 186.500 45.800 ;
        RECT 189.400 43.200 189.700 85.800 ;
        RECT 190.200 66.100 190.600 66.200 ;
        RECT 191.000 66.100 191.400 66.200 ;
        RECT 190.200 65.800 191.400 66.100 ;
        RECT 189.400 42.800 189.800 43.200 ;
        RECT 191.800 38.200 192.100 120.800 ;
        RECT 192.600 83.800 193.000 84.200 ;
        RECT 192.600 67.200 192.900 83.800 ;
        RECT 194.200 75.800 194.600 76.200 ;
        RECT 194.200 75.200 194.500 75.800 ;
        RECT 195.000 75.200 195.300 127.800 ;
        RECT 195.800 121.200 196.100 162.800 ;
        RECT 195.800 120.800 196.200 121.200 ;
        RECT 195.800 115.800 196.200 116.200 ;
        RECT 195.800 98.200 196.100 115.800 ;
        RECT 196.600 106.200 196.900 174.800 ;
        RECT 197.400 136.200 197.700 225.800 ;
        RECT 211.800 218.800 212.200 219.200 ;
        RECT 199.800 205.800 200.200 206.200 ;
        RECT 199.800 186.200 200.100 205.800 ;
        RECT 200.600 194.800 201.000 195.200 ;
        RECT 199.800 185.800 200.200 186.200 ;
        RECT 200.600 174.200 200.900 194.800 ;
        RECT 210.200 190.800 210.600 191.200 ;
        RECT 209.400 185.800 209.800 186.200 ;
        RECT 209.400 183.200 209.700 185.800 ;
        RECT 209.400 182.800 209.800 183.200 ;
        RECT 210.200 179.200 210.500 190.800 ;
        RECT 210.200 178.800 210.600 179.200 ;
        RECT 209.400 177.100 209.800 177.200 ;
        RECT 210.200 177.100 210.600 177.200 ;
        RECT 209.400 176.800 210.600 177.100 ;
        RECT 200.600 173.800 201.000 174.200 ;
        RECT 204.600 173.800 205.000 174.200 ;
        RECT 210.200 174.100 210.600 174.200 ;
        RECT 211.000 174.100 211.400 174.200 ;
        RECT 210.200 173.800 211.400 174.100 ;
        RECT 198.200 152.100 198.600 152.200 ;
        RECT 198.200 151.800 199.300 152.100 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 199.000 126.200 199.300 151.800 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 202.200 146.200 202.500 146.800 ;
        RECT 202.200 145.800 202.600 146.200 ;
        RECT 199.000 125.800 199.400 126.200 ;
        RECT 197.400 114.800 197.800 115.200 ;
        RECT 196.600 105.800 197.000 106.200 ;
        RECT 195.800 97.800 196.200 98.200 ;
        RECT 197.400 77.200 197.700 114.800 ;
        RECT 198.200 108.800 198.600 109.200 ;
        RECT 197.400 76.800 197.800 77.200 ;
        RECT 194.200 74.800 194.600 75.200 ;
        RECT 195.000 74.800 195.400 75.200 ;
        RECT 192.600 66.800 193.000 67.200 ;
        RECT 195.000 65.800 195.400 66.200 ;
        RECT 195.000 45.200 195.300 65.800 ;
        RECT 195.000 44.800 195.400 45.200 ;
        RECT 191.800 37.800 192.200 38.200 ;
        RECT 198.200 36.200 198.500 108.800 ;
        RECT 204.600 106.200 204.900 173.800 ;
        RECT 211.000 171.800 211.400 172.200 ;
        RECT 211.000 165.200 211.300 171.800 ;
        RECT 211.000 164.800 211.400 165.200 ;
        RECT 209.400 157.800 209.800 158.200 ;
        RECT 200.600 106.100 201.000 106.200 ;
        RECT 201.400 106.100 201.800 106.200 ;
        RECT 200.600 105.800 201.800 106.100 ;
        RECT 204.600 105.800 205.000 106.200 ;
        RECT 207.800 106.100 208.200 106.200 ;
        RECT 208.600 106.100 209.000 106.200 ;
        RECT 207.800 105.800 209.000 106.100 ;
        RECT 200.600 73.800 201.000 74.200 ;
        RECT 204.600 74.100 204.900 105.800 ;
        RECT 207.800 103.800 208.200 104.200 ;
        RECT 207.800 83.200 208.100 103.800 ;
        RECT 209.400 101.200 209.700 157.800 ;
        RECT 209.400 100.800 209.800 101.200 ;
        RECT 208.600 83.800 209.000 84.200 ;
        RECT 207.800 82.800 208.200 83.200 ;
        RECT 206.200 75.100 206.600 75.200 ;
        RECT 207.000 75.100 207.400 75.200 ;
        RECT 206.200 74.800 207.400 75.100 ;
        RECT 205.400 74.100 205.800 74.200 ;
        RECT 204.600 73.800 205.800 74.100 ;
        RECT 199.000 66.100 199.400 66.200 ;
        RECT 199.800 66.100 200.200 66.200 ;
        RECT 199.000 65.800 200.200 66.100 ;
        RECT 200.600 53.200 200.900 73.800 ;
        RECT 205.400 72.800 205.800 73.200 ;
        RECT 203.800 69.800 204.200 70.200 ;
        RECT 203.800 67.200 204.100 69.800 ;
        RECT 203.800 66.800 204.200 67.200 ;
        RECT 205.400 66.200 205.700 72.800 ;
        RECT 205.400 65.800 205.800 66.200 ;
        RECT 200.600 52.800 201.000 53.200 ;
        RECT 198.200 35.800 198.600 36.200 ;
        RECT 208.600 33.200 208.900 83.800 ;
        RECT 211.000 81.200 211.300 164.800 ;
        RECT 211.800 125.200 212.100 218.800 ;
        RECT 212.600 216.800 213.000 217.200 ;
        RECT 212.600 141.200 212.900 216.800 ;
        RECT 215.800 195.200 216.100 225.800 ;
        RECT 219.800 195.800 220.200 196.200 ;
        RECT 215.800 194.800 216.200 195.200 ;
        RECT 218.200 191.800 218.600 192.200 ;
        RECT 218.200 186.200 218.500 191.800 ;
        RECT 218.200 186.100 218.600 186.200 ;
        RECT 217.400 185.800 218.600 186.100 ;
        RECT 215.800 175.100 216.200 175.200 ;
        RECT 216.600 175.100 217.000 175.200 ;
        RECT 215.800 174.800 217.000 175.100 ;
        RECT 216.600 157.800 217.000 158.200 ;
        RECT 213.400 146.100 213.800 146.200 ;
        RECT 214.200 146.100 214.600 146.200 ;
        RECT 213.400 145.800 214.600 146.100 ;
        RECT 212.600 140.800 213.000 141.200 ;
        RECT 211.800 124.800 212.200 125.200 ;
        RECT 215.000 123.800 215.400 124.200 ;
        RECT 212.600 101.800 213.000 102.200 ;
        RECT 211.000 80.800 211.400 81.200 ;
        RECT 212.600 67.200 212.900 101.800 ;
        RECT 212.600 66.800 213.000 67.200 ;
        RECT 214.200 66.800 214.600 67.200 ;
        RECT 214.200 65.200 214.500 66.800 ;
        RECT 214.200 64.800 214.600 65.200 ;
        RECT 208.600 32.800 209.000 33.200 ;
        RECT 186.200 29.800 186.600 30.200 ;
        RECT 160.600 26.100 161.000 26.200 ;
        RECT 161.400 26.100 161.800 26.200 ;
        RECT 160.600 25.800 161.800 26.100 ;
        RECT 196.600 23.800 197.000 24.200 ;
        RECT 159.800 20.800 160.200 21.200 ;
        RECT 157.400 15.800 157.800 16.200 ;
        RECT 196.600 7.200 196.900 23.800 ;
        RECT 215.000 18.200 215.300 123.800 ;
        RECT 215.800 105.800 216.200 106.200 ;
        RECT 215.800 105.200 216.100 105.800 ;
        RECT 215.800 104.800 216.200 105.200 ;
        RECT 215.800 99.800 216.200 100.200 ;
        RECT 215.000 17.800 215.400 18.200 ;
        RECT 215.800 15.200 216.100 99.800 ;
        RECT 216.600 68.200 216.900 157.800 ;
        RECT 216.600 67.800 217.000 68.200 ;
        RECT 216.600 27.200 216.900 67.800 ;
        RECT 217.400 47.200 217.700 185.800 ;
        RECT 219.800 185.200 220.100 195.800 ;
        RECT 218.200 184.800 218.600 185.200 ;
        RECT 219.800 184.800 220.200 185.200 ;
        RECT 218.200 104.200 218.500 184.800 ;
        RECT 219.800 127.100 220.100 184.800 ;
        RECT 221.400 148.200 221.700 233.800 ;
        RECT 223.800 233.800 224.200 234.200 ;
        RECT 230.200 233.800 230.600 234.200 ;
        RECT 222.200 198.800 222.600 199.200 ;
        RECT 222.200 167.200 222.500 198.800 ;
        RECT 223.000 179.800 223.400 180.200 ;
        RECT 222.200 166.800 222.600 167.200 ;
        RECT 221.400 147.800 221.800 148.200 ;
        RECT 222.200 146.200 222.500 166.800 ;
        RECT 222.200 145.800 222.600 146.200 ;
        RECT 220.600 127.100 221.000 127.200 ;
        RECT 219.800 126.800 221.000 127.100 ;
        RECT 220.600 125.200 220.900 126.800 ;
        RECT 220.600 124.800 221.000 125.200 ;
        RECT 218.200 103.800 218.600 104.200 ;
        RECT 219.800 103.800 220.200 104.200 ;
        RECT 217.400 46.800 217.800 47.200 ;
        RECT 219.800 34.200 220.100 103.800 ;
        RECT 220.600 84.200 220.900 124.800 ;
        RECT 222.200 104.200 222.500 145.800 ;
        RECT 222.200 103.800 222.600 104.200 ;
        RECT 220.600 83.800 221.000 84.200 ;
        RECT 223.000 36.200 223.300 179.800 ;
        RECT 223.800 68.200 224.100 233.800 ;
        RECT 226.200 225.800 226.600 226.200 ;
        RECT 226.200 225.200 226.500 225.800 ;
        RECT 226.200 224.800 226.600 225.200 ;
        RECT 228.600 224.800 229.000 225.200 ;
        RECT 225.400 174.800 225.800 175.200 ;
        RECT 225.400 118.200 225.700 174.800 ;
        RECT 228.600 146.100 228.900 224.800 ;
        RECT 229.400 146.100 229.800 146.200 ;
        RECT 228.600 145.800 229.800 146.100 ;
        RECT 228.600 131.800 229.000 132.200 ;
        RECT 225.400 117.800 225.800 118.200 ;
        RECT 223.800 67.800 224.200 68.200 ;
        RECT 224.600 67.800 225.000 68.200 ;
        RECT 224.600 66.200 224.900 67.800 ;
        RECT 224.600 65.800 225.000 66.200 ;
        RECT 225.400 46.200 225.700 117.800 ;
        RECT 228.600 68.200 228.900 131.800 ;
        RECT 229.400 109.200 229.700 145.800 ;
        RECT 230.200 113.200 230.500 233.800 ;
        RECT 230.200 112.800 230.600 113.200 ;
        RECT 229.400 108.800 229.800 109.200 ;
        RECT 229.400 105.100 229.800 105.200 ;
        RECT 230.200 105.100 230.600 105.200 ;
        RECT 229.400 104.800 230.600 105.100 ;
        RECT 230.200 103.800 230.600 104.200 ;
        RECT 228.600 67.800 229.000 68.200 ;
        RECT 230.200 58.200 230.500 103.800 ;
        RECT 231.000 86.200 231.300 234.800 ;
        RECT 233.400 231.800 233.800 232.200 ;
        RECT 232.600 194.800 233.000 195.200 ;
        RECT 231.800 190.800 232.200 191.200 ;
        RECT 231.800 136.200 232.100 190.800 ;
        RECT 231.800 135.800 232.200 136.200 ;
        RECT 232.600 135.100 232.900 194.800 ;
        RECT 231.800 134.800 232.900 135.100 ;
        RECT 231.800 104.200 232.100 134.800 ;
        RECT 232.600 118.800 233.000 119.200 ;
        RECT 231.800 103.800 232.200 104.200 ;
        RECT 231.000 85.800 231.400 86.200 ;
        RECT 231.000 68.100 231.400 68.200 ;
        RECT 231.000 67.800 232.100 68.100 ;
        RECT 230.200 57.800 230.600 58.200 ;
        RECT 231.800 55.200 232.100 67.800 ;
        RECT 232.600 58.200 232.900 118.800 ;
        RECT 233.400 94.200 233.700 231.800 ;
        RECT 235.800 227.800 236.200 228.200 ;
        RECT 235.000 222.800 235.400 223.200 ;
        RECT 235.000 175.200 235.300 222.800 ;
        RECT 235.000 174.800 235.400 175.200 ;
        RECT 235.000 95.200 235.300 174.800 ;
        RECT 235.800 145.200 236.100 227.800 ;
        RECT 237.400 215.800 237.800 216.200 ;
        RECT 237.400 213.200 237.700 215.800 ;
        RECT 237.400 212.800 237.800 213.200 ;
        RECT 236.600 197.800 237.000 198.200 ;
        RECT 235.800 144.800 236.200 145.200 ;
        RECT 235.000 94.800 235.400 95.200 ;
        RECT 233.400 93.800 233.800 94.200 ;
        RECT 232.600 57.800 233.000 58.200 ;
        RECT 231.800 54.800 232.200 55.200 ;
        RECT 234.200 48.800 234.600 49.200 ;
        RECT 234.200 46.200 234.500 48.800 ;
        RECT 225.400 45.800 225.800 46.200 ;
        RECT 234.200 45.800 234.600 46.200 ;
        RECT 223.000 35.800 223.400 36.200 ;
        RECT 219.800 33.800 220.200 34.200 ;
        RECT 236.600 27.200 236.900 197.800 ;
        RECT 237.400 175.800 237.800 176.200 ;
        RECT 237.400 162.200 237.700 175.800 ;
        RECT 237.400 161.800 237.800 162.200 ;
        RECT 237.400 160.800 237.800 161.200 ;
        RECT 237.400 107.200 237.700 160.800 ;
        RECT 238.200 146.200 238.500 235.800 ;
        RECT 241.400 234.800 241.800 235.200 ;
        RECT 239.000 231.800 239.400 232.200 ;
        RECT 239.000 161.200 239.300 231.800 ;
        RECT 241.400 185.200 241.700 234.800 ;
        RECT 246.200 233.800 246.600 234.200 ;
        RECT 244.600 231.800 245.000 232.200 ;
        RECT 244.600 224.200 244.900 231.800 ;
        RECT 244.600 223.800 245.000 224.200 ;
        RECT 244.600 203.200 244.900 223.800 ;
        RECT 245.400 218.800 245.800 219.200 ;
        RECT 244.600 202.800 245.000 203.200 ;
        RECT 242.200 195.800 242.600 196.200 ;
        RECT 241.400 184.800 241.800 185.200 ;
        RECT 242.200 184.100 242.500 195.800 ;
        RECT 241.400 183.800 242.500 184.100 ;
        RECT 244.600 193.800 245.000 194.200 ;
        RECT 239.800 181.800 240.200 182.200 ;
        RECT 239.000 160.800 239.400 161.200 ;
        RECT 239.000 159.800 239.400 160.200 ;
        RECT 238.200 145.800 238.600 146.200 ;
        RECT 237.400 106.800 237.800 107.200 ;
        RECT 238.200 61.200 238.500 145.800 ;
        RECT 239.000 144.200 239.300 159.800 ;
        RECT 239.000 143.800 239.400 144.200 ;
        RECT 239.000 142.800 239.400 143.200 ;
        RECT 239.000 127.200 239.300 142.800 ;
        RECT 239.000 126.800 239.400 127.200 ;
        RECT 239.000 126.200 239.300 126.800 ;
        RECT 239.000 125.800 239.400 126.200 ;
        RECT 239.800 116.200 240.100 181.800 ;
        RECT 240.600 171.800 241.000 172.200 ;
        RECT 239.800 116.100 240.200 116.200 ;
        RECT 239.000 115.800 240.200 116.100 ;
        RECT 238.200 60.800 238.600 61.200 ;
        RECT 239.000 45.200 239.300 115.800 ;
        RECT 239.800 73.800 240.200 74.200 ;
        RECT 239.000 44.800 239.400 45.200 ;
        RECT 239.800 36.200 240.100 73.800 ;
        RECT 239.800 35.800 240.200 36.200 ;
        RECT 216.600 26.800 217.000 27.200 ;
        RECT 236.600 26.800 237.000 27.200 ;
        RECT 240.600 24.200 240.900 171.800 ;
        RECT 241.400 160.200 241.700 183.800 ;
        RECT 243.800 169.800 244.200 170.200 ;
        RECT 242.200 160.800 242.600 161.200 ;
        RECT 241.400 159.800 241.800 160.200 ;
        RECT 241.400 149.800 241.800 150.200 ;
        RECT 241.400 128.200 241.700 149.800 ;
        RECT 241.400 127.800 241.800 128.200 ;
        RECT 241.400 126.800 241.800 127.200 ;
        RECT 241.400 112.200 241.700 126.800 ;
        RECT 241.400 111.800 241.800 112.200 ;
        RECT 241.400 108.800 241.800 109.200 ;
        RECT 241.400 87.200 241.700 108.800 ;
        RECT 241.400 86.800 241.800 87.200 ;
        RECT 242.200 54.200 242.500 160.800 ;
        RECT 243.000 148.800 243.400 149.200 ;
        RECT 243.000 115.200 243.300 148.800 ;
        RECT 243.000 114.800 243.400 115.200 ;
        RECT 243.800 107.200 244.100 169.800 ;
        RECT 244.600 109.200 244.900 193.800 ;
        RECT 244.600 108.800 245.000 109.200 ;
        RECT 243.800 106.800 244.200 107.200 ;
        RECT 243.000 96.100 243.400 96.200 ;
        RECT 243.000 95.800 244.100 96.100 ;
        RECT 243.800 95.200 244.100 95.800 ;
        RECT 243.000 94.800 243.400 95.200 ;
        RECT 243.800 94.800 244.200 95.200 ;
        RECT 242.200 53.800 242.600 54.200 ;
        RECT 243.000 52.200 243.300 94.800 ;
        RECT 245.400 66.200 245.700 218.800 ;
        RECT 246.200 194.200 246.500 233.800 ;
        RECT 247.000 226.100 247.400 226.200 ;
        RECT 247.800 226.100 248.200 226.200 ;
        RECT 247.000 225.800 248.200 226.100 ;
        RECT 249.400 208.800 249.800 209.200 ;
        RECT 246.200 193.800 246.600 194.200 ;
        RECT 248.600 181.800 249.000 182.200 ;
        RECT 247.800 173.800 248.200 174.200 ;
        RECT 247.000 126.800 247.400 127.200 ;
        RECT 246.200 119.800 246.600 120.200 ;
        RECT 245.400 65.800 245.800 66.200 ;
        RECT 243.000 51.800 243.400 52.200 ;
        RECT 240.600 23.800 241.000 24.200 ;
        RECT 215.800 14.800 216.200 15.200 ;
        RECT 246.200 9.200 246.500 119.800 ;
        RECT 247.000 87.200 247.300 126.800 ;
        RECT 247.800 106.200 248.100 173.800 ;
        RECT 248.600 155.200 248.900 181.800 ;
        RECT 248.600 154.800 249.000 155.200 ;
        RECT 248.600 125.200 248.900 154.800 ;
        RECT 248.600 124.800 249.000 125.200 ;
        RECT 248.600 123.800 249.000 124.200 ;
        RECT 247.800 105.800 248.200 106.200 ;
        RECT 247.000 86.800 247.400 87.200 ;
        RECT 246.200 8.800 246.600 9.200 ;
        RECT 247.000 7.200 247.300 86.800 ;
        RECT 248.600 29.200 248.900 123.800 ;
        RECT 249.400 110.200 249.700 208.800 ;
        RECT 251.800 196.800 252.200 197.200 ;
        RECT 251.000 175.800 251.400 176.200 ;
        RECT 250.200 149.800 250.600 150.200 ;
        RECT 249.400 109.800 249.800 110.200 ;
        RECT 250.200 107.100 250.500 149.800 ;
        RECT 249.400 106.800 250.500 107.100 ;
        RECT 249.400 76.200 249.700 106.800 ;
        RECT 251.000 106.100 251.300 175.800 ;
        RECT 250.200 105.800 251.300 106.100 ;
        RECT 249.400 75.800 249.800 76.200 ;
        RECT 250.200 36.200 250.500 105.800 ;
        RECT 251.000 87.800 251.400 88.200 ;
        RECT 251.000 69.200 251.300 87.800 ;
        RECT 251.000 68.800 251.400 69.200 ;
        RECT 250.200 35.800 250.600 36.200 ;
        RECT 248.600 28.800 249.000 29.200 ;
        RECT 251.800 25.200 252.100 196.800 ;
        RECT 251.800 24.800 252.200 25.200 ;
        RECT 196.600 6.800 197.000 7.200 ;
        RECT 247.000 6.800 247.400 7.200 ;
        RECT 140.600 6.100 141.000 6.200 ;
        RECT 139.800 5.800 141.000 6.100 ;
        RECT 143.800 5.800 144.200 6.200 ;
      LAYER via4 ;
        RECT 236.600 234.800 237.000 235.200 ;
        RECT 5.400 233.800 5.800 234.200 ;
        RECT 39.800 225.800 40.200 226.200 ;
        RECT 12.600 74.800 13.000 75.200 ;
        RECT 33.400 75.800 33.800 76.200 ;
        RECT 31.800 73.800 32.200 74.200 ;
        RECT 34.200 66.800 34.600 67.200 ;
        RECT 28.600 65.800 29.000 66.200 ;
        RECT 58.200 185.800 58.600 186.200 ;
        RECT 49.400 66.800 49.800 67.200 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 63.800 194.800 64.200 195.200 ;
        RECT 56.600 63.800 57.000 64.200 ;
        RECT 60.600 63.800 61.000 64.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 79.000 114.800 79.400 115.200 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 82.200 65.800 82.600 66.200 ;
        RECT 91.800 85.800 92.200 86.200 ;
        RECT 155.000 226.800 155.400 227.200 ;
        RECT 113.400 205.800 113.800 206.200 ;
        RECT 110.200 104.800 110.600 105.200 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 135.000 103.800 135.400 104.200 ;
        RECT 145.400 192.800 145.800 193.200 ;
        RECT 150.200 186.800 150.600 187.200 ;
        RECT 159.000 184.800 159.400 185.200 ;
        RECT 160.600 86.800 161.000 87.200 ;
        RECT 171.800 86.800 172.200 87.200 ;
        RECT 201.400 105.800 201.800 106.200 ;
        RECT 208.600 105.800 209.000 106.200 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 161.400 25.800 161.800 26.200 ;
        RECT 247.800 225.800 248.200 226.200 ;
      LAYER metal5 ;
        RECT 236.600 234.800 237.000 235.200 ;
        RECT 236.600 234.200 236.900 234.800 ;
        RECT 5.400 234.100 5.800 234.200 ;
        RECT 122.200 234.100 122.600 234.200 ;
        RECT 5.400 233.800 122.600 234.100 ;
        RECT 236.500 233.700 237.000 234.200 ;
        RECT 135.800 227.100 136.200 227.200 ;
        RECT 155.000 227.100 155.400 227.200 ;
        RECT 135.800 226.800 155.400 227.100 ;
        RECT 39.800 226.100 40.200 226.200 ;
        RECT 59.000 226.100 59.400 226.200 ;
        RECT 39.800 225.800 59.400 226.100 ;
        RECT 247.800 225.800 248.200 226.200 ;
        RECT 247.800 225.200 248.100 225.800 ;
        RECT 43.800 225.100 44.200 225.200 ;
        RECT 124.600 225.100 125.000 225.200 ;
        RECT 43.800 224.800 125.000 225.100 ;
        RECT 144.600 225.100 145.000 225.200 ;
        RECT 226.200 225.100 226.600 225.200 ;
        RECT 144.600 224.800 226.600 225.100 ;
        RECT 247.700 224.700 248.200 225.200 ;
        RECT 75.800 224.100 76.200 224.200 ;
        RECT 115.000 224.100 115.400 224.200 ;
        RECT 75.800 223.800 115.400 224.100 ;
        RECT 59.800 213.100 60.200 213.200 ;
        RECT 131.000 213.100 131.400 213.200 ;
        RECT 237.400 213.100 237.800 213.200 ;
        RECT 59.800 212.800 237.800 213.100 ;
        RECT 113.400 206.100 113.800 206.200 ;
        RECT 190.200 206.100 190.600 206.200 ;
        RECT 113.400 205.800 190.600 206.100 ;
        RECT 85.400 202.100 85.800 202.200 ;
        RECT 111.800 202.100 112.200 202.200 ;
        RECT 85.400 201.800 112.200 202.100 ;
        RECT 82.200 196.100 82.600 196.200 ;
        RECT 95.000 196.100 95.400 196.200 ;
        RECT 144.600 196.100 145.000 196.200 ;
        RECT 82.200 195.800 145.000 196.100 ;
        RECT 63.800 195.100 64.200 195.200 ;
        RECT 70.200 195.100 70.600 195.200 ;
        RECT 63.800 194.800 70.600 195.100 ;
        RECT 51.800 194.100 52.200 194.200 ;
        RECT 130.200 194.100 130.600 194.200 ;
        RECT 51.800 193.800 130.600 194.100 ;
        RECT 145.400 193.100 145.800 193.200 ;
        RECT 191.000 193.100 191.400 193.200 ;
        RECT 145.400 192.800 191.400 193.100 ;
        RECT 74.200 187.100 74.600 187.200 ;
        RECT 150.200 187.100 150.600 187.200 ;
        RECT 187.800 187.100 188.200 187.200 ;
        RECT 74.200 186.800 188.200 187.100 ;
        RECT 58.200 186.100 58.600 186.200 ;
        RECT 134.200 186.100 134.600 186.200 ;
        RECT 58.200 185.800 134.600 186.100 ;
        RECT 159.000 185.100 159.400 185.200 ;
        RECT 219.800 185.100 220.200 185.200 ;
        RECT 159.000 184.800 220.200 185.100 ;
        RECT 154.200 184.100 154.600 184.200 ;
        RECT 184.600 184.100 185.000 184.200 ;
        RECT 154.200 183.800 185.000 184.100 ;
        RECT 117.400 183.100 117.800 183.200 ;
        RECT 209.400 183.100 209.800 183.200 ;
        RECT 117.400 182.800 209.800 183.100 ;
        RECT 60.600 177.100 61.000 177.200 ;
        RECT 150.200 177.100 150.600 177.200 ;
        RECT 209.400 177.100 209.800 177.200 ;
        RECT 60.600 176.800 209.800 177.100 ;
        RECT 133.400 175.100 133.800 175.200 ;
        RECT 215.800 175.100 216.200 175.200 ;
        RECT 133.400 174.800 216.200 175.100 ;
        RECT 185.400 174.100 185.800 174.200 ;
        RECT 210.200 174.100 210.600 174.200 ;
        RECT 185.400 173.800 210.600 174.100 ;
        RECT 19.000 166.800 19.400 167.200 ;
        RECT 159.800 167.100 160.200 167.200 ;
        RECT 193.400 167.100 193.800 167.200 ;
        RECT 159.800 166.800 193.800 167.100 ;
        RECT 19.000 166.100 19.300 166.800 ;
        RECT 107.800 166.100 108.200 166.200 ;
        RECT 19.000 165.800 108.200 166.100 ;
        RECT 167.800 166.100 168.200 166.200 ;
        RECT 176.600 166.100 177.000 166.200 ;
        RECT 167.800 165.800 177.000 166.100 ;
        RECT 123.800 165.100 124.200 165.200 ;
        RECT 175.000 165.100 175.400 165.200 ;
        RECT 123.800 164.800 175.400 165.100 ;
        RECT 237.400 161.100 237.800 161.200 ;
        RECT 239.000 161.100 239.400 161.200 ;
        RECT 237.400 160.800 239.400 161.100 ;
        RECT 239.000 160.100 239.400 160.200 ;
        RECT 241.400 160.100 241.800 160.200 ;
        RECT 239.000 159.800 241.800 160.100 ;
        RECT 47.800 145.800 48.200 146.200 ;
        RECT 202.200 146.100 202.600 146.200 ;
        RECT 213.400 146.100 213.800 146.200 ;
        RECT 202.200 145.800 213.800 146.100 ;
        RECT 37.400 145.100 37.800 145.200 ;
        RECT 47.800 145.100 48.100 145.800 ;
        RECT 37.400 144.800 48.100 145.100 ;
        RECT 187.800 139.100 188.200 139.200 ;
        RECT 191.800 139.100 192.200 139.200 ;
        RECT 187.800 138.800 192.200 139.100 ;
        RECT 236.500 127.100 237.000 127.200 ;
        RECT 241.400 127.100 241.800 127.200 ;
        RECT 236.500 126.800 241.800 127.100 ;
        RECT 236.500 126.700 237.000 126.800 ;
        RECT 247.700 124.100 248.200 124.200 ;
        RECT 248.600 124.100 249.000 124.200 ;
        RECT 247.700 123.800 249.000 124.100 ;
        RECT 247.700 123.700 248.200 123.800 ;
        RECT 79.000 115.100 79.400 115.200 ;
        RECT 96.600 115.100 97.000 115.200 ;
        RECT 79.000 114.800 97.000 115.100 ;
        RECT 94.200 108.100 94.600 108.200 ;
        RECT 143.800 108.100 144.200 108.200 ;
        RECT 94.200 107.800 144.200 108.100 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 119.000 106.100 119.400 106.200 ;
        RECT 68.600 105.800 119.400 106.100 ;
        RECT 131.000 105.800 131.400 106.200 ;
        RECT 131.800 106.100 132.200 106.200 ;
        RECT 201.400 106.100 201.800 106.200 ;
        RECT 204.600 106.100 205.000 106.200 ;
        RECT 131.800 105.800 205.000 106.100 ;
        RECT 208.600 106.100 209.000 106.200 ;
        RECT 215.800 106.100 216.200 106.200 ;
        RECT 208.600 105.800 216.200 106.100 ;
        RECT 92.600 105.100 93.000 105.200 ;
        RECT 110.200 105.100 110.600 105.200 ;
        RECT 131.000 105.100 131.300 105.800 ;
        RECT 229.400 105.100 229.800 105.200 ;
        RECT 92.600 104.800 131.300 105.100 ;
        RECT 191.000 104.800 229.800 105.100 ;
        RECT 191.000 104.200 191.300 104.800 ;
        RECT 121.400 104.100 121.800 104.200 ;
        RECT 135.000 104.100 135.400 104.200 ;
        RECT 121.400 103.800 135.400 104.100 ;
        RECT 191.000 103.800 191.400 104.200 ;
        RECT 114.200 95.100 114.600 95.200 ;
        RECT 243.800 95.100 244.200 95.200 ;
        RECT 114.200 94.800 244.200 95.100 ;
        RECT 67.800 94.100 68.200 94.200 ;
        RECT 135.800 94.100 136.200 94.200 ;
        RECT 67.800 93.800 136.200 94.100 ;
        RECT 64.600 87.100 65.000 87.200 ;
        RECT 129.400 87.100 129.800 87.200 ;
        RECT 64.600 86.800 129.800 87.100 ;
        RECT 160.600 87.100 161.000 87.200 ;
        RECT 171.800 87.100 172.200 87.200 ;
        RECT 160.600 86.800 172.200 87.100 ;
        RECT 91.800 86.100 92.200 86.200 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 91.800 85.800 125.800 86.100 ;
        RECT 111.800 85.100 112.200 85.200 ;
        RECT 149.400 85.100 149.800 85.200 ;
        RECT 111.800 84.800 149.800 85.100 ;
        RECT 33.400 84.100 33.800 84.200 ;
        RECT 139.000 84.100 139.400 84.200 ;
        RECT 33.400 83.800 139.400 84.100 ;
        RECT 15.800 78.100 16.200 78.200 ;
        RECT 122.200 78.100 122.600 78.200 ;
        RECT 15.800 77.800 122.600 78.100 ;
        RECT 33.400 76.100 33.800 76.200 ;
        RECT 111.000 76.100 111.400 76.200 ;
        RECT 33.400 75.800 111.400 76.100 ;
        RECT 12.600 75.100 13.000 75.200 ;
        RECT 131.800 75.100 132.200 75.200 ;
        RECT 12.600 74.800 132.200 75.100 ;
        RECT 160.600 74.800 161.000 75.200 ;
        RECT 194.200 75.100 194.600 75.200 ;
        RECT 206.200 75.100 206.600 75.200 ;
        RECT 194.200 74.800 206.600 75.100 ;
        RECT 31.800 74.100 32.200 74.200 ;
        RECT 105.400 74.100 105.800 74.200 ;
        RECT 31.800 73.800 105.800 74.100 ;
        RECT 160.600 74.100 160.900 74.800 ;
        RECT 169.400 74.100 169.800 74.200 ;
        RECT 160.600 73.800 169.800 74.100 ;
        RECT 75.000 73.100 75.400 73.200 ;
        RECT 100.600 73.100 101.000 73.200 ;
        RECT 123.800 73.100 124.200 73.200 ;
        RECT 164.600 73.100 165.000 73.200 ;
        RECT 205.400 73.100 205.800 73.200 ;
        RECT 75.000 72.800 205.800 73.100 ;
        RECT 115.800 69.800 116.200 70.200 ;
        RECT 35.000 69.100 35.400 69.200 ;
        RECT 115.800 69.100 116.100 69.800 ;
        RECT 35.000 68.800 116.100 69.100 ;
        RECT 53.400 68.100 53.800 68.200 ;
        RECT 83.000 68.100 83.400 68.200 ;
        RECT 53.400 67.800 84.100 68.100 ;
        RECT 34.200 67.100 34.600 67.200 ;
        RECT 40.600 67.100 41.000 67.200 ;
        RECT 34.200 66.800 41.000 67.100 ;
        RECT 49.400 67.100 49.800 67.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 49.400 66.800 65.000 67.100 ;
        RECT 173.400 67.100 173.800 67.200 ;
        RECT 203.800 67.100 204.200 67.200 ;
        RECT 173.400 66.800 204.200 67.100 ;
        RECT 28.600 66.100 29.000 66.200 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 28.600 65.800 37.800 66.100 ;
        RECT 46.200 66.100 46.600 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 46.200 65.800 77.000 66.100 ;
        RECT 82.200 66.100 82.600 66.200 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 82.200 65.800 110.600 66.100 ;
        RECT 137.400 66.100 137.800 66.200 ;
        RECT 190.200 66.100 190.600 66.200 ;
        RECT 137.400 65.800 190.600 66.100 ;
        RECT 199.800 66.100 200.200 66.200 ;
        RECT 224.600 66.100 225.000 66.200 ;
        RECT 199.800 65.800 225.000 66.100 ;
        RECT 4.600 65.100 5.000 65.200 ;
        RECT 114.200 65.100 114.600 65.200 ;
        RECT 4.600 64.800 114.600 65.100 ;
        RECT 56.600 64.100 57.000 64.200 ;
        RECT 60.600 64.100 61.000 64.200 ;
        RECT 56.600 63.800 61.000 64.100 ;
        RECT 59.000 58.100 59.400 58.200 ;
        RECT 114.200 58.100 114.600 58.200 ;
        RECT 59.000 57.800 114.600 58.100 ;
        RECT 45.400 56.100 45.800 56.200 ;
        RECT 119.800 56.100 120.200 56.200 ;
        RECT 45.400 55.800 120.200 56.100 ;
        RECT 115.000 37.100 115.400 37.200 ;
        RECT 159.800 37.100 160.200 37.200 ;
        RECT 115.000 36.800 160.200 37.100 ;
        RECT 69.400 35.800 69.800 36.200 ;
        RECT 69.400 35.100 69.700 35.800 ;
        RECT 114.200 35.100 114.600 35.200 ;
        RECT 69.400 34.800 114.600 35.100 ;
        RECT 80.600 26.100 81.000 26.200 ;
        RECT 161.400 26.100 161.800 26.200 ;
        RECT 80.600 25.800 161.800 26.100 ;
        RECT 59.800 24.100 60.200 24.200 ;
        RECT 138.200 24.100 138.600 24.200 ;
        RECT 59.800 23.800 138.600 24.100 ;
        RECT 103.000 16.100 103.400 16.200 ;
        RECT 157.400 16.100 157.800 16.200 ;
        RECT 103.000 15.800 157.800 16.100 ;
        RECT 67.800 6.100 68.200 6.200 ;
        RECT 109.400 6.100 109.800 6.200 ;
        RECT 67.800 5.800 109.800 6.100 ;
      LAYER metal6 ;
        RECT 236.500 126.700 237.000 234.200 ;
        RECT 247.700 123.700 248.200 225.200 ;
  END
END ram32_sram
END LIBRARY

